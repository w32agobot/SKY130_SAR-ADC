* SPICE3 file created from extract2.ext - technology: sky130A

C0 extract_0/dummy_top extract_0/top_16 2.87fF
C1 extract_0/dummy_bot extract_0/bot_4 6.96fF
C2 extract_0/bot_2 extract_0/dummy_bot 6.95fF
C3 extract_0/top_4 extract_0/bot_4 4.72fF
C4 extract_0/dummy_top extract_0/dummy_bot 38.44fF
C5 extract_0/dummy_bot extract_0/bot_1 6.95fF
C6 extract_0/dummy_bot extract_0/bot_8 6.95fF
C7 extract_0/dummy_top extract_0/top_4 2.49fF
C8 extract_0/bot_16 extract_0/top_16 4.42fF
C9 extract_0/top_2 extract_0/bot_2 4.68fF
C10 extract_0/dummy_top extract_0/top_8 2.59fF
C11 extract_0/top_2 extract_0/dummy_top 2.44fF
C12 extract_0/top_8 extract_0/bot_8 4.83fF
C13 extract_0/bot_16 extract_0/dummy_bot 6.10fF
C14 extract_0/top_1 extract_0/dummy_top 2.39fF
C15 extract_0/top_1 extract_0/bot_1 4.66fF
C16 extract_0/dummy_top VSUBS 7.32fF
C17 extract_0/bot_1 VSUBS 2.65fF
C18 extract_0/bot_2 VSUBS 2.64fF
C19 extract_0/bot_4 VSUBS 2.64fF
C20 extract_0/bot_8 VSUBS 2.64fF
C21 extract_0/bot_16 VSUBS 2.01fF
C22 extract_0/dummy_bot VSUBS 36.54fF
