magic
tech sky130A
timestamp 1659968763
<< metal2 >>
rect 44 1674 414 1719
rect 44 1646 89 1674
rect 117 1646 175 1674
rect 203 1646 261 1674
rect 289 1646 347 1674
rect 375 1646 414 1674
rect 44 1588 414 1646
rect 44 1560 89 1588
rect 117 1560 175 1588
rect 203 1560 261 1588
rect 289 1560 347 1588
rect 375 1560 414 1588
rect 44 1553 414 1560
rect 442 1674 812 1719
rect 442 1646 487 1674
rect 515 1646 573 1674
rect 601 1646 659 1674
rect 687 1646 745 1674
rect 773 1646 812 1674
rect 442 1588 812 1646
rect 442 1560 487 1588
rect 515 1560 573 1588
rect 601 1560 659 1588
rect 687 1560 745 1588
rect 773 1560 812 1588
rect 442 1553 812 1560
rect 840 1674 1210 1719
rect 840 1646 885 1674
rect 913 1646 971 1674
rect 999 1646 1057 1674
rect 1085 1646 1143 1674
rect 1171 1646 1210 1674
rect 840 1588 1210 1646
rect 840 1560 885 1588
rect 913 1560 971 1588
rect 999 1560 1057 1588
rect 1085 1560 1143 1588
rect 1171 1560 1210 1588
rect 840 1553 1210 1560
rect 1238 1674 1608 1719
rect 1238 1646 1283 1674
rect 1311 1646 1369 1674
rect 1397 1646 1455 1674
rect 1483 1646 1541 1674
rect 1569 1646 1608 1674
rect 1238 1588 1608 1646
rect 1238 1560 1283 1588
rect 1311 1560 1369 1588
rect 1397 1560 1455 1588
rect 1483 1560 1541 1588
rect 1569 1560 1608 1588
rect 1238 1553 1608 1560
rect 1636 1674 2006 1719
rect 1636 1646 1681 1674
rect 1709 1646 1767 1674
rect 1795 1646 1853 1674
rect 1881 1646 1939 1674
rect 1967 1646 2006 1674
rect 1636 1588 2006 1646
rect 1636 1560 1681 1588
rect 1709 1560 1767 1588
rect 1795 1560 1853 1588
rect 1881 1560 1939 1588
rect 1967 1560 2006 1588
rect 1636 1553 2006 1560
rect 2034 1674 2404 1719
rect 2034 1646 2079 1674
rect 2107 1646 2165 1674
rect 2193 1646 2251 1674
rect 2279 1646 2337 1674
rect 2365 1646 2404 1674
rect 2034 1588 2404 1646
rect 2034 1560 2079 1588
rect 2107 1560 2165 1588
rect 2193 1560 2251 1588
rect 2279 1560 2337 1588
rect 2365 1560 2404 1588
rect 2034 1553 2404 1560
rect 2432 1674 2802 1719
rect 2432 1646 2477 1674
rect 2505 1646 2563 1674
rect 2591 1646 2649 1674
rect 2677 1646 2735 1674
rect 2763 1646 2802 1674
rect 2432 1588 2802 1646
rect 2432 1560 2477 1588
rect 2505 1560 2563 1588
rect 2591 1560 2649 1588
rect 2677 1560 2735 1588
rect 2763 1560 2802 1588
rect 2432 1553 2802 1560
rect 2830 1674 3200 1719
rect 2830 1646 2875 1674
rect 2903 1646 2961 1674
rect 2989 1646 3047 1674
rect 3075 1646 3133 1674
rect 3161 1646 3200 1674
rect 2830 1588 3200 1646
rect 2830 1560 2875 1588
rect 2903 1560 2961 1588
rect 2989 1560 3047 1588
rect 3075 1560 3133 1588
rect 3161 1560 3200 1588
rect 2830 1553 3200 1560
rect 3228 1674 3598 1719
rect 3228 1646 3273 1674
rect 3301 1646 3359 1674
rect 3387 1646 3445 1674
rect 3473 1646 3531 1674
rect 3559 1646 3598 1674
rect 3228 1588 3598 1646
rect 3228 1560 3273 1588
rect 3301 1560 3359 1588
rect 3387 1560 3445 1588
rect 3473 1560 3531 1588
rect 3559 1560 3598 1588
rect 3228 1553 3598 1560
rect 3626 1674 3996 1719
rect 3626 1646 3671 1674
rect 3699 1646 3757 1674
rect 3785 1646 3843 1674
rect 3871 1646 3929 1674
rect 3957 1646 3996 1674
rect 3626 1588 3996 1646
rect 3626 1560 3671 1588
rect 3699 1560 3757 1588
rect 3785 1560 3843 1588
rect 3871 1560 3929 1588
rect 3957 1560 3996 1588
rect 3626 1553 3996 1560
rect 4024 1674 4394 1719
rect 4024 1646 4069 1674
rect 4097 1646 4155 1674
rect 4183 1646 4241 1674
rect 4269 1646 4327 1674
rect 4355 1646 4394 1674
rect 4024 1588 4394 1646
rect 4024 1560 4069 1588
rect 4097 1560 4155 1588
rect 4183 1560 4241 1588
rect 4269 1560 4327 1588
rect 4355 1560 4394 1588
rect 4024 1553 4394 1560
rect 4422 1674 4792 1719
rect 4422 1646 4467 1674
rect 4495 1646 4553 1674
rect 4581 1646 4639 1674
rect 4667 1646 4725 1674
rect 4753 1646 4792 1674
rect 4422 1588 4792 1646
rect 4422 1560 4467 1588
rect 4495 1560 4553 1588
rect 4581 1560 4639 1588
rect 4667 1560 4725 1588
rect 4753 1560 4792 1588
rect 4422 1553 4792 1560
rect 4820 1674 5190 1719
rect 4820 1646 4865 1674
rect 4893 1646 4951 1674
rect 4979 1646 5037 1674
rect 5065 1646 5123 1674
rect 5151 1646 5190 1674
rect 4820 1588 5190 1646
rect 4820 1560 4865 1588
rect 4893 1560 4951 1588
rect 4979 1560 5037 1588
rect 5065 1560 5123 1588
rect 5151 1560 5190 1588
rect 4820 1553 5190 1560
rect 5218 1674 5588 1719
rect 5218 1646 5263 1674
rect 5291 1646 5349 1674
rect 5377 1646 5435 1674
rect 5463 1646 5521 1674
rect 5549 1646 5588 1674
rect 5218 1588 5588 1646
rect 5218 1560 5263 1588
rect 5291 1560 5349 1588
rect 5377 1560 5435 1588
rect 5463 1560 5521 1588
rect 5549 1560 5588 1588
rect 5218 1553 5588 1560
rect 5616 1674 5986 1719
rect 5616 1646 5661 1674
rect 5689 1646 5747 1674
rect 5775 1646 5833 1674
rect 5861 1646 5919 1674
rect 5947 1646 5986 1674
rect 5616 1588 5986 1646
rect 5616 1560 5661 1588
rect 5689 1560 5747 1588
rect 5775 1560 5833 1588
rect 5861 1560 5919 1588
rect 5947 1560 5986 1588
rect 5616 1553 5986 1560
rect 6014 1674 6384 1719
rect 6014 1646 6059 1674
rect 6087 1646 6145 1674
rect 6173 1646 6231 1674
rect 6259 1646 6317 1674
rect 6345 1646 6384 1674
rect 6014 1588 6384 1646
rect 6014 1560 6059 1588
rect 6087 1560 6145 1588
rect 6173 1560 6231 1588
rect 6259 1560 6317 1588
rect 6345 1560 6384 1588
rect 6014 1553 6384 1560
rect 6412 1674 6782 1719
rect 6412 1646 6457 1674
rect 6485 1646 6543 1674
rect 6571 1646 6629 1674
rect 6657 1646 6715 1674
rect 6743 1646 6782 1674
rect 6412 1588 6782 1646
rect 6412 1560 6457 1588
rect 6485 1560 6543 1588
rect 6571 1560 6629 1588
rect 6657 1560 6715 1588
rect 6743 1560 6782 1588
rect 6412 1553 6782 1560
rect 6810 1674 7180 1719
rect 6810 1646 6855 1674
rect 6883 1646 6941 1674
rect 6969 1646 7027 1674
rect 7055 1646 7113 1674
rect 7141 1646 7180 1674
rect 6810 1588 7180 1646
rect 6810 1560 6855 1588
rect 6883 1560 6941 1588
rect 6969 1560 7027 1588
rect 7055 1560 7113 1588
rect 7141 1560 7180 1588
rect 6810 1553 7180 1560
rect 7208 1674 7578 1719
rect 7208 1646 7253 1674
rect 7281 1646 7339 1674
rect 7367 1646 7425 1674
rect 7453 1646 7511 1674
rect 7539 1646 7578 1674
rect 7208 1588 7578 1646
rect 7208 1560 7253 1588
rect 7281 1560 7339 1588
rect 7367 1560 7425 1588
rect 7453 1560 7511 1588
rect 7539 1560 7578 1588
rect 7208 1553 7578 1560
rect 7606 1674 7976 1719
rect 7606 1646 7651 1674
rect 7679 1646 7737 1674
rect 7765 1646 7823 1674
rect 7851 1646 7909 1674
rect 7937 1646 7976 1674
rect 7606 1588 7976 1646
rect 7606 1560 7651 1588
rect 7679 1560 7737 1588
rect 7765 1560 7823 1588
rect 7851 1560 7909 1588
rect 7937 1560 7976 1588
rect 7606 1553 7976 1560
rect 8004 1674 8374 1719
rect 8004 1646 8049 1674
rect 8077 1646 8135 1674
rect 8163 1646 8221 1674
rect 8249 1646 8307 1674
rect 8335 1646 8374 1674
rect 8004 1588 8374 1646
rect 8004 1560 8049 1588
rect 8077 1560 8135 1588
rect 8163 1560 8221 1588
rect 8249 1560 8307 1588
rect 8335 1560 8374 1588
rect 8004 1553 8374 1560
rect 8402 1674 8772 1719
rect 8402 1646 8447 1674
rect 8475 1646 8533 1674
rect 8561 1646 8619 1674
rect 8647 1646 8705 1674
rect 8733 1646 8772 1674
rect 8402 1588 8772 1646
rect 8402 1560 8447 1588
rect 8475 1560 8533 1588
rect 8561 1560 8619 1588
rect 8647 1560 8705 1588
rect 8733 1560 8772 1588
rect 8402 1553 8772 1560
rect 8800 1674 9170 1719
rect 8800 1646 8845 1674
rect 8873 1646 8931 1674
rect 8959 1646 9017 1674
rect 9045 1646 9103 1674
rect 9131 1646 9170 1674
rect 8800 1588 9170 1646
rect 8800 1560 8845 1588
rect 8873 1560 8931 1588
rect 8959 1560 9017 1588
rect 9045 1560 9103 1588
rect 9131 1560 9170 1588
rect 8800 1553 9170 1560
rect 9198 1674 9568 1719
rect 9198 1646 9243 1674
rect 9271 1646 9329 1674
rect 9357 1646 9415 1674
rect 9443 1646 9501 1674
rect 9529 1646 9568 1674
rect 9198 1588 9568 1646
rect 9198 1560 9243 1588
rect 9271 1560 9329 1588
rect 9357 1560 9415 1588
rect 9443 1560 9501 1588
rect 9529 1560 9568 1588
rect 9198 1553 9568 1560
rect 9596 1674 9966 1719
rect 9596 1646 9641 1674
rect 9669 1646 9727 1674
rect 9755 1646 9813 1674
rect 9841 1646 9899 1674
rect 9927 1646 9966 1674
rect 9596 1588 9966 1646
rect 9596 1560 9641 1588
rect 9669 1560 9727 1588
rect 9755 1560 9813 1588
rect 9841 1560 9899 1588
rect 9927 1560 9966 1588
rect 9596 1553 9966 1560
rect 44 1533 9966 1553
rect 44 1502 414 1533
rect 44 1474 89 1502
rect 117 1474 175 1502
rect 203 1474 261 1502
rect 289 1474 347 1502
rect 375 1474 414 1502
rect 44 1416 414 1474
rect 44 1388 89 1416
rect 117 1388 175 1416
rect 203 1388 261 1416
rect 289 1388 347 1416
rect 375 1388 414 1416
rect 44 1349 414 1388
rect 442 1502 812 1533
rect 442 1474 487 1502
rect 515 1474 573 1502
rect 601 1474 659 1502
rect 687 1474 745 1502
rect 773 1474 812 1502
rect 442 1416 812 1474
rect 442 1388 487 1416
rect 515 1388 573 1416
rect 601 1388 659 1416
rect 687 1388 745 1416
rect 773 1388 812 1416
rect 442 1349 812 1388
rect 840 1502 1210 1533
rect 840 1474 885 1502
rect 913 1474 971 1502
rect 999 1474 1057 1502
rect 1085 1474 1143 1502
rect 1171 1474 1210 1502
rect 840 1416 1210 1474
rect 840 1388 885 1416
rect 913 1388 971 1416
rect 999 1388 1057 1416
rect 1085 1388 1143 1416
rect 1171 1388 1210 1416
rect 840 1349 1210 1388
rect 1238 1502 1608 1533
rect 1238 1474 1283 1502
rect 1311 1474 1369 1502
rect 1397 1474 1455 1502
rect 1483 1474 1541 1502
rect 1569 1474 1608 1502
rect 1238 1416 1608 1474
rect 1238 1388 1283 1416
rect 1311 1388 1369 1416
rect 1397 1388 1455 1416
rect 1483 1388 1541 1416
rect 1569 1388 1608 1416
rect 1238 1349 1608 1388
rect 1636 1502 2006 1533
rect 1636 1474 1681 1502
rect 1709 1474 1767 1502
rect 1795 1474 1853 1502
rect 1881 1474 1939 1502
rect 1967 1474 2006 1502
rect 1636 1416 2006 1474
rect 1636 1388 1681 1416
rect 1709 1388 1767 1416
rect 1795 1388 1853 1416
rect 1881 1388 1939 1416
rect 1967 1388 2006 1416
rect 1636 1349 2006 1388
rect 2034 1502 2404 1533
rect 2034 1474 2079 1502
rect 2107 1474 2165 1502
rect 2193 1474 2251 1502
rect 2279 1474 2337 1502
rect 2365 1474 2404 1502
rect 2034 1416 2404 1474
rect 2034 1388 2079 1416
rect 2107 1388 2165 1416
rect 2193 1388 2251 1416
rect 2279 1388 2337 1416
rect 2365 1388 2404 1416
rect 2034 1349 2404 1388
rect 2432 1502 2802 1533
rect 2432 1474 2477 1502
rect 2505 1474 2563 1502
rect 2591 1474 2649 1502
rect 2677 1474 2735 1502
rect 2763 1474 2802 1502
rect 2432 1416 2802 1474
rect 2432 1388 2477 1416
rect 2505 1388 2563 1416
rect 2591 1388 2649 1416
rect 2677 1388 2735 1416
rect 2763 1388 2802 1416
rect 2432 1349 2802 1388
rect 2830 1502 3200 1533
rect 2830 1474 2875 1502
rect 2903 1474 2961 1502
rect 2989 1474 3047 1502
rect 3075 1474 3133 1502
rect 3161 1474 3200 1502
rect 2830 1416 3200 1474
rect 2830 1388 2875 1416
rect 2903 1388 2961 1416
rect 2989 1388 3047 1416
rect 3075 1388 3133 1416
rect 3161 1388 3200 1416
rect 2830 1349 3200 1388
rect 3228 1502 3598 1533
rect 3228 1474 3273 1502
rect 3301 1474 3359 1502
rect 3387 1474 3445 1502
rect 3473 1474 3531 1502
rect 3559 1474 3598 1502
rect 3228 1416 3598 1474
rect 3228 1388 3273 1416
rect 3301 1388 3359 1416
rect 3387 1388 3445 1416
rect 3473 1388 3531 1416
rect 3559 1388 3598 1416
rect 3228 1349 3598 1388
rect 3626 1502 3996 1533
rect 3626 1474 3671 1502
rect 3699 1474 3757 1502
rect 3785 1474 3843 1502
rect 3871 1474 3929 1502
rect 3957 1474 3996 1502
rect 3626 1416 3996 1474
rect 3626 1388 3671 1416
rect 3699 1388 3757 1416
rect 3785 1388 3843 1416
rect 3871 1388 3929 1416
rect 3957 1388 3996 1416
rect 3626 1349 3996 1388
rect 4024 1502 4394 1533
rect 4024 1474 4069 1502
rect 4097 1474 4155 1502
rect 4183 1474 4241 1502
rect 4269 1474 4327 1502
rect 4355 1474 4394 1502
rect 4024 1416 4394 1474
rect 4024 1388 4069 1416
rect 4097 1388 4155 1416
rect 4183 1388 4241 1416
rect 4269 1388 4327 1416
rect 4355 1388 4394 1416
rect 4024 1349 4394 1388
rect 4422 1502 4792 1533
rect 4422 1474 4467 1502
rect 4495 1474 4553 1502
rect 4581 1474 4639 1502
rect 4667 1474 4725 1502
rect 4753 1474 4792 1502
rect 4422 1416 4792 1474
rect 4422 1388 4467 1416
rect 4495 1388 4553 1416
rect 4581 1388 4639 1416
rect 4667 1388 4725 1416
rect 4753 1388 4792 1416
rect 4422 1349 4792 1388
rect 4820 1502 5190 1533
rect 4820 1474 4865 1502
rect 4893 1474 4951 1502
rect 4979 1474 5037 1502
rect 5065 1474 5123 1502
rect 5151 1474 5190 1502
rect 4820 1416 5190 1474
rect 4820 1388 4865 1416
rect 4893 1388 4951 1416
rect 4979 1388 5037 1416
rect 5065 1388 5123 1416
rect 5151 1388 5190 1416
rect 4820 1349 5190 1388
rect 5218 1502 5588 1533
rect 5218 1474 5263 1502
rect 5291 1474 5349 1502
rect 5377 1474 5435 1502
rect 5463 1474 5521 1502
rect 5549 1474 5588 1502
rect 5218 1416 5588 1474
rect 5218 1388 5263 1416
rect 5291 1388 5349 1416
rect 5377 1388 5435 1416
rect 5463 1388 5521 1416
rect 5549 1388 5588 1416
rect 5218 1349 5588 1388
rect 5616 1502 5986 1533
rect 5616 1474 5661 1502
rect 5689 1474 5747 1502
rect 5775 1474 5833 1502
rect 5861 1474 5919 1502
rect 5947 1474 5986 1502
rect 5616 1416 5986 1474
rect 5616 1388 5661 1416
rect 5689 1388 5747 1416
rect 5775 1388 5833 1416
rect 5861 1388 5919 1416
rect 5947 1388 5986 1416
rect 5616 1349 5986 1388
rect 6014 1502 6384 1533
rect 6014 1474 6059 1502
rect 6087 1474 6145 1502
rect 6173 1474 6231 1502
rect 6259 1474 6317 1502
rect 6345 1474 6384 1502
rect 6014 1416 6384 1474
rect 6014 1388 6059 1416
rect 6087 1388 6145 1416
rect 6173 1388 6231 1416
rect 6259 1388 6317 1416
rect 6345 1388 6384 1416
rect 6014 1349 6384 1388
rect 6412 1502 6782 1533
rect 6412 1474 6457 1502
rect 6485 1474 6543 1502
rect 6571 1474 6629 1502
rect 6657 1474 6715 1502
rect 6743 1474 6782 1502
rect 6412 1416 6782 1474
rect 6412 1388 6457 1416
rect 6485 1388 6543 1416
rect 6571 1388 6629 1416
rect 6657 1388 6715 1416
rect 6743 1388 6782 1416
rect 6412 1349 6782 1388
rect 6810 1502 7180 1533
rect 6810 1474 6855 1502
rect 6883 1474 6941 1502
rect 6969 1474 7027 1502
rect 7055 1474 7113 1502
rect 7141 1474 7180 1502
rect 6810 1416 7180 1474
rect 6810 1388 6855 1416
rect 6883 1388 6941 1416
rect 6969 1388 7027 1416
rect 7055 1388 7113 1416
rect 7141 1388 7180 1416
rect 6810 1349 7180 1388
rect 7208 1502 7578 1533
rect 7208 1474 7253 1502
rect 7281 1474 7339 1502
rect 7367 1474 7425 1502
rect 7453 1474 7511 1502
rect 7539 1474 7578 1502
rect 7208 1416 7578 1474
rect 7208 1388 7253 1416
rect 7281 1388 7339 1416
rect 7367 1388 7425 1416
rect 7453 1388 7511 1416
rect 7539 1388 7578 1416
rect 7208 1349 7578 1388
rect 7606 1502 7976 1533
rect 7606 1474 7651 1502
rect 7679 1474 7737 1502
rect 7765 1474 7823 1502
rect 7851 1474 7909 1502
rect 7937 1474 7976 1502
rect 7606 1416 7976 1474
rect 7606 1388 7651 1416
rect 7679 1388 7737 1416
rect 7765 1388 7823 1416
rect 7851 1388 7909 1416
rect 7937 1388 7976 1416
rect 7606 1349 7976 1388
rect 8004 1502 8374 1533
rect 8004 1474 8049 1502
rect 8077 1474 8135 1502
rect 8163 1474 8221 1502
rect 8249 1474 8307 1502
rect 8335 1474 8374 1502
rect 8004 1416 8374 1474
rect 8004 1388 8049 1416
rect 8077 1388 8135 1416
rect 8163 1388 8221 1416
rect 8249 1388 8307 1416
rect 8335 1388 8374 1416
rect 8004 1349 8374 1388
rect 8402 1502 8772 1533
rect 8402 1474 8447 1502
rect 8475 1474 8533 1502
rect 8561 1474 8619 1502
rect 8647 1474 8705 1502
rect 8733 1474 8772 1502
rect 8402 1416 8772 1474
rect 8402 1388 8447 1416
rect 8475 1388 8533 1416
rect 8561 1388 8619 1416
rect 8647 1388 8705 1416
rect 8733 1388 8772 1416
rect 8402 1349 8772 1388
rect 8800 1502 9170 1533
rect 8800 1474 8845 1502
rect 8873 1474 8931 1502
rect 8959 1474 9017 1502
rect 9045 1474 9103 1502
rect 9131 1474 9170 1502
rect 8800 1416 9170 1474
rect 8800 1388 8845 1416
rect 8873 1388 8931 1416
rect 8959 1388 9017 1416
rect 9045 1388 9103 1416
rect 9131 1388 9170 1416
rect 8800 1349 9170 1388
rect 9198 1502 9568 1533
rect 9198 1474 9243 1502
rect 9271 1474 9329 1502
rect 9357 1474 9415 1502
rect 9443 1474 9501 1502
rect 9529 1474 9568 1502
rect 9198 1416 9568 1474
rect 9198 1388 9243 1416
rect 9271 1388 9329 1416
rect 9357 1388 9415 1416
rect 9443 1388 9501 1416
rect 9529 1388 9568 1416
rect 9198 1349 9568 1388
rect 9596 1502 9966 1533
rect 9596 1474 9641 1502
rect 9669 1474 9727 1502
rect 9755 1474 9813 1502
rect 9841 1474 9899 1502
rect 9927 1474 9966 1502
rect 9596 1416 9966 1474
rect 9596 1388 9641 1416
rect 9669 1388 9727 1416
rect 9755 1388 9813 1416
rect 9841 1388 9899 1416
rect 9927 1388 9966 1416
rect 9596 1349 9966 1388
rect 215 1285 232 1349
rect 1814 1285 1831 1349
rect 2213 1285 2230 1349
rect 3804 1285 3821 1349
rect 4199 1285 4216 1349
rect 5784 1285 5801 1349
rect 6192 1285 6209 1349
rect 7788 1285 7805 1349
rect 8182 1285 8199 1349
rect 9770 1285 9787 1349
rect 44 1240 414 1285
rect 44 1212 89 1240
rect 117 1212 175 1240
rect 203 1212 261 1240
rect 289 1212 347 1240
rect 375 1212 414 1240
rect 44 1154 414 1212
rect 44 1126 89 1154
rect 117 1126 175 1154
rect 203 1126 261 1154
rect 289 1126 347 1154
rect 375 1126 414 1154
rect 44 1068 414 1126
rect 44 1040 89 1068
rect 117 1040 175 1068
rect 203 1040 261 1068
rect 289 1040 347 1068
rect 375 1040 414 1068
rect 44 982 414 1040
rect 44 954 89 982
rect 117 954 175 982
rect 203 954 261 982
rect 289 954 347 982
rect 375 954 414 982
rect 44 915 414 954
rect 442 1240 812 1285
rect 442 1212 487 1240
rect 515 1212 573 1240
rect 601 1212 659 1240
rect 687 1212 745 1240
rect 773 1212 812 1240
rect 442 1154 812 1212
rect 442 1126 487 1154
rect 515 1126 573 1154
rect 601 1126 659 1154
rect 687 1126 745 1154
rect 773 1126 812 1154
rect 442 1103 812 1126
rect 840 1240 1210 1285
rect 840 1212 885 1240
rect 913 1212 971 1240
rect 999 1212 1057 1240
rect 1085 1212 1143 1240
rect 1171 1212 1210 1240
rect 840 1154 1210 1212
rect 840 1126 885 1154
rect 913 1126 971 1154
rect 999 1126 1057 1154
rect 1085 1126 1143 1154
rect 1171 1126 1210 1154
rect 840 1103 1210 1126
rect 1238 1240 1608 1285
rect 1238 1212 1283 1240
rect 1311 1212 1369 1240
rect 1397 1212 1455 1240
rect 1483 1212 1541 1240
rect 1569 1212 1608 1240
rect 1238 1154 1608 1212
rect 1238 1126 1283 1154
rect 1311 1126 1369 1154
rect 1397 1126 1455 1154
rect 1483 1126 1541 1154
rect 1569 1126 1608 1154
rect 1238 1103 1608 1126
rect 442 1087 1608 1103
rect 442 1068 812 1087
rect 442 1040 487 1068
rect 515 1040 573 1068
rect 601 1040 659 1068
rect 687 1040 745 1068
rect 773 1040 812 1068
rect 442 982 812 1040
rect 442 954 487 982
rect 515 954 573 982
rect 601 954 659 982
rect 687 954 745 982
rect 773 954 812 982
rect 442 915 812 954
rect 840 1068 1210 1087
rect 840 1040 885 1068
rect 913 1040 971 1068
rect 999 1040 1057 1068
rect 1085 1040 1143 1068
rect 1171 1040 1210 1068
rect 840 982 1210 1040
rect 840 954 885 982
rect 913 954 971 982
rect 999 954 1057 982
rect 1085 954 1143 982
rect 1171 954 1210 982
rect 840 915 1210 954
rect 1238 1068 1608 1087
rect 1238 1040 1283 1068
rect 1311 1040 1369 1068
rect 1397 1040 1455 1068
rect 1483 1040 1541 1068
rect 1569 1040 1608 1068
rect 1238 982 1608 1040
rect 1238 954 1283 982
rect 1311 954 1369 982
rect 1397 954 1455 982
rect 1483 954 1541 982
rect 1569 954 1608 982
rect 1238 915 1608 954
rect 1636 1240 2006 1285
rect 1636 1212 1681 1240
rect 1709 1212 1767 1240
rect 1795 1212 1853 1240
rect 1881 1212 1939 1240
rect 1967 1212 2006 1240
rect 1636 1154 2006 1212
rect 1636 1126 1681 1154
rect 1709 1126 1767 1154
rect 1795 1126 1853 1154
rect 1881 1126 1939 1154
rect 1967 1126 2006 1154
rect 1636 1068 2006 1126
rect 1636 1040 1681 1068
rect 1709 1040 1767 1068
rect 1795 1040 1853 1068
rect 1881 1040 1939 1068
rect 1967 1040 2006 1068
rect 1636 982 2006 1040
rect 1636 954 1681 982
rect 1709 954 1767 982
rect 1795 954 1853 982
rect 1881 954 1939 982
rect 1967 954 2006 982
rect 1636 915 2006 954
rect 2034 1240 2404 1285
rect 2034 1212 2079 1240
rect 2107 1212 2165 1240
rect 2193 1212 2251 1240
rect 2279 1212 2337 1240
rect 2365 1212 2404 1240
rect 2034 1154 2404 1212
rect 2034 1126 2079 1154
rect 2107 1126 2165 1154
rect 2193 1126 2251 1154
rect 2279 1126 2337 1154
rect 2365 1126 2404 1154
rect 2034 1068 2404 1126
rect 2034 1040 2079 1068
rect 2107 1040 2165 1068
rect 2193 1040 2251 1068
rect 2279 1040 2337 1068
rect 2365 1040 2404 1068
rect 2034 982 2404 1040
rect 2034 954 2079 982
rect 2107 954 2165 982
rect 2193 954 2251 982
rect 2279 954 2337 982
rect 2365 954 2404 982
rect 2034 915 2404 954
rect 2432 1240 2802 1285
rect 2432 1212 2477 1240
rect 2505 1212 2563 1240
rect 2591 1212 2649 1240
rect 2677 1212 2735 1240
rect 2763 1212 2802 1240
rect 2432 1154 2802 1212
rect 2432 1126 2477 1154
rect 2505 1126 2563 1154
rect 2591 1126 2649 1154
rect 2677 1126 2735 1154
rect 2763 1126 2802 1154
rect 2432 1102 2802 1126
rect 2830 1240 3200 1285
rect 2830 1212 2875 1240
rect 2903 1212 2961 1240
rect 2989 1212 3047 1240
rect 3075 1212 3133 1240
rect 3161 1212 3200 1240
rect 2830 1154 3200 1212
rect 2830 1126 2875 1154
rect 2903 1126 2961 1154
rect 2989 1126 3047 1154
rect 3075 1126 3133 1154
rect 3161 1126 3200 1154
rect 2830 1102 3200 1126
rect 3228 1240 3598 1285
rect 3228 1212 3273 1240
rect 3301 1212 3359 1240
rect 3387 1212 3445 1240
rect 3473 1212 3531 1240
rect 3559 1212 3598 1240
rect 3228 1154 3598 1212
rect 3228 1126 3273 1154
rect 3301 1126 3359 1154
rect 3387 1126 3445 1154
rect 3473 1126 3531 1154
rect 3559 1126 3598 1154
rect 3228 1102 3598 1126
rect 2432 1086 3598 1102
rect 2432 1068 2802 1086
rect 2432 1040 2477 1068
rect 2505 1040 2563 1068
rect 2591 1040 2649 1068
rect 2677 1040 2735 1068
rect 2763 1040 2802 1068
rect 2432 982 2802 1040
rect 2432 954 2477 982
rect 2505 954 2563 982
rect 2591 954 2649 982
rect 2677 954 2735 982
rect 2763 954 2802 982
rect 2432 915 2802 954
rect 2830 1068 3200 1086
rect 2830 1040 2875 1068
rect 2903 1040 2961 1068
rect 2989 1040 3047 1068
rect 3075 1040 3133 1068
rect 3161 1040 3200 1068
rect 2830 982 3200 1040
rect 2830 954 2875 982
rect 2903 954 2961 982
rect 2989 954 3047 982
rect 3075 954 3133 982
rect 3161 954 3200 982
rect 2830 915 3200 954
rect 3228 1068 3598 1086
rect 3228 1040 3273 1068
rect 3301 1040 3359 1068
rect 3387 1040 3445 1068
rect 3473 1040 3531 1068
rect 3559 1040 3598 1068
rect 3228 982 3598 1040
rect 3228 954 3273 982
rect 3301 954 3359 982
rect 3387 954 3445 982
rect 3473 954 3531 982
rect 3559 954 3598 982
rect 3228 915 3598 954
rect 3626 1240 3996 1285
rect 3626 1212 3671 1240
rect 3699 1212 3757 1240
rect 3785 1212 3843 1240
rect 3871 1212 3929 1240
rect 3957 1212 3996 1240
rect 3626 1154 3996 1212
rect 3626 1126 3671 1154
rect 3699 1126 3757 1154
rect 3785 1126 3843 1154
rect 3871 1126 3929 1154
rect 3957 1126 3996 1154
rect 3626 1068 3996 1126
rect 3626 1040 3671 1068
rect 3699 1040 3757 1068
rect 3785 1040 3843 1068
rect 3871 1040 3929 1068
rect 3957 1040 3996 1068
rect 3626 982 3996 1040
rect 3626 954 3671 982
rect 3699 954 3757 982
rect 3785 954 3843 982
rect 3871 954 3929 982
rect 3957 954 3996 982
rect 3626 915 3996 954
rect 4024 1240 4394 1285
rect 4024 1212 4069 1240
rect 4097 1212 4155 1240
rect 4183 1212 4241 1240
rect 4269 1212 4327 1240
rect 4355 1212 4394 1240
rect 4024 1154 4394 1212
rect 4024 1126 4069 1154
rect 4097 1126 4155 1154
rect 4183 1126 4241 1154
rect 4269 1126 4327 1154
rect 4355 1126 4394 1154
rect 4024 1068 4394 1126
rect 4024 1040 4069 1068
rect 4097 1040 4155 1068
rect 4183 1040 4241 1068
rect 4269 1040 4327 1068
rect 4355 1040 4394 1068
rect 4024 982 4394 1040
rect 4024 954 4069 982
rect 4097 954 4155 982
rect 4183 954 4241 982
rect 4269 954 4327 982
rect 4355 954 4394 982
rect 4024 915 4394 954
rect 4422 1240 4792 1285
rect 4422 1212 4467 1240
rect 4495 1212 4553 1240
rect 4581 1212 4639 1240
rect 4667 1212 4725 1240
rect 4753 1212 4792 1240
rect 4422 1154 4792 1212
rect 4422 1126 4467 1154
rect 4495 1126 4553 1154
rect 4581 1126 4639 1154
rect 4667 1126 4725 1154
rect 4753 1126 4792 1154
rect 4422 1109 4792 1126
rect 4820 1240 5190 1285
rect 4820 1212 4865 1240
rect 4893 1212 4951 1240
rect 4979 1212 5037 1240
rect 5065 1212 5123 1240
rect 5151 1212 5190 1240
rect 4820 1154 5190 1212
rect 4820 1126 4865 1154
rect 4893 1126 4951 1154
rect 4979 1126 5037 1154
rect 5065 1126 5123 1154
rect 5151 1126 5190 1154
rect 4820 1109 5190 1126
rect 5218 1240 5588 1285
rect 5218 1212 5263 1240
rect 5291 1212 5349 1240
rect 5377 1212 5435 1240
rect 5463 1212 5521 1240
rect 5549 1212 5588 1240
rect 5218 1154 5588 1212
rect 5218 1126 5263 1154
rect 5291 1126 5349 1154
rect 5377 1126 5435 1154
rect 5463 1126 5521 1154
rect 5549 1126 5588 1154
rect 5218 1109 5588 1126
rect 4422 1093 5588 1109
rect 4422 1068 4792 1093
rect 4422 1040 4467 1068
rect 4495 1040 4553 1068
rect 4581 1040 4639 1068
rect 4667 1040 4725 1068
rect 4753 1040 4792 1068
rect 4422 982 4792 1040
rect 4422 954 4467 982
rect 4495 954 4553 982
rect 4581 954 4639 982
rect 4667 954 4725 982
rect 4753 954 4792 982
rect 4422 915 4792 954
rect 4820 1068 5190 1093
rect 4820 1040 4865 1068
rect 4893 1040 4951 1068
rect 4979 1040 5037 1068
rect 5065 1040 5123 1068
rect 5151 1040 5190 1068
rect 4820 982 5190 1040
rect 4820 954 4865 982
rect 4893 954 4951 982
rect 4979 954 5037 982
rect 5065 954 5123 982
rect 5151 954 5190 982
rect 4820 915 5190 954
rect 5218 1068 5588 1093
rect 5218 1040 5263 1068
rect 5291 1040 5349 1068
rect 5377 1040 5435 1068
rect 5463 1040 5521 1068
rect 5549 1040 5588 1068
rect 5218 982 5588 1040
rect 5218 954 5263 982
rect 5291 954 5349 982
rect 5377 954 5435 982
rect 5463 954 5521 982
rect 5549 954 5588 982
rect 5218 915 5588 954
rect 5616 1240 5986 1285
rect 5616 1212 5661 1240
rect 5689 1212 5747 1240
rect 5775 1212 5833 1240
rect 5861 1212 5919 1240
rect 5947 1212 5986 1240
rect 5616 1154 5986 1212
rect 5616 1126 5661 1154
rect 5689 1126 5747 1154
rect 5775 1126 5833 1154
rect 5861 1126 5919 1154
rect 5947 1126 5986 1154
rect 5616 1068 5986 1126
rect 5616 1040 5661 1068
rect 5689 1040 5747 1068
rect 5775 1040 5833 1068
rect 5861 1040 5919 1068
rect 5947 1040 5986 1068
rect 5616 982 5986 1040
rect 5616 954 5661 982
rect 5689 954 5747 982
rect 5775 954 5833 982
rect 5861 954 5919 982
rect 5947 954 5986 982
rect 5616 915 5986 954
rect 6014 1240 6384 1285
rect 6014 1212 6059 1240
rect 6087 1212 6145 1240
rect 6173 1212 6231 1240
rect 6259 1212 6317 1240
rect 6345 1212 6384 1240
rect 6014 1154 6384 1212
rect 6014 1126 6059 1154
rect 6087 1126 6145 1154
rect 6173 1126 6231 1154
rect 6259 1126 6317 1154
rect 6345 1126 6384 1154
rect 6014 1068 6384 1126
rect 6014 1040 6059 1068
rect 6087 1040 6145 1068
rect 6173 1040 6231 1068
rect 6259 1040 6317 1068
rect 6345 1040 6384 1068
rect 6014 982 6384 1040
rect 6014 954 6059 982
rect 6087 954 6145 982
rect 6173 954 6231 982
rect 6259 954 6317 982
rect 6345 954 6384 982
rect 6014 915 6384 954
rect 6412 1240 6782 1285
rect 6412 1212 6457 1240
rect 6485 1212 6543 1240
rect 6571 1212 6629 1240
rect 6657 1212 6715 1240
rect 6743 1212 6782 1240
rect 6412 1154 6782 1212
rect 6412 1126 6457 1154
rect 6485 1126 6543 1154
rect 6571 1126 6629 1154
rect 6657 1126 6715 1154
rect 6743 1126 6782 1154
rect 6412 1102 6782 1126
rect 6810 1240 7180 1285
rect 6810 1212 6855 1240
rect 6883 1212 6941 1240
rect 6969 1212 7027 1240
rect 7055 1212 7113 1240
rect 7141 1212 7180 1240
rect 6810 1154 7180 1212
rect 6810 1126 6855 1154
rect 6883 1126 6941 1154
rect 6969 1126 7027 1154
rect 7055 1126 7113 1154
rect 7141 1126 7180 1154
rect 6810 1102 7180 1126
rect 7208 1240 7578 1285
rect 7208 1212 7253 1240
rect 7281 1212 7339 1240
rect 7367 1212 7425 1240
rect 7453 1212 7511 1240
rect 7539 1212 7578 1240
rect 7208 1154 7578 1212
rect 7208 1126 7253 1154
rect 7281 1126 7339 1154
rect 7367 1126 7425 1154
rect 7453 1126 7511 1154
rect 7539 1126 7578 1154
rect 7208 1102 7578 1126
rect 6412 1086 7578 1102
rect 6412 1068 6782 1086
rect 6412 1040 6457 1068
rect 6485 1040 6543 1068
rect 6571 1040 6629 1068
rect 6657 1040 6715 1068
rect 6743 1040 6782 1068
rect 6412 982 6782 1040
rect 6412 954 6457 982
rect 6485 954 6543 982
rect 6571 954 6629 982
rect 6657 954 6715 982
rect 6743 954 6782 982
rect 6412 915 6782 954
rect 6810 1068 7180 1086
rect 6810 1040 6855 1068
rect 6883 1040 6941 1068
rect 6969 1040 7027 1068
rect 7055 1040 7113 1068
rect 7141 1040 7180 1068
rect 6810 982 7180 1040
rect 6810 954 6855 982
rect 6883 954 6941 982
rect 6969 954 7027 982
rect 7055 954 7113 982
rect 7141 954 7180 982
rect 6810 915 7180 954
rect 7208 1068 7578 1086
rect 7208 1040 7253 1068
rect 7281 1040 7339 1068
rect 7367 1040 7425 1068
rect 7453 1040 7511 1068
rect 7539 1040 7578 1068
rect 7208 982 7578 1040
rect 7208 954 7253 982
rect 7281 954 7339 982
rect 7367 954 7425 982
rect 7453 954 7511 982
rect 7539 954 7578 982
rect 7208 915 7578 954
rect 7606 1240 7976 1285
rect 7606 1212 7651 1240
rect 7679 1212 7737 1240
rect 7765 1212 7823 1240
rect 7851 1212 7909 1240
rect 7937 1212 7976 1240
rect 7606 1154 7976 1212
rect 7606 1126 7651 1154
rect 7679 1126 7737 1154
rect 7765 1126 7823 1154
rect 7851 1126 7909 1154
rect 7937 1126 7976 1154
rect 7606 1068 7976 1126
rect 7606 1040 7651 1068
rect 7679 1040 7737 1068
rect 7765 1040 7823 1068
rect 7851 1040 7909 1068
rect 7937 1040 7976 1068
rect 7606 982 7976 1040
rect 7606 954 7651 982
rect 7679 954 7737 982
rect 7765 954 7823 982
rect 7851 954 7909 982
rect 7937 954 7976 982
rect 7606 915 7976 954
rect 8004 1240 8374 1285
rect 8004 1212 8049 1240
rect 8077 1212 8135 1240
rect 8163 1212 8221 1240
rect 8249 1212 8307 1240
rect 8335 1212 8374 1240
rect 8004 1154 8374 1212
rect 8004 1126 8049 1154
rect 8077 1126 8135 1154
rect 8163 1126 8221 1154
rect 8249 1126 8307 1154
rect 8335 1126 8374 1154
rect 8004 1068 8374 1126
rect 8004 1040 8049 1068
rect 8077 1040 8135 1068
rect 8163 1040 8221 1068
rect 8249 1040 8307 1068
rect 8335 1040 8374 1068
rect 8004 982 8374 1040
rect 8004 954 8049 982
rect 8077 954 8135 982
rect 8163 954 8221 982
rect 8249 954 8307 982
rect 8335 954 8374 982
rect 8004 915 8374 954
rect 8402 1240 8772 1285
rect 8402 1212 8447 1240
rect 8475 1212 8533 1240
rect 8561 1212 8619 1240
rect 8647 1212 8705 1240
rect 8733 1212 8772 1240
rect 8402 1154 8772 1212
rect 8402 1126 8447 1154
rect 8475 1126 8533 1154
rect 8561 1126 8619 1154
rect 8647 1126 8705 1154
rect 8733 1126 8772 1154
rect 8402 1108 8772 1126
rect 8800 1240 9170 1285
rect 8800 1212 8845 1240
rect 8873 1212 8931 1240
rect 8959 1212 9017 1240
rect 9045 1212 9103 1240
rect 9131 1212 9170 1240
rect 8800 1154 9170 1212
rect 8800 1126 8845 1154
rect 8873 1126 8931 1154
rect 8959 1126 9017 1154
rect 9045 1126 9103 1154
rect 9131 1126 9170 1154
rect 8800 1108 9170 1126
rect 9198 1240 9568 1285
rect 9198 1212 9243 1240
rect 9271 1212 9329 1240
rect 9357 1212 9415 1240
rect 9443 1212 9501 1240
rect 9529 1212 9568 1240
rect 9198 1154 9568 1212
rect 9198 1126 9243 1154
rect 9271 1126 9329 1154
rect 9357 1126 9415 1154
rect 9443 1126 9501 1154
rect 9529 1126 9568 1154
rect 9198 1108 9568 1126
rect 8402 1092 9568 1108
rect 8402 1068 8772 1092
rect 8402 1040 8447 1068
rect 8475 1040 8533 1068
rect 8561 1040 8619 1068
rect 8647 1040 8705 1068
rect 8733 1040 8772 1068
rect 8402 982 8772 1040
rect 8402 954 8447 982
rect 8475 954 8533 982
rect 8561 954 8619 982
rect 8647 954 8705 982
rect 8733 954 8772 982
rect 8402 915 8772 954
rect 8800 1068 9170 1092
rect 8800 1040 8845 1068
rect 8873 1040 8931 1068
rect 8959 1040 9017 1068
rect 9045 1040 9103 1068
rect 9131 1040 9170 1068
rect 8800 982 9170 1040
rect 8800 954 8845 982
rect 8873 954 8931 982
rect 8959 954 9017 982
rect 9045 954 9103 982
rect 9131 954 9170 982
rect 8800 915 9170 954
rect 9198 1068 9568 1092
rect 9198 1040 9243 1068
rect 9271 1040 9329 1068
rect 9357 1040 9415 1068
rect 9443 1040 9501 1068
rect 9529 1040 9568 1068
rect 9198 982 9568 1040
rect 9198 954 9243 982
rect 9271 954 9329 982
rect 9357 954 9415 982
rect 9443 954 9501 982
rect 9529 954 9568 982
rect 9198 915 9568 954
rect 9596 1240 9966 1285
rect 9596 1212 9641 1240
rect 9669 1212 9727 1240
rect 9755 1212 9813 1240
rect 9841 1212 9899 1240
rect 9927 1212 9966 1240
rect 9596 1154 9966 1212
rect 9596 1126 9641 1154
rect 9669 1126 9727 1154
rect 9755 1126 9813 1154
rect 9841 1126 9899 1154
rect 9927 1126 9966 1154
rect 9596 1068 9966 1126
rect 9596 1040 9641 1068
rect 9669 1040 9727 1068
rect 9755 1040 9813 1068
rect 9841 1040 9899 1068
rect 9927 1040 9966 1068
rect 9596 982 9966 1040
rect 9596 954 9641 982
rect 9669 954 9727 982
rect 9755 954 9813 982
rect 9841 954 9899 982
rect 9927 954 9966 982
rect 9596 915 9966 954
rect 215 851 232 915
rect 1015 851 1030 915
rect 1814 851 1831 915
rect 2213 851 2230 915
rect 3010 851 3027 915
rect 3804 851 3821 915
rect 4199 851 4216 915
rect 4999 851 5016 915
rect 5784 851 5801 915
rect 6192 851 6209 915
rect 6992 851 7009 915
rect 7788 851 7805 915
rect 8182 851 8199 915
rect 8975 851 8992 915
rect 9770 851 9787 915
rect 44 806 414 851
rect 44 778 89 806
rect 117 778 175 806
rect 203 778 261 806
rect 289 778 347 806
rect 375 778 414 806
rect 44 720 414 778
rect 44 692 89 720
rect 117 692 175 720
rect 203 692 261 720
rect 289 692 347 720
rect 375 692 414 720
rect 44 634 414 692
rect 44 606 89 634
rect 117 606 175 634
rect 203 606 261 634
rect 289 606 347 634
rect 375 606 414 634
rect 44 548 414 606
rect 44 520 89 548
rect 117 520 175 548
rect 203 520 261 548
rect 289 520 347 548
rect 375 520 414 548
rect 44 481 414 520
rect 442 806 812 851
rect 442 778 487 806
rect 515 778 573 806
rect 601 778 659 806
rect 687 778 745 806
rect 773 778 812 806
rect 442 720 812 778
rect 442 692 487 720
rect 515 692 573 720
rect 601 692 659 720
rect 687 692 745 720
rect 773 692 812 720
rect 442 668 812 692
rect 840 806 1210 851
rect 840 778 885 806
rect 913 778 971 806
rect 999 778 1057 806
rect 1085 778 1143 806
rect 1171 778 1210 806
rect 840 720 1210 778
rect 840 692 885 720
rect 913 692 971 720
rect 999 692 1057 720
rect 1085 692 1143 720
rect 1171 692 1210 720
rect 840 668 1210 692
rect 1238 806 1608 851
rect 1238 778 1283 806
rect 1311 778 1369 806
rect 1397 778 1455 806
rect 1483 778 1541 806
rect 1569 778 1608 806
rect 1238 720 1608 778
rect 1238 692 1283 720
rect 1311 692 1369 720
rect 1397 692 1455 720
rect 1483 692 1541 720
rect 1569 692 1608 720
rect 1238 668 1608 692
rect 442 652 1608 668
rect 442 634 812 652
rect 442 606 487 634
rect 515 606 573 634
rect 601 606 659 634
rect 687 606 745 634
rect 773 606 812 634
rect 442 548 812 606
rect 442 520 487 548
rect 515 520 573 548
rect 601 520 659 548
rect 687 520 745 548
rect 773 520 812 548
rect 442 481 812 520
rect 840 634 1210 652
rect 840 606 885 634
rect 913 606 971 634
rect 999 606 1057 634
rect 1085 606 1143 634
rect 1171 606 1210 634
rect 840 548 1210 606
rect 840 520 885 548
rect 913 520 971 548
rect 999 520 1057 548
rect 1085 520 1143 548
rect 1171 520 1210 548
rect 840 481 1210 520
rect 1238 634 1608 652
rect 1238 606 1283 634
rect 1311 606 1369 634
rect 1397 606 1455 634
rect 1483 606 1541 634
rect 1569 606 1608 634
rect 1238 548 1608 606
rect 1238 520 1283 548
rect 1311 520 1369 548
rect 1397 520 1455 548
rect 1483 520 1541 548
rect 1569 520 1608 548
rect 1238 481 1608 520
rect 1636 806 2006 851
rect 1636 778 1681 806
rect 1709 778 1767 806
rect 1795 778 1853 806
rect 1881 778 1939 806
rect 1967 778 2006 806
rect 1636 720 2006 778
rect 1636 692 1681 720
rect 1709 692 1767 720
rect 1795 692 1853 720
rect 1881 692 1939 720
rect 1967 692 2006 720
rect 1636 634 2006 692
rect 1636 606 1681 634
rect 1709 606 1767 634
rect 1795 606 1853 634
rect 1881 606 1939 634
rect 1967 606 2006 634
rect 1636 548 2006 606
rect 1636 520 1681 548
rect 1709 520 1767 548
rect 1795 520 1853 548
rect 1881 520 1939 548
rect 1967 520 2006 548
rect 1636 481 2006 520
rect 2034 806 2404 851
rect 2034 778 2079 806
rect 2107 778 2165 806
rect 2193 778 2251 806
rect 2279 778 2337 806
rect 2365 778 2404 806
rect 2034 720 2404 778
rect 2034 692 2079 720
rect 2107 692 2165 720
rect 2193 692 2251 720
rect 2279 692 2337 720
rect 2365 692 2404 720
rect 2034 634 2404 692
rect 2034 606 2079 634
rect 2107 606 2165 634
rect 2193 606 2251 634
rect 2279 606 2337 634
rect 2365 606 2404 634
rect 2034 548 2404 606
rect 2034 520 2079 548
rect 2107 520 2165 548
rect 2193 520 2251 548
rect 2279 520 2337 548
rect 2365 520 2404 548
rect 2034 481 2404 520
rect 2432 806 2802 851
rect 2432 778 2477 806
rect 2505 778 2563 806
rect 2591 778 2649 806
rect 2677 778 2735 806
rect 2763 778 2802 806
rect 2432 720 2802 778
rect 2432 692 2477 720
rect 2505 692 2563 720
rect 2591 692 2649 720
rect 2677 692 2735 720
rect 2763 692 2802 720
rect 2432 674 2802 692
rect 2830 806 3200 851
rect 2830 778 2875 806
rect 2903 778 2961 806
rect 2989 778 3047 806
rect 3075 778 3133 806
rect 3161 778 3200 806
rect 2830 720 3200 778
rect 2830 692 2875 720
rect 2903 692 2961 720
rect 2989 692 3047 720
rect 3075 692 3133 720
rect 3161 692 3200 720
rect 2830 674 3200 692
rect 3228 806 3598 851
rect 3228 778 3273 806
rect 3301 778 3359 806
rect 3387 778 3445 806
rect 3473 778 3531 806
rect 3559 778 3598 806
rect 3228 720 3598 778
rect 3228 692 3273 720
rect 3301 692 3359 720
rect 3387 692 3445 720
rect 3473 692 3531 720
rect 3559 692 3598 720
rect 3228 674 3598 692
rect 2432 658 3598 674
rect 2432 634 2802 658
rect 2432 606 2477 634
rect 2505 606 2563 634
rect 2591 606 2649 634
rect 2677 606 2735 634
rect 2763 606 2802 634
rect 2432 548 2802 606
rect 2432 520 2477 548
rect 2505 520 2563 548
rect 2591 520 2649 548
rect 2677 520 2735 548
rect 2763 520 2802 548
rect 2432 481 2802 520
rect 2830 634 3200 658
rect 2830 606 2875 634
rect 2903 606 2961 634
rect 2989 606 3047 634
rect 3075 606 3133 634
rect 3161 606 3200 634
rect 2830 548 3200 606
rect 2830 520 2875 548
rect 2903 520 2961 548
rect 2989 520 3047 548
rect 3075 520 3133 548
rect 3161 520 3200 548
rect 2830 481 3200 520
rect 3228 634 3598 658
rect 3228 606 3273 634
rect 3301 606 3359 634
rect 3387 606 3445 634
rect 3473 606 3531 634
rect 3559 606 3598 634
rect 3228 548 3598 606
rect 3228 520 3273 548
rect 3301 520 3359 548
rect 3387 520 3445 548
rect 3473 520 3531 548
rect 3559 520 3598 548
rect 3228 481 3598 520
rect 3626 806 3996 851
rect 3626 778 3671 806
rect 3699 778 3757 806
rect 3785 778 3843 806
rect 3871 778 3929 806
rect 3957 778 3996 806
rect 3626 720 3996 778
rect 3626 692 3671 720
rect 3699 692 3757 720
rect 3785 692 3843 720
rect 3871 692 3929 720
rect 3957 692 3996 720
rect 3626 634 3996 692
rect 3626 606 3671 634
rect 3699 606 3757 634
rect 3785 606 3843 634
rect 3871 606 3929 634
rect 3957 606 3996 634
rect 3626 548 3996 606
rect 3626 520 3671 548
rect 3699 520 3757 548
rect 3785 520 3843 548
rect 3871 520 3929 548
rect 3957 520 3996 548
rect 3626 481 3996 520
rect 4024 806 4394 851
rect 4024 778 4069 806
rect 4097 778 4155 806
rect 4183 778 4241 806
rect 4269 778 4327 806
rect 4355 778 4394 806
rect 4024 720 4394 778
rect 4024 692 4069 720
rect 4097 692 4155 720
rect 4183 692 4241 720
rect 4269 692 4327 720
rect 4355 692 4394 720
rect 4024 634 4394 692
rect 4024 606 4069 634
rect 4097 606 4155 634
rect 4183 606 4241 634
rect 4269 606 4327 634
rect 4355 606 4394 634
rect 4024 548 4394 606
rect 4024 520 4069 548
rect 4097 520 4155 548
rect 4183 520 4241 548
rect 4269 520 4327 548
rect 4355 520 4394 548
rect 4024 481 4394 520
rect 4422 806 4792 851
rect 4422 778 4467 806
rect 4495 778 4553 806
rect 4581 778 4639 806
rect 4667 778 4725 806
rect 4753 778 4792 806
rect 4422 720 4792 778
rect 4422 692 4467 720
rect 4495 692 4553 720
rect 4581 692 4639 720
rect 4667 692 4725 720
rect 4753 692 4792 720
rect 4422 674 4792 692
rect 4820 806 5190 851
rect 4820 778 4865 806
rect 4893 778 4951 806
rect 4979 778 5037 806
rect 5065 778 5123 806
rect 5151 778 5190 806
rect 4820 720 5190 778
rect 4820 692 4865 720
rect 4893 692 4951 720
rect 4979 692 5037 720
rect 5065 692 5123 720
rect 5151 692 5190 720
rect 4820 674 5190 692
rect 5218 806 5588 851
rect 5218 778 5263 806
rect 5291 778 5349 806
rect 5377 778 5435 806
rect 5463 778 5521 806
rect 5549 778 5588 806
rect 5218 720 5588 778
rect 5218 692 5263 720
rect 5291 692 5349 720
rect 5377 692 5435 720
rect 5463 692 5521 720
rect 5549 692 5588 720
rect 5218 674 5588 692
rect 4422 658 5588 674
rect 4422 634 4792 658
rect 4422 606 4467 634
rect 4495 606 4553 634
rect 4581 606 4639 634
rect 4667 606 4725 634
rect 4753 606 4792 634
rect 4422 548 4792 606
rect 4422 520 4467 548
rect 4495 520 4553 548
rect 4581 520 4639 548
rect 4667 520 4725 548
rect 4753 520 4792 548
rect 4422 481 4792 520
rect 4820 634 5190 658
rect 4820 606 4865 634
rect 4893 606 4951 634
rect 4979 606 5037 634
rect 5065 606 5123 634
rect 5151 606 5190 634
rect 4820 548 5190 606
rect 4820 520 4865 548
rect 4893 520 4951 548
rect 4979 520 5037 548
rect 5065 520 5123 548
rect 5151 520 5190 548
rect 4820 481 5190 520
rect 5218 634 5588 658
rect 5218 606 5263 634
rect 5291 606 5349 634
rect 5377 606 5435 634
rect 5463 606 5521 634
rect 5549 606 5588 634
rect 5218 548 5588 606
rect 5218 520 5263 548
rect 5291 520 5349 548
rect 5377 520 5435 548
rect 5463 520 5521 548
rect 5549 520 5588 548
rect 5218 481 5588 520
rect 5616 806 5986 851
rect 5616 778 5661 806
rect 5689 778 5747 806
rect 5775 778 5833 806
rect 5861 778 5919 806
rect 5947 778 5986 806
rect 5616 720 5986 778
rect 5616 692 5661 720
rect 5689 692 5747 720
rect 5775 692 5833 720
rect 5861 692 5919 720
rect 5947 692 5986 720
rect 5616 634 5986 692
rect 5616 606 5661 634
rect 5689 606 5747 634
rect 5775 606 5833 634
rect 5861 606 5919 634
rect 5947 606 5986 634
rect 5616 548 5986 606
rect 5616 520 5661 548
rect 5689 520 5747 548
rect 5775 520 5833 548
rect 5861 520 5919 548
rect 5947 520 5986 548
rect 5616 481 5986 520
rect 6014 806 6384 851
rect 6014 778 6059 806
rect 6087 778 6145 806
rect 6173 778 6231 806
rect 6259 778 6317 806
rect 6345 778 6384 806
rect 6014 720 6384 778
rect 6014 692 6059 720
rect 6087 692 6145 720
rect 6173 692 6231 720
rect 6259 692 6317 720
rect 6345 692 6384 720
rect 6014 634 6384 692
rect 6014 606 6059 634
rect 6087 606 6145 634
rect 6173 606 6231 634
rect 6259 606 6317 634
rect 6345 606 6384 634
rect 6014 548 6384 606
rect 6014 520 6059 548
rect 6087 520 6145 548
rect 6173 520 6231 548
rect 6259 520 6317 548
rect 6345 520 6384 548
rect 6014 481 6384 520
rect 6412 806 6782 851
rect 6412 778 6457 806
rect 6485 778 6543 806
rect 6571 778 6629 806
rect 6657 778 6715 806
rect 6743 778 6782 806
rect 6412 720 6782 778
rect 6412 692 6457 720
rect 6485 692 6543 720
rect 6571 692 6629 720
rect 6657 692 6715 720
rect 6743 692 6782 720
rect 6412 672 6782 692
rect 6810 806 7180 851
rect 6810 778 6855 806
rect 6883 778 6941 806
rect 6969 778 7027 806
rect 7055 778 7113 806
rect 7141 778 7180 806
rect 6810 720 7180 778
rect 6810 692 6855 720
rect 6883 692 6941 720
rect 6969 692 7027 720
rect 7055 692 7113 720
rect 7141 692 7180 720
rect 6810 672 7180 692
rect 7208 806 7578 851
rect 7208 778 7253 806
rect 7281 778 7339 806
rect 7367 778 7425 806
rect 7453 778 7511 806
rect 7539 778 7578 806
rect 7208 720 7578 778
rect 7208 692 7253 720
rect 7281 692 7339 720
rect 7367 692 7425 720
rect 7453 692 7511 720
rect 7539 692 7578 720
rect 7208 672 7578 692
rect 6412 656 7578 672
rect 6412 634 6782 656
rect 6412 606 6457 634
rect 6485 606 6543 634
rect 6571 606 6629 634
rect 6657 606 6715 634
rect 6743 606 6782 634
rect 6412 548 6782 606
rect 6412 520 6457 548
rect 6485 520 6543 548
rect 6571 520 6629 548
rect 6657 520 6715 548
rect 6743 520 6782 548
rect 6412 481 6782 520
rect 6810 634 7180 656
rect 6810 606 6855 634
rect 6883 606 6941 634
rect 6969 606 7027 634
rect 7055 606 7113 634
rect 7141 606 7180 634
rect 6810 548 7180 606
rect 6810 520 6855 548
rect 6883 520 6941 548
rect 6969 520 7027 548
rect 7055 520 7113 548
rect 7141 520 7180 548
rect 6810 481 7180 520
rect 7208 634 7578 656
rect 7208 606 7253 634
rect 7281 606 7339 634
rect 7367 606 7425 634
rect 7453 606 7511 634
rect 7539 606 7578 634
rect 7208 548 7578 606
rect 7208 520 7253 548
rect 7281 520 7339 548
rect 7367 520 7425 548
rect 7453 520 7511 548
rect 7539 520 7578 548
rect 7208 481 7578 520
rect 7606 806 7976 851
rect 7606 778 7651 806
rect 7679 778 7737 806
rect 7765 778 7823 806
rect 7851 778 7909 806
rect 7937 778 7976 806
rect 7606 720 7976 778
rect 7606 692 7651 720
rect 7679 692 7737 720
rect 7765 692 7823 720
rect 7851 692 7909 720
rect 7937 692 7976 720
rect 7606 634 7976 692
rect 7606 606 7651 634
rect 7679 606 7737 634
rect 7765 606 7823 634
rect 7851 606 7909 634
rect 7937 606 7976 634
rect 7606 548 7976 606
rect 7606 520 7651 548
rect 7679 520 7737 548
rect 7765 520 7823 548
rect 7851 520 7909 548
rect 7937 520 7976 548
rect 7606 481 7976 520
rect 8004 806 8374 851
rect 8004 778 8049 806
rect 8077 778 8135 806
rect 8163 778 8221 806
rect 8249 778 8307 806
rect 8335 778 8374 806
rect 8004 720 8374 778
rect 8004 692 8049 720
rect 8077 692 8135 720
rect 8163 692 8221 720
rect 8249 692 8307 720
rect 8335 692 8374 720
rect 8004 634 8374 692
rect 8004 606 8049 634
rect 8077 606 8135 634
rect 8163 606 8221 634
rect 8249 606 8307 634
rect 8335 606 8374 634
rect 8004 548 8374 606
rect 8004 520 8049 548
rect 8077 520 8135 548
rect 8163 520 8221 548
rect 8249 520 8307 548
rect 8335 520 8374 548
rect 8004 481 8374 520
rect 8402 806 8772 851
rect 8402 778 8447 806
rect 8475 778 8533 806
rect 8561 778 8619 806
rect 8647 778 8705 806
rect 8733 778 8772 806
rect 8402 720 8772 778
rect 8402 692 8447 720
rect 8475 692 8533 720
rect 8561 692 8619 720
rect 8647 692 8705 720
rect 8733 692 8772 720
rect 8402 674 8772 692
rect 8800 806 9170 851
rect 8800 778 8845 806
rect 8873 778 8931 806
rect 8959 778 9017 806
rect 9045 778 9103 806
rect 9131 778 9170 806
rect 8800 720 9170 778
rect 8800 692 8845 720
rect 8873 692 8931 720
rect 8959 692 9017 720
rect 9045 692 9103 720
rect 9131 692 9170 720
rect 8800 674 9170 692
rect 9198 806 9568 851
rect 9198 778 9243 806
rect 9271 778 9329 806
rect 9357 778 9415 806
rect 9443 778 9501 806
rect 9529 778 9568 806
rect 9198 720 9568 778
rect 9198 692 9243 720
rect 9271 692 9329 720
rect 9357 692 9415 720
rect 9443 692 9501 720
rect 9529 692 9568 720
rect 9198 674 9568 692
rect 8402 658 9568 674
rect 8402 634 8772 658
rect 8402 606 8447 634
rect 8475 606 8533 634
rect 8561 606 8619 634
rect 8647 606 8705 634
rect 8733 606 8772 634
rect 8402 548 8772 606
rect 8402 520 8447 548
rect 8475 520 8533 548
rect 8561 520 8619 548
rect 8647 520 8705 548
rect 8733 520 8772 548
rect 8402 481 8772 520
rect 8800 634 9170 658
rect 8800 606 8845 634
rect 8873 606 8931 634
rect 8959 606 9017 634
rect 9045 606 9103 634
rect 9131 606 9170 634
rect 8800 548 9170 606
rect 8800 520 8845 548
rect 8873 520 8931 548
rect 8959 520 9017 548
rect 9045 520 9103 548
rect 9131 520 9170 548
rect 8800 481 9170 520
rect 9198 634 9568 658
rect 9198 606 9243 634
rect 9271 606 9329 634
rect 9357 606 9415 634
rect 9443 606 9501 634
rect 9529 606 9568 634
rect 9198 548 9568 606
rect 9198 520 9243 548
rect 9271 520 9329 548
rect 9357 520 9415 548
rect 9443 520 9501 548
rect 9529 520 9568 548
rect 9198 481 9568 520
rect 9596 806 9966 851
rect 9596 778 9641 806
rect 9669 778 9727 806
rect 9755 778 9813 806
rect 9841 778 9899 806
rect 9927 778 9966 806
rect 9596 720 9966 778
rect 9596 692 9641 720
rect 9669 692 9727 720
rect 9755 692 9813 720
rect 9841 692 9899 720
rect 9927 692 9966 720
rect 9596 634 9966 692
rect 9596 606 9641 634
rect 9669 606 9727 634
rect 9755 606 9813 634
rect 9841 606 9899 634
rect 9927 606 9966 634
rect 9596 548 9966 606
rect 9596 520 9641 548
rect 9669 520 9727 548
rect 9755 520 9813 548
rect 9841 520 9899 548
rect 9927 520 9966 548
rect 9596 481 9966 520
rect 215 417 232 481
rect 1814 417 1831 481
rect 2213 417 2230 481
rect 3010 417 3027 481
rect 3804 417 3821 481
rect 4199 417 4216 481
rect 4999 417 5016 481
rect 5784 417 5801 481
rect 6192 417 6209 481
rect 6992 417 7009 481
rect 7788 417 7805 481
rect 8182 417 8199 481
rect 8975 417 8992 481
rect 9770 417 9787 481
rect 44 372 414 417
rect 44 344 89 372
rect 117 344 175 372
rect 203 344 261 372
rect 289 344 347 372
rect 375 344 414 372
rect 44 286 414 344
rect 44 258 89 286
rect 117 258 175 286
rect 203 258 261 286
rect 289 258 347 286
rect 375 258 414 286
rect 44 236 414 258
rect 442 372 812 417
rect 442 344 487 372
rect 515 344 573 372
rect 601 344 659 372
rect 687 344 745 372
rect 773 344 812 372
rect 442 286 812 344
rect 442 258 487 286
rect 515 258 573 286
rect 601 258 659 286
rect 687 258 745 286
rect 773 258 812 286
rect 442 236 812 258
rect 840 372 1210 417
rect 840 344 885 372
rect 913 344 971 372
rect 999 344 1057 372
rect 1085 344 1143 372
rect 1171 344 1210 372
rect 840 286 1210 344
rect 840 258 885 286
rect 913 258 971 286
rect 999 258 1057 286
rect 1085 258 1143 286
rect 1171 258 1210 286
rect 840 236 1210 258
rect 1238 372 1608 417
rect 1238 344 1283 372
rect 1311 344 1369 372
rect 1397 344 1455 372
rect 1483 344 1541 372
rect 1569 344 1608 372
rect 1238 286 1608 344
rect 1238 258 1283 286
rect 1311 258 1369 286
rect 1397 258 1455 286
rect 1483 258 1541 286
rect 1569 258 1608 286
rect 1238 236 1608 258
rect 1636 372 2006 417
rect 1636 344 1681 372
rect 1709 344 1767 372
rect 1795 344 1853 372
rect 1881 344 1939 372
rect 1967 344 2006 372
rect 1636 286 2006 344
rect 1636 258 1681 286
rect 1709 258 1767 286
rect 1795 258 1853 286
rect 1881 258 1939 286
rect 1967 258 2006 286
rect 1636 236 2006 258
rect 2034 372 2404 417
rect 2034 344 2079 372
rect 2107 344 2165 372
rect 2193 344 2251 372
rect 2279 344 2337 372
rect 2365 344 2404 372
rect 2034 286 2404 344
rect 2034 258 2079 286
rect 2107 258 2165 286
rect 2193 258 2251 286
rect 2279 258 2337 286
rect 2365 258 2404 286
rect 2034 236 2404 258
rect 2432 372 2802 417
rect 2432 344 2477 372
rect 2505 344 2563 372
rect 2591 344 2649 372
rect 2677 344 2735 372
rect 2763 344 2802 372
rect 2432 286 2802 344
rect 2432 258 2477 286
rect 2505 258 2563 286
rect 2591 258 2649 286
rect 2677 258 2735 286
rect 2763 258 2802 286
rect 2432 236 2802 258
rect 44 209 2802 236
rect 44 200 414 209
rect 44 172 89 200
rect 117 172 175 200
rect 203 172 261 200
rect 289 172 347 200
rect 375 172 414 200
rect 44 114 414 172
rect 44 86 89 114
rect 117 86 175 114
rect 203 86 261 114
rect 289 86 347 114
rect 375 86 414 114
rect 44 47 414 86
rect 442 200 812 209
rect 442 172 487 200
rect 515 172 573 200
rect 601 172 659 200
rect 687 172 745 200
rect 773 172 812 200
rect 442 114 812 172
rect 442 86 487 114
rect 515 86 573 114
rect 601 86 659 114
rect 687 86 745 114
rect 773 86 812 114
rect 442 47 812 86
rect 840 200 1210 209
rect 840 172 885 200
rect 913 172 971 200
rect 999 172 1057 200
rect 1085 172 1143 200
rect 1171 172 1210 200
rect 840 114 1210 172
rect 840 86 885 114
rect 913 86 971 114
rect 999 86 1057 114
rect 1085 86 1143 114
rect 1171 86 1210 114
rect 840 47 1210 86
rect 1238 200 1608 209
rect 1238 172 1283 200
rect 1311 172 1369 200
rect 1397 172 1455 200
rect 1483 172 1541 200
rect 1569 172 1608 200
rect 1238 114 1608 172
rect 1238 86 1283 114
rect 1311 86 1369 114
rect 1397 86 1455 114
rect 1483 86 1541 114
rect 1569 86 1608 114
rect 1238 47 1608 86
rect 1636 200 2006 209
rect 1636 172 1681 200
rect 1709 172 1767 200
rect 1795 172 1853 200
rect 1881 172 1939 200
rect 1967 172 2006 200
rect 1636 114 2006 172
rect 1636 86 1681 114
rect 1709 86 1767 114
rect 1795 86 1853 114
rect 1881 86 1939 114
rect 1967 86 2006 114
rect 1636 47 2006 86
rect 2034 200 2404 209
rect 2034 172 2079 200
rect 2107 172 2165 200
rect 2193 172 2251 200
rect 2279 172 2337 200
rect 2365 172 2404 200
rect 2034 114 2404 172
rect 2034 86 2079 114
rect 2107 86 2165 114
rect 2193 86 2251 114
rect 2279 86 2337 114
rect 2365 86 2404 114
rect 2034 47 2404 86
rect 2432 200 2802 209
rect 2432 172 2477 200
rect 2505 172 2563 200
rect 2591 172 2649 200
rect 2677 172 2735 200
rect 2763 172 2802 200
rect 2432 114 2802 172
rect 2432 86 2477 114
rect 2505 86 2563 114
rect 2591 86 2649 114
rect 2677 86 2735 114
rect 2763 86 2802 114
rect 2432 47 2802 86
rect 2830 372 3200 417
rect 2830 344 2875 372
rect 2903 344 2961 372
rect 2989 344 3047 372
rect 3075 344 3133 372
rect 3161 344 3200 372
rect 2830 286 3200 344
rect 2830 258 2875 286
rect 2903 258 2961 286
rect 2989 258 3047 286
rect 3075 258 3133 286
rect 3161 258 3200 286
rect 2830 200 3200 258
rect 2830 172 2875 200
rect 2903 172 2961 200
rect 2989 172 3047 200
rect 3075 172 3133 200
rect 3161 172 3200 200
rect 2830 114 3200 172
rect 2830 86 2875 114
rect 2903 86 2961 114
rect 2989 86 3047 114
rect 3075 86 3133 114
rect 3161 86 3200 114
rect 2830 47 3200 86
rect 3228 372 3598 417
rect 3228 344 3273 372
rect 3301 344 3359 372
rect 3387 344 3445 372
rect 3473 344 3531 372
rect 3559 344 3598 372
rect 3228 286 3598 344
rect 3228 258 3273 286
rect 3301 258 3359 286
rect 3387 258 3445 286
rect 3473 258 3531 286
rect 3559 258 3598 286
rect 3228 236 3598 258
rect 3626 372 3996 417
rect 3626 344 3671 372
rect 3699 344 3757 372
rect 3785 344 3843 372
rect 3871 344 3929 372
rect 3957 344 3996 372
rect 3626 286 3996 344
rect 3626 258 3671 286
rect 3699 258 3757 286
rect 3785 258 3843 286
rect 3871 258 3929 286
rect 3957 258 3996 286
rect 3626 236 3996 258
rect 4024 372 4394 417
rect 4024 344 4069 372
rect 4097 344 4155 372
rect 4183 344 4241 372
rect 4269 344 4327 372
rect 4355 344 4394 372
rect 4024 286 4394 344
rect 4024 258 4069 286
rect 4097 258 4155 286
rect 4183 258 4241 286
rect 4269 258 4327 286
rect 4355 258 4394 286
rect 4024 236 4394 258
rect 4422 372 4792 417
rect 4422 344 4467 372
rect 4495 344 4553 372
rect 4581 344 4639 372
rect 4667 344 4725 372
rect 4753 344 4792 372
rect 4422 286 4792 344
rect 4422 258 4467 286
rect 4495 258 4553 286
rect 4581 258 4639 286
rect 4667 258 4725 286
rect 4753 258 4792 286
rect 4422 236 4792 258
rect 3228 209 4792 236
rect 3228 200 3598 209
rect 3228 172 3273 200
rect 3301 172 3359 200
rect 3387 172 3445 200
rect 3473 172 3531 200
rect 3559 172 3598 200
rect 3228 114 3598 172
rect 3228 86 3273 114
rect 3301 86 3359 114
rect 3387 86 3445 114
rect 3473 86 3531 114
rect 3559 86 3598 114
rect 3228 47 3598 86
rect 3626 200 3996 209
rect 3626 172 3671 200
rect 3699 172 3757 200
rect 3785 172 3843 200
rect 3871 172 3929 200
rect 3957 172 3996 200
rect 3626 114 3996 172
rect 3626 86 3671 114
rect 3699 86 3757 114
rect 3785 86 3843 114
rect 3871 86 3929 114
rect 3957 86 3996 114
rect 3626 47 3996 86
rect 4024 200 4394 209
rect 4024 172 4069 200
rect 4097 172 4155 200
rect 4183 172 4241 200
rect 4269 172 4327 200
rect 4355 172 4394 200
rect 4024 114 4394 172
rect 4024 86 4069 114
rect 4097 86 4155 114
rect 4183 86 4241 114
rect 4269 86 4327 114
rect 4355 86 4394 114
rect 4024 47 4394 86
rect 4422 200 4792 209
rect 4422 172 4467 200
rect 4495 172 4553 200
rect 4581 172 4639 200
rect 4667 172 4725 200
rect 4753 172 4792 200
rect 4422 114 4792 172
rect 4422 86 4467 114
rect 4495 86 4553 114
rect 4581 86 4639 114
rect 4667 86 4725 114
rect 4753 86 4792 114
rect 4422 47 4792 86
rect 4820 372 5190 417
rect 4820 344 4865 372
rect 4893 344 4951 372
rect 4979 344 5037 372
rect 5065 344 5123 372
rect 5151 344 5190 372
rect 4820 286 5190 344
rect 4820 258 4865 286
rect 4893 258 4951 286
rect 4979 258 5037 286
rect 5065 258 5123 286
rect 5151 258 5190 286
rect 4820 200 5190 258
rect 4820 172 4865 200
rect 4893 172 4951 200
rect 4979 172 5037 200
rect 5065 172 5123 200
rect 5151 172 5190 200
rect 4820 114 5190 172
rect 4820 86 4865 114
rect 4893 86 4951 114
rect 4979 86 5037 114
rect 5065 86 5123 114
rect 5151 86 5190 114
rect 4820 47 5190 86
rect 5218 372 5588 417
rect 5218 344 5263 372
rect 5291 344 5349 372
rect 5377 344 5435 372
rect 5463 344 5521 372
rect 5549 344 5588 372
rect 5218 286 5588 344
rect 5218 258 5263 286
rect 5291 258 5349 286
rect 5377 258 5435 286
rect 5463 258 5521 286
rect 5549 258 5588 286
rect 5218 236 5588 258
rect 5616 372 5986 417
rect 5616 344 5661 372
rect 5689 344 5747 372
rect 5775 344 5833 372
rect 5861 344 5919 372
rect 5947 344 5986 372
rect 5616 286 5986 344
rect 5616 258 5661 286
rect 5689 258 5747 286
rect 5775 258 5833 286
rect 5861 258 5919 286
rect 5947 258 5986 286
rect 5616 236 5986 258
rect 6014 372 6384 417
rect 6014 344 6059 372
rect 6087 344 6145 372
rect 6173 344 6231 372
rect 6259 344 6317 372
rect 6345 344 6384 372
rect 6014 286 6384 344
rect 6014 258 6059 286
rect 6087 258 6145 286
rect 6173 258 6231 286
rect 6259 258 6317 286
rect 6345 258 6384 286
rect 6014 236 6384 258
rect 6412 372 6782 417
rect 6412 344 6457 372
rect 6485 344 6543 372
rect 6571 344 6629 372
rect 6657 344 6715 372
rect 6743 344 6782 372
rect 6412 286 6782 344
rect 6412 258 6457 286
rect 6485 258 6543 286
rect 6571 258 6629 286
rect 6657 258 6715 286
rect 6743 258 6782 286
rect 6412 236 6782 258
rect 5218 209 6782 236
rect 5218 200 5588 209
rect 5218 172 5263 200
rect 5291 172 5349 200
rect 5377 172 5435 200
rect 5463 172 5521 200
rect 5549 172 5588 200
rect 5218 114 5588 172
rect 5218 86 5263 114
rect 5291 86 5349 114
rect 5377 86 5435 114
rect 5463 86 5521 114
rect 5549 86 5588 114
rect 5218 47 5588 86
rect 5616 200 5986 209
rect 5616 172 5661 200
rect 5689 172 5747 200
rect 5775 172 5833 200
rect 5861 172 5919 200
rect 5947 172 5986 200
rect 5616 114 5986 172
rect 5616 86 5661 114
rect 5689 86 5747 114
rect 5775 86 5833 114
rect 5861 86 5919 114
rect 5947 86 5986 114
rect 5616 47 5986 86
rect 6014 200 6384 209
rect 6014 172 6059 200
rect 6087 172 6145 200
rect 6173 172 6231 200
rect 6259 172 6317 200
rect 6345 172 6384 200
rect 6014 114 6384 172
rect 6014 86 6059 114
rect 6087 86 6145 114
rect 6173 86 6231 114
rect 6259 86 6317 114
rect 6345 86 6384 114
rect 6014 47 6384 86
rect 6412 200 6782 209
rect 6412 172 6457 200
rect 6485 172 6543 200
rect 6571 172 6629 200
rect 6657 172 6715 200
rect 6743 172 6782 200
rect 6412 114 6782 172
rect 6412 86 6457 114
rect 6485 86 6543 114
rect 6571 86 6629 114
rect 6657 86 6715 114
rect 6743 86 6782 114
rect 6412 47 6782 86
rect 6810 372 7180 417
rect 6810 344 6855 372
rect 6883 344 6941 372
rect 6969 344 7027 372
rect 7055 344 7113 372
rect 7141 344 7180 372
rect 6810 286 7180 344
rect 6810 258 6855 286
rect 6883 258 6941 286
rect 6969 258 7027 286
rect 7055 258 7113 286
rect 7141 258 7180 286
rect 6810 200 7180 258
rect 6810 172 6855 200
rect 6883 172 6941 200
rect 6969 172 7027 200
rect 7055 172 7113 200
rect 7141 172 7180 200
rect 6810 114 7180 172
rect 6810 86 6855 114
rect 6883 86 6941 114
rect 6969 86 7027 114
rect 7055 86 7113 114
rect 7141 86 7180 114
rect 6810 47 7180 86
rect 7208 372 7578 417
rect 7208 344 7253 372
rect 7281 344 7339 372
rect 7367 344 7425 372
rect 7453 344 7511 372
rect 7539 344 7578 372
rect 7208 286 7578 344
rect 7208 258 7253 286
rect 7281 258 7339 286
rect 7367 258 7425 286
rect 7453 258 7511 286
rect 7539 258 7578 286
rect 7208 236 7578 258
rect 7606 372 7976 417
rect 7606 344 7651 372
rect 7679 344 7737 372
rect 7765 344 7823 372
rect 7851 344 7909 372
rect 7937 344 7976 372
rect 7606 286 7976 344
rect 7606 258 7651 286
rect 7679 258 7737 286
rect 7765 258 7823 286
rect 7851 258 7909 286
rect 7937 258 7976 286
rect 7606 236 7976 258
rect 8004 372 8374 417
rect 8004 344 8049 372
rect 8077 344 8135 372
rect 8163 344 8221 372
rect 8249 344 8307 372
rect 8335 344 8374 372
rect 8004 286 8374 344
rect 8004 258 8049 286
rect 8077 258 8135 286
rect 8163 258 8221 286
rect 8249 258 8307 286
rect 8335 258 8374 286
rect 8004 236 8374 258
rect 8402 372 8772 417
rect 8402 344 8447 372
rect 8475 344 8533 372
rect 8561 344 8619 372
rect 8647 344 8705 372
rect 8733 344 8772 372
rect 8402 286 8772 344
rect 8402 258 8447 286
rect 8475 258 8533 286
rect 8561 258 8619 286
rect 8647 258 8705 286
rect 8733 258 8772 286
rect 8402 236 8772 258
rect 7208 209 8772 236
rect 7208 200 7578 209
rect 7208 172 7253 200
rect 7281 172 7339 200
rect 7367 172 7425 200
rect 7453 172 7511 200
rect 7539 172 7578 200
rect 7208 114 7578 172
rect 7208 86 7253 114
rect 7281 86 7339 114
rect 7367 86 7425 114
rect 7453 86 7511 114
rect 7539 86 7578 114
rect 7208 47 7578 86
rect 7606 200 7976 209
rect 7606 172 7651 200
rect 7679 172 7737 200
rect 7765 172 7823 200
rect 7851 172 7909 200
rect 7937 172 7976 200
rect 7606 114 7976 172
rect 7606 86 7651 114
rect 7679 86 7737 114
rect 7765 86 7823 114
rect 7851 86 7909 114
rect 7937 86 7976 114
rect 7606 47 7976 86
rect 8004 200 8374 209
rect 8004 172 8049 200
rect 8077 172 8135 200
rect 8163 172 8221 200
rect 8249 172 8307 200
rect 8335 172 8374 200
rect 8004 114 8374 172
rect 8004 86 8049 114
rect 8077 86 8135 114
rect 8163 86 8221 114
rect 8249 86 8307 114
rect 8335 86 8374 114
rect 8004 47 8374 86
rect 8402 200 8772 209
rect 8402 172 8447 200
rect 8475 172 8533 200
rect 8561 172 8619 200
rect 8647 172 8705 200
rect 8733 172 8772 200
rect 8402 114 8772 172
rect 8402 86 8447 114
rect 8475 86 8533 114
rect 8561 86 8619 114
rect 8647 86 8705 114
rect 8733 86 8772 114
rect 8402 47 8772 86
rect 8800 372 9170 417
rect 8800 344 8845 372
rect 8873 344 8931 372
rect 8959 344 9017 372
rect 9045 344 9103 372
rect 9131 344 9170 372
rect 8800 286 9170 344
rect 8800 258 8845 286
rect 8873 258 8931 286
rect 8959 258 9017 286
rect 9045 258 9103 286
rect 9131 258 9170 286
rect 8800 200 9170 258
rect 8800 172 8845 200
rect 8873 172 8931 200
rect 8959 172 9017 200
rect 9045 172 9103 200
rect 9131 172 9170 200
rect 8800 114 9170 172
rect 8800 86 8845 114
rect 8873 86 8931 114
rect 8959 86 9017 114
rect 9045 86 9103 114
rect 9131 86 9170 114
rect 8800 47 9170 86
rect 9198 372 9568 417
rect 9198 344 9243 372
rect 9271 344 9329 372
rect 9357 344 9415 372
rect 9443 344 9501 372
rect 9529 344 9568 372
rect 9198 286 9568 344
rect 9198 258 9243 286
rect 9271 258 9329 286
rect 9357 258 9415 286
rect 9443 258 9501 286
rect 9529 258 9568 286
rect 9198 236 9568 258
rect 9596 372 9966 417
rect 9596 344 9641 372
rect 9669 344 9727 372
rect 9755 344 9813 372
rect 9841 344 9899 372
rect 9927 344 9966 372
rect 9596 286 9966 344
rect 9596 258 9641 286
rect 9669 258 9727 286
rect 9755 258 9813 286
rect 9841 258 9899 286
rect 9927 258 9966 286
rect 9596 236 9966 258
rect 9198 209 9966 236
rect 9198 200 9568 209
rect 9198 172 9243 200
rect 9271 172 9329 200
rect 9357 172 9415 200
rect 9443 172 9501 200
rect 9529 172 9568 200
rect 9198 114 9568 172
rect 9198 86 9243 114
rect 9271 86 9329 114
rect 9357 86 9415 114
rect 9443 86 9501 114
rect 9529 86 9568 114
rect 9198 47 9568 86
rect 9596 200 9966 209
rect 9596 172 9641 200
rect 9669 172 9727 200
rect 9755 172 9813 200
rect 9841 172 9899 200
rect 9927 172 9966 200
rect 9596 114 9966 172
rect 9596 86 9641 114
rect 9669 86 9727 114
rect 9755 86 9813 114
rect 9841 86 9899 114
rect 9927 86 9966 114
rect 9596 47 9966 86
<< via2 >>
rect 89 1646 117 1674
rect 175 1646 203 1674
rect 261 1646 289 1674
rect 347 1646 375 1674
rect 89 1560 117 1588
rect 175 1560 203 1588
rect 261 1560 289 1588
rect 347 1560 375 1588
rect 487 1646 515 1674
rect 573 1646 601 1674
rect 659 1646 687 1674
rect 745 1646 773 1674
rect 487 1560 515 1588
rect 573 1560 601 1588
rect 659 1560 687 1588
rect 745 1560 773 1588
rect 885 1646 913 1674
rect 971 1646 999 1674
rect 1057 1646 1085 1674
rect 1143 1646 1171 1674
rect 885 1560 913 1588
rect 971 1560 999 1588
rect 1057 1560 1085 1588
rect 1143 1560 1171 1588
rect 1283 1646 1311 1674
rect 1369 1646 1397 1674
rect 1455 1646 1483 1674
rect 1541 1646 1569 1674
rect 1283 1560 1311 1588
rect 1369 1560 1397 1588
rect 1455 1560 1483 1588
rect 1541 1560 1569 1588
rect 1681 1646 1709 1674
rect 1767 1646 1795 1674
rect 1853 1646 1881 1674
rect 1939 1646 1967 1674
rect 1681 1560 1709 1588
rect 1767 1560 1795 1588
rect 1853 1560 1881 1588
rect 1939 1560 1967 1588
rect 2079 1646 2107 1674
rect 2165 1646 2193 1674
rect 2251 1646 2279 1674
rect 2337 1646 2365 1674
rect 2079 1560 2107 1588
rect 2165 1560 2193 1588
rect 2251 1560 2279 1588
rect 2337 1560 2365 1588
rect 2477 1646 2505 1674
rect 2563 1646 2591 1674
rect 2649 1646 2677 1674
rect 2735 1646 2763 1674
rect 2477 1560 2505 1588
rect 2563 1560 2591 1588
rect 2649 1560 2677 1588
rect 2735 1560 2763 1588
rect 2875 1646 2903 1674
rect 2961 1646 2989 1674
rect 3047 1646 3075 1674
rect 3133 1646 3161 1674
rect 2875 1560 2903 1588
rect 2961 1560 2989 1588
rect 3047 1560 3075 1588
rect 3133 1560 3161 1588
rect 3273 1646 3301 1674
rect 3359 1646 3387 1674
rect 3445 1646 3473 1674
rect 3531 1646 3559 1674
rect 3273 1560 3301 1588
rect 3359 1560 3387 1588
rect 3445 1560 3473 1588
rect 3531 1560 3559 1588
rect 3671 1646 3699 1674
rect 3757 1646 3785 1674
rect 3843 1646 3871 1674
rect 3929 1646 3957 1674
rect 3671 1560 3699 1588
rect 3757 1560 3785 1588
rect 3843 1560 3871 1588
rect 3929 1560 3957 1588
rect 4069 1646 4097 1674
rect 4155 1646 4183 1674
rect 4241 1646 4269 1674
rect 4327 1646 4355 1674
rect 4069 1560 4097 1588
rect 4155 1560 4183 1588
rect 4241 1560 4269 1588
rect 4327 1560 4355 1588
rect 4467 1646 4495 1674
rect 4553 1646 4581 1674
rect 4639 1646 4667 1674
rect 4725 1646 4753 1674
rect 4467 1560 4495 1588
rect 4553 1560 4581 1588
rect 4639 1560 4667 1588
rect 4725 1560 4753 1588
rect 4865 1646 4893 1674
rect 4951 1646 4979 1674
rect 5037 1646 5065 1674
rect 5123 1646 5151 1674
rect 4865 1560 4893 1588
rect 4951 1560 4979 1588
rect 5037 1560 5065 1588
rect 5123 1560 5151 1588
rect 5263 1646 5291 1674
rect 5349 1646 5377 1674
rect 5435 1646 5463 1674
rect 5521 1646 5549 1674
rect 5263 1560 5291 1588
rect 5349 1560 5377 1588
rect 5435 1560 5463 1588
rect 5521 1560 5549 1588
rect 5661 1646 5689 1674
rect 5747 1646 5775 1674
rect 5833 1646 5861 1674
rect 5919 1646 5947 1674
rect 5661 1560 5689 1588
rect 5747 1560 5775 1588
rect 5833 1560 5861 1588
rect 5919 1560 5947 1588
rect 6059 1646 6087 1674
rect 6145 1646 6173 1674
rect 6231 1646 6259 1674
rect 6317 1646 6345 1674
rect 6059 1560 6087 1588
rect 6145 1560 6173 1588
rect 6231 1560 6259 1588
rect 6317 1560 6345 1588
rect 6457 1646 6485 1674
rect 6543 1646 6571 1674
rect 6629 1646 6657 1674
rect 6715 1646 6743 1674
rect 6457 1560 6485 1588
rect 6543 1560 6571 1588
rect 6629 1560 6657 1588
rect 6715 1560 6743 1588
rect 6855 1646 6883 1674
rect 6941 1646 6969 1674
rect 7027 1646 7055 1674
rect 7113 1646 7141 1674
rect 6855 1560 6883 1588
rect 6941 1560 6969 1588
rect 7027 1560 7055 1588
rect 7113 1560 7141 1588
rect 7253 1646 7281 1674
rect 7339 1646 7367 1674
rect 7425 1646 7453 1674
rect 7511 1646 7539 1674
rect 7253 1560 7281 1588
rect 7339 1560 7367 1588
rect 7425 1560 7453 1588
rect 7511 1560 7539 1588
rect 7651 1646 7679 1674
rect 7737 1646 7765 1674
rect 7823 1646 7851 1674
rect 7909 1646 7937 1674
rect 7651 1560 7679 1588
rect 7737 1560 7765 1588
rect 7823 1560 7851 1588
rect 7909 1560 7937 1588
rect 8049 1646 8077 1674
rect 8135 1646 8163 1674
rect 8221 1646 8249 1674
rect 8307 1646 8335 1674
rect 8049 1560 8077 1588
rect 8135 1560 8163 1588
rect 8221 1560 8249 1588
rect 8307 1560 8335 1588
rect 8447 1646 8475 1674
rect 8533 1646 8561 1674
rect 8619 1646 8647 1674
rect 8705 1646 8733 1674
rect 8447 1560 8475 1588
rect 8533 1560 8561 1588
rect 8619 1560 8647 1588
rect 8705 1560 8733 1588
rect 8845 1646 8873 1674
rect 8931 1646 8959 1674
rect 9017 1646 9045 1674
rect 9103 1646 9131 1674
rect 8845 1560 8873 1588
rect 8931 1560 8959 1588
rect 9017 1560 9045 1588
rect 9103 1560 9131 1588
rect 9243 1646 9271 1674
rect 9329 1646 9357 1674
rect 9415 1646 9443 1674
rect 9501 1646 9529 1674
rect 9243 1560 9271 1588
rect 9329 1560 9357 1588
rect 9415 1560 9443 1588
rect 9501 1560 9529 1588
rect 9641 1646 9669 1674
rect 9727 1646 9755 1674
rect 9813 1646 9841 1674
rect 9899 1646 9927 1674
rect 9641 1560 9669 1588
rect 9727 1560 9755 1588
rect 9813 1560 9841 1588
rect 9899 1560 9927 1588
rect 89 1474 117 1502
rect 175 1474 203 1502
rect 261 1474 289 1502
rect 347 1474 375 1502
rect 89 1388 117 1416
rect 175 1388 203 1416
rect 261 1388 289 1416
rect 347 1388 375 1416
rect 487 1474 515 1502
rect 573 1474 601 1502
rect 659 1474 687 1502
rect 745 1474 773 1502
rect 487 1388 515 1416
rect 573 1388 601 1416
rect 659 1388 687 1416
rect 745 1388 773 1416
rect 885 1474 913 1502
rect 971 1474 999 1502
rect 1057 1474 1085 1502
rect 1143 1474 1171 1502
rect 885 1388 913 1416
rect 971 1388 999 1416
rect 1057 1388 1085 1416
rect 1143 1388 1171 1416
rect 1283 1474 1311 1502
rect 1369 1474 1397 1502
rect 1455 1474 1483 1502
rect 1541 1474 1569 1502
rect 1283 1388 1311 1416
rect 1369 1388 1397 1416
rect 1455 1388 1483 1416
rect 1541 1388 1569 1416
rect 1681 1474 1709 1502
rect 1767 1474 1795 1502
rect 1853 1474 1881 1502
rect 1939 1474 1967 1502
rect 1681 1388 1709 1416
rect 1767 1388 1795 1416
rect 1853 1388 1881 1416
rect 1939 1388 1967 1416
rect 2079 1474 2107 1502
rect 2165 1474 2193 1502
rect 2251 1474 2279 1502
rect 2337 1474 2365 1502
rect 2079 1388 2107 1416
rect 2165 1388 2193 1416
rect 2251 1388 2279 1416
rect 2337 1388 2365 1416
rect 2477 1474 2505 1502
rect 2563 1474 2591 1502
rect 2649 1474 2677 1502
rect 2735 1474 2763 1502
rect 2477 1388 2505 1416
rect 2563 1388 2591 1416
rect 2649 1388 2677 1416
rect 2735 1388 2763 1416
rect 2875 1474 2903 1502
rect 2961 1474 2989 1502
rect 3047 1474 3075 1502
rect 3133 1474 3161 1502
rect 2875 1388 2903 1416
rect 2961 1388 2989 1416
rect 3047 1388 3075 1416
rect 3133 1388 3161 1416
rect 3273 1474 3301 1502
rect 3359 1474 3387 1502
rect 3445 1474 3473 1502
rect 3531 1474 3559 1502
rect 3273 1388 3301 1416
rect 3359 1388 3387 1416
rect 3445 1388 3473 1416
rect 3531 1388 3559 1416
rect 3671 1474 3699 1502
rect 3757 1474 3785 1502
rect 3843 1474 3871 1502
rect 3929 1474 3957 1502
rect 3671 1388 3699 1416
rect 3757 1388 3785 1416
rect 3843 1388 3871 1416
rect 3929 1388 3957 1416
rect 4069 1474 4097 1502
rect 4155 1474 4183 1502
rect 4241 1474 4269 1502
rect 4327 1474 4355 1502
rect 4069 1388 4097 1416
rect 4155 1388 4183 1416
rect 4241 1388 4269 1416
rect 4327 1388 4355 1416
rect 4467 1474 4495 1502
rect 4553 1474 4581 1502
rect 4639 1474 4667 1502
rect 4725 1474 4753 1502
rect 4467 1388 4495 1416
rect 4553 1388 4581 1416
rect 4639 1388 4667 1416
rect 4725 1388 4753 1416
rect 4865 1474 4893 1502
rect 4951 1474 4979 1502
rect 5037 1474 5065 1502
rect 5123 1474 5151 1502
rect 4865 1388 4893 1416
rect 4951 1388 4979 1416
rect 5037 1388 5065 1416
rect 5123 1388 5151 1416
rect 5263 1474 5291 1502
rect 5349 1474 5377 1502
rect 5435 1474 5463 1502
rect 5521 1474 5549 1502
rect 5263 1388 5291 1416
rect 5349 1388 5377 1416
rect 5435 1388 5463 1416
rect 5521 1388 5549 1416
rect 5661 1474 5689 1502
rect 5747 1474 5775 1502
rect 5833 1474 5861 1502
rect 5919 1474 5947 1502
rect 5661 1388 5689 1416
rect 5747 1388 5775 1416
rect 5833 1388 5861 1416
rect 5919 1388 5947 1416
rect 6059 1474 6087 1502
rect 6145 1474 6173 1502
rect 6231 1474 6259 1502
rect 6317 1474 6345 1502
rect 6059 1388 6087 1416
rect 6145 1388 6173 1416
rect 6231 1388 6259 1416
rect 6317 1388 6345 1416
rect 6457 1474 6485 1502
rect 6543 1474 6571 1502
rect 6629 1474 6657 1502
rect 6715 1474 6743 1502
rect 6457 1388 6485 1416
rect 6543 1388 6571 1416
rect 6629 1388 6657 1416
rect 6715 1388 6743 1416
rect 6855 1474 6883 1502
rect 6941 1474 6969 1502
rect 7027 1474 7055 1502
rect 7113 1474 7141 1502
rect 6855 1388 6883 1416
rect 6941 1388 6969 1416
rect 7027 1388 7055 1416
rect 7113 1388 7141 1416
rect 7253 1474 7281 1502
rect 7339 1474 7367 1502
rect 7425 1474 7453 1502
rect 7511 1474 7539 1502
rect 7253 1388 7281 1416
rect 7339 1388 7367 1416
rect 7425 1388 7453 1416
rect 7511 1388 7539 1416
rect 7651 1474 7679 1502
rect 7737 1474 7765 1502
rect 7823 1474 7851 1502
rect 7909 1474 7937 1502
rect 7651 1388 7679 1416
rect 7737 1388 7765 1416
rect 7823 1388 7851 1416
rect 7909 1388 7937 1416
rect 8049 1474 8077 1502
rect 8135 1474 8163 1502
rect 8221 1474 8249 1502
rect 8307 1474 8335 1502
rect 8049 1388 8077 1416
rect 8135 1388 8163 1416
rect 8221 1388 8249 1416
rect 8307 1388 8335 1416
rect 8447 1474 8475 1502
rect 8533 1474 8561 1502
rect 8619 1474 8647 1502
rect 8705 1474 8733 1502
rect 8447 1388 8475 1416
rect 8533 1388 8561 1416
rect 8619 1388 8647 1416
rect 8705 1388 8733 1416
rect 8845 1474 8873 1502
rect 8931 1474 8959 1502
rect 9017 1474 9045 1502
rect 9103 1474 9131 1502
rect 8845 1388 8873 1416
rect 8931 1388 8959 1416
rect 9017 1388 9045 1416
rect 9103 1388 9131 1416
rect 9243 1474 9271 1502
rect 9329 1474 9357 1502
rect 9415 1474 9443 1502
rect 9501 1474 9529 1502
rect 9243 1388 9271 1416
rect 9329 1388 9357 1416
rect 9415 1388 9443 1416
rect 9501 1388 9529 1416
rect 9641 1474 9669 1502
rect 9727 1474 9755 1502
rect 9813 1474 9841 1502
rect 9899 1474 9927 1502
rect 9641 1388 9669 1416
rect 9727 1388 9755 1416
rect 9813 1388 9841 1416
rect 9899 1388 9927 1416
rect 89 1212 117 1240
rect 175 1212 203 1240
rect 261 1212 289 1240
rect 347 1212 375 1240
rect 89 1126 117 1154
rect 175 1126 203 1154
rect 261 1126 289 1154
rect 347 1126 375 1154
rect 89 1040 117 1068
rect 175 1040 203 1068
rect 261 1040 289 1068
rect 347 1040 375 1068
rect 89 954 117 982
rect 175 954 203 982
rect 261 954 289 982
rect 347 954 375 982
rect 487 1212 515 1240
rect 573 1212 601 1240
rect 659 1212 687 1240
rect 745 1212 773 1240
rect 487 1126 515 1154
rect 573 1126 601 1154
rect 659 1126 687 1154
rect 745 1126 773 1154
rect 885 1212 913 1240
rect 971 1212 999 1240
rect 1057 1212 1085 1240
rect 1143 1212 1171 1240
rect 885 1126 913 1154
rect 971 1126 999 1154
rect 1057 1126 1085 1154
rect 1143 1126 1171 1154
rect 1283 1212 1311 1240
rect 1369 1212 1397 1240
rect 1455 1212 1483 1240
rect 1541 1212 1569 1240
rect 1283 1126 1311 1154
rect 1369 1126 1397 1154
rect 1455 1126 1483 1154
rect 1541 1126 1569 1154
rect 487 1040 515 1068
rect 573 1040 601 1068
rect 659 1040 687 1068
rect 745 1040 773 1068
rect 487 954 515 982
rect 573 954 601 982
rect 659 954 687 982
rect 745 954 773 982
rect 885 1040 913 1068
rect 971 1040 999 1068
rect 1057 1040 1085 1068
rect 1143 1040 1171 1068
rect 885 954 913 982
rect 971 954 999 982
rect 1057 954 1085 982
rect 1143 954 1171 982
rect 1283 1040 1311 1068
rect 1369 1040 1397 1068
rect 1455 1040 1483 1068
rect 1541 1040 1569 1068
rect 1283 954 1311 982
rect 1369 954 1397 982
rect 1455 954 1483 982
rect 1541 954 1569 982
rect 1681 1212 1709 1240
rect 1767 1212 1795 1240
rect 1853 1212 1881 1240
rect 1939 1212 1967 1240
rect 1681 1126 1709 1154
rect 1767 1126 1795 1154
rect 1853 1126 1881 1154
rect 1939 1126 1967 1154
rect 1681 1040 1709 1068
rect 1767 1040 1795 1068
rect 1853 1040 1881 1068
rect 1939 1040 1967 1068
rect 1681 954 1709 982
rect 1767 954 1795 982
rect 1853 954 1881 982
rect 1939 954 1967 982
rect 2079 1212 2107 1240
rect 2165 1212 2193 1240
rect 2251 1212 2279 1240
rect 2337 1212 2365 1240
rect 2079 1126 2107 1154
rect 2165 1126 2193 1154
rect 2251 1126 2279 1154
rect 2337 1126 2365 1154
rect 2079 1040 2107 1068
rect 2165 1040 2193 1068
rect 2251 1040 2279 1068
rect 2337 1040 2365 1068
rect 2079 954 2107 982
rect 2165 954 2193 982
rect 2251 954 2279 982
rect 2337 954 2365 982
rect 2477 1212 2505 1240
rect 2563 1212 2591 1240
rect 2649 1212 2677 1240
rect 2735 1212 2763 1240
rect 2477 1126 2505 1154
rect 2563 1126 2591 1154
rect 2649 1126 2677 1154
rect 2735 1126 2763 1154
rect 2875 1212 2903 1240
rect 2961 1212 2989 1240
rect 3047 1212 3075 1240
rect 3133 1212 3161 1240
rect 2875 1126 2903 1154
rect 2961 1126 2989 1154
rect 3047 1126 3075 1154
rect 3133 1126 3161 1154
rect 3273 1212 3301 1240
rect 3359 1212 3387 1240
rect 3445 1212 3473 1240
rect 3531 1212 3559 1240
rect 3273 1126 3301 1154
rect 3359 1126 3387 1154
rect 3445 1126 3473 1154
rect 3531 1126 3559 1154
rect 2477 1040 2505 1068
rect 2563 1040 2591 1068
rect 2649 1040 2677 1068
rect 2735 1040 2763 1068
rect 2477 954 2505 982
rect 2563 954 2591 982
rect 2649 954 2677 982
rect 2735 954 2763 982
rect 2875 1040 2903 1068
rect 2961 1040 2989 1068
rect 3047 1040 3075 1068
rect 3133 1040 3161 1068
rect 2875 954 2903 982
rect 2961 954 2989 982
rect 3047 954 3075 982
rect 3133 954 3161 982
rect 3273 1040 3301 1068
rect 3359 1040 3387 1068
rect 3445 1040 3473 1068
rect 3531 1040 3559 1068
rect 3273 954 3301 982
rect 3359 954 3387 982
rect 3445 954 3473 982
rect 3531 954 3559 982
rect 3671 1212 3699 1240
rect 3757 1212 3785 1240
rect 3843 1212 3871 1240
rect 3929 1212 3957 1240
rect 3671 1126 3699 1154
rect 3757 1126 3785 1154
rect 3843 1126 3871 1154
rect 3929 1126 3957 1154
rect 3671 1040 3699 1068
rect 3757 1040 3785 1068
rect 3843 1040 3871 1068
rect 3929 1040 3957 1068
rect 3671 954 3699 982
rect 3757 954 3785 982
rect 3843 954 3871 982
rect 3929 954 3957 982
rect 4069 1212 4097 1240
rect 4155 1212 4183 1240
rect 4241 1212 4269 1240
rect 4327 1212 4355 1240
rect 4069 1126 4097 1154
rect 4155 1126 4183 1154
rect 4241 1126 4269 1154
rect 4327 1126 4355 1154
rect 4069 1040 4097 1068
rect 4155 1040 4183 1068
rect 4241 1040 4269 1068
rect 4327 1040 4355 1068
rect 4069 954 4097 982
rect 4155 954 4183 982
rect 4241 954 4269 982
rect 4327 954 4355 982
rect 4467 1212 4495 1240
rect 4553 1212 4581 1240
rect 4639 1212 4667 1240
rect 4725 1212 4753 1240
rect 4467 1126 4495 1154
rect 4553 1126 4581 1154
rect 4639 1126 4667 1154
rect 4725 1126 4753 1154
rect 4865 1212 4893 1240
rect 4951 1212 4979 1240
rect 5037 1212 5065 1240
rect 5123 1212 5151 1240
rect 4865 1126 4893 1154
rect 4951 1126 4979 1154
rect 5037 1126 5065 1154
rect 5123 1126 5151 1154
rect 5263 1212 5291 1240
rect 5349 1212 5377 1240
rect 5435 1212 5463 1240
rect 5521 1212 5549 1240
rect 5263 1126 5291 1154
rect 5349 1126 5377 1154
rect 5435 1126 5463 1154
rect 5521 1126 5549 1154
rect 4467 1040 4495 1068
rect 4553 1040 4581 1068
rect 4639 1040 4667 1068
rect 4725 1040 4753 1068
rect 4467 954 4495 982
rect 4553 954 4581 982
rect 4639 954 4667 982
rect 4725 954 4753 982
rect 4865 1040 4893 1068
rect 4951 1040 4979 1068
rect 5037 1040 5065 1068
rect 5123 1040 5151 1068
rect 4865 954 4893 982
rect 4951 954 4979 982
rect 5037 954 5065 982
rect 5123 954 5151 982
rect 5263 1040 5291 1068
rect 5349 1040 5377 1068
rect 5435 1040 5463 1068
rect 5521 1040 5549 1068
rect 5263 954 5291 982
rect 5349 954 5377 982
rect 5435 954 5463 982
rect 5521 954 5549 982
rect 5661 1212 5689 1240
rect 5747 1212 5775 1240
rect 5833 1212 5861 1240
rect 5919 1212 5947 1240
rect 5661 1126 5689 1154
rect 5747 1126 5775 1154
rect 5833 1126 5861 1154
rect 5919 1126 5947 1154
rect 5661 1040 5689 1068
rect 5747 1040 5775 1068
rect 5833 1040 5861 1068
rect 5919 1040 5947 1068
rect 5661 954 5689 982
rect 5747 954 5775 982
rect 5833 954 5861 982
rect 5919 954 5947 982
rect 6059 1212 6087 1240
rect 6145 1212 6173 1240
rect 6231 1212 6259 1240
rect 6317 1212 6345 1240
rect 6059 1126 6087 1154
rect 6145 1126 6173 1154
rect 6231 1126 6259 1154
rect 6317 1126 6345 1154
rect 6059 1040 6087 1068
rect 6145 1040 6173 1068
rect 6231 1040 6259 1068
rect 6317 1040 6345 1068
rect 6059 954 6087 982
rect 6145 954 6173 982
rect 6231 954 6259 982
rect 6317 954 6345 982
rect 6457 1212 6485 1240
rect 6543 1212 6571 1240
rect 6629 1212 6657 1240
rect 6715 1212 6743 1240
rect 6457 1126 6485 1154
rect 6543 1126 6571 1154
rect 6629 1126 6657 1154
rect 6715 1126 6743 1154
rect 6855 1212 6883 1240
rect 6941 1212 6969 1240
rect 7027 1212 7055 1240
rect 7113 1212 7141 1240
rect 6855 1126 6883 1154
rect 6941 1126 6969 1154
rect 7027 1126 7055 1154
rect 7113 1126 7141 1154
rect 7253 1212 7281 1240
rect 7339 1212 7367 1240
rect 7425 1212 7453 1240
rect 7511 1212 7539 1240
rect 7253 1126 7281 1154
rect 7339 1126 7367 1154
rect 7425 1126 7453 1154
rect 7511 1126 7539 1154
rect 6457 1040 6485 1068
rect 6543 1040 6571 1068
rect 6629 1040 6657 1068
rect 6715 1040 6743 1068
rect 6457 954 6485 982
rect 6543 954 6571 982
rect 6629 954 6657 982
rect 6715 954 6743 982
rect 6855 1040 6883 1068
rect 6941 1040 6969 1068
rect 7027 1040 7055 1068
rect 7113 1040 7141 1068
rect 6855 954 6883 982
rect 6941 954 6969 982
rect 7027 954 7055 982
rect 7113 954 7141 982
rect 7253 1040 7281 1068
rect 7339 1040 7367 1068
rect 7425 1040 7453 1068
rect 7511 1040 7539 1068
rect 7253 954 7281 982
rect 7339 954 7367 982
rect 7425 954 7453 982
rect 7511 954 7539 982
rect 7651 1212 7679 1240
rect 7737 1212 7765 1240
rect 7823 1212 7851 1240
rect 7909 1212 7937 1240
rect 7651 1126 7679 1154
rect 7737 1126 7765 1154
rect 7823 1126 7851 1154
rect 7909 1126 7937 1154
rect 7651 1040 7679 1068
rect 7737 1040 7765 1068
rect 7823 1040 7851 1068
rect 7909 1040 7937 1068
rect 7651 954 7679 982
rect 7737 954 7765 982
rect 7823 954 7851 982
rect 7909 954 7937 982
rect 8049 1212 8077 1240
rect 8135 1212 8163 1240
rect 8221 1212 8249 1240
rect 8307 1212 8335 1240
rect 8049 1126 8077 1154
rect 8135 1126 8163 1154
rect 8221 1126 8249 1154
rect 8307 1126 8335 1154
rect 8049 1040 8077 1068
rect 8135 1040 8163 1068
rect 8221 1040 8249 1068
rect 8307 1040 8335 1068
rect 8049 954 8077 982
rect 8135 954 8163 982
rect 8221 954 8249 982
rect 8307 954 8335 982
rect 8447 1212 8475 1240
rect 8533 1212 8561 1240
rect 8619 1212 8647 1240
rect 8705 1212 8733 1240
rect 8447 1126 8475 1154
rect 8533 1126 8561 1154
rect 8619 1126 8647 1154
rect 8705 1126 8733 1154
rect 8845 1212 8873 1240
rect 8931 1212 8959 1240
rect 9017 1212 9045 1240
rect 9103 1212 9131 1240
rect 8845 1126 8873 1154
rect 8931 1126 8959 1154
rect 9017 1126 9045 1154
rect 9103 1126 9131 1154
rect 9243 1212 9271 1240
rect 9329 1212 9357 1240
rect 9415 1212 9443 1240
rect 9501 1212 9529 1240
rect 9243 1126 9271 1154
rect 9329 1126 9357 1154
rect 9415 1126 9443 1154
rect 9501 1126 9529 1154
rect 8447 1040 8475 1068
rect 8533 1040 8561 1068
rect 8619 1040 8647 1068
rect 8705 1040 8733 1068
rect 8447 954 8475 982
rect 8533 954 8561 982
rect 8619 954 8647 982
rect 8705 954 8733 982
rect 8845 1040 8873 1068
rect 8931 1040 8959 1068
rect 9017 1040 9045 1068
rect 9103 1040 9131 1068
rect 8845 954 8873 982
rect 8931 954 8959 982
rect 9017 954 9045 982
rect 9103 954 9131 982
rect 9243 1040 9271 1068
rect 9329 1040 9357 1068
rect 9415 1040 9443 1068
rect 9501 1040 9529 1068
rect 9243 954 9271 982
rect 9329 954 9357 982
rect 9415 954 9443 982
rect 9501 954 9529 982
rect 9641 1212 9669 1240
rect 9727 1212 9755 1240
rect 9813 1212 9841 1240
rect 9899 1212 9927 1240
rect 9641 1126 9669 1154
rect 9727 1126 9755 1154
rect 9813 1126 9841 1154
rect 9899 1126 9927 1154
rect 9641 1040 9669 1068
rect 9727 1040 9755 1068
rect 9813 1040 9841 1068
rect 9899 1040 9927 1068
rect 9641 954 9669 982
rect 9727 954 9755 982
rect 9813 954 9841 982
rect 9899 954 9927 982
rect 89 778 117 806
rect 175 778 203 806
rect 261 778 289 806
rect 347 778 375 806
rect 89 692 117 720
rect 175 692 203 720
rect 261 692 289 720
rect 347 692 375 720
rect 89 606 117 634
rect 175 606 203 634
rect 261 606 289 634
rect 347 606 375 634
rect 89 520 117 548
rect 175 520 203 548
rect 261 520 289 548
rect 347 520 375 548
rect 487 778 515 806
rect 573 778 601 806
rect 659 778 687 806
rect 745 778 773 806
rect 487 692 515 720
rect 573 692 601 720
rect 659 692 687 720
rect 745 692 773 720
rect 885 778 913 806
rect 971 778 999 806
rect 1057 778 1085 806
rect 1143 778 1171 806
rect 885 692 913 720
rect 971 692 999 720
rect 1057 692 1085 720
rect 1143 692 1171 720
rect 1283 778 1311 806
rect 1369 778 1397 806
rect 1455 778 1483 806
rect 1541 778 1569 806
rect 1283 692 1311 720
rect 1369 692 1397 720
rect 1455 692 1483 720
rect 1541 692 1569 720
rect 487 606 515 634
rect 573 606 601 634
rect 659 606 687 634
rect 745 606 773 634
rect 487 520 515 548
rect 573 520 601 548
rect 659 520 687 548
rect 745 520 773 548
rect 885 606 913 634
rect 971 606 999 634
rect 1057 606 1085 634
rect 1143 606 1171 634
rect 885 520 913 548
rect 971 520 999 548
rect 1057 520 1085 548
rect 1143 520 1171 548
rect 1283 606 1311 634
rect 1369 606 1397 634
rect 1455 606 1483 634
rect 1541 606 1569 634
rect 1283 520 1311 548
rect 1369 520 1397 548
rect 1455 520 1483 548
rect 1541 520 1569 548
rect 1681 778 1709 806
rect 1767 778 1795 806
rect 1853 778 1881 806
rect 1939 778 1967 806
rect 1681 692 1709 720
rect 1767 692 1795 720
rect 1853 692 1881 720
rect 1939 692 1967 720
rect 1681 606 1709 634
rect 1767 606 1795 634
rect 1853 606 1881 634
rect 1939 606 1967 634
rect 1681 520 1709 548
rect 1767 520 1795 548
rect 1853 520 1881 548
rect 1939 520 1967 548
rect 2079 778 2107 806
rect 2165 778 2193 806
rect 2251 778 2279 806
rect 2337 778 2365 806
rect 2079 692 2107 720
rect 2165 692 2193 720
rect 2251 692 2279 720
rect 2337 692 2365 720
rect 2079 606 2107 634
rect 2165 606 2193 634
rect 2251 606 2279 634
rect 2337 606 2365 634
rect 2079 520 2107 548
rect 2165 520 2193 548
rect 2251 520 2279 548
rect 2337 520 2365 548
rect 2477 778 2505 806
rect 2563 778 2591 806
rect 2649 778 2677 806
rect 2735 778 2763 806
rect 2477 692 2505 720
rect 2563 692 2591 720
rect 2649 692 2677 720
rect 2735 692 2763 720
rect 2875 778 2903 806
rect 2961 778 2989 806
rect 3047 778 3075 806
rect 3133 778 3161 806
rect 2875 692 2903 720
rect 2961 692 2989 720
rect 3047 692 3075 720
rect 3133 692 3161 720
rect 3273 778 3301 806
rect 3359 778 3387 806
rect 3445 778 3473 806
rect 3531 778 3559 806
rect 3273 692 3301 720
rect 3359 692 3387 720
rect 3445 692 3473 720
rect 3531 692 3559 720
rect 2477 606 2505 634
rect 2563 606 2591 634
rect 2649 606 2677 634
rect 2735 606 2763 634
rect 2477 520 2505 548
rect 2563 520 2591 548
rect 2649 520 2677 548
rect 2735 520 2763 548
rect 2875 606 2903 634
rect 2961 606 2989 634
rect 3047 606 3075 634
rect 3133 606 3161 634
rect 2875 520 2903 548
rect 2961 520 2989 548
rect 3047 520 3075 548
rect 3133 520 3161 548
rect 3273 606 3301 634
rect 3359 606 3387 634
rect 3445 606 3473 634
rect 3531 606 3559 634
rect 3273 520 3301 548
rect 3359 520 3387 548
rect 3445 520 3473 548
rect 3531 520 3559 548
rect 3671 778 3699 806
rect 3757 778 3785 806
rect 3843 778 3871 806
rect 3929 778 3957 806
rect 3671 692 3699 720
rect 3757 692 3785 720
rect 3843 692 3871 720
rect 3929 692 3957 720
rect 3671 606 3699 634
rect 3757 606 3785 634
rect 3843 606 3871 634
rect 3929 606 3957 634
rect 3671 520 3699 548
rect 3757 520 3785 548
rect 3843 520 3871 548
rect 3929 520 3957 548
rect 4069 778 4097 806
rect 4155 778 4183 806
rect 4241 778 4269 806
rect 4327 778 4355 806
rect 4069 692 4097 720
rect 4155 692 4183 720
rect 4241 692 4269 720
rect 4327 692 4355 720
rect 4069 606 4097 634
rect 4155 606 4183 634
rect 4241 606 4269 634
rect 4327 606 4355 634
rect 4069 520 4097 548
rect 4155 520 4183 548
rect 4241 520 4269 548
rect 4327 520 4355 548
rect 4467 778 4495 806
rect 4553 778 4581 806
rect 4639 778 4667 806
rect 4725 778 4753 806
rect 4467 692 4495 720
rect 4553 692 4581 720
rect 4639 692 4667 720
rect 4725 692 4753 720
rect 4865 778 4893 806
rect 4951 778 4979 806
rect 5037 778 5065 806
rect 5123 778 5151 806
rect 4865 692 4893 720
rect 4951 692 4979 720
rect 5037 692 5065 720
rect 5123 692 5151 720
rect 5263 778 5291 806
rect 5349 778 5377 806
rect 5435 778 5463 806
rect 5521 778 5549 806
rect 5263 692 5291 720
rect 5349 692 5377 720
rect 5435 692 5463 720
rect 5521 692 5549 720
rect 4467 606 4495 634
rect 4553 606 4581 634
rect 4639 606 4667 634
rect 4725 606 4753 634
rect 4467 520 4495 548
rect 4553 520 4581 548
rect 4639 520 4667 548
rect 4725 520 4753 548
rect 4865 606 4893 634
rect 4951 606 4979 634
rect 5037 606 5065 634
rect 5123 606 5151 634
rect 4865 520 4893 548
rect 4951 520 4979 548
rect 5037 520 5065 548
rect 5123 520 5151 548
rect 5263 606 5291 634
rect 5349 606 5377 634
rect 5435 606 5463 634
rect 5521 606 5549 634
rect 5263 520 5291 548
rect 5349 520 5377 548
rect 5435 520 5463 548
rect 5521 520 5549 548
rect 5661 778 5689 806
rect 5747 778 5775 806
rect 5833 778 5861 806
rect 5919 778 5947 806
rect 5661 692 5689 720
rect 5747 692 5775 720
rect 5833 692 5861 720
rect 5919 692 5947 720
rect 5661 606 5689 634
rect 5747 606 5775 634
rect 5833 606 5861 634
rect 5919 606 5947 634
rect 5661 520 5689 548
rect 5747 520 5775 548
rect 5833 520 5861 548
rect 5919 520 5947 548
rect 6059 778 6087 806
rect 6145 778 6173 806
rect 6231 778 6259 806
rect 6317 778 6345 806
rect 6059 692 6087 720
rect 6145 692 6173 720
rect 6231 692 6259 720
rect 6317 692 6345 720
rect 6059 606 6087 634
rect 6145 606 6173 634
rect 6231 606 6259 634
rect 6317 606 6345 634
rect 6059 520 6087 548
rect 6145 520 6173 548
rect 6231 520 6259 548
rect 6317 520 6345 548
rect 6457 778 6485 806
rect 6543 778 6571 806
rect 6629 778 6657 806
rect 6715 778 6743 806
rect 6457 692 6485 720
rect 6543 692 6571 720
rect 6629 692 6657 720
rect 6715 692 6743 720
rect 6855 778 6883 806
rect 6941 778 6969 806
rect 7027 778 7055 806
rect 7113 778 7141 806
rect 6855 692 6883 720
rect 6941 692 6969 720
rect 7027 692 7055 720
rect 7113 692 7141 720
rect 7253 778 7281 806
rect 7339 778 7367 806
rect 7425 778 7453 806
rect 7511 778 7539 806
rect 7253 692 7281 720
rect 7339 692 7367 720
rect 7425 692 7453 720
rect 7511 692 7539 720
rect 6457 606 6485 634
rect 6543 606 6571 634
rect 6629 606 6657 634
rect 6715 606 6743 634
rect 6457 520 6485 548
rect 6543 520 6571 548
rect 6629 520 6657 548
rect 6715 520 6743 548
rect 6855 606 6883 634
rect 6941 606 6969 634
rect 7027 606 7055 634
rect 7113 606 7141 634
rect 6855 520 6883 548
rect 6941 520 6969 548
rect 7027 520 7055 548
rect 7113 520 7141 548
rect 7253 606 7281 634
rect 7339 606 7367 634
rect 7425 606 7453 634
rect 7511 606 7539 634
rect 7253 520 7281 548
rect 7339 520 7367 548
rect 7425 520 7453 548
rect 7511 520 7539 548
rect 7651 778 7679 806
rect 7737 778 7765 806
rect 7823 778 7851 806
rect 7909 778 7937 806
rect 7651 692 7679 720
rect 7737 692 7765 720
rect 7823 692 7851 720
rect 7909 692 7937 720
rect 7651 606 7679 634
rect 7737 606 7765 634
rect 7823 606 7851 634
rect 7909 606 7937 634
rect 7651 520 7679 548
rect 7737 520 7765 548
rect 7823 520 7851 548
rect 7909 520 7937 548
rect 8049 778 8077 806
rect 8135 778 8163 806
rect 8221 778 8249 806
rect 8307 778 8335 806
rect 8049 692 8077 720
rect 8135 692 8163 720
rect 8221 692 8249 720
rect 8307 692 8335 720
rect 8049 606 8077 634
rect 8135 606 8163 634
rect 8221 606 8249 634
rect 8307 606 8335 634
rect 8049 520 8077 548
rect 8135 520 8163 548
rect 8221 520 8249 548
rect 8307 520 8335 548
rect 8447 778 8475 806
rect 8533 778 8561 806
rect 8619 778 8647 806
rect 8705 778 8733 806
rect 8447 692 8475 720
rect 8533 692 8561 720
rect 8619 692 8647 720
rect 8705 692 8733 720
rect 8845 778 8873 806
rect 8931 778 8959 806
rect 9017 778 9045 806
rect 9103 778 9131 806
rect 8845 692 8873 720
rect 8931 692 8959 720
rect 9017 692 9045 720
rect 9103 692 9131 720
rect 9243 778 9271 806
rect 9329 778 9357 806
rect 9415 778 9443 806
rect 9501 778 9529 806
rect 9243 692 9271 720
rect 9329 692 9357 720
rect 9415 692 9443 720
rect 9501 692 9529 720
rect 8447 606 8475 634
rect 8533 606 8561 634
rect 8619 606 8647 634
rect 8705 606 8733 634
rect 8447 520 8475 548
rect 8533 520 8561 548
rect 8619 520 8647 548
rect 8705 520 8733 548
rect 8845 606 8873 634
rect 8931 606 8959 634
rect 9017 606 9045 634
rect 9103 606 9131 634
rect 8845 520 8873 548
rect 8931 520 8959 548
rect 9017 520 9045 548
rect 9103 520 9131 548
rect 9243 606 9271 634
rect 9329 606 9357 634
rect 9415 606 9443 634
rect 9501 606 9529 634
rect 9243 520 9271 548
rect 9329 520 9357 548
rect 9415 520 9443 548
rect 9501 520 9529 548
rect 9641 778 9669 806
rect 9727 778 9755 806
rect 9813 778 9841 806
rect 9899 778 9927 806
rect 9641 692 9669 720
rect 9727 692 9755 720
rect 9813 692 9841 720
rect 9899 692 9927 720
rect 9641 606 9669 634
rect 9727 606 9755 634
rect 9813 606 9841 634
rect 9899 606 9927 634
rect 9641 520 9669 548
rect 9727 520 9755 548
rect 9813 520 9841 548
rect 9899 520 9927 548
rect 89 344 117 372
rect 175 344 203 372
rect 261 344 289 372
rect 347 344 375 372
rect 89 258 117 286
rect 175 258 203 286
rect 261 258 289 286
rect 347 258 375 286
rect 487 344 515 372
rect 573 344 601 372
rect 659 344 687 372
rect 745 344 773 372
rect 487 258 515 286
rect 573 258 601 286
rect 659 258 687 286
rect 745 258 773 286
rect 885 344 913 372
rect 971 344 999 372
rect 1057 344 1085 372
rect 1143 344 1171 372
rect 885 258 913 286
rect 971 258 999 286
rect 1057 258 1085 286
rect 1143 258 1171 286
rect 1283 344 1311 372
rect 1369 344 1397 372
rect 1455 344 1483 372
rect 1541 344 1569 372
rect 1283 258 1311 286
rect 1369 258 1397 286
rect 1455 258 1483 286
rect 1541 258 1569 286
rect 1681 344 1709 372
rect 1767 344 1795 372
rect 1853 344 1881 372
rect 1939 344 1967 372
rect 1681 258 1709 286
rect 1767 258 1795 286
rect 1853 258 1881 286
rect 1939 258 1967 286
rect 2079 344 2107 372
rect 2165 344 2193 372
rect 2251 344 2279 372
rect 2337 344 2365 372
rect 2079 258 2107 286
rect 2165 258 2193 286
rect 2251 258 2279 286
rect 2337 258 2365 286
rect 2477 344 2505 372
rect 2563 344 2591 372
rect 2649 344 2677 372
rect 2735 344 2763 372
rect 2477 258 2505 286
rect 2563 258 2591 286
rect 2649 258 2677 286
rect 2735 258 2763 286
rect 89 172 117 200
rect 175 172 203 200
rect 261 172 289 200
rect 347 172 375 200
rect 89 86 117 114
rect 175 86 203 114
rect 261 86 289 114
rect 347 86 375 114
rect 487 172 515 200
rect 573 172 601 200
rect 659 172 687 200
rect 745 172 773 200
rect 487 86 515 114
rect 573 86 601 114
rect 659 86 687 114
rect 745 86 773 114
rect 885 172 913 200
rect 971 172 999 200
rect 1057 172 1085 200
rect 1143 172 1171 200
rect 885 86 913 114
rect 971 86 999 114
rect 1057 86 1085 114
rect 1143 86 1171 114
rect 1283 172 1311 200
rect 1369 172 1397 200
rect 1455 172 1483 200
rect 1541 172 1569 200
rect 1283 86 1311 114
rect 1369 86 1397 114
rect 1455 86 1483 114
rect 1541 86 1569 114
rect 1681 172 1709 200
rect 1767 172 1795 200
rect 1853 172 1881 200
rect 1939 172 1967 200
rect 1681 86 1709 114
rect 1767 86 1795 114
rect 1853 86 1881 114
rect 1939 86 1967 114
rect 2079 172 2107 200
rect 2165 172 2193 200
rect 2251 172 2279 200
rect 2337 172 2365 200
rect 2079 86 2107 114
rect 2165 86 2193 114
rect 2251 86 2279 114
rect 2337 86 2365 114
rect 2477 172 2505 200
rect 2563 172 2591 200
rect 2649 172 2677 200
rect 2735 172 2763 200
rect 2477 86 2505 114
rect 2563 86 2591 114
rect 2649 86 2677 114
rect 2735 86 2763 114
rect 2875 344 2903 372
rect 2961 344 2989 372
rect 3047 344 3075 372
rect 3133 344 3161 372
rect 2875 258 2903 286
rect 2961 258 2989 286
rect 3047 258 3075 286
rect 3133 258 3161 286
rect 2875 172 2903 200
rect 2961 172 2989 200
rect 3047 172 3075 200
rect 3133 172 3161 200
rect 2875 86 2903 114
rect 2961 86 2989 114
rect 3047 86 3075 114
rect 3133 86 3161 114
rect 3273 344 3301 372
rect 3359 344 3387 372
rect 3445 344 3473 372
rect 3531 344 3559 372
rect 3273 258 3301 286
rect 3359 258 3387 286
rect 3445 258 3473 286
rect 3531 258 3559 286
rect 3671 344 3699 372
rect 3757 344 3785 372
rect 3843 344 3871 372
rect 3929 344 3957 372
rect 3671 258 3699 286
rect 3757 258 3785 286
rect 3843 258 3871 286
rect 3929 258 3957 286
rect 4069 344 4097 372
rect 4155 344 4183 372
rect 4241 344 4269 372
rect 4327 344 4355 372
rect 4069 258 4097 286
rect 4155 258 4183 286
rect 4241 258 4269 286
rect 4327 258 4355 286
rect 4467 344 4495 372
rect 4553 344 4581 372
rect 4639 344 4667 372
rect 4725 344 4753 372
rect 4467 258 4495 286
rect 4553 258 4581 286
rect 4639 258 4667 286
rect 4725 258 4753 286
rect 3273 172 3301 200
rect 3359 172 3387 200
rect 3445 172 3473 200
rect 3531 172 3559 200
rect 3273 86 3301 114
rect 3359 86 3387 114
rect 3445 86 3473 114
rect 3531 86 3559 114
rect 3671 172 3699 200
rect 3757 172 3785 200
rect 3843 172 3871 200
rect 3929 172 3957 200
rect 3671 86 3699 114
rect 3757 86 3785 114
rect 3843 86 3871 114
rect 3929 86 3957 114
rect 4069 172 4097 200
rect 4155 172 4183 200
rect 4241 172 4269 200
rect 4327 172 4355 200
rect 4069 86 4097 114
rect 4155 86 4183 114
rect 4241 86 4269 114
rect 4327 86 4355 114
rect 4467 172 4495 200
rect 4553 172 4581 200
rect 4639 172 4667 200
rect 4725 172 4753 200
rect 4467 86 4495 114
rect 4553 86 4581 114
rect 4639 86 4667 114
rect 4725 86 4753 114
rect 4865 344 4893 372
rect 4951 344 4979 372
rect 5037 344 5065 372
rect 5123 344 5151 372
rect 4865 258 4893 286
rect 4951 258 4979 286
rect 5037 258 5065 286
rect 5123 258 5151 286
rect 4865 172 4893 200
rect 4951 172 4979 200
rect 5037 172 5065 200
rect 5123 172 5151 200
rect 4865 86 4893 114
rect 4951 86 4979 114
rect 5037 86 5065 114
rect 5123 86 5151 114
rect 5263 344 5291 372
rect 5349 344 5377 372
rect 5435 344 5463 372
rect 5521 344 5549 372
rect 5263 258 5291 286
rect 5349 258 5377 286
rect 5435 258 5463 286
rect 5521 258 5549 286
rect 5661 344 5689 372
rect 5747 344 5775 372
rect 5833 344 5861 372
rect 5919 344 5947 372
rect 5661 258 5689 286
rect 5747 258 5775 286
rect 5833 258 5861 286
rect 5919 258 5947 286
rect 6059 344 6087 372
rect 6145 344 6173 372
rect 6231 344 6259 372
rect 6317 344 6345 372
rect 6059 258 6087 286
rect 6145 258 6173 286
rect 6231 258 6259 286
rect 6317 258 6345 286
rect 6457 344 6485 372
rect 6543 344 6571 372
rect 6629 344 6657 372
rect 6715 344 6743 372
rect 6457 258 6485 286
rect 6543 258 6571 286
rect 6629 258 6657 286
rect 6715 258 6743 286
rect 5263 172 5291 200
rect 5349 172 5377 200
rect 5435 172 5463 200
rect 5521 172 5549 200
rect 5263 86 5291 114
rect 5349 86 5377 114
rect 5435 86 5463 114
rect 5521 86 5549 114
rect 5661 172 5689 200
rect 5747 172 5775 200
rect 5833 172 5861 200
rect 5919 172 5947 200
rect 5661 86 5689 114
rect 5747 86 5775 114
rect 5833 86 5861 114
rect 5919 86 5947 114
rect 6059 172 6087 200
rect 6145 172 6173 200
rect 6231 172 6259 200
rect 6317 172 6345 200
rect 6059 86 6087 114
rect 6145 86 6173 114
rect 6231 86 6259 114
rect 6317 86 6345 114
rect 6457 172 6485 200
rect 6543 172 6571 200
rect 6629 172 6657 200
rect 6715 172 6743 200
rect 6457 86 6485 114
rect 6543 86 6571 114
rect 6629 86 6657 114
rect 6715 86 6743 114
rect 6855 344 6883 372
rect 6941 344 6969 372
rect 7027 344 7055 372
rect 7113 344 7141 372
rect 6855 258 6883 286
rect 6941 258 6969 286
rect 7027 258 7055 286
rect 7113 258 7141 286
rect 6855 172 6883 200
rect 6941 172 6969 200
rect 7027 172 7055 200
rect 7113 172 7141 200
rect 6855 86 6883 114
rect 6941 86 6969 114
rect 7027 86 7055 114
rect 7113 86 7141 114
rect 7253 344 7281 372
rect 7339 344 7367 372
rect 7425 344 7453 372
rect 7511 344 7539 372
rect 7253 258 7281 286
rect 7339 258 7367 286
rect 7425 258 7453 286
rect 7511 258 7539 286
rect 7651 344 7679 372
rect 7737 344 7765 372
rect 7823 344 7851 372
rect 7909 344 7937 372
rect 7651 258 7679 286
rect 7737 258 7765 286
rect 7823 258 7851 286
rect 7909 258 7937 286
rect 8049 344 8077 372
rect 8135 344 8163 372
rect 8221 344 8249 372
rect 8307 344 8335 372
rect 8049 258 8077 286
rect 8135 258 8163 286
rect 8221 258 8249 286
rect 8307 258 8335 286
rect 8447 344 8475 372
rect 8533 344 8561 372
rect 8619 344 8647 372
rect 8705 344 8733 372
rect 8447 258 8475 286
rect 8533 258 8561 286
rect 8619 258 8647 286
rect 8705 258 8733 286
rect 7253 172 7281 200
rect 7339 172 7367 200
rect 7425 172 7453 200
rect 7511 172 7539 200
rect 7253 86 7281 114
rect 7339 86 7367 114
rect 7425 86 7453 114
rect 7511 86 7539 114
rect 7651 172 7679 200
rect 7737 172 7765 200
rect 7823 172 7851 200
rect 7909 172 7937 200
rect 7651 86 7679 114
rect 7737 86 7765 114
rect 7823 86 7851 114
rect 7909 86 7937 114
rect 8049 172 8077 200
rect 8135 172 8163 200
rect 8221 172 8249 200
rect 8307 172 8335 200
rect 8049 86 8077 114
rect 8135 86 8163 114
rect 8221 86 8249 114
rect 8307 86 8335 114
rect 8447 172 8475 200
rect 8533 172 8561 200
rect 8619 172 8647 200
rect 8705 172 8733 200
rect 8447 86 8475 114
rect 8533 86 8561 114
rect 8619 86 8647 114
rect 8705 86 8733 114
rect 8845 344 8873 372
rect 8931 344 8959 372
rect 9017 344 9045 372
rect 9103 344 9131 372
rect 8845 258 8873 286
rect 8931 258 8959 286
rect 9017 258 9045 286
rect 9103 258 9131 286
rect 8845 172 8873 200
rect 8931 172 8959 200
rect 9017 172 9045 200
rect 9103 172 9131 200
rect 8845 86 8873 114
rect 8931 86 8959 114
rect 9017 86 9045 114
rect 9103 86 9131 114
rect 9243 344 9271 372
rect 9329 344 9357 372
rect 9415 344 9443 372
rect 9501 344 9529 372
rect 9243 258 9271 286
rect 9329 258 9357 286
rect 9415 258 9443 286
rect 9501 258 9529 286
rect 9641 344 9669 372
rect 9727 344 9755 372
rect 9813 344 9841 372
rect 9899 344 9927 372
rect 9641 258 9669 286
rect 9727 258 9755 286
rect 9813 258 9841 286
rect 9899 258 9927 286
rect 9243 172 9271 200
rect 9329 172 9357 200
rect 9415 172 9443 200
rect 9501 172 9529 200
rect 9243 86 9271 114
rect 9329 86 9357 114
rect 9415 86 9443 114
rect 9501 86 9529 114
rect 9641 172 9669 200
rect 9727 172 9755 200
rect 9813 172 9841 200
rect 9899 172 9927 200
rect 9641 86 9669 114
rect 9727 86 9755 114
rect 9813 86 9841 114
rect 9899 86 9927 114
<< metal3 >>
rect 52 1674 406 1677
rect 52 1646 89 1674
rect 117 1646 175 1674
rect 203 1646 261 1674
rect 289 1646 347 1674
rect 375 1646 406 1674
rect 52 1643 406 1646
rect 450 1674 804 1677
rect 450 1646 487 1674
rect 515 1646 573 1674
rect 601 1646 659 1674
rect 687 1646 745 1674
rect 773 1646 804 1674
rect 450 1643 804 1646
rect 848 1674 1202 1677
rect 848 1646 885 1674
rect 913 1646 971 1674
rect 999 1646 1057 1674
rect 1085 1646 1143 1674
rect 1171 1646 1202 1674
rect 848 1643 1202 1646
rect 1246 1674 1600 1677
rect 1246 1646 1283 1674
rect 1311 1646 1369 1674
rect 1397 1646 1455 1674
rect 1483 1646 1541 1674
rect 1569 1646 1600 1674
rect 1246 1643 1600 1646
rect 1644 1674 1998 1677
rect 1644 1646 1681 1674
rect 1709 1646 1767 1674
rect 1795 1646 1853 1674
rect 1881 1646 1939 1674
rect 1967 1646 1998 1674
rect 1644 1643 1998 1646
rect 2042 1674 2396 1677
rect 2042 1646 2079 1674
rect 2107 1646 2165 1674
rect 2193 1646 2251 1674
rect 2279 1646 2337 1674
rect 2365 1646 2396 1674
rect 2042 1643 2396 1646
rect 2440 1674 2794 1677
rect 2440 1646 2477 1674
rect 2505 1646 2563 1674
rect 2591 1646 2649 1674
rect 2677 1646 2735 1674
rect 2763 1646 2794 1674
rect 2440 1643 2794 1646
rect 2838 1674 3192 1677
rect 2838 1646 2875 1674
rect 2903 1646 2961 1674
rect 2989 1646 3047 1674
rect 3075 1646 3133 1674
rect 3161 1646 3192 1674
rect 2838 1643 3192 1646
rect 3236 1674 3590 1677
rect 3236 1646 3273 1674
rect 3301 1646 3359 1674
rect 3387 1646 3445 1674
rect 3473 1646 3531 1674
rect 3559 1646 3590 1674
rect 3236 1643 3590 1646
rect 3634 1674 3988 1677
rect 3634 1646 3671 1674
rect 3699 1646 3757 1674
rect 3785 1646 3843 1674
rect 3871 1646 3929 1674
rect 3957 1646 3988 1674
rect 3634 1643 3988 1646
rect 4032 1674 4386 1677
rect 4032 1646 4069 1674
rect 4097 1646 4155 1674
rect 4183 1646 4241 1674
rect 4269 1646 4327 1674
rect 4355 1646 4386 1674
rect 4032 1643 4386 1646
rect 4430 1674 4784 1677
rect 4430 1646 4467 1674
rect 4495 1646 4553 1674
rect 4581 1646 4639 1674
rect 4667 1646 4725 1674
rect 4753 1646 4784 1674
rect 4430 1643 4784 1646
rect 4828 1674 5182 1677
rect 4828 1646 4865 1674
rect 4893 1646 4951 1674
rect 4979 1646 5037 1674
rect 5065 1646 5123 1674
rect 5151 1646 5182 1674
rect 4828 1643 5182 1646
rect 5226 1674 5580 1677
rect 5226 1646 5263 1674
rect 5291 1646 5349 1674
rect 5377 1646 5435 1674
rect 5463 1646 5521 1674
rect 5549 1646 5580 1674
rect 5226 1643 5580 1646
rect 5624 1674 5978 1677
rect 5624 1646 5661 1674
rect 5689 1646 5747 1674
rect 5775 1646 5833 1674
rect 5861 1646 5919 1674
rect 5947 1646 5978 1674
rect 5624 1643 5978 1646
rect 6022 1674 6376 1677
rect 6022 1646 6059 1674
rect 6087 1646 6145 1674
rect 6173 1646 6231 1674
rect 6259 1646 6317 1674
rect 6345 1646 6376 1674
rect 6022 1643 6376 1646
rect 6420 1674 6774 1677
rect 6420 1646 6457 1674
rect 6485 1646 6543 1674
rect 6571 1646 6629 1674
rect 6657 1646 6715 1674
rect 6743 1646 6774 1674
rect 6420 1643 6774 1646
rect 6818 1674 7172 1677
rect 6818 1646 6855 1674
rect 6883 1646 6941 1674
rect 6969 1646 7027 1674
rect 7055 1646 7113 1674
rect 7141 1646 7172 1674
rect 6818 1643 7172 1646
rect 7216 1674 7570 1677
rect 7216 1646 7253 1674
rect 7281 1646 7339 1674
rect 7367 1646 7425 1674
rect 7453 1646 7511 1674
rect 7539 1646 7570 1674
rect 7216 1643 7570 1646
rect 7614 1674 7968 1677
rect 7614 1646 7651 1674
rect 7679 1646 7737 1674
rect 7765 1646 7823 1674
rect 7851 1646 7909 1674
rect 7937 1646 7968 1674
rect 7614 1643 7968 1646
rect 8012 1674 8366 1677
rect 8012 1646 8049 1674
rect 8077 1646 8135 1674
rect 8163 1646 8221 1674
rect 8249 1646 8307 1674
rect 8335 1646 8366 1674
rect 8012 1643 8366 1646
rect 8410 1674 8764 1677
rect 8410 1646 8447 1674
rect 8475 1646 8533 1674
rect 8561 1646 8619 1674
rect 8647 1646 8705 1674
rect 8733 1646 8764 1674
rect 8410 1643 8764 1646
rect 8808 1674 9162 1677
rect 8808 1646 8845 1674
rect 8873 1646 8931 1674
rect 8959 1646 9017 1674
rect 9045 1646 9103 1674
rect 9131 1646 9162 1674
rect 8808 1643 9162 1646
rect 9206 1674 9560 1677
rect 9206 1646 9243 1674
rect 9271 1646 9329 1674
rect 9357 1646 9415 1674
rect 9443 1646 9501 1674
rect 9529 1646 9560 1674
rect 9206 1643 9560 1646
rect 9604 1674 9958 1677
rect 9604 1646 9641 1674
rect 9669 1646 9727 1674
rect 9755 1646 9813 1674
rect 9841 1646 9899 1674
rect 9927 1646 9958 1674
rect 9604 1643 9958 1646
rect 52 1588 406 1591
rect 52 1560 89 1588
rect 117 1560 175 1588
rect 203 1560 261 1588
rect 289 1560 347 1588
rect 375 1560 406 1588
rect 52 1557 406 1560
rect 450 1588 804 1591
rect 450 1560 487 1588
rect 515 1560 573 1588
rect 601 1560 659 1588
rect 687 1560 745 1588
rect 773 1560 804 1588
rect 450 1557 804 1560
rect 848 1588 1202 1591
rect 848 1560 885 1588
rect 913 1560 971 1588
rect 999 1560 1057 1588
rect 1085 1560 1143 1588
rect 1171 1560 1202 1588
rect 848 1557 1202 1560
rect 1246 1588 1600 1591
rect 1246 1560 1283 1588
rect 1311 1560 1369 1588
rect 1397 1560 1455 1588
rect 1483 1560 1541 1588
rect 1569 1560 1600 1588
rect 1246 1557 1600 1560
rect 1644 1588 1998 1591
rect 1644 1560 1681 1588
rect 1709 1560 1767 1588
rect 1795 1560 1853 1588
rect 1881 1560 1939 1588
rect 1967 1560 1998 1588
rect 1644 1557 1998 1560
rect 2042 1588 2396 1591
rect 2042 1560 2079 1588
rect 2107 1560 2165 1588
rect 2193 1560 2251 1588
rect 2279 1560 2337 1588
rect 2365 1560 2396 1588
rect 2042 1557 2396 1560
rect 2440 1588 2794 1591
rect 2440 1560 2477 1588
rect 2505 1560 2563 1588
rect 2591 1560 2649 1588
rect 2677 1560 2735 1588
rect 2763 1560 2794 1588
rect 2440 1557 2794 1560
rect 2838 1588 3192 1591
rect 2838 1560 2875 1588
rect 2903 1560 2961 1588
rect 2989 1560 3047 1588
rect 3075 1560 3133 1588
rect 3161 1560 3192 1588
rect 2838 1557 3192 1560
rect 3236 1588 3590 1591
rect 3236 1560 3273 1588
rect 3301 1560 3359 1588
rect 3387 1560 3445 1588
rect 3473 1560 3531 1588
rect 3559 1560 3590 1588
rect 3236 1557 3590 1560
rect 3634 1588 3988 1591
rect 3634 1560 3671 1588
rect 3699 1560 3757 1588
rect 3785 1560 3843 1588
rect 3871 1560 3929 1588
rect 3957 1560 3988 1588
rect 3634 1557 3988 1560
rect 4032 1588 4386 1591
rect 4032 1560 4069 1588
rect 4097 1560 4155 1588
rect 4183 1560 4241 1588
rect 4269 1560 4327 1588
rect 4355 1560 4386 1588
rect 4032 1557 4386 1560
rect 4430 1588 4784 1591
rect 4430 1560 4467 1588
rect 4495 1560 4553 1588
rect 4581 1560 4639 1588
rect 4667 1560 4725 1588
rect 4753 1560 4784 1588
rect 4430 1557 4784 1560
rect 4828 1588 5182 1591
rect 4828 1560 4865 1588
rect 4893 1560 4951 1588
rect 4979 1560 5037 1588
rect 5065 1560 5123 1588
rect 5151 1560 5182 1588
rect 4828 1557 5182 1560
rect 5226 1588 5580 1591
rect 5226 1560 5263 1588
rect 5291 1560 5349 1588
rect 5377 1560 5435 1588
rect 5463 1560 5521 1588
rect 5549 1560 5580 1588
rect 5226 1557 5580 1560
rect 5624 1588 5978 1591
rect 5624 1560 5661 1588
rect 5689 1560 5747 1588
rect 5775 1560 5833 1588
rect 5861 1560 5919 1588
rect 5947 1560 5978 1588
rect 5624 1557 5978 1560
rect 6022 1588 6376 1591
rect 6022 1560 6059 1588
rect 6087 1560 6145 1588
rect 6173 1560 6231 1588
rect 6259 1560 6317 1588
rect 6345 1560 6376 1588
rect 6022 1557 6376 1560
rect 6420 1588 6774 1591
rect 6420 1560 6457 1588
rect 6485 1560 6543 1588
rect 6571 1560 6629 1588
rect 6657 1560 6715 1588
rect 6743 1560 6774 1588
rect 6420 1557 6774 1560
rect 6818 1588 7172 1591
rect 6818 1560 6855 1588
rect 6883 1560 6941 1588
rect 6969 1560 7027 1588
rect 7055 1560 7113 1588
rect 7141 1560 7172 1588
rect 6818 1557 7172 1560
rect 7216 1588 7570 1591
rect 7216 1560 7253 1588
rect 7281 1560 7339 1588
rect 7367 1560 7425 1588
rect 7453 1560 7511 1588
rect 7539 1560 7570 1588
rect 7216 1557 7570 1560
rect 7614 1588 7968 1591
rect 7614 1560 7651 1588
rect 7679 1560 7737 1588
rect 7765 1560 7823 1588
rect 7851 1560 7909 1588
rect 7937 1560 7968 1588
rect 7614 1557 7968 1560
rect 8012 1588 8366 1591
rect 8012 1560 8049 1588
rect 8077 1560 8135 1588
rect 8163 1560 8221 1588
rect 8249 1560 8307 1588
rect 8335 1560 8366 1588
rect 8012 1557 8366 1560
rect 8410 1588 8764 1591
rect 8410 1560 8447 1588
rect 8475 1560 8533 1588
rect 8561 1560 8619 1588
rect 8647 1560 8705 1588
rect 8733 1560 8764 1588
rect 8410 1557 8764 1560
rect 8808 1588 9162 1591
rect 8808 1560 8845 1588
rect 8873 1560 8931 1588
rect 8959 1560 9017 1588
rect 9045 1560 9103 1588
rect 9131 1560 9162 1588
rect 8808 1557 9162 1560
rect 9206 1588 9560 1591
rect 9206 1560 9243 1588
rect 9271 1560 9329 1588
rect 9357 1560 9415 1588
rect 9443 1560 9501 1588
rect 9529 1560 9560 1588
rect 9206 1557 9560 1560
rect 9604 1588 9958 1591
rect 9604 1560 9641 1588
rect 9669 1560 9727 1588
rect 9755 1560 9813 1588
rect 9841 1560 9899 1588
rect 9927 1560 9958 1588
rect 9604 1557 9958 1560
rect 52 1502 406 1505
rect 52 1474 89 1502
rect 117 1474 175 1502
rect 203 1474 261 1502
rect 289 1474 347 1502
rect 375 1474 406 1502
rect 52 1471 406 1474
rect 450 1502 804 1505
rect 450 1474 487 1502
rect 515 1474 573 1502
rect 601 1474 659 1502
rect 687 1474 745 1502
rect 773 1474 804 1502
rect 450 1471 804 1474
rect 848 1502 1202 1505
rect 848 1474 885 1502
rect 913 1474 971 1502
rect 999 1474 1057 1502
rect 1085 1474 1143 1502
rect 1171 1474 1202 1502
rect 848 1471 1202 1474
rect 1246 1502 1600 1505
rect 1246 1474 1283 1502
rect 1311 1474 1369 1502
rect 1397 1474 1455 1502
rect 1483 1474 1541 1502
rect 1569 1474 1600 1502
rect 1246 1471 1600 1474
rect 1644 1502 1998 1505
rect 1644 1474 1681 1502
rect 1709 1474 1767 1502
rect 1795 1474 1853 1502
rect 1881 1474 1939 1502
rect 1967 1474 1998 1502
rect 1644 1471 1998 1474
rect 2042 1502 2396 1505
rect 2042 1474 2079 1502
rect 2107 1474 2165 1502
rect 2193 1474 2251 1502
rect 2279 1474 2337 1502
rect 2365 1474 2396 1502
rect 2042 1471 2396 1474
rect 2440 1502 2794 1505
rect 2440 1474 2477 1502
rect 2505 1474 2563 1502
rect 2591 1474 2649 1502
rect 2677 1474 2735 1502
rect 2763 1474 2794 1502
rect 2440 1471 2794 1474
rect 2838 1502 3192 1505
rect 2838 1474 2875 1502
rect 2903 1474 2961 1502
rect 2989 1474 3047 1502
rect 3075 1474 3133 1502
rect 3161 1474 3192 1502
rect 2838 1471 3192 1474
rect 3236 1502 3590 1505
rect 3236 1474 3273 1502
rect 3301 1474 3359 1502
rect 3387 1474 3445 1502
rect 3473 1474 3531 1502
rect 3559 1474 3590 1502
rect 3236 1471 3590 1474
rect 3634 1502 3988 1505
rect 3634 1474 3671 1502
rect 3699 1474 3757 1502
rect 3785 1474 3843 1502
rect 3871 1474 3929 1502
rect 3957 1474 3988 1502
rect 3634 1471 3988 1474
rect 4032 1502 4386 1505
rect 4032 1474 4069 1502
rect 4097 1474 4155 1502
rect 4183 1474 4241 1502
rect 4269 1474 4327 1502
rect 4355 1474 4386 1502
rect 4032 1471 4386 1474
rect 4430 1502 4784 1505
rect 4430 1474 4467 1502
rect 4495 1474 4553 1502
rect 4581 1474 4639 1502
rect 4667 1474 4725 1502
rect 4753 1474 4784 1502
rect 4430 1471 4784 1474
rect 4828 1502 5182 1505
rect 4828 1474 4865 1502
rect 4893 1474 4951 1502
rect 4979 1474 5037 1502
rect 5065 1474 5123 1502
rect 5151 1474 5182 1502
rect 4828 1471 5182 1474
rect 5226 1502 5580 1505
rect 5226 1474 5263 1502
rect 5291 1474 5349 1502
rect 5377 1474 5435 1502
rect 5463 1474 5521 1502
rect 5549 1474 5580 1502
rect 5226 1471 5580 1474
rect 5624 1502 5978 1505
rect 5624 1474 5661 1502
rect 5689 1474 5747 1502
rect 5775 1474 5833 1502
rect 5861 1474 5919 1502
rect 5947 1474 5978 1502
rect 5624 1471 5978 1474
rect 6022 1502 6376 1505
rect 6022 1474 6059 1502
rect 6087 1474 6145 1502
rect 6173 1474 6231 1502
rect 6259 1474 6317 1502
rect 6345 1474 6376 1502
rect 6022 1471 6376 1474
rect 6420 1502 6774 1505
rect 6420 1474 6457 1502
rect 6485 1474 6543 1502
rect 6571 1474 6629 1502
rect 6657 1474 6715 1502
rect 6743 1474 6774 1502
rect 6420 1471 6774 1474
rect 6818 1502 7172 1505
rect 6818 1474 6855 1502
rect 6883 1474 6941 1502
rect 6969 1474 7027 1502
rect 7055 1474 7113 1502
rect 7141 1474 7172 1502
rect 6818 1471 7172 1474
rect 7216 1502 7570 1505
rect 7216 1474 7253 1502
rect 7281 1474 7339 1502
rect 7367 1474 7425 1502
rect 7453 1474 7511 1502
rect 7539 1474 7570 1502
rect 7216 1471 7570 1474
rect 7614 1502 7968 1505
rect 7614 1474 7651 1502
rect 7679 1474 7737 1502
rect 7765 1474 7823 1502
rect 7851 1474 7909 1502
rect 7937 1474 7968 1502
rect 7614 1471 7968 1474
rect 8012 1502 8366 1505
rect 8012 1474 8049 1502
rect 8077 1474 8135 1502
rect 8163 1474 8221 1502
rect 8249 1474 8307 1502
rect 8335 1474 8366 1502
rect 8012 1471 8366 1474
rect 8410 1502 8764 1505
rect 8410 1474 8447 1502
rect 8475 1474 8533 1502
rect 8561 1474 8619 1502
rect 8647 1474 8705 1502
rect 8733 1474 8764 1502
rect 8410 1471 8764 1474
rect 8808 1502 9162 1505
rect 8808 1474 8845 1502
rect 8873 1474 8931 1502
rect 8959 1474 9017 1502
rect 9045 1474 9103 1502
rect 9131 1474 9162 1502
rect 8808 1471 9162 1474
rect 9206 1502 9560 1505
rect 9206 1474 9243 1502
rect 9271 1474 9329 1502
rect 9357 1474 9415 1502
rect 9443 1474 9501 1502
rect 9529 1474 9560 1502
rect 9206 1471 9560 1474
rect 9604 1502 9958 1505
rect 9604 1474 9641 1502
rect 9669 1474 9727 1502
rect 9755 1474 9813 1502
rect 9841 1474 9899 1502
rect 9927 1474 9958 1502
rect 9604 1471 9958 1474
rect 52 1416 406 1419
rect 52 1388 89 1416
rect 117 1388 175 1416
rect 203 1388 261 1416
rect 289 1388 347 1416
rect 375 1388 406 1416
rect 52 1385 406 1388
rect 450 1416 804 1419
rect 450 1388 487 1416
rect 515 1388 573 1416
rect 601 1388 659 1416
rect 687 1388 745 1416
rect 773 1388 804 1416
rect 450 1385 804 1388
rect 848 1416 1202 1419
rect 848 1388 885 1416
rect 913 1388 971 1416
rect 999 1388 1057 1416
rect 1085 1388 1143 1416
rect 1171 1388 1202 1416
rect 848 1385 1202 1388
rect 1246 1416 1600 1419
rect 1246 1388 1283 1416
rect 1311 1388 1369 1416
rect 1397 1388 1455 1416
rect 1483 1388 1541 1416
rect 1569 1388 1600 1416
rect 1246 1385 1600 1388
rect 1644 1416 1998 1419
rect 1644 1388 1681 1416
rect 1709 1388 1767 1416
rect 1795 1388 1853 1416
rect 1881 1388 1939 1416
rect 1967 1388 1998 1416
rect 1644 1385 1998 1388
rect 2042 1416 2396 1419
rect 2042 1388 2079 1416
rect 2107 1388 2165 1416
rect 2193 1388 2251 1416
rect 2279 1388 2337 1416
rect 2365 1388 2396 1416
rect 2042 1385 2396 1388
rect 2440 1416 2794 1419
rect 2440 1388 2477 1416
rect 2505 1388 2563 1416
rect 2591 1388 2649 1416
rect 2677 1388 2735 1416
rect 2763 1388 2794 1416
rect 2440 1385 2794 1388
rect 2838 1416 3192 1419
rect 2838 1388 2875 1416
rect 2903 1388 2961 1416
rect 2989 1388 3047 1416
rect 3075 1388 3133 1416
rect 3161 1388 3192 1416
rect 2838 1385 3192 1388
rect 3236 1416 3590 1419
rect 3236 1388 3273 1416
rect 3301 1388 3359 1416
rect 3387 1388 3445 1416
rect 3473 1388 3531 1416
rect 3559 1388 3590 1416
rect 3236 1385 3590 1388
rect 3634 1416 3988 1419
rect 3634 1388 3671 1416
rect 3699 1388 3757 1416
rect 3785 1388 3843 1416
rect 3871 1388 3929 1416
rect 3957 1388 3988 1416
rect 3634 1385 3988 1388
rect 4032 1416 4386 1419
rect 4032 1388 4069 1416
rect 4097 1388 4155 1416
rect 4183 1388 4241 1416
rect 4269 1388 4327 1416
rect 4355 1388 4386 1416
rect 4032 1385 4386 1388
rect 4430 1416 4784 1419
rect 4430 1388 4467 1416
rect 4495 1388 4553 1416
rect 4581 1388 4639 1416
rect 4667 1388 4725 1416
rect 4753 1388 4784 1416
rect 4430 1385 4784 1388
rect 4828 1416 5182 1419
rect 4828 1388 4865 1416
rect 4893 1388 4951 1416
rect 4979 1388 5037 1416
rect 5065 1388 5123 1416
rect 5151 1388 5182 1416
rect 4828 1385 5182 1388
rect 5226 1416 5580 1419
rect 5226 1388 5263 1416
rect 5291 1388 5349 1416
rect 5377 1388 5435 1416
rect 5463 1388 5521 1416
rect 5549 1388 5580 1416
rect 5226 1385 5580 1388
rect 5624 1416 5978 1419
rect 5624 1388 5661 1416
rect 5689 1388 5747 1416
rect 5775 1388 5833 1416
rect 5861 1388 5919 1416
rect 5947 1388 5978 1416
rect 5624 1385 5978 1388
rect 6022 1416 6376 1419
rect 6022 1388 6059 1416
rect 6087 1388 6145 1416
rect 6173 1388 6231 1416
rect 6259 1388 6317 1416
rect 6345 1388 6376 1416
rect 6022 1385 6376 1388
rect 6420 1416 6774 1419
rect 6420 1388 6457 1416
rect 6485 1388 6543 1416
rect 6571 1388 6629 1416
rect 6657 1388 6715 1416
rect 6743 1388 6774 1416
rect 6420 1385 6774 1388
rect 6818 1416 7172 1419
rect 6818 1388 6855 1416
rect 6883 1388 6941 1416
rect 6969 1388 7027 1416
rect 7055 1388 7113 1416
rect 7141 1388 7172 1416
rect 6818 1385 7172 1388
rect 7216 1416 7570 1419
rect 7216 1388 7253 1416
rect 7281 1388 7339 1416
rect 7367 1388 7425 1416
rect 7453 1388 7511 1416
rect 7539 1388 7570 1416
rect 7216 1385 7570 1388
rect 7614 1416 7968 1419
rect 7614 1388 7651 1416
rect 7679 1388 7737 1416
rect 7765 1388 7823 1416
rect 7851 1388 7909 1416
rect 7937 1388 7968 1416
rect 7614 1385 7968 1388
rect 8012 1416 8366 1419
rect 8012 1388 8049 1416
rect 8077 1388 8135 1416
rect 8163 1388 8221 1416
rect 8249 1388 8307 1416
rect 8335 1388 8366 1416
rect 8012 1385 8366 1388
rect 8410 1416 8764 1419
rect 8410 1388 8447 1416
rect 8475 1388 8533 1416
rect 8561 1388 8619 1416
rect 8647 1388 8705 1416
rect 8733 1388 8764 1416
rect 8410 1385 8764 1388
rect 8808 1416 9162 1419
rect 8808 1388 8845 1416
rect 8873 1388 8931 1416
rect 8959 1388 9017 1416
rect 9045 1388 9103 1416
rect 9131 1388 9162 1416
rect 8808 1385 9162 1388
rect 9206 1416 9560 1419
rect 9206 1388 9243 1416
rect 9271 1388 9329 1416
rect 9357 1388 9415 1416
rect 9443 1388 9501 1416
rect 9529 1388 9560 1416
rect 9206 1385 9560 1388
rect 9604 1416 9958 1419
rect 9604 1388 9641 1416
rect 9669 1388 9727 1416
rect 9755 1388 9813 1416
rect 9841 1388 9899 1416
rect 9927 1388 9958 1416
rect 9604 1385 9958 1388
rect 52 1240 406 1243
rect 52 1212 89 1240
rect 117 1212 175 1240
rect 203 1212 261 1240
rect 289 1212 347 1240
rect 375 1212 406 1240
rect 52 1209 406 1212
rect 450 1240 804 1243
rect 450 1212 487 1240
rect 515 1212 573 1240
rect 601 1212 659 1240
rect 687 1212 745 1240
rect 773 1212 804 1240
rect 450 1209 804 1212
rect 848 1240 1202 1243
rect 848 1212 885 1240
rect 913 1212 971 1240
rect 999 1212 1057 1240
rect 1085 1212 1143 1240
rect 1171 1212 1202 1240
rect 848 1209 1202 1212
rect 1246 1240 1600 1243
rect 1246 1212 1283 1240
rect 1311 1212 1369 1240
rect 1397 1212 1455 1240
rect 1483 1212 1541 1240
rect 1569 1212 1600 1240
rect 1246 1209 1600 1212
rect 1644 1240 1998 1243
rect 1644 1212 1681 1240
rect 1709 1212 1767 1240
rect 1795 1212 1853 1240
rect 1881 1212 1939 1240
rect 1967 1212 1998 1240
rect 1644 1209 1998 1212
rect 2042 1240 2396 1243
rect 2042 1212 2079 1240
rect 2107 1212 2165 1240
rect 2193 1212 2251 1240
rect 2279 1212 2337 1240
rect 2365 1212 2396 1240
rect 2042 1209 2396 1212
rect 2440 1240 2794 1243
rect 2440 1212 2477 1240
rect 2505 1212 2563 1240
rect 2591 1212 2649 1240
rect 2677 1212 2735 1240
rect 2763 1212 2794 1240
rect 2440 1209 2794 1212
rect 2838 1240 3192 1243
rect 2838 1212 2875 1240
rect 2903 1212 2961 1240
rect 2989 1212 3047 1240
rect 3075 1212 3133 1240
rect 3161 1212 3192 1240
rect 2838 1209 3192 1212
rect 3236 1240 3590 1243
rect 3236 1212 3273 1240
rect 3301 1212 3359 1240
rect 3387 1212 3445 1240
rect 3473 1212 3531 1240
rect 3559 1212 3590 1240
rect 3236 1209 3590 1212
rect 3634 1240 3988 1243
rect 3634 1212 3671 1240
rect 3699 1212 3757 1240
rect 3785 1212 3843 1240
rect 3871 1212 3929 1240
rect 3957 1212 3988 1240
rect 3634 1209 3988 1212
rect 4032 1240 4386 1243
rect 4032 1212 4069 1240
rect 4097 1212 4155 1240
rect 4183 1212 4241 1240
rect 4269 1212 4327 1240
rect 4355 1212 4386 1240
rect 4032 1209 4386 1212
rect 4430 1240 4784 1243
rect 4430 1212 4467 1240
rect 4495 1212 4553 1240
rect 4581 1212 4639 1240
rect 4667 1212 4725 1240
rect 4753 1212 4784 1240
rect 4430 1209 4784 1212
rect 4828 1240 5182 1243
rect 4828 1212 4865 1240
rect 4893 1212 4951 1240
rect 4979 1212 5037 1240
rect 5065 1212 5123 1240
rect 5151 1212 5182 1240
rect 4828 1209 5182 1212
rect 5226 1240 5580 1243
rect 5226 1212 5263 1240
rect 5291 1212 5349 1240
rect 5377 1212 5435 1240
rect 5463 1212 5521 1240
rect 5549 1212 5580 1240
rect 5226 1209 5580 1212
rect 5624 1240 5978 1243
rect 5624 1212 5661 1240
rect 5689 1212 5747 1240
rect 5775 1212 5833 1240
rect 5861 1212 5919 1240
rect 5947 1212 5978 1240
rect 5624 1209 5978 1212
rect 6022 1240 6376 1243
rect 6022 1212 6059 1240
rect 6087 1212 6145 1240
rect 6173 1212 6231 1240
rect 6259 1212 6317 1240
rect 6345 1212 6376 1240
rect 6022 1209 6376 1212
rect 6420 1240 6774 1243
rect 6420 1212 6457 1240
rect 6485 1212 6543 1240
rect 6571 1212 6629 1240
rect 6657 1212 6715 1240
rect 6743 1212 6774 1240
rect 6420 1209 6774 1212
rect 6818 1240 7172 1243
rect 6818 1212 6855 1240
rect 6883 1212 6941 1240
rect 6969 1212 7027 1240
rect 7055 1212 7113 1240
rect 7141 1212 7172 1240
rect 6818 1209 7172 1212
rect 7216 1240 7570 1243
rect 7216 1212 7253 1240
rect 7281 1212 7339 1240
rect 7367 1212 7425 1240
rect 7453 1212 7511 1240
rect 7539 1212 7570 1240
rect 7216 1209 7570 1212
rect 7614 1240 7968 1243
rect 7614 1212 7651 1240
rect 7679 1212 7737 1240
rect 7765 1212 7823 1240
rect 7851 1212 7909 1240
rect 7937 1212 7968 1240
rect 7614 1209 7968 1212
rect 8012 1240 8366 1243
rect 8012 1212 8049 1240
rect 8077 1212 8135 1240
rect 8163 1212 8221 1240
rect 8249 1212 8307 1240
rect 8335 1212 8366 1240
rect 8012 1209 8366 1212
rect 8410 1240 8764 1243
rect 8410 1212 8447 1240
rect 8475 1212 8533 1240
rect 8561 1212 8619 1240
rect 8647 1212 8705 1240
rect 8733 1212 8764 1240
rect 8410 1209 8764 1212
rect 8808 1240 9162 1243
rect 8808 1212 8845 1240
rect 8873 1212 8931 1240
rect 8959 1212 9017 1240
rect 9045 1212 9103 1240
rect 9131 1212 9162 1240
rect 8808 1209 9162 1212
rect 9206 1240 9560 1243
rect 9206 1212 9243 1240
rect 9271 1212 9329 1240
rect 9357 1212 9415 1240
rect 9443 1212 9501 1240
rect 9529 1212 9560 1240
rect 9206 1209 9560 1212
rect 9604 1240 9958 1243
rect 9604 1212 9641 1240
rect 9669 1212 9727 1240
rect 9755 1212 9813 1240
rect 9841 1212 9899 1240
rect 9927 1212 9958 1240
rect 9604 1209 9958 1212
rect 52 1154 406 1157
rect 52 1126 89 1154
rect 117 1126 175 1154
rect 203 1126 261 1154
rect 289 1126 347 1154
rect 375 1126 406 1154
rect 52 1123 406 1126
rect 450 1154 804 1157
rect 450 1126 487 1154
rect 515 1126 573 1154
rect 601 1126 659 1154
rect 687 1126 745 1154
rect 773 1126 804 1154
rect 450 1123 804 1126
rect 848 1154 1202 1157
rect 848 1126 885 1154
rect 913 1126 971 1154
rect 999 1126 1057 1154
rect 1085 1126 1143 1154
rect 1171 1126 1202 1154
rect 848 1123 1202 1126
rect 1246 1154 1600 1157
rect 1246 1126 1283 1154
rect 1311 1126 1369 1154
rect 1397 1126 1455 1154
rect 1483 1126 1541 1154
rect 1569 1126 1600 1154
rect 1246 1123 1600 1126
rect 1644 1154 1998 1157
rect 1644 1126 1681 1154
rect 1709 1126 1767 1154
rect 1795 1126 1853 1154
rect 1881 1126 1939 1154
rect 1967 1126 1998 1154
rect 1644 1123 1998 1126
rect 2042 1154 2396 1157
rect 2042 1126 2079 1154
rect 2107 1126 2165 1154
rect 2193 1126 2251 1154
rect 2279 1126 2337 1154
rect 2365 1126 2396 1154
rect 2042 1123 2396 1126
rect 2440 1154 2794 1157
rect 2440 1126 2477 1154
rect 2505 1126 2563 1154
rect 2591 1126 2649 1154
rect 2677 1126 2735 1154
rect 2763 1126 2794 1154
rect 2440 1123 2794 1126
rect 2838 1154 3192 1157
rect 2838 1126 2875 1154
rect 2903 1126 2961 1154
rect 2989 1126 3047 1154
rect 3075 1126 3133 1154
rect 3161 1126 3192 1154
rect 2838 1123 3192 1126
rect 3236 1154 3590 1157
rect 3236 1126 3273 1154
rect 3301 1126 3359 1154
rect 3387 1126 3445 1154
rect 3473 1126 3531 1154
rect 3559 1126 3590 1154
rect 3236 1123 3590 1126
rect 3634 1154 3988 1157
rect 3634 1126 3671 1154
rect 3699 1126 3757 1154
rect 3785 1126 3843 1154
rect 3871 1126 3929 1154
rect 3957 1126 3988 1154
rect 3634 1123 3988 1126
rect 4032 1154 4386 1157
rect 4032 1126 4069 1154
rect 4097 1126 4155 1154
rect 4183 1126 4241 1154
rect 4269 1126 4327 1154
rect 4355 1126 4386 1154
rect 4032 1123 4386 1126
rect 4430 1154 4784 1157
rect 4430 1126 4467 1154
rect 4495 1126 4553 1154
rect 4581 1126 4639 1154
rect 4667 1126 4725 1154
rect 4753 1126 4784 1154
rect 4430 1123 4784 1126
rect 4828 1154 5182 1157
rect 4828 1126 4865 1154
rect 4893 1126 4951 1154
rect 4979 1126 5037 1154
rect 5065 1126 5123 1154
rect 5151 1126 5182 1154
rect 4828 1123 5182 1126
rect 5226 1154 5580 1157
rect 5226 1126 5263 1154
rect 5291 1126 5349 1154
rect 5377 1126 5435 1154
rect 5463 1126 5521 1154
rect 5549 1126 5580 1154
rect 5226 1123 5580 1126
rect 5624 1154 5978 1157
rect 5624 1126 5661 1154
rect 5689 1126 5747 1154
rect 5775 1126 5833 1154
rect 5861 1126 5919 1154
rect 5947 1126 5978 1154
rect 5624 1123 5978 1126
rect 6022 1154 6376 1157
rect 6022 1126 6059 1154
rect 6087 1126 6145 1154
rect 6173 1126 6231 1154
rect 6259 1126 6317 1154
rect 6345 1126 6376 1154
rect 6022 1123 6376 1126
rect 6420 1154 6774 1157
rect 6420 1126 6457 1154
rect 6485 1126 6543 1154
rect 6571 1126 6629 1154
rect 6657 1126 6715 1154
rect 6743 1126 6774 1154
rect 6420 1123 6774 1126
rect 6818 1154 7172 1157
rect 6818 1126 6855 1154
rect 6883 1126 6941 1154
rect 6969 1126 7027 1154
rect 7055 1126 7113 1154
rect 7141 1126 7172 1154
rect 6818 1123 7172 1126
rect 7216 1154 7570 1157
rect 7216 1126 7253 1154
rect 7281 1126 7339 1154
rect 7367 1126 7425 1154
rect 7453 1126 7511 1154
rect 7539 1126 7570 1154
rect 7216 1123 7570 1126
rect 7614 1154 7968 1157
rect 7614 1126 7651 1154
rect 7679 1126 7737 1154
rect 7765 1126 7823 1154
rect 7851 1126 7909 1154
rect 7937 1126 7968 1154
rect 7614 1123 7968 1126
rect 8012 1154 8366 1157
rect 8012 1126 8049 1154
rect 8077 1126 8135 1154
rect 8163 1126 8221 1154
rect 8249 1126 8307 1154
rect 8335 1126 8366 1154
rect 8012 1123 8366 1126
rect 8410 1154 8764 1157
rect 8410 1126 8447 1154
rect 8475 1126 8533 1154
rect 8561 1126 8619 1154
rect 8647 1126 8705 1154
rect 8733 1126 8764 1154
rect 8410 1123 8764 1126
rect 8808 1154 9162 1157
rect 8808 1126 8845 1154
rect 8873 1126 8931 1154
rect 8959 1126 9017 1154
rect 9045 1126 9103 1154
rect 9131 1126 9162 1154
rect 8808 1123 9162 1126
rect 9206 1154 9560 1157
rect 9206 1126 9243 1154
rect 9271 1126 9329 1154
rect 9357 1126 9415 1154
rect 9443 1126 9501 1154
rect 9529 1126 9560 1154
rect 9206 1123 9560 1126
rect 9604 1154 9958 1157
rect 9604 1126 9641 1154
rect 9669 1126 9727 1154
rect 9755 1126 9813 1154
rect 9841 1126 9899 1154
rect 9927 1126 9958 1154
rect 9604 1123 9958 1126
rect 52 1068 406 1071
rect 52 1040 89 1068
rect 117 1040 175 1068
rect 203 1040 261 1068
rect 289 1040 347 1068
rect 375 1040 406 1068
rect 52 1037 406 1040
rect 450 1068 804 1071
rect 450 1040 487 1068
rect 515 1040 573 1068
rect 601 1040 659 1068
rect 687 1040 745 1068
rect 773 1040 804 1068
rect 450 1037 804 1040
rect 848 1068 1202 1071
rect 848 1040 885 1068
rect 913 1040 971 1068
rect 999 1040 1057 1068
rect 1085 1040 1143 1068
rect 1171 1040 1202 1068
rect 848 1037 1202 1040
rect 1246 1068 1600 1071
rect 1246 1040 1283 1068
rect 1311 1040 1369 1068
rect 1397 1040 1455 1068
rect 1483 1040 1541 1068
rect 1569 1040 1600 1068
rect 1246 1037 1600 1040
rect 1644 1068 1998 1071
rect 1644 1040 1681 1068
rect 1709 1040 1767 1068
rect 1795 1040 1853 1068
rect 1881 1040 1939 1068
rect 1967 1040 1998 1068
rect 1644 1037 1998 1040
rect 2042 1068 2396 1071
rect 2042 1040 2079 1068
rect 2107 1040 2165 1068
rect 2193 1040 2251 1068
rect 2279 1040 2337 1068
rect 2365 1040 2396 1068
rect 2042 1037 2396 1040
rect 2440 1068 2794 1071
rect 2440 1040 2477 1068
rect 2505 1040 2563 1068
rect 2591 1040 2649 1068
rect 2677 1040 2735 1068
rect 2763 1040 2794 1068
rect 2440 1037 2794 1040
rect 2838 1068 3192 1071
rect 2838 1040 2875 1068
rect 2903 1040 2961 1068
rect 2989 1040 3047 1068
rect 3075 1040 3133 1068
rect 3161 1040 3192 1068
rect 2838 1037 3192 1040
rect 3236 1068 3590 1071
rect 3236 1040 3273 1068
rect 3301 1040 3359 1068
rect 3387 1040 3445 1068
rect 3473 1040 3531 1068
rect 3559 1040 3590 1068
rect 3236 1037 3590 1040
rect 3634 1068 3988 1071
rect 3634 1040 3671 1068
rect 3699 1040 3757 1068
rect 3785 1040 3843 1068
rect 3871 1040 3929 1068
rect 3957 1040 3988 1068
rect 3634 1037 3988 1040
rect 4032 1068 4386 1071
rect 4032 1040 4069 1068
rect 4097 1040 4155 1068
rect 4183 1040 4241 1068
rect 4269 1040 4327 1068
rect 4355 1040 4386 1068
rect 4032 1037 4386 1040
rect 4430 1068 4784 1071
rect 4430 1040 4467 1068
rect 4495 1040 4553 1068
rect 4581 1040 4639 1068
rect 4667 1040 4725 1068
rect 4753 1040 4784 1068
rect 4430 1037 4784 1040
rect 4828 1068 5182 1071
rect 4828 1040 4865 1068
rect 4893 1040 4951 1068
rect 4979 1040 5037 1068
rect 5065 1040 5123 1068
rect 5151 1040 5182 1068
rect 4828 1037 5182 1040
rect 5226 1068 5580 1071
rect 5226 1040 5263 1068
rect 5291 1040 5349 1068
rect 5377 1040 5435 1068
rect 5463 1040 5521 1068
rect 5549 1040 5580 1068
rect 5226 1037 5580 1040
rect 5624 1068 5978 1071
rect 5624 1040 5661 1068
rect 5689 1040 5747 1068
rect 5775 1040 5833 1068
rect 5861 1040 5919 1068
rect 5947 1040 5978 1068
rect 5624 1037 5978 1040
rect 6022 1068 6376 1071
rect 6022 1040 6059 1068
rect 6087 1040 6145 1068
rect 6173 1040 6231 1068
rect 6259 1040 6317 1068
rect 6345 1040 6376 1068
rect 6022 1037 6376 1040
rect 6420 1068 6774 1071
rect 6420 1040 6457 1068
rect 6485 1040 6543 1068
rect 6571 1040 6629 1068
rect 6657 1040 6715 1068
rect 6743 1040 6774 1068
rect 6420 1037 6774 1040
rect 6818 1068 7172 1071
rect 6818 1040 6855 1068
rect 6883 1040 6941 1068
rect 6969 1040 7027 1068
rect 7055 1040 7113 1068
rect 7141 1040 7172 1068
rect 6818 1037 7172 1040
rect 7216 1068 7570 1071
rect 7216 1040 7253 1068
rect 7281 1040 7339 1068
rect 7367 1040 7425 1068
rect 7453 1040 7511 1068
rect 7539 1040 7570 1068
rect 7216 1037 7570 1040
rect 7614 1068 7968 1071
rect 7614 1040 7651 1068
rect 7679 1040 7737 1068
rect 7765 1040 7823 1068
rect 7851 1040 7909 1068
rect 7937 1040 7968 1068
rect 7614 1037 7968 1040
rect 8012 1068 8366 1071
rect 8012 1040 8049 1068
rect 8077 1040 8135 1068
rect 8163 1040 8221 1068
rect 8249 1040 8307 1068
rect 8335 1040 8366 1068
rect 8012 1037 8366 1040
rect 8410 1068 8764 1071
rect 8410 1040 8447 1068
rect 8475 1040 8533 1068
rect 8561 1040 8619 1068
rect 8647 1040 8705 1068
rect 8733 1040 8764 1068
rect 8410 1037 8764 1040
rect 8808 1068 9162 1071
rect 8808 1040 8845 1068
rect 8873 1040 8931 1068
rect 8959 1040 9017 1068
rect 9045 1040 9103 1068
rect 9131 1040 9162 1068
rect 8808 1037 9162 1040
rect 9206 1068 9560 1071
rect 9206 1040 9243 1068
rect 9271 1040 9329 1068
rect 9357 1040 9415 1068
rect 9443 1040 9501 1068
rect 9529 1040 9560 1068
rect 9206 1037 9560 1040
rect 9604 1068 9958 1071
rect 9604 1040 9641 1068
rect 9669 1040 9727 1068
rect 9755 1040 9813 1068
rect 9841 1040 9899 1068
rect 9927 1040 9958 1068
rect 9604 1037 9958 1040
rect 52 982 406 985
rect 52 954 89 982
rect 117 954 175 982
rect 203 954 261 982
rect 289 954 347 982
rect 375 954 406 982
rect 52 951 406 954
rect 450 982 804 985
rect 450 954 487 982
rect 515 954 573 982
rect 601 954 659 982
rect 687 954 745 982
rect 773 954 804 982
rect 450 951 804 954
rect 848 982 1202 985
rect 848 954 885 982
rect 913 954 971 982
rect 999 954 1057 982
rect 1085 954 1143 982
rect 1171 954 1202 982
rect 848 951 1202 954
rect 1246 982 1600 985
rect 1246 954 1283 982
rect 1311 954 1369 982
rect 1397 954 1455 982
rect 1483 954 1541 982
rect 1569 954 1600 982
rect 1246 951 1600 954
rect 1644 982 1998 985
rect 1644 954 1681 982
rect 1709 954 1767 982
rect 1795 954 1853 982
rect 1881 954 1939 982
rect 1967 954 1998 982
rect 1644 951 1998 954
rect 2042 982 2396 985
rect 2042 954 2079 982
rect 2107 954 2165 982
rect 2193 954 2251 982
rect 2279 954 2337 982
rect 2365 954 2396 982
rect 2042 951 2396 954
rect 2440 982 2794 985
rect 2440 954 2477 982
rect 2505 954 2563 982
rect 2591 954 2649 982
rect 2677 954 2735 982
rect 2763 954 2794 982
rect 2440 951 2794 954
rect 2838 982 3192 985
rect 2838 954 2875 982
rect 2903 954 2961 982
rect 2989 954 3047 982
rect 3075 954 3133 982
rect 3161 954 3192 982
rect 2838 951 3192 954
rect 3236 982 3590 985
rect 3236 954 3273 982
rect 3301 954 3359 982
rect 3387 954 3445 982
rect 3473 954 3531 982
rect 3559 954 3590 982
rect 3236 951 3590 954
rect 3634 982 3988 985
rect 3634 954 3671 982
rect 3699 954 3757 982
rect 3785 954 3843 982
rect 3871 954 3929 982
rect 3957 954 3988 982
rect 3634 951 3988 954
rect 4032 982 4386 985
rect 4032 954 4069 982
rect 4097 954 4155 982
rect 4183 954 4241 982
rect 4269 954 4327 982
rect 4355 954 4386 982
rect 4032 951 4386 954
rect 4430 982 4784 985
rect 4430 954 4467 982
rect 4495 954 4553 982
rect 4581 954 4639 982
rect 4667 954 4725 982
rect 4753 954 4784 982
rect 4430 951 4784 954
rect 4828 982 5182 985
rect 4828 954 4865 982
rect 4893 954 4951 982
rect 4979 954 5037 982
rect 5065 954 5123 982
rect 5151 954 5182 982
rect 4828 951 5182 954
rect 5226 982 5580 985
rect 5226 954 5263 982
rect 5291 954 5349 982
rect 5377 954 5435 982
rect 5463 954 5521 982
rect 5549 954 5580 982
rect 5226 951 5580 954
rect 5624 982 5978 985
rect 5624 954 5661 982
rect 5689 954 5747 982
rect 5775 954 5833 982
rect 5861 954 5919 982
rect 5947 954 5978 982
rect 5624 951 5978 954
rect 6022 982 6376 985
rect 6022 954 6059 982
rect 6087 954 6145 982
rect 6173 954 6231 982
rect 6259 954 6317 982
rect 6345 954 6376 982
rect 6022 951 6376 954
rect 6420 982 6774 985
rect 6420 954 6457 982
rect 6485 954 6543 982
rect 6571 954 6629 982
rect 6657 954 6715 982
rect 6743 954 6774 982
rect 6420 951 6774 954
rect 6818 982 7172 985
rect 6818 954 6855 982
rect 6883 954 6941 982
rect 6969 954 7027 982
rect 7055 954 7113 982
rect 7141 954 7172 982
rect 6818 951 7172 954
rect 7216 982 7570 985
rect 7216 954 7253 982
rect 7281 954 7339 982
rect 7367 954 7425 982
rect 7453 954 7511 982
rect 7539 954 7570 982
rect 7216 951 7570 954
rect 7614 982 7968 985
rect 7614 954 7651 982
rect 7679 954 7737 982
rect 7765 954 7823 982
rect 7851 954 7909 982
rect 7937 954 7968 982
rect 7614 951 7968 954
rect 8012 982 8366 985
rect 8012 954 8049 982
rect 8077 954 8135 982
rect 8163 954 8221 982
rect 8249 954 8307 982
rect 8335 954 8366 982
rect 8012 951 8366 954
rect 8410 982 8764 985
rect 8410 954 8447 982
rect 8475 954 8533 982
rect 8561 954 8619 982
rect 8647 954 8705 982
rect 8733 954 8764 982
rect 8410 951 8764 954
rect 8808 982 9162 985
rect 8808 954 8845 982
rect 8873 954 8931 982
rect 8959 954 9017 982
rect 9045 954 9103 982
rect 9131 954 9162 982
rect 8808 951 9162 954
rect 9206 982 9560 985
rect 9206 954 9243 982
rect 9271 954 9329 982
rect 9357 954 9415 982
rect 9443 954 9501 982
rect 9529 954 9560 982
rect 9206 951 9560 954
rect 9604 982 9958 985
rect 9604 954 9641 982
rect 9669 954 9727 982
rect 9755 954 9813 982
rect 9841 954 9899 982
rect 9927 954 9958 982
rect 9604 951 9958 954
rect 52 806 406 809
rect 52 778 89 806
rect 117 778 175 806
rect 203 778 261 806
rect 289 778 347 806
rect 375 778 406 806
rect 52 775 406 778
rect 450 806 804 809
rect 450 778 487 806
rect 515 778 573 806
rect 601 778 659 806
rect 687 778 745 806
rect 773 778 804 806
rect 450 775 804 778
rect 848 806 1202 809
rect 848 778 885 806
rect 913 778 971 806
rect 999 778 1057 806
rect 1085 778 1143 806
rect 1171 778 1202 806
rect 848 775 1202 778
rect 1246 806 1600 809
rect 1246 778 1283 806
rect 1311 778 1369 806
rect 1397 778 1455 806
rect 1483 778 1541 806
rect 1569 778 1600 806
rect 1246 775 1600 778
rect 1644 806 1998 809
rect 1644 778 1681 806
rect 1709 778 1767 806
rect 1795 778 1853 806
rect 1881 778 1939 806
rect 1967 778 1998 806
rect 1644 775 1998 778
rect 2042 806 2396 809
rect 2042 778 2079 806
rect 2107 778 2165 806
rect 2193 778 2251 806
rect 2279 778 2337 806
rect 2365 778 2396 806
rect 2042 775 2396 778
rect 2440 806 2794 809
rect 2440 778 2477 806
rect 2505 778 2563 806
rect 2591 778 2649 806
rect 2677 778 2735 806
rect 2763 778 2794 806
rect 2440 775 2794 778
rect 2838 806 3192 809
rect 2838 778 2875 806
rect 2903 778 2961 806
rect 2989 778 3047 806
rect 3075 778 3133 806
rect 3161 778 3192 806
rect 2838 775 3192 778
rect 3236 806 3590 809
rect 3236 778 3273 806
rect 3301 778 3359 806
rect 3387 778 3445 806
rect 3473 778 3531 806
rect 3559 778 3590 806
rect 3236 775 3590 778
rect 3634 806 3988 809
rect 3634 778 3671 806
rect 3699 778 3757 806
rect 3785 778 3843 806
rect 3871 778 3929 806
rect 3957 778 3988 806
rect 3634 775 3988 778
rect 4032 806 4386 809
rect 4032 778 4069 806
rect 4097 778 4155 806
rect 4183 778 4241 806
rect 4269 778 4327 806
rect 4355 778 4386 806
rect 4032 775 4386 778
rect 4430 806 4784 809
rect 4430 778 4467 806
rect 4495 778 4553 806
rect 4581 778 4639 806
rect 4667 778 4725 806
rect 4753 778 4784 806
rect 4430 775 4784 778
rect 4828 806 5182 809
rect 4828 778 4865 806
rect 4893 778 4951 806
rect 4979 778 5037 806
rect 5065 778 5123 806
rect 5151 778 5182 806
rect 4828 775 5182 778
rect 5226 806 5580 809
rect 5226 778 5263 806
rect 5291 778 5349 806
rect 5377 778 5435 806
rect 5463 778 5521 806
rect 5549 778 5580 806
rect 5226 775 5580 778
rect 5624 806 5978 809
rect 5624 778 5661 806
rect 5689 778 5747 806
rect 5775 778 5833 806
rect 5861 778 5919 806
rect 5947 778 5978 806
rect 5624 775 5978 778
rect 6022 806 6376 809
rect 6022 778 6059 806
rect 6087 778 6145 806
rect 6173 778 6231 806
rect 6259 778 6317 806
rect 6345 778 6376 806
rect 6022 775 6376 778
rect 6420 806 6774 809
rect 6420 778 6457 806
rect 6485 778 6543 806
rect 6571 778 6629 806
rect 6657 778 6715 806
rect 6743 778 6774 806
rect 6420 775 6774 778
rect 6818 806 7172 809
rect 6818 778 6855 806
rect 6883 778 6941 806
rect 6969 778 7027 806
rect 7055 778 7113 806
rect 7141 778 7172 806
rect 6818 775 7172 778
rect 7216 806 7570 809
rect 7216 778 7253 806
rect 7281 778 7339 806
rect 7367 778 7425 806
rect 7453 778 7511 806
rect 7539 778 7570 806
rect 7216 775 7570 778
rect 7614 806 7968 809
rect 7614 778 7651 806
rect 7679 778 7737 806
rect 7765 778 7823 806
rect 7851 778 7909 806
rect 7937 778 7968 806
rect 7614 775 7968 778
rect 8012 806 8366 809
rect 8012 778 8049 806
rect 8077 778 8135 806
rect 8163 778 8221 806
rect 8249 778 8307 806
rect 8335 778 8366 806
rect 8012 775 8366 778
rect 8410 806 8764 809
rect 8410 778 8447 806
rect 8475 778 8533 806
rect 8561 778 8619 806
rect 8647 778 8705 806
rect 8733 778 8764 806
rect 8410 775 8764 778
rect 8808 806 9162 809
rect 8808 778 8845 806
rect 8873 778 8931 806
rect 8959 778 9017 806
rect 9045 778 9103 806
rect 9131 778 9162 806
rect 8808 775 9162 778
rect 9206 806 9560 809
rect 9206 778 9243 806
rect 9271 778 9329 806
rect 9357 778 9415 806
rect 9443 778 9501 806
rect 9529 778 9560 806
rect 9206 775 9560 778
rect 9604 806 9958 809
rect 9604 778 9641 806
rect 9669 778 9727 806
rect 9755 778 9813 806
rect 9841 778 9899 806
rect 9927 778 9958 806
rect 9604 775 9958 778
rect 52 720 406 723
rect 52 692 89 720
rect 117 692 175 720
rect 203 692 261 720
rect 289 692 347 720
rect 375 692 406 720
rect 52 689 406 692
rect 450 720 804 723
rect 450 692 487 720
rect 515 692 573 720
rect 601 692 659 720
rect 687 692 745 720
rect 773 692 804 720
rect 450 689 804 692
rect 848 720 1202 723
rect 848 692 885 720
rect 913 692 971 720
rect 999 692 1057 720
rect 1085 692 1143 720
rect 1171 692 1202 720
rect 848 689 1202 692
rect 1246 720 1600 723
rect 1246 692 1283 720
rect 1311 692 1369 720
rect 1397 692 1455 720
rect 1483 692 1541 720
rect 1569 692 1600 720
rect 1246 689 1600 692
rect 1644 720 1998 723
rect 1644 692 1681 720
rect 1709 692 1767 720
rect 1795 692 1853 720
rect 1881 692 1939 720
rect 1967 692 1998 720
rect 1644 689 1998 692
rect 2042 720 2396 723
rect 2042 692 2079 720
rect 2107 692 2165 720
rect 2193 692 2251 720
rect 2279 692 2337 720
rect 2365 692 2396 720
rect 2042 689 2396 692
rect 2440 720 2794 723
rect 2440 692 2477 720
rect 2505 692 2563 720
rect 2591 692 2649 720
rect 2677 692 2735 720
rect 2763 692 2794 720
rect 2440 689 2794 692
rect 2838 720 3192 723
rect 2838 692 2875 720
rect 2903 692 2961 720
rect 2989 692 3047 720
rect 3075 692 3133 720
rect 3161 692 3192 720
rect 2838 689 3192 692
rect 3236 720 3590 723
rect 3236 692 3273 720
rect 3301 692 3359 720
rect 3387 692 3445 720
rect 3473 692 3531 720
rect 3559 692 3590 720
rect 3236 689 3590 692
rect 3634 720 3988 723
rect 3634 692 3671 720
rect 3699 692 3757 720
rect 3785 692 3843 720
rect 3871 692 3929 720
rect 3957 692 3988 720
rect 3634 689 3988 692
rect 4032 720 4386 723
rect 4032 692 4069 720
rect 4097 692 4155 720
rect 4183 692 4241 720
rect 4269 692 4327 720
rect 4355 692 4386 720
rect 4032 689 4386 692
rect 4430 720 4784 723
rect 4430 692 4467 720
rect 4495 692 4553 720
rect 4581 692 4639 720
rect 4667 692 4725 720
rect 4753 692 4784 720
rect 4430 689 4784 692
rect 4828 720 5182 723
rect 4828 692 4865 720
rect 4893 692 4951 720
rect 4979 692 5037 720
rect 5065 692 5123 720
rect 5151 692 5182 720
rect 4828 689 5182 692
rect 5226 720 5580 723
rect 5226 692 5263 720
rect 5291 692 5349 720
rect 5377 692 5435 720
rect 5463 692 5521 720
rect 5549 692 5580 720
rect 5226 689 5580 692
rect 5624 720 5978 723
rect 5624 692 5661 720
rect 5689 692 5747 720
rect 5775 692 5833 720
rect 5861 692 5919 720
rect 5947 692 5978 720
rect 5624 689 5978 692
rect 6022 720 6376 723
rect 6022 692 6059 720
rect 6087 692 6145 720
rect 6173 692 6231 720
rect 6259 692 6317 720
rect 6345 692 6376 720
rect 6022 689 6376 692
rect 6420 720 6774 723
rect 6420 692 6457 720
rect 6485 692 6543 720
rect 6571 692 6629 720
rect 6657 692 6715 720
rect 6743 692 6774 720
rect 6420 689 6774 692
rect 6818 720 7172 723
rect 6818 692 6855 720
rect 6883 692 6941 720
rect 6969 692 7027 720
rect 7055 692 7113 720
rect 7141 692 7172 720
rect 6818 689 7172 692
rect 7216 720 7570 723
rect 7216 692 7253 720
rect 7281 692 7339 720
rect 7367 692 7425 720
rect 7453 692 7511 720
rect 7539 692 7570 720
rect 7216 689 7570 692
rect 7614 720 7968 723
rect 7614 692 7651 720
rect 7679 692 7737 720
rect 7765 692 7823 720
rect 7851 692 7909 720
rect 7937 692 7968 720
rect 7614 689 7968 692
rect 8012 720 8366 723
rect 8012 692 8049 720
rect 8077 692 8135 720
rect 8163 692 8221 720
rect 8249 692 8307 720
rect 8335 692 8366 720
rect 8012 689 8366 692
rect 8410 720 8764 723
rect 8410 692 8447 720
rect 8475 692 8533 720
rect 8561 692 8619 720
rect 8647 692 8705 720
rect 8733 692 8764 720
rect 8410 689 8764 692
rect 8808 720 9162 723
rect 8808 692 8845 720
rect 8873 692 8931 720
rect 8959 692 9017 720
rect 9045 692 9103 720
rect 9131 692 9162 720
rect 8808 689 9162 692
rect 9206 720 9560 723
rect 9206 692 9243 720
rect 9271 692 9329 720
rect 9357 692 9415 720
rect 9443 692 9501 720
rect 9529 692 9560 720
rect 9206 689 9560 692
rect 9604 720 9958 723
rect 9604 692 9641 720
rect 9669 692 9727 720
rect 9755 692 9813 720
rect 9841 692 9899 720
rect 9927 692 9958 720
rect 9604 689 9958 692
rect 52 634 406 637
rect 52 606 89 634
rect 117 606 175 634
rect 203 606 261 634
rect 289 606 347 634
rect 375 606 406 634
rect 52 603 406 606
rect 450 634 804 637
rect 450 606 487 634
rect 515 606 573 634
rect 601 606 659 634
rect 687 606 745 634
rect 773 606 804 634
rect 450 603 804 606
rect 848 634 1202 637
rect 848 606 885 634
rect 913 606 971 634
rect 999 606 1057 634
rect 1085 606 1143 634
rect 1171 606 1202 634
rect 848 603 1202 606
rect 1246 634 1600 637
rect 1246 606 1283 634
rect 1311 606 1369 634
rect 1397 606 1455 634
rect 1483 606 1541 634
rect 1569 606 1600 634
rect 1246 603 1600 606
rect 1644 634 1998 637
rect 1644 606 1681 634
rect 1709 606 1767 634
rect 1795 606 1853 634
rect 1881 606 1939 634
rect 1967 606 1998 634
rect 1644 603 1998 606
rect 2042 634 2396 637
rect 2042 606 2079 634
rect 2107 606 2165 634
rect 2193 606 2251 634
rect 2279 606 2337 634
rect 2365 606 2396 634
rect 2042 603 2396 606
rect 2440 634 2794 637
rect 2440 606 2477 634
rect 2505 606 2563 634
rect 2591 606 2649 634
rect 2677 606 2735 634
rect 2763 606 2794 634
rect 2440 603 2794 606
rect 2838 634 3192 637
rect 2838 606 2875 634
rect 2903 606 2961 634
rect 2989 606 3047 634
rect 3075 606 3133 634
rect 3161 606 3192 634
rect 2838 603 3192 606
rect 3236 634 3590 637
rect 3236 606 3273 634
rect 3301 606 3359 634
rect 3387 606 3445 634
rect 3473 606 3531 634
rect 3559 606 3590 634
rect 3236 603 3590 606
rect 3634 634 3988 637
rect 3634 606 3671 634
rect 3699 606 3757 634
rect 3785 606 3843 634
rect 3871 606 3929 634
rect 3957 606 3988 634
rect 3634 603 3988 606
rect 4032 634 4386 637
rect 4032 606 4069 634
rect 4097 606 4155 634
rect 4183 606 4241 634
rect 4269 606 4327 634
rect 4355 606 4386 634
rect 4032 603 4386 606
rect 4430 634 4784 637
rect 4430 606 4467 634
rect 4495 606 4553 634
rect 4581 606 4639 634
rect 4667 606 4725 634
rect 4753 606 4784 634
rect 4430 603 4784 606
rect 4828 634 5182 637
rect 4828 606 4865 634
rect 4893 606 4951 634
rect 4979 606 5037 634
rect 5065 606 5123 634
rect 5151 606 5182 634
rect 4828 603 5182 606
rect 5226 634 5580 637
rect 5226 606 5263 634
rect 5291 606 5349 634
rect 5377 606 5435 634
rect 5463 606 5521 634
rect 5549 606 5580 634
rect 5226 603 5580 606
rect 5624 634 5978 637
rect 5624 606 5661 634
rect 5689 606 5747 634
rect 5775 606 5833 634
rect 5861 606 5919 634
rect 5947 606 5978 634
rect 5624 603 5978 606
rect 6022 634 6376 637
rect 6022 606 6059 634
rect 6087 606 6145 634
rect 6173 606 6231 634
rect 6259 606 6317 634
rect 6345 606 6376 634
rect 6022 603 6376 606
rect 6420 634 6774 637
rect 6420 606 6457 634
rect 6485 606 6543 634
rect 6571 606 6629 634
rect 6657 606 6715 634
rect 6743 606 6774 634
rect 6420 603 6774 606
rect 6818 634 7172 637
rect 6818 606 6855 634
rect 6883 606 6941 634
rect 6969 606 7027 634
rect 7055 606 7113 634
rect 7141 606 7172 634
rect 6818 603 7172 606
rect 7216 634 7570 637
rect 7216 606 7253 634
rect 7281 606 7339 634
rect 7367 606 7425 634
rect 7453 606 7511 634
rect 7539 606 7570 634
rect 7216 603 7570 606
rect 7614 634 7968 637
rect 7614 606 7651 634
rect 7679 606 7737 634
rect 7765 606 7823 634
rect 7851 606 7909 634
rect 7937 606 7968 634
rect 7614 603 7968 606
rect 8012 634 8366 637
rect 8012 606 8049 634
rect 8077 606 8135 634
rect 8163 606 8221 634
rect 8249 606 8307 634
rect 8335 606 8366 634
rect 8012 603 8366 606
rect 8410 634 8764 637
rect 8410 606 8447 634
rect 8475 606 8533 634
rect 8561 606 8619 634
rect 8647 606 8705 634
rect 8733 606 8764 634
rect 8410 603 8764 606
rect 8808 634 9162 637
rect 8808 606 8845 634
rect 8873 606 8931 634
rect 8959 606 9017 634
rect 9045 606 9103 634
rect 9131 606 9162 634
rect 8808 603 9162 606
rect 9206 634 9560 637
rect 9206 606 9243 634
rect 9271 606 9329 634
rect 9357 606 9415 634
rect 9443 606 9501 634
rect 9529 606 9560 634
rect 9206 603 9560 606
rect 9604 634 9958 637
rect 9604 606 9641 634
rect 9669 606 9727 634
rect 9755 606 9813 634
rect 9841 606 9899 634
rect 9927 606 9958 634
rect 9604 603 9958 606
rect 52 548 406 551
rect 52 520 89 548
rect 117 520 175 548
rect 203 520 261 548
rect 289 520 347 548
rect 375 520 406 548
rect 52 517 406 520
rect 450 548 804 551
rect 450 520 487 548
rect 515 520 573 548
rect 601 520 659 548
rect 687 520 745 548
rect 773 520 804 548
rect 450 517 804 520
rect 848 548 1202 551
rect 848 520 885 548
rect 913 520 971 548
rect 999 520 1057 548
rect 1085 520 1143 548
rect 1171 520 1202 548
rect 848 517 1202 520
rect 1246 548 1600 551
rect 1246 520 1283 548
rect 1311 520 1369 548
rect 1397 520 1455 548
rect 1483 520 1541 548
rect 1569 520 1600 548
rect 1246 517 1600 520
rect 1644 548 1998 551
rect 1644 520 1681 548
rect 1709 520 1767 548
rect 1795 520 1853 548
rect 1881 520 1939 548
rect 1967 520 1998 548
rect 1644 517 1998 520
rect 2042 548 2396 551
rect 2042 520 2079 548
rect 2107 520 2165 548
rect 2193 520 2251 548
rect 2279 520 2337 548
rect 2365 520 2396 548
rect 2042 517 2396 520
rect 2440 548 2794 551
rect 2440 520 2477 548
rect 2505 520 2563 548
rect 2591 520 2649 548
rect 2677 520 2735 548
rect 2763 520 2794 548
rect 2440 517 2794 520
rect 2838 548 3192 551
rect 2838 520 2875 548
rect 2903 520 2961 548
rect 2989 520 3047 548
rect 3075 520 3133 548
rect 3161 520 3192 548
rect 2838 517 3192 520
rect 3236 548 3590 551
rect 3236 520 3273 548
rect 3301 520 3359 548
rect 3387 520 3445 548
rect 3473 520 3531 548
rect 3559 520 3590 548
rect 3236 517 3590 520
rect 3634 548 3988 551
rect 3634 520 3671 548
rect 3699 520 3757 548
rect 3785 520 3843 548
rect 3871 520 3929 548
rect 3957 520 3988 548
rect 3634 517 3988 520
rect 4032 548 4386 551
rect 4032 520 4069 548
rect 4097 520 4155 548
rect 4183 520 4241 548
rect 4269 520 4327 548
rect 4355 520 4386 548
rect 4032 517 4386 520
rect 4430 548 4784 551
rect 4430 520 4467 548
rect 4495 520 4553 548
rect 4581 520 4639 548
rect 4667 520 4725 548
rect 4753 520 4784 548
rect 4430 517 4784 520
rect 4828 548 5182 551
rect 4828 520 4865 548
rect 4893 520 4951 548
rect 4979 520 5037 548
rect 5065 520 5123 548
rect 5151 520 5182 548
rect 4828 517 5182 520
rect 5226 548 5580 551
rect 5226 520 5263 548
rect 5291 520 5349 548
rect 5377 520 5435 548
rect 5463 520 5521 548
rect 5549 520 5580 548
rect 5226 517 5580 520
rect 5624 548 5978 551
rect 5624 520 5661 548
rect 5689 520 5747 548
rect 5775 520 5833 548
rect 5861 520 5919 548
rect 5947 520 5978 548
rect 5624 517 5978 520
rect 6022 548 6376 551
rect 6022 520 6059 548
rect 6087 520 6145 548
rect 6173 520 6231 548
rect 6259 520 6317 548
rect 6345 520 6376 548
rect 6022 517 6376 520
rect 6420 548 6774 551
rect 6420 520 6457 548
rect 6485 520 6543 548
rect 6571 520 6629 548
rect 6657 520 6715 548
rect 6743 520 6774 548
rect 6420 517 6774 520
rect 6818 548 7172 551
rect 6818 520 6855 548
rect 6883 520 6941 548
rect 6969 520 7027 548
rect 7055 520 7113 548
rect 7141 520 7172 548
rect 6818 517 7172 520
rect 7216 548 7570 551
rect 7216 520 7253 548
rect 7281 520 7339 548
rect 7367 520 7425 548
rect 7453 520 7511 548
rect 7539 520 7570 548
rect 7216 517 7570 520
rect 7614 548 7968 551
rect 7614 520 7651 548
rect 7679 520 7737 548
rect 7765 520 7823 548
rect 7851 520 7909 548
rect 7937 520 7968 548
rect 7614 517 7968 520
rect 8012 548 8366 551
rect 8012 520 8049 548
rect 8077 520 8135 548
rect 8163 520 8221 548
rect 8249 520 8307 548
rect 8335 520 8366 548
rect 8012 517 8366 520
rect 8410 548 8764 551
rect 8410 520 8447 548
rect 8475 520 8533 548
rect 8561 520 8619 548
rect 8647 520 8705 548
rect 8733 520 8764 548
rect 8410 517 8764 520
rect 8808 548 9162 551
rect 8808 520 8845 548
rect 8873 520 8931 548
rect 8959 520 9017 548
rect 9045 520 9103 548
rect 9131 520 9162 548
rect 8808 517 9162 520
rect 9206 548 9560 551
rect 9206 520 9243 548
rect 9271 520 9329 548
rect 9357 520 9415 548
rect 9443 520 9501 548
rect 9529 520 9560 548
rect 9206 517 9560 520
rect 9604 548 9958 551
rect 9604 520 9641 548
rect 9669 520 9727 548
rect 9755 520 9813 548
rect 9841 520 9899 548
rect 9927 520 9958 548
rect 9604 517 9958 520
rect 52 372 406 375
rect 52 344 89 372
rect 117 344 175 372
rect 203 344 261 372
rect 289 344 347 372
rect 375 344 406 372
rect 52 341 406 344
rect 450 372 804 375
rect 450 344 487 372
rect 515 344 573 372
rect 601 344 659 372
rect 687 344 745 372
rect 773 344 804 372
rect 450 341 804 344
rect 848 372 1202 375
rect 848 344 885 372
rect 913 344 971 372
rect 999 344 1057 372
rect 1085 344 1143 372
rect 1171 344 1202 372
rect 848 341 1202 344
rect 1246 372 1600 375
rect 1246 344 1283 372
rect 1311 344 1369 372
rect 1397 344 1455 372
rect 1483 344 1541 372
rect 1569 344 1600 372
rect 1246 341 1600 344
rect 1644 372 1998 375
rect 1644 344 1681 372
rect 1709 344 1767 372
rect 1795 344 1853 372
rect 1881 344 1939 372
rect 1967 344 1998 372
rect 1644 341 1998 344
rect 2042 372 2396 375
rect 2042 344 2079 372
rect 2107 344 2165 372
rect 2193 344 2251 372
rect 2279 344 2337 372
rect 2365 344 2396 372
rect 2042 341 2396 344
rect 2440 372 2794 375
rect 2440 344 2477 372
rect 2505 344 2563 372
rect 2591 344 2649 372
rect 2677 344 2735 372
rect 2763 344 2794 372
rect 2440 341 2794 344
rect 2838 372 3192 375
rect 2838 344 2875 372
rect 2903 344 2961 372
rect 2989 344 3047 372
rect 3075 344 3133 372
rect 3161 344 3192 372
rect 2838 341 3192 344
rect 3236 372 3590 375
rect 3236 344 3273 372
rect 3301 344 3359 372
rect 3387 344 3445 372
rect 3473 344 3531 372
rect 3559 344 3590 372
rect 3236 341 3590 344
rect 3634 372 3988 375
rect 3634 344 3671 372
rect 3699 344 3757 372
rect 3785 344 3843 372
rect 3871 344 3929 372
rect 3957 344 3988 372
rect 3634 341 3988 344
rect 4032 372 4386 375
rect 4032 344 4069 372
rect 4097 344 4155 372
rect 4183 344 4241 372
rect 4269 344 4327 372
rect 4355 344 4386 372
rect 4032 341 4386 344
rect 4430 372 4784 375
rect 4430 344 4467 372
rect 4495 344 4553 372
rect 4581 344 4639 372
rect 4667 344 4725 372
rect 4753 344 4784 372
rect 4430 341 4784 344
rect 4828 372 5182 375
rect 4828 344 4865 372
rect 4893 344 4951 372
rect 4979 344 5037 372
rect 5065 344 5123 372
rect 5151 344 5182 372
rect 4828 341 5182 344
rect 5226 372 5580 375
rect 5226 344 5263 372
rect 5291 344 5349 372
rect 5377 344 5435 372
rect 5463 344 5521 372
rect 5549 344 5580 372
rect 5226 341 5580 344
rect 5624 372 5978 375
rect 5624 344 5661 372
rect 5689 344 5747 372
rect 5775 344 5833 372
rect 5861 344 5919 372
rect 5947 344 5978 372
rect 5624 341 5978 344
rect 6022 372 6376 375
rect 6022 344 6059 372
rect 6087 344 6145 372
rect 6173 344 6231 372
rect 6259 344 6317 372
rect 6345 344 6376 372
rect 6022 341 6376 344
rect 6420 372 6774 375
rect 6420 344 6457 372
rect 6485 344 6543 372
rect 6571 344 6629 372
rect 6657 344 6715 372
rect 6743 344 6774 372
rect 6420 341 6774 344
rect 6818 372 7172 375
rect 6818 344 6855 372
rect 6883 344 6941 372
rect 6969 344 7027 372
rect 7055 344 7113 372
rect 7141 344 7172 372
rect 6818 341 7172 344
rect 7216 372 7570 375
rect 7216 344 7253 372
rect 7281 344 7339 372
rect 7367 344 7425 372
rect 7453 344 7511 372
rect 7539 344 7570 372
rect 7216 341 7570 344
rect 7614 372 7968 375
rect 7614 344 7651 372
rect 7679 344 7737 372
rect 7765 344 7823 372
rect 7851 344 7909 372
rect 7937 344 7968 372
rect 7614 341 7968 344
rect 8012 372 8366 375
rect 8012 344 8049 372
rect 8077 344 8135 372
rect 8163 344 8221 372
rect 8249 344 8307 372
rect 8335 344 8366 372
rect 8012 341 8366 344
rect 8410 372 8764 375
rect 8410 344 8447 372
rect 8475 344 8533 372
rect 8561 344 8619 372
rect 8647 344 8705 372
rect 8733 344 8764 372
rect 8410 341 8764 344
rect 8808 372 9162 375
rect 8808 344 8845 372
rect 8873 344 8931 372
rect 8959 344 9017 372
rect 9045 344 9103 372
rect 9131 344 9162 372
rect 8808 341 9162 344
rect 9206 372 9560 375
rect 9206 344 9243 372
rect 9271 344 9329 372
rect 9357 344 9415 372
rect 9443 344 9501 372
rect 9529 344 9560 372
rect 9206 341 9560 344
rect 9604 372 9958 375
rect 9604 344 9641 372
rect 9669 344 9727 372
rect 9755 344 9813 372
rect 9841 344 9899 372
rect 9927 344 9958 372
rect 9604 341 9958 344
rect 52 286 406 289
rect 52 258 89 286
rect 117 258 175 286
rect 203 258 261 286
rect 289 258 347 286
rect 375 258 406 286
rect 52 255 406 258
rect 450 286 804 289
rect 450 258 487 286
rect 515 258 573 286
rect 601 258 659 286
rect 687 258 745 286
rect 773 258 804 286
rect 450 255 804 258
rect 848 286 1202 289
rect 848 258 885 286
rect 913 258 971 286
rect 999 258 1057 286
rect 1085 258 1143 286
rect 1171 258 1202 286
rect 848 255 1202 258
rect 1246 286 1600 289
rect 1246 258 1283 286
rect 1311 258 1369 286
rect 1397 258 1455 286
rect 1483 258 1541 286
rect 1569 258 1600 286
rect 1246 255 1600 258
rect 1644 286 1998 289
rect 1644 258 1681 286
rect 1709 258 1767 286
rect 1795 258 1853 286
rect 1881 258 1939 286
rect 1967 258 1998 286
rect 1644 255 1998 258
rect 2042 286 2396 289
rect 2042 258 2079 286
rect 2107 258 2165 286
rect 2193 258 2251 286
rect 2279 258 2337 286
rect 2365 258 2396 286
rect 2042 255 2396 258
rect 2440 286 2794 289
rect 2440 258 2477 286
rect 2505 258 2563 286
rect 2591 258 2649 286
rect 2677 258 2735 286
rect 2763 258 2794 286
rect 2440 255 2794 258
rect 2838 286 3192 289
rect 2838 258 2875 286
rect 2903 258 2961 286
rect 2989 258 3047 286
rect 3075 258 3133 286
rect 3161 258 3192 286
rect 2838 255 3192 258
rect 3236 286 3590 289
rect 3236 258 3273 286
rect 3301 258 3359 286
rect 3387 258 3445 286
rect 3473 258 3531 286
rect 3559 258 3590 286
rect 3236 255 3590 258
rect 3634 286 3988 289
rect 3634 258 3671 286
rect 3699 258 3757 286
rect 3785 258 3843 286
rect 3871 258 3929 286
rect 3957 258 3988 286
rect 3634 255 3988 258
rect 4032 286 4386 289
rect 4032 258 4069 286
rect 4097 258 4155 286
rect 4183 258 4241 286
rect 4269 258 4327 286
rect 4355 258 4386 286
rect 4032 255 4386 258
rect 4430 286 4784 289
rect 4430 258 4467 286
rect 4495 258 4553 286
rect 4581 258 4639 286
rect 4667 258 4725 286
rect 4753 258 4784 286
rect 4430 255 4784 258
rect 4828 286 5182 289
rect 4828 258 4865 286
rect 4893 258 4951 286
rect 4979 258 5037 286
rect 5065 258 5123 286
rect 5151 258 5182 286
rect 4828 255 5182 258
rect 5226 286 5580 289
rect 5226 258 5263 286
rect 5291 258 5349 286
rect 5377 258 5435 286
rect 5463 258 5521 286
rect 5549 258 5580 286
rect 5226 255 5580 258
rect 5624 286 5978 289
rect 5624 258 5661 286
rect 5689 258 5747 286
rect 5775 258 5833 286
rect 5861 258 5919 286
rect 5947 258 5978 286
rect 5624 255 5978 258
rect 6022 286 6376 289
rect 6022 258 6059 286
rect 6087 258 6145 286
rect 6173 258 6231 286
rect 6259 258 6317 286
rect 6345 258 6376 286
rect 6022 255 6376 258
rect 6420 286 6774 289
rect 6420 258 6457 286
rect 6485 258 6543 286
rect 6571 258 6629 286
rect 6657 258 6715 286
rect 6743 258 6774 286
rect 6420 255 6774 258
rect 6818 286 7172 289
rect 6818 258 6855 286
rect 6883 258 6941 286
rect 6969 258 7027 286
rect 7055 258 7113 286
rect 7141 258 7172 286
rect 6818 255 7172 258
rect 7216 286 7570 289
rect 7216 258 7253 286
rect 7281 258 7339 286
rect 7367 258 7425 286
rect 7453 258 7511 286
rect 7539 258 7570 286
rect 7216 255 7570 258
rect 7614 286 7968 289
rect 7614 258 7651 286
rect 7679 258 7737 286
rect 7765 258 7823 286
rect 7851 258 7909 286
rect 7937 258 7968 286
rect 7614 255 7968 258
rect 8012 286 8366 289
rect 8012 258 8049 286
rect 8077 258 8135 286
rect 8163 258 8221 286
rect 8249 258 8307 286
rect 8335 258 8366 286
rect 8012 255 8366 258
rect 8410 286 8764 289
rect 8410 258 8447 286
rect 8475 258 8533 286
rect 8561 258 8619 286
rect 8647 258 8705 286
rect 8733 258 8764 286
rect 8410 255 8764 258
rect 8808 286 9162 289
rect 8808 258 8845 286
rect 8873 258 8931 286
rect 8959 258 9017 286
rect 9045 258 9103 286
rect 9131 258 9162 286
rect 8808 255 9162 258
rect 9206 286 9560 289
rect 9206 258 9243 286
rect 9271 258 9329 286
rect 9357 258 9415 286
rect 9443 258 9501 286
rect 9529 258 9560 286
rect 9206 255 9560 258
rect 9604 286 9958 289
rect 9604 258 9641 286
rect 9669 258 9727 286
rect 9755 258 9813 286
rect 9841 258 9899 286
rect 9927 258 9958 286
rect 9604 255 9958 258
rect 52 200 406 203
rect 52 172 89 200
rect 117 172 175 200
rect 203 172 261 200
rect 289 172 347 200
rect 375 172 406 200
rect 52 169 406 172
rect 450 200 804 203
rect 450 172 487 200
rect 515 172 573 200
rect 601 172 659 200
rect 687 172 745 200
rect 773 172 804 200
rect 450 169 804 172
rect 848 200 1202 203
rect 848 172 885 200
rect 913 172 971 200
rect 999 172 1057 200
rect 1085 172 1143 200
rect 1171 172 1202 200
rect 848 169 1202 172
rect 1246 200 1600 203
rect 1246 172 1283 200
rect 1311 172 1369 200
rect 1397 172 1455 200
rect 1483 172 1541 200
rect 1569 172 1600 200
rect 1246 169 1600 172
rect 1644 200 1998 203
rect 1644 172 1681 200
rect 1709 172 1767 200
rect 1795 172 1853 200
rect 1881 172 1939 200
rect 1967 172 1998 200
rect 1644 169 1998 172
rect 2042 200 2396 203
rect 2042 172 2079 200
rect 2107 172 2165 200
rect 2193 172 2251 200
rect 2279 172 2337 200
rect 2365 172 2396 200
rect 2042 169 2396 172
rect 2440 200 2794 203
rect 2440 172 2477 200
rect 2505 172 2563 200
rect 2591 172 2649 200
rect 2677 172 2735 200
rect 2763 172 2794 200
rect 2440 169 2794 172
rect 2838 200 3192 203
rect 2838 172 2875 200
rect 2903 172 2961 200
rect 2989 172 3047 200
rect 3075 172 3133 200
rect 3161 172 3192 200
rect 2838 169 3192 172
rect 3236 200 3590 203
rect 3236 172 3273 200
rect 3301 172 3359 200
rect 3387 172 3445 200
rect 3473 172 3531 200
rect 3559 172 3590 200
rect 3236 169 3590 172
rect 3634 200 3988 203
rect 3634 172 3671 200
rect 3699 172 3757 200
rect 3785 172 3843 200
rect 3871 172 3929 200
rect 3957 172 3988 200
rect 3634 169 3988 172
rect 4032 200 4386 203
rect 4032 172 4069 200
rect 4097 172 4155 200
rect 4183 172 4241 200
rect 4269 172 4327 200
rect 4355 172 4386 200
rect 4032 169 4386 172
rect 4430 200 4784 203
rect 4430 172 4467 200
rect 4495 172 4553 200
rect 4581 172 4639 200
rect 4667 172 4725 200
rect 4753 172 4784 200
rect 4430 169 4784 172
rect 4828 200 5182 203
rect 4828 172 4865 200
rect 4893 172 4951 200
rect 4979 172 5037 200
rect 5065 172 5123 200
rect 5151 172 5182 200
rect 4828 169 5182 172
rect 5226 200 5580 203
rect 5226 172 5263 200
rect 5291 172 5349 200
rect 5377 172 5435 200
rect 5463 172 5521 200
rect 5549 172 5580 200
rect 5226 169 5580 172
rect 5624 200 5978 203
rect 5624 172 5661 200
rect 5689 172 5747 200
rect 5775 172 5833 200
rect 5861 172 5919 200
rect 5947 172 5978 200
rect 5624 169 5978 172
rect 6022 200 6376 203
rect 6022 172 6059 200
rect 6087 172 6145 200
rect 6173 172 6231 200
rect 6259 172 6317 200
rect 6345 172 6376 200
rect 6022 169 6376 172
rect 6420 200 6774 203
rect 6420 172 6457 200
rect 6485 172 6543 200
rect 6571 172 6629 200
rect 6657 172 6715 200
rect 6743 172 6774 200
rect 6420 169 6774 172
rect 6818 200 7172 203
rect 6818 172 6855 200
rect 6883 172 6941 200
rect 6969 172 7027 200
rect 7055 172 7113 200
rect 7141 172 7172 200
rect 6818 169 7172 172
rect 7216 200 7570 203
rect 7216 172 7253 200
rect 7281 172 7339 200
rect 7367 172 7425 200
rect 7453 172 7511 200
rect 7539 172 7570 200
rect 7216 169 7570 172
rect 7614 200 7968 203
rect 7614 172 7651 200
rect 7679 172 7737 200
rect 7765 172 7823 200
rect 7851 172 7909 200
rect 7937 172 7968 200
rect 7614 169 7968 172
rect 8012 200 8366 203
rect 8012 172 8049 200
rect 8077 172 8135 200
rect 8163 172 8221 200
rect 8249 172 8307 200
rect 8335 172 8366 200
rect 8012 169 8366 172
rect 8410 200 8764 203
rect 8410 172 8447 200
rect 8475 172 8533 200
rect 8561 172 8619 200
rect 8647 172 8705 200
rect 8733 172 8764 200
rect 8410 169 8764 172
rect 8808 200 9162 203
rect 8808 172 8845 200
rect 8873 172 8931 200
rect 8959 172 9017 200
rect 9045 172 9103 200
rect 9131 172 9162 200
rect 8808 169 9162 172
rect 9206 200 9560 203
rect 9206 172 9243 200
rect 9271 172 9329 200
rect 9357 172 9415 200
rect 9443 172 9501 200
rect 9529 172 9560 200
rect 9206 169 9560 172
rect 9604 200 9958 203
rect 9604 172 9641 200
rect 9669 172 9727 200
rect 9755 172 9813 200
rect 9841 172 9899 200
rect 9927 172 9958 200
rect 9604 169 9958 172
rect 52 114 406 117
rect 52 86 89 114
rect 117 86 175 114
rect 203 86 261 114
rect 289 86 347 114
rect 375 86 406 114
rect 52 83 406 86
rect 450 114 804 117
rect 450 86 487 114
rect 515 86 573 114
rect 601 86 659 114
rect 687 86 745 114
rect 773 86 804 114
rect 450 83 804 86
rect 848 114 1202 117
rect 848 86 885 114
rect 913 86 971 114
rect 999 86 1057 114
rect 1085 86 1143 114
rect 1171 86 1202 114
rect 848 83 1202 86
rect 1246 114 1600 117
rect 1246 86 1283 114
rect 1311 86 1369 114
rect 1397 86 1455 114
rect 1483 86 1541 114
rect 1569 86 1600 114
rect 1246 83 1600 86
rect 1644 114 1998 117
rect 1644 86 1681 114
rect 1709 86 1767 114
rect 1795 86 1853 114
rect 1881 86 1939 114
rect 1967 86 1998 114
rect 1644 83 1998 86
rect 2042 114 2396 117
rect 2042 86 2079 114
rect 2107 86 2165 114
rect 2193 86 2251 114
rect 2279 86 2337 114
rect 2365 86 2396 114
rect 2042 83 2396 86
rect 2440 114 2794 117
rect 2440 86 2477 114
rect 2505 86 2563 114
rect 2591 86 2649 114
rect 2677 86 2735 114
rect 2763 86 2794 114
rect 2440 83 2794 86
rect 2838 114 3192 117
rect 2838 86 2875 114
rect 2903 86 2961 114
rect 2989 86 3047 114
rect 3075 86 3133 114
rect 3161 86 3192 114
rect 2838 83 3192 86
rect 3236 114 3590 117
rect 3236 86 3273 114
rect 3301 86 3359 114
rect 3387 86 3445 114
rect 3473 86 3531 114
rect 3559 86 3590 114
rect 3236 83 3590 86
rect 3634 114 3988 117
rect 3634 86 3671 114
rect 3699 86 3757 114
rect 3785 86 3843 114
rect 3871 86 3929 114
rect 3957 86 3988 114
rect 3634 83 3988 86
rect 4032 114 4386 117
rect 4032 86 4069 114
rect 4097 86 4155 114
rect 4183 86 4241 114
rect 4269 86 4327 114
rect 4355 86 4386 114
rect 4032 83 4386 86
rect 4430 114 4784 117
rect 4430 86 4467 114
rect 4495 86 4553 114
rect 4581 86 4639 114
rect 4667 86 4725 114
rect 4753 86 4784 114
rect 4430 83 4784 86
rect 4828 114 5182 117
rect 4828 86 4865 114
rect 4893 86 4951 114
rect 4979 86 5037 114
rect 5065 86 5123 114
rect 5151 86 5182 114
rect 4828 83 5182 86
rect 5226 114 5580 117
rect 5226 86 5263 114
rect 5291 86 5349 114
rect 5377 86 5435 114
rect 5463 86 5521 114
rect 5549 86 5580 114
rect 5226 83 5580 86
rect 5624 114 5978 117
rect 5624 86 5661 114
rect 5689 86 5747 114
rect 5775 86 5833 114
rect 5861 86 5919 114
rect 5947 86 5978 114
rect 5624 83 5978 86
rect 6022 114 6376 117
rect 6022 86 6059 114
rect 6087 86 6145 114
rect 6173 86 6231 114
rect 6259 86 6317 114
rect 6345 86 6376 114
rect 6022 83 6376 86
rect 6420 114 6774 117
rect 6420 86 6457 114
rect 6485 86 6543 114
rect 6571 86 6629 114
rect 6657 86 6715 114
rect 6743 86 6774 114
rect 6420 83 6774 86
rect 6818 114 7172 117
rect 6818 86 6855 114
rect 6883 86 6941 114
rect 6969 86 7027 114
rect 7055 86 7113 114
rect 7141 86 7172 114
rect 6818 83 7172 86
rect 7216 114 7570 117
rect 7216 86 7253 114
rect 7281 86 7339 114
rect 7367 86 7425 114
rect 7453 86 7511 114
rect 7539 86 7570 114
rect 7216 83 7570 86
rect 7614 114 7968 117
rect 7614 86 7651 114
rect 7679 86 7737 114
rect 7765 86 7823 114
rect 7851 86 7909 114
rect 7937 86 7968 114
rect 7614 83 7968 86
rect 8012 114 8366 117
rect 8012 86 8049 114
rect 8077 86 8135 114
rect 8163 86 8221 114
rect 8249 86 8307 114
rect 8335 86 8366 114
rect 8012 83 8366 86
rect 8410 114 8764 117
rect 8410 86 8447 114
rect 8475 86 8533 114
rect 8561 86 8619 114
rect 8647 86 8705 114
rect 8733 86 8764 114
rect 8410 83 8764 86
rect 8808 114 9162 117
rect 8808 86 8845 114
rect 8873 86 8931 114
rect 8959 86 9017 114
rect 9045 86 9103 114
rect 9131 86 9162 114
rect 8808 83 9162 86
rect 9206 114 9560 117
rect 9206 86 9243 114
rect 9271 86 9329 114
rect 9357 86 9415 114
rect 9443 86 9501 114
rect 9529 86 9560 114
rect 9206 83 9560 86
rect 9604 114 9958 117
rect 9604 86 9641 114
rect 9669 86 9727 114
rect 9755 86 9813 114
rect 9841 86 9899 114
rect 9927 86 9958 114
rect 9604 83 9958 86
<< metal4 >>
rect 0 1736 413 1766
rect 443 1736 1607 1766
rect 1637 1736 2403 1766
rect 2433 1736 3597 1766
rect 3627 1736 4393 1766
rect 4423 1736 5587 1766
rect 5617 1736 6383 1766
rect 6413 1736 7577 1766
rect 7607 1736 8373 1766
rect 8403 1736 9567 1766
rect 9597 1736 10010 1766
rect 0 1332 30 1736
rect 86 1677 120 1736
rect 172 1677 206 1736
rect 258 1677 292 1736
rect 344 1677 378 1736
rect 484 1677 518 1736
rect 570 1677 604 1736
rect 656 1677 690 1736
rect 742 1677 776 1736
rect 882 1677 916 1736
rect 968 1677 1002 1736
rect 1054 1677 1088 1736
rect 1140 1677 1174 1736
rect 1280 1677 1314 1736
rect 1366 1677 1400 1736
rect 1452 1677 1486 1736
rect 1538 1677 1572 1736
rect 1678 1677 1712 1736
rect 1764 1677 1798 1736
rect 1850 1677 1884 1736
rect 1936 1677 1970 1736
rect 2076 1677 2110 1736
rect 2162 1677 2196 1736
rect 2248 1677 2282 1736
rect 2334 1677 2368 1736
rect 2474 1677 2508 1736
rect 2560 1677 2594 1736
rect 2646 1677 2680 1736
rect 2732 1677 2766 1736
rect 2872 1677 2906 1736
rect 2958 1677 2992 1736
rect 3044 1677 3078 1736
rect 3130 1677 3164 1736
rect 3270 1677 3304 1736
rect 3356 1677 3390 1736
rect 3442 1677 3476 1736
rect 3528 1677 3562 1736
rect 3668 1677 3702 1736
rect 3754 1677 3788 1736
rect 3840 1677 3874 1736
rect 3926 1677 3960 1736
rect 4066 1677 4100 1736
rect 4152 1677 4186 1736
rect 4238 1677 4272 1736
rect 4324 1677 4358 1736
rect 4464 1677 4498 1736
rect 4550 1677 4584 1736
rect 4636 1677 4670 1736
rect 4722 1677 4756 1736
rect 4862 1677 4896 1736
rect 4948 1677 4982 1736
rect 5034 1677 5068 1736
rect 5120 1677 5154 1736
rect 5260 1677 5294 1736
rect 5346 1677 5380 1736
rect 5432 1677 5466 1736
rect 5518 1677 5552 1736
rect 5658 1677 5692 1736
rect 5744 1677 5778 1736
rect 5830 1677 5864 1736
rect 5916 1677 5950 1736
rect 6056 1677 6090 1736
rect 6142 1677 6176 1736
rect 6228 1677 6262 1736
rect 6314 1677 6348 1736
rect 6454 1677 6488 1736
rect 6540 1677 6574 1736
rect 6626 1677 6660 1736
rect 6712 1677 6746 1736
rect 6852 1677 6886 1736
rect 6938 1677 6972 1736
rect 7024 1677 7058 1736
rect 7110 1677 7144 1736
rect 7250 1677 7284 1736
rect 7336 1677 7370 1736
rect 7422 1677 7456 1736
rect 7508 1677 7542 1736
rect 7648 1677 7682 1736
rect 7734 1677 7768 1736
rect 7820 1677 7854 1736
rect 7906 1677 7940 1736
rect 8046 1677 8080 1736
rect 8132 1677 8166 1736
rect 8218 1677 8252 1736
rect 8304 1677 8338 1736
rect 8444 1677 8478 1736
rect 8530 1677 8564 1736
rect 8616 1677 8650 1736
rect 8702 1677 8736 1736
rect 8842 1677 8876 1736
rect 8928 1677 8962 1736
rect 9014 1677 9048 1736
rect 9100 1677 9134 1736
rect 9240 1677 9274 1736
rect 9326 1677 9360 1736
rect 9412 1677 9446 1736
rect 9498 1677 9532 1736
rect 9638 1677 9672 1736
rect 9724 1677 9758 1736
rect 9810 1677 9844 1736
rect 9896 1677 9930 1736
rect 75 1643 131 1677
rect 161 1643 217 1677
rect 247 1643 303 1677
rect 333 1643 389 1677
rect 473 1643 529 1677
rect 559 1643 615 1677
rect 645 1643 701 1677
rect 731 1643 787 1677
rect 871 1643 927 1677
rect 957 1643 1013 1677
rect 1043 1643 1099 1677
rect 1129 1643 1185 1677
rect 1269 1643 1325 1677
rect 1355 1643 1411 1677
rect 1441 1643 1497 1677
rect 1527 1643 1583 1677
rect 1667 1643 1723 1677
rect 1753 1643 1809 1677
rect 1839 1643 1895 1677
rect 1925 1643 1981 1677
rect 2065 1643 2121 1677
rect 2151 1643 2207 1677
rect 2237 1643 2293 1677
rect 2323 1643 2379 1677
rect 2463 1643 2519 1677
rect 2549 1643 2605 1677
rect 2635 1643 2691 1677
rect 2721 1643 2777 1677
rect 2861 1643 2917 1677
rect 2947 1643 3003 1677
rect 3033 1643 3089 1677
rect 3119 1643 3175 1677
rect 3259 1643 3315 1677
rect 3345 1643 3401 1677
rect 3431 1643 3487 1677
rect 3517 1643 3573 1677
rect 3657 1643 3713 1677
rect 3743 1643 3799 1677
rect 3829 1643 3885 1677
rect 3915 1643 3971 1677
rect 4055 1643 4111 1677
rect 4141 1643 4197 1677
rect 4227 1643 4283 1677
rect 4313 1643 4369 1677
rect 4453 1643 4509 1677
rect 4539 1643 4595 1677
rect 4625 1643 4681 1677
rect 4711 1643 4767 1677
rect 4851 1643 4907 1677
rect 4937 1643 4993 1677
rect 5023 1643 5079 1677
rect 5109 1643 5165 1677
rect 5249 1643 5305 1677
rect 5335 1643 5391 1677
rect 5421 1643 5477 1677
rect 5507 1643 5563 1677
rect 5647 1643 5703 1677
rect 5733 1643 5789 1677
rect 5819 1643 5875 1677
rect 5905 1643 5961 1677
rect 6045 1643 6101 1677
rect 6131 1643 6187 1677
rect 6217 1643 6273 1677
rect 6303 1643 6359 1677
rect 6443 1643 6499 1677
rect 6529 1643 6585 1677
rect 6615 1643 6671 1677
rect 6701 1643 6757 1677
rect 6841 1643 6897 1677
rect 6927 1643 6983 1677
rect 7013 1643 7069 1677
rect 7099 1643 7155 1677
rect 7239 1643 7295 1677
rect 7325 1643 7381 1677
rect 7411 1643 7467 1677
rect 7497 1643 7553 1677
rect 7637 1643 7693 1677
rect 7723 1643 7779 1677
rect 7809 1643 7865 1677
rect 7895 1643 7951 1677
rect 8035 1643 8091 1677
rect 8121 1643 8177 1677
rect 8207 1643 8263 1677
rect 8293 1643 8349 1677
rect 8433 1643 8489 1677
rect 8519 1643 8575 1677
rect 8605 1643 8661 1677
rect 8691 1643 8747 1677
rect 8831 1643 8887 1677
rect 8917 1643 8973 1677
rect 9003 1643 9059 1677
rect 9089 1643 9145 1677
rect 9229 1643 9285 1677
rect 9315 1643 9371 1677
rect 9401 1643 9457 1677
rect 9487 1643 9543 1677
rect 9627 1643 9683 1677
rect 9713 1643 9769 1677
rect 9799 1643 9855 1677
rect 9885 1643 9941 1677
rect 86 1591 120 1643
rect 172 1591 206 1643
rect 258 1591 292 1643
rect 344 1591 378 1643
rect 484 1591 518 1643
rect 570 1591 604 1643
rect 656 1591 690 1643
rect 742 1591 776 1643
rect 882 1591 916 1643
rect 968 1591 1002 1643
rect 1054 1591 1088 1643
rect 1140 1591 1174 1643
rect 1280 1591 1314 1643
rect 1366 1591 1400 1643
rect 1452 1591 1486 1643
rect 1538 1591 1572 1643
rect 1678 1591 1712 1643
rect 1764 1591 1798 1643
rect 1850 1591 1884 1643
rect 1936 1591 1970 1643
rect 2076 1591 2110 1643
rect 2162 1591 2196 1643
rect 2248 1591 2282 1643
rect 2334 1591 2368 1643
rect 2474 1591 2508 1643
rect 2560 1591 2594 1643
rect 2646 1591 2680 1643
rect 2732 1591 2766 1643
rect 2872 1591 2906 1643
rect 2958 1591 2992 1643
rect 3044 1591 3078 1643
rect 3130 1591 3164 1643
rect 3270 1591 3304 1643
rect 3356 1591 3390 1643
rect 3442 1591 3476 1643
rect 3528 1591 3562 1643
rect 3668 1591 3702 1643
rect 3754 1591 3788 1643
rect 3840 1591 3874 1643
rect 3926 1591 3960 1643
rect 4066 1591 4100 1643
rect 4152 1591 4186 1643
rect 4238 1591 4272 1643
rect 4324 1591 4358 1643
rect 4464 1591 4498 1643
rect 4550 1591 4584 1643
rect 4636 1591 4670 1643
rect 4722 1591 4756 1643
rect 4862 1591 4896 1643
rect 4948 1591 4982 1643
rect 5034 1591 5068 1643
rect 5120 1591 5154 1643
rect 5260 1591 5294 1643
rect 5346 1591 5380 1643
rect 5432 1591 5466 1643
rect 5518 1591 5552 1643
rect 5658 1591 5692 1643
rect 5744 1591 5778 1643
rect 5830 1591 5864 1643
rect 5916 1591 5950 1643
rect 6056 1591 6090 1643
rect 6142 1591 6176 1643
rect 6228 1591 6262 1643
rect 6314 1591 6348 1643
rect 6454 1591 6488 1643
rect 6540 1591 6574 1643
rect 6626 1591 6660 1643
rect 6712 1591 6746 1643
rect 6852 1591 6886 1643
rect 6938 1591 6972 1643
rect 7024 1591 7058 1643
rect 7110 1591 7144 1643
rect 7250 1591 7284 1643
rect 7336 1591 7370 1643
rect 7422 1591 7456 1643
rect 7508 1591 7542 1643
rect 7648 1591 7682 1643
rect 7734 1591 7768 1643
rect 7820 1591 7854 1643
rect 7906 1591 7940 1643
rect 8046 1591 8080 1643
rect 8132 1591 8166 1643
rect 8218 1591 8252 1643
rect 8304 1591 8338 1643
rect 8444 1591 8478 1643
rect 8530 1591 8564 1643
rect 8616 1591 8650 1643
rect 8702 1591 8736 1643
rect 8842 1591 8876 1643
rect 8928 1591 8962 1643
rect 9014 1591 9048 1643
rect 9100 1591 9134 1643
rect 9240 1591 9274 1643
rect 9326 1591 9360 1643
rect 9412 1591 9446 1643
rect 9498 1591 9532 1643
rect 9638 1591 9672 1643
rect 9724 1591 9758 1643
rect 9810 1591 9844 1643
rect 9896 1591 9930 1643
rect 75 1557 131 1591
rect 161 1557 217 1591
rect 247 1557 303 1591
rect 333 1557 389 1591
rect 473 1557 529 1591
rect 559 1557 615 1591
rect 645 1557 701 1591
rect 731 1557 787 1591
rect 871 1557 927 1591
rect 957 1557 1013 1591
rect 1043 1557 1099 1591
rect 1129 1557 1185 1591
rect 1269 1557 1325 1591
rect 1355 1557 1411 1591
rect 1441 1557 1497 1591
rect 1527 1557 1583 1591
rect 1667 1557 1723 1591
rect 1753 1557 1809 1591
rect 1839 1557 1895 1591
rect 1925 1557 1981 1591
rect 2065 1557 2121 1591
rect 2151 1557 2207 1591
rect 2237 1557 2293 1591
rect 2323 1557 2379 1591
rect 2463 1557 2519 1591
rect 2549 1557 2605 1591
rect 2635 1557 2691 1591
rect 2721 1557 2777 1591
rect 2861 1557 2917 1591
rect 2947 1557 3003 1591
rect 3033 1557 3089 1591
rect 3119 1557 3175 1591
rect 3259 1557 3315 1591
rect 3345 1557 3401 1591
rect 3431 1557 3487 1591
rect 3517 1557 3573 1591
rect 3657 1557 3713 1591
rect 3743 1557 3799 1591
rect 3829 1557 3885 1591
rect 3915 1557 3971 1591
rect 4055 1557 4111 1591
rect 4141 1557 4197 1591
rect 4227 1557 4283 1591
rect 4313 1557 4369 1591
rect 4453 1557 4509 1591
rect 4539 1557 4595 1591
rect 4625 1557 4681 1591
rect 4711 1557 4767 1591
rect 4851 1557 4907 1591
rect 4937 1557 4993 1591
rect 5023 1557 5079 1591
rect 5109 1557 5165 1591
rect 5249 1557 5305 1591
rect 5335 1557 5391 1591
rect 5421 1557 5477 1591
rect 5507 1557 5563 1591
rect 5647 1557 5703 1591
rect 5733 1557 5789 1591
rect 5819 1557 5875 1591
rect 5905 1557 5961 1591
rect 6045 1557 6101 1591
rect 6131 1557 6187 1591
rect 6217 1557 6273 1591
rect 6303 1557 6359 1591
rect 6443 1557 6499 1591
rect 6529 1557 6585 1591
rect 6615 1557 6671 1591
rect 6701 1557 6757 1591
rect 6841 1557 6897 1591
rect 6927 1557 6983 1591
rect 7013 1557 7069 1591
rect 7099 1557 7155 1591
rect 7239 1557 7295 1591
rect 7325 1557 7381 1591
rect 7411 1557 7467 1591
rect 7497 1557 7553 1591
rect 7637 1557 7693 1591
rect 7723 1557 7779 1591
rect 7809 1557 7865 1591
rect 7895 1557 7951 1591
rect 8035 1557 8091 1591
rect 8121 1557 8177 1591
rect 8207 1557 8263 1591
rect 8293 1557 8349 1591
rect 8433 1557 8489 1591
rect 8519 1557 8575 1591
rect 8605 1557 8661 1591
rect 8691 1557 8747 1591
rect 8831 1557 8887 1591
rect 8917 1557 8973 1591
rect 9003 1557 9059 1591
rect 9089 1557 9145 1591
rect 9229 1557 9285 1591
rect 9315 1557 9371 1591
rect 9401 1557 9457 1591
rect 9487 1557 9543 1591
rect 9627 1557 9683 1591
rect 9713 1557 9769 1591
rect 9799 1557 9855 1591
rect 9885 1557 9941 1591
rect 86 1505 120 1557
rect 172 1505 206 1557
rect 258 1505 292 1557
rect 344 1505 378 1557
rect 484 1505 518 1557
rect 570 1505 604 1557
rect 656 1505 690 1557
rect 742 1505 776 1557
rect 882 1505 916 1557
rect 968 1505 1002 1557
rect 1054 1505 1088 1557
rect 1140 1505 1174 1557
rect 1280 1505 1314 1557
rect 1366 1505 1400 1557
rect 1452 1505 1486 1557
rect 1538 1505 1572 1557
rect 1678 1505 1712 1557
rect 1764 1505 1798 1557
rect 1850 1505 1884 1557
rect 1936 1505 1970 1557
rect 2076 1505 2110 1557
rect 2162 1505 2196 1557
rect 2248 1505 2282 1557
rect 2334 1505 2368 1557
rect 2474 1505 2508 1557
rect 2560 1505 2594 1557
rect 2646 1505 2680 1557
rect 2732 1505 2766 1557
rect 2872 1505 2906 1557
rect 2958 1505 2992 1557
rect 3044 1505 3078 1557
rect 3130 1505 3164 1557
rect 3270 1505 3304 1557
rect 3356 1505 3390 1557
rect 3442 1505 3476 1557
rect 3528 1505 3562 1557
rect 3668 1505 3702 1557
rect 3754 1505 3788 1557
rect 3840 1505 3874 1557
rect 3926 1505 3960 1557
rect 4066 1505 4100 1557
rect 4152 1505 4186 1557
rect 4238 1505 4272 1557
rect 4324 1505 4358 1557
rect 4464 1505 4498 1557
rect 4550 1505 4584 1557
rect 4636 1505 4670 1557
rect 4722 1505 4756 1557
rect 4862 1505 4896 1557
rect 4948 1505 4982 1557
rect 5034 1505 5068 1557
rect 5120 1505 5154 1557
rect 5260 1505 5294 1557
rect 5346 1505 5380 1557
rect 5432 1505 5466 1557
rect 5518 1505 5552 1557
rect 5658 1505 5692 1557
rect 5744 1505 5778 1557
rect 5830 1505 5864 1557
rect 5916 1505 5950 1557
rect 6056 1505 6090 1557
rect 6142 1505 6176 1557
rect 6228 1505 6262 1557
rect 6314 1505 6348 1557
rect 6454 1505 6488 1557
rect 6540 1505 6574 1557
rect 6626 1505 6660 1557
rect 6712 1505 6746 1557
rect 6852 1505 6886 1557
rect 6938 1505 6972 1557
rect 7024 1505 7058 1557
rect 7110 1505 7144 1557
rect 7250 1505 7284 1557
rect 7336 1505 7370 1557
rect 7422 1505 7456 1557
rect 7508 1505 7542 1557
rect 7648 1505 7682 1557
rect 7734 1505 7768 1557
rect 7820 1505 7854 1557
rect 7906 1505 7940 1557
rect 8046 1505 8080 1557
rect 8132 1505 8166 1557
rect 8218 1505 8252 1557
rect 8304 1505 8338 1557
rect 8444 1505 8478 1557
rect 8530 1505 8564 1557
rect 8616 1505 8650 1557
rect 8702 1505 8736 1557
rect 8842 1505 8876 1557
rect 8928 1505 8962 1557
rect 9014 1505 9048 1557
rect 9100 1505 9134 1557
rect 9240 1505 9274 1557
rect 9326 1505 9360 1557
rect 9412 1505 9446 1557
rect 9498 1505 9532 1557
rect 9638 1505 9672 1557
rect 9724 1505 9758 1557
rect 9810 1505 9844 1557
rect 9896 1505 9930 1557
rect 75 1471 131 1505
rect 161 1471 217 1505
rect 247 1471 303 1505
rect 333 1471 389 1505
rect 473 1471 529 1505
rect 559 1471 615 1505
rect 645 1471 701 1505
rect 731 1471 787 1505
rect 871 1471 927 1505
rect 957 1471 1013 1505
rect 1043 1471 1099 1505
rect 1129 1471 1185 1505
rect 1269 1471 1325 1505
rect 1355 1471 1411 1505
rect 1441 1471 1497 1505
rect 1527 1471 1583 1505
rect 1667 1471 1723 1505
rect 1753 1471 1809 1505
rect 1839 1471 1895 1505
rect 1925 1471 1981 1505
rect 2065 1471 2121 1505
rect 2151 1471 2207 1505
rect 2237 1471 2293 1505
rect 2323 1471 2379 1505
rect 2463 1471 2519 1505
rect 2549 1471 2605 1505
rect 2635 1471 2691 1505
rect 2721 1471 2777 1505
rect 2861 1471 2917 1505
rect 2947 1471 3003 1505
rect 3033 1471 3089 1505
rect 3119 1471 3175 1505
rect 3259 1471 3315 1505
rect 3345 1471 3401 1505
rect 3431 1471 3487 1505
rect 3517 1471 3573 1505
rect 3657 1471 3713 1505
rect 3743 1471 3799 1505
rect 3829 1471 3885 1505
rect 3915 1471 3971 1505
rect 4055 1471 4111 1505
rect 4141 1471 4197 1505
rect 4227 1471 4283 1505
rect 4313 1471 4369 1505
rect 4453 1471 4509 1505
rect 4539 1471 4595 1505
rect 4625 1471 4681 1505
rect 4711 1471 4767 1505
rect 4851 1471 4907 1505
rect 4937 1471 4993 1505
rect 5023 1471 5079 1505
rect 5109 1471 5165 1505
rect 5249 1471 5305 1505
rect 5335 1471 5391 1505
rect 5421 1471 5477 1505
rect 5507 1471 5563 1505
rect 5647 1471 5703 1505
rect 5733 1471 5789 1505
rect 5819 1471 5875 1505
rect 5905 1471 5961 1505
rect 6045 1471 6101 1505
rect 6131 1471 6187 1505
rect 6217 1471 6273 1505
rect 6303 1471 6359 1505
rect 6443 1471 6499 1505
rect 6529 1471 6585 1505
rect 6615 1471 6671 1505
rect 6701 1471 6757 1505
rect 6841 1471 6897 1505
rect 6927 1471 6983 1505
rect 7013 1471 7069 1505
rect 7099 1471 7155 1505
rect 7239 1471 7295 1505
rect 7325 1471 7381 1505
rect 7411 1471 7467 1505
rect 7497 1471 7553 1505
rect 7637 1471 7693 1505
rect 7723 1471 7779 1505
rect 7809 1471 7865 1505
rect 7895 1471 7951 1505
rect 8035 1471 8091 1505
rect 8121 1471 8177 1505
rect 8207 1471 8263 1505
rect 8293 1471 8349 1505
rect 8433 1471 8489 1505
rect 8519 1471 8575 1505
rect 8605 1471 8661 1505
rect 8691 1471 8747 1505
rect 8831 1471 8887 1505
rect 8917 1471 8973 1505
rect 9003 1471 9059 1505
rect 9089 1471 9145 1505
rect 9229 1471 9285 1505
rect 9315 1471 9371 1505
rect 9401 1471 9457 1505
rect 9487 1471 9543 1505
rect 9627 1471 9683 1505
rect 9713 1471 9769 1505
rect 9799 1471 9855 1505
rect 9885 1471 9941 1505
rect 86 1419 120 1471
rect 172 1419 206 1471
rect 258 1419 292 1471
rect 344 1419 378 1471
rect 484 1419 518 1471
rect 570 1419 604 1471
rect 656 1419 690 1471
rect 742 1419 776 1471
rect 882 1419 916 1471
rect 968 1419 1002 1471
rect 1054 1419 1088 1471
rect 1140 1419 1174 1471
rect 1280 1419 1314 1471
rect 1366 1419 1400 1471
rect 1452 1419 1486 1471
rect 1538 1419 1572 1471
rect 1678 1419 1712 1471
rect 1764 1419 1798 1471
rect 1850 1419 1884 1471
rect 1936 1419 1970 1471
rect 2076 1419 2110 1471
rect 2162 1419 2196 1471
rect 2248 1419 2282 1471
rect 2334 1419 2368 1471
rect 2474 1419 2508 1471
rect 2560 1419 2594 1471
rect 2646 1419 2680 1471
rect 2732 1419 2766 1471
rect 2872 1419 2906 1471
rect 2958 1419 2992 1471
rect 3044 1419 3078 1471
rect 3130 1419 3164 1471
rect 3270 1419 3304 1471
rect 3356 1419 3390 1471
rect 3442 1419 3476 1471
rect 3528 1419 3562 1471
rect 3668 1419 3702 1471
rect 3754 1419 3788 1471
rect 3840 1419 3874 1471
rect 3926 1419 3960 1471
rect 4066 1419 4100 1471
rect 4152 1419 4186 1471
rect 4238 1419 4272 1471
rect 4324 1419 4358 1471
rect 4464 1419 4498 1471
rect 4550 1419 4584 1471
rect 4636 1419 4670 1471
rect 4722 1419 4756 1471
rect 4862 1419 4896 1471
rect 4948 1419 4982 1471
rect 5034 1419 5068 1471
rect 5120 1419 5154 1471
rect 5260 1419 5294 1471
rect 5346 1419 5380 1471
rect 5432 1419 5466 1471
rect 5518 1419 5552 1471
rect 5658 1419 5692 1471
rect 5744 1419 5778 1471
rect 5830 1419 5864 1471
rect 5916 1419 5950 1471
rect 6056 1419 6090 1471
rect 6142 1419 6176 1471
rect 6228 1419 6262 1471
rect 6314 1419 6348 1471
rect 6454 1419 6488 1471
rect 6540 1419 6574 1471
rect 6626 1419 6660 1471
rect 6712 1419 6746 1471
rect 6852 1419 6886 1471
rect 6938 1419 6972 1471
rect 7024 1419 7058 1471
rect 7110 1419 7144 1471
rect 7250 1419 7284 1471
rect 7336 1419 7370 1471
rect 7422 1419 7456 1471
rect 7508 1419 7542 1471
rect 7648 1419 7682 1471
rect 7734 1419 7768 1471
rect 7820 1419 7854 1471
rect 7906 1419 7940 1471
rect 8046 1419 8080 1471
rect 8132 1419 8166 1471
rect 8218 1419 8252 1471
rect 8304 1419 8338 1471
rect 8444 1419 8478 1471
rect 8530 1419 8564 1471
rect 8616 1419 8650 1471
rect 8702 1419 8736 1471
rect 8842 1419 8876 1471
rect 8928 1419 8962 1471
rect 9014 1419 9048 1471
rect 9100 1419 9134 1471
rect 9240 1419 9274 1471
rect 9326 1419 9360 1471
rect 9412 1419 9446 1471
rect 9498 1419 9532 1471
rect 9638 1419 9672 1471
rect 9724 1419 9758 1471
rect 9810 1419 9844 1471
rect 9896 1419 9930 1471
rect 75 1385 131 1419
rect 161 1385 217 1419
rect 247 1385 303 1419
rect 333 1385 389 1419
rect 473 1385 529 1419
rect 559 1385 615 1419
rect 645 1385 701 1419
rect 731 1385 787 1419
rect 871 1385 927 1419
rect 957 1385 1013 1419
rect 1043 1385 1099 1419
rect 1129 1385 1185 1419
rect 1269 1385 1325 1419
rect 1355 1385 1411 1419
rect 1441 1385 1497 1419
rect 1527 1385 1583 1419
rect 1667 1385 1723 1419
rect 1753 1385 1809 1419
rect 1839 1385 1895 1419
rect 1925 1385 1981 1419
rect 2065 1385 2121 1419
rect 2151 1385 2207 1419
rect 2237 1385 2293 1419
rect 2323 1385 2379 1419
rect 2463 1385 2519 1419
rect 2549 1385 2605 1419
rect 2635 1385 2691 1419
rect 2721 1385 2777 1419
rect 2861 1385 2917 1419
rect 2947 1385 3003 1419
rect 3033 1385 3089 1419
rect 3119 1385 3175 1419
rect 3259 1385 3315 1419
rect 3345 1385 3401 1419
rect 3431 1385 3487 1419
rect 3517 1385 3573 1419
rect 3657 1385 3713 1419
rect 3743 1385 3799 1419
rect 3829 1385 3885 1419
rect 3915 1385 3971 1419
rect 4055 1385 4111 1419
rect 4141 1385 4197 1419
rect 4227 1385 4283 1419
rect 4313 1385 4369 1419
rect 4453 1385 4509 1419
rect 4539 1385 4595 1419
rect 4625 1385 4681 1419
rect 4711 1385 4767 1419
rect 4851 1385 4907 1419
rect 4937 1385 4993 1419
rect 5023 1385 5079 1419
rect 5109 1385 5165 1419
rect 5249 1385 5305 1419
rect 5335 1385 5391 1419
rect 5421 1385 5477 1419
rect 5507 1385 5563 1419
rect 5647 1385 5703 1419
rect 5733 1385 5789 1419
rect 5819 1385 5875 1419
rect 5905 1385 5961 1419
rect 6045 1385 6101 1419
rect 6131 1385 6187 1419
rect 6217 1385 6273 1419
rect 6303 1385 6359 1419
rect 6443 1385 6499 1419
rect 6529 1385 6585 1419
rect 6615 1385 6671 1419
rect 6701 1385 6757 1419
rect 6841 1385 6897 1419
rect 6927 1385 6983 1419
rect 7013 1385 7069 1419
rect 7099 1385 7155 1419
rect 7239 1385 7295 1419
rect 7325 1385 7381 1419
rect 7411 1385 7467 1419
rect 7497 1385 7553 1419
rect 7637 1385 7693 1419
rect 7723 1385 7779 1419
rect 7809 1385 7865 1419
rect 7895 1385 7951 1419
rect 8035 1385 8091 1419
rect 8121 1385 8177 1419
rect 8207 1385 8263 1419
rect 8293 1385 8349 1419
rect 8433 1385 8489 1419
rect 8519 1385 8575 1419
rect 8605 1385 8661 1419
rect 8691 1385 8747 1419
rect 8831 1385 8887 1419
rect 8917 1385 8973 1419
rect 9003 1385 9059 1419
rect 9089 1385 9145 1419
rect 9229 1385 9285 1419
rect 9315 1385 9371 1419
rect 9401 1385 9457 1419
rect 9487 1385 9543 1419
rect 9627 1385 9683 1419
rect 9713 1385 9769 1419
rect 9799 1385 9855 1419
rect 9885 1385 9941 1419
rect 86 1332 120 1385
rect 172 1332 206 1385
rect 258 1332 292 1385
rect 344 1332 378 1385
rect 484 1362 518 1385
rect 570 1362 604 1385
rect 656 1362 690 1385
rect 742 1362 776 1385
rect 882 1362 916 1385
rect 968 1362 1002 1385
rect 1054 1362 1088 1385
rect 1140 1362 1174 1385
rect 1280 1362 1314 1385
rect 1366 1362 1400 1385
rect 1452 1362 1486 1385
rect 1538 1362 1572 1385
rect 1678 1332 1712 1385
rect 1764 1332 1798 1385
rect 1850 1332 1884 1385
rect 1936 1332 1970 1385
rect 2076 1332 2110 1385
rect 2162 1332 2196 1385
rect 2248 1332 2282 1385
rect 2334 1332 2368 1385
rect 2474 1362 2508 1385
rect 2560 1362 2594 1385
rect 2646 1362 2680 1385
rect 2732 1362 2766 1385
rect 2872 1362 2906 1385
rect 2958 1362 2992 1385
rect 3044 1362 3078 1385
rect 3130 1362 3164 1385
rect 3270 1362 3304 1385
rect 3356 1362 3390 1385
rect 3442 1362 3476 1385
rect 3528 1362 3562 1385
rect 3668 1332 3702 1385
rect 3754 1332 3788 1385
rect 3840 1332 3874 1385
rect 3926 1332 3960 1385
rect 4066 1332 4100 1385
rect 4152 1332 4186 1385
rect 4238 1332 4272 1385
rect 4324 1332 4358 1385
rect 4464 1362 4498 1385
rect 4550 1362 4584 1385
rect 4636 1362 4670 1385
rect 4722 1362 4756 1385
rect 4862 1362 4896 1385
rect 4948 1362 4982 1385
rect 5034 1362 5068 1385
rect 5120 1362 5154 1385
rect 5260 1362 5294 1385
rect 5346 1362 5380 1385
rect 5432 1362 5466 1385
rect 5518 1362 5552 1385
rect 5658 1332 5692 1385
rect 5744 1332 5778 1385
rect 5830 1332 5864 1385
rect 5916 1332 5950 1385
rect 6056 1332 6090 1385
rect 6142 1332 6176 1385
rect 6228 1332 6262 1385
rect 6314 1332 6348 1385
rect 6454 1362 6488 1385
rect 6540 1362 6574 1385
rect 6626 1362 6660 1385
rect 6712 1362 6746 1385
rect 6852 1362 6886 1385
rect 6938 1362 6972 1385
rect 7024 1362 7058 1385
rect 7110 1362 7144 1385
rect 7250 1362 7284 1385
rect 7336 1362 7370 1385
rect 7422 1362 7456 1385
rect 7508 1362 7542 1385
rect 7648 1332 7682 1385
rect 7734 1332 7768 1385
rect 7820 1332 7854 1385
rect 7906 1332 7940 1385
rect 8046 1332 8080 1385
rect 8132 1332 8166 1385
rect 8218 1332 8252 1385
rect 8304 1332 8338 1385
rect 8444 1362 8478 1385
rect 8530 1362 8564 1385
rect 8616 1362 8650 1385
rect 8702 1362 8736 1385
rect 8842 1362 8876 1385
rect 8928 1362 8962 1385
rect 9014 1362 9048 1385
rect 9100 1362 9134 1385
rect 9240 1362 9274 1385
rect 9326 1362 9360 1385
rect 9412 1362 9446 1385
rect 9498 1362 9532 1385
rect 9638 1332 9672 1385
rect 9724 1332 9758 1385
rect 9810 1332 9844 1385
rect 9896 1332 9930 1385
rect 9980 1332 10010 1736
rect 0 1302 413 1332
rect 443 1302 1607 1332
rect 1637 1302 2403 1332
rect 2433 1302 3597 1332
rect 3627 1302 4393 1332
rect 4423 1302 5587 1332
rect 5617 1302 6383 1332
rect 6413 1302 7577 1332
rect 7607 1302 8373 1332
rect 8403 1302 9567 1332
rect 9597 1302 10010 1332
rect 0 898 30 1302
rect 86 1243 120 1302
rect 172 1243 206 1302
rect 258 1243 292 1302
rect 344 1243 378 1302
rect 484 1243 518 1302
rect 570 1243 604 1302
rect 656 1243 690 1302
rect 742 1243 776 1302
rect 882 1243 916 1302
rect 968 1243 1002 1302
rect 1054 1243 1088 1302
rect 1140 1243 1174 1302
rect 1280 1243 1314 1302
rect 1366 1243 1400 1302
rect 1452 1243 1486 1302
rect 1538 1243 1572 1302
rect 1678 1243 1712 1302
rect 1764 1243 1798 1302
rect 1850 1243 1884 1302
rect 1936 1243 1970 1302
rect 2076 1243 2110 1302
rect 2162 1243 2196 1302
rect 2248 1243 2282 1302
rect 2334 1243 2368 1302
rect 2474 1243 2508 1302
rect 2560 1243 2594 1302
rect 2646 1243 2680 1302
rect 2732 1243 2766 1302
rect 2872 1243 2906 1302
rect 2958 1243 2992 1302
rect 3044 1243 3078 1302
rect 3130 1243 3164 1302
rect 3270 1243 3304 1302
rect 3356 1243 3390 1302
rect 3442 1243 3476 1302
rect 3528 1243 3562 1302
rect 3668 1243 3702 1302
rect 3754 1243 3788 1302
rect 3840 1243 3874 1302
rect 3926 1243 3960 1302
rect 4066 1243 4100 1302
rect 4152 1243 4186 1302
rect 4238 1243 4272 1302
rect 4324 1243 4358 1302
rect 4464 1243 4498 1302
rect 4550 1243 4584 1302
rect 4636 1243 4670 1302
rect 4722 1243 4756 1302
rect 4862 1243 4896 1302
rect 4948 1243 4982 1302
rect 5034 1243 5068 1302
rect 5120 1243 5154 1302
rect 5260 1243 5294 1302
rect 5346 1243 5380 1302
rect 5432 1243 5466 1302
rect 5518 1243 5552 1302
rect 5658 1243 5692 1302
rect 5744 1243 5778 1302
rect 5830 1243 5864 1302
rect 5916 1243 5950 1302
rect 6056 1243 6090 1302
rect 6142 1243 6176 1302
rect 6228 1243 6262 1302
rect 6314 1243 6348 1302
rect 6454 1243 6488 1302
rect 6540 1243 6574 1302
rect 6626 1243 6660 1302
rect 6712 1243 6746 1302
rect 6852 1243 6886 1302
rect 6938 1243 6972 1302
rect 7024 1243 7058 1302
rect 7110 1243 7144 1302
rect 7250 1243 7284 1302
rect 7336 1243 7370 1302
rect 7422 1243 7456 1302
rect 7508 1243 7542 1302
rect 7648 1243 7682 1302
rect 7734 1243 7768 1302
rect 7820 1243 7854 1302
rect 7906 1243 7940 1302
rect 8046 1243 8080 1302
rect 8132 1243 8166 1302
rect 8218 1243 8252 1302
rect 8304 1243 8338 1302
rect 8444 1243 8478 1302
rect 8530 1243 8564 1302
rect 8616 1243 8650 1302
rect 8702 1243 8736 1302
rect 8842 1243 8876 1302
rect 8928 1243 8962 1302
rect 9014 1243 9048 1302
rect 9100 1243 9134 1302
rect 9240 1243 9274 1302
rect 9326 1243 9360 1302
rect 9412 1243 9446 1302
rect 9498 1243 9532 1302
rect 9638 1243 9672 1302
rect 9724 1243 9758 1302
rect 9810 1243 9844 1302
rect 9896 1243 9930 1302
rect 75 1209 131 1243
rect 161 1209 217 1243
rect 247 1209 303 1243
rect 333 1209 389 1243
rect 473 1209 529 1243
rect 559 1209 615 1243
rect 645 1209 701 1243
rect 731 1209 787 1243
rect 871 1209 927 1243
rect 957 1209 1013 1243
rect 1043 1209 1099 1243
rect 1129 1209 1185 1243
rect 1269 1209 1325 1243
rect 1355 1209 1411 1243
rect 1441 1209 1497 1243
rect 1527 1209 1583 1243
rect 1667 1209 1723 1243
rect 1753 1209 1809 1243
rect 1839 1209 1895 1243
rect 1925 1209 1981 1243
rect 2065 1209 2121 1243
rect 2151 1209 2207 1243
rect 2237 1209 2293 1243
rect 2323 1209 2379 1243
rect 2463 1209 2519 1243
rect 2549 1209 2605 1243
rect 2635 1209 2691 1243
rect 2721 1209 2777 1243
rect 2861 1209 2917 1243
rect 2947 1209 3003 1243
rect 3033 1209 3089 1243
rect 3119 1209 3175 1243
rect 3259 1209 3315 1243
rect 3345 1209 3401 1243
rect 3431 1209 3487 1243
rect 3517 1209 3573 1243
rect 3657 1209 3713 1243
rect 3743 1209 3799 1243
rect 3829 1209 3885 1243
rect 3915 1209 3971 1243
rect 4055 1209 4111 1243
rect 4141 1209 4197 1243
rect 4227 1209 4283 1243
rect 4313 1209 4369 1243
rect 4453 1209 4509 1243
rect 4539 1209 4595 1243
rect 4625 1209 4681 1243
rect 4711 1209 4767 1243
rect 4851 1209 4907 1243
rect 4937 1209 4993 1243
rect 5023 1209 5079 1243
rect 5109 1209 5165 1243
rect 5249 1209 5305 1243
rect 5335 1209 5391 1243
rect 5421 1209 5477 1243
rect 5507 1209 5563 1243
rect 5647 1209 5703 1243
rect 5733 1209 5789 1243
rect 5819 1209 5875 1243
rect 5905 1209 5961 1243
rect 6045 1209 6101 1243
rect 6131 1209 6187 1243
rect 6217 1209 6273 1243
rect 6303 1209 6359 1243
rect 6443 1209 6499 1243
rect 6529 1209 6585 1243
rect 6615 1209 6671 1243
rect 6701 1209 6757 1243
rect 6841 1209 6897 1243
rect 6927 1209 6983 1243
rect 7013 1209 7069 1243
rect 7099 1209 7155 1243
rect 7239 1209 7295 1243
rect 7325 1209 7381 1243
rect 7411 1209 7467 1243
rect 7497 1209 7553 1243
rect 7637 1209 7693 1243
rect 7723 1209 7779 1243
rect 7809 1209 7865 1243
rect 7895 1209 7951 1243
rect 8035 1209 8091 1243
rect 8121 1209 8177 1243
rect 8207 1209 8263 1243
rect 8293 1209 8349 1243
rect 8433 1209 8489 1243
rect 8519 1209 8575 1243
rect 8605 1209 8661 1243
rect 8691 1209 8747 1243
rect 8831 1209 8887 1243
rect 8917 1209 8973 1243
rect 9003 1209 9059 1243
rect 9089 1209 9145 1243
rect 9229 1209 9285 1243
rect 9315 1209 9371 1243
rect 9401 1209 9457 1243
rect 9487 1209 9543 1243
rect 9627 1209 9683 1243
rect 9713 1209 9769 1243
rect 9799 1209 9855 1243
rect 9885 1209 9941 1243
rect 86 1157 120 1209
rect 172 1157 206 1209
rect 258 1157 292 1209
rect 344 1157 378 1209
rect 484 1157 518 1209
rect 570 1157 604 1209
rect 656 1157 690 1209
rect 742 1157 776 1209
rect 882 1157 916 1209
rect 968 1157 1002 1209
rect 1054 1157 1088 1209
rect 1140 1157 1174 1209
rect 1280 1157 1314 1209
rect 1366 1157 1400 1209
rect 1452 1157 1486 1209
rect 1538 1157 1572 1209
rect 1678 1157 1712 1209
rect 1764 1157 1798 1209
rect 1850 1157 1884 1209
rect 1936 1157 1970 1209
rect 2076 1157 2110 1209
rect 2162 1157 2196 1209
rect 2248 1157 2282 1209
rect 2334 1157 2368 1209
rect 2474 1157 2508 1209
rect 2560 1157 2594 1209
rect 2646 1157 2680 1209
rect 2732 1157 2766 1209
rect 2872 1157 2906 1209
rect 2958 1157 2992 1209
rect 3044 1157 3078 1209
rect 3130 1157 3164 1209
rect 3270 1157 3304 1209
rect 3356 1157 3390 1209
rect 3442 1157 3476 1209
rect 3528 1157 3562 1209
rect 3668 1157 3702 1209
rect 3754 1157 3788 1209
rect 3840 1157 3874 1209
rect 3926 1157 3960 1209
rect 4066 1157 4100 1209
rect 4152 1157 4186 1209
rect 4238 1157 4272 1209
rect 4324 1157 4358 1209
rect 4464 1157 4498 1209
rect 4550 1157 4584 1209
rect 4636 1157 4670 1209
rect 4722 1157 4756 1209
rect 4862 1157 4896 1209
rect 4948 1157 4982 1209
rect 5034 1157 5068 1209
rect 5120 1157 5154 1209
rect 5260 1157 5294 1209
rect 5346 1157 5380 1209
rect 5432 1157 5466 1209
rect 5518 1157 5552 1209
rect 5658 1157 5692 1209
rect 5744 1157 5778 1209
rect 5830 1157 5864 1209
rect 5916 1157 5950 1209
rect 6056 1157 6090 1209
rect 6142 1157 6176 1209
rect 6228 1157 6262 1209
rect 6314 1157 6348 1209
rect 6454 1157 6488 1209
rect 6540 1157 6574 1209
rect 6626 1157 6660 1209
rect 6712 1157 6746 1209
rect 6852 1157 6886 1209
rect 6938 1157 6972 1209
rect 7024 1157 7058 1209
rect 7110 1157 7144 1209
rect 7250 1157 7284 1209
rect 7336 1157 7370 1209
rect 7422 1157 7456 1209
rect 7508 1157 7542 1209
rect 7648 1157 7682 1209
rect 7734 1157 7768 1209
rect 7820 1157 7854 1209
rect 7906 1157 7940 1209
rect 8046 1157 8080 1209
rect 8132 1157 8166 1209
rect 8218 1157 8252 1209
rect 8304 1157 8338 1209
rect 8444 1157 8478 1209
rect 8530 1157 8564 1209
rect 8616 1157 8650 1209
rect 8702 1157 8736 1209
rect 8842 1157 8876 1209
rect 8928 1157 8962 1209
rect 9014 1157 9048 1209
rect 9100 1157 9134 1209
rect 9240 1157 9274 1209
rect 9326 1157 9360 1209
rect 9412 1157 9446 1209
rect 9498 1157 9532 1209
rect 9638 1157 9672 1209
rect 9724 1157 9758 1209
rect 9810 1157 9844 1209
rect 9896 1157 9930 1209
rect 75 1123 131 1157
rect 161 1123 217 1157
rect 247 1123 303 1157
rect 333 1123 389 1157
rect 473 1123 529 1157
rect 559 1123 615 1157
rect 645 1123 701 1157
rect 731 1123 787 1157
rect 871 1123 927 1157
rect 957 1123 1013 1157
rect 1043 1123 1099 1157
rect 1129 1123 1185 1157
rect 1269 1123 1325 1157
rect 1355 1123 1411 1157
rect 1441 1123 1497 1157
rect 1527 1123 1583 1157
rect 1667 1123 1723 1157
rect 1753 1123 1809 1157
rect 1839 1123 1895 1157
rect 1925 1123 1981 1157
rect 2065 1123 2121 1157
rect 2151 1123 2207 1157
rect 2237 1123 2293 1157
rect 2323 1123 2379 1157
rect 2463 1123 2519 1157
rect 2549 1123 2605 1157
rect 2635 1123 2691 1157
rect 2721 1123 2777 1157
rect 2861 1123 2917 1157
rect 2947 1123 3003 1157
rect 3033 1123 3089 1157
rect 3119 1123 3175 1157
rect 3259 1123 3315 1157
rect 3345 1123 3401 1157
rect 3431 1123 3487 1157
rect 3517 1123 3573 1157
rect 3657 1123 3713 1157
rect 3743 1123 3799 1157
rect 3829 1123 3885 1157
rect 3915 1123 3971 1157
rect 4055 1123 4111 1157
rect 4141 1123 4197 1157
rect 4227 1123 4283 1157
rect 4313 1123 4369 1157
rect 4453 1123 4509 1157
rect 4539 1123 4595 1157
rect 4625 1123 4681 1157
rect 4711 1123 4767 1157
rect 4851 1123 4907 1157
rect 4937 1123 4993 1157
rect 5023 1123 5079 1157
rect 5109 1123 5165 1157
rect 5249 1123 5305 1157
rect 5335 1123 5391 1157
rect 5421 1123 5477 1157
rect 5507 1123 5563 1157
rect 5647 1123 5703 1157
rect 5733 1123 5789 1157
rect 5819 1123 5875 1157
rect 5905 1123 5961 1157
rect 6045 1123 6101 1157
rect 6131 1123 6187 1157
rect 6217 1123 6273 1157
rect 6303 1123 6359 1157
rect 6443 1123 6499 1157
rect 6529 1123 6585 1157
rect 6615 1123 6671 1157
rect 6701 1123 6757 1157
rect 6841 1123 6897 1157
rect 6927 1123 6983 1157
rect 7013 1123 7069 1157
rect 7099 1123 7155 1157
rect 7239 1123 7295 1157
rect 7325 1123 7381 1157
rect 7411 1123 7467 1157
rect 7497 1123 7553 1157
rect 7637 1123 7693 1157
rect 7723 1123 7779 1157
rect 7809 1123 7865 1157
rect 7895 1123 7951 1157
rect 8035 1123 8091 1157
rect 8121 1123 8177 1157
rect 8207 1123 8263 1157
rect 8293 1123 8349 1157
rect 8433 1123 8489 1157
rect 8519 1123 8575 1157
rect 8605 1123 8661 1157
rect 8691 1123 8747 1157
rect 8831 1123 8887 1157
rect 8917 1123 8973 1157
rect 9003 1123 9059 1157
rect 9089 1123 9145 1157
rect 9229 1123 9285 1157
rect 9315 1123 9371 1157
rect 9401 1123 9457 1157
rect 9487 1123 9543 1157
rect 9627 1123 9683 1157
rect 9713 1123 9769 1157
rect 9799 1123 9855 1157
rect 9885 1123 9941 1157
rect 86 1071 120 1123
rect 172 1071 206 1123
rect 258 1071 292 1123
rect 344 1071 378 1123
rect 484 1071 518 1123
rect 570 1071 604 1123
rect 656 1071 690 1123
rect 742 1071 776 1123
rect 882 1071 916 1123
rect 968 1071 1002 1123
rect 1054 1071 1088 1123
rect 1140 1071 1174 1123
rect 1280 1071 1314 1123
rect 1366 1071 1400 1123
rect 1452 1071 1486 1123
rect 1538 1071 1572 1123
rect 1678 1071 1712 1123
rect 1764 1071 1798 1123
rect 1850 1071 1884 1123
rect 1936 1071 1970 1123
rect 2076 1071 2110 1123
rect 2162 1071 2196 1123
rect 2248 1071 2282 1123
rect 2334 1071 2368 1123
rect 2474 1071 2508 1123
rect 2560 1071 2594 1123
rect 2646 1071 2680 1123
rect 2732 1071 2766 1123
rect 2872 1071 2906 1123
rect 2958 1071 2992 1123
rect 3044 1071 3078 1123
rect 3130 1071 3164 1123
rect 3270 1071 3304 1123
rect 3356 1071 3390 1123
rect 3442 1071 3476 1123
rect 3528 1071 3562 1123
rect 3668 1071 3702 1123
rect 3754 1071 3788 1123
rect 3840 1071 3874 1123
rect 3926 1071 3960 1123
rect 4066 1071 4100 1123
rect 4152 1071 4186 1123
rect 4238 1071 4272 1123
rect 4324 1071 4358 1123
rect 4464 1071 4498 1123
rect 4550 1071 4584 1123
rect 4636 1071 4670 1123
rect 4722 1071 4756 1123
rect 4862 1071 4896 1123
rect 4948 1071 4982 1123
rect 5034 1071 5068 1123
rect 5120 1071 5154 1123
rect 5260 1071 5294 1123
rect 5346 1071 5380 1123
rect 5432 1071 5466 1123
rect 5518 1071 5552 1123
rect 5658 1071 5692 1123
rect 5744 1071 5778 1123
rect 5830 1071 5864 1123
rect 5916 1071 5950 1123
rect 6056 1071 6090 1123
rect 6142 1071 6176 1123
rect 6228 1071 6262 1123
rect 6314 1071 6348 1123
rect 6454 1071 6488 1123
rect 6540 1071 6574 1123
rect 6626 1071 6660 1123
rect 6712 1071 6746 1123
rect 6852 1071 6886 1123
rect 6938 1071 6972 1123
rect 7024 1071 7058 1123
rect 7110 1071 7144 1123
rect 7250 1071 7284 1123
rect 7336 1071 7370 1123
rect 7422 1071 7456 1123
rect 7508 1071 7542 1123
rect 7648 1071 7682 1123
rect 7734 1071 7768 1123
rect 7820 1071 7854 1123
rect 7906 1071 7940 1123
rect 8046 1071 8080 1123
rect 8132 1071 8166 1123
rect 8218 1071 8252 1123
rect 8304 1071 8338 1123
rect 8444 1071 8478 1123
rect 8530 1071 8564 1123
rect 8616 1071 8650 1123
rect 8702 1071 8736 1123
rect 8842 1071 8876 1123
rect 8928 1071 8962 1123
rect 9014 1071 9048 1123
rect 9100 1071 9134 1123
rect 9240 1071 9274 1123
rect 9326 1071 9360 1123
rect 9412 1071 9446 1123
rect 9498 1071 9532 1123
rect 9638 1071 9672 1123
rect 9724 1071 9758 1123
rect 9810 1071 9844 1123
rect 9896 1071 9930 1123
rect 75 1037 131 1071
rect 161 1037 217 1071
rect 247 1037 303 1071
rect 333 1037 389 1071
rect 473 1037 529 1071
rect 559 1037 615 1071
rect 645 1037 701 1071
rect 731 1037 787 1071
rect 871 1037 927 1071
rect 957 1037 1013 1071
rect 1043 1037 1099 1071
rect 1129 1037 1185 1071
rect 1269 1037 1325 1071
rect 1355 1037 1411 1071
rect 1441 1037 1497 1071
rect 1527 1037 1583 1071
rect 1667 1037 1723 1071
rect 1753 1037 1809 1071
rect 1839 1037 1895 1071
rect 1925 1037 1981 1071
rect 2065 1037 2121 1071
rect 2151 1037 2207 1071
rect 2237 1037 2293 1071
rect 2323 1037 2379 1071
rect 2463 1037 2519 1071
rect 2549 1037 2605 1071
rect 2635 1037 2691 1071
rect 2721 1037 2777 1071
rect 2861 1037 2917 1071
rect 2947 1037 3003 1071
rect 3033 1037 3089 1071
rect 3119 1037 3175 1071
rect 3259 1037 3315 1071
rect 3345 1037 3401 1071
rect 3431 1037 3487 1071
rect 3517 1037 3573 1071
rect 3657 1037 3713 1071
rect 3743 1037 3799 1071
rect 3829 1037 3885 1071
rect 3915 1037 3971 1071
rect 4055 1037 4111 1071
rect 4141 1037 4197 1071
rect 4227 1037 4283 1071
rect 4313 1037 4369 1071
rect 4453 1037 4509 1071
rect 4539 1037 4595 1071
rect 4625 1037 4681 1071
rect 4711 1037 4767 1071
rect 4851 1037 4907 1071
rect 4937 1037 4993 1071
rect 5023 1037 5079 1071
rect 5109 1037 5165 1071
rect 5249 1037 5305 1071
rect 5335 1037 5391 1071
rect 5421 1037 5477 1071
rect 5507 1037 5563 1071
rect 5647 1037 5703 1071
rect 5733 1037 5789 1071
rect 5819 1037 5875 1071
rect 5905 1037 5961 1071
rect 6045 1037 6101 1071
rect 6131 1037 6187 1071
rect 6217 1037 6273 1071
rect 6303 1037 6359 1071
rect 6443 1037 6499 1071
rect 6529 1037 6585 1071
rect 6615 1037 6671 1071
rect 6701 1037 6757 1071
rect 6841 1037 6897 1071
rect 6927 1037 6983 1071
rect 7013 1037 7069 1071
rect 7099 1037 7155 1071
rect 7239 1037 7295 1071
rect 7325 1037 7381 1071
rect 7411 1037 7467 1071
rect 7497 1037 7553 1071
rect 7637 1037 7693 1071
rect 7723 1037 7779 1071
rect 7809 1037 7865 1071
rect 7895 1037 7951 1071
rect 8035 1037 8091 1071
rect 8121 1037 8177 1071
rect 8207 1037 8263 1071
rect 8293 1037 8349 1071
rect 8433 1037 8489 1071
rect 8519 1037 8575 1071
rect 8605 1037 8661 1071
rect 8691 1037 8747 1071
rect 8831 1037 8887 1071
rect 8917 1037 8973 1071
rect 9003 1037 9059 1071
rect 9089 1037 9145 1071
rect 9229 1037 9285 1071
rect 9315 1037 9371 1071
rect 9401 1037 9457 1071
rect 9487 1037 9543 1071
rect 9627 1037 9683 1071
rect 9713 1037 9769 1071
rect 9799 1037 9855 1071
rect 9885 1037 9941 1071
rect 86 985 120 1037
rect 172 985 206 1037
rect 258 985 292 1037
rect 344 985 378 1037
rect 484 985 518 1037
rect 570 985 604 1037
rect 656 985 690 1037
rect 742 985 776 1037
rect 882 985 916 1037
rect 968 985 1002 1037
rect 1054 985 1088 1037
rect 1140 985 1174 1037
rect 1280 985 1314 1037
rect 1366 985 1400 1037
rect 1452 985 1486 1037
rect 1538 985 1572 1037
rect 1678 985 1712 1037
rect 1764 985 1798 1037
rect 1850 985 1884 1037
rect 1936 985 1970 1037
rect 2076 985 2110 1037
rect 2162 985 2196 1037
rect 2248 985 2282 1037
rect 2334 985 2368 1037
rect 2474 985 2508 1037
rect 2560 985 2594 1037
rect 2646 985 2680 1037
rect 2732 985 2766 1037
rect 2872 985 2906 1037
rect 2958 985 2992 1037
rect 3044 985 3078 1037
rect 3130 985 3164 1037
rect 3270 985 3304 1037
rect 3356 985 3390 1037
rect 3442 985 3476 1037
rect 3528 985 3562 1037
rect 3668 985 3702 1037
rect 3754 985 3788 1037
rect 3840 985 3874 1037
rect 3926 985 3960 1037
rect 4066 985 4100 1037
rect 4152 985 4186 1037
rect 4238 985 4272 1037
rect 4324 985 4358 1037
rect 4464 985 4498 1037
rect 4550 985 4584 1037
rect 4636 985 4670 1037
rect 4722 985 4756 1037
rect 4862 985 4896 1037
rect 4948 985 4982 1037
rect 5034 985 5068 1037
rect 5120 985 5154 1037
rect 5260 985 5294 1037
rect 5346 985 5380 1037
rect 5432 985 5466 1037
rect 5518 985 5552 1037
rect 5658 985 5692 1037
rect 5744 985 5778 1037
rect 5830 985 5864 1037
rect 5916 985 5950 1037
rect 6056 985 6090 1037
rect 6142 985 6176 1037
rect 6228 985 6262 1037
rect 6314 985 6348 1037
rect 6454 985 6488 1037
rect 6540 985 6574 1037
rect 6626 985 6660 1037
rect 6712 985 6746 1037
rect 6852 985 6886 1037
rect 6938 985 6972 1037
rect 7024 985 7058 1037
rect 7110 985 7144 1037
rect 7250 985 7284 1037
rect 7336 985 7370 1037
rect 7422 985 7456 1037
rect 7508 985 7542 1037
rect 7648 985 7682 1037
rect 7734 985 7768 1037
rect 7820 985 7854 1037
rect 7906 985 7940 1037
rect 8046 985 8080 1037
rect 8132 985 8166 1037
rect 8218 985 8252 1037
rect 8304 985 8338 1037
rect 8444 985 8478 1037
rect 8530 985 8564 1037
rect 8616 985 8650 1037
rect 8702 985 8736 1037
rect 8842 985 8876 1037
rect 8928 985 8962 1037
rect 9014 985 9048 1037
rect 9100 985 9134 1037
rect 9240 985 9274 1037
rect 9326 985 9360 1037
rect 9412 985 9446 1037
rect 9498 985 9532 1037
rect 9638 985 9672 1037
rect 9724 985 9758 1037
rect 9810 985 9844 1037
rect 9896 985 9930 1037
rect 75 951 131 985
rect 161 951 217 985
rect 247 951 303 985
rect 333 951 389 985
rect 473 951 529 985
rect 559 951 615 985
rect 645 951 701 985
rect 731 951 787 985
rect 871 951 927 985
rect 957 951 1013 985
rect 1043 951 1099 985
rect 1129 951 1185 985
rect 1269 951 1325 985
rect 1355 951 1411 985
rect 1441 951 1497 985
rect 1527 951 1583 985
rect 1667 951 1723 985
rect 1753 951 1809 985
rect 1839 951 1895 985
rect 1925 951 1981 985
rect 2065 951 2121 985
rect 2151 951 2207 985
rect 2237 951 2293 985
rect 2323 951 2379 985
rect 2463 951 2519 985
rect 2549 951 2605 985
rect 2635 951 2691 985
rect 2721 951 2777 985
rect 2861 951 2917 985
rect 2947 951 3003 985
rect 3033 951 3089 985
rect 3119 951 3175 985
rect 3259 951 3315 985
rect 3345 951 3401 985
rect 3431 951 3487 985
rect 3517 951 3573 985
rect 3657 951 3713 985
rect 3743 951 3799 985
rect 3829 951 3885 985
rect 3915 951 3971 985
rect 4055 951 4111 985
rect 4141 951 4197 985
rect 4227 951 4283 985
rect 4313 951 4369 985
rect 4453 951 4509 985
rect 4539 951 4595 985
rect 4625 951 4681 985
rect 4711 951 4767 985
rect 4851 951 4907 985
rect 4937 951 4993 985
rect 5023 951 5079 985
rect 5109 951 5165 985
rect 5249 951 5305 985
rect 5335 951 5391 985
rect 5421 951 5477 985
rect 5507 951 5563 985
rect 5647 951 5703 985
rect 5733 951 5789 985
rect 5819 951 5875 985
rect 5905 951 5961 985
rect 6045 951 6101 985
rect 6131 951 6187 985
rect 6217 951 6273 985
rect 6303 951 6359 985
rect 6443 951 6499 985
rect 6529 951 6585 985
rect 6615 951 6671 985
rect 6701 951 6757 985
rect 6841 951 6897 985
rect 6927 951 6983 985
rect 7013 951 7069 985
rect 7099 951 7155 985
rect 7239 951 7295 985
rect 7325 951 7381 985
rect 7411 951 7467 985
rect 7497 951 7553 985
rect 7637 951 7693 985
rect 7723 951 7779 985
rect 7809 951 7865 985
rect 7895 951 7951 985
rect 8035 951 8091 985
rect 8121 951 8177 985
rect 8207 951 8263 985
rect 8293 951 8349 985
rect 8433 951 8489 985
rect 8519 951 8575 985
rect 8605 951 8661 985
rect 8691 951 8747 985
rect 8831 951 8887 985
rect 8917 951 8973 985
rect 9003 951 9059 985
rect 9089 951 9145 985
rect 9229 951 9285 985
rect 9315 951 9371 985
rect 9401 951 9457 985
rect 9487 951 9543 985
rect 9627 951 9683 985
rect 9713 951 9769 985
rect 9799 951 9855 985
rect 9885 951 9941 985
rect 86 898 120 951
rect 172 898 206 951
rect 258 898 292 951
rect 344 898 378 951
rect 484 898 518 951
rect 570 898 604 951
rect 656 898 690 951
rect 742 898 776 951
rect 882 898 916 951
rect 968 898 1002 951
rect 1054 898 1088 951
rect 1140 898 1174 951
rect 1280 898 1314 951
rect 1366 898 1400 951
rect 1452 898 1486 951
rect 1538 898 1572 951
rect 1678 898 1712 951
rect 1764 898 1798 951
rect 1850 898 1884 951
rect 1936 898 1970 951
rect 2076 898 2110 951
rect 2162 898 2196 951
rect 2248 898 2282 951
rect 2334 898 2368 951
rect 2474 898 2508 951
rect 2560 898 2594 951
rect 2646 898 2680 951
rect 2732 898 2766 951
rect 2872 898 2906 951
rect 2958 898 2992 951
rect 3044 898 3078 951
rect 3130 898 3164 951
rect 3270 898 3304 951
rect 3356 898 3390 951
rect 3442 898 3476 951
rect 3528 898 3562 951
rect 3668 898 3702 951
rect 3754 898 3788 951
rect 3840 898 3874 951
rect 3926 898 3960 951
rect 4066 898 4100 951
rect 4152 898 4186 951
rect 4238 898 4272 951
rect 4324 898 4358 951
rect 4464 898 4498 951
rect 4550 898 4584 951
rect 4636 898 4670 951
rect 4722 898 4756 951
rect 4862 898 4896 951
rect 4948 898 4982 951
rect 5034 898 5068 951
rect 5120 898 5154 951
rect 5260 898 5294 951
rect 5346 898 5380 951
rect 5432 898 5466 951
rect 5518 898 5552 951
rect 5658 898 5692 951
rect 5744 898 5778 951
rect 5830 898 5864 951
rect 5916 898 5950 951
rect 6056 898 6090 951
rect 6142 898 6176 951
rect 6228 898 6262 951
rect 6314 898 6348 951
rect 6454 898 6488 951
rect 6540 898 6574 951
rect 6626 898 6660 951
rect 6712 898 6746 951
rect 6852 898 6886 951
rect 6938 898 6972 951
rect 7024 898 7058 951
rect 7110 898 7144 951
rect 7250 898 7284 951
rect 7336 898 7370 951
rect 7422 898 7456 951
rect 7508 898 7542 951
rect 7648 898 7682 951
rect 7734 898 7768 951
rect 7820 898 7854 951
rect 7906 898 7940 951
rect 8046 898 8080 951
rect 8132 898 8166 951
rect 8218 898 8252 951
rect 8304 898 8338 951
rect 8444 898 8478 951
rect 8530 898 8564 951
rect 8616 898 8650 951
rect 8702 898 8736 951
rect 8842 898 8876 951
rect 8928 898 8962 951
rect 9014 898 9048 951
rect 9100 898 9134 951
rect 9240 898 9274 951
rect 9326 898 9360 951
rect 9412 898 9446 951
rect 9498 898 9532 951
rect 9638 898 9672 951
rect 9724 898 9758 951
rect 9810 898 9844 951
rect 9896 898 9930 951
rect 9980 898 10010 1302
rect 0 868 413 898
rect 443 868 1607 898
rect 1637 868 2403 898
rect 2433 868 3597 898
rect 3627 868 4393 898
rect 4423 868 5587 898
rect 5617 868 6383 898
rect 6413 868 7577 898
rect 7607 868 8373 898
rect 8403 868 9567 898
rect 9597 868 10010 898
rect 0 464 30 868
rect 86 809 120 868
rect 172 809 206 868
rect 258 809 292 868
rect 344 809 378 868
rect 484 809 518 868
rect 570 809 604 868
rect 656 809 690 868
rect 742 809 776 868
rect 882 809 916 868
rect 968 809 1002 868
rect 1054 809 1088 868
rect 1140 809 1174 868
rect 1280 809 1314 868
rect 1366 809 1400 868
rect 1452 809 1486 868
rect 1538 809 1572 868
rect 1678 809 1712 868
rect 1764 809 1798 868
rect 1850 809 1884 868
rect 1936 809 1970 868
rect 2076 809 2110 868
rect 2162 809 2196 868
rect 2248 809 2282 868
rect 2334 809 2368 868
rect 2474 809 2508 868
rect 2560 809 2594 868
rect 2646 809 2680 868
rect 2732 809 2766 868
rect 2872 809 2906 868
rect 2958 809 2992 868
rect 3044 809 3078 868
rect 3130 809 3164 868
rect 3270 809 3304 868
rect 3356 809 3390 868
rect 3442 809 3476 868
rect 3528 809 3562 868
rect 3668 809 3702 868
rect 3754 809 3788 868
rect 3840 809 3874 868
rect 3926 809 3960 868
rect 4066 809 4100 868
rect 4152 809 4186 868
rect 4238 809 4272 868
rect 4324 809 4358 868
rect 4464 809 4498 868
rect 4550 809 4584 868
rect 4636 809 4670 868
rect 4722 809 4756 868
rect 4862 809 4896 868
rect 4948 809 4982 868
rect 5034 809 5068 868
rect 5120 809 5154 868
rect 5260 809 5294 868
rect 5346 809 5380 868
rect 5432 809 5466 868
rect 5518 809 5552 868
rect 5658 809 5692 868
rect 5744 809 5778 868
rect 5830 809 5864 868
rect 5916 809 5950 868
rect 6056 809 6090 868
rect 6142 809 6176 868
rect 6228 809 6262 868
rect 6314 809 6348 868
rect 6454 809 6488 868
rect 6540 809 6574 868
rect 6626 809 6660 868
rect 6712 809 6746 868
rect 6852 809 6886 868
rect 6938 809 6972 868
rect 7024 809 7058 868
rect 7110 809 7144 868
rect 7250 809 7284 868
rect 7336 809 7370 868
rect 7422 809 7456 868
rect 7508 809 7542 868
rect 7648 809 7682 868
rect 7734 809 7768 868
rect 7820 809 7854 868
rect 7906 809 7940 868
rect 8046 809 8080 868
rect 8132 809 8166 868
rect 8218 809 8252 868
rect 8304 809 8338 868
rect 8444 809 8478 868
rect 8530 809 8564 868
rect 8616 809 8650 868
rect 8702 809 8736 868
rect 8842 809 8876 868
rect 8928 809 8962 868
rect 9014 809 9048 868
rect 9100 809 9134 868
rect 9240 809 9274 868
rect 9326 809 9360 868
rect 9412 809 9446 868
rect 9498 809 9532 868
rect 9638 809 9672 868
rect 9724 809 9758 868
rect 9810 809 9844 868
rect 9896 809 9930 868
rect 75 775 131 809
rect 161 775 217 809
rect 247 775 303 809
rect 333 775 389 809
rect 473 775 529 809
rect 559 775 615 809
rect 645 775 701 809
rect 731 775 787 809
rect 871 775 927 809
rect 957 775 1013 809
rect 1043 775 1099 809
rect 1129 775 1185 809
rect 1269 775 1325 809
rect 1355 775 1411 809
rect 1441 775 1497 809
rect 1527 775 1583 809
rect 1667 775 1723 809
rect 1753 775 1809 809
rect 1839 775 1895 809
rect 1925 775 1981 809
rect 2065 775 2121 809
rect 2151 775 2207 809
rect 2237 775 2293 809
rect 2323 775 2379 809
rect 2463 775 2519 809
rect 2549 775 2605 809
rect 2635 775 2691 809
rect 2721 775 2777 809
rect 2861 775 2917 809
rect 2947 775 3003 809
rect 3033 775 3089 809
rect 3119 775 3175 809
rect 3259 775 3315 809
rect 3345 775 3401 809
rect 3431 775 3487 809
rect 3517 775 3573 809
rect 3657 775 3713 809
rect 3743 775 3799 809
rect 3829 775 3885 809
rect 3915 775 3971 809
rect 4055 775 4111 809
rect 4141 775 4197 809
rect 4227 775 4283 809
rect 4313 775 4369 809
rect 4453 775 4509 809
rect 4539 775 4595 809
rect 4625 775 4681 809
rect 4711 775 4767 809
rect 4851 775 4907 809
rect 4937 775 4993 809
rect 5023 775 5079 809
rect 5109 775 5165 809
rect 5249 775 5305 809
rect 5335 775 5391 809
rect 5421 775 5477 809
rect 5507 775 5563 809
rect 5647 775 5703 809
rect 5733 775 5789 809
rect 5819 775 5875 809
rect 5905 775 5961 809
rect 6045 775 6101 809
rect 6131 775 6187 809
rect 6217 775 6273 809
rect 6303 775 6359 809
rect 6443 775 6499 809
rect 6529 775 6585 809
rect 6615 775 6671 809
rect 6701 775 6757 809
rect 6841 775 6897 809
rect 6927 775 6983 809
rect 7013 775 7069 809
rect 7099 775 7155 809
rect 7239 775 7295 809
rect 7325 775 7381 809
rect 7411 775 7467 809
rect 7497 775 7553 809
rect 7637 775 7693 809
rect 7723 775 7779 809
rect 7809 775 7865 809
rect 7895 775 7951 809
rect 8035 775 8091 809
rect 8121 775 8177 809
rect 8207 775 8263 809
rect 8293 775 8349 809
rect 8433 775 8489 809
rect 8519 775 8575 809
rect 8605 775 8661 809
rect 8691 775 8747 809
rect 8831 775 8887 809
rect 8917 775 8973 809
rect 9003 775 9059 809
rect 9089 775 9145 809
rect 9229 775 9285 809
rect 9315 775 9371 809
rect 9401 775 9457 809
rect 9487 775 9543 809
rect 9627 775 9683 809
rect 9713 775 9769 809
rect 9799 775 9855 809
rect 9885 775 9941 809
rect 86 723 120 775
rect 172 723 206 775
rect 258 723 292 775
rect 344 723 378 775
rect 484 723 518 775
rect 570 723 604 775
rect 656 723 690 775
rect 742 723 776 775
rect 882 723 916 775
rect 968 723 1002 775
rect 1054 723 1088 775
rect 1140 723 1174 775
rect 1280 723 1314 775
rect 1366 723 1400 775
rect 1452 723 1486 775
rect 1538 723 1572 775
rect 1678 723 1712 775
rect 1764 723 1798 775
rect 1850 723 1884 775
rect 1936 723 1970 775
rect 2076 723 2110 775
rect 2162 723 2196 775
rect 2248 723 2282 775
rect 2334 723 2368 775
rect 2474 723 2508 775
rect 2560 723 2594 775
rect 2646 723 2680 775
rect 2732 723 2766 775
rect 2872 723 2906 775
rect 2958 723 2992 775
rect 3044 723 3078 775
rect 3130 723 3164 775
rect 3270 723 3304 775
rect 3356 723 3390 775
rect 3442 723 3476 775
rect 3528 723 3562 775
rect 3668 723 3702 775
rect 3754 723 3788 775
rect 3840 723 3874 775
rect 3926 723 3960 775
rect 4066 723 4100 775
rect 4152 723 4186 775
rect 4238 723 4272 775
rect 4324 723 4358 775
rect 4464 723 4498 775
rect 4550 723 4584 775
rect 4636 723 4670 775
rect 4722 723 4756 775
rect 4862 723 4896 775
rect 4948 723 4982 775
rect 5034 723 5068 775
rect 5120 723 5154 775
rect 5260 723 5294 775
rect 5346 723 5380 775
rect 5432 723 5466 775
rect 5518 723 5552 775
rect 5658 723 5692 775
rect 5744 723 5778 775
rect 5830 723 5864 775
rect 5916 723 5950 775
rect 6056 723 6090 775
rect 6142 723 6176 775
rect 6228 723 6262 775
rect 6314 723 6348 775
rect 6454 723 6488 775
rect 6540 723 6574 775
rect 6626 723 6660 775
rect 6712 723 6746 775
rect 6852 723 6886 775
rect 6938 723 6972 775
rect 7024 723 7058 775
rect 7110 723 7144 775
rect 7250 723 7284 775
rect 7336 723 7370 775
rect 7422 723 7456 775
rect 7508 723 7542 775
rect 7648 723 7682 775
rect 7734 723 7768 775
rect 7820 723 7854 775
rect 7906 723 7940 775
rect 8046 723 8080 775
rect 8132 723 8166 775
rect 8218 723 8252 775
rect 8304 723 8338 775
rect 8444 723 8478 775
rect 8530 723 8564 775
rect 8616 723 8650 775
rect 8702 723 8736 775
rect 8842 723 8876 775
rect 8928 723 8962 775
rect 9014 723 9048 775
rect 9100 723 9134 775
rect 9240 723 9274 775
rect 9326 723 9360 775
rect 9412 723 9446 775
rect 9498 723 9532 775
rect 9638 723 9672 775
rect 9724 723 9758 775
rect 9810 723 9844 775
rect 9896 723 9930 775
rect 75 689 131 723
rect 161 689 217 723
rect 247 689 303 723
rect 333 689 389 723
rect 473 689 529 723
rect 559 689 615 723
rect 645 689 701 723
rect 731 689 787 723
rect 871 689 927 723
rect 957 689 1013 723
rect 1043 689 1099 723
rect 1129 689 1185 723
rect 1269 689 1325 723
rect 1355 689 1411 723
rect 1441 689 1497 723
rect 1527 689 1583 723
rect 1667 689 1723 723
rect 1753 689 1809 723
rect 1839 689 1895 723
rect 1925 689 1981 723
rect 2065 689 2121 723
rect 2151 689 2207 723
rect 2237 689 2293 723
rect 2323 689 2379 723
rect 2463 689 2519 723
rect 2549 689 2605 723
rect 2635 689 2691 723
rect 2721 689 2777 723
rect 2861 689 2917 723
rect 2947 689 3003 723
rect 3033 689 3089 723
rect 3119 689 3175 723
rect 3259 689 3315 723
rect 3345 689 3401 723
rect 3431 689 3487 723
rect 3517 689 3573 723
rect 3657 689 3713 723
rect 3743 689 3799 723
rect 3829 689 3885 723
rect 3915 689 3971 723
rect 4055 689 4111 723
rect 4141 689 4197 723
rect 4227 689 4283 723
rect 4313 689 4369 723
rect 4453 689 4509 723
rect 4539 689 4595 723
rect 4625 689 4681 723
rect 4711 689 4767 723
rect 4851 689 4907 723
rect 4937 689 4993 723
rect 5023 689 5079 723
rect 5109 689 5165 723
rect 5249 689 5305 723
rect 5335 689 5391 723
rect 5421 689 5477 723
rect 5507 689 5563 723
rect 5647 689 5703 723
rect 5733 689 5789 723
rect 5819 689 5875 723
rect 5905 689 5961 723
rect 6045 689 6101 723
rect 6131 689 6187 723
rect 6217 689 6273 723
rect 6303 689 6359 723
rect 6443 689 6499 723
rect 6529 689 6585 723
rect 6615 689 6671 723
rect 6701 689 6757 723
rect 6841 689 6897 723
rect 6927 689 6983 723
rect 7013 689 7069 723
rect 7099 689 7155 723
rect 7239 689 7295 723
rect 7325 689 7381 723
rect 7411 689 7467 723
rect 7497 689 7553 723
rect 7637 689 7693 723
rect 7723 689 7779 723
rect 7809 689 7865 723
rect 7895 689 7951 723
rect 8035 689 8091 723
rect 8121 689 8177 723
rect 8207 689 8263 723
rect 8293 689 8349 723
rect 8433 689 8489 723
rect 8519 689 8575 723
rect 8605 689 8661 723
rect 8691 689 8747 723
rect 8831 689 8887 723
rect 8917 689 8973 723
rect 9003 689 9059 723
rect 9089 689 9145 723
rect 9229 689 9285 723
rect 9315 689 9371 723
rect 9401 689 9457 723
rect 9487 689 9543 723
rect 9627 689 9683 723
rect 9713 689 9769 723
rect 9799 689 9855 723
rect 9885 689 9941 723
rect 86 637 120 689
rect 172 637 206 689
rect 258 637 292 689
rect 344 637 378 689
rect 484 637 518 689
rect 570 637 604 689
rect 656 637 690 689
rect 742 637 776 689
rect 882 637 916 689
rect 968 637 1002 689
rect 1054 637 1088 689
rect 1140 637 1174 689
rect 1280 637 1314 689
rect 1366 637 1400 689
rect 1452 637 1486 689
rect 1538 637 1572 689
rect 1678 637 1712 689
rect 1764 637 1798 689
rect 1850 637 1884 689
rect 1936 637 1970 689
rect 2076 637 2110 689
rect 2162 637 2196 689
rect 2248 637 2282 689
rect 2334 637 2368 689
rect 2474 637 2508 689
rect 2560 637 2594 689
rect 2646 637 2680 689
rect 2732 637 2766 689
rect 2872 637 2906 689
rect 2958 637 2992 689
rect 3044 637 3078 689
rect 3130 637 3164 689
rect 3270 637 3304 689
rect 3356 637 3390 689
rect 3442 637 3476 689
rect 3528 637 3562 689
rect 3668 637 3702 689
rect 3754 637 3788 689
rect 3840 637 3874 689
rect 3926 637 3960 689
rect 4066 637 4100 689
rect 4152 637 4186 689
rect 4238 637 4272 689
rect 4324 637 4358 689
rect 4464 637 4498 689
rect 4550 637 4584 689
rect 4636 637 4670 689
rect 4722 637 4756 689
rect 4862 637 4896 689
rect 4948 637 4982 689
rect 5034 637 5068 689
rect 5120 637 5154 689
rect 5260 637 5294 689
rect 5346 637 5380 689
rect 5432 637 5466 689
rect 5518 637 5552 689
rect 5658 637 5692 689
rect 5744 637 5778 689
rect 5830 637 5864 689
rect 5916 637 5950 689
rect 6056 637 6090 689
rect 6142 637 6176 689
rect 6228 637 6262 689
rect 6314 637 6348 689
rect 6454 637 6488 689
rect 6540 637 6574 689
rect 6626 637 6660 689
rect 6712 637 6746 689
rect 6852 637 6886 689
rect 6938 637 6972 689
rect 7024 637 7058 689
rect 7110 637 7144 689
rect 7250 637 7284 689
rect 7336 637 7370 689
rect 7422 637 7456 689
rect 7508 637 7542 689
rect 7648 637 7682 689
rect 7734 637 7768 689
rect 7820 637 7854 689
rect 7906 637 7940 689
rect 8046 637 8080 689
rect 8132 637 8166 689
rect 8218 637 8252 689
rect 8304 637 8338 689
rect 8444 637 8478 689
rect 8530 637 8564 689
rect 8616 637 8650 689
rect 8702 637 8736 689
rect 8842 637 8876 689
rect 8928 637 8962 689
rect 9014 637 9048 689
rect 9100 637 9134 689
rect 9240 637 9274 689
rect 9326 637 9360 689
rect 9412 637 9446 689
rect 9498 637 9532 689
rect 9638 637 9672 689
rect 9724 637 9758 689
rect 9810 637 9844 689
rect 9896 637 9930 689
rect 75 603 131 637
rect 161 603 217 637
rect 247 603 303 637
rect 333 603 389 637
rect 473 603 529 637
rect 559 603 615 637
rect 645 603 701 637
rect 731 603 787 637
rect 871 603 927 637
rect 957 603 1013 637
rect 1043 603 1099 637
rect 1129 603 1185 637
rect 1269 603 1325 637
rect 1355 603 1411 637
rect 1441 603 1497 637
rect 1527 603 1583 637
rect 1667 603 1723 637
rect 1753 603 1809 637
rect 1839 603 1895 637
rect 1925 603 1981 637
rect 2065 603 2121 637
rect 2151 603 2207 637
rect 2237 603 2293 637
rect 2323 603 2379 637
rect 2463 603 2519 637
rect 2549 603 2605 637
rect 2635 603 2691 637
rect 2721 603 2777 637
rect 2861 603 2917 637
rect 2947 603 3003 637
rect 3033 603 3089 637
rect 3119 603 3175 637
rect 3259 603 3315 637
rect 3345 603 3401 637
rect 3431 603 3487 637
rect 3517 603 3573 637
rect 3657 603 3713 637
rect 3743 603 3799 637
rect 3829 603 3885 637
rect 3915 603 3971 637
rect 4055 603 4111 637
rect 4141 603 4197 637
rect 4227 603 4283 637
rect 4313 603 4369 637
rect 4453 603 4509 637
rect 4539 603 4595 637
rect 4625 603 4681 637
rect 4711 603 4767 637
rect 4851 603 4907 637
rect 4937 603 4993 637
rect 5023 603 5079 637
rect 5109 603 5165 637
rect 5249 603 5305 637
rect 5335 603 5391 637
rect 5421 603 5477 637
rect 5507 603 5563 637
rect 5647 603 5703 637
rect 5733 603 5789 637
rect 5819 603 5875 637
rect 5905 603 5961 637
rect 6045 603 6101 637
rect 6131 603 6187 637
rect 6217 603 6273 637
rect 6303 603 6359 637
rect 6443 603 6499 637
rect 6529 603 6585 637
rect 6615 603 6671 637
rect 6701 603 6757 637
rect 6841 603 6897 637
rect 6927 603 6983 637
rect 7013 603 7069 637
rect 7099 603 7155 637
rect 7239 603 7295 637
rect 7325 603 7381 637
rect 7411 603 7467 637
rect 7497 603 7553 637
rect 7637 603 7693 637
rect 7723 603 7779 637
rect 7809 603 7865 637
rect 7895 603 7951 637
rect 8035 603 8091 637
rect 8121 603 8177 637
rect 8207 603 8263 637
rect 8293 603 8349 637
rect 8433 603 8489 637
rect 8519 603 8575 637
rect 8605 603 8661 637
rect 8691 603 8747 637
rect 8831 603 8887 637
rect 8917 603 8973 637
rect 9003 603 9059 637
rect 9089 603 9145 637
rect 9229 603 9285 637
rect 9315 603 9371 637
rect 9401 603 9457 637
rect 9487 603 9543 637
rect 9627 603 9683 637
rect 9713 603 9769 637
rect 9799 603 9855 637
rect 9885 603 9941 637
rect 86 551 120 603
rect 172 551 206 603
rect 258 551 292 603
rect 344 551 378 603
rect 484 551 518 603
rect 570 551 604 603
rect 656 551 690 603
rect 742 551 776 603
rect 882 551 916 603
rect 968 551 1002 603
rect 1054 551 1088 603
rect 1140 551 1174 603
rect 1280 551 1314 603
rect 1366 551 1400 603
rect 1452 551 1486 603
rect 1538 551 1572 603
rect 1678 551 1712 603
rect 1764 551 1798 603
rect 1850 551 1884 603
rect 1936 551 1970 603
rect 2076 551 2110 603
rect 2162 551 2196 603
rect 2248 551 2282 603
rect 2334 551 2368 603
rect 2474 551 2508 603
rect 2560 551 2594 603
rect 2646 551 2680 603
rect 2732 551 2766 603
rect 2872 551 2906 603
rect 2958 551 2992 603
rect 3044 551 3078 603
rect 3130 551 3164 603
rect 3270 551 3304 603
rect 3356 551 3390 603
rect 3442 551 3476 603
rect 3528 551 3562 603
rect 3668 551 3702 603
rect 3754 551 3788 603
rect 3840 551 3874 603
rect 3926 551 3960 603
rect 4066 551 4100 603
rect 4152 551 4186 603
rect 4238 551 4272 603
rect 4324 551 4358 603
rect 4464 551 4498 603
rect 4550 551 4584 603
rect 4636 551 4670 603
rect 4722 551 4756 603
rect 4862 551 4896 603
rect 4948 551 4982 603
rect 5034 551 5068 603
rect 5120 551 5154 603
rect 5260 551 5294 603
rect 5346 551 5380 603
rect 5432 551 5466 603
rect 5518 551 5552 603
rect 5658 551 5692 603
rect 5744 551 5778 603
rect 5830 551 5864 603
rect 5916 551 5950 603
rect 6056 551 6090 603
rect 6142 551 6176 603
rect 6228 551 6262 603
rect 6314 551 6348 603
rect 6454 551 6488 603
rect 6540 551 6574 603
rect 6626 551 6660 603
rect 6712 551 6746 603
rect 6852 551 6886 603
rect 6938 551 6972 603
rect 7024 551 7058 603
rect 7110 551 7144 603
rect 7250 551 7284 603
rect 7336 551 7370 603
rect 7422 551 7456 603
rect 7508 551 7542 603
rect 7648 551 7682 603
rect 7734 551 7768 603
rect 7820 551 7854 603
rect 7906 551 7940 603
rect 8046 551 8080 603
rect 8132 551 8166 603
rect 8218 551 8252 603
rect 8304 551 8338 603
rect 8444 551 8478 603
rect 8530 551 8564 603
rect 8616 551 8650 603
rect 8702 551 8736 603
rect 8842 551 8876 603
rect 8928 551 8962 603
rect 9014 551 9048 603
rect 9100 551 9134 603
rect 9240 551 9274 603
rect 9326 551 9360 603
rect 9412 551 9446 603
rect 9498 551 9532 603
rect 9638 551 9672 603
rect 9724 551 9758 603
rect 9810 551 9844 603
rect 9896 551 9930 603
rect 75 517 131 551
rect 161 517 217 551
rect 247 517 303 551
rect 333 517 389 551
rect 473 517 529 551
rect 559 517 615 551
rect 645 517 701 551
rect 731 517 787 551
rect 871 517 927 551
rect 957 517 1013 551
rect 1043 517 1099 551
rect 1129 517 1185 551
rect 1269 517 1325 551
rect 1355 517 1411 551
rect 1441 517 1497 551
rect 1527 517 1583 551
rect 1667 517 1723 551
rect 1753 517 1809 551
rect 1839 517 1895 551
rect 1925 517 1981 551
rect 2065 517 2121 551
rect 2151 517 2207 551
rect 2237 517 2293 551
rect 2323 517 2379 551
rect 2463 517 2519 551
rect 2549 517 2605 551
rect 2635 517 2691 551
rect 2721 517 2777 551
rect 2861 517 2917 551
rect 2947 517 3003 551
rect 3033 517 3089 551
rect 3119 517 3175 551
rect 3259 517 3315 551
rect 3345 517 3401 551
rect 3431 517 3487 551
rect 3517 517 3573 551
rect 3657 517 3713 551
rect 3743 517 3799 551
rect 3829 517 3885 551
rect 3915 517 3971 551
rect 4055 517 4111 551
rect 4141 517 4197 551
rect 4227 517 4283 551
rect 4313 517 4369 551
rect 4453 517 4509 551
rect 4539 517 4595 551
rect 4625 517 4681 551
rect 4711 517 4767 551
rect 4851 517 4907 551
rect 4937 517 4993 551
rect 5023 517 5079 551
rect 5109 517 5165 551
rect 5249 517 5305 551
rect 5335 517 5391 551
rect 5421 517 5477 551
rect 5507 517 5563 551
rect 5647 517 5703 551
rect 5733 517 5789 551
rect 5819 517 5875 551
rect 5905 517 5961 551
rect 6045 517 6101 551
rect 6131 517 6187 551
rect 6217 517 6273 551
rect 6303 517 6359 551
rect 6443 517 6499 551
rect 6529 517 6585 551
rect 6615 517 6671 551
rect 6701 517 6757 551
rect 6841 517 6897 551
rect 6927 517 6983 551
rect 7013 517 7069 551
rect 7099 517 7155 551
rect 7239 517 7295 551
rect 7325 517 7381 551
rect 7411 517 7467 551
rect 7497 517 7553 551
rect 7637 517 7693 551
rect 7723 517 7779 551
rect 7809 517 7865 551
rect 7895 517 7951 551
rect 8035 517 8091 551
rect 8121 517 8177 551
rect 8207 517 8263 551
rect 8293 517 8349 551
rect 8433 517 8489 551
rect 8519 517 8575 551
rect 8605 517 8661 551
rect 8691 517 8747 551
rect 8831 517 8887 551
rect 8917 517 8973 551
rect 9003 517 9059 551
rect 9089 517 9145 551
rect 9229 517 9285 551
rect 9315 517 9371 551
rect 9401 517 9457 551
rect 9487 517 9543 551
rect 9627 517 9683 551
rect 9713 517 9769 551
rect 9799 517 9855 551
rect 9885 517 9941 551
rect 86 464 120 517
rect 172 464 206 517
rect 258 464 292 517
rect 344 464 378 517
rect 484 464 518 517
rect 570 464 604 517
rect 656 464 690 517
rect 742 464 776 517
rect 882 464 916 517
rect 968 464 1002 517
rect 1054 464 1088 517
rect 1140 464 1174 517
rect 1280 464 1314 517
rect 1366 464 1400 517
rect 1452 464 1486 517
rect 1538 464 1572 517
rect 1678 464 1712 517
rect 1764 464 1798 517
rect 1850 464 1884 517
rect 1936 464 1970 517
rect 2076 464 2110 517
rect 2162 464 2196 517
rect 2248 464 2282 517
rect 2334 464 2368 517
rect 2474 464 2508 517
rect 2560 464 2594 517
rect 2646 464 2680 517
rect 2732 464 2766 517
rect 2872 464 2906 517
rect 2958 464 2992 517
rect 3044 464 3078 517
rect 3130 464 3164 517
rect 3270 464 3304 517
rect 3356 464 3390 517
rect 3442 464 3476 517
rect 3528 464 3562 517
rect 3668 464 3702 517
rect 3754 464 3788 517
rect 3840 464 3874 517
rect 3926 464 3960 517
rect 4066 464 4100 517
rect 4152 464 4186 517
rect 4238 464 4272 517
rect 4324 464 4358 517
rect 4464 464 4498 517
rect 4550 464 4584 517
rect 4636 464 4670 517
rect 4722 464 4756 517
rect 4862 464 4896 517
rect 4948 464 4982 517
rect 5034 464 5068 517
rect 5120 464 5154 517
rect 5260 464 5294 517
rect 5346 464 5380 517
rect 5432 464 5466 517
rect 5518 464 5552 517
rect 5658 464 5692 517
rect 5744 464 5778 517
rect 5830 464 5864 517
rect 5916 464 5950 517
rect 6056 464 6090 517
rect 6142 464 6176 517
rect 6228 464 6262 517
rect 6314 464 6348 517
rect 6454 464 6488 517
rect 6540 464 6574 517
rect 6626 464 6660 517
rect 6712 464 6746 517
rect 6852 464 6886 517
rect 6938 464 6972 517
rect 7024 464 7058 517
rect 7110 464 7144 517
rect 7250 464 7284 517
rect 7336 464 7370 517
rect 7422 464 7456 517
rect 7508 464 7542 517
rect 7648 464 7682 517
rect 7734 464 7768 517
rect 7820 464 7854 517
rect 7906 464 7940 517
rect 8046 464 8080 517
rect 8132 464 8166 517
rect 8218 464 8252 517
rect 8304 464 8338 517
rect 8444 464 8478 517
rect 8530 464 8564 517
rect 8616 464 8650 517
rect 8702 464 8736 517
rect 8842 464 8876 517
rect 8928 464 8962 517
rect 9014 464 9048 517
rect 9100 464 9134 517
rect 9240 464 9274 517
rect 9326 464 9360 517
rect 9412 464 9446 517
rect 9498 464 9532 517
rect 9638 464 9672 517
rect 9724 464 9758 517
rect 9810 464 9844 517
rect 9896 464 9930 517
rect 9980 464 10010 868
rect 0 434 413 464
rect 443 434 1607 464
rect 1637 434 2403 464
rect 2433 434 3597 464
rect 3627 434 4393 464
rect 4423 434 5587 464
rect 5617 434 6383 464
rect 6413 434 7577 464
rect 7607 434 8373 464
rect 8403 434 9567 464
rect 9597 434 10010 464
rect 0 30 30 434
rect 86 375 120 434
rect 172 375 206 434
rect 258 375 292 434
rect 344 375 378 434
rect 484 375 518 404
rect 570 375 604 404
rect 656 375 690 404
rect 742 375 776 404
rect 882 375 916 404
rect 968 375 1002 404
rect 1054 375 1088 404
rect 1140 375 1174 404
rect 1280 375 1314 404
rect 1366 375 1400 404
rect 1452 375 1486 404
rect 1538 375 1572 404
rect 1678 375 1712 434
rect 1764 375 1798 434
rect 1850 375 1884 434
rect 1936 375 1970 434
rect 2076 375 2110 434
rect 2162 375 2196 434
rect 2248 375 2282 434
rect 2334 375 2368 434
rect 2474 375 2508 404
rect 2560 375 2594 404
rect 2646 375 2680 404
rect 2732 375 2766 404
rect 2872 375 2906 434
rect 2958 375 2992 434
rect 3044 375 3078 434
rect 3130 375 3164 434
rect 3270 375 3304 404
rect 3356 375 3390 404
rect 3442 375 3476 404
rect 3528 375 3562 404
rect 3668 375 3702 434
rect 3754 375 3788 434
rect 3840 375 3874 434
rect 3926 375 3960 434
rect 4066 375 4100 434
rect 4152 375 4186 434
rect 4238 375 4272 434
rect 4324 375 4358 434
rect 4464 375 4498 404
rect 4550 375 4584 404
rect 4636 375 4670 404
rect 4722 375 4756 404
rect 4862 375 4896 434
rect 4948 375 4982 434
rect 5034 375 5068 434
rect 5120 375 5154 434
rect 5260 375 5294 404
rect 5346 375 5380 404
rect 5432 375 5466 404
rect 5518 375 5552 404
rect 5658 375 5692 434
rect 5744 375 5778 434
rect 5830 375 5864 434
rect 5916 375 5950 434
rect 6056 375 6090 434
rect 6142 375 6176 434
rect 6228 375 6262 434
rect 6314 375 6348 434
rect 6454 375 6488 404
rect 6540 375 6574 404
rect 6626 375 6660 404
rect 6712 375 6746 404
rect 6852 375 6886 434
rect 6938 375 6972 434
rect 7024 375 7058 404
rect 7110 375 7144 404
rect 7250 375 7284 404
rect 7336 375 7370 404
rect 7422 375 7456 404
rect 7508 375 7542 404
rect 7648 375 7682 434
rect 7734 375 7768 434
rect 7820 375 7854 434
rect 7906 375 7940 434
rect 8046 375 8080 434
rect 8132 375 8166 434
rect 8218 375 8252 434
rect 8304 375 8338 434
rect 8444 375 8478 404
rect 8530 375 8564 404
rect 8616 375 8650 404
rect 8702 375 8736 404
rect 8842 375 8876 404
rect 8928 375 8962 434
rect 9014 375 9048 404
rect 9100 375 9134 404
rect 9240 375 9274 404
rect 9326 375 9360 404
rect 9412 375 9446 404
rect 9498 375 9532 404
rect 9638 375 9672 434
rect 9724 375 9758 434
rect 9810 375 9844 434
rect 9896 375 9930 434
rect 75 341 131 375
rect 161 341 217 375
rect 247 341 303 375
rect 333 341 389 375
rect 473 341 529 375
rect 559 341 615 375
rect 645 341 701 375
rect 731 341 787 375
rect 871 341 927 375
rect 957 341 1013 375
rect 1043 341 1099 375
rect 1129 341 1185 375
rect 1269 341 1325 375
rect 1355 341 1411 375
rect 1441 341 1497 375
rect 1527 341 1583 375
rect 1667 341 1723 375
rect 1753 341 1809 375
rect 1839 341 1895 375
rect 1925 341 1981 375
rect 2065 341 2121 375
rect 2151 341 2207 375
rect 2237 341 2293 375
rect 2323 341 2379 375
rect 2463 341 2519 375
rect 2549 341 2605 375
rect 2635 341 2691 375
rect 2721 341 2777 375
rect 2861 341 2917 375
rect 2947 341 3003 375
rect 3033 341 3089 375
rect 3119 341 3175 375
rect 3259 341 3315 375
rect 3345 341 3401 375
rect 3431 341 3487 375
rect 3517 341 3573 375
rect 3657 341 3713 375
rect 3743 341 3799 375
rect 3829 341 3885 375
rect 3915 341 3971 375
rect 4055 341 4111 375
rect 4141 341 4197 375
rect 4227 341 4283 375
rect 4313 341 4369 375
rect 4453 341 4509 375
rect 4539 341 4595 375
rect 4625 341 4681 375
rect 4711 341 4767 375
rect 4851 341 4907 375
rect 4937 341 4993 375
rect 5023 341 5079 375
rect 5109 341 5165 375
rect 5249 341 5305 375
rect 5335 341 5391 375
rect 5421 341 5477 375
rect 5507 341 5563 375
rect 5647 341 5703 375
rect 5733 341 5789 375
rect 5819 341 5875 375
rect 5905 341 5961 375
rect 6045 341 6101 375
rect 6131 341 6187 375
rect 6217 341 6273 375
rect 6303 341 6359 375
rect 6443 341 6499 375
rect 6529 341 6585 375
rect 6615 341 6671 375
rect 6701 341 6757 375
rect 6841 341 6897 375
rect 6927 341 6983 375
rect 7013 341 7069 375
rect 7099 341 7155 375
rect 7239 341 7295 375
rect 7325 341 7381 375
rect 7411 341 7467 375
rect 7497 341 7553 375
rect 7637 341 7693 375
rect 7723 341 7779 375
rect 7809 341 7865 375
rect 7895 341 7951 375
rect 8035 341 8091 375
rect 8121 341 8177 375
rect 8207 341 8263 375
rect 8293 341 8349 375
rect 8433 341 8489 375
rect 8519 341 8575 375
rect 8605 341 8661 375
rect 8691 341 8747 375
rect 8831 341 8887 375
rect 8917 341 8973 375
rect 9003 341 9059 375
rect 9089 341 9145 375
rect 9229 341 9285 375
rect 9315 341 9371 375
rect 9401 341 9457 375
rect 9487 341 9543 375
rect 9627 341 9683 375
rect 9713 341 9769 375
rect 9799 341 9855 375
rect 9885 341 9941 375
rect 86 289 120 341
rect 172 289 206 341
rect 258 289 292 341
rect 344 289 378 341
rect 484 289 518 341
rect 570 289 604 341
rect 656 289 690 341
rect 742 289 776 341
rect 882 289 916 341
rect 968 289 1002 341
rect 1054 289 1088 341
rect 1140 289 1174 341
rect 1280 289 1314 341
rect 1366 289 1400 341
rect 1452 289 1486 341
rect 1538 289 1572 341
rect 1678 289 1712 341
rect 1764 289 1798 341
rect 1850 289 1884 341
rect 1936 289 1970 341
rect 2076 289 2110 341
rect 2162 289 2196 341
rect 2248 289 2282 341
rect 2334 289 2368 341
rect 2474 289 2508 341
rect 2560 289 2594 341
rect 2646 289 2680 341
rect 2732 289 2766 341
rect 2872 289 2906 341
rect 2958 289 2992 341
rect 3044 289 3078 341
rect 3130 289 3164 341
rect 3270 289 3304 341
rect 3356 289 3390 341
rect 3442 289 3476 341
rect 3528 289 3562 341
rect 3668 289 3702 341
rect 3754 289 3788 341
rect 3840 289 3874 341
rect 3926 289 3960 341
rect 4066 289 4100 341
rect 4152 289 4186 341
rect 4238 289 4272 341
rect 4324 289 4358 341
rect 4464 289 4498 341
rect 4550 289 4584 341
rect 4636 289 4670 341
rect 4722 289 4756 341
rect 4862 325 4896 341
rect 4948 325 4982 341
rect 5034 325 5068 341
rect 5120 325 5154 341
rect 5260 289 5294 341
rect 5346 289 5380 341
rect 5432 289 5466 341
rect 5518 289 5552 341
rect 5658 289 5692 341
rect 5744 289 5778 341
rect 5830 289 5864 341
rect 5916 289 5950 341
rect 6056 289 6090 341
rect 6142 289 6176 341
rect 6228 289 6262 341
rect 6314 289 6348 341
rect 6454 289 6488 341
rect 6540 289 6574 341
rect 6626 289 6660 341
rect 6712 289 6746 341
rect 6852 325 6886 341
rect 6938 325 6972 341
rect 7024 289 7058 341
rect 7110 289 7144 341
rect 7250 289 7284 341
rect 7336 289 7370 341
rect 7422 289 7456 341
rect 7508 289 7542 341
rect 7648 289 7682 341
rect 7734 289 7768 341
rect 7820 289 7854 341
rect 7906 289 7940 341
rect 8046 289 8080 341
rect 8132 289 8166 341
rect 8218 289 8252 341
rect 8304 289 8338 341
rect 8444 289 8478 341
rect 8530 289 8564 341
rect 8616 289 8650 341
rect 8702 289 8736 341
rect 8842 289 8876 341
rect 8928 325 8962 341
rect 9014 289 9048 341
rect 9100 289 9134 341
rect 9240 289 9274 341
rect 9326 289 9360 341
rect 9412 289 9446 341
rect 9498 289 9532 341
rect 9638 289 9672 341
rect 9724 289 9758 341
rect 9810 289 9844 341
rect 9896 289 9930 341
rect 75 255 131 289
rect 161 255 217 289
rect 247 255 303 289
rect 333 255 389 289
rect 473 255 529 289
rect 559 255 615 289
rect 645 255 701 289
rect 731 255 787 289
rect 871 255 927 289
rect 957 255 1013 289
rect 1043 255 1099 289
rect 1129 255 1185 289
rect 1269 255 1325 289
rect 1355 255 1411 289
rect 1441 255 1497 289
rect 1527 255 1583 289
rect 1667 255 1723 289
rect 1753 255 1809 289
rect 1839 255 1895 289
rect 1925 255 1981 289
rect 2065 255 2121 289
rect 2151 255 2207 289
rect 2237 255 2293 289
rect 2323 255 2379 289
rect 2463 255 2519 289
rect 2549 255 2605 289
rect 2635 255 2691 289
rect 2721 255 2777 289
rect 2861 255 2917 289
rect 2947 255 3003 289
rect 3033 255 3089 289
rect 3119 255 3175 289
rect 3259 255 3315 289
rect 3345 255 3401 289
rect 3431 255 3487 289
rect 3517 255 3573 289
rect 3657 255 3713 289
rect 3743 255 3799 289
rect 3829 255 3885 289
rect 3915 255 3971 289
rect 4055 255 4111 289
rect 4141 255 4197 289
rect 4227 255 4283 289
rect 4313 255 4369 289
rect 4453 255 4509 289
rect 4539 255 4595 289
rect 4625 255 4681 289
rect 4711 255 4767 289
rect 4851 255 4907 289
rect 4937 255 4993 289
rect 5023 255 5079 289
rect 5109 255 5165 289
rect 5249 255 5305 289
rect 5335 255 5391 289
rect 5421 255 5477 289
rect 5507 255 5563 289
rect 5647 255 5703 289
rect 5733 255 5789 289
rect 5819 255 5875 289
rect 5905 255 5961 289
rect 6045 255 6101 289
rect 6131 255 6187 289
rect 6217 255 6273 289
rect 6303 255 6359 289
rect 6443 255 6499 289
rect 6529 255 6585 289
rect 6615 255 6671 289
rect 6701 255 6757 289
rect 6841 255 6897 289
rect 6927 255 6983 289
rect 7013 255 7069 289
rect 7099 255 7155 289
rect 7239 255 7295 289
rect 7325 255 7381 289
rect 7411 255 7467 289
rect 7497 255 7553 289
rect 7637 255 7693 289
rect 7723 255 7779 289
rect 7809 255 7865 289
rect 7895 255 7951 289
rect 8035 255 8091 289
rect 8121 255 8177 289
rect 8207 255 8263 289
rect 8293 255 8349 289
rect 8433 255 8489 289
rect 8519 255 8575 289
rect 8605 255 8661 289
rect 8691 255 8747 289
rect 8831 255 8887 289
rect 8917 255 8973 289
rect 9003 255 9059 289
rect 9089 255 9145 289
rect 9229 255 9285 289
rect 9315 255 9371 289
rect 9401 255 9457 289
rect 9487 255 9543 289
rect 9627 255 9683 289
rect 9713 255 9769 289
rect 9799 255 9855 289
rect 9885 255 9941 289
rect 86 203 120 255
rect 172 203 206 255
rect 258 203 292 255
rect 344 203 378 255
rect 484 203 518 255
rect 570 203 604 255
rect 656 203 690 255
rect 742 203 776 255
rect 882 203 916 255
rect 968 203 1002 255
rect 1054 203 1088 255
rect 1140 203 1174 255
rect 1280 203 1314 255
rect 1366 203 1400 255
rect 1452 203 1486 255
rect 1538 203 1572 255
rect 1678 203 1712 255
rect 1764 203 1798 255
rect 1850 203 1884 255
rect 1936 203 1970 255
rect 2076 203 2110 255
rect 2162 203 2196 255
rect 2248 203 2282 255
rect 2334 203 2368 255
rect 2474 203 2508 255
rect 2560 203 2594 255
rect 2646 203 2680 255
rect 2732 203 2766 255
rect 2872 239 2906 255
rect 2958 239 2992 255
rect 3044 239 3078 255
rect 3130 239 3164 255
rect 3270 203 3304 255
rect 3356 203 3390 255
rect 3442 203 3476 255
rect 3528 203 3562 255
rect 3668 203 3702 255
rect 3754 203 3788 255
rect 3840 203 3874 255
rect 3926 203 3960 255
rect 4066 203 4100 255
rect 4152 203 4186 255
rect 4238 203 4272 255
rect 4324 203 4358 255
rect 4464 203 4498 255
rect 4550 203 4584 255
rect 4636 203 4670 255
rect 4722 203 4756 255
rect 4862 203 4896 255
rect 4948 203 4982 255
rect 5034 203 5068 255
rect 5120 203 5154 255
rect 5260 203 5294 255
rect 5346 203 5380 255
rect 5432 203 5466 255
rect 5518 203 5552 255
rect 5658 203 5692 255
rect 5744 203 5778 255
rect 5830 203 5864 255
rect 5916 203 5950 255
rect 6056 203 6090 255
rect 6142 203 6176 255
rect 6228 203 6262 255
rect 6314 203 6348 255
rect 6454 203 6488 255
rect 6540 203 6574 255
rect 6626 203 6660 255
rect 6712 203 6746 255
rect 6852 203 6886 255
rect 6938 203 6972 255
rect 7024 203 7058 255
rect 7110 203 7144 255
rect 7250 203 7284 255
rect 7336 203 7370 255
rect 7422 203 7456 255
rect 7508 203 7542 255
rect 7648 203 7682 255
rect 7734 203 7768 255
rect 7820 203 7854 255
rect 7906 203 7940 255
rect 8046 203 8080 255
rect 8132 203 8166 255
rect 8218 203 8252 255
rect 8304 203 8338 255
rect 8444 203 8478 255
rect 8530 203 8564 255
rect 8616 203 8650 255
rect 8702 203 8736 255
rect 8842 203 8876 255
rect 8928 203 8962 255
rect 9014 203 9048 255
rect 9100 203 9134 255
rect 9240 203 9274 255
rect 9326 203 9360 255
rect 9412 203 9446 255
rect 9498 203 9532 255
rect 9638 203 9672 255
rect 9724 203 9758 255
rect 9810 203 9844 255
rect 9896 203 9930 255
rect 75 169 131 203
rect 161 169 217 203
rect 247 169 303 203
rect 333 169 389 203
rect 473 169 529 203
rect 559 169 615 203
rect 645 169 701 203
rect 731 169 787 203
rect 871 169 927 203
rect 957 169 1013 203
rect 1043 169 1099 203
rect 1129 169 1185 203
rect 1269 169 1325 203
rect 1355 169 1411 203
rect 1441 169 1497 203
rect 1527 169 1583 203
rect 1667 169 1723 203
rect 1753 169 1809 203
rect 1839 169 1895 203
rect 1925 169 1981 203
rect 2065 169 2121 203
rect 2151 169 2207 203
rect 2237 169 2293 203
rect 2323 169 2379 203
rect 2463 169 2519 203
rect 2549 169 2605 203
rect 2635 169 2691 203
rect 2721 169 2777 203
rect 2861 169 2917 203
rect 2947 169 3003 203
rect 3033 169 3089 203
rect 3119 169 3175 203
rect 3259 169 3315 203
rect 3345 169 3401 203
rect 3431 169 3487 203
rect 3517 169 3573 203
rect 3657 169 3713 203
rect 3743 169 3799 203
rect 3829 169 3885 203
rect 3915 169 3971 203
rect 4055 169 4111 203
rect 4141 169 4197 203
rect 4227 169 4283 203
rect 4313 169 4369 203
rect 4453 169 4509 203
rect 4539 169 4595 203
rect 4625 169 4681 203
rect 4711 169 4767 203
rect 4851 169 4907 203
rect 4937 169 4993 203
rect 5023 169 5079 203
rect 5109 169 5165 203
rect 5249 169 5305 203
rect 5335 169 5391 203
rect 5421 169 5477 203
rect 5507 169 5563 203
rect 5647 169 5703 203
rect 5733 169 5789 203
rect 5819 169 5875 203
rect 5905 169 5961 203
rect 6045 169 6101 203
rect 6131 169 6187 203
rect 6217 169 6273 203
rect 6303 169 6359 203
rect 6443 169 6499 203
rect 6529 169 6585 203
rect 6615 169 6671 203
rect 6701 169 6757 203
rect 6841 169 6897 203
rect 6927 169 6983 203
rect 7013 169 7069 203
rect 7099 169 7155 203
rect 7239 169 7295 203
rect 7325 169 7381 203
rect 7411 169 7467 203
rect 7497 169 7553 203
rect 7637 169 7693 203
rect 7723 169 7779 203
rect 7809 169 7865 203
rect 7895 169 7951 203
rect 8035 169 8091 203
rect 8121 169 8177 203
rect 8207 169 8263 203
rect 8293 169 8349 203
rect 8433 169 8489 203
rect 8519 169 8575 203
rect 8605 169 8661 203
rect 8691 169 8747 203
rect 8831 169 8887 203
rect 8917 169 8973 203
rect 9003 169 9059 203
rect 9089 169 9145 203
rect 9229 169 9285 203
rect 9315 169 9371 203
rect 9401 169 9457 203
rect 9487 169 9543 203
rect 9627 169 9683 203
rect 9713 169 9769 203
rect 9799 169 9855 203
rect 9885 169 9941 203
rect 86 117 120 169
rect 172 117 206 169
rect 258 117 292 169
rect 344 117 378 169
rect 484 117 518 169
rect 570 117 604 169
rect 656 117 690 169
rect 742 117 776 169
rect 882 117 916 169
rect 968 117 1002 169
rect 1054 117 1088 169
rect 1140 117 1174 169
rect 1280 117 1314 169
rect 1366 117 1400 169
rect 1452 117 1486 169
rect 1538 117 1572 169
rect 1678 117 1712 169
rect 1764 117 1798 169
rect 1850 117 1884 169
rect 1936 117 1970 169
rect 2076 117 2110 169
rect 2162 117 2196 169
rect 2248 117 2282 169
rect 2334 117 2368 169
rect 2474 117 2508 169
rect 2560 117 2594 169
rect 2646 117 2680 169
rect 2732 117 2766 169
rect 2872 117 2906 169
rect 2958 117 2992 169
rect 3044 117 3078 169
rect 3130 117 3164 169
rect 3270 117 3304 169
rect 3356 117 3390 169
rect 3442 117 3476 169
rect 3528 117 3562 169
rect 3668 117 3702 169
rect 3754 117 3788 169
rect 3840 117 3874 169
rect 3926 117 3960 169
rect 4066 117 4100 169
rect 4152 117 4186 169
rect 4238 117 4272 169
rect 4324 117 4358 169
rect 4464 117 4498 169
rect 4550 117 4584 169
rect 4636 117 4670 169
rect 4722 117 4756 169
rect 4862 117 4896 169
rect 4948 117 4982 169
rect 5034 117 5068 169
rect 5120 117 5154 169
rect 5260 117 5294 169
rect 5346 117 5380 169
rect 5432 117 5466 169
rect 5518 117 5552 169
rect 5658 117 5692 169
rect 5744 117 5778 169
rect 5830 117 5864 169
rect 5916 117 5950 169
rect 6056 117 6090 169
rect 6142 117 6176 169
rect 6228 117 6262 169
rect 6314 117 6348 169
rect 6454 117 6488 169
rect 6540 117 6574 169
rect 6626 117 6660 169
rect 6712 117 6746 169
rect 6852 117 6886 169
rect 6938 117 6972 169
rect 7024 117 7058 169
rect 7110 117 7144 169
rect 7250 117 7284 169
rect 7336 117 7370 169
rect 7422 117 7456 169
rect 7508 117 7542 169
rect 7648 117 7682 169
rect 7734 117 7768 169
rect 7820 117 7854 169
rect 7906 117 7940 169
rect 8046 117 8080 169
rect 8132 117 8166 169
rect 8218 117 8252 169
rect 8304 117 8338 169
rect 8444 117 8478 169
rect 8530 117 8564 169
rect 8616 117 8650 169
rect 8702 117 8736 169
rect 8842 117 8876 169
rect 8928 117 8962 169
rect 9014 117 9048 169
rect 9100 117 9134 169
rect 9240 117 9274 169
rect 9326 117 9360 169
rect 9412 117 9446 169
rect 9498 117 9532 169
rect 9638 117 9672 169
rect 9724 117 9758 169
rect 9810 117 9844 169
rect 9896 117 9930 169
rect 75 83 131 117
rect 161 83 217 117
rect 247 83 303 117
rect 333 83 389 117
rect 473 83 529 117
rect 559 83 615 117
rect 645 83 701 117
rect 731 83 787 117
rect 871 83 927 117
rect 957 83 1013 117
rect 1043 83 1099 117
rect 1129 83 1185 117
rect 1269 83 1325 117
rect 1355 83 1411 117
rect 1441 83 1497 117
rect 1527 83 1583 117
rect 1667 83 1723 117
rect 1753 83 1809 117
rect 1839 83 1895 117
rect 1925 83 1981 117
rect 2065 83 2121 117
rect 2151 83 2207 117
rect 2237 83 2293 117
rect 2323 83 2379 117
rect 2463 83 2519 117
rect 2549 83 2605 117
rect 2635 83 2691 117
rect 2721 83 2777 117
rect 2861 83 2917 117
rect 2947 83 3003 117
rect 3033 83 3089 117
rect 3119 83 3175 117
rect 3259 83 3315 117
rect 3345 83 3401 117
rect 3431 83 3487 117
rect 3517 83 3573 117
rect 3657 83 3713 117
rect 3743 83 3799 117
rect 3829 83 3885 117
rect 3915 83 3971 117
rect 4055 83 4111 117
rect 4141 83 4197 117
rect 4227 83 4283 117
rect 4313 83 4369 117
rect 4453 83 4509 117
rect 4539 83 4595 117
rect 4625 83 4681 117
rect 4711 83 4767 117
rect 4851 83 4907 117
rect 4937 83 4993 117
rect 5023 83 5079 117
rect 5109 83 5165 117
rect 5249 83 5305 117
rect 5335 83 5391 117
rect 5421 83 5477 117
rect 5507 83 5563 117
rect 5647 83 5703 117
rect 5733 83 5789 117
rect 5819 83 5875 117
rect 5905 83 5961 117
rect 6045 83 6101 117
rect 6131 83 6187 117
rect 6217 83 6273 117
rect 6303 83 6359 117
rect 6443 83 6499 117
rect 6529 83 6585 117
rect 6615 83 6671 117
rect 6701 83 6757 117
rect 6841 83 6897 117
rect 6927 83 6983 117
rect 7013 83 7069 117
rect 7099 83 7155 117
rect 7239 83 7295 117
rect 7325 83 7381 117
rect 7411 83 7467 117
rect 7497 83 7553 117
rect 7637 83 7693 117
rect 7723 83 7779 117
rect 7809 83 7865 117
rect 7895 83 7951 117
rect 8035 83 8091 117
rect 8121 83 8177 117
rect 8207 83 8263 117
rect 8293 83 8349 117
rect 8433 83 8489 117
rect 8519 83 8575 117
rect 8605 83 8661 117
rect 8691 83 8747 117
rect 8831 83 8887 117
rect 8917 83 8973 117
rect 9003 83 9059 117
rect 9089 83 9145 117
rect 9229 83 9285 117
rect 9315 83 9371 117
rect 9401 83 9457 117
rect 9487 83 9543 117
rect 9627 83 9683 117
rect 9713 83 9769 117
rect 9799 83 9855 117
rect 9885 83 9941 117
rect 86 30 120 83
rect 172 30 206 83
rect 258 30 292 83
rect 344 30 378 83
rect 484 30 518 83
rect 570 30 604 83
rect 656 30 690 83
rect 742 30 776 83
rect 882 30 916 83
rect 968 30 1002 83
rect 1054 30 1088 83
rect 1140 30 1174 83
rect 1280 30 1314 83
rect 1366 30 1400 83
rect 1452 30 1486 83
rect 1538 30 1572 83
rect 1678 30 1712 83
rect 1764 30 1798 83
rect 1850 30 1884 83
rect 1936 30 1970 83
rect 2076 30 2110 83
rect 2162 30 2196 83
rect 2248 30 2282 83
rect 2334 30 2368 83
rect 2474 30 2508 83
rect 2560 30 2594 83
rect 2646 30 2680 83
rect 2732 30 2766 83
rect 2872 66 2906 83
rect 2958 66 2992 83
rect 3044 66 3078 83
rect 3130 66 3164 83
rect 3270 30 3304 83
rect 3356 30 3390 83
rect 3442 30 3476 83
rect 3528 30 3562 83
rect 3668 30 3702 83
rect 3754 30 3788 83
rect 3840 30 3874 83
rect 3926 30 3960 83
rect 4066 30 4100 83
rect 4152 30 4186 83
rect 4238 30 4272 83
rect 4324 30 4358 83
rect 4464 30 4498 83
rect 4550 30 4584 83
rect 4636 30 4670 83
rect 4722 30 4756 83
rect 4862 66 4896 83
rect 4948 66 4982 83
rect 5034 66 5068 83
rect 5120 66 5154 83
rect 5260 30 5294 83
rect 5346 30 5380 83
rect 5432 30 5466 83
rect 5518 30 5552 83
rect 5658 30 5692 83
rect 5744 30 5778 83
rect 5830 30 5864 83
rect 5916 30 5950 83
rect 6056 30 6090 83
rect 6142 30 6176 83
rect 6228 30 6262 83
rect 6314 30 6348 83
rect 6454 30 6488 83
rect 6540 30 6574 83
rect 6626 30 6660 83
rect 6712 30 6746 83
rect 6852 66 6886 83
rect 6938 66 6972 83
rect 7024 66 7058 83
rect 7110 66 7144 83
rect 7250 30 7284 83
rect 7336 30 7370 83
rect 7422 30 7456 83
rect 7508 30 7542 83
rect 7648 30 7682 83
rect 7734 30 7768 83
rect 7820 30 7854 83
rect 7906 30 7940 83
rect 8046 30 8080 83
rect 8132 30 8166 83
rect 8218 30 8252 83
rect 8304 30 8338 83
rect 8444 30 8478 83
rect 8530 30 8564 83
rect 8616 30 8650 83
rect 8702 30 8736 83
rect 8842 66 8876 83
rect 8928 66 8962 83
rect 9014 66 9048 83
rect 9100 66 9134 83
rect 9240 30 9274 83
rect 9326 30 9360 83
rect 9412 30 9446 83
rect 9498 30 9532 83
rect 9638 30 9672 83
rect 9724 30 9758 83
rect 9810 30 9844 83
rect 9896 30 9930 83
rect 9980 30 10010 434
rect 0 0 10010 30
<< comment >>
rect 413 1736 428 1751
rect 811 1736 826 1751
rect 1209 1736 1224 1751
rect 1607 1736 1622 1751
rect 2005 1736 2020 1751
rect 2403 1736 2418 1751
rect 2801 1736 2816 1751
rect 3199 1736 3214 1751
rect 3597 1736 3612 1751
rect 3995 1736 4010 1751
rect 4393 1736 4408 1751
rect 4791 1736 4806 1751
rect 5189 1736 5204 1751
rect 5587 1736 5602 1751
rect 5985 1736 6000 1751
rect 6383 1736 6398 1751
rect 6781 1736 6796 1751
rect 7179 1736 7194 1751
rect 7577 1736 7592 1751
rect 7975 1736 7990 1751
rect 8373 1736 8388 1751
rect 8771 1736 8786 1751
rect 9169 1736 9184 1751
rect 9567 1736 9582 1751
rect 9965 1736 9980 1751
rect 30 1719 44 1726
rect 414 1719 442 1726
rect 812 1719 840 1726
rect 1210 1719 1238 1726
rect 1608 1719 1636 1726
rect 2006 1719 2034 1726
rect 2404 1719 2432 1726
rect 2802 1719 2830 1726
rect 3200 1719 3228 1726
rect 3598 1719 3626 1726
rect 3996 1719 4024 1726
rect 4394 1719 4422 1726
rect 4792 1719 4820 1726
rect 5190 1719 5218 1726
rect 5588 1719 5616 1726
rect 5986 1719 6014 1726
rect 6384 1719 6412 1726
rect 6782 1719 6810 1726
rect 7180 1719 7208 1726
rect 7578 1719 7606 1726
rect 7976 1719 8004 1726
rect 8374 1719 8402 1726
rect 8772 1719 8800 1726
rect 9170 1719 9198 1726
rect 9568 1719 9596 1726
rect 9966 1719 9980 1726
rect 30 1342 44 1349
rect 414 1342 442 1349
rect 812 1342 840 1349
rect 1210 1342 1238 1349
rect 1608 1342 1636 1349
rect 2006 1342 2034 1349
rect 2404 1342 2432 1349
rect 2802 1342 2830 1349
rect 3200 1342 3228 1349
rect 3598 1342 3626 1349
rect 3996 1342 4024 1349
rect 4394 1342 4422 1349
rect 4792 1342 4820 1349
rect 5190 1342 5218 1349
rect 5588 1342 5616 1349
rect 5986 1342 6014 1349
rect 6384 1342 6412 1349
rect 6782 1342 6810 1349
rect 7180 1342 7208 1349
rect 7578 1342 7606 1349
rect 7976 1342 8004 1349
rect 8374 1342 8402 1349
rect 8772 1342 8800 1349
rect 9170 1342 9198 1349
rect 9568 1342 9596 1349
rect 9966 1342 9980 1349
rect 413 1302 428 1317
rect 811 1302 826 1317
rect 1209 1302 1224 1317
rect 1607 1302 1622 1317
rect 2005 1302 2020 1317
rect 2403 1302 2418 1317
rect 2801 1302 2816 1317
rect 3199 1302 3214 1317
rect 3597 1302 3612 1317
rect 3995 1302 4010 1317
rect 4393 1302 4408 1317
rect 4791 1302 4806 1317
rect 5189 1302 5204 1317
rect 5587 1302 5602 1317
rect 5985 1302 6000 1317
rect 6383 1302 6398 1317
rect 6781 1302 6796 1317
rect 7179 1302 7194 1317
rect 7577 1302 7592 1317
rect 7975 1302 7990 1317
rect 8373 1302 8388 1317
rect 8771 1302 8786 1317
rect 9169 1302 9184 1317
rect 9567 1302 9582 1317
rect 9965 1302 9980 1317
rect 30 1285 44 1292
rect 414 1285 442 1292
rect 812 1285 840 1292
rect 1210 1285 1238 1292
rect 1608 1285 1636 1292
rect 2006 1285 2034 1292
rect 2404 1285 2432 1292
rect 2802 1285 2830 1292
rect 3200 1285 3228 1292
rect 3598 1285 3626 1292
rect 3996 1285 4024 1292
rect 4394 1285 4422 1292
rect 4792 1285 4820 1292
rect 5190 1285 5218 1292
rect 5588 1285 5616 1292
rect 5986 1285 6014 1292
rect 6384 1285 6412 1292
rect 6782 1285 6810 1292
rect 7180 1285 7208 1292
rect 7578 1285 7606 1292
rect 7976 1285 8004 1292
rect 8374 1285 8402 1292
rect 8772 1285 8800 1292
rect 9170 1285 9198 1292
rect 9568 1285 9596 1292
rect 9966 1285 9980 1292
rect 30 908 44 915
rect 414 908 442 915
rect 812 908 840 915
rect 1210 908 1238 915
rect 1608 908 1636 915
rect 2006 908 2034 915
rect 2404 908 2432 915
rect 2802 908 2830 915
rect 3200 908 3228 915
rect 3598 908 3626 915
rect 3996 908 4024 915
rect 4394 908 4422 915
rect 4792 908 4820 915
rect 5190 908 5218 915
rect 5588 908 5616 915
rect 5986 908 6014 915
rect 6384 908 6412 915
rect 6782 908 6810 915
rect 7180 908 7208 915
rect 7578 908 7606 915
rect 7976 908 8004 915
rect 8374 908 8402 915
rect 8772 908 8800 915
rect 9170 908 9198 915
rect 9568 908 9596 915
rect 9966 908 9980 915
rect 413 868 428 883
rect 811 868 826 883
rect 1209 868 1224 883
rect 1607 868 1622 883
rect 2005 868 2020 883
rect 2403 868 2418 883
rect 2801 868 2816 883
rect 3199 868 3214 883
rect 3597 868 3612 883
rect 3995 868 4010 883
rect 4393 868 4408 883
rect 4791 868 4806 883
rect 5189 868 5204 883
rect 5587 868 5602 883
rect 5985 868 6000 883
rect 6383 868 6398 883
rect 6781 868 6796 883
rect 7179 868 7194 883
rect 7577 868 7592 883
rect 7975 868 7990 883
rect 8373 868 8388 883
rect 8771 868 8786 883
rect 9169 868 9184 883
rect 9567 868 9582 883
rect 9965 868 9980 883
rect 30 851 44 858
rect 414 851 442 858
rect 812 851 840 858
rect 1210 851 1238 858
rect 1608 851 1636 858
rect 2006 851 2034 858
rect 2404 851 2432 858
rect 2802 851 2830 858
rect 3200 851 3228 858
rect 3598 851 3626 858
rect 3996 851 4024 858
rect 4394 851 4422 858
rect 4792 851 4820 858
rect 5190 851 5218 858
rect 5588 851 5616 858
rect 5986 851 6014 858
rect 6384 851 6412 858
rect 6782 851 6810 858
rect 7180 851 7208 858
rect 7578 851 7606 858
rect 7976 851 8004 858
rect 8374 851 8402 858
rect 8772 851 8800 858
rect 9170 851 9198 858
rect 9568 851 9596 858
rect 9966 851 9980 858
rect 30 474 44 481
rect 414 474 442 481
rect 812 474 840 481
rect 1210 474 1238 481
rect 1608 474 1636 481
rect 2006 474 2034 481
rect 2404 474 2432 481
rect 2802 474 2830 481
rect 3200 474 3228 481
rect 3598 474 3626 481
rect 3996 474 4024 481
rect 4394 474 4422 481
rect 4792 474 4820 481
rect 5190 474 5218 481
rect 5588 474 5616 481
rect 5986 474 6014 481
rect 6384 474 6412 481
rect 6782 474 6810 481
rect 7180 474 7208 481
rect 7578 474 7606 481
rect 7976 474 8004 481
rect 8374 474 8402 481
rect 8772 474 8800 481
rect 9170 474 9198 481
rect 9568 474 9596 481
rect 9966 474 9980 481
rect 428 449 443 464
rect 413 434 428 449
rect 811 434 826 449
rect 1209 434 1224 449
rect 1607 434 1622 449
rect 2005 434 2020 449
rect 2403 434 2418 449
rect 2801 434 2816 449
rect 3199 434 3214 449
rect 3597 434 3612 449
rect 3995 434 4010 449
rect 4393 434 4408 449
rect 4791 434 4806 449
rect 5189 434 5204 449
rect 5587 434 5602 449
rect 5985 434 6000 449
rect 6383 434 6398 449
rect 6781 434 6796 449
rect 7179 434 7194 449
rect 7577 434 7592 449
rect 7975 434 7990 449
rect 8373 434 8388 449
rect 8771 434 8786 449
rect 9169 434 9184 449
rect 9567 434 9582 449
rect 9965 434 9980 449
rect 30 417 44 424
rect 414 417 442 424
rect 812 417 840 424
rect 1210 417 1238 424
rect 1608 417 1636 424
rect 2006 417 2034 424
rect 2404 417 2432 424
rect 2802 417 2830 424
rect 3200 417 3228 424
rect 3598 417 3626 424
rect 3996 417 4024 424
rect 4394 417 4422 424
rect 4792 417 4820 424
rect 5190 417 5218 424
rect 5588 417 5616 424
rect 5986 417 6014 424
rect 6384 417 6412 424
rect 6782 417 6810 424
rect 7180 417 7208 424
rect 7578 417 7606 424
rect 7976 417 8004 424
rect 8374 417 8402 424
rect 8772 417 8800 424
rect 9170 417 9198 424
rect 9568 417 9596 424
rect 9966 417 9980 424
rect 30 40 44 47
rect 414 40 442 47
rect 812 40 840 47
rect 1210 40 1238 47
rect 1608 40 1636 47
rect 2006 40 2034 47
rect 2404 40 2432 47
rect 2802 40 2830 47
rect 3200 40 3228 47
rect 3598 40 3626 47
rect 3996 40 4024 47
rect 4394 40 4422 47
rect 4792 40 4820 47
rect 5190 40 5218 47
rect 5588 40 5616 47
rect 5986 40 6014 47
rect 6384 40 6412 47
rect 6782 40 6810 47
rect 7180 40 7208 47
rect 7578 40 7606 47
rect 7976 40 8004 47
rect 8374 40 8402 47
rect 8772 40 8800 47
rect 9170 40 9198 47
rect 9568 40 9596 47
rect 9966 40 9980 47
rect 15 15 30 30
rect 0 0 15 15
<< labels >>
rlabel metal4 0 63 0 86 7 extract_0/dummy_top
rlabel metal2 44 57 44 80 7 extract_0/dummy_bot
rlabel metal4 443 434 443 464 7 extract_0/top_16
rlabel metal2 442 481 442 511 7 extract_0/bot_16
rlabel metal4 2433 434 2433 464 7 extract_0/top_8
rlabel metal2 2432 481 2432 511 7 extract_0/bot_8
rlabel metal4 4423 434 4423 464 7 extract_0/top_4
rlabel metal2 4422 481 4422 511 7 extract_0/bot_4
rlabel metal4 6413 434 6413 464 7 extract_0/top_2
rlabel metal2 6412 481 6412 511 7 extract_0/bot_2
rlabel metal4 8403 434 8403 464 7 extract_0/top_1
rlabel metal2 8402 481 8402 511 7 extract_0/bot_1
<< end >>
