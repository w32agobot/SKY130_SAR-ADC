magic
tech sky130A
timestamp 1661167023
<< metal2 >>
rect 16 2431 432 2449
rect 16 2400 201 2431
rect 247 2400 432 2431
rect 16 2306 432 2400
rect 16 2275 201 2306
rect 247 2275 432 2306
rect 16 2182 432 2275
rect 16 2151 201 2182
rect 247 2176 432 2182
rect 464 2431 880 2449
rect 464 2400 649 2431
rect 695 2400 880 2431
rect 464 2306 880 2400
rect 464 2275 649 2306
rect 695 2275 880 2306
rect 464 2182 880 2275
rect 464 2176 649 2182
rect 247 2153 649 2176
rect 247 2151 432 2153
rect 16 2058 432 2151
rect 16 2027 201 2058
rect 247 2027 432 2058
rect 16 1934 432 2027
rect 16 1903 201 1934
rect 247 1903 432 1934
rect 16 1884 432 1903
rect 464 2151 649 2153
rect 695 2175 880 2182
rect 912 2431 1328 2449
rect 912 2400 1097 2431
rect 1143 2400 1328 2431
rect 912 2306 1328 2400
rect 912 2275 1097 2306
rect 1143 2275 1328 2306
rect 912 2182 1328 2275
rect 912 2175 1097 2182
rect 695 2152 1097 2175
rect 695 2151 880 2152
rect 464 2058 880 2151
rect 464 2027 649 2058
rect 695 2027 880 2058
rect 464 1934 880 2027
rect 464 1903 649 1934
rect 695 1903 880 1934
rect 464 1884 880 1903
rect 912 2151 1097 2152
rect 1143 2180 1328 2182
rect 1360 2431 1776 2449
rect 1360 2400 1545 2431
rect 1591 2400 1776 2431
rect 1360 2306 1776 2400
rect 1360 2275 1545 2306
rect 1591 2275 1776 2306
rect 1360 2182 1776 2275
rect 1360 2180 1545 2182
rect 1143 2157 1545 2180
rect 1143 2151 1328 2157
rect 912 2058 1328 2151
rect 912 2027 1097 2058
rect 1143 2027 1328 2058
rect 912 1934 1328 2027
rect 912 1903 1097 1934
rect 1143 1903 1328 1934
rect 912 1884 1328 1903
rect 1360 2151 1545 2157
rect 1591 2179 1776 2182
rect 1808 2431 2224 2449
rect 1808 2400 1993 2431
rect 2039 2400 2224 2431
rect 1808 2306 2224 2400
rect 1808 2275 1993 2306
rect 2039 2275 2224 2306
rect 1808 2182 2224 2275
rect 1808 2179 1993 2182
rect 1591 2156 1993 2179
rect 1591 2151 1776 2156
rect 1360 2058 1776 2151
rect 1360 2027 1545 2058
rect 1591 2027 1776 2058
rect 1360 1934 1776 2027
rect 1360 1903 1545 1934
rect 1591 1903 1776 1934
rect 1360 1884 1776 1903
rect 1808 2151 1993 2156
rect 2039 2177 2224 2182
rect 2256 2431 2672 2449
rect 2256 2400 2441 2431
rect 2487 2400 2672 2431
rect 2256 2306 2672 2400
rect 2256 2275 2441 2306
rect 2487 2275 2672 2306
rect 2256 2182 2672 2275
rect 2256 2177 2441 2182
rect 2039 2154 2441 2177
rect 2039 2151 2224 2154
rect 1808 2058 2224 2151
rect 1808 2027 1993 2058
rect 2039 2027 2224 2058
rect 1808 1934 2224 2027
rect 1808 1903 1993 1934
rect 2039 1903 2224 1934
rect 1808 1884 2224 1903
rect 2256 2151 2441 2154
rect 2487 2176 2672 2182
rect 2704 2431 3120 2449
rect 2704 2400 2889 2431
rect 2935 2400 3120 2431
rect 2704 2306 3120 2400
rect 2704 2275 2889 2306
rect 2935 2275 3120 2306
rect 2704 2182 3120 2275
rect 2704 2176 2889 2182
rect 2487 2153 2889 2176
rect 2487 2151 2672 2153
rect 2256 2058 2672 2151
rect 2256 2027 2441 2058
rect 2487 2027 2672 2058
rect 2256 1934 2672 2027
rect 2256 1903 2441 1934
rect 2487 1903 2672 1934
rect 2256 1884 2672 1903
rect 2704 2151 2889 2153
rect 2935 2175 3120 2182
rect 3152 2431 3568 2449
rect 3152 2400 3337 2431
rect 3383 2400 3568 2431
rect 3152 2306 3568 2400
rect 3152 2275 3337 2306
rect 3383 2275 3568 2306
rect 3152 2182 3568 2275
rect 3152 2175 3337 2182
rect 2935 2152 3337 2175
rect 2935 2151 3120 2152
rect 2704 2058 3120 2151
rect 2704 2027 2889 2058
rect 2935 2027 3120 2058
rect 2704 1934 3120 2027
rect 2704 1903 2889 1934
rect 2935 1903 3120 1934
rect 2704 1884 3120 1903
rect 3152 2151 3337 2152
rect 3383 2180 3568 2182
rect 3600 2431 4016 2449
rect 3600 2400 3785 2431
rect 3831 2400 4016 2431
rect 3600 2306 4016 2400
rect 3600 2275 3785 2306
rect 3831 2275 4016 2306
rect 3600 2182 4016 2275
rect 3600 2180 3785 2182
rect 3383 2157 3785 2180
rect 3383 2151 3568 2157
rect 3152 2058 3568 2151
rect 3152 2027 3337 2058
rect 3383 2027 3568 2058
rect 3152 1934 3568 2027
rect 3152 1903 3337 1934
rect 3383 1903 3568 1934
rect 3152 1884 3568 1903
rect 3600 2151 3785 2157
rect 3831 2179 4016 2182
rect 4048 2431 4464 2449
rect 4048 2400 4233 2431
rect 4279 2400 4464 2431
rect 4048 2306 4464 2400
rect 4048 2275 4233 2306
rect 4279 2275 4464 2306
rect 4048 2182 4464 2275
rect 4048 2179 4233 2182
rect 3831 2156 4233 2179
rect 3831 2151 4016 2156
rect 3600 2058 4016 2151
rect 3600 2027 3785 2058
rect 3831 2027 4016 2058
rect 3600 1934 4016 2027
rect 3600 1903 3785 1934
rect 3831 1903 4016 1934
rect 3600 1884 4016 1903
rect 4048 2151 4233 2156
rect 4279 2178 4464 2182
rect 4496 2431 4912 2449
rect 4496 2400 4681 2431
rect 4727 2400 4912 2431
rect 4496 2306 4912 2400
rect 4496 2275 4681 2306
rect 4727 2275 4912 2306
rect 4496 2182 4912 2275
rect 4496 2178 4681 2182
rect 4279 2154 4681 2178
rect 4279 2151 4464 2154
rect 4048 2058 4464 2151
rect 4048 2027 4233 2058
rect 4279 2027 4464 2058
rect 4048 1934 4464 2027
rect 4048 1903 4233 1934
rect 4279 1903 4464 1934
rect 4048 1884 4464 1903
rect 4496 2151 4681 2154
rect 4727 2176 4912 2182
rect 4944 2431 5360 2449
rect 4944 2400 5129 2431
rect 5175 2400 5360 2431
rect 4944 2306 5360 2400
rect 4944 2275 5129 2306
rect 5175 2275 5360 2306
rect 4944 2182 5360 2275
rect 4944 2176 5129 2182
rect 4727 2153 5129 2176
rect 4727 2151 4912 2153
rect 4496 2058 4912 2151
rect 4496 2027 4681 2058
rect 4727 2027 4912 2058
rect 4496 1934 4912 2027
rect 4496 1903 4681 1934
rect 4727 1903 4912 1934
rect 4496 1884 4912 1903
rect 4944 2151 5129 2153
rect 5175 2175 5360 2182
rect 5392 2431 5808 2449
rect 5392 2400 5577 2431
rect 5623 2400 5808 2431
rect 5392 2306 5808 2400
rect 5392 2275 5577 2306
rect 5623 2275 5808 2306
rect 5392 2182 5808 2275
rect 5392 2175 5577 2182
rect 5175 2152 5577 2175
rect 5175 2151 5360 2152
rect 4944 2058 5360 2151
rect 4944 2027 5129 2058
rect 5175 2027 5360 2058
rect 4944 1934 5360 2027
rect 4944 1903 5129 1934
rect 5175 1903 5360 1934
rect 4944 1884 5360 1903
rect 5392 2151 5577 2152
rect 5623 2180 5808 2182
rect 5840 2431 6256 2449
rect 5840 2400 6025 2431
rect 6071 2400 6256 2431
rect 5840 2306 6256 2400
rect 5840 2275 6025 2306
rect 6071 2275 6256 2306
rect 5840 2182 6256 2275
rect 5840 2180 6025 2182
rect 5623 2157 6025 2180
rect 5623 2151 5808 2157
rect 5392 2058 5808 2151
rect 5392 2027 5577 2058
rect 5623 2027 5808 2058
rect 5392 1934 5808 2027
rect 5392 1903 5577 1934
rect 5623 1903 5808 1934
rect 5392 1884 5808 1903
rect 5840 2151 6025 2157
rect 6071 2179 6256 2182
rect 6288 2431 6704 2449
rect 6288 2400 6473 2431
rect 6519 2400 6704 2431
rect 6288 2306 6704 2400
rect 6288 2275 6473 2306
rect 6519 2275 6704 2306
rect 6288 2182 6704 2275
rect 6288 2179 6473 2182
rect 6071 2156 6473 2179
rect 6071 2151 6256 2156
rect 5840 2058 6256 2151
rect 5840 2027 6025 2058
rect 6071 2027 6256 2058
rect 5840 1934 6256 2027
rect 5840 1903 6025 1934
rect 6071 1903 6256 1934
rect 5840 1884 6256 1903
rect 6288 2151 6473 2156
rect 6519 2177 6704 2182
rect 6736 2431 7152 2449
rect 6736 2400 6921 2431
rect 6967 2400 7152 2431
rect 6736 2306 7152 2400
rect 6736 2275 6921 2306
rect 6967 2275 7152 2306
rect 6736 2182 7152 2275
rect 6736 2177 6921 2182
rect 6519 2154 6921 2177
rect 6519 2151 6704 2154
rect 6288 2058 6704 2151
rect 6288 2027 6473 2058
rect 6519 2027 6704 2058
rect 6288 1934 6704 2027
rect 6288 1903 6473 1934
rect 6519 1903 6704 1934
rect 6288 1884 6704 1903
rect 6736 2151 6921 2154
rect 6967 2176 7152 2182
rect 7184 2431 7600 2449
rect 7184 2400 7369 2431
rect 7415 2400 7600 2431
rect 7184 2306 7600 2400
rect 7184 2275 7369 2306
rect 7415 2275 7600 2306
rect 7184 2182 7600 2275
rect 7184 2176 7369 2182
rect 6967 2153 7369 2176
rect 6967 2151 7152 2153
rect 6736 2058 7152 2151
rect 6736 2027 6921 2058
rect 6967 2027 7152 2058
rect 6736 1934 7152 2027
rect 6736 1903 6921 1934
rect 6967 1903 7152 1934
rect 6736 1884 7152 1903
rect 7184 2151 7369 2153
rect 7415 2175 7600 2182
rect 7632 2431 8048 2449
rect 7632 2400 7817 2431
rect 7863 2400 8048 2431
rect 7632 2306 8048 2400
rect 7632 2275 7817 2306
rect 7863 2275 8048 2306
rect 7632 2182 8048 2275
rect 7632 2175 7817 2182
rect 7415 2152 7817 2175
rect 7415 2151 7600 2152
rect 7184 2058 7600 2151
rect 7184 2027 7369 2058
rect 7415 2027 7600 2058
rect 7184 1934 7600 2027
rect 7184 1903 7369 1934
rect 7415 1903 7600 1934
rect 7184 1884 7600 1903
rect 7632 2151 7817 2152
rect 7863 2180 8048 2182
rect 8080 2431 8496 2449
rect 8080 2400 8265 2431
rect 8311 2400 8496 2431
rect 8080 2306 8496 2400
rect 8080 2275 8265 2306
rect 8311 2275 8496 2306
rect 8080 2182 8496 2275
rect 8080 2180 8265 2182
rect 7863 2157 8265 2180
rect 7863 2151 8048 2157
rect 7632 2058 8048 2151
rect 7632 2027 7817 2058
rect 7863 2027 8048 2058
rect 7632 1934 8048 2027
rect 7632 1903 7817 1934
rect 7863 1903 8048 1934
rect 7632 1884 8048 1903
rect 8080 2151 8265 2157
rect 8311 2179 8496 2182
rect 8528 2431 8944 2449
rect 8528 2400 8713 2431
rect 8759 2400 8944 2431
rect 8528 2306 8944 2400
rect 8528 2275 8713 2306
rect 8759 2275 8944 2306
rect 8528 2182 8944 2275
rect 8528 2179 8713 2182
rect 8311 2156 8713 2179
rect 8311 2151 8496 2156
rect 8080 2058 8496 2151
rect 8080 2027 8265 2058
rect 8311 2027 8496 2058
rect 8080 1934 8496 2027
rect 8080 1903 8265 1934
rect 8311 1903 8496 1934
rect 8080 1884 8496 1903
rect 8528 2151 8713 2156
rect 8759 2177 8944 2182
rect 8759 2154 8960 2177
rect 8759 2151 8944 2154
rect 8528 2058 8944 2151
rect 8528 2027 8713 2058
rect 8759 2027 8944 2058
rect 8528 1934 8944 2027
rect 8528 1903 8713 1934
rect 8759 1903 8944 1934
rect 8528 1884 8944 1903
rect 216 1830 237 1884
rect 2005 1830 2028 1884
rect 2456 1830 2477 1884
rect 4245 1830 4268 1884
rect 4696 1830 4717 1884
rect 6485 1830 6508 1884
rect 6936 1830 6957 1884
rect 8725 1830 8748 1884
rect 16 1812 432 1830
rect 16 1781 201 1812
rect 247 1781 432 1812
rect 16 1687 432 1781
rect 16 1656 201 1687
rect 247 1656 432 1687
rect 16 1563 432 1656
rect 16 1532 201 1563
rect 247 1532 432 1563
rect 16 1439 432 1532
rect 16 1408 201 1439
rect 247 1408 432 1439
rect 16 1315 432 1408
rect 16 1284 201 1315
rect 247 1284 432 1315
rect 16 1265 432 1284
rect 464 1812 880 1830
rect 464 1781 649 1812
rect 695 1781 880 1812
rect 464 1687 880 1781
rect 464 1656 649 1687
rect 695 1656 880 1687
rect 464 1563 880 1656
rect 464 1532 649 1563
rect 695 1551 880 1563
rect 912 1812 1328 1830
rect 912 1781 1097 1812
rect 1143 1781 1328 1812
rect 912 1687 1328 1781
rect 912 1656 1097 1687
rect 1143 1656 1328 1687
rect 912 1563 1328 1656
rect 912 1551 1097 1563
rect 695 1532 1097 1551
rect 1143 1556 1328 1563
rect 1360 1812 1776 1830
rect 1360 1781 1545 1812
rect 1591 1781 1776 1812
rect 1360 1687 1776 1781
rect 1360 1656 1545 1687
rect 1591 1656 1776 1687
rect 1360 1563 1776 1656
rect 1360 1556 1545 1563
rect 1143 1537 1545 1556
rect 1143 1532 1328 1537
rect 464 1439 880 1532
rect 464 1408 649 1439
rect 695 1408 880 1439
rect 464 1315 880 1408
rect 464 1284 649 1315
rect 695 1284 880 1315
rect 464 1265 880 1284
rect 912 1439 1328 1532
rect 912 1408 1097 1439
rect 1143 1408 1328 1439
rect 912 1315 1328 1408
rect 912 1284 1097 1315
rect 1143 1284 1328 1315
rect 912 1265 1328 1284
rect 1360 1532 1545 1537
rect 1591 1532 1776 1563
rect 1360 1439 1776 1532
rect 1360 1408 1545 1439
rect 1591 1408 1776 1439
rect 1360 1315 1776 1408
rect 1360 1284 1545 1315
rect 1591 1284 1776 1315
rect 1360 1265 1776 1284
rect 1808 1812 2224 1830
rect 1808 1781 1993 1812
rect 2039 1781 2224 1812
rect 1808 1687 2224 1781
rect 1808 1656 1993 1687
rect 2039 1656 2224 1687
rect 1808 1563 2224 1656
rect 1808 1532 1993 1563
rect 2039 1532 2224 1563
rect 1808 1439 2224 1532
rect 1808 1408 1993 1439
rect 2039 1408 2224 1439
rect 1808 1315 2224 1408
rect 1808 1284 1993 1315
rect 2039 1284 2224 1315
rect 1808 1265 2224 1284
rect 2256 1812 2672 1830
rect 2256 1781 2441 1812
rect 2487 1781 2672 1812
rect 2256 1687 2672 1781
rect 2256 1656 2441 1687
rect 2487 1656 2672 1687
rect 2256 1563 2672 1656
rect 2256 1532 2441 1563
rect 2487 1532 2672 1563
rect 2256 1439 2672 1532
rect 2256 1408 2441 1439
rect 2487 1408 2672 1439
rect 2256 1315 2672 1408
rect 2256 1284 2441 1315
rect 2487 1284 2672 1315
rect 2256 1265 2672 1284
rect 2704 1812 3120 1830
rect 2704 1781 2889 1812
rect 2935 1781 3120 1812
rect 2704 1687 3120 1781
rect 2704 1656 2889 1687
rect 2935 1656 3120 1687
rect 2704 1563 3120 1656
rect 2704 1532 2889 1563
rect 2935 1551 3120 1563
rect 3152 1812 3568 1830
rect 3152 1781 3337 1812
rect 3383 1781 3568 1812
rect 3152 1687 3568 1781
rect 3152 1656 3337 1687
rect 3383 1656 3568 1687
rect 3152 1563 3568 1656
rect 3152 1551 3337 1563
rect 2935 1532 3337 1551
rect 3383 1556 3568 1563
rect 3600 1812 4016 1830
rect 3600 1781 3785 1812
rect 3831 1781 4016 1812
rect 3600 1687 4016 1781
rect 3600 1656 3785 1687
rect 3831 1656 4016 1687
rect 3600 1563 4016 1656
rect 3600 1556 3785 1563
rect 3383 1537 3785 1556
rect 3383 1532 3568 1537
rect 2704 1439 3120 1532
rect 2704 1408 2889 1439
rect 2935 1408 3120 1439
rect 2704 1315 3120 1408
rect 2704 1284 2889 1315
rect 2935 1284 3120 1315
rect 2704 1265 3120 1284
rect 3152 1439 3568 1532
rect 3152 1408 3337 1439
rect 3383 1408 3568 1439
rect 3152 1315 3568 1408
rect 3152 1284 3337 1315
rect 3383 1284 3568 1315
rect 3152 1265 3568 1284
rect 3600 1532 3785 1537
rect 3831 1532 4016 1563
rect 3600 1439 4016 1532
rect 3600 1408 3785 1439
rect 3831 1408 4016 1439
rect 3600 1315 4016 1408
rect 3600 1284 3785 1315
rect 3831 1284 4016 1315
rect 3600 1265 4016 1284
rect 4048 1812 4464 1830
rect 4048 1781 4233 1812
rect 4279 1781 4464 1812
rect 4048 1687 4464 1781
rect 4048 1656 4233 1687
rect 4279 1656 4464 1687
rect 4048 1563 4464 1656
rect 4048 1532 4233 1563
rect 4279 1532 4464 1563
rect 4048 1439 4464 1532
rect 4048 1408 4233 1439
rect 4279 1408 4464 1439
rect 4048 1315 4464 1408
rect 4048 1284 4233 1315
rect 4279 1284 4464 1315
rect 4048 1265 4464 1284
rect 4496 1812 4912 1830
rect 4496 1781 4681 1812
rect 4727 1781 4912 1812
rect 4496 1687 4912 1781
rect 4496 1656 4681 1687
rect 4727 1656 4912 1687
rect 4496 1563 4912 1656
rect 4496 1532 4681 1563
rect 4727 1532 4912 1563
rect 4496 1439 4912 1532
rect 4496 1408 4681 1439
rect 4727 1408 4912 1439
rect 4496 1315 4912 1408
rect 4496 1284 4681 1315
rect 4727 1284 4912 1315
rect 4496 1265 4912 1284
rect 4944 1812 5360 1830
rect 4944 1781 5129 1812
rect 5175 1781 5360 1812
rect 4944 1687 5360 1781
rect 4944 1656 5129 1687
rect 5175 1656 5360 1687
rect 4944 1563 5360 1656
rect 4944 1532 5129 1563
rect 5175 1551 5360 1563
rect 5392 1812 5808 1830
rect 5392 1781 5577 1812
rect 5623 1781 5808 1812
rect 5392 1687 5808 1781
rect 5392 1656 5577 1687
rect 5623 1656 5808 1687
rect 5392 1563 5808 1656
rect 5392 1551 5577 1563
rect 5175 1532 5577 1551
rect 5623 1556 5808 1563
rect 5840 1812 6256 1830
rect 5840 1781 6025 1812
rect 6071 1781 6256 1812
rect 5840 1687 6256 1781
rect 5840 1656 6025 1687
rect 6071 1656 6256 1687
rect 5840 1563 6256 1656
rect 5840 1556 6025 1563
rect 5623 1537 6025 1556
rect 5623 1532 5808 1537
rect 4944 1439 5360 1532
rect 4944 1408 5129 1439
rect 5175 1408 5360 1439
rect 4944 1315 5360 1408
rect 4944 1284 5129 1315
rect 5175 1284 5360 1315
rect 4944 1265 5360 1284
rect 5392 1439 5808 1532
rect 5392 1408 5577 1439
rect 5623 1408 5808 1439
rect 5392 1315 5808 1408
rect 5392 1284 5577 1315
rect 5623 1284 5808 1315
rect 5392 1265 5808 1284
rect 5840 1532 6025 1537
rect 6071 1532 6256 1563
rect 5840 1439 6256 1532
rect 5840 1408 6025 1439
rect 6071 1408 6256 1439
rect 5840 1315 6256 1408
rect 5840 1284 6025 1315
rect 6071 1284 6256 1315
rect 5840 1265 6256 1284
rect 6288 1812 6704 1830
rect 6288 1781 6473 1812
rect 6519 1781 6704 1812
rect 6288 1687 6704 1781
rect 6288 1656 6473 1687
rect 6519 1656 6704 1687
rect 6288 1563 6704 1656
rect 6288 1532 6473 1563
rect 6519 1532 6704 1563
rect 6288 1439 6704 1532
rect 6288 1408 6473 1439
rect 6519 1408 6704 1439
rect 6288 1315 6704 1408
rect 6288 1284 6473 1315
rect 6519 1284 6704 1315
rect 6288 1265 6704 1284
rect 6736 1812 7152 1830
rect 6736 1781 6921 1812
rect 6967 1781 7152 1812
rect 6736 1687 7152 1781
rect 6736 1656 6921 1687
rect 6967 1656 7152 1687
rect 6736 1563 7152 1656
rect 6736 1532 6921 1563
rect 6967 1532 7152 1563
rect 6736 1439 7152 1532
rect 6736 1408 6921 1439
rect 6967 1408 7152 1439
rect 6736 1315 7152 1408
rect 6736 1284 6921 1315
rect 6967 1284 7152 1315
rect 6736 1265 7152 1284
rect 7184 1812 7600 1830
rect 7184 1781 7369 1812
rect 7415 1781 7600 1812
rect 7184 1687 7600 1781
rect 7184 1656 7369 1687
rect 7415 1656 7600 1687
rect 7184 1563 7600 1656
rect 7184 1532 7369 1563
rect 7415 1551 7600 1563
rect 7632 1812 8048 1830
rect 7632 1781 7817 1812
rect 7863 1781 8048 1812
rect 7632 1687 8048 1781
rect 7632 1656 7817 1687
rect 7863 1656 8048 1687
rect 7632 1563 8048 1656
rect 7632 1551 7817 1563
rect 7415 1532 7817 1551
rect 7863 1556 8048 1563
rect 8080 1812 8496 1830
rect 8080 1781 8265 1812
rect 8311 1781 8496 1812
rect 8080 1687 8496 1781
rect 8080 1656 8265 1687
rect 8311 1656 8496 1687
rect 8080 1563 8496 1656
rect 8080 1556 8265 1563
rect 7863 1537 8265 1556
rect 7863 1532 8048 1537
rect 7184 1439 7600 1532
rect 7184 1408 7369 1439
rect 7415 1408 7600 1439
rect 7184 1315 7600 1408
rect 7184 1284 7369 1315
rect 7415 1284 7600 1315
rect 7184 1265 7600 1284
rect 7632 1439 8048 1532
rect 7632 1408 7817 1439
rect 7863 1408 8048 1439
rect 7632 1315 8048 1408
rect 7632 1284 7817 1315
rect 7863 1284 8048 1315
rect 7632 1265 8048 1284
rect 8080 1532 8265 1537
rect 8311 1532 8496 1563
rect 8080 1439 8496 1532
rect 8080 1408 8265 1439
rect 8311 1408 8496 1439
rect 8080 1315 8496 1408
rect 8080 1284 8265 1315
rect 8311 1284 8496 1315
rect 8080 1265 8496 1284
rect 8528 1812 8944 1830
rect 8528 1781 8713 1812
rect 8759 1781 8944 1812
rect 8528 1687 8944 1781
rect 8528 1656 8713 1687
rect 8759 1656 8944 1687
rect 8528 1563 8944 1656
rect 8528 1532 8713 1563
rect 8759 1532 8944 1563
rect 8528 1439 8944 1532
rect 8528 1408 8713 1439
rect 8759 1408 8944 1439
rect 8528 1315 8944 1408
rect 8528 1284 8713 1315
rect 8759 1284 8944 1315
rect 8528 1265 8944 1284
rect 212 1211 233 1265
rect 1113 1211 1127 1265
rect 2004 1211 2027 1265
rect 2452 1211 2473 1265
rect 3353 1211 3367 1265
rect 4244 1211 4267 1265
rect 4692 1211 4713 1265
rect 5593 1211 5607 1265
rect 6484 1211 6507 1265
rect 6932 1211 6953 1265
rect 7833 1211 7847 1265
rect 8724 1211 8747 1265
rect 16 1193 432 1211
rect 16 1162 201 1193
rect 247 1162 432 1193
rect 16 1068 432 1162
rect 16 1037 201 1068
rect 247 1037 432 1068
rect 16 944 432 1037
rect 16 913 201 944
rect 247 913 432 944
rect 16 820 432 913
rect 16 789 201 820
rect 247 789 432 820
rect 16 696 432 789
rect 16 665 201 696
rect 247 665 432 696
rect 16 646 432 665
rect 464 1193 880 1211
rect 464 1162 649 1193
rect 695 1162 880 1193
rect 464 1068 880 1162
rect 464 1037 649 1068
rect 695 1037 880 1068
rect 464 944 880 1037
rect 464 913 649 944
rect 695 936 880 944
rect 912 1193 1328 1211
rect 912 1162 1097 1193
rect 1143 1162 1328 1193
rect 912 1068 1328 1162
rect 912 1037 1097 1068
rect 1143 1037 1328 1068
rect 912 944 1328 1037
rect 912 936 1097 944
rect 695 915 1097 936
rect 695 913 880 915
rect 464 820 880 913
rect 464 789 649 820
rect 695 789 880 820
rect 464 696 880 789
rect 464 665 649 696
rect 695 665 880 696
rect 464 646 880 665
rect 912 913 1097 915
rect 1143 938 1328 944
rect 1360 1193 1776 1211
rect 1360 1162 1545 1193
rect 1591 1162 1776 1193
rect 1360 1068 1776 1162
rect 1360 1037 1545 1068
rect 1591 1037 1776 1068
rect 1360 944 1776 1037
rect 1360 938 1545 944
rect 1143 917 1545 938
rect 1143 913 1328 917
rect 912 820 1328 913
rect 912 789 1097 820
rect 1143 789 1328 820
rect 912 696 1328 789
rect 912 665 1097 696
rect 1143 665 1328 696
rect 912 646 1328 665
rect 1360 913 1545 917
rect 1591 913 1776 944
rect 1360 820 1776 913
rect 1360 789 1545 820
rect 1591 789 1776 820
rect 1360 696 1776 789
rect 1360 665 1545 696
rect 1591 665 1776 696
rect 1360 646 1776 665
rect 1808 1193 2224 1211
rect 1808 1162 1993 1193
rect 2039 1162 2224 1193
rect 1808 1068 2224 1162
rect 1808 1037 1993 1068
rect 2039 1037 2224 1068
rect 1808 944 2224 1037
rect 1808 913 1993 944
rect 2039 913 2224 944
rect 1808 820 2224 913
rect 1808 789 1993 820
rect 2039 789 2224 820
rect 1808 696 2224 789
rect 1808 665 1993 696
rect 2039 665 2224 696
rect 1808 646 2224 665
rect 2256 1193 2672 1211
rect 2256 1162 2441 1193
rect 2487 1162 2672 1193
rect 2256 1068 2672 1162
rect 2256 1037 2441 1068
rect 2487 1037 2672 1068
rect 2256 944 2672 1037
rect 2256 913 2441 944
rect 2487 913 2672 944
rect 2256 820 2672 913
rect 2256 789 2441 820
rect 2487 789 2672 820
rect 2256 696 2672 789
rect 2256 665 2441 696
rect 2487 665 2672 696
rect 2256 646 2672 665
rect 2704 1193 3120 1211
rect 2704 1162 2889 1193
rect 2935 1162 3120 1193
rect 2704 1068 3120 1162
rect 2704 1037 2889 1068
rect 2935 1037 3120 1068
rect 2704 944 3120 1037
rect 2704 913 2889 944
rect 2935 936 3120 944
rect 3152 1193 3568 1211
rect 3152 1162 3337 1193
rect 3383 1162 3568 1193
rect 3152 1068 3568 1162
rect 3152 1037 3337 1068
rect 3383 1037 3568 1068
rect 3152 944 3568 1037
rect 3152 936 3337 944
rect 2935 915 3337 936
rect 2935 913 3120 915
rect 2704 820 3120 913
rect 2704 789 2889 820
rect 2935 789 3120 820
rect 2704 696 3120 789
rect 2704 665 2889 696
rect 2935 665 3120 696
rect 2704 646 3120 665
rect 3152 913 3337 915
rect 3383 938 3568 944
rect 3600 1193 4016 1211
rect 3600 1162 3785 1193
rect 3831 1162 4016 1193
rect 3600 1068 4016 1162
rect 3600 1037 3785 1068
rect 3831 1037 4016 1068
rect 3600 944 4016 1037
rect 3600 938 3785 944
rect 3383 917 3785 938
rect 3383 913 3568 917
rect 3152 820 3568 913
rect 3152 789 3337 820
rect 3383 789 3568 820
rect 3152 696 3568 789
rect 3152 665 3337 696
rect 3383 665 3568 696
rect 3152 646 3568 665
rect 3600 913 3785 917
rect 3831 913 4016 944
rect 3600 820 4016 913
rect 3600 789 3785 820
rect 3831 789 4016 820
rect 3600 696 4016 789
rect 3600 665 3785 696
rect 3831 665 4016 696
rect 3600 646 4016 665
rect 4048 1193 4464 1211
rect 4048 1162 4233 1193
rect 4279 1162 4464 1193
rect 4048 1068 4464 1162
rect 4048 1037 4233 1068
rect 4279 1037 4464 1068
rect 4048 944 4464 1037
rect 4048 913 4233 944
rect 4279 913 4464 944
rect 4048 820 4464 913
rect 4048 789 4233 820
rect 4279 789 4464 820
rect 4048 696 4464 789
rect 4048 665 4233 696
rect 4279 665 4464 696
rect 4048 646 4464 665
rect 4496 1193 4912 1211
rect 4496 1162 4681 1193
rect 4727 1162 4912 1193
rect 4496 1068 4912 1162
rect 4496 1037 4681 1068
rect 4727 1037 4912 1068
rect 4496 944 4912 1037
rect 4496 913 4681 944
rect 4727 913 4912 944
rect 4496 820 4912 913
rect 4496 789 4681 820
rect 4727 789 4912 820
rect 4496 696 4912 789
rect 4496 665 4681 696
rect 4727 665 4912 696
rect 4496 646 4912 665
rect 4944 1193 5360 1211
rect 4944 1162 5129 1193
rect 5175 1162 5360 1193
rect 4944 1068 5360 1162
rect 4944 1037 5129 1068
rect 5175 1037 5360 1068
rect 4944 944 5360 1037
rect 4944 913 5129 944
rect 5175 936 5360 944
rect 5392 1193 5808 1211
rect 5392 1162 5577 1193
rect 5623 1162 5808 1193
rect 5392 1068 5808 1162
rect 5392 1037 5577 1068
rect 5623 1037 5808 1068
rect 5392 944 5808 1037
rect 5392 936 5577 944
rect 5175 915 5577 936
rect 5175 913 5360 915
rect 4944 820 5360 913
rect 4944 789 5129 820
rect 5175 789 5360 820
rect 4944 696 5360 789
rect 4944 665 5129 696
rect 5175 665 5360 696
rect 4944 646 5360 665
rect 5392 913 5577 915
rect 5623 938 5808 944
rect 5840 1193 6256 1211
rect 5840 1162 6025 1193
rect 6071 1162 6256 1193
rect 5840 1068 6256 1162
rect 5840 1037 6025 1068
rect 6071 1037 6256 1068
rect 5840 944 6256 1037
rect 5840 938 6025 944
rect 5623 917 6025 938
rect 5623 913 5808 917
rect 5392 820 5808 913
rect 5392 789 5577 820
rect 5623 789 5808 820
rect 5392 696 5808 789
rect 5392 665 5577 696
rect 5623 665 5808 696
rect 5392 646 5808 665
rect 5840 913 6025 917
rect 6071 913 6256 944
rect 5840 820 6256 913
rect 5840 789 6025 820
rect 6071 789 6256 820
rect 5840 696 6256 789
rect 5840 665 6025 696
rect 6071 665 6256 696
rect 5840 646 6256 665
rect 6288 1193 6704 1211
rect 6288 1162 6473 1193
rect 6519 1162 6704 1193
rect 6288 1068 6704 1162
rect 6288 1037 6473 1068
rect 6519 1037 6704 1068
rect 6288 944 6704 1037
rect 6288 913 6473 944
rect 6519 913 6704 944
rect 6288 820 6704 913
rect 6288 789 6473 820
rect 6519 789 6704 820
rect 6288 696 6704 789
rect 6288 665 6473 696
rect 6519 665 6704 696
rect 6288 646 6704 665
rect 6736 1193 7152 1211
rect 6736 1162 6921 1193
rect 6967 1162 7152 1193
rect 6736 1068 7152 1162
rect 6736 1037 6921 1068
rect 6967 1037 7152 1068
rect 6736 944 7152 1037
rect 6736 913 6921 944
rect 6967 913 7152 944
rect 6736 820 7152 913
rect 6736 789 6921 820
rect 6967 789 7152 820
rect 6736 696 7152 789
rect 6736 665 6921 696
rect 6967 665 7152 696
rect 6736 646 7152 665
rect 7184 1193 7600 1211
rect 7184 1162 7369 1193
rect 7415 1162 7600 1193
rect 7184 1068 7600 1162
rect 7184 1037 7369 1068
rect 7415 1037 7600 1068
rect 7184 944 7600 1037
rect 7184 913 7369 944
rect 7415 936 7600 944
rect 7632 1193 8048 1211
rect 7632 1162 7817 1193
rect 7863 1162 8048 1193
rect 7632 1068 8048 1162
rect 7632 1037 7817 1068
rect 7863 1037 8048 1068
rect 7632 944 8048 1037
rect 7632 936 7817 944
rect 7415 915 7817 936
rect 7415 913 7600 915
rect 7184 820 7600 913
rect 7184 789 7369 820
rect 7415 789 7600 820
rect 7184 696 7600 789
rect 7184 665 7369 696
rect 7415 665 7600 696
rect 7184 646 7600 665
rect 7632 913 7817 915
rect 7863 938 8048 944
rect 8080 1193 8496 1211
rect 8080 1162 8265 1193
rect 8311 1162 8496 1193
rect 8080 1068 8496 1162
rect 8080 1037 8265 1068
rect 8311 1037 8496 1068
rect 8080 944 8496 1037
rect 8080 938 8265 944
rect 7863 917 8265 938
rect 7863 913 8048 917
rect 7632 820 8048 913
rect 7632 789 7817 820
rect 7863 789 8048 820
rect 7632 696 8048 789
rect 7632 665 7817 696
rect 7863 665 8048 696
rect 7632 646 8048 665
rect 8080 913 8265 917
rect 8311 913 8496 944
rect 8080 820 8496 913
rect 8080 789 8265 820
rect 8311 789 8496 820
rect 8080 696 8496 789
rect 8080 665 8265 696
rect 8311 665 8496 696
rect 8080 646 8496 665
rect 8528 1193 8944 1211
rect 8528 1162 8713 1193
rect 8759 1162 8944 1193
rect 8528 1068 8944 1162
rect 8528 1037 8713 1068
rect 8759 1037 8944 1068
rect 8528 944 8944 1037
rect 8528 913 8713 944
rect 8759 913 8944 944
rect 8528 820 8944 913
rect 8528 789 8713 820
rect 8759 789 8944 820
rect 8528 696 8944 789
rect 8528 665 8713 696
rect 8759 665 8944 696
rect 8528 646 8944 665
rect 212 592 233 646
rect 2007 592 2030 646
rect 2452 592 2473 646
rect 3348 592 3375 646
rect 4247 592 4270 646
rect 4692 592 4713 646
rect 5586 592 5607 646
rect 6487 592 6510 646
rect 6932 592 6953 646
rect 7831 592 7847 646
rect 8727 592 8750 646
rect 16 574 432 592
rect 16 543 201 574
rect 247 543 432 574
rect 16 449 432 543
rect 16 418 201 449
rect 247 418 432 449
rect 16 325 432 418
rect 16 294 201 325
rect 247 312 432 325
rect 464 574 880 592
rect 464 543 649 574
rect 695 543 880 574
rect 464 449 880 543
rect 464 418 649 449
rect 695 418 880 449
rect 464 325 880 418
rect 464 312 649 325
rect 247 294 649 312
rect 695 317 880 325
rect 912 574 1328 592
rect 912 543 1097 574
rect 1143 543 1328 574
rect 912 449 1328 543
rect 912 418 1097 449
rect 1143 418 1328 449
rect 912 325 1328 418
rect 912 317 1097 325
rect 695 299 1097 317
rect 695 294 880 299
rect 16 292 880 294
rect 16 201 432 292
rect 16 170 201 201
rect 247 170 432 201
rect 16 77 432 170
rect 16 46 201 77
rect 247 46 432 77
rect 16 27 432 46
rect 464 201 880 292
rect 464 170 649 201
rect 695 170 880 201
rect 464 77 880 170
rect 464 46 649 77
rect 695 46 880 77
rect 464 27 880 46
rect 912 294 1097 299
rect 1143 316 1328 325
rect 1360 574 1776 592
rect 1360 543 1545 574
rect 1591 543 1776 574
rect 1360 449 1776 543
rect 1360 418 1545 449
rect 1591 418 1776 449
rect 1360 325 1776 418
rect 1360 316 1545 325
rect 1143 298 1545 316
rect 1143 294 1328 298
rect 912 201 1328 294
rect 912 170 1097 201
rect 1143 170 1328 201
rect 912 77 1328 170
rect 912 46 1097 77
rect 1143 46 1328 77
rect 912 27 1328 46
rect 1360 294 1545 298
rect 1591 294 1776 325
rect 1360 257 1776 294
rect 1808 574 2224 592
rect 1808 543 1993 574
rect 2039 543 2224 574
rect 1808 449 2224 543
rect 1808 418 1993 449
rect 2039 418 2224 449
rect 1808 325 2224 418
rect 1808 294 1993 325
rect 2039 294 2224 325
rect 1808 257 2224 294
rect 1360 237 2224 257
rect 1360 201 1776 237
rect 1360 170 1545 201
rect 1591 170 1776 201
rect 1360 77 1776 170
rect 1360 46 1545 77
rect 1591 46 1776 77
rect 1360 27 1776 46
rect 1808 201 2224 237
rect 1808 170 1993 201
rect 2039 170 2224 201
rect 1808 77 2224 170
rect 1808 46 1993 77
rect 2039 46 2224 77
rect 1808 27 2224 46
rect 2256 574 2672 592
rect 2256 543 2441 574
rect 2487 543 2672 574
rect 2256 449 2672 543
rect 2256 418 2441 449
rect 2487 418 2672 449
rect 2256 325 2672 418
rect 2256 294 2441 325
rect 2487 312 2672 325
rect 2704 574 3120 592
rect 2704 543 2889 574
rect 2935 543 3120 574
rect 2704 449 3120 543
rect 2704 418 2889 449
rect 2935 418 3120 449
rect 2704 325 3120 418
rect 2704 312 2889 325
rect 2487 294 2889 312
rect 2935 294 3120 325
rect 2256 292 3120 294
rect 2256 201 2672 292
rect 2256 170 2441 201
rect 2487 170 2672 201
rect 2256 77 2672 170
rect 2256 46 2441 77
rect 2487 46 2672 77
rect 2256 27 2672 46
rect 2704 201 3120 292
rect 2704 170 2889 201
rect 2935 170 3120 201
rect 2704 77 3120 170
rect 2704 46 2889 77
rect 2935 46 3120 77
rect 2704 27 3120 46
rect 3152 574 3568 592
rect 3152 543 3337 574
rect 3383 543 3568 574
rect 3152 449 3568 543
rect 3152 418 3337 449
rect 3383 418 3568 449
rect 3152 325 3568 418
rect 3152 294 3337 325
rect 3383 294 3568 325
rect 3152 201 3568 294
rect 3152 170 3337 201
rect 3383 170 3568 201
rect 3152 77 3568 170
rect 3152 46 3337 77
rect 3383 46 3568 77
rect 3152 27 3568 46
rect 3600 574 4016 592
rect 3600 543 3785 574
rect 3831 543 4016 574
rect 3600 449 4016 543
rect 3600 418 3785 449
rect 3831 418 4016 449
rect 3600 325 4016 418
rect 3600 294 3785 325
rect 3831 294 4016 325
rect 3600 257 4016 294
rect 4048 574 4464 592
rect 4048 543 4233 574
rect 4279 543 4464 574
rect 4048 449 4464 543
rect 4048 418 4233 449
rect 4279 418 4464 449
rect 4048 325 4464 418
rect 4048 294 4233 325
rect 4279 294 4464 325
rect 4048 257 4464 294
rect 3600 237 4464 257
rect 3600 201 4016 237
rect 3600 170 3785 201
rect 3831 170 4016 201
rect 3600 77 4016 170
rect 3600 46 3785 77
rect 3831 46 4016 77
rect 3600 27 4016 46
rect 4048 201 4464 237
rect 4048 170 4233 201
rect 4279 170 4464 201
rect 4048 77 4464 170
rect 4048 46 4233 77
rect 4279 46 4464 77
rect 4048 27 4464 46
rect 4496 574 4912 592
rect 4496 543 4681 574
rect 4727 543 4912 574
rect 4496 449 4912 543
rect 4496 418 4681 449
rect 4727 418 4912 449
rect 4496 325 4912 418
rect 4496 294 4681 325
rect 4727 312 4912 325
rect 4944 574 5360 592
rect 4944 543 5129 574
rect 5175 543 5360 574
rect 4944 449 5360 543
rect 4944 418 5129 449
rect 5175 418 5360 449
rect 4944 325 5360 418
rect 4944 312 5129 325
rect 4727 294 5129 312
rect 5175 294 5360 325
rect 4496 292 5360 294
rect 4496 201 4912 292
rect 4496 170 4681 201
rect 4727 170 4912 201
rect 4496 77 4912 170
rect 4496 46 4681 77
rect 4727 46 4912 77
rect 4496 27 4912 46
rect 4944 201 5360 292
rect 4944 170 5129 201
rect 5175 170 5360 201
rect 4944 77 5360 170
rect 4944 46 5129 77
rect 5175 46 5360 77
rect 4944 27 5360 46
rect 5392 574 5808 592
rect 5392 543 5577 574
rect 5623 543 5808 574
rect 5392 449 5808 543
rect 5392 418 5577 449
rect 5623 418 5808 449
rect 5392 325 5808 418
rect 5392 294 5577 325
rect 5623 294 5808 325
rect 5392 201 5808 294
rect 5392 170 5577 201
rect 5623 170 5808 201
rect 5392 77 5808 170
rect 5392 46 5577 77
rect 5623 46 5808 77
rect 5392 27 5808 46
rect 5840 574 6256 592
rect 5840 543 6025 574
rect 6071 543 6256 574
rect 5840 449 6256 543
rect 5840 418 6025 449
rect 6071 418 6256 449
rect 5840 325 6256 418
rect 5840 294 6025 325
rect 6071 294 6256 325
rect 5840 257 6256 294
rect 6288 574 6704 592
rect 6288 543 6473 574
rect 6519 543 6704 574
rect 6288 449 6704 543
rect 6288 418 6473 449
rect 6519 418 6704 449
rect 6288 325 6704 418
rect 6288 294 6473 325
rect 6519 294 6704 325
rect 6288 257 6704 294
rect 5840 237 6704 257
rect 5840 201 6256 237
rect 5840 170 6025 201
rect 6071 170 6256 201
rect 5840 77 6256 170
rect 5840 46 6025 77
rect 6071 46 6256 77
rect 5840 27 6256 46
rect 6288 201 6704 237
rect 6288 170 6473 201
rect 6519 170 6704 201
rect 6288 77 6704 170
rect 6288 46 6473 77
rect 6519 46 6704 77
rect 6288 27 6704 46
rect 6736 574 7152 592
rect 6736 543 6921 574
rect 6967 543 7152 574
rect 6736 449 7152 543
rect 6736 418 6921 449
rect 6967 418 7152 449
rect 6736 325 7152 418
rect 6736 294 6921 325
rect 6967 312 7152 325
rect 7184 574 7600 592
rect 7184 543 7369 574
rect 7415 543 7600 574
rect 7184 449 7600 543
rect 7184 418 7369 449
rect 7415 418 7600 449
rect 7184 325 7600 418
rect 7184 312 7369 325
rect 6967 294 7369 312
rect 7415 294 7600 325
rect 6736 292 7600 294
rect 6736 201 7152 292
rect 6736 170 6921 201
rect 6967 170 7152 201
rect 6736 77 7152 170
rect 6736 46 6921 77
rect 6967 46 7152 77
rect 6736 27 7152 46
rect 7184 201 7600 292
rect 7184 170 7369 201
rect 7415 170 7600 201
rect 7184 77 7600 170
rect 7184 46 7369 77
rect 7415 46 7600 77
rect 7184 27 7600 46
rect 7632 574 8048 592
rect 7632 543 7817 574
rect 7863 543 8048 574
rect 7632 449 8048 543
rect 7632 418 7817 449
rect 7863 418 8048 449
rect 7632 325 8048 418
rect 7632 294 7817 325
rect 7863 294 8048 325
rect 7632 201 8048 294
rect 7632 170 7817 201
rect 7863 170 8048 201
rect 7632 77 8048 170
rect 7632 46 7817 77
rect 7863 46 8048 77
rect 7632 27 8048 46
rect 8080 574 8496 592
rect 8080 543 8265 574
rect 8311 543 8496 574
rect 8080 449 8496 543
rect 8080 418 8265 449
rect 8311 418 8496 449
rect 8080 325 8496 418
rect 8080 294 8265 325
rect 8311 294 8496 325
rect 8080 257 8496 294
rect 8528 574 8944 592
rect 8528 543 8713 574
rect 8759 543 8944 574
rect 8528 449 8944 543
rect 8528 418 8713 449
rect 8759 418 8944 449
rect 8528 325 8944 418
rect 8528 294 8713 325
rect 8759 294 8944 325
rect 8528 257 8944 294
rect 8080 237 8944 257
rect 8080 201 8496 237
rect 8080 170 8265 201
rect 8311 170 8496 201
rect 8080 77 8496 170
rect 8080 46 8265 77
rect 8311 46 8496 77
rect 8080 27 8496 46
rect 8528 201 8944 237
rect 8528 170 8713 201
rect 8759 170 8944 201
rect 8528 77 8944 170
rect 8528 46 8713 77
rect 8759 46 8944 77
rect 8528 27 8944 46
<< via2 >>
rect 201 2400 247 2431
rect 201 2275 247 2306
rect 201 2151 247 2182
rect 649 2400 695 2431
rect 649 2275 695 2306
rect 201 2027 247 2058
rect 201 1903 247 1934
rect 649 2151 695 2182
rect 1097 2400 1143 2431
rect 1097 2275 1143 2306
rect 649 2027 695 2058
rect 649 1903 695 1934
rect 1097 2151 1143 2182
rect 1545 2400 1591 2431
rect 1545 2275 1591 2306
rect 1097 2027 1143 2058
rect 1097 1903 1143 1934
rect 1545 2151 1591 2182
rect 1993 2400 2039 2431
rect 1993 2275 2039 2306
rect 1545 2027 1591 2058
rect 1545 1903 1591 1934
rect 1993 2151 2039 2182
rect 2441 2400 2487 2431
rect 2441 2275 2487 2306
rect 1993 2027 2039 2058
rect 1993 1903 2039 1934
rect 2441 2151 2487 2182
rect 2889 2400 2935 2431
rect 2889 2275 2935 2306
rect 2441 2027 2487 2058
rect 2441 1903 2487 1934
rect 2889 2151 2935 2182
rect 3337 2400 3383 2431
rect 3337 2275 3383 2306
rect 2889 2027 2935 2058
rect 2889 1903 2935 1934
rect 3337 2151 3383 2182
rect 3785 2400 3831 2431
rect 3785 2275 3831 2306
rect 3337 2027 3383 2058
rect 3337 1903 3383 1934
rect 3785 2151 3831 2182
rect 4233 2400 4279 2431
rect 4233 2275 4279 2306
rect 3785 2027 3831 2058
rect 3785 1903 3831 1934
rect 4233 2151 4279 2182
rect 4681 2400 4727 2431
rect 4681 2275 4727 2306
rect 4233 2027 4279 2058
rect 4233 1903 4279 1934
rect 4681 2151 4727 2182
rect 5129 2400 5175 2431
rect 5129 2275 5175 2306
rect 4681 2027 4727 2058
rect 4681 1903 4727 1934
rect 5129 2151 5175 2182
rect 5577 2400 5623 2431
rect 5577 2275 5623 2306
rect 5129 2027 5175 2058
rect 5129 1903 5175 1934
rect 5577 2151 5623 2182
rect 6025 2400 6071 2431
rect 6025 2275 6071 2306
rect 5577 2027 5623 2058
rect 5577 1903 5623 1934
rect 6025 2151 6071 2182
rect 6473 2400 6519 2431
rect 6473 2275 6519 2306
rect 6025 2027 6071 2058
rect 6025 1903 6071 1934
rect 6473 2151 6519 2182
rect 6921 2400 6967 2431
rect 6921 2275 6967 2306
rect 6473 2027 6519 2058
rect 6473 1903 6519 1934
rect 6921 2151 6967 2182
rect 7369 2400 7415 2431
rect 7369 2275 7415 2306
rect 6921 2027 6967 2058
rect 6921 1903 6967 1934
rect 7369 2151 7415 2182
rect 7817 2400 7863 2431
rect 7817 2275 7863 2306
rect 7369 2027 7415 2058
rect 7369 1903 7415 1934
rect 7817 2151 7863 2182
rect 8265 2400 8311 2431
rect 8265 2275 8311 2306
rect 7817 2027 7863 2058
rect 7817 1903 7863 1934
rect 8265 2151 8311 2182
rect 8713 2400 8759 2431
rect 8713 2275 8759 2306
rect 8265 2027 8311 2058
rect 8265 1903 8311 1934
rect 8713 2151 8759 2182
rect 8713 2027 8759 2058
rect 8713 1903 8759 1934
rect 201 1781 247 1812
rect 201 1656 247 1687
rect 201 1532 247 1563
rect 201 1408 247 1439
rect 201 1284 247 1315
rect 649 1781 695 1812
rect 649 1656 695 1687
rect 649 1532 695 1563
rect 1097 1781 1143 1812
rect 1097 1656 1143 1687
rect 1097 1532 1143 1563
rect 1545 1781 1591 1812
rect 1545 1656 1591 1687
rect 649 1408 695 1439
rect 649 1284 695 1315
rect 1097 1408 1143 1439
rect 1097 1284 1143 1315
rect 1545 1532 1591 1563
rect 1545 1408 1591 1439
rect 1545 1284 1591 1315
rect 1993 1781 2039 1812
rect 1993 1656 2039 1687
rect 1993 1532 2039 1563
rect 1993 1408 2039 1439
rect 1993 1284 2039 1315
rect 2441 1781 2487 1812
rect 2441 1656 2487 1687
rect 2441 1532 2487 1563
rect 2441 1408 2487 1439
rect 2441 1284 2487 1315
rect 2889 1781 2935 1812
rect 2889 1656 2935 1687
rect 2889 1532 2935 1563
rect 3337 1781 3383 1812
rect 3337 1656 3383 1687
rect 3337 1532 3383 1563
rect 3785 1781 3831 1812
rect 3785 1656 3831 1687
rect 2889 1408 2935 1439
rect 2889 1284 2935 1315
rect 3337 1408 3383 1439
rect 3337 1284 3383 1315
rect 3785 1532 3831 1563
rect 3785 1408 3831 1439
rect 3785 1284 3831 1315
rect 4233 1781 4279 1812
rect 4233 1656 4279 1687
rect 4233 1532 4279 1563
rect 4233 1408 4279 1439
rect 4233 1284 4279 1315
rect 4681 1781 4727 1812
rect 4681 1656 4727 1687
rect 4681 1532 4727 1563
rect 4681 1408 4727 1439
rect 4681 1284 4727 1315
rect 5129 1781 5175 1812
rect 5129 1656 5175 1687
rect 5129 1532 5175 1563
rect 5577 1781 5623 1812
rect 5577 1656 5623 1687
rect 5577 1532 5623 1563
rect 6025 1781 6071 1812
rect 6025 1656 6071 1687
rect 5129 1408 5175 1439
rect 5129 1284 5175 1315
rect 5577 1408 5623 1439
rect 5577 1284 5623 1315
rect 6025 1532 6071 1563
rect 6025 1408 6071 1439
rect 6025 1284 6071 1315
rect 6473 1781 6519 1812
rect 6473 1656 6519 1687
rect 6473 1532 6519 1563
rect 6473 1408 6519 1439
rect 6473 1284 6519 1315
rect 6921 1781 6967 1812
rect 6921 1656 6967 1687
rect 6921 1532 6967 1563
rect 6921 1408 6967 1439
rect 6921 1284 6967 1315
rect 7369 1781 7415 1812
rect 7369 1656 7415 1687
rect 7369 1532 7415 1563
rect 7817 1781 7863 1812
rect 7817 1656 7863 1687
rect 7817 1532 7863 1563
rect 8265 1781 8311 1812
rect 8265 1656 8311 1687
rect 7369 1408 7415 1439
rect 7369 1284 7415 1315
rect 7817 1408 7863 1439
rect 7817 1284 7863 1315
rect 8265 1532 8311 1563
rect 8265 1408 8311 1439
rect 8265 1284 8311 1315
rect 8713 1781 8759 1812
rect 8713 1656 8759 1687
rect 8713 1532 8759 1563
rect 8713 1408 8759 1439
rect 8713 1284 8759 1315
rect 201 1162 247 1193
rect 201 1037 247 1068
rect 201 913 247 944
rect 201 789 247 820
rect 201 665 247 696
rect 649 1162 695 1193
rect 649 1037 695 1068
rect 649 913 695 944
rect 1097 1162 1143 1193
rect 1097 1037 1143 1068
rect 649 789 695 820
rect 649 665 695 696
rect 1097 913 1143 944
rect 1545 1162 1591 1193
rect 1545 1037 1591 1068
rect 1097 789 1143 820
rect 1097 665 1143 696
rect 1545 913 1591 944
rect 1545 789 1591 820
rect 1545 665 1591 696
rect 1993 1162 2039 1193
rect 1993 1037 2039 1068
rect 1993 913 2039 944
rect 1993 789 2039 820
rect 1993 665 2039 696
rect 2441 1162 2487 1193
rect 2441 1037 2487 1068
rect 2441 913 2487 944
rect 2441 789 2487 820
rect 2441 665 2487 696
rect 2889 1162 2935 1193
rect 2889 1037 2935 1068
rect 2889 913 2935 944
rect 3337 1162 3383 1193
rect 3337 1037 3383 1068
rect 2889 789 2935 820
rect 2889 665 2935 696
rect 3337 913 3383 944
rect 3785 1162 3831 1193
rect 3785 1037 3831 1068
rect 3337 789 3383 820
rect 3337 665 3383 696
rect 3785 913 3831 944
rect 3785 789 3831 820
rect 3785 665 3831 696
rect 4233 1162 4279 1193
rect 4233 1037 4279 1068
rect 4233 913 4279 944
rect 4233 789 4279 820
rect 4233 665 4279 696
rect 4681 1162 4727 1193
rect 4681 1037 4727 1068
rect 4681 913 4727 944
rect 4681 789 4727 820
rect 4681 665 4727 696
rect 5129 1162 5175 1193
rect 5129 1037 5175 1068
rect 5129 913 5175 944
rect 5577 1162 5623 1193
rect 5577 1037 5623 1068
rect 5129 789 5175 820
rect 5129 665 5175 696
rect 5577 913 5623 944
rect 6025 1162 6071 1193
rect 6025 1037 6071 1068
rect 5577 789 5623 820
rect 5577 665 5623 696
rect 6025 913 6071 944
rect 6025 789 6071 820
rect 6025 665 6071 696
rect 6473 1162 6519 1193
rect 6473 1037 6519 1068
rect 6473 913 6519 944
rect 6473 789 6519 820
rect 6473 665 6519 696
rect 6921 1162 6967 1193
rect 6921 1037 6967 1068
rect 6921 913 6967 944
rect 6921 789 6967 820
rect 6921 665 6967 696
rect 7369 1162 7415 1193
rect 7369 1037 7415 1068
rect 7369 913 7415 944
rect 7817 1162 7863 1193
rect 7817 1037 7863 1068
rect 7369 789 7415 820
rect 7369 665 7415 696
rect 7817 913 7863 944
rect 8265 1162 8311 1193
rect 8265 1037 8311 1068
rect 7817 789 7863 820
rect 7817 665 7863 696
rect 8265 913 8311 944
rect 8265 789 8311 820
rect 8265 665 8311 696
rect 8713 1162 8759 1193
rect 8713 1037 8759 1068
rect 8713 913 8759 944
rect 8713 789 8759 820
rect 8713 665 8759 696
rect 201 543 247 574
rect 201 418 247 449
rect 201 294 247 325
rect 649 543 695 574
rect 649 418 695 449
rect 649 294 695 325
rect 1097 543 1143 574
rect 1097 418 1143 449
rect 201 170 247 201
rect 201 46 247 77
rect 649 170 695 201
rect 649 46 695 77
rect 1097 294 1143 325
rect 1545 543 1591 574
rect 1545 418 1591 449
rect 1097 170 1143 201
rect 1097 46 1143 77
rect 1545 294 1591 325
rect 1993 543 2039 574
rect 1993 418 2039 449
rect 1993 294 2039 325
rect 1545 170 1591 201
rect 1545 46 1591 77
rect 1993 170 2039 201
rect 1993 46 2039 77
rect 2441 543 2487 574
rect 2441 418 2487 449
rect 2441 294 2487 325
rect 2889 543 2935 574
rect 2889 418 2935 449
rect 2889 294 2935 325
rect 2441 170 2487 201
rect 2441 46 2487 77
rect 2889 170 2935 201
rect 2889 46 2935 77
rect 3337 543 3383 574
rect 3337 418 3383 449
rect 3337 294 3383 325
rect 3337 170 3383 201
rect 3337 46 3383 77
rect 3785 543 3831 574
rect 3785 418 3831 449
rect 3785 294 3831 325
rect 4233 543 4279 574
rect 4233 418 4279 449
rect 4233 294 4279 325
rect 3785 170 3831 201
rect 3785 46 3831 77
rect 4233 170 4279 201
rect 4233 46 4279 77
rect 4681 543 4727 574
rect 4681 418 4727 449
rect 4681 294 4727 325
rect 5129 543 5175 574
rect 5129 418 5175 449
rect 5129 294 5175 325
rect 4681 170 4727 201
rect 4681 46 4727 77
rect 5129 170 5175 201
rect 5129 46 5175 77
rect 5577 543 5623 574
rect 5577 418 5623 449
rect 5577 294 5623 325
rect 5577 170 5623 201
rect 5577 46 5623 77
rect 6025 543 6071 574
rect 6025 418 6071 449
rect 6025 294 6071 325
rect 6473 543 6519 574
rect 6473 418 6519 449
rect 6473 294 6519 325
rect 6025 170 6071 201
rect 6025 46 6071 77
rect 6473 170 6519 201
rect 6473 46 6519 77
rect 6921 543 6967 574
rect 6921 418 6967 449
rect 6921 294 6967 325
rect 7369 543 7415 574
rect 7369 418 7415 449
rect 7369 294 7415 325
rect 6921 170 6967 201
rect 6921 46 6967 77
rect 7369 170 7415 201
rect 7369 46 7415 77
rect 7817 543 7863 574
rect 7817 418 7863 449
rect 7817 294 7863 325
rect 7817 170 7863 201
rect 7817 46 7863 77
rect 8265 543 8311 574
rect 8265 418 8311 449
rect 8265 294 8311 325
rect 8713 543 8759 574
rect 8713 418 8759 449
rect 8713 294 8759 325
rect 8265 170 8311 201
rect 8265 46 8311 77
rect 8713 170 8759 201
rect 8713 46 8759 77
<< metal3 >>
rect 196 2431 252 2434
rect 196 2430 201 2431
rect 35 2400 201 2430
rect 247 2430 252 2431
rect 644 2431 700 2434
rect 644 2430 649 2431
rect 247 2400 413 2430
rect 483 2400 649 2430
rect 695 2430 700 2431
rect 1092 2431 1148 2434
rect 1092 2430 1097 2431
rect 695 2400 861 2430
rect 931 2400 1097 2430
rect 1143 2430 1148 2431
rect 1540 2431 1596 2434
rect 1540 2430 1545 2431
rect 1143 2400 1309 2430
rect 1379 2400 1545 2430
rect 1591 2430 1596 2431
rect 1988 2431 2044 2434
rect 1988 2430 1993 2431
rect 1591 2400 1757 2430
rect 1827 2400 1993 2430
rect 2039 2430 2044 2431
rect 2436 2431 2492 2434
rect 2436 2430 2441 2431
rect 2039 2400 2205 2430
rect 2275 2400 2441 2430
rect 2487 2430 2492 2431
rect 2884 2431 2940 2434
rect 2884 2430 2889 2431
rect 2487 2400 2653 2430
rect 2723 2400 2889 2430
rect 2935 2430 2940 2431
rect 3332 2431 3388 2434
rect 3332 2430 3337 2431
rect 2935 2400 3101 2430
rect 3171 2400 3337 2430
rect 3383 2430 3388 2431
rect 3780 2431 3836 2434
rect 3780 2430 3785 2431
rect 3383 2400 3549 2430
rect 3619 2400 3785 2430
rect 3831 2430 3836 2431
rect 4228 2431 4284 2434
rect 4228 2430 4233 2431
rect 3831 2400 3997 2430
rect 4067 2400 4233 2430
rect 4279 2430 4284 2431
rect 4676 2431 4732 2434
rect 4676 2430 4681 2431
rect 4279 2400 4445 2430
rect 4515 2400 4681 2430
rect 4727 2430 4732 2431
rect 5124 2431 5180 2434
rect 5124 2430 5129 2431
rect 4727 2400 4893 2430
rect 4963 2400 5129 2430
rect 5175 2430 5180 2431
rect 5572 2431 5628 2434
rect 5572 2430 5577 2431
rect 5175 2400 5341 2430
rect 5411 2400 5577 2430
rect 5623 2430 5628 2431
rect 6020 2431 6076 2434
rect 6020 2430 6025 2431
rect 5623 2400 5789 2430
rect 5859 2400 6025 2430
rect 6071 2430 6076 2431
rect 6468 2431 6524 2434
rect 6468 2430 6473 2431
rect 6071 2400 6237 2430
rect 6307 2400 6473 2430
rect 6519 2430 6524 2431
rect 6916 2431 6972 2434
rect 6916 2430 6921 2431
rect 6519 2400 6685 2430
rect 6755 2400 6921 2430
rect 6967 2430 6972 2431
rect 7364 2431 7420 2434
rect 7364 2430 7369 2431
rect 6967 2400 7133 2430
rect 7203 2400 7369 2430
rect 7415 2430 7420 2431
rect 7812 2431 7868 2434
rect 7812 2430 7817 2431
rect 7415 2400 7581 2430
rect 7651 2400 7817 2430
rect 7863 2430 7868 2431
rect 8260 2431 8316 2434
rect 8260 2430 8265 2431
rect 7863 2400 8029 2430
rect 8099 2400 8265 2430
rect 8311 2430 8316 2431
rect 8708 2431 8764 2434
rect 8708 2430 8713 2431
rect 8311 2400 8477 2430
rect 8547 2400 8713 2430
rect 8759 2430 8764 2431
rect 8759 2400 8925 2430
rect 196 2396 252 2400
rect 644 2396 700 2400
rect 1092 2396 1148 2400
rect 1540 2396 1596 2400
rect 1988 2396 2044 2400
rect 2436 2396 2492 2400
rect 2884 2396 2940 2400
rect 3332 2396 3388 2400
rect 3780 2396 3836 2400
rect 4228 2396 4284 2400
rect 4676 2396 4732 2400
rect 5124 2396 5180 2400
rect 5572 2396 5628 2400
rect 6020 2396 6076 2400
rect 6468 2396 6524 2400
rect 6916 2396 6972 2400
rect 7364 2396 7420 2400
rect 7812 2396 7868 2400
rect 8260 2396 8316 2400
rect 8708 2396 8764 2400
rect 99 2368 137 2369
rect 99 2367 102 2368
rect 54 2337 102 2367
rect 99 2336 102 2337
rect 134 2367 137 2368
rect 311 2368 349 2369
rect 311 2367 314 2368
rect 134 2337 181 2367
rect 267 2337 314 2367
rect 134 2336 137 2337
rect 99 2335 137 2336
rect 311 2336 314 2337
rect 346 2367 349 2368
rect 547 2368 585 2369
rect 547 2367 550 2368
rect 346 2337 394 2367
rect 502 2337 550 2367
rect 346 2336 349 2337
rect 311 2335 349 2336
rect 547 2336 550 2337
rect 582 2367 585 2368
rect 759 2368 797 2369
rect 759 2367 762 2368
rect 582 2337 629 2367
rect 715 2337 762 2367
rect 582 2336 585 2337
rect 547 2335 585 2336
rect 759 2336 762 2337
rect 794 2367 797 2368
rect 995 2368 1033 2369
rect 995 2367 998 2368
rect 794 2337 842 2367
rect 950 2337 998 2367
rect 794 2336 797 2337
rect 759 2335 797 2336
rect 995 2336 998 2337
rect 1030 2367 1033 2368
rect 1207 2368 1245 2369
rect 1207 2367 1210 2368
rect 1030 2337 1077 2367
rect 1163 2337 1210 2367
rect 1030 2336 1033 2337
rect 995 2335 1033 2336
rect 1207 2336 1210 2337
rect 1242 2367 1245 2368
rect 1443 2368 1481 2369
rect 1443 2367 1446 2368
rect 1242 2337 1290 2367
rect 1398 2337 1446 2367
rect 1242 2336 1245 2337
rect 1207 2335 1245 2336
rect 1443 2336 1446 2337
rect 1478 2367 1481 2368
rect 1655 2368 1693 2369
rect 1655 2367 1658 2368
rect 1478 2337 1525 2367
rect 1611 2337 1658 2367
rect 1478 2336 1481 2337
rect 1443 2335 1481 2336
rect 1655 2336 1658 2337
rect 1690 2367 1693 2368
rect 1891 2368 1929 2369
rect 1891 2367 1894 2368
rect 1690 2337 1738 2367
rect 1846 2337 1894 2367
rect 1690 2336 1693 2337
rect 1655 2335 1693 2336
rect 1891 2336 1894 2337
rect 1926 2367 1929 2368
rect 2103 2368 2141 2369
rect 2103 2367 2106 2368
rect 1926 2337 1973 2367
rect 2059 2337 2106 2367
rect 1926 2336 1929 2337
rect 1891 2335 1929 2336
rect 2103 2336 2106 2337
rect 2138 2367 2141 2368
rect 2339 2368 2377 2369
rect 2339 2367 2342 2368
rect 2138 2337 2186 2367
rect 2294 2337 2342 2367
rect 2138 2336 2141 2337
rect 2103 2335 2141 2336
rect 2339 2336 2342 2337
rect 2374 2367 2377 2368
rect 2551 2368 2589 2369
rect 2551 2367 2554 2368
rect 2374 2337 2421 2367
rect 2507 2337 2554 2367
rect 2374 2336 2377 2337
rect 2339 2335 2377 2336
rect 2551 2336 2554 2337
rect 2586 2367 2589 2368
rect 2787 2368 2825 2369
rect 2787 2367 2790 2368
rect 2586 2337 2634 2367
rect 2742 2337 2790 2367
rect 2586 2336 2589 2337
rect 2551 2335 2589 2336
rect 2787 2336 2790 2337
rect 2822 2367 2825 2368
rect 2999 2368 3037 2369
rect 2999 2367 3002 2368
rect 2822 2337 2869 2367
rect 2955 2337 3002 2367
rect 2822 2336 2825 2337
rect 2787 2335 2825 2336
rect 2999 2336 3002 2337
rect 3034 2367 3037 2368
rect 3235 2368 3273 2369
rect 3235 2367 3238 2368
rect 3034 2337 3082 2367
rect 3190 2337 3238 2367
rect 3034 2336 3037 2337
rect 2999 2335 3037 2336
rect 3235 2336 3238 2337
rect 3270 2367 3273 2368
rect 3447 2368 3485 2369
rect 3447 2367 3450 2368
rect 3270 2337 3317 2367
rect 3403 2337 3450 2367
rect 3270 2336 3273 2337
rect 3235 2335 3273 2336
rect 3447 2336 3450 2337
rect 3482 2367 3485 2368
rect 3683 2368 3721 2369
rect 3683 2367 3686 2368
rect 3482 2337 3530 2367
rect 3638 2337 3686 2367
rect 3482 2336 3485 2337
rect 3447 2335 3485 2336
rect 3683 2336 3686 2337
rect 3718 2367 3721 2368
rect 3895 2368 3933 2369
rect 3895 2367 3898 2368
rect 3718 2337 3765 2367
rect 3851 2337 3898 2367
rect 3718 2336 3721 2337
rect 3683 2335 3721 2336
rect 3895 2336 3898 2337
rect 3930 2367 3933 2368
rect 4131 2368 4169 2369
rect 4131 2367 4134 2368
rect 3930 2337 3978 2367
rect 4086 2337 4134 2367
rect 3930 2336 3933 2337
rect 3895 2335 3933 2336
rect 4131 2336 4134 2337
rect 4166 2367 4169 2368
rect 4343 2368 4381 2369
rect 4343 2367 4346 2368
rect 4166 2337 4213 2367
rect 4299 2337 4346 2367
rect 4166 2336 4169 2337
rect 4131 2335 4169 2336
rect 4343 2336 4346 2337
rect 4378 2367 4381 2368
rect 4579 2368 4617 2369
rect 4579 2367 4582 2368
rect 4378 2337 4426 2367
rect 4534 2337 4582 2367
rect 4378 2336 4381 2337
rect 4343 2335 4381 2336
rect 4579 2336 4582 2337
rect 4614 2367 4617 2368
rect 4791 2368 4829 2369
rect 4791 2367 4794 2368
rect 4614 2337 4661 2367
rect 4747 2337 4794 2367
rect 4614 2336 4617 2337
rect 4579 2335 4617 2336
rect 4791 2336 4794 2337
rect 4826 2367 4829 2368
rect 5027 2368 5065 2369
rect 5027 2367 5030 2368
rect 4826 2337 4874 2367
rect 4982 2337 5030 2367
rect 4826 2336 4829 2337
rect 4791 2335 4829 2336
rect 5027 2336 5030 2337
rect 5062 2367 5065 2368
rect 5239 2368 5277 2369
rect 5239 2367 5242 2368
rect 5062 2337 5109 2367
rect 5195 2337 5242 2367
rect 5062 2336 5065 2337
rect 5027 2335 5065 2336
rect 5239 2336 5242 2337
rect 5274 2367 5277 2368
rect 5475 2368 5513 2369
rect 5475 2367 5478 2368
rect 5274 2337 5322 2367
rect 5430 2337 5478 2367
rect 5274 2336 5277 2337
rect 5239 2335 5277 2336
rect 5475 2336 5478 2337
rect 5510 2367 5513 2368
rect 5687 2368 5725 2369
rect 5687 2367 5690 2368
rect 5510 2337 5557 2367
rect 5643 2337 5690 2367
rect 5510 2336 5513 2337
rect 5475 2335 5513 2336
rect 5687 2336 5690 2337
rect 5722 2367 5725 2368
rect 5923 2368 5961 2369
rect 5923 2367 5926 2368
rect 5722 2337 5770 2367
rect 5878 2337 5926 2367
rect 5722 2336 5725 2337
rect 5687 2335 5725 2336
rect 5923 2336 5926 2337
rect 5958 2367 5961 2368
rect 6135 2368 6173 2369
rect 6135 2367 6138 2368
rect 5958 2337 6005 2367
rect 6091 2337 6138 2367
rect 5958 2336 5961 2337
rect 5923 2335 5961 2336
rect 6135 2336 6138 2337
rect 6170 2367 6173 2368
rect 6371 2368 6409 2369
rect 6371 2367 6374 2368
rect 6170 2337 6218 2367
rect 6326 2337 6374 2367
rect 6170 2336 6173 2337
rect 6135 2335 6173 2336
rect 6371 2336 6374 2337
rect 6406 2367 6409 2368
rect 6583 2368 6621 2369
rect 6583 2367 6586 2368
rect 6406 2337 6453 2367
rect 6539 2337 6586 2367
rect 6406 2336 6409 2337
rect 6371 2335 6409 2336
rect 6583 2336 6586 2337
rect 6618 2367 6621 2368
rect 6819 2368 6857 2369
rect 6819 2367 6822 2368
rect 6618 2337 6666 2367
rect 6774 2337 6822 2367
rect 6618 2336 6621 2337
rect 6583 2335 6621 2336
rect 6819 2336 6822 2337
rect 6854 2367 6857 2368
rect 7031 2368 7069 2369
rect 7031 2367 7034 2368
rect 6854 2337 6901 2367
rect 6987 2337 7034 2367
rect 6854 2336 6857 2337
rect 6819 2335 6857 2336
rect 7031 2336 7034 2337
rect 7066 2367 7069 2368
rect 7267 2368 7305 2369
rect 7267 2367 7270 2368
rect 7066 2337 7114 2367
rect 7222 2337 7270 2367
rect 7066 2336 7069 2337
rect 7031 2335 7069 2336
rect 7267 2336 7270 2337
rect 7302 2367 7305 2368
rect 7479 2368 7517 2369
rect 7479 2367 7482 2368
rect 7302 2337 7349 2367
rect 7435 2337 7482 2367
rect 7302 2336 7305 2337
rect 7267 2335 7305 2336
rect 7479 2336 7482 2337
rect 7514 2367 7517 2368
rect 7715 2368 7753 2369
rect 7715 2367 7718 2368
rect 7514 2337 7562 2367
rect 7670 2337 7718 2367
rect 7514 2336 7517 2337
rect 7479 2335 7517 2336
rect 7715 2336 7718 2337
rect 7750 2367 7753 2368
rect 7927 2368 7965 2369
rect 7927 2367 7930 2368
rect 7750 2337 7797 2367
rect 7883 2337 7930 2367
rect 7750 2336 7753 2337
rect 7715 2335 7753 2336
rect 7927 2336 7930 2337
rect 7962 2367 7965 2368
rect 8163 2368 8201 2369
rect 8163 2367 8166 2368
rect 7962 2337 8010 2367
rect 8118 2337 8166 2367
rect 7962 2336 7965 2337
rect 7927 2335 7965 2336
rect 8163 2336 8166 2337
rect 8198 2367 8201 2368
rect 8375 2368 8413 2369
rect 8375 2367 8378 2368
rect 8198 2337 8245 2367
rect 8331 2337 8378 2367
rect 8198 2336 8201 2337
rect 8163 2335 8201 2336
rect 8375 2336 8378 2337
rect 8410 2367 8413 2368
rect 8611 2368 8649 2369
rect 8611 2367 8614 2368
rect 8410 2337 8458 2367
rect 8566 2337 8614 2367
rect 8410 2336 8413 2337
rect 8375 2335 8413 2336
rect 8611 2336 8614 2337
rect 8646 2367 8649 2368
rect 8823 2368 8861 2369
rect 8823 2367 8826 2368
rect 8646 2337 8693 2367
rect 8779 2337 8826 2367
rect 8646 2336 8649 2337
rect 8611 2335 8649 2336
rect 8823 2336 8826 2337
rect 8858 2367 8861 2368
rect 8858 2337 8906 2367
rect 8858 2336 8861 2337
rect 8823 2335 8861 2336
rect 196 2306 252 2309
rect 196 2305 201 2306
rect 35 2275 201 2305
rect 247 2305 252 2306
rect 644 2306 700 2309
rect 644 2305 649 2306
rect 247 2275 413 2305
rect 483 2275 649 2305
rect 695 2305 700 2306
rect 1092 2306 1148 2309
rect 1092 2305 1097 2306
rect 695 2275 861 2305
rect 931 2275 1097 2305
rect 1143 2305 1148 2306
rect 1540 2306 1596 2309
rect 1540 2305 1545 2306
rect 1143 2275 1309 2305
rect 1379 2275 1545 2305
rect 1591 2305 1596 2306
rect 1988 2306 2044 2309
rect 1988 2305 1993 2306
rect 1591 2275 1757 2305
rect 1827 2275 1993 2305
rect 2039 2305 2044 2306
rect 2436 2306 2492 2309
rect 2436 2305 2441 2306
rect 2039 2275 2205 2305
rect 2275 2275 2441 2305
rect 2487 2305 2492 2306
rect 2884 2306 2940 2309
rect 2884 2305 2889 2306
rect 2487 2275 2653 2305
rect 2723 2275 2889 2305
rect 2935 2305 2940 2306
rect 3332 2306 3388 2309
rect 3332 2305 3337 2306
rect 2935 2275 3101 2305
rect 3171 2275 3337 2305
rect 3383 2305 3388 2306
rect 3780 2306 3836 2309
rect 3780 2305 3785 2306
rect 3383 2275 3549 2305
rect 3619 2275 3785 2305
rect 3831 2305 3836 2306
rect 4228 2306 4284 2309
rect 4228 2305 4233 2306
rect 3831 2275 3997 2305
rect 4067 2275 4233 2305
rect 4279 2305 4284 2306
rect 4676 2306 4732 2309
rect 4676 2305 4681 2306
rect 4279 2275 4445 2305
rect 4515 2275 4681 2305
rect 4727 2305 4732 2306
rect 5124 2306 5180 2309
rect 5124 2305 5129 2306
rect 4727 2275 4893 2305
rect 4963 2275 5129 2305
rect 5175 2305 5180 2306
rect 5572 2306 5628 2309
rect 5572 2305 5577 2306
rect 5175 2275 5341 2305
rect 5411 2275 5577 2305
rect 5623 2305 5628 2306
rect 6020 2306 6076 2309
rect 6020 2305 6025 2306
rect 5623 2275 5789 2305
rect 5859 2275 6025 2305
rect 6071 2305 6076 2306
rect 6468 2306 6524 2309
rect 6468 2305 6473 2306
rect 6071 2275 6237 2305
rect 6307 2275 6473 2305
rect 6519 2305 6524 2306
rect 6916 2306 6972 2309
rect 6916 2305 6921 2306
rect 6519 2275 6685 2305
rect 6755 2275 6921 2305
rect 6967 2305 6972 2306
rect 7364 2306 7420 2309
rect 7364 2305 7369 2306
rect 6967 2275 7133 2305
rect 7203 2275 7369 2305
rect 7415 2305 7420 2306
rect 7812 2306 7868 2309
rect 7812 2305 7817 2306
rect 7415 2275 7581 2305
rect 7651 2275 7817 2305
rect 7863 2305 7868 2306
rect 8260 2306 8316 2309
rect 8260 2305 8265 2306
rect 7863 2275 8029 2305
rect 8099 2275 8265 2305
rect 8311 2305 8316 2306
rect 8708 2306 8764 2309
rect 8708 2305 8713 2306
rect 8311 2275 8477 2305
rect 8547 2275 8713 2305
rect 8759 2305 8764 2306
rect 8759 2275 8925 2305
rect 196 2271 252 2275
rect 644 2271 700 2275
rect 1092 2271 1148 2275
rect 1540 2271 1596 2275
rect 1988 2271 2044 2275
rect 2436 2271 2492 2275
rect 2884 2271 2940 2275
rect 3332 2271 3388 2275
rect 3780 2271 3836 2275
rect 4228 2271 4284 2275
rect 4676 2271 4732 2275
rect 5124 2271 5180 2275
rect 5572 2271 5628 2275
rect 6020 2271 6076 2275
rect 6468 2271 6524 2275
rect 6916 2271 6972 2275
rect 7364 2271 7420 2275
rect 7812 2271 7868 2275
rect 8260 2271 8316 2275
rect 8708 2271 8764 2275
rect 99 2244 137 2245
rect 99 2243 102 2244
rect 54 2213 102 2243
rect 99 2212 102 2213
rect 134 2243 137 2244
rect 311 2244 349 2245
rect 311 2243 314 2244
rect 134 2213 181 2243
rect 267 2213 314 2243
rect 134 2212 137 2213
rect 99 2211 137 2212
rect 311 2212 314 2213
rect 346 2243 349 2244
rect 547 2244 585 2245
rect 547 2243 550 2244
rect 346 2213 394 2243
rect 502 2213 550 2243
rect 346 2212 349 2213
rect 311 2211 349 2212
rect 547 2212 550 2213
rect 582 2243 585 2244
rect 759 2244 797 2245
rect 759 2243 762 2244
rect 582 2213 629 2243
rect 715 2213 762 2243
rect 582 2212 585 2213
rect 547 2211 585 2212
rect 759 2212 762 2213
rect 794 2243 797 2244
rect 995 2244 1033 2245
rect 995 2243 998 2244
rect 794 2213 842 2243
rect 950 2213 998 2243
rect 794 2212 797 2213
rect 759 2211 797 2212
rect 995 2212 998 2213
rect 1030 2243 1033 2244
rect 1207 2244 1245 2245
rect 1207 2243 1210 2244
rect 1030 2213 1077 2243
rect 1163 2213 1210 2243
rect 1030 2212 1033 2213
rect 995 2211 1033 2212
rect 1207 2212 1210 2213
rect 1242 2243 1245 2244
rect 1443 2244 1481 2245
rect 1443 2243 1446 2244
rect 1242 2213 1290 2243
rect 1398 2213 1446 2243
rect 1242 2212 1245 2213
rect 1207 2211 1245 2212
rect 1443 2212 1446 2213
rect 1478 2243 1481 2244
rect 1655 2244 1693 2245
rect 1655 2243 1658 2244
rect 1478 2213 1525 2243
rect 1611 2213 1658 2243
rect 1478 2212 1481 2213
rect 1443 2211 1481 2212
rect 1655 2212 1658 2213
rect 1690 2243 1693 2244
rect 1891 2244 1929 2245
rect 1891 2243 1894 2244
rect 1690 2213 1738 2243
rect 1846 2213 1894 2243
rect 1690 2212 1693 2213
rect 1655 2211 1693 2212
rect 1891 2212 1894 2213
rect 1926 2243 1929 2244
rect 2103 2244 2141 2245
rect 2103 2243 2106 2244
rect 1926 2213 1973 2243
rect 2059 2213 2106 2243
rect 1926 2212 1929 2213
rect 1891 2211 1929 2212
rect 2103 2212 2106 2213
rect 2138 2243 2141 2244
rect 2339 2244 2377 2245
rect 2339 2243 2342 2244
rect 2138 2213 2186 2243
rect 2294 2213 2342 2243
rect 2138 2212 2141 2213
rect 2103 2211 2141 2212
rect 2339 2212 2342 2213
rect 2374 2243 2377 2244
rect 2551 2244 2589 2245
rect 2551 2243 2554 2244
rect 2374 2213 2421 2243
rect 2507 2213 2554 2243
rect 2374 2212 2377 2213
rect 2339 2211 2377 2212
rect 2551 2212 2554 2213
rect 2586 2243 2589 2244
rect 2787 2244 2825 2245
rect 2787 2243 2790 2244
rect 2586 2213 2634 2243
rect 2742 2213 2790 2243
rect 2586 2212 2589 2213
rect 2551 2211 2589 2212
rect 2787 2212 2790 2213
rect 2822 2243 2825 2244
rect 2999 2244 3037 2245
rect 2999 2243 3002 2244
rect 2822 2213 2869 2243
rect 2955 2213 3002 2243
rect 2822 2212 2825 2213
rect 2787 2211 2825 2212
rect 2999 2212 3002 2213
rect 3034 2243 3037 2244
rect 3235 2244 3273 2245
rect 3235 2243 3238 2244
rect 3034 2213 3082 2243
rect 3190 2213 3238 2243
rect 3034 2212 3037 2213
rect 2999 2211 3037 2212
rect 3235 2212 3238 2213
rect 3270 2243 3273 2244
rect 3447 2244 3485 2245
rect 3447 2243 3450 2244
rect 3270 2213 3317 2243
rect 3403 2213 3450 2243
rect 3270 2212 3273 2213
rect 3235 2211 3273 2212
rect 3447 2212 3450 2213
rect 3482 2243 3485 2244
rect 3683 2244 3721 2245
rect 3683 2243 3686 2244
rect 3482 2213 3530 2243
rect 3638 2213 3686 2243
rect 3482 2212 3485 2213
rect 3447 2211 3485 2212
rect 3683 2212 3686 2213
rect 3718 2243 3721 2244
rect 3895 2244 3933 2245
rect 3895 2243 3898 2244
rect 3718 2213 3765 2243
rect 3851 2213 3898 2243
rect 3718 2212 3721 2213
rect 3683 2211 3721 2212
rect 3895 2212 3898 2213
rect 3930 2243 3933 2244
rect 4131 2244 4169 2245
rect 4131 2243 4134 2244
rect 3930 2213 3978 2243
rect 4086 2213 4134 2243
rect 3930 2212 3933 2213
rect 3895 2211 3933 2212
rect 4131 2212 4134 2213
rect 4166 2243 4169 2244
rect 4343 2244 4381 2245
rect 4343 2243 4346 2244
rect 4166 2213 4213 2243
rect 4299 2213 4346 2243
rect 4166 2212 4169 2213
rect 4131 2211 4169 2212
rect 4343 2212 4346 2213
rect 4378 2243 4381 2244
rect 4579 2244 4617 2245
rect 4579 2243 4582 2244
rect 4378 2213 4426 2243
rect 4534 2213 4582 2243
rect 4378 2212 4381 2213
rect 4343 2211 4381 2212
rect 4579 2212 4582 2213
rect 4614 2243 4617 2244
rect 4791 2244 4829 2245
rect 4791 2243 4794 2244
rect 4614 2213 4661 2243
rect 4747 2213 4794 2243
rect 4614 2212 4617 2213
rect 4579 2211 4617 2212
rect 4791 2212 4794 2213
rect 4826 2243 4829 2244
rect 5027 2244 5065 2245
rect 5027 2243 5030 2244
rect 4826 2213 4874 2243
rect 4982 2213 5030 2243
rect 4826 2212 4829 2213
rect 4791 2211 4829 2212
rect 5027 2212 5030 2213
rect 5062 2243 5065 2244
rect 5239 2244 5277 2245
rect 5239 2243 5242 2244
rect 5062 2213 5109 2243
rect 5195 2213 5242 2243
rect 5062 2212 5065 2213
rect 5027 2211 5065 2212
rect 5239 2212 5242 2213
rect 5274 2243 5277 2244
rect 5475 2244 5513 2245
rect 5475 2243 5478 2244
rect 5274 2213 5322 2243
rect 5430 2213 5478 2243
rect 5274 2212 5277 2213
rect 5239 2211 5277 2212
rect 5475 2212 5478 2213
rect 5510 2243 5513 2244
rect 5687 2244 5725 2245
rect 5687 2243 5690 2244
rect 5510 2213 5557 2243
rect 5643 2213 5690 2243
rect 5510 2212 5513 2213
rect 5475 2211 5513 2212
rect 5687 2212 5690 2213
rect 5722 2243 5725 2244
rect 5923 2244 5961 2245
rect 5923 2243 5926 2244
rect 5722 2213 5770 2243
rect 5878 2213 5926 2243
rect 5722 2212 5725 2213
rect 5687 2211 5725 2212
rect 5923 2212 5926 2213
rect 5958 2243 5961 2244
rect 6135 2244 6173 2245
rect 6135 2243 6138 2244
rect 5958 2213 6005 2243
rect 6091 2213 6138 2243
rect 5958 2212 5961 2213
rect 5923 2211 5961 2212
rect 6135 2212 6138 2213
rect 6170 2243 6173 2244
rect 6371 2244 6409 2245
rect 6371 2243 6374 2244
rect 6170 2213 6218 2243
rect 6326 2213 6374 2243
rect 6170 2212 6173 2213
rect 6135 2211 6173 2212
rect 6371 2212 6374 2213
rect 6406 2243 6409 2244
rect 6583 2244 6621 2245
rect 6583 2243 6586 2244
rect 6406 2213 6453 2243
rect 6539 2213 6586 2243
rect 6406 2212 6409 2213
rect 6371 2211 6409 2212
rect 6583 2212 6586 2213
rect 6618 2243 6621 2244
rect 6819 2244 6857 2245
rect 6819 2243 6822 2244
rect 6618 2213 6666 2243
rect 6774 2213 6822 2243
rect 6618 2212 6621 2213
rect 6583 2211 6621 2212
rect 6819 2212 6822 2213
rect 6854 2243 6857 2244
rect 7031 2244 7069 2245
rect 7031 2243 7034 2244
rect 6854 2213 6901 2243
rect 6987 2213 7034 2243
rect 6854 2212 6857 2213
rect 6819 2211 6857 2212
rect 7031 2212 7034 2213
rect 7066 2243 7069 2244
rect 7267 2244 7305 2245
rect 7267 2243 7270 2244
rect 7066 2213 7114 2243
rect 7222 2213 7270 2243
rect 7066 2212 7069 2213
rect 7031 2211 7069 2212
rect 7267 2212 7270 2213
rect 7302 2243 7305 2244
rect 7479 2244 7517 2245
rect 7479 2243 7482 2244
rect 7302 2213 7349 2243
rect 7435 2213 7482 2243
rect 7302 2212 7305 2213
rect 7267 2211 7305 2212
rect 7479 2212 7482 2213
rect 7514 2243 7517 2244
rect 7715 2244 7753 2245
rect 7715 2243 7718 2244
rect 7514 2213 7562 2243
rect 7670 2213 7718 2243
rect 7514 2212 7517 2213
rect 7479 2211 7517 2212
rect 7715 2212 7718 2213
rect 7750 2243 7753 2244
rect 7927 2244 7965 2245
rect 7927 2243 7930 2244
rect 7750 2213 7797 2243
rect 7883 2213 7930 2243
rect 7750 2212 7753 2213
rect 7715 2211 7753 2212
rect 7927 2212 7930 2213
rect 7962 2243 7965 2244
rect 8163 2244 8201 2245
rect 8163 2243 8166 2244
rect 7962 2213 8010 2243
rect 8118 2213 8166 2243
rect 7962 2212 7965 2213
rect 7927 2211 7965 2212
rect 8163 2212 8166 2213
rect 8198 2243 8201 2244
rect 8375 2244 8413 2245
rect 8375 2243 8378 2244
rect 8198 2213 8245 2243
rect 8331 2213 8378 2243
rect 8198 2212 8201 2213
rect 8163 2211 8201 2212
rect 8375 2212 8378 2213
rect 8410 2243 8413 2244
rect 8611 2244 8649 2245
rect 8611 2243 8614 2244
rect 8410 2213 8458 2243
rect 8566 2213 8614 2243
rect 8410 2212 8413 2213
rect 8375 2211 8413 2212
rect 8611 2212 8614 2213
rect 8646 2243 8649 2244
rect 8823 2244 8861 2245
rect 8823 2243 8826 2244
rect 8646 2213 8693 2243
rect 8779 2213 8826 2243
rect 8646 2212 8649 2213
rect 8611 2211 8649 2212
rect 8823 2212 8826 2213
rect 8858 2243 8861 2244
rect 8858 2213 8906 2243
rect 8858 2212 8861 2213
rect 8823 2211 8861 2212
rect 196 2182 252 2185
rect 196 2181 201 2182
rect 35 2151 201 2181
rect 247 2181 252 2182
rect 644 2182 700 2185
rect 644 2181 649 2182
rect 247 2151 413 2181
rect 483 2151 649 2181
rect 695 2181 700 2182
rect 1092 2182 1148 2185
rect 1092 2181 1097 2182
rect 695 2151 861 2181
rect 931 2151 1097 2181
rect 1143 2181 1148 2182
rect 1540 2182 1596 2185
rect 1540 2181 1545 2182
rect 1143 2151 1309 2181
rect 1379 2151 1545 2181
rect 1591 2181 1596 2182
rect 1988 2182 2044 2185
rect 1988 2181 1993 2182
rect 1591 2151 1757 2181
rect 1827 2151 1993 2181
rect 2039 2181 2044 2182
rect 2436 2182 2492 2185
rect 2436 2181 2441 2182
rect 2039 2151 2205 2181
rect 2275 2151 2441 2181
rect 2487 2181 2492 2182
rect 2884 2182 2940 2185
rect 2884 2181 2889 2182
rect 2487 2151 2653 2181
rect 2723 2151 2889 2181
rect 2935 2181 2940 2182
rect 3332 2182 3388 2185
rect 3332 2181 3337 2182
rect 2935 2151 3101 2181
rect 3171 2151 3337 2181
rect 3383 2181 3388 2182
rect 3780 2182 3836 2185
rect 3780 2181 3785 2182
rect 3383 2151 3549 2181
rect 3619 2151 3785 2181
rect 3831 2181 3836 2182
rect 4228 2182 4284 2185
rect 4228 2181 4233 2182
rect 3831 2151 3997 2181
rect 4067 2151 4233 2181
rect 4279 2181 4284 2182
rect 4676 2182 4732 2185
rect 4676 2181 4681 2182
rect 4279 2151 4445 2181
rect 4515 2151 4681 2181
rect 4727 2181 4732 2182
rect 5124 2182 5180 2185
rect 5124 2181 5129 2182
rect 4727 2151 4893 2181
rect 4963 2151 5129 2181
rect 5175 2181 5180 2182
rect 5572 2182 5628 2185
rect 5572 2181 5577 2182
rect 5175 2151 5341 2181
rect 5411 2151 5577 2181
rect 5623 2181 5628 2182
rect 6020 2182 6076 2185
rect 6020 2181 6025 2182
rect 5623 2151 5789 2181
rect 5859 2151 6025 2181
rect 6071 2181 6076 2182
rect 6468 2182 6524 2185
rect 6468 2181 6473 2182
rect 6071 2151 6237 2181
rect 6307 2151 6473 2181
rect 6519 2181 6524 2182
rect 6916 2182 6972 2185
rect 6916 2181 6921 2182
rect 6519 2151 6685 2181
rect 6755 2151 6921 2181
rect 6967 2181 6972 2182
rect 7364 2182 7420 2185
rect 7364 2181 7369 2182
rect 6967 2151 7133 2181
rect 7203 2151 7369 2181
rect 7415 2181 7420 2182
rect 7812 2182 7868 2185
rect 7812 2181 7817 2182
rect 7415 2151 7581 2181
rect 7651 2151 7817 2181
rect 7863 2181 7868 2182
rect 8260 2182 8316 2185
rect 8260 2181 8265 2182
rect 7863 2151 8029 2181
rect 8099 2151 8265 2181
rect 8311 2181 8316 2182
rect 8708 2182 8764 2185
rect 8708 2181 8713 2182
rect 8311 2151 8477 2181
rect 8547 2151 8713 2181
rect 8759 2181 8764 2182
rect 8759 2151 8925 2181
rect 196 2147 252 2151
rect 644 2147 700 2151
rect 1092 2147 1148 2151
rect 1540 2147 1596 2151
rect 1988 2147 2044 2151
rect 2436 2147 2492 2151
rect 2884 2147 2940 2151
rect 3332 2147 3388 2151
rect 3780 2147 3836 2151
rect 4228 2147 4284 2151
rect 4676 2147 4732 2151
rect 5124 2147 5180 2151
rect 5572 2147 5628 2151
rect 6020 2147 6076 2151
rect 6468 2147 6524 2151
rect 6916 2147 6972 2151
rect 7364 2147 7420 2151
rect 7812 2147 7868 2151
rect 8260 2147 8316 2151
rect 8708 2147 8764 2151
rect 99 2120 137 2121
rect 99 2119 102 2120
rect 54 2089 102 2119
rect 99 2088 102 2089
rect 134 2119 137 2120
rect 311 2120 349 2121
rect 311 2119 314 2120
rect 134 2089 181 2119
rect 267 2089 314 2119
rect 134 2088 137 2089
rect 99 2087 137 2088
rect 311 2088 314 2089
rect 346 2119 349 2120
rect 547 2120 585 2121
rect 547 2119 550 2120
rect 346 2089 394 2119
rect 502 2089 550 2119
rect 346 2088 349 2089
rect 311 2087 349 2088
rect 547 2088 550 2089
rect 582 2119 585 2120
rect 759 2120 797 2121
rect 759 2119 762 2120
rect 582 2089 629 2119
rect 715 2089 762 2119
rect 582 2088 585 2089
rect 547 2087 585 2088
rect 759 2088 762 2089
rect 794 2119 797 2120
rect 995 2120 1033 2121
rect 995 2119 998 2120
rect 794 2089 842 2119
rect 950 2089 998 2119
rect 794 2088 797 2089
rect 759 2087 797 2088
rect 995 2088 998 2089
rect 1030 2119 1033 2120
rect 1207 2120 1245 2121
rect 1207 2119 1210 2120
rect 1030 2089 1077 2119
rect 1163 2089 1210 2119
rect 1030 2088 1033 2089
rect 995 2087 1033 2088
rect 1207 2088 1210 2089
rect 1242 2119 1245 2120
rect 1443 2120 1481 2121
rect 1443 2119 1446 2120
rect 1242 2089 1290 2119
rect 1398 2089 1446 2119
rect 1242 2088 1245 2089
rect 1207 2087 1245 2088
rect 1443 2088 1446 2089
rect 1478 2119 1481 2120
rect 1655 2120 1693 2121
rect 1655 2119 1658 2120
rect 1478 2089 1525 2119
rect 1611 2089 1658 2119
rect 1478 2088 1481 2089
rect 1443 2087 1481 2088
rect 1655 2088 1658 2089
rect 1690 2119 1693 2120
rect 1891 2120 1929 2121
rect 1891 2119 1894 2120
rect 1690 2089 1738 2119
rect 1846 2089 1894 2119
rect 1690 2088 1693 2089
rect 1655 2087 1693 2088
rect 1891 2088 1894 2089
rect 1926 2119 1929 2120
rect 2103 2120 2141 2121
rect 2103 2119 2106 2120
rect 1926 2089 1973 2119
rect 2059 2089 2106 2119
rect 1926 2088 1929 2089
rect 1891 2087 1929 2088
rect 2103 2088 2106 2089
rect 2138 2119 2141 2120
rect 2339 2120 2377 2121
rect 2339 2119 2342 2120
rect 2138 2089 2186 2119
rect 2294 2089 2342 2119
rect 2138 2088 2141 2089
rect 2103 2087 2141 2088
rect 2339 2088 2342 2089
rect 2374 2119 2377 2120
rect 2551 2120 2589 2121
rect 2551 2119 2554 2120
rect 2374 2089 2421 2119
rect 2507 2089 2554 2119
rect 2374 2088 2377 2089
rect 2339 2087 2377 2088
rect 2551 2088 2554 2089
rect 2586 2119 2589 2120
rect 2787 2120 2825 2121
rect 2787 2119 2790 2120
rect 2586 2089 2634 2119
rect 2742 2089 2790 2119
rect 2586 2088 2589 2089
rect 2551 2087 2589 2088
rect 2787 2088 2790 2089
rect 2822 2119 2825 2120
rect 2999 2120 3037 2121
rect 2999 2119 3002 2120
rect 2822 2089 2869 2119
rect 2955 2089 3002 2119
rect 2822 2088 2825 2089
rect 2787 2087 2825 2088
rect 2999 2088 3002 2089
rect 3034 2119 3037 2120
rect 3235 2120 3273 2121
rect 3235 2119 3238 2120
rect 3034 2089 3082 2119
rect 3190 2089 3238 2119
rect 3034 2088 3037 2089
rect 2999 2087 3037 2088
rect 3235 2088 3238 2089
rect 3270 2119 3273 2120
rect 3447 2120 3485 2121
rect 3447 2119 3450 2120
rect 3270 2089 3317 2119
rect 3403 2089 3450 2119
rect 3270 2088 3273 2089
rect 3235 2087 3273 2088
rect 3447 2088 3450 2089
rect 3482 2119 3485 2120
rect 3683 2120 3721 2121
rect 3683 2119 3686 2120
rect 3482 2089 3530 2119
rect 3638 2089 3686 2119
rect 3482 2088 3485 2089
rect 3447 2087 3485 2088
rect 3683 2088 3686 2089
rect 3718 2119 3721 2120
rect 3895 2120 3933 2121
rect 3895 2119 3898 2120
rect 3718 2089 3765 2119
rect 3851 2089 3898 2119
rect 3718 2088 3721 2089
rect 3683 2087 3721 2088
rect 3895 2088 3898 2089
rect 3930 2119 3933 2120
rect 4131 2120 4169 2121
rect 4131 2119 4134 2120
rect 3930 2089 3978 2119
rect 4086 2089 4134 2119
rect 3930 2088 3933 2089
rect 3895 2087 3933 2088
rect 4131 2088 4134 2089
rect 4166 2119 4169 2120
rect 4343 2120 4381 2121
rect 4343 2119 4346 2120
rect 4166 2089 4213 2119
rect 4299 2089 4346 2119
rect 4166 2088 4169 2089
rect 4131 2087 4169 2088
rect 4343 2088 4346 2089
rect 4378 2119 4381 2120
rect 4579 2120 4617 2121
rect 4579 2119 4582 2120
rect 4378 2089 4426 2119
rect 4534 2089 4582 2119
rect 4378 2088 4381 2089
rect 4343 2087 4381 2088
rect 4579 2088 4582 2089
rect 4614 2119 4617 2120
rect 4791 2120 4829 2121
rect 4791 2119 4794 2120
rect 4614 2089 4661 2119
rect 4747 2089 4794 2119
rect 4614 2088 4617 2089
rect 4579 2087 4617 2088
rect 4791 2088 4794 2089
rect 4826 2119 4829 2120
rect 5027 2120 5065 2121
rect 5027 2119 5030 2120
rect 4826 2089 4874 2119
rect 4982 2089 5030 2119
rect 4826 2088 4829 2089
rect 4791 2087 4829 2088
rect 5027 2088 5030 2089
rect 5062 2119 5065 2120
rect 5239 2120 5277 2121
rect 5239 2119 5242 2120
rect 5062 2089 5109 2119
rect 5195 2089 5242 2119
rect 5062 2088 5065 2089
rect 5027 2087 5065 2088
rect 5239 2088 5242 2089
rect 5274 2119 5277 2120
rect 5475 2120 5513 2121
rect 5475 2119 5478 2120
rect 5274 2089 5322 2119
rect 5430 2089 5478 2119
rect 5274 2088 5277 2089
rect 5239 2087 5277 2088
rect 5475 2088 5478 2089
rect 5510 2119 5513 2120
rect 5687 2120 5725 2121
rect 5687 2119 5690 2120
rect 5510 2089 5557 2119
rect 5643 2089 5690 2119
rect 5510 2088 5513 2089
rect 5475 2087 5513 2088
rect 5687 2088 5690 2089
rect 5722 2119 5725 2120
rect 5923 2120 5961 2121
rect 5923 2119 5926 2120
rect 5722 2089 5770 2119
rect 5878 2089 5926 2119
rect 5722 2088 5725 2089
rect 5687 2087 5725 2088
rect 5923 2088 5926 2089
rect 5958 2119 5961 2120
rect 6135 2120 6173 2121
rect 6135 2119 6138 2120
rect 5958 2089 6005 2119
rect 6091 2089 6138 2119
rect 5958 2088 5961 2089
rect 5923 2087 5961 2088
rect 6135 2088 6138 2089
rect 6170 2119 6173 2120
rect 6371 2120 6409 2121
rect 6371 2119 6374 2120
rect 6170 2089 6218 2119
rect 6326 2089 6374 2119
rect 6170 2088 6173 2089
rect 6135 2087 6173 2088
rect 6371 2088 6374 2089
rect 6406 2119 6409 2120
rect 6583 2120 6621 2121
rect 6583 2119 6586 2120
rect 6406 2089 6453 2119
rect 6539 2089 6586 2119
rect 6406 2088 6409 2089
rect 6371 2087 6409 2088
rect 6583 2088 6586 2089
rect 6618 2119 6621 2120
rect 6819 2120 6857 2121
rect 6819 2119 6822 2120
rect 6618 2089 6666 2119
rect 6774 2089 6822 2119
rect 6618 2088 6621 2089
rect 6583 2087 6621 2088
rect 6819 2088 6822 2089
rect 6854 2119 6857 2120
rect 7031 2120 7069 2121
rect 7031 2119 7034 2120
rect 6854 2089 6901 2119
rect 6987 2089 7034 2119
rect 6854 2088 6857 2089
rect 6819 2087 6857 2088
rect 7031 2088 7034 2089
rect 7066 2119 7069 2120
rect 7267 2120 7305 2121
rect 7267 2119 7270 2120
rect 7066 2089 7114 2119
rect 7222 2089 7270 2119
rect 7066 2088 7069 2089
rect 7031 2087 7069 2088
rect 7267 2088 7270 2089
rect 7302 2119 7305 2120
rect 7479 2120 7517 2121
rect 7479 2119 7482 2120
rect 7302 2089 7349 2119
rect 7435 2089 7482 2119
rect 7302 2088 7305 2089
rect 7267 2087 7305 2088
rect 7479 2088 7482 2089
rect 7514 2119 7517 2120
rect 7715 2120 7753 2121
rect 7715 2119 7718 2120
rect 7514 2089 7562 2119
rect 7670 2089 7718 2119
rect 7514 2088 7517 2089
rect 7479 2087 7517 2088
rect 7715 2088 7718 2089
rect 7750 2119 7753 2120
rect 7927 2120 7965 2121
rect 7927 2119 7930 2120
rect 7750 2089 7797 2119
rect 7883 2089 7930 2119
rect 7750 2088 7753 2089
rect 7715 2087 7753 2088
rect 7927 2088 7930 2089
rect 7962 2119 7965 2120
rect 8163 2120 8201 2121
rect 8163 2119 8166 2120
rect 7962 2089 8010 2119
rect 8118 2089 8166 2119
rect 7962 2088 7965 2089
rect 7927 2087 7965 2088
rect 8163 2088 8166 2089
rect 8198 2119 8201 2120
rect 8375 2120 8413 2121
rect 8375 2119 8378 2120
rect 8198 2089 8245 2119
rect 8331 2089 8378 2119
rect 8198 2088 8201 2089
rect 8163 2087 8201 2088
rect 8375 2088 8378 2089
rect 8410 2119 8413 2120
rect 8611 2120 8649 2121
rect 8611 2119 8614 2120
rect 8410 2089 8458 2119
rect 8566 2089 8614 2119
rect 8410 2088 8413 2089
rect 8375 2087 8413 2088
rect 8611 2088 8614 2089
rect 8646 2119 8649 2120
rect 8823 2120 8861 2121
rect 8823 2119 8826 2120
rect 8646 2089 8693 2119
rect 8779 2089 8826 2119
rect 8646 2088 8649 2089
rect 8611 2087 8649 2088
rect 8823 2088 8826 2089
rect 8858 2119 8861 2120
rect 8858 2089 8906 2119
rect 8858 2088 8861 2089
rect 8823 2087 8861 2088
rect 196 2058 252 2061
rect 196 2057 201 2058
rect 35 2027 201 2057
rect 247 2057 252 2058
rect 644 2058 700 2061
rect 644 2057 649 2058
rect 247 2027 413 2057
rect 483 2027 649 2057
rect 695 2057 700 2058
rect 1092 2058 1148 2061
rect 1092 2057 1097 2058
rect 695 2027 861 2057
rect 931 2027 1097 2057
rect 1143 2057 1148 2058
rect 1540 2058 1596 2061
rect 1540 2057 1545 2058
rect 1143 2027 1309 2057
rect 1379 2027 1545 2057
rect 1591 2057 1596 2058
rect 1988 2058 2044 2061
rect 1988 2057 1993 2058
rect 1591 2027 1757 2057
rect 1827 2027 1993 2057
rect 2039 2057 2044 2058
rect 2436 2058 2492 2061
rect 2436 2057 2441 2058
rect 2039 2027 2205 2057
rect 2275 2027 2441 2057
rect 2487 2057 2492 2058
rect 2884 2058 2940 2061
rect 2884 2057 2889 2058
rect 2487 2027 2653 2057
rect 2723 2027 2889 2057
rect 2935 2057 2940 2058
rect 3332 2058 3388 2061
rect 3332 2057 3337 2058
rect 2935 2027 3101 2057
rect 3171 2027 3337 2057
rect 3383 2057 3388 2058
rect 3780 2058 3836 2061
rect 3780 2057 3785 2058
rect 3383 2027 3549 2057
rect 3619 2027 3785 2057
rect 3831 2057 3836 2058
rect 4228 2058 4284 2061
rect 4228 2057 4233 2058
rect 3831 2027 3997 2057
rect 4067 2027 4233 2057
rect 4279 2057 4284 2058
rect 4676 2058 4732 2061
rect 4676 2057 4681 2058
rect 4279 2027 4445 2057
rect 4515 2027 4681 2057
rect 4727 2057 4732 2058
rect 5124 2058 5180 2061
rect 5124 2057 5129 2058
rect 4727 2027 4893 2057
rect 4963 2027 5129 2057
rect 5175 2057 5180 2058
rect 5572 2058 5628 2061
rect 5572 2057 5577 2058
rect 5175 2027 5341 2057
rect 5411 2027 5577 2057
rect 5623 2057 5628 2058
rect 6020 2058 6076 2061
rect 6020 2057 6025 2058
rect 5623 2027 5789 2057
rect 5859 2027 6025 2057
rect 6071 2057 6076 2058
rect 6468 2058 6524 2061
rect 6468 2057 6473 2058
rect 6071 2027 6237 2057
rect 6307 2027 6473 2057
rect 6519 2057 6524 2058
rect 6916 2058 6972 2061
rect 6916 2057 6921 2058
rect 6519 2027 6685 2057
rect 6755 2027 6921 2057
rect 6967 2057 6972 2058
rect 7364 2058 7420 2061
rect 7364 2057 7369 2058
rect 6967 2027 7133 2057
rect 7203 2027 7369 2057
rect 7415 2057 7420 2058
rect 7812 2058 7868 2061
rect 7812 2057 7817 2058
rect 7415 2027 7581 2057
rect 7651 2027 7817 2057
rect 7863 2057 7868 2058
rect 8260 2058 8316 2061
rect 8260 2057 8265 2058
rect 7863 2027 8029 2057
rect 8099 2027 8265 2057
rect 8311 2057 8316 2058
rect 8708 2058 8764 2061
rect 8708 2057 8713 2058
rect 8311 2027 8477 2057
rect 8547 2027 8713 2057
rect 8759 2057 8764 2058
rect 8759 2027 8925 2057
rect 196 2023 252 2027
rect 644 2023 700 2027
rect 1092 2023 1148 2027
rect 1540 2023 1596 2027
rect 1988 2023 2044 2027
rect 2436 2023 2492 2027
rect 2884 2023 2940 2027
rect 3332 2023 3388 2027
rect 3780 2023 3836 2027
rect 4228 2023 4284 2027
rect 4676 2023 4732 2027
rect 5124 2023 5180 2027
rect 5572 2023 5628 2027
rect 6020 2023 6076 2027
rect 6468 2023 6524 2027
rect 6916 2023 6972 2027
rect 7364 2023 7420 2027
rect 7812 2023 7868 2027
rect 8260 2023 8316 2027
rect 8708 2023 8764 2027
rect 99 1996 137 1997
rect 99 1995 102 1996
rect 54 1965 102 1995
rect 99 1964 102 1965
rect 134 1995 137 1996
rect 311 1996 349 1997
rect 311 1995 314 1996
rect 134 1965 181 1995
rect 267 1965 314 1995
rect 134 1964 137 1965
rect 99 1963 137 1964
rect 311 1964 314 1965
rect 346 1995 349 1996
rect 547 1996 585 1997
rect 547 1995 550 1996
rect 346 1965 394 1995
rect 502 1965 550 1995
rect 346 1964 349 1965
rect 311 1963 349 1964
rect 547 1964 550 1965
rect 582 1995 585 1996
rect 759 1996 797 1997
rect 759 1995 762 1996
rect 582 1965 629 1995
rect 715 1965 762 1995
rect 582 1964 585 1965
rect 547 1963 585 1964
rect 759 1964 762 1965
rect 794 1995 797 1996
rect 995 1996 1033 1997
rect 995 1995 998 1996
rect 794 1965 842 1995
rect 950 1965 998 1995
rect 794 1964 797 1965
rect 759 1963 797 1964
rect 995 1964 998 1965
rect 1030 1995 1033 1996
rect 1207 1996 1245 1997
rect 1207 1995 1210 1996
rect 1030 1965 1077 1995
rect 1163 1965 1210 1995
rect 1030 1964 1033 1965
rect 995 1963 1033 1964
rect 1207 1964 1210 1965
rect 1242 1995 1245 1996
rect 1443 1996 1481 1997
rect 1443 1995 1446 1996
rect 1242 1965 1290 1995
rect 1398 1965 1446 1995
rect 1242 1964 1245 1965
rect 1207 1963 1245 1964
rect 1443 1964 1446 1965
rect 1478 1995 1481 1996
rect 1655 1996 1693 1997
rect 1655 1995 1658 1996
rect 1478 1965 1525 1995
rect 1611 1965 1658 1995
rect 1478 1964 1481 1965
rect 1443 1963 1481 1964
rect 1655 1964 1658 1965
rect 1690 1995 1693 1996
rect 1891 1996 1929 1997
rect 1891 1995 1894 1996
rect 1690 1965 1738 1995
rect 1846 1965 1894 1995
rect 1690 1964 1693 1965
rect 1655 1963 1693 1964
rect 1891 1964 1894 1965
rect 1926 1995 1929 1996
rect 2103 1996 2141 1997
rect 2103 1995 2106 1996
rect 1926 1965 1973 1995
rect 2059 1965 2106 1995
rect 1926 1964 1929 1965
rect 1891 1963 1929 1964
rect 2103 1964 2106 1965
rect 2138 1995 2141 1996
rect 2339 1996 2377 1997
rect 2339 1995 2342 1996
rect 2138 1965 2186 1995
rect 2294 1965 2342 1995
rect 2138 1964 2141 1965
rect 2103 1963 2141 1964
rect 2339 1964 2342 1965
rect 2374 1995 2377 1996
rect 2551 1996 2589 1997
rect 2551 1995 2554 1996
rect 2374 1965 2421 1995
rect 2507 1965 2554 1995
rect 2374 1964 2377 1965
rect 2339 1963 2377 1964
rect 2551 1964 2554 1965
rect 2586 1995 2589 1996
rect 2787 1996 2825 1997
rect 2787 1995 2790 1996
rect 2586 1965 2634 1995
rect 2742 1965 2790 1995
rect 2586 1964 2589 1965
rect 2551 1963 2589 1964
rect 2787 1964 2790 1965
rect 2822 1995 2825 1996
rect 2999 1996 3037 1997
rect 2999 1995 3002 1996
rect 2822 1965 2869 1995
rect 2955 1965 3002 1995
rect 2822 1964 2825 1965
rect 2787 1963 2825 1964
rect 2999 1964 3002 1965
rect 3034 1995 3037 1996
rect 3235 1996 3273 1997
rect 3235 1995 3238 1996
rect 3034 1965 3082 1995
rect 3190 1965 3238 1995
rect 3034 1964 3037 1965
rect 2999 1963 3037 1964
rect 3235 1964 3238 1965
rect 3270 1995 3273 1996
rect 3447 1996 3485 1997
rect 3447 1995 3450 1996
rect 3270 1965 3317 1995
rect 3403 1965 3450 1995
rect 3270 1964 3273 1965
rect 3235 1963 3273 1964
rect 3447 1964 3450 1965
rect 3482 1995 3485 1996
rect 3683 1996 3721 1997
rect 3683 1995 3686 1996
rect 3482 1965 3530 1995
rect 3638 1965 3686 1995
rect 3482 1964 3485 1965
rect 3447 1963 3485 1964
rect 3683 1964 3686 1965
rect 3718 1995 3721 1996
rect 3895 1996 3933 1997
rect 3895 1995 3898 1996
rect 3718 1965 3765 1995
rect 3851 1965 3898 1995
rect 3718 1964 3721 1965
rect 3683 1963 3721 1964
rect 3895 1964 3898 1965
rect 3930 1995 3933 1996
rect 4131 1996 4169 1997
rect 4131 1995 4134 1996
rect 3930 1965 3978 1995
rect 4086 1965 4134 1995
rect 3930 1964 3933 1965
rect 3895 1963 3933 1964
rect 4131 1964 4134 1965
rect 4166 1995 4169 1996
rect 4343 1996 4381 1997
rect 4343 1995 4346 1996
rect 4166 1965 4213 1995
rect 4299 1965 4346 1995
rect 4166 1964 4169 1965
rect 4131 1963 4169 1964
rect 4343 1964 4346 1965
rect 4378 1995 4381 1996
rect 4579 1996 4617 1997
rect 4579 1995 4582 1996
rect 4378 1965 4426 1995
rect 4534 1965 4582 1995
rect 4378 1964 4381 1965
rect 4343 1963 4381 1964
rect 4579 1964 4582 1965
rect 4614 1995 4617 1996
rect 4791 1996 4829 1997
rect 4791 1995 4794 1996
rect 4614 1965 4661 1995
rect 4747 1965 4794 1995
rect 4614 1964 4617 1965
rect 4579 1963 4617 1964
rect 4791 1964 4794 1965
rect 4826 1995 4829 1996
rect 5027 1996 5065 1997
rect 5027 1995 5030 1996
rect 4826 1965 4874 1995
rect 4982 1965 5030 1995
rect 4826 1964 4829 1965
rect 4791 1963 4829 1964
rect 5027 1964 5030 1965
rect 5062 1995 5065 1996
rect 5239 1996 5277 1997
rect 5239 1995 5242 1996
rect 5062 1965 5109 1995
rect 5195 1965 5242 1995
rect 5062 1964 5065 1965
rect 5027 1963 5065 1964
rect 5239 1964 5242 1965
rect 5274 1995 5277 1996
rect 5475 1996 5513 1997
rect 5475 1995 5478 1996
rect 5274 1965 5322 1995
rect 5430 1965 5478 1995
rect 5274 1964 5277 1965
rect 5239 1963 5277 1964
rect 5475 1964 5478 1965
rect 5510 1995 5513 1996
rect 5687 1996 5725 1997
rect 5687 1995 5690 1996
rect 5510 1965 5557 1995
rect 5643 1965 5690 1995
rect 5510 1964 5513 1965
rect 5475 1963 5513 1964
rect 5687 1964 5690 1965
rect 5722 1995 5725 1996
rect 5923 1996 5961 1997
rect 5923 1995 5926 1996
rect 5722 1965 5770 1995
rect 5878 1965 5926 1995
rect 5722 1964 5725 1965
rect 5687 1963 5725 1964
rect 5923 1964 5926 1965
rect 5958 1995 5961 1996
rect 6135 1996 6173 1997
rect 6135 1995 6138 1996
rect 5958 1965 6005 1995
rect 6091 1965 6138 1995
rect 5958 1964 5961 1965
rect 5923 1963 5961 1964
rect 6135 1964 6138 1965
rect 6170 1995 6173 1996
rect 6371 1996 6409 1997
rect 6371 1995 6374 1996
rect 6170 1965 6218 1995
rect 6326 1965 6374 1995
rect 6170 1964 6173 1965
rect 6135 1963 6173 1964
rect 6371 1964 6374 1965
rect 6406 1995 6409 1996
rect 6583 1996 6621 1997
rect 6583 1995 6586 1996
rect 6406 1965 6453 1995
rect 6539 1965 6586 1995
rect 6406 1964 6409 1965
rect 6371 1963 6409 1964
rect 6583 1964 6586 1965
rect 6618 1995 6621 1996
rect 6819 1996 6857 1997
rect 6819 1995 6822 1996
rect 6618 1965 6666 1995
rect 6774 1965 6822 1995
rect 6618 1964 6621 1965
rect 6583 1963 6621 1964
rect 6819 1964 6822 1965
rect 6854 1995 6857 1996
rect 7031 1996 7069 1997
rect 7031 1995 7034 1996
rect 6854 1965 6901 1995
rect 6987 1965 7034 1995
rect 6854 1964 6857 1965
rect 6819 1963 6857 1964
rect 7031 1964 7034 1965
rect 7066 1995 7069 1996
rect 7267 1996 7305 1997
rect 7267 1995 7270 1996
rect 7066 1965 7114 1995
rect 7222 1965 7270 1995
rect 7066 1964 7069 1965
rect 7031 1963 7069 1964
rect 7267 1964 7270 1965
rect 7302 1995 7305 1996
rect 7479 1996 7517 1997
rect 7479 1995 7482 1996
rect 7302 1965 7349 1995
rect 7435 1965 7482 1995
rect 7302 1964 7305 1965
rect 7267 1963 7305 1964
rect 7479 1964 7482 1965
rect 7514 1995 7517 1996
rect 7715 1996 7753 1997
rect 7715 1995 7718 1996
rect 7514 1965 7562 1995
rect 7670 1965 7718 1995
rect 7514 1964 7517 1965
rect 7479 1963 7517 1964
rect 7715 1964 7718 1965
rect 7750 1995 7753 1996
rect 7927 1996 7965 1997
rect 7927 1995 7930 1996
rect 7750 1965 7797 1995
rect 7883 1965 7930 1995
rect 7750 1964 7753 1965
rect 7715 1963 7753 1964
rect 7927 1964 7930 1965
rect 7962 1995 7965 1996
rect 8163 1996 8201 1997
rect 8163 1995 8166 1996
rect 7962 1965 8010 1995
rect 8118 1965 8166 1995
rect 7962 1964 7965 1965
rect 7927 1963 7965 1964
rect 8163 1964 8166 1965
rect 8198 1995 8201 1996
rect 8375 1996 8413 1997
rect 8375 1995 8378 1996
rect 8198 1965 8245 1995
rect 8331 1965 8378 1995
rect 8198 1964 8201 1965
rect 8163 1963 8201 1964
rect 8375 1964 8378 1965
rect 8410 1995 8413 1996
rect 8611 1996 8649 1997
rect 8611 1995 8614 1996
rect 8410 1965 8458 1995
rect 8566 1965 8614 1995
rect 8410 1964 8413 1965
rect 8375 1963 8413 1964
rect 8611 1964 8614 1965
rect 8646 1995 8649 1996
rect 8823 1996 8861 1997
rect 8823 1995 8826 1996
rect 8646 1965 8693 1995
rect 8779 1965 8826 1995
rect 8646 1964 8649 1965
rect 8611 1963 8649 1964
rect 8823 1964 8826 1965
rect 8858 1995 8861 1996
rect 8858 1965 8906 1995
rect 8858 1964 8861 1965
rect 8823 1963 8861 1964
rect 196 1934 252 1937
rect 196 1933 201 1934
rect 35 1903 201 1933
rect 247 1933 252 1934
rect 644 1934 700 1937
rect 644 1933 649 1934
rect 247 1903 413 1933
rect 483 1903 649 1933
rect 695 1933 700 1934
rect 1092 1934 1148 1937
rect 1092 1933 1097 1934
rect 695 1903 861 1933
rect 931 1903 1097 1933
rect 1143 1933 1148 1934
rect 1540 1934 1596 1937
rect 1540 1933 1545 1934
rect 1143 1903 1309 1933
rect 1379 1903 1545 1933
rect 1591 1933 1596 1934
rect 1988 1934 2044 1937
rect 1988 1933 1993 1934
rect 1591 1903 1757 1933
rect 1827 1903 1993 1933
rect 2039 1933 2044 1934
rect 2436 1934 2492 1937
rect 2436 1933 2441 1934
rect 2039 1903 2205 1933
rect 2275 1903 2441 1933
rect 2487 1933 2492 1934
rect 2884 1934 2940 1937
rect 2884 1933 2889 1934
rect 2487 1903 2653 1933
rect 2723 1903 2889 1933
rect 2935 1933 2940 1934
rect 3332 1934 3388 1937
rect 3332 1933 3337 1934
rect 2935 1903 3101 1933
rect 3171 1903 3337 1933
rect 3383 1933 3388 1934
rect 3780 1934 3836 1937
rect 3780 1933 3785 1934
rect 3383 1903 3549 1933
rect 3619 1903 3785 1933
rect 3831 1933 3836 1934
rect 4228 1934 4284 1937
rect 4228 1933 4233 1934
rect 3831 1903 3997 1933
rect 4067 1903 4233 1933
rect 4279 1933 4284 1934
rect 4676 1934 4732 1937
rect 4676 1933 4681 1934
rect 4279 1903 4445 1933
rect 4515 1903 4681 1933
rect 4727 1933 4732 1934
rect 5124 1934 5180 1937
rect 5124 1933 5129 1934
rect 4727 1903 4893 1933
rect 4963 1903 5129 1933
rect 5175 1933 5180 1934
rect 5572 1934 5628 1937
rect 5572 1933 5577 1934
rect 5175 1903 5341 1933
rect 5411 1903 5577 1933
rect 5623 1933 5628 1934
rect 6020 1934 6076 1937
rect 6020 1933 6025 1934
rect 5623 1903 5789 1933
rect 5859 1903 6025 1933
rect 6071 1933 6076 1934
rect 6468 1934 6524 1937
rect 6468 1933 6473 1934
rect 6071 1903 6237 1933
rect 6307 1903 6473 1933
rect 6519 1933 6524 1934
rect 6916 1934 6972 1937
rect 6916 1933 6921 1934
rect 6519 1903 6685 1933
rect 6755 1903 6921 1933
rect 6967 1933 6972 1934
rect 7364 1934 7420 1937
rect 7364 1933 7369 1934
rect 6967 1903 7133 1933
rect 7203 1903 7369 1933
rect 7415 1933 7420 1934
rect 7812 1934 7868 1937
rect 7812 1933 7817 1934
rect 7415 1903 7581 1933
rect 7651 1903 7817 1933
rect 7863 1933 7868 1934
rect 8260 1934 8316 1937
rect 8260 1933 8265 1934
rect 7863 1903 8029 1933
rect 8099 1903 8265 1933
rect 8311 1933 8316 1934
rect 8708 1934 8764 1937
rect 8708 1933 8713 1934
rect 8311 1903 8477 1933
rect 8547 1903 8713 1933
rect 8759 1933 8764 1934
rect 8759 1903 8925 1933
rect 196 1899 252 1903
rect 644 1899 700 1903
rect 1092 1899 1148 1903
rect 1540 1899 1596 1903
rect 1988 1899 2044 1903
rect 2436 1899 2492 1903
rect 2884 1899 2940 1903
rect 3332 1899 3388 1903
rect 3780 1899 3836 1903
rect 4228 1899 4284 1903
rect 4676 1899 4732 1903
rect 5124 1899 5180 1903
rect 5572 1899 5628 1903
rect 6020 1899 6076 1903
rect 6468 1899 6524 1903
rect 6916 1899 6972 1903
rect 7364 1899 7420 1903
rect 7812 1899 7868 1903
rect 8260 1899 8316 1903
rect 8708 1899 8764 1903
rect 196 1812 252 1815
rect 196 1811 201 1812
rect 35 1781 201 1811
rect 247 1811 252 1812
rect 644 1812 700 1815
rect 644 1811 649 1812
rect 247 1781 413 1811
rect 483 1781 649 1811
rect 695 1811 700 1812
rect 1092 1812 1148 1815
rect 1092 1811 1097 1812
rect 695 1781 861 1811
rect 931 1781 1097 1811
rect 1143 1811 1148 1812
rect 1540 1812 1596 1815
rect 1540 1811 1545 1812
rect 1143 1781 1309 1811
rect 1379 1781 1545 1811
rect 1591 1811 1596 1812
rect 1988 1812 2044 1815
rect 1988 1811 1993 1812
rect 1591 1781 1757 1811
rect 1827 1781 1993 1811
rect 2039 1811 2044 1812
rect 2436 1812 2492 1815
rect 2436 1811 2441 1812
rect 2039 1781 2205 1811
rect 2275 1781 2441 1811
rect 2487 1811 2492 1812
rect 2884 1812 2940 1815
rect 2884 1811 2889 1812
rect 2487 1781 2653 1811
rect 2723 1781 2889 1811
rect 2935 1811 2940 1812
rect 3332 1812 3388 1815
rect 3332 1811 3337 1812
rect 2935 1781 3101 1811
rect 3171 1781 3337 1811
rect 3383 1811 3388 1812
rect 3780 1812 3836 1815
rect 3780 1811 3785 1812
rect 3383 1781 3549 1811
rect 3619 1781 3785 1811
rect 3831 1811 3836 1812
rect 4228 1812 4284 1815
rect 4228 1811 4233 1812
rect 3831 1781 3997 1811
rect 4067 1781 4233 1811
rect 4279 1811 4284 1812
rect 4676 1812 4732 1815
rect 4676 1811 4681 1812
rect 4279 1781 4445 1811
rect 4515 1781 4681 1811
rect 4727 1811 4732 1812
rect 5124 1812 5180 1815
rect 5124 1811 5129 1812
rect 4727 1781 4893 1811
rect 4963 1781 5129 1811
rect 5175 1811 5180 1812
rect 5572 1812 5628 1815
rect 5572 1811 5577 1812
rect 5175 1781 5341 1811
rect 5411 1781 5577 1811
rect 5623 1811 5628 1812
rect 6020 1812 6076 1815
rect 6020 1811 6025 1812
rect 5623 1781 5789 1811
rect 5859 1781 6025 1811
rect 6071 1811 6076 1812
rect 6468 1812 6524 1815
rect 6468 1811 6473 1812
rect 6071 1781 6237 1811
rect 6307 1781 6473 1811
rect 6519 1811 6524 1812
rect 6916 1812 6972 1815
rect 6916 1811 6921 1812
rect 6519 1781 6685 1811
rect 6755 1781 6921 1811
rect 6967 1811 6972 1812
rect 7364 1812 7420 1815
rect 7364 1811 7369 1812
rect 6967 1781 7133 1811
rect 7203 1781 7369 1811
rect 7415 1811 7420 1812
rect 7812 1812 7868 1815
rect 7812 1811 7817 1812
rect 7415 1781 7581 1811
rect 7651 1781 7817 1811
rect 7863 1811 7868 1812
rect 8260 1812 8316 1815
rect 8260 1811 8265 1812
rect 7863 1781 8029 1811
rect 8099 1781 8265 1811
rect 8311 1811 8316 1812
rect 8708 1812 8764 1815
rect 8708 1811 8713 1812
rect 8311 1781 8477 1811
rect 8547 1781 8713 1811
rect 8759 1811 8764 1812
rect 8759 1781 8925 1811
rect 196 1777 252 1781
rect 644 1777 700 1781
rect 1092 1777 1148 1781
rect 1540 1777 1596 1781
rect 1988 1777 2044 1781
rect 2436 1777 2492 1781
rect 2884 1777 2940 1781
rect 3332 1777 3388 1781
rect 3780 1777 3836 1781
rect 4228 1777 4284 1781
rect 4676 1777 4732 1781
rect 5124 1777 5180 1781
rect 5572 1777 5628 1781
rect 6020 1777 6076 1781
rect 6468 1777 6524 1781
rect 6916 1777 6972 1781
rect 7364 1777 7420 1781
rect 7812 1777 7868 1781
rect 8260 1777 8316 1781
rect 8708 1777 8764 1781
rect 99 1749 137 1750
rect 99 1748 102 1749
rect 54 1718 102 1748
rect 99 1717 102 1718
rect 134 1748 137 1749
rect 311 1749 349 1750
rect 311 1748 314 1749
rect 134 1718 181 1748
rect 267 1718 314 1748
rect 134 1717 137 1718
rect 99 1716 137 1717
rect 311 1717 314 1718
rect 346 1748 349 1749
rect 547 1749 585 1750
rect 547 1748 550 1749
rect 346 1718 394 1748
rect 502 1718 550 1748
rect 346 1717 349 1718
rect 311 1716 349 1717
rect 547 1717 550 1718
rect 582 1748 585 1749
rect 759 1749 797 1750
rect 759 1748 762 1749
rect 582 1718 629 1748
rect 715 1718 762 1748
rect 582 1717 585 1718
rect 547 1716 585 1717
rect 759 1717 762 1718
rect 794 1748 797 1749
rect 995 1749 1033 1750
rect 995 1748 998 1749
rect 794 1718 842 1748
rect 950 1718 998 1748
rect 794 1717 797 1718
rect 759 1716 797 1717
rect 995 1717 998 1718
rect 1030 1748 1033 1749
rect 1207 1749 1245 1750
rect 1207 1748 1210 1749
rect 1030 1718 1077 1748
rect 1163 1718 1210 1748
rect 1030 1717 1033 1718
rect 995 1716 1033 1717
rect 1207 1717 1210 1718
rect 1242 1748 1245 1749
rect 1443 1749 1481 1750
rect 1443 1748 1446 1749
rect 1242 1718 1290 1748
rect 1398 1718 1446 1748
rect 1242 1717 1245 1718
rect 1207 1716 1245 1717
rect 1443 1717 1446 1718
rect 1478 1748 1481 1749
rect 1655 1749 1693 1750
rect 1655 1748 1658 1749
rect 1478 1718 1525 1748
rect 1611 1718 1658 1748
rect 1478 1717 1481 1718
rect 1443 1716 1481 1717
rect 1655 1717 1658 1718
rect 1690 1748 1693 1749
rect 1891 1749 1929 1750
rect 1891 1748 1894 1749
rect 1690 1718 1738 1748
rect 1846 1718 1894 1748
rect 1690 1717 1693 1718
rect 1655 1716 1693 1717
rect 1891 1717 1894 1718
rect 1926 1748 1929 1749
rect 2103 1749 2141 1750
rect 2103 1748 2106 1749
rect 1926 1718 1973 1748
rect 2059 1718 2106 1748
rect 1926 1717 1929 1718
rect 1891 1716 1929 1717
rect 2103 1717 2106 1718
rect 2138 1748 2141 1749
rect 2339 1749 2377 1750
rect 2339 1748 2342 1749
rect 2138 1718 2186 1748
rect 2294 1718 2342 1748
rect 2138 1717 2141 1718
rect 2103 1716 2141 1717
rect 2339 1717 2342 1718
rect 2374 1748 2377 1749
rect 2551 1749 2589 1750
rect 2551 1748 2554 1749
rect 2374 1718 2421 1748
rect 2507 1718 2554 1748
rect 2374 1717 2377 1718
rect 2339 1716 2377 1717
rect 2551 1717 2554 1718
rect 2586 1748 2589 1749
rect 2787 1749 2825 1750
rect 2787 1748 2790 1749
rect 2586 1718 2634 1748
rect 2742 1718 2790 1748
rect 2586 1717 2589 1718
rect 2551 1716 2589 1717
rect 2787 1717 2790 1718
rect 2822 1748 2825 1749
rect 2999 1749 3037 1750
rect 2999 1748 3002 1749
rect 2822 1718 2869 1748
rect 2955 1718 3002 1748
rect 2822 1717 2825 1718
rect 2787 1716 2825 1717
rect 2999 1717 3002 1718
rect 3034 1748 3037 1749
rect 3235 1749 3273 1750
rect 3235 1748 3238 1749
rect 3034 1718 3082 1748
rect 3190 1718 3238 1748
rect 3034 1717 3037 1718
rect 2999 1716 3037 1717
rect 3235 1717 3238 1718
rect 3270 1748 3273 1749
rect 3447 1749 3485 1750
rect 3447 1748 3450 1749
rect 3270 1718 3317 1748
rect 3403 1718 3450 1748
rect 3270 1717 3273 1718
rect 3235 1716 3273 1717
rect 3447 1717 3450 1718
rect 3482 1748 3485 1749
rect 3683 1749 3721 1750
rect 3683 1748 3686 1749
rect 3482 1718 3530 1748
rect 3638 1718 3686 1748
rect 3482 1717 3485 1718
rect 3447 1716 3485 1717
rect 3683 1717 3686 1718
rect 3718 1748 3721 1749
rect 3895 1749 3933 1750
rect 3895 1748 3898 1749
rect 3718 1718 3765 1748
rect 3851 1718 3898 1748
rect 3718 1717 3721 1718
rect 3683 1716 3721 1717
rect 3895 1717 3898 1718
rect 3930 1748 3933 1749
rect 4131 1749 4169 1750
rect 4131 1748 4134 1749
rect 3930 1718 3978 1748
rect 4086 1718 4134 1748
rect 3930 1717 3933 1718
rect 3895 1716 3933 1717
rect 4131 1717 4134 1718
rect 4166 1748 4169 1749
rect 4343 1749 4381 1750
rect 4343 1748 4346 1749
rect 4166 1718 4213 1748
rect 4299 1718 4346 1748
rect 4166 1717 4169 1718
rect 4131 1716 4169 1717
rect 4343 1717 4346 1718
rect 4378 1748 4381 1749
rect 4579 1749 4617 1750
rect 4579 1748 4582 1749
rect 4378 1718 4426 1748
rect 4534 1718 4582 1748
rect 4378 1717 4381 1718
rect 4343 1716 4381 1717
rect 4579 1717 4582 1718
rect 4614 1748 4617 1749
rect 4791 1749 4829 1750
rect 4791 1748 4794 1749
rect 4614 1718 4661 1748
rect 4747 1718 4794 1748
rect 4614 1717 4617 1718
rect 4579 1716 4617 1717
rect 4791 1717 4794 1718
rect 4826 1748 4829 1749
rect 5027 1749 5065 1750
rect 5027 1748 5030 1749
rect 4826 1718 4874 1748
rect 4982 1718 5030 1748
rect 4826 1717 4829 1718
rect 4791 1716 4829 1717
rect 5027 1717 5030 1718
rect 5062 1748 5065 1749
rect 5239 1749 5277 1750
rect 5239 1748 5242 1749
rect 5062 1718 5109 1748
rect 5195 1718 5242 1748
rect 5062 1717 5065 1718
rect 5027 1716 5065 1717
rect 5239 1717 5242 1718
rect 5274 1748 5277 1749
rect 5475 1749 5513 1750
rect 5475 1748 5478 1749
rect 5274 1718 5322 1748
rect 5430 1718 5478 1748
rect 5274 1717 5277 1718
rect 5239 1716 5277 1717
rect 5475 1717 5478 1718
rect 5510 1748 5513 1749
rect 5687 1749 5725 1750
rect 5687 1748 5690 1749
rect 5510 1718 5557 1748
rect 5643 1718 5690 1748
rect 5510 1717 5513 1718
rect 5475 1716 5513 1717
rect 5687 1717 5690 1718
rect 5722 1748 5725 1749
rect 5923 1749 5961 1750
rect 5923 1748 5926 1749
rect 5722 1718 5770 1748
rect 5878 1718 5926 1748
rect 5722 1717 5725 1718
rect 5687 1716 5725 1717
rect 5923 1717 5926 1718
rect 5958 1748 5961 1749
rect 6135 1749 6173 1750
rect 6135 1748 6138 1749
rect 5958 1718 6005 1748
rect 6091 1718 6138 1748
rect 5958 1717 5961 1718
rect 5923 1716 5961 1717
rect 6135 1717 6138 1718
rect 6170 1748 6173 1749
rect 6371 1749 6409 1750
rect 6371 1748 6374 1749
rect 6170 1718 6218 1748
rect 6326 1718 6374 1748
rect 6170 1717 6173 1718
rect 6135 1716 6173 1717
rect 6371 1717 6374 1718
rect 6406 1748 6409 1749
rect 6583 1749 6621 1750
rect 6583 1748 6586 1749
rect 6406 1718 6453 1748
rect 6539 1718 6586 1748
rect 6406 1717 6409 1718
rect 6371 1716 6409 1717
rect 6583 1717 6586 1718
rect 6618 1748 6621 1749
rect 6819 1749 6857 1750
rect 6819 1748 6822 1749
rect 6618 1718 6666 1748
rect 6774 1718 6822 1748
rect 6618 1717 6621 1718
rect 6583 1716 6621 1717
rect 6819 1717 6822 1718
rect 6854 1748 6857 1749
rect 7031 1749 7069 1750
rect 7031 1748 7034 1749
rect 6854 1718 6901 1748
rect 6987 1718 7034 1748
rect 6854 1717 6857 1718
rect 6819 1716 6857 1717
rect 7031 1717 7034 1718
rect 7066 1748 7069 1749
rect 7267 1749 7305 1750
rect 7267 1748 7270 1749
rect 7066 1718 7114 1748
rect 7222 1718 7270 1748
rect 7066 1717 7069 1718
rect 7031 1716 7069 1717
rect 7267 1717 7270 1718
rect 7302 1748 7305 1749
rect 7479 1749 7517 1750
rect 7479 1748 7482 1749
rect 7302 1718 7349 1748
rect 7435 1718 7482 1748
rect 7302 1717 7305 1718
rect 7267 1716 7305 1717
rect 7479 1717 7482 1718
rect 7514 1748 7517 1749
rect 7715 1749 7753 1750
rect 7715 1748 7718 1749
rect 7514 1718 7562 1748
rect 7670 1718 7718 1748
rect 7514 1717 7517 1718
rect 7479 1716 7517 1717
rect 7715 1717 7718 1718
rect 7750 1748 7753 1749
rect 7927 1749 7965 1750
rect 7927 1748 7930 1749
rect 7750 1718 7797 1748
rect 7883 1718 7930 1748
rect 7750 1717 7753 1718
rect 7715 1716 7753 1717
rect 7927 1717 7930 1718
rect 7962 1748 7965 1749
rect 8163 1749 8201 1750
rect 8163 1748 8166 1749
rect 7962 1718 8010 1748
rect 8118 1718 8166 1748
rect 7962 1717 7965 1718
rect 7927 1716 7965 1717
rect 8163 1717 8166 1718
rect 8198 1748 8201 1749
rect 8375 1749 8413 1750
rect 8375 1748 8378 1749
rect 8198 1718 8245 1748
rect 8331 1718 8378 1748
rect 8198 1717 8201 1718
rect 8163 1716 8201 1717
rect 8375 1717 8378 1718
rect 8410 1748 8413 1749
rect 8611 1749 8649 1750
rect 8611 1748 8614 1749
rect 8410 1718 8458 1748
rect 8566 1718 8614 1748
rect 8410 1717 8413 1718
rect 8375 1716 8413 1717
rect 8611 1717 8614 1718
rect 8646 1748 8649 1749
rect 8823 1749 8861 1750
rect 8823 1748 8826 1749
rect 8646 1718 8693 1748
rect 8779 1718 8826 1748
rect 8646 1717 8649 1718
rect 8611 1716 8649 1717
rect 8823 1717 8826 1718
rect 8858 1748 8861 1749
rect 8858 1718 8906 1748
rect 8858 1717 8861 1718
rect 8823 1716 8861 1717
rect 196 1687 252 1690
rect 196 1686 201 1687
rect 35 1656 201 1686
rect 247 1686 252 1687
rect 644 1687 700 1690
rect 644 1686 649 1687
rect 247 1656 413 1686
rect 483 1656 649 1686
rect 695 1686 700 1687
rect 1092 1687 1148 1690
rect 1092 1686 1097 1687
rect 695 1656 861 1686
rect 931 1656 1097 1686
rect 1143 1686 1148 1687
rect 1540 1687 1596 1690
rect 1540 1686 1545 1687
rect 1143 1656 1309 1686
rect 1379 1656 1545 1686
rect 1591 1686 1596 1687
rect 1988 1687 2044 1690
rect 1988 1686 1993 1687
rect 1591 1656 1757 1686
rect 1827 1656 1993 1686
rect 2039 1686 2044 1687
rect 2436 1687 2492 1690
rect 2436 1686 2441 1687
rect 2039 1656 2205 1686
rect 2275 1656 2441 1686
rect 2487 1686 2492 1687
rect 2884 1687 2940 1690
rect 2884 1686 2889 1687
rect 2487 1656 2653 1686
rect 2723 1656 2889 1686
rect 2935 1686 2940 1687
rect 3332 1687 3388 1690
rect 3332 1686 3337 1687
rect 2935 1656 3101 1686
rect 3171 1656 3337 1686
rect 3383 1686 3388 1687
rect 3780 1687 3836 1690
rect 3780 1686 3785 1687
rect 3383 1656 3549 1686
rect 3619 1656 3785 1686
rect 3831 1686 3836 1687
rect 4228 1687 4284 1690
rect 4228 1686 4233 1687
rect 3831 1656 3997 1686
rect 4067 1656 4233 1686
rect 4279 1686 4284 1687
rect 4676 1687 4732 1690
rect 4676 1686 4681 1687
rect 4279 1656 4445 1686
rect 4515 1656 4681 1686
rect 4727 1686 4732 1687
rect 5124 1687 5180 1690
rect 5124 1686 5129 1687
rect 4727 1656 4893 1686
rect 4963 1656 5129 1686
rect 5175 1686 5180 1687
rect 5572 1687 5628 1690
rect 5572 1686 5577 1687
rect 5175 1656 5341 1686
rect 5411 1656 5577 1686
rect 5623 1686 5628 1687
rect 6020 1687 6076 1690
rect 6020 1686 6025 1687
rect 5623 1656 5789 1686
rect 5859 1656 6025 1686
rect 6071 1686 6076 1687
rect 6468 1687 6524 1690
rect 6468 1686 6473 1687
rect 6071 1656 6237 1686
rect 6307 1656 6473 1686
rect 6519 1686 6524 1687
rect 6916 1687 6972 1690
rect 6916 1686 6921 1687
rect 6519 1656 6685 1686
rect 6755 1656 6921 1686
rect 6967 1686 6972 1687
rect 7364 1687 7420 1690
rect 7364 1686 7369 1687
rect 6967 1656 7133 1686
rect 7203 1656 7369 1686
rect 7415 1686 7420 1687
rect 7812 1687 7868 1690
rect 7812 1686 7817 1687
rect 7415 1656 7581 1686
rect 7651 1656 7817 1686
rect 7863 1686 7868 1687
rect 8260 1687 8316 1690
rect 8260 1686 8265 1687
rect 7863 1656 8029 1686
rect 8099 1656 8265 1686
rect 8311 1686 8316 1687
rect 8708 1687 8764 1690
rect 8708 1686 8713 1687
rect 8311 1656 8477 1686
rect 8547 1656 8713 1686
rect 8759 1686 8764 1687
rect 8759 1656 8925 1686
rect 196 1652 252 1656
rect 644 1652 700 1656
rect 1092 1652 1148 1656
rect 1540 1652 1596 1656
rect 1988 1652 2044 1656
rect 2436 1652 2492 1656
rect 2884 1652 2940 1656
rect 3332 1652 3388 1656
rect 3780 1652 3836 1656
rect 4228 1652 4284 1656
rect 4676 1652 4732 1656
rect 5124 1652 5180 1656
rect 5572 1652 5628 1656
rect 6020 1652 6076 1656
rect 6468 1652 6524 1656
rect 6916 1652 6972 1656
rect 7364 1652 7420 1656
rect 7812 1652 7868 1656
rect 8260 1652 8316 1656
rect 8708 1652 8764 1656
rect 99 1625 137 1626
rect 99 1624 102 1625
rect 54 1594 102 1624
rect 99 1593 102 1594
rect 134 1624 137 1625
rect 311 1625 349 1626
rect 311 1624 314 1625
rect 134 1594 181 1624
rect 267 1594 314 1624
rect 134 1593 137 1594
rect 99 1592 137 1593
rect 311 1593 314 1594
rect 346 1624 349 1625
rect 547 1625 585 1626
rect 547 1624 550 1625
rect 346 1594 394 1624
rect 502 1594 550 1624
rect 346 1593 349 1594
rect 311 1592 349 1593
rect 547 1593 550 1594
rect 582 1624 585 1625
rect 759 1625 797 1626
rect 759 1624 762 1625
rect 582 1594 629 1624
rect 715 1594 762 1624
rect 582 1593 585 1594
rect 547 1592 585 1593
rect 759 1593 762 1594
rect 794 1624 797 1625
rect 995 1625 1033 1626
rect 995 1624 998 1625
rect 794 1594 842 1624
rect 950 1594 998 1624
rect 794 1593 797 1594
rect 759 1592 797 1593
rect 995 1593 998 1594
rect 1030 1624 1033 1625
rect 1207 1625 1245 1626
rect 1207 1624 1210 1625
rect 1030 1594 1077 1624
rect 1163 1594 1210 1624
rect 1030 1593 1033 1594
rect 995 1592 1033 1593
rect 1207 1593 1210 1594
rect 1242 1624 1245 1625
rect 1443 1625 1481 1626
rect 1443 1624 1446 1625
rect 1242 1594 1290 1624
rect 1398 1594 1446 1624
rect 1242 1593 1245 1594
rect 1207 1592 1245 1593
rect 1443 1593 1446 1594
rect 1478 1624 1481 1625
rect 1655 1625 1693 1626
rect 1655 1624 1658 1625
rect 1478 1594 1525 1624
rect 1611 1594 1658 1624
rect 1478 1593 1481 1594
rect 1443 1592 1481 1593
rect 1655 1593 1658 1594
rect 1690 1624 1693 1625
rect 1891 1625 1929 1626
rect 1891 1624 1894 1625
rect 1690 1594 1738 1624
rect 1846 1594 1894 1624
rect 1690 1593 1693 1594
rect 1655 1592 1693 1593
rect 1891 1593 1894 1594
rect 1926 1624 1929 1625
rect 2103 1625 2141 1626
rect 2103 1624 2106 1625
rect 1926 1594 1973 1624
rect 2059 1594 2106 1624
rect 1926 1593 1929 1594
rect 1891 1592 1929 1593
rect 2103 1593 2106 1594
rect 2138 1624 2141 1625
rect 2339 1625 2377 1626
rect 2339 1624 2342 1625
rect 2138 1594 2186 1624
rect 2294 1594 2342 1624
rect 2138 1593 2141 1594
rect 2103 1592 2141 1593
rect 2339 1593 2342 1594
rect 2374 1624 2377 1625
rect 2551 1625 2589 1626
rect 2551 1624 2554 1625
rect 2374 1594 2421 1624
rect 2507 1594 2554 1624
rect 2374 1593 2377 1594
rect 2339 1592 2377 1593
rect 2551 1593 2554 1594
rect 2586 1624 2589 1625
rect 2787 1625 2825 1626
rect 2787 1624 2790 1625
rect 2586 1594 2634 1624
rect 2742 1594 2790 1624
rect 2586 1593 2589 1594
rect 2551 1592 2589 1593
rect 2787 1593 2790 1594
rect 2822 1624 2825 1625
rect 2999 1625 3037 1626
rect 2999 1624 3002 1625
rect 2822 1594 2869 1624
rect 2955 1594 3002 1624
rect 2822 1593 2825 1594
rect 2787 1592 2825 1593
rect 2999 1593 3002 1594
rect 3034 1624 3037 1625
rect 3235 1625 3273 1626
rect 3235 1624 3238 1625
rect 3034 1594 3082 1624
rect 3190 1594 3238 1624
rect 3034 1593 3037 1594
rect 2999 1592 3037 1593
rect 3235 1593 3238 1594
rect 3270 1624 3273 1625
rect 3447 1625 3485 1626
rect 3447 1624 3450 1625
rect 3270 1594 3317 1624
rect 3403 1594 3450 1624
rect 3270 1593 3273 1594
rect 3235 1592 3273 1593
rect 3447 1593 3450 1594
rect 3482 1624 3485 1625
rect 3683 1625 3721 1626
rect 3683 1624 3686 1625
rect 3482 1594 3530 1624
rect 3638 1594 3686 1624
rect 3482 1593 3485 1594
rect 3447 1592 3485 1593
rect 3683 1593 3686 1594
rect 3718 1624 3721 1625
rect 3895 1625 3933 1626
rect 3895 1624 3898 1625
rect 3718 1594 3765 1624
rect 3851 1594 3898 1624
rect 3718 1593 3721 1594
rect 3683 1592 3721 1593
rect 3895 1593 3898 1594
rect 3930 1624 3933 1625
rect 4131 1625 4169 1626
rect 4131 1624 4134 1625
rect 3930 1594 3978 1624
rect 4086 1594 4134 1624
rect 3930 1593 3933 1594
rect 3895 1592 3933 1593
rect 4131 1593 4134 1594
rect 4166 1624 4169 1625
rect 4343 1625 4381 1626
rect 4343 1624 4346 1625
rect 4166 1594 4213 1624
rect 4299 1594 4346 1624
rect 4166 1593 4169 1594
rect 4131 1592 4169 1593
rect 4343 1593 4346 1594
rect 4378 1624 4381 1625
rect 4579 1625 4617 1626
rect 4579 1624 4582 1625
rect 4378 1594 4426 1624
rect 4534 1594 4582 1624
rect 4378 1593 4381 1594
rect 4343 1592 4381 1593
rect 4579 1593 4582 1594
rect 4614 1624 4617 1625
rect 4791 1625 4829 1626
rect 4791 1624 4794 1625
rect 4614 1594 4661 1624
rect 4747 1594 4794 1624
rect 4614 1593 4617 1594
rect 4579 1592 4617 1593
rect 4791 1593 4794 1594
rect 4826 1624 4829 1625
rect 5027 1625 5065 1626
rect 5027 1624 5030 1625
rect 4826 1594 4874 1624
rect 4982 1594 5030 1624
rect 4826 1593 4829 1594
rect 4791 1592 4829 1593
rect 5027 1593 5030 1594
rect 5062 1624 5065 1625
rect 5239 1625 5277 1626
rect 5239 1624 5242 1625
rect 5062 1594 5109 1624
rect 5195 1594 5242 1624
rect 5062 1593 5065 1594
rect 5027 1592 5065 1593
rect 5239 1593 5242 1594
rect 5274 1624 5277 1625
rect 5475 1625 5513 1626
rect 5475 1624 5478 1625
rect 5274 1594 5322 1624
rect 5430 1594 5478 1624
rect 5274 1593 5277 1594
rect 5239 1592 5277 1593
rect 5475 1593 5478 1594
rect 5510 1624 5513 1625
rect 5687 1625 5725 1626
rect 5687 1624 5690 1625
rect 5510 1594 5557 1624
rect 5643 1594 5690 1624
rect 5510 1593 5513 1594
rect 5475 1592 5513 1593
rect 5687 1593 5690 1594
rect 5722 1624 5725 1625
rect 5923 1625 5961 1626
rect 5923 1624 5926 1625
rect 5722 1594 5770 1624
rect 5878 1594 5926 1624
rect 5722 1593 5725 1594
rect 5687 1592 5725 1593
rect 5923 1593 5926 1594
rect 5958 1624 5961 1625
rect 6135 1625 6173 1626
rect 6135 1624 6138 1625
rect 5958 1594 6005 1624
rect 6091 1594 6138 1624
rect 5958 1593 5961 1594
rect 5923 1592 5961 1593
rect 6135 1593 6138 1594
rect 6170 1624 6173 1625
rect 6371 1625 6409 1626
rect 6371 1624 6374 1625
rect 6170 1594 6218 1624
rect 6326 1594 6374 1624
rect 6170 1593 6173 1594
rect 6135 1592 6173 1593
rect 6371 1593 6374 1594
rect 6406 1624 6409 1625
rect 6583 1625 6621 1626
rect 6583 1624 6586 1625
rect 6406 1594 6453 1624
rect 6539 1594 6586 1624
rect 6406 1593 6409 1594
rect 6371 1592 6409 1593
rect 6583 1593 6586 1594
rect 6618 1624 6621 1625
rect 6819 1625 6857 1626
rect 6819 1624 6822 1625
rect 6618 1594 6666 1624
rect 6774 1594 6822 1624
rect 6618 1593 6621 1594
rect 6583 1592 6621 1593
rect 6819 1593 6822 1594
rect 6854 1624 6857 1625
rect 7031 1625 7069 1626
rect 7031 1624 7034 1625
rect 6854 1594 6901 1624
rect 6987 1594 7034 1624
rect 6854 1593 6857 1594
rect 6819 1592 6857 1593
rect 7031 1593 7034 1594
rect 7066 1624 7069 1625
rect 7267 1625 7305 1626
rect 7267 1624 7270 1625
rect 7066 1594 7114 1624
rect 7222 1594 7270 1624
rect 7066 1593 7069 1594
rect 7031 1592 7069 1593
rect 7267 1593 7270 1594
rect 7302 1624 7305 1625
rect 7479 1625 7517 1626
rect 7479 1624 7482 1625
rect 7302 1594 7349 1624
rect 7435 1594 7482 1624
rect 7302 1593 7305 1594
rect 7267 1592 7305 1593
rect 7479 1593 7482 1594
rect 7514 1624 7517 1625
rect 7715 1625 7753 1626
rect 7715 1624 7718 1625
rect 7514 1594 7562 1624
rect 7670 1594 7718 1624
rect 7514 1593 7517 1594
rect 7479 1592 7517 1593
rect 7715 1593 7718 1594
rect 7750 1624 7753 1625
rect 7927 1625 7965 1626
rect 7927 1624 7930 1625
rect 7750 1594 7797 1624
rect 7883 1594 7930 1624
rect 7750 1593 7753 1594
rect 7715 1592 7753 1593
rect 7927 1593 7930 1594
rect 7962 1624 7965 1625
rect 8163 1625 8201 1626
rect 8163 1624 8166 1625
rect 7962 1594 8010 1624
rect 8118 1594 8166 1624
rect 7962 1593 7965 1594
rect 7927 1592 7965 1593
rect 8163 1593 8166 1594
rect 8198 1624 8201 1625
rect 8375 1625 8413 1626
rect 8375 1624 8378 1625
rect 8198 1594 8245 1624
rect 8331 1594 8378 1624
rect 8198 1593 8201 1594
rect 8163 1592 8201 1593
rect 8375 1593 8378 1594
rect 8410 1624 8413 1625
rect 8611 1625 8649 1626
rect 8611 1624 8614 1625
rect 8410 1594 8458 1624
rect 8566 1594 8614 1624
rect 8410 1593 8413 1594
rect 8375 1592 8413 1593
rect 8611 1593 8614 1594
rect 8646 1624 8649 1625
rect 8823 1625 8861 1626
rect 8823 1624 8826 1625
rect 8646 1594 8693 1624
rect 8779 1594 8826 1624
rect 8646 1593 8649 1594
rect 8611 1592 8649 1593
rect 8823 1593 8826 1594
rect 8858 1624 8861 1625
rect 8858 1594 8906 1624
rect 8858 1593 8861 1594
rect 8823 1592 8861 1593
rect 196 1563 252 1566
rect 196 1562 201 1563
rect 35 1532 201 1562
rect 247 1562 252 1563
rect 644 1563 700 1566
rect 644 1562 649 1563
rect 247 1532 413 1562
rect 483 1532 649 1562
rect 695 1562 700 1563
rect 1092 1563 1148 1566
rect 1092 1562 1097 1563
rect 695 1532 861 1562
rect 931 1532 1097 1562
rect 1143 1562 1148 1563
rect 1540 1563 1596 1566
rect 1540 1562 1545 1563
rect 1143 1532 1309 1562
rect 1379 1532 1545 1562
rect 1591 1562 1596 1563
rect 1988 1563 2044 1566
rect 1988 1562 1993 1563
rect 1591 1532 1757 1562
rect 1827 1532 1993 1562
rect 2039 1562 2044 1563
rect 2436 1563 2492 1566
rect 2436 1562 2441 1563
rect 2039 1532 2205 1562
rect 2275 1532 2441 1562
rect 2487 1562 2492 1563
rect 2884 1563 2940 1566
rect 2884 1562 2889 1563
rect 2487 1532 2653 1562
rect 2723 1532 2889 1562
rect 2935 1562 2940 1563
rect 3332 1563 3388 1566
rect 3332 1562 3337 1563
rect 2935 1532 3101 1562
rect 3171 1532 3337 1562
rect 3383 1562 3388 1563
rect 3780 1563 3836 1566
rect 3780 1562 3785 1563
rect 3383 1532 3549 1562
rect 3619 1532 3785 1562
rect 3831 1562 3836 1563
rect 4228 1563 4284 1566
rect 4228 1562 4233 1563
rect 3831 1532 3997 1562
rect 4067 1532 4233 1562
rect 4279 1562 4284 1563
rect 4676 1563 4732 1566
rect 4676 1562 4681 1563
rect 4279 1532 4445 1562
rect 4515 1532 4681 1562
rect 4727 1562 4732 1563
rect 5124 1563 5180 1566
rect 5124 1562 5129 1563
rect 4727 1532 4893 1562
rect 4963 1532 5129 1562
rect 5175 1562 5180 1563
rect 5572 1563 5628 1566
rect 5572 1562 5577 1563
rect 5175 1532 5341 1562
rect 5411 1532 5577 1562
rect 5623 1562 5628 1563
rect 6020 1563 6076 1566
rect 6020 1562 6025 1563
rect 5623 1532 5789 1562
rect 5859 1532 6025 1562
rect 6071 1562 6076 1563
rect 6468 1563 6524 1566
rect 6468 1562 6473 1563
rect 6071 1532 6237 1562
rect 6307 1532 6473 1562
rect 6519 1562 6524 1563
rect 6916 1563 6972 1566
rect 6916 1562 6921 1563
rect 6519 1532 6685 1562
rect 6755 1532 6921 1562
rect 6967 1562 6972 1563
rect 7364 1563 7420 1566
rect 7364 1562 7369 1563
rect 6967 1532 7133 1562
rect 7203 1532 7369 1562
rect 7415 1562 7420 1563
rect 7812 1563 7868 1566
rect 7812 1562 7817 1563
rect 7415 1532 7581 1562
rect 7651 1532 7817 1562
rect 7863 1562 7868 1563
rect 8260 1563 8316 1566
rect 8260 1562 8265 1563
rect 7863 1532 8029 1562
rect 8099 1532 8265 1562
rect 8311 1562 8316 1563
rect 8708 1563 8764 1566
rect 8708 1562 8713 1563
rect 8311 1532 8477 1562
rect 8547 1532 8713 1562
rect 8759 1562 8764 1563
rect 8759 1532 8925 1562
rect 196 1528 252 1532
rect 644 1528 700 1532
rect 1092 1528 1148 1532
rect 1540 1528 1596 1532
rect 1988 1528 2044 1532
rect 2436 1528 2492 1532
rect 2884 1528 2940 1532
rect 3332 1528 3388 1532
rect 3780 1528 3836 1532
rect 4228 1528 4284 1532
rect 4676 1528 4732 1532
rect 5124 1528 5180 1532
rect 5572 1528 5628 1532
rect 6020 1528 6076 1532
rect 6468 1528 6524 1532
rect 6916 1528 6972 1532
rect 7364 1528 7420 1532
rect 7812 1528 7868 1532
rect 8260 1528 8316 1532
rect 8708 1528 8764 1532
rect 99 1501 137 1502
rect 99 1500 102 1501
rect 54 1470 102 1500
rect 99 1469 102 1470
rect 134 1500 137 1501
rect 311 1501 349 1502
rect 311 1500 314 1501
rect 134 1470 181 1500
rect 267 1470 314 1500
rect 134 1469 137 1470
rect 99 1468 137 1469
rect 311 1469 314 1470
rect 346 1500 349 1501
rect 547 1501 585 1502
rect 547 1500 550 1501
rect 346 1470 394 1500
rect 502 1470 550 1500
rect 346 1469 349 1470
rect 311 1468 349 1469
rect 547 1469 550 1470
rect 582 1500 585 1501
rect 759 1501 797 1502
rect 759 1500 762 1501
rect 582 1470 629 1500
rect 715 1470 762 1500
rect 582 1469 585 1470
rect 547 1468 585 1469
rect 759 1469 762 1470
rect 794 1500 797 1501
rect 995 1501 1033 1502
rect 995 1500 998 1501
rect 794 1470 842 1500
rect 950 1470 998 1500
rect 794 1469 797 1470
rect 759 1468 797 1469
rect 995 1469 998 1470
rect 1030 1500 1033 1501
rect 1207 1501 1245 1502
rect 1207 1500 1210 1501
rect 1030 1470 1077 1500
rect 1163 1470 1210 1500
rect 1030 1469 1033 1470
rect 995 1468 1033 1469
rect 1207 1469 1210 1470
rect 1242 1500 1245 1501
rect 1443 1501 1481 1502
rect 1443 1500 1446 1501
rect 1242 1470 1290 1500
rect 1398 1470 1446 1500
rect 1242 1469 1245 1470
rect 1207 1468 1245 1469
rect 1443 1469 1446 1470
rect 1478 1500 1481 1501
rect 1655 1501 1693 1502
rect 1655 1500 1658 1501
rect 1478 1470 1525 1500
rect 1611 1470 1658 1500
rect 1478 1469 1481 1470
rect 1443 1468 1481 1469
rect 1655 1469 1658 1470
rect 1690 1500 1693 1501
rect 1891 1501 1929 1502
rect 1891 1500 1894 1501
rect 1690 1470 1738 1500
rect 1846 1470 1894 1500
rect 1690 1469 1693 1470
rect 1655 1468 1693 1469
rect 1891 1469 1894 1470
rect 1926 1500 1929 1501
rect 2103 1501 2141 1502
rect 2103 1500 2106 1501
rect 1926 1470 1973 1500
rect 2059 1470 2106 1500
rect 1926 1469 1929 1470
rect 1891 1468 1929 1469
rect 2103 1469 2106 1470
rect 2138 1500 2141 1501
rect 2339 1501 2377 1502
rect 2339 1500 2342 1501
rect 2138 1470 2186 1500
rect 2294 1470 2342 1500
rect 2138 1469 2141 1470
rect 2103 1468 2141 1469
rect 2339 1469 2342 1470
rect 2374 1500 2377 1501
rect 2551 1501 2589 1502
rect 2551 1500 2554 1501
rect 2374 1470 2421 1500
rect 2507 1470 2554 1500
rect 2374 1469 2377 1470
rect 2339 1468 2377 1469
rect 2551 1469 2554 1470
rect 2586 1500 2589 1501
rect 2787 1501 2825 1502
rect 2787 1500 2790 1501
rect 2586 1470 2634 1500
rect 2742 1470 2790 1500
rect 2586 1469 2589 1470
rect 2551 1468 2589 1469
rect 2787 1469 2790 1470
rect 2822 1500 2825 1501
rect 2999 1501 3037 1502
rect 2999 1500 3002 1501
rect 2822 1470 2869 1500
rect 2955 1470 3002 1500
rect 2822 1469 2825 1470
rect 2787 1468 2825 1469
rect 2999 1469 3002 1470
rect 3034 1500 3037 1501
rect 3235 1501 3273 1502
rect 3235 1500 3238 1501
rect 3034 1470 3082 1500
rect 3190 1470 3238 1500
rect 3034 1469 3037 1470
rect 2999 1468 3037 1469
rect 3235 1469 3238 1470
rect 3270 1500 3273 1501
rect 3447 1501 3485 1502
rect 3447 1500 3450 1501
rect 3270 1470 3317 1500
rect 3403 1470 3450 1500
rect 3270 1469 3273 1470
rect 3235 1468 3273 1469
rect 3447 1469 3450 1470
rect 3482 1500 3485 1501
rect 3683 1501 3721 1502
rect 3683 1500 3686 1501
rect 3482 1470 3530 1500
rect 3638 1470 3686 1500
rect 3482 1469 3485 1470
rect 3447 1468 3485 1469
rect 3683 1469 3686 1470
rect 3718 1500 3721 1501
rect 3895 1501 3933 1502
rect 3895 1500 3898 1501
rect 3718 1470 3765 1500
rect 3851 1470 3898 1500
rect 3718 1469 3721 1470
rect 3683 1468 3721 1469
rect 3895 1469 3898 1470
rect 3930 1500 3933 1501
rect 4131 1501 4169 1502
rect 4131 1500 4134 1501
rect 3930 1470 3978 1500
rect 4086 1470 4134 1500
rect 3930 1469 3933 1470
rect 3895 1468 3933 1469
rect 4131 1469 4134 1470
rect 4166 1500 4169 1501
rect 4343 1501 4381 1502
rect 4343 1500 4346 1501
rect 4166 1470 4213 1500
rect 4299 1470 4346 1500
rect 4166 1469 4169 1470
rect 4131 1468 4169 1469
rect 4343 1469 4346 1470
rect 4378 1500 4381 1501
rect 4579 1501 4617 1502
rect 4579 1500 4582 1501
rect 4378 1470 4426 1500
rect 4534 1470 4582 1500
rect 4378 1469 4381 1470
rect 4343 1468 4381 1469
rect 4579 1469 4582 1470
rect 4614 1500 4617 1501
rect 4791 1501 4829 1502
rect 4791 1500 4794 1501
rect 4614 1470 4661 1500
rect 4747 1470 4794 1500
rect 4614 1469 4617 1470
rect 4579 1468 4617 1469
rect 4791 1469 4794 1470
rect 4826 1500 4829 1501
rect 5027 1501 5065 1502
rect 5027 1500 5030 1501
rect 4826 1470 4874 1500
rect 4982 1470 5030 1500
rect 4826 1469 4829 1470
rect 4791 1468 4829 1469
rect 5027 1469 5030 1470
rect 5062 1500 5065 1501
rect 5239 1501 5277 1502
rect 5239 1500 5242 1501
rect 5062 1470 5109 1500
rect 5195 1470 5242 1500
rect 5062 1469 5065 1470
rect 5027 1468 5065 1469
rect 5239 1469 5242 1470
rect 5274 1500 5277 1501
rect 5475 1501 5513 1502
rect 5475 1500 5478 1501
rect 5274 1470 5322 1500
rect 5430 1470 5478 1500
rect 5274 1469 5277 1470
rect 5239 1468 5277 1469
rect 5475 1469 5478 1470
rect 5510 1500 5513 1501
rect 5687 1501 5725 1502
rect 5687 1500 5690 1501
rect 5510 1470 5557 1500
rect 5643 1470 5690 1500
rect 5510 1469 5513 1470
rect 5475 1468 5513 1469
rect 5687 1469 5690 1470
rect 5722 1500 5725 1501
rect 5923 1501 5961 1502
rect 5923 1500 5926 1501
rect 5722 1470 5770 1500
rect 5878 1470 5926 1500
rect 5722 1469 5725 1470
rect 5687 1468 5725 1469
rect 5923 1469 5926 1470
rect 5958 1500 5961 1501
rect 6135 1501 6173 1502
rect 6135 1500 6138 1501
rect 5958 1470 6005 1500
rect 6091 1470 6138 1500
rect 5958 1469 5961 1470
rect 5923 1468 5961 1469
rect 6135 1469 6138 1470
rect 6170 1500 6173 1501
rect 6371 1501 6409 1502
rect 6371 1500 6374 1501
rect 6170 1470 6218 1500
rect 6326 1470 6374 1500
rect 6170 1469 6173 1470
rect 6135 1468 6173 1469
rect 6371 1469 6374 1470
rect 6406 1500 6409 1501
rect 6583 1501 6621 1502
rect 6583 1500 6586 1501
rect 6406 1470 6453 1500
rect 6539 1470 6586 1500
rect 6406 1469 6409 1470
rect 6371 1468 6409 1469
rect 6583 1469 6586 1470
rect 6618 1500 6621 1501
rect 6819 1501 6857 1502
rect 6819 1500 6822 1501
rect 6618 1470 6666 1500
rect 6774 1470 6822 1500
rect 6618 1469 6621 1470
rect 6583 1468 6621 1469
rect 6819 1469 6822 1470
rect 6854 1500 6857 1501
rect 7031 1501 7069 1502
rect 7031 1500 7034 1501
rect 6854 1470 6901 1500
rect 6987 1470 7034 1500
rect 6854 1469 6857 1470
rect 6819 1468 6857 1469
rect 7031 1469 7034 1470
rect 7066 1500 7069 1501
rect 7267 1501 7305 1502
rect 7267 1500 7270 1501
rect 7066 1470 7114 1500
rect 7222 1470 7270 1500
rect 7066 1469 7069 1470
rect 7031 1468 7069 1469
rect 7267 1469 7270 1470
rect 7302 1500 7305 1501
rect 7479 1501 7517 1502
rect 7479 1500 7482 1501
rect 7302 1470 7349 1500
rect 7435 1470 7482 1500
rect 7302 1469 7305 1470
rect 7267 1468 7305 1469
rect 7479 1469 7482 1470
rect 7514 1500 7517 1501
rect 7715 1501 7753 1502
rect 7715 1500 7718 1501
rect 7514 1470 7562 1500
rect 7670 1470 7718 1500
rect 7514 1469 7517 1470
rect 7479 1468 7517 1469
rect 7715 1469 7718 1470
rect 7750 1500 7753 1501
rect 7927 1501 7965 1502
rect 7927 1500 7930 1501
rect 7750 1470 7797 1500
rect 7883 1470 7930 1500
rect 7750 1469 7753 1470
rect 7715 1468 7753 1469
rect 7927 1469 7930 1470
rect 7962 1500 7965 1501
rect 8163 1501 8201 1502
rect 8163 1500 8166 1501
rect 7962 1470 8010 1500
rect 8118 1470 8166 1500
rect 7962 1469 7965 1470
rect 7927 1468 7965 1469
rect 8163 1469 8166 1470
rect 8198 1500 8201 1501
rect 8375 1501 8413 1502
rect 8375 1500 8378 1501
rect 8198 1470 8245 1500
rect 8331 1470 8378 1500
rect 8198 1469 8201 1470
rect 8163 1468 8201 1469
rect 8375 1469 8378 1470
rect 8410 1500 8413 1501
rect 8611 1501 8649 1502
rect 8611 1500 8614 1501
rect 8410 1470 8458 1500
rect 8566 1470 8614 1500
rect 8410 1469 8413 1470
rect 8375 1468 8413 1469
rect 8611 1469 8614 1470
rect 8646 1500 8649 1501
rect 8823 1501 8861 1502
rect 8823 1500 8826 1501
rect 8646 1470 8693 1500
rect 8779 1470 8826 1500
rect 8646 1469 8649 1470
rect 8611 1468 8649 1469
rect 8823 1469 8826 1470
rect 8858 1500 8861 1501
rect 8858 1470 8906 1500
rect 8858 1469 8861 1470
rect 8823 1468 8861 1469
rect 196 1439 252 1442
rect 196 1438 201 1439
rect 35 1408 201 1438
rect 247 1438 252 1439
rect 644 1439 700 1442
rect 644 1438 649 1439
rect 247 1408 413 1438
rect 483 1408 649 1438
rect 695 1438 700 1439
rect 1092 1439 1148 1442
rect 1092 1438 1097 1439
rect 695 1408 861 1438
rect 931 1408 1097 1438
rect 1143 1438 1148 1439
rect 1540 1439 1596 1442
rect 1540 1438 1545 1439
rect 1143 1408 1309 1438
rect 1379 1408 1545 1438
rect 1591 1438 1596 1439
rect 1988 1439 2044 1442
rect 1988 1438 1993 1439
rect 1591 1408 1757 1438
rect 1827 1408 1993 1438
rect 2039 1438 2044 1439
rect 2436 1439 2492 1442
rect 2436 1438 2441 1439
rect 2039 1408 2205 1438
rect 2275 1408 2441 1438
rect 2487 1438 2492 1439
rect 2884 1439 2940 1442
rect 2884 1438 2889 1439
rect 2487 1408 2653 1438
rect 2723 1408 2889 1438
rect 2935 1438 2940 1439
rect 3332 1439 3388 1442
rect 3332 1438 3337 1439
rect 2935 1408 3101 1438
rect 3171 1408 3337 1438
rect 3383 1438 3388 1439
rect 3780 1439 3836 1442
rect 3780 1438 3785 1439
rect 3383 1408 3549 1438
rect 3619 1408 3785 1438
rect 3831 1438 3836 1439
rect 4228 1439 4284 1442
rect 4228 1438 4233 1439
rect 3831 1408 3997 1438
rect 4067 1408 4233 1438
rect 4279 1438 4284 1439
rect 4676 1439 4732 1442
rect 4676 1438 4681 1439
rect 4279 1408 4445 1438
rect 4515 1408 4681 1438
rect 4727 1438 4732 1439
rect 5124 1439 5180 1442
rect 5124 1438 5129 1439
rect 4727 1408 4893 1438
rect 4963 1408 5129 1438
rect 5175 1438 5180 1439
rect 5572 1439 5628 1442
rect 5572 1438 5577 1439
rect 5175 1408 5341 1438
rect 5411 1408 5577 1438
rect 5623 1438 5628 1439
rect 6020 1439 6076 1442
rect 6020 1438 6025 1439
rect 5623 1408 5789 1438
rect 5859 1408 6025 1438
rect 6071 1438 6076 1439
rect 6468 1439 6524 1442
rect 6468 1438 6473 1439
rect 6071 1408 6237 1438
rect 6307 1408 6473 1438
rect 6519 1438 6524 1439
rect 6916 1439 6972 1442
rect 6916 1438 6921 1439
rect 6519 1408 6685 1438
rect 6755 1408 6921 1438
rect 6967 1438 6972 1439
rect 7364 1439 7420 1442
rect 7364 1438 7369 1439
rect 6967 1408 7133 1438
rect 7203 1408 7369 1438
rect 7415 1438 7420 1439
rect 7812 1439 7868 1442
rect 7812 1438 7817 1439
rect 7415 1408 7581 1438
rect 7651 1408 7817 1438
rect 7863 1438 7868 1439
rect 8260 1439 8316 1442
rect 8260 1438 8265 1439
rect 7863 1408 8029 1438
rect 8099 1408 8265 1438
rect 8311 1438 8316 1439
rect 8708 1439 8764 1442
rect 8708 1438 8713 1439
rect 8311 1408 8477 1438
rect 8547 1408 8713 1438
rect 8759 1438 8764 1439
rect 8759 1408 8925 1438
rect 196 1404 252 1408
rect 644 1404 700 1408
rect 1092 1404 1148 1408
rect 1540 1404 1596 1408
rect 1988 1404 2044 1408
rect 2436 1404 2492 1408
rect 2884 1404 2940 1408
rect 3332 1404 3388 1408
rect 3780 1404 3836 1408
rect 4228 1404 4284 1408
rect 4676 1404 4732 1408
rect 5124 1404 5180 1408
rect 5572 1404 5628 1408
rect 6020 1404 6076 1408
rect 6468 1404 6524 1408
rect 6916 1404 6972 1408
rect 7364 1404 7420 1408
rect 7812 1404 7868 1408
rect 8260 1404 8316 1408
rect 8708 1404 8764 1408
rect 99 1377 137 1378
rect 99 1376 102 1377
rect 54 1346 102 1376
rect 99 1345 102 1346
rect 134 1376 137 1377
rect 311 1377 349 1378
rect 311 1376 314 1377
rect 134 1346 181 1376
rect 267 1346 314 1376
rect 134 1345 137 1346
rect 99 1344 137 1345
rect 311 1345 314 1346
rect 346 1376 349 1377
rect 547 1377 585 1378
rect 547 1376 550 1377
rect 346 1346 394 1376
rect 502 1346 550 1376
rect 346 1345 349 1346
rect 311 1344 349 1345
rect 547 1345 550 1346
rect 582 1376 585 1377
rect 759 1377 797 1378
rect 759 1376 762 1377
rect 582 1346 629 1376
rect 715 1346 762 1376
rect 582 1345 585 1346
rect 547 1344 585 1345
rect 759 1345 762 1346
rect 794 1376 797 1377
rect 995 1377 1033 1378
rect 995 1376 998 1377
rect 794 1346 842 1376
rect 950 1346 998 1376
rect 794 1345 797 1346
rect 759 1344 797 1345
rect 995 1345 998 1346
rect 1030 1376 1033 1377
rect 1207 1377 1245 1378
rect 1207 1376 1210 1377
rect 1030 1346 1077 1376
rect 1163 1346 1210 1376
rect 1030 1345 1033 1346
rect 995 1344 1033 1345
rect 1207 1345 1210 1346
rect 1242 1376 1245 1377
rect 1443 1377 1481 1378
rect 1443 1376 1446 1377
rect 1242 1346 1290 1376
rect 1398 1346 1446 1376
rect 1242 1345 1245 1346
rect 1207 1344 1245 1345
rect 1443 1345 1446 1346
rect 1478 1376 1481 1377
rect 1655 1377 1693 1378
rect 1655 1376 1658 1377
rect 1478 1346 1525 1376
rect 1611 1346 1658 1376
rect 1478 1345 1481 1346
rect 1443 1344 1481 1345
rect 1655 1345 1658 1346
rect 1690 1376 1693 1377
rect 1891 1377 1929 1378
rect 1891 1376 1894 1377
rect 1690 1346 1738 1376
rect 1846 1346 1894 1376
rect 1690 1345 1693 1346
rect 1655 1344 1693 1345
rect 1891 1345 1894 1346
rect 1926 1376 1929 1377
rect 2103 1377 2141 1378
rect 2103 1376 2106 1377
rect 1926 1346 1973 1376
rect 2059 1346 2106 1376
rect 1926 1345 1929 1346
rect 1891 1344 1929 1345
rect 2103 1345 2106 1346
rect 2138 1376 2141 1377
rect 2339 1377 2377 1378
rect 2339 1376 2342 1377
rect 2138 1346 2186 1376
rect 2294 1346 2342 1376
rect 2138 1345 2141 1346
rect 2103 1344 2141 1345
rect 2339 1345 2342 1346
rect 2374 1376 2377 1377
rect 2551 1377 2589 1378
rect 2551 1376 2554 1377
rect 2374 1346 2421 1376
rect 2507 1346 2554 1376
rect 2374 1345 2377 1346
rect 2339 1344 2377 1345
rect 2551 1345 2554 1346
rect 2586 1376 2589 1377
rect 2787 1377 2825 1378
rect 2787 1376 2790 1377
rect 2586 1346 2634 1376
rect 2742 1346 2790 1376
rect 2586 1345 2589 1346
rect 2551 1344 2589 1345
rect 2787 1345 2790 1346
rect 2822 1376 2825 1377
rect 2999 1377 3037 1378
rect 2999 1376 3002 1377
rect 2822 1346 2869 1376
rect 2955 1346 3002 1376
rect 2822 1345 2825 1346
rect 2787 1344 2825 1345
rect 2999 1345 3002 1346
rect 3034 1376 3037 1377
rect 3235 1377 3273 1378
rect 3235 1376 3238 1377
rect 3034 1346 3082 1376
rect 3190 1346 3238 1376
rect 3034 1345 3037 1346
rect 2999 1344 3037 1345
rect 3235 1345 3238 1346
rect 3270 1376 3273 1377
rect 3447 1377 3485 1378
rect 3447 1376 3450 1377
rect 3270 1346 3317 1376
rect 3403 1346 3450 1376
rect 3270 1345 3273 1346
rect 3235 1344 3273 1345
rect 3447 1345 3450 1346
rect 3482 1376 3485 1377
rect 3683 1377 3721 1378
rect 3683 1376 3686 1377
rect 3482 1346 3530 1376
rect 3638 1346 3686 1376
rect 3482 1345 3485 1346
rect 3447 1344 3485 1345
rect 3683 1345 3686 1346
rect 3718 1376 3721 1377
rect 3895 1377 3933 1378
rect 3895 1376 3898 1377
rect 3718 1346 3765 1376
rect 3851 1346 3898 1376
rect 3718 1345 3721 1346
rect 3683 1344 3721 1345
rect 3895 1345 3898 1346
rect 3930 1376 3933 1377
rect 4131 1377 4169 1378
rect 4131 1376 4134 1377
rect 3930 1346 3978 1376
rect 4086 1346 4134 1376
rect 3930 1345 3933 1346
rect 3895 1344 3933 1345
rect 4131 1345 4134 1346
rect 4166 1376 4169 1377
rect 4343 1377 4381 1378
rect 4343 1376 4346 1377
rect 4166 1346 4213 1376
rect 4299 1346 4346 1376
rect 4166 1345 4169 1346
rect 4131 1344 4169 1345
rect 4343 1345 4346 1346
rect 4378 1376 4381 1377
rect 4579 1377 4617 1378
rect 4579 1376 4582 1377
rect 4378 1346 4426 1376
rect 4534 1346 4582 1376
rect 4378 1345 4381 1346
rect 4343 1344 4381 1345
rect 4579 1345 4582 1346
rect 4614 1376 4617 1377
rect 4791 1377 4829 1378
rect 4791 1376 4794 1377
rect 4614 1346 4661 1376
rect 4747 1346 4794 1376
rect 4614 1345 4617 1346
rect 4579 1344 4617 1345
rect 4791 1345 4794 1346
rect 4826 1376 4829 1377
rect 5027 1377 5065 1378
rect 5027 1376 5030 1377
rect 4826 1346 4874 1376
rect 4982 1346 5030 1376
rect 4826 1345 4829 1346
rect 4791 1344 4829 1345
rect 5027 1345 5030 1346
rect 5062 1376 5065 1377
rect 5239 1377 5277 1378
rect 5239 1376 5242 1377
rect 5062 1346 5109 1376
rect 5195 1346 5242 1376
rect 5062 1345 5065 1346
rect 5027 1344 5065 1345
rect 5239 1345 5242 1346
rect 5274 1376 5277 1377
rect 5475 1377 5513 1378
rect 5475 1376 5478 1377
rect 5274 1346 5322 1376
rect 5430 1346 5478 1376
rect 5274 1345 5277 1346
rect 5239 1344 5277 1345
rect 5475 1345 5478 1346
rect 5510 1376 5513 1377
rect 5687 1377 5725 1378
rect 5687 1376 5690 1377
rect 5510 1346 5557 1376
rect 5643 1346 5690 1376
rect 5510 1345 5513 1346
rect 5475 1344 5513 1345
rect 5687 1345 5690 1346
rect 5722 1376 5725 1377
rect 5923 1377 5961 1378
rect 5923 1376 5926 1377
rect 5722 1346 5770 1376
rect 5878 1346 5926 1376
rect 5722 1345 5725 1346
rect 5687 1344 5725 1345
rect 5923 1345 5926 1346
rect 5958 1376 5961 1377
rect 6135 1377 6173 1378
rect 6135 1376 6138 1377
rect 5958 1346 6005 1376
rect 6091 1346 6138 1376
rect 5958 1345 5961 1346
rect 5923 1344 5961 1345
rect 6135 1345 6138 1346
rect 6170 1376 6173 1377
rect 6371 1377 6409 1378
rect 6371 1376 6374 1377
rect 6170 1346 6218 1376
rect 6326 1346 6374 1376
rect 6170 1345 6173 1346
rect 6135 1344 6173 1345
rect 6371 1345 6374 1346
rect 6406 1376 6409 1377
rect 6583 1377 6621 1378
rect 6583 1376 6586 1377
rect 6406 1346 6453 1376
rect 6539 1346 6586 1376
rect 6406 1345 6409 1346
rect 6371 1344 6409 1345
rect 6583 1345 6586 1346
rect 6618 1376 6621 1377
rect 6819 1377 6857 1378
rect 6819 1376 6822 1377
rect 6618 1346 6666 1376
rect 6774 1346 6822 1376
rect 6618 1345 6621 1346
rect 6583 1344 6621 1345
rect 6819 1345 6822 1346
rect 6854 1376 6857 1377
rect 7031 1377 7069 1378
rect 7031 1376 7034 1377
rect 6854 1346 6901 1376
rect 6987 1346 7034 1376
rect 6854 1345 6857 1346
rect 6819 1344 6857 1345
rect 7031 1345 7034 1346
rect 7066 1376 7069 1377
rect 7267 1377 7305 1378
rect 7267 1376 7270 1377
rect 7066 1346 7114 1376
rect 7222 1346 7270 1376
rect 7066 1345 7069 1346
rect 7031 1344 7069 1345
rect 7267 1345 7270 1346
rect 7302 1376 7305 1377
rect 7479 1377 7517 1378
rect 7479 1376 7482 1377
rect 7302 1346 7349 1376
rect 7435 1346 7482 1376
rect 7302 1345 7305 1346
rect 7267 1344 7305 1345
rect 7479 1345 7482 1346
rect 7514 1376 7517 1377
rect 7715 1377 7753 1378
rect 7715 1376 7718 1377
rect 7514 1346 7562 1376
rect 7670 1346 7718 1376
rect 7514 1345 7517 1346
rect 7479 1344 7517 1345
rect 7715 1345 7718 1346
rect 7750 1376 7753 1377
rect 7927 1377 7965 1378
rect 7927 1376 7930 1377
rect 7750 1346 7797 1376
rect 7883 1346 7930 1376
rect 7750 1345 7753 1346
rect 7715 1344 7753 1345
rect 7927 1345 7930 1346
rect 7962 1376 7965 1377
rect 8163 1377 8201 1378
rect 8163 1376 8166 1377
rect 7962 1346 8010 1376
rect 8118 1346 8166 1376
rect 7962 1345 7965 1346
rect 7927 1344 7965 1345
rect 8163 1345 8166 1346
rect 8198 1376 8201 1377
rect 8375 1377 8413 1378
rect 8375 1376 8378 1377
rect 8198 1346 8245 1376
rect 8331 1346 8378 1376
rect 8198 1345 8201 1346
rect 8163 1344 8201 1345
rect 8375 1345 8378 1346
rect 8410 1376 8413 1377
rect 8611 1377 8649 1378
rect 8611 1376 8614 1377
rect 8410 1346 8458 1376
rect 8566 1346 8614 1376
rect 8410 1345 8413 1346
rect 8375 1344 8413 1345
rect 8611 1345 8614 1346
rect 8646 1376 8649 1377
rect 8823 1377 8861 1378
rect 8823 1376 8826 1377
rect 8646 1346 8693 1376
rect 8779 1346 8826 1376
rect 8646 1345 8649 1346
rect 8611 1344 8649 1345
rect 8823 1345 8826 1346
rect 8858 1376 8861 1377
rect 8858 1346 8906 1376
rect 8858 1345 8861 1346
rect 8823 1344 8861 1345
rect 196 1315 252 1318
rect 196 1314 201 1315
rect 35 1284 201 1314
rect 247 1314 252 1315
rect 644 1315 700 1318
rect 644 1314 649 1315
rect 247 1284 413 1314
rect 483 1284 649 1314
rect 695 1314 700 1315
rect 1092 1315 1148 1318
rect 1092 1314 1097 1315
rect 695 1284 861 1314
rect 931 1284 1097 1314
rect 1143 1314 1148 1315
rect 1540 1315 1596 1318
rect 1540 1314 1545 1315
rect 1143 1284 1309 1314
rect 1379 1284 1545 1314
rect 1591 1314 1596 1315
rect 1988 1315 2044 1318
rect 1988 1314 1993 1315
rect 1591 1284 1757 1314
rect 1827 1284 1993 1314
rect 2039 1314 2044 1315
rect 2436 1315 2492 1318
rect 2436 1314 2441 1315
rect 2039 1284 2205 1314
rect 2275 1284 2441 1314
rect 2487 1314 2492 1315
rect 2884 1315 2940 1318
rect 2884 1314 2889 1315
rect 2487 1284 2653 1314
rect 2723 1284 2889 1314
rect 2935 1314 2940 1315
rect 3332 1315 3388 1318
rect 3332 1314 3337 1315
rect 2935 1284 3101 1314
rect 3171 1284 3337 1314
rect 3383 1314 3388 1315
rect 3780 1315 3836 1318
rect 3780 1314 3785 1315
rect 3383 1284 3549 1314
rect 3619 1284 3785 1314
rect 3831 1314 3836 1315
rect 4228 1315 4284 1318
rect 4228 1314 4233 1315
rect 3831 1284 3997 1314
rect 4067 1284 4233 1314
rect 4279 1314 4284 1315
rect 4676 1315 4732 1318
rect 4676 1314 4681 1315
rect 4279 1284 4445 1314
rect 4515 1284 4681 1314
rect 4727 1314 4732 1315
rect 5124 1315 5180 1318
rect 5124 1314 5129 1315
rect 4727 1284 4893 1314
rect 4963 1284 5129 1314
rect 5175 1314 5180 1315
rect 5572 1315 5628 1318
rect 5572 1314 5577 1315
rect 5175 1284 5341 1314
rect 5411 1284 5577 1314
rect 5623 1314 5628 1315
rect 6020 1315 6076 1318
rect 6020 1314 6025 1315
rect 5623 1284 5789 1314
rect 5859 1284 6025 1314
rect 6071 1314 6076 1315
rect 6468 1315 6524 1318
rect 6468 1314 6473 1315
rect 6071 1284 6237 1314
rect 6307 1284 6473 1314
rect 6519 1314 6524 1315
rect 6916 1315 6972 1318
rect 6916 1314 6921 1315
rect 6519 1284 6685 1314
rect 6755 1284 6921 1314
rect 6967 1314 6972 1315
rect 7364 1315 7420 1318
rect 7364 1314 7369 1315
rect 6967 1284 7133 1314
rect 7203 1284 7369 1314
rect 7415 1314 7420 1315
rect 7812 1315 7868 1318
rect 7812 1314 7817 1315
rect 7415 1284 7581 1314
rect 7651 1284 7817 1314
rect 7863 1314 7868 1315
rect 8260 1315 8316 1318
rect 8260 1314 8265 1315
rect 7863 1284 8029 1314
rect 8099 1284 8265 1314
rect 8311 1314 8316 1315
rect 8708 1315 8764 1318
rect 8708 1314 8713 1315
rect 8311 1284 8477 1314
rect 8547 1284 8713 1314
rect 8759 1314 8764 1315
rect 8759 1284 8925 1314
rect 196 1280 252 1284
rect 644 1280 700 1284
rect 1092 1280 1148 1284
rect 1540 1280 1596 1284
rect 1988 1280 2044 1284
rect 2436 1280 2492 1284
rect 2884 1280 2940 1284
rect 3332 1280 3388 1284
rect 3780 1280 3836 1284
rect 4228 1280 4284 1284
rect 4676 1280 4732 1284
rect 5124 1280 5180 1284
rect 5572 1280 5628 1284
rect 6020 1280 6076 1284
rect 6468 1280 6524 1284
rect 6916 1280 6972 1284
rect 7364 1280 7420 1284
rect 7812 1280 7868 1284
rect 8260 1280 8316 1284
rect 8708 1280 8764 1284
rect 196 1193 252 1196
rect 196 1192 201 1193
rect 35 1162 201 1192
rect 247 1192 252 1193
rect 644 1193 700 1196
rect 644 1192 649 1193
rect 247 1162 413 1192
rect 483 1162 649 1192
rect 695 1192 700 1193
rect 1092 1193 1148 1196
rect 1092 1192 1097 1193
rect 695 1162 861 1192
rect 931 1162 1097 1192
rect 1143 1192 1148 1193
rect 1540 1193 1596 1196
rect 1540 1192 1545 1193
rect 1143 1162 1309 1192
rect 1379 1162 1545 1192
rect 1591 1192 1596 1193
rect 1988 1193 2044 1196
rect 1988 1192 1993 1193
rect 1591 1162 1757 1192
rect 1827 1162 1993 1192
rect 2039 1192 2044 1193
rect 2436 1193 2492 1196
rect 2436 1192 2441 1193
rect 2039 1162 2205 1192
rect 2275 1162 2441 1192
rect 2487 1192 2492 1193
rect 2884 1193 2940 1196
rect 2884 1192 2889 1193
rect 2487 1162 2653 1192
rect 2723 1162 2889 1192
rect 2935 1192 2940 1193
rect 3332 1193 3388 1196
rect 3332 1192 3337 1193
rect 2935 1162 3101 1192
rect 3171 1162 3337 1192
rect 3383 1192 3388 1193
rect 3780 1193 3836 1196
rect 3780 1192 3785 1193
rect 3383 1162 3549 1192
rect 3619 1162 3785 1192
rect 3831 1192 3836 1193
rect 4228 1193 4284 1196
rect 4228 1192 4233 1193
rect 3831 1162 3997 1192
rect 4067 1162 4233 1192
rect 4279 1192 4284 1193
rect 4676 1193 4732 1196
rect 4676 1192 4681 1193
rect 4279 1162 4445 1192
rect 4515 1162 4681 1192
rect 4727 1192 4732 1193
rect 5124 1193 5180 1196
rect 5124 1192 5129 1193
rect 4727 1162 4893 1192
rect 4963 1162 5129 1192
rect 5175 1192 5180 1193
rect 5572 1193 5628 1196
rect 5572 1192 5577 1193
rect 5175 1162 5341 1192
rect 5411 1162 5577 1192
rect 5623 1192 5628 1193
rect 6020 1193 6076 1196
rect 6020 1192 6025 1193
rect 5623 1162 5789 1192
rect 5859 1162 6025 1192
rect 6071 1192 6076 1193
rect 6468 1193 6524 1196
rect 6468 1192 6473 1193
rect 6071 1162 6237 1192
rect 6307 1162 6473 1192
rect 6519 1192 6524 1193
rect 6916 1193 6972 1196
rect 6916 1192 6921 1193
rect 6519 1162 6685 1192
rect 6755 1162 6921 1192
rect 6967 1192 6972 1193
rect 7364 1193 7420 1196
rect 7364 1192 7369 1193
rect 6967 1162 7133 1192
rect 7203 1162 7369 1192
rect 7415 1192 7420 1193
rect 7812 1193 7868 1196
rect 7812 1192 7817 1193
rect 7415 1162 7581 1192
rect 7651 1162 7817 1192
rect 7863 1192 7868 1193
rect 8260 1193 8316 1196
rect 8260 1192 8265 1193
rect 7863 1162 8029 1192
rect 8099 1162 8265 1192
rect 8311 1192 8316 1193
rect 8708 1193 8764 1196
rect 8708 1192 8713 1193
rect 8311 1162 8477 1192
rect 8547 1162 8713 1192
rect 8759 1192 8764 1193
rect 8759 1162 8925 1192
rect 196 1158 252 1162
rect 644 1158 700 1162
rect 1092 1158 1148 1162
rect 1540 1158 1596 1162
rect 1988 1158 2044 1162
rect 2436 1158 2492 1162
rect 2884 1158 2940 1162
rect 3332 1158 3388 1162
rect 3780 1158 3836 1162
rect 4228 1158 4284 1162
rect 4676 1158 4732 1162
rect 5124 1158 5180 1162
rect 5572 1158 5628 1162
rect 6020 1158 6076 1162
rect 6468 1158 6524 1162
rect 6916 1158 6972 1162
rect 7364 1158 7420 1162
rect 7812 1158 7868 1162
rect 8260 1158 8316 1162
rect 8708 1158 8764 1162
rect 99 1130 137 1131
rect 99 1129 102 1130
rect 54 1099 102 1129
rect 99 1098 102 1099
rect 134 1129 137 1130
rect 311 1130 349 1131
rect 311 1129 314 1130
rect 134 1099 181 1129
rect 267 1099 314 1129
rect 134 1098 137 1099
rect 99 1097 137 1098
rect 311 1098 314 1099
rect 346 1129 349 1130
rect 547 1130 585 1131
rect 547 1129 550 1130
rect 346 1099 394 1129
rect 502 1099 550 1129
rect 346 1098 349 1099
rect 311 1097 349 1098
rect 547 1098 550 1099
rect 582 1129 585 1130
rect 759 1130 797 1131
rect 759 1129 762 1130
rect 582 1099 629 1129
rect 715 1099 762 1129
rect 582 1098 585 1099
rect 547 1097 585 1098
rect 759 1098 762 1099
rect 794 1129 797 1130
rect 995 1130 1033 1131
rect 995 1129 998 1130
rect 794 1099 842 1129
rect 950 1099 998 1129
rect 794 1098 797 1099
rect 759 1097 797 1098
rect 995 1098 998 1099
rect 1030 1129 1033 1130
rect 1207 1130 1245 1131
rect 1207 1129 1210 1130
rect 1030 1099 1077 1129
rect 1163 1099 1210 1129
rect 1030 1098 1033 1099
rect 995 1097 1033 1098
rect 1207 1098 1210 1099
rect 1242 1129 1245 1130
rect 1443 1130 1481 1131
rect 1443 1129 1446 1130
rect 1242 1099 1290 1129
rect 1398 1099 1446 1129
rect 1242 1098 1245 1099
rect 1207 1097 1245 1098
rect 1443 1098 1446 1099
rect 1478 1129 1481 1130
rect 1655 1130 1693 1131
rect 1655 1129 1658 1130
rect 1478 1099 1525 1129
rect 1611 1099 1658 1129
rect 1478 1098 1481 1099
rect 1443 1097 1481 1098
rect 1655 1098 1658 1099
rect 1690 1129 1693 1130
rect 1891 1130 1929 1131
rect 1891 1129 1894 1130
rect 1690 1099 1738 1129
rect 1846 1099 1894 1129
rect 1690 1098 1693 1099
rect 1655 1097 1693 1098
rect 1891 1098 1894 1099
rect 1926 1129 1929 1130
rect 2103 1130 2141 1131
rect 2103 1129 2106 1130
rect 1926 1099 1973 1129
rect 2059 1099 2106 1129
rect 1926 1098 1929 1099
rect 1891 1097 1929 1098
rect 2103 1098 2106 1099
rect 2138 1129 2141 1130
rect 2339 1130 2377 1131
rect 2339 1129 2342 1130
rect 2138 1099 2186 1129
rect 2294 1099 2342 1129
rect 2138 1098 2141 1099
rect 2103 1097 2141 1098
rect 2339 1098 2342 1099
rect 2374 1129 2377 1130
rect 2551 1130 2589 1131
rect 2551 1129 2554 1130
rect 2374 1099 2421 1129
rect 2507 1099 2554 1129
rect 2374 1098 2377 1099
rect 2339 1097 2377 1098
rect 2551 1098 2554 1099
rect 2586 1129 2589 1130
rect 2787 1130 2825 1131
rect 2787 1129 2790 1130
rect 2586 1099 2634 1129
rect 2742 1099 2790 1129
rect 2586 1098 2589 1099
rect 2551 1097 2589 1098
rect 2787 1098 2790 1099
rect 2822 1129 2825 1130
rect 2999 1130 3037 1131
rect 2999 1129 3002 1130
rect 2822 1099 2869 1129
rect 2955 1099 3002 1129
rect 2822 1098 2825 1099
rect 2787 1097 2825 1098
rect 2999 1098 3002 1099
rect 3034 1129 3037 1130
rect 3235 1130 3273 1131
rect 3235 1129 3238 1130
rect 3034 1099 3082 1129
rect 3190 1099 3238 1129
rect 3034 1098 3037 1099
rect 2999 1097 3037 1098
rect 3235 1098 3238 1099
rect 3270 1129 3273 1130
rect 3447 1130 3485 1131
rect 3447 1129 3450 1130
rect 3270 1099 3317 1129
rect 3403 1099 3450 1129
rect 3270 1098 3273 1099
rect 3235 1097 3273 1098
rect 3447 1098 3450 1099
rect 3482 1129 3485 1130
rect 3683 1130 3721 1131
rect 3683 1129 3686 1130
rect 3482 1099 3530 1129
rect 3638 1099 3686 1129
rect 3482 1098 3485 1099
rect 3447 1097 3485 1098
rect 3683 1098 3686 1099
rect 3718 1129 3721 1130
rect 3895 1130 3933 1131
rect 3895 1129 3898 1130
rect 3718 1099 3765 1129
rect 3851 1099 3898 1129
rect 3718 1098 3721 1099
rect 3683 1097 3721 1098
rect 3895 1098 3898 1099
rect 3930 1129 3933 1130
rect 4131 1130 4169 1131
rect 4131 1129 4134 1130
rect 3930 1099 3978 1129
rect 4086 1099 4134 1129
rect 3930 1098 3933 1099
rect 3895 1097 3933 1098
rect 4131 1098 4134 1099
rect 4166 1129 4169 1130
rect 4343 1130 4381 1131
rect 4343 1129 4346 1130
rect 4166 1099 4213 1129
rect 4299 1099 4346 1129
rect 4166 1098 4169 1099
rect 4131 1097 4169 1098
rect 4343 1098 4346 1099
rect 4378 1129 4381 1130
rect 4579 1130 4617 1131
rect 4579 1129 4582 1130
rect 4378 1099 4426 1129
rect 4534 1099 4582 1129
rect 4378 1098 4381 1099
rect 4343 1097 4381 1098
rect 4579 1098 4582 1099
rect 4614 1129 4617 1130
rect 4791 1130 4829 1131
rect 4791 1129 4794 1130
rect 4614 1099 4661 1129
rect 4747 1099 4794 1129
rect 4614 1098 4617 1099
rect 4579 1097 4617 1098
rect 4791 1098 4794 1099
rect 4826 1129 4829 1130
rect 5027 1130 5065 1131
rect 5027 1129 5030 1130
rect 4826 1099 4874 1129
rect 4982 1099 5030 1129
rect 4826 1098 4829 1099
rect 4791 1097 4829 1098
rect 5027 1098 5030 1099
rect 5062 1129 5065 1130
rect 5239 1130 5277 1131
rect 5239 1129 5242 1130
rect 5062 1099 5109 1129
rect 5195 1099 5242 1129
rect 5062 1098 5065 1099
rect 5027 1097 5065 1098
rect 5239 1098 5242 1099
rect 5274 1129 5277 1130
rect 5475 1130 5513 1131
rect 5475 1129 5478 1130
rect 5274 1099 5322 1129
rect 5430 1099 5478 1129
rect 5274 1098 5277 1099
rect 5239 1097 5277 1098
rect 5475 1098 5478 1099
rect 5510 1129 5513 1130
rect 5687 1130 5725 1131
rect 5687 1129 5690 1130
rect 5510 1099 5557 1129
rect 5643 1099 5690 1129
rect 5510 1098 5513 1099
rect 5475 1097 5513 1098
rect 5687 1098 5690 1099
rect 5722 1129 5725 1130
rect 5923 1130 5961 1131
rect 5923 1129 5926 1130
rect 5722 1099 5770 1129
rect 5878 1099 5926 1129
rect 5722 1098 5725 1099
rect 5687 1097 5725 1098
rect 5923 1098 5926 1099
rect 5958 1129 5961 1130
rect 6135 1130 6173 1131
rect 6135 1129 6138 1130
rect 5958 1099 6005 1129
rect 6091 1099 6138 1129
rect 5958 1098 5961 1099
rect 5923 1097 5961 1098
rect 6135 1098 6138 1099
rect 6170 1129 6173 1130
rect 6371 1130 6409 1131
rect 6371 1129 6374 1130
rect 6170 1099 6218 1129
rect 6326 1099 6374 1129
rect 6170 1098 6173 1099
rect 6135 1097 6173 1098
rect 6371 1098 6374 1099
rect 6406 1129 6409 1130
rect 6583 1130 6621 1131
rect 6583 1129 6586 1130
rect 6406 1099 6453 1129
rect 6539 1099 6586 1129
rect 6406 1098 6409 1099
rect 6371 1097 6409 1098
rect 6583 1098 6586 1099
rect 6618 1129 6621 1130
rect 6819 1130 6857 1131
rect 6819 1129 6822 1130
rect 6618 1099 6666 1129
rect 6774 1099 6822 1129
rect 6618 1098 6621 1099
rect 6583 1097 6621 1098
rect 6819 1098 6822 1099
rect 6854 1129 6857 1130
rect 7031 1130 7069 1131
rect 7031 1129 7034 1130
rect 6854 1099 6901 1129
rect 6987 1099 7034 1129
rect 6854 1098 6857 1099
rect 6819 1097 6857 1098
rect 7031 1098 7034 1099
rect 7066 1129 7069 1130
rect 7267 1130 7305 1131
rect 7267 1129 7270 1130
rect 7066 1099 7114 1129
rect 7222 1099 7270 1129
rect 7066 1098 7069 1099
rect 7031 1097 7069 1098
rect 7267 1098 7270 1099
rect 7302 1129 7305 1130
rect 7479 1130 7517 1131
rect 7479 1129 7482 1130
rect 7302 1099 7349 1129
rect 7435 1099 7482 1129
rect 7302 1098 7305 1099
rect 7267 1097 7305 1098
rect 7479 1098 7482 1099
rect 7514 1129 7517 1130
rect 7715 1130 7753 1131
rect 7715 1129 7718 1130
rect 7514 1099 7562 1129
rect 7670 1099 7718 1129
rect 7514 1098 7517 1099
rect 7479 1097 7517 1098
rect 7715 1098 7718 1099
rect 7750 1129 7753 1130
rect 7927 1130 7965 1131
rect 7927 1129 7930 1130
rect 7750 1099 7797 1129
rect 7883 1099 7930 1129
rect 7750 1098 7753 1099
rect 7715 1097 7753 1098
rect 7927 1098 7930 1099
rect 7962 1129 7965 1130
rect 8163 1130 8201 1131
rect 8163 1129 8166 1130
rect 7962 1099 8010 1129
rect 8118 1099 8166 1129
rect 7962 1098 7965 1099
rect 7927 1097 7965 1098
rect 8163 1098 8166 1099
rect 8198 1129 8201 1130
rect 8375 1130 8413 1131
rect 8375 1129 8378 1130
rect 8198 1099 8245 1129
rect 8331 1099 8378 1129
rect 8198 1098 8201 1099
rect 8163 1097 8201 1098
rect 8375 1098 8378 1099
rect 8410 1129 8413 1130
rect 8611 1130 8649 1131
rect 8611 1129 8614 1130
rect 8410 1099 8458 1129
rect 8566 1099 8614 1129
rect 8410 1098 8413 1099
rect 8375 1097 8413 1098
rect 8611 1098 8614 1099
rect 8646 1129 8649 1130
rect 8823 1130 8861 1131
rect 8823 1129 8826 1130
rect 8646 1099 8693 1129
rect 8779 1099 8826 1129
rect 8646 1098 8649 1099
rect 8611 1097 8649 1098
rect 8823 1098 8826 1099
rect 8858 1129 8861 1130
rect 8858 1099 8906 1129
rect 8858 1098 8861 1099
rect 8823 1097 8861 1098
rect 196 1068 252 1071
rect 196 1067 201 1068
rect 35 1037 201 1067
rect 247 1067 252 1068
rect 644 1068 700 1071
rect 644 1067 649 1068
rect 247 1037 413 1067
rect 483 1037 649 1067
rect 695 1067 700 1068
rect 1092 1068 1148 1071
rect 1092 1067 1097 1068
rect 695 1037 861 1067
rect 931 1037 1097 1067
rect 1143 1067 1148 1068
rect 1540 1068 1596 1071
rect 1540 1067 1545 1068
rect 1143 1037 1309 1067
rect 1379 1037 1545 1067
rect 1591 1067 1596 1068
rect 1988 1068 2044 1071
rect 1988 1067 1993 1068
rect 1591 1037 1757 1067
rect 1827 1037 1993 1067
rect 2039 1067 2044 1068
rect 2436 1068 2492 1071
rect 2436 1067 2441 1068
rect 2039 1037 2205 1067
rect 2275 1037 2441 1067
rect 2487 1067 2492 1068
rect 2884 1068 2940 1071
rect 2884 1067 2889 1068
rect 2487 1037 2653 1067
rect 2723 1037 2889 1067
rect 2935 1067 2940 1068
rect 3332 1068 3388 1071
rect 3332 1067 3337 1068
rect 2935 1037 3101 1067
rect 3171 1037 3337 1067
rect 3383 1067 3388 1068
rect 3780 1068 3836 1071
rect 3780 1067 3785 1068
rect 3383 1037 3549 1067
rect 3619 1037 3785 1067
rect 3831 1067 3836 1068
rect 4228 1068 4284 1071
rect 4228 1067 4233 1068
rect 3831 1037 3997 1067
rect 4067 1037 4233 1067
rect 4279 1067 4284 1068
rect 4676 1068 4732 1071
rect 4676 1067 4681 1068
rect 4279 1037 4445 1067
rect 4515 1037 4681 1067
rect 4727 1067 4732 1068
rect 5124 1068 5180 1071
rect 5124 1067 5129 1068
rect 4727 1037 4893 1067
rect 4963 1037 5129 1067
rect 5175 1067 5180 1068
rect 5572 1068 5628 1071
rect 5572 1067 5577 1068
rect 5175 1037 5341 1067
rect 5411 1037 5577 1067
rect 5623 1067 5628 1068
rect 6020 1068 6076 1071
rect 6020 1067 6025 1068
rect 5623 1037 5789 1067
rect 5859 1037 6025 1067
rect 6071 1067 6076 1068
rect 6468 1068 6524 1071
rect 6468 1067 6473 1068
rect 6071 1037 6237 1067
rect 6307 1037 6473 1067
rect 6519 1067 6524 1068
rect 6916 1068 6972 1071
rect 6916 1067 6921 1068
rect 6519 1037 6685 1067
rect 6755 1037 6921 1067
rect 6967 1067 6972 1068
rect 7364 1068 7420 1071
rect 7364 1067 7369 1068
rect 6967 1037 7133 1067
rect 7203 1037 7369 1067
rect 7415 1067 7420 1068
rect 7812 1068 7868 1071
rect 7812 1067 7817 1068
rect 7415 1037 7581 1067
rect 7651 1037 7817 1067
rect 7863 1067 7868 1068
rect 8260 1068 8316 1071
rect 8260 1067 8265 1068
rect 7863 1037 8029 1067
rect 8099 1037 8265 1067
rect 8311 1067 8316 1068
rect 8708 1068 8764 1071
rect 8708 1067 8713 1068
rect 8311 1037 8477 1067
rect 8547 1037 8713 1067
rect 8759 1067 8764 1068
rect 8759 1037 8925 1067
rect 196 1033 252 1037
rect 644 1033 700 1037
rect 1092 1033 1148 1037
rect 1540 1033 1596 1037
rect 1988 1033 2044 1037
rect 2436 1033 2492 1037
rect 2884 1033 2940 1037
rect 3332 1033 3388 1037
rect 3780 1033 3836 1037
rect 4228 1033 4284 1037
rect 4676 1033 4732 1037
rect 5124 1033 5180 1037
rect 5572 1033 5628 1037
rect 6020 1033 6076 1037
rect 6468 1033 6524 1037
rect 6916 1033 6972 1037
rect 7364 1033 7420 1037
rect 7812 1033 7868 1037
rect 8260 1033 8316 1037
rect 8708 1033 8764 1037
rect 99 1006 137 1007
rect 99 1005 102 1006
rect 54 975 102 1005
rect 99 974 102 975
rect 134 1005 137 1006
rect 311 1006 349 1007
rect 311 1005 314 1006
rect 134 975 181 1005
rect 267 975 314 1005
rect 134 974 137 975
rect 99 973 137 974
rect 311 974 314 975
rect 346 1005 349 1006
rect 547 1006 585 1007
rect 547 1005 550 1006
rect 346 975 394 1005
rect 502 975 550 1005
rect 346 974 349 975
rect 311 973 349 974
rect 547 974 550 975
rect 582 1005 585 1006
rect 759 1006 797 1007
rect 759 1005 762 1006
rect 582 975 629 1005
rect 715 975 762 1005
rect 582 974 585 975
rect 547 973 585 974
rect 759 974 762 975
rect 794 1005 797 1006
rect 995 1006 1033 1007
rect 995 1005 998 1006
rect 794 975 842 1005
rect 950 975 998 1005
rect 794 974 797 975
rect 759 973 797 974
rect 995 974 998 975
rect 1030 1005 1033 1006
rect 1207 1006 1245 1007
rect 1207 1005 1210 1006
rect 1030 975 1077 1005
rect 1163 975 1210 1005
rect 1030 974 1033 975
rect 995 973 1033 974
rect 1207 974 1210 975
rect 1242 1005 1245 1006
rect 1443 1006 1481 1007
rect 1443 1005 1446 1006
rect 1242 975 1290 1005
rect 1398 975 1446 1005
rect 1242 974 1245 975
rect 1207 973 1245 974
rect 1443 974 1446 975
rect 1478 1005 1481 1006
rect 1655 1006 1693 1007
rect 1655 1005 1658 1006
rect 1478 975 1525 1005
rect 1611 975 1658 1005
rect 1478 974 1481 975
rect 1443 973 1481 974
rect 1655 974 1658 975
rect 1690 1005 1693 1006
rect 1891 1006 1929 1007
rect 1891 1005 1894 1006
rect 1690 975 1738 1005
rect 1846 975 1894 1005
rect 1690 974 1693 975
rect 1655 973 1693 974
rect 1891 974 1894 975
rect 1926 1005 1929 1006
rect 2103 1006 2141 1007
rect 2103 1005 2106 1006
rect 1926 975 1973 1005
rect 2059 975 2106 1005
rect 1926 974 1929 975
rect 1891 973 1929 974
rect 2103 974 2106 975
rect 2138 1005 2141 1006
rect 2339 1006 2377 1007
rect 2339 1005 2342 1006
rect 2138 975 2186 1005
rect 2294 975 2342 1005
rect 2138 974 2141 975
rect 2103 973 2141 974
rect 2339 974 2342 975
rect 2374 1005 2377 1006
rect 2551 1006 2589 1007
rect 2551 1005 2554 1006
rect 2374 975 2421 1005
rect 2507 975 2554 1005
rect 2374 974 2377 975
rect 2339 973 2377 974
rect 2551 974 2554 975
rect 2586 1005 2589 1006
rect 2787 1006 2825 1007
rect 2787 1005 2790 1006
rect 2586 975 2634 1005
rect 2742 975 2790 1005
rect 2586 974 2589 975
rect 2551 973 2589 974
rect 2787 974 2790 975
rect 2822 1005 2825 1006
rect 2999 1006 3037 1007
rect 2999 1005 3002 1006
rect 2822 975 2869 1005
rect 2955 975 3002 1005
rect 2822 974 2825 975
rect 2787 973 2825 974
rect 2999 974 3002 975
rect 3034 1005 3037 1006
rect 3235 1006 3273 1007
rect 3235 1005 3238 1006
rect 3034 975 3082 1005
rect 3190 975 3238 1005
rect 3034 974 3037 975
rect 2999 973 3037 974
rect 3235 974 3238 975
rect 3270 1005 3273 1006
rect 3447 1006 3485 1007
rect 3447 1005 3450 1006
rect 3270 975 3317 1005
rect 3403 975 3450 1005
rect 3270 974 3273 975
rect 3235 973 3273 974
rect 3447 974 3450 975
rect 3482 1005 3485 1006
rect 3683 1006 3721 1007
rect 3683 1005 3686 1006
rect 3482 975 3530 1005
rect 3638 975 3686 1005
rect 3482 974 3485 975
rect 3447 973 3485 974
rect 3683 974 3686 975
rect 3718 1005 3721 1006
rect 3895 1006 3933 1007
rect 3895 1005 3898 1006
rect 3718 975 3765 1005
rect 3851 975 3898 1005
rect 3718 974 3721 975
rect 3683 973 3721 974
rect 3895 974 3898 975
rect 3930 1005 3933 1006
rect 4131 1006 4169 1007
rect 4131 1005 4134 1006
rect 3930 975 3978 1005
rect 4086 975 4134 1005
rect 3930 974 3933 975
rect 3895 973 3933 974
rect 4131 974 4134 975
rect 4166 1005 4169 1006
rect 4343 1006 4381 1007
rect 4343 1005 4346 1006
rect 4166 975 4213 1005
rect 4299 975 4346 1005
rect 4166 974 4169 975
rect 4131 973 4169 974
rect 4343 974 4346 975
rect 4378 1005 4381 1006
rect 4579 1006 4617 1007
rect 4579 1005 4582 1006
rect 4378 975 4426 1005
rect 4534 975 4582 1005
rect 4378 974 4381 975
rect 4343 973 4381 974
rect 4579 974 4582 975
rect 4614 1005 4617 1006
rect 4791 1006 4829 1007
rect 4791 1005 4794 1006
rect 4614 975 4661 1005
rect 4747 975 4794 1005
rect 4614 974 4617 975
rect 4579 973 4617 974
rect 4791 974 4794 975
rect 4826 1005 4829 1006
rect 5027 1006 5065 1007
rect 5027 1005 5030 1006
rect 4826 975 4874 1005
rect 4982 975 5030 1005
rect 4826 974 4829 975
rect 4791 973 4829 974
rect 5027 974 5030 975
rect 5062 1005 5065 1006
rect 5239 1006 5277 1007
rect 5239 1005 5242 1006
rect 5062 975 5109 1005
rect 5195 975 5242 1005
rect 5062 974 5065 975
rect 5027 973 5065 974
rect 5239 974 5242 975
rect 5274 1005 5277 1006
rect 5475 1006 5513 1007
rect 5475 1005 5478 1006
rect 5274 975 5322 1005
rect 5430 975 5478 1005
rect 5274 974 5277 975
rect 5239 973 5277 974
rect 5475 974 5478 975
rect 5510 1005 5513 1006
rect 5687 1006 5725 1007
rect 5687 1005 5690 1006
rect 5510 975 5557 1005
rect 5643 975 5690 1005
rect 5510 974 5513 975
rect 5475 973 5513 974
rect 5687 974 5690 975
rect 5722 1005 5725 1006
rect 5923 1006 5961 1007
rect 5923 1005 5926 1006
rect 5722 975 5770 1005
rect 5878 975 5926 1005
rect 5722 974 5725 975
rect 5687 973 5725 974
rect 5923 974 5926 975
rect 5958 1005 5961 1006
rect 6135 1006 6173 1007
rect 6135 1005 6138 1006
rect 5958 975 6005 1005
rect 6091 975 6138 1005
rect 5958 974 5961 975
rect 5923 973 5961 974
rect 6135 974 6138 975
rect 6170 1005 6173 1006
rect 6371 1006 6409 1007
rect 6371 1005 6374 1006
rect 6170 975 6218 1005
rect 6326 975 6374 1005
rect 6170 974 6173 975
rect 6135 973 6173 974
rect 6371 974 6374 975
rect 6406 1005 6409 1006
rect 6583 1006 6621 1007
rect 6583 1005 6586 1006
rect 6406 975 6453 1005
rect 6539 975 6586 1005
rect 6406 974 6409 975
rect 6371 973 6409 974
rect 6583 974 6586 975
rect 6618 1005 6621 1006
rect 6819 1006 6857 1007
rect 6819 1005 6822 1006
rect 6618 975 6666 1005
rect 6774 975 6822 1005
rect 6618 974 6621 975
rect 6583 973 6621 974
rect 6819 974 6822 975
rect 6854 1005 6857 1006
rect 7031 1006 7069 1007
rect 7031 1005 7034 1006
rect 6854 975 6901 1005
rect 6987 975 7034 1005
rect 6854 974 6857 975
rect 6819 973 6857 974
rect 7031 974 7034 975
rect 7066 1005 7069 1006
rect 7267 1006 7305 1007
rect 7267 1005 7270 1006
rect 7066 975 7114 1005
rect 7222 975 7270 1005
rect 7066 974 7069 975
rect 7031 973 7069 974
rect 7267 974 7270 975
rect 7302 1005 7305 1006
rect 7479 1006 7517 1007
rect 7479 1005 7482 1006
rect 7302 975 7349 1005
rect 7435 975 7482 1005
rect 7302 974 7305 975
rect 7267 973 7305 974
rect 7479 974 7482 975
rect 7514 1005 7517 1006
rect 7715 1006 7753 1007
rect 7715 1005 7718 1006
rect 7514 975 7562 1005
rect 7670 975 7718 1005
rect 7514 974 7517 975
rect 7479 973 7517 974
rect 7715 974 7718 975
rect 7750 1005 7753 1006
rect 7927 1006 7965 1007
rect 7927 1005 7930 1006
rect 7750 975 7797 1005
rect 7883 975 7930 1005
rect 7750 974 7753 975
rect 7715 973 7753 974
rect 7927 974 7930 975
rect 7962 1005 7965 1006
rect 8163 1006 8201 1007
rect 8163 1005 8166 1006
rect 7962 975 8010 1005
rect 8118 975 8166 1005
rect 7962 974 7965 975
rect 7927 973 7965 974
rect 8163 974 8166 975
rect 8198 1005 8201 1006
rect 8375 1006 8413 1007
rect 8375 1005 8378 1006
rect 8198 975 8245 1005
rect 8331 975 8378 1005
rect 8198 974 8201 975
rect 8163 973 8201 974
rect 8375 974 8378 975
rect 8410 1005 8413 1006
rect 8611 1006 8649 1007
rect 8611 1005 8614 1006
rect 8410 975 8458 1005
rect 8566 975 8614 1005
rect 8410 974 8413 975
rect 8375 973 8413 974
rect 8611 974 8614 975
rect 8646 1005 8649 1006
rect 8823 1006 8861 1007
rect 8823 1005 8826 1006
rect 8646 975 8693 1005
rect 8779 975 8826 1005
rect 8646 974 8649 975
rect 8611 973 8649 974
rect 8823 974 8826 975
rect 8858 1005 8861 1006
rect 8858 975 8906 1005
rect 8858 974 8861 975
rect 8823 973 8861 974
rect 196 944 252 947
rect 196 943 201 944
rect 35 913 201 943
rect 247 943 252 944
rect 644 944 700 947
rect 644 943 649 944
rect 247 913 413 943
rect 483 913 649 943
rect 695 943 700 944
rect 1092 944 1148 947
rect 1092 943 1097 944
rect 695 913 861 943
rect 931 913 1097 943
rect 1143 943 1148 944
rect 1540 944 1596 947
rect 1540 943 1545 944
rect 1143 913 1309 943
rect 1379 913 1545 943
rect 1591 943 1596 944
rect 1988 944 2044 947
rect 1988 943 1993 944
rect 1591 913 1757 943
rect 1827 913 1993 943
rect 2039 943 2044 944
rect 2436 944 2492 947
rect 2436 943 2441 944
rect 2039 913 2205 943
rect 2275 913 2441 943
rect 2487 943 2492 944
rect 2884 944 2940 947
rect 2884 943 2889 944
rect 2487 913 2653 943
rect 2723 913 2889 943
rect 2935 943 2940 944
rect 3332 944 3388 947
rect 3332 943 3337 944
rect 2935 913 3101 943
rect 3171 913 3337 943
rect 3383 943 3388 944
rect 3780 944 3836 947
rect 3780 943 3785 944
rect 3383 913 3549 943
rect 3619 913 3785 943
rect 3831 943 3836 944
rect 4228 944 4284 947
rect 4228 943 4233 944
rect 3831 913 3997 943
rect 4067 913 4233 943
rect 4279 943 4284 944
rect 4676 944 4732 947
rect 4676 943 4681 944
rect 4279 913 4445 943
rect 4515 913 4681 943
rect 4727 943 4732 944
rect 5124 944 5180 947
rect 5124 943 5129 944
rect 4727 913 4893 943
rect 4963 913 5129 943
rect 5175 943 5180 944
rect 5572 944 5628 947
rect 5572 943 5577 944
rect 5175 913 5341 943
rect 5411 913 5577 943
rect 5623 943 5628 944
rect 6020 944 6076 947
rect 6020 943 6025 944
rect 5623 913 5789 943
rect 5859 913 6025 943
rect 6071 943 6076 944
rect 6468 944 6524 947
rect 6468 943 6473 944
rect 6071 913 6237 943
rect 6307 913 6473 943
rect 6519 943 6524 944
rect 6916 944 6972 947
rect 6916 943 6921 944
rect 6519 913 6685 943
rect 6755 913 6921 943
rect 6967 943 6972 944
rect 7364 944 7420 947
rect 7364 943 7369 944
rect 6967 913 7133 943
rect 7203 913 7369 943
rect 7415 943 7420 944
rect 7812 944 7868 947
rect 7812 943 7817 944
rect 7415 913 7581 943
rect 7651 913 7817 943
rect 7863 943 7868 944
rect 8260 944 8316 947
rect 8260 943 8265 944
rect 7863 913 8029 943
rect 8099 913 8265 943
rect 8311 943 8316 944
rect 8708 944 8764 947
rect 8708 943 8713 944
rect 8311 913 8477 943
rect 8547 913 8713 943
rect 8759 943 8764 944
rect 8759 913 8925 943
rect 196 909 252 913
rect 644 909 700 913
rect 1092 909 1148 913
rect 1540 909 1596 913
rect 1988 909 2044 913
rect 2436 909 2492 913
rect 2884 909 2940 913
rect 3332 909 3388 913
rect 3780 909 3836 913
rect 4228 909 4284 913
rect 4676 909 4732 913
rect 5124 909 5180 913
rect 5572 909 5628 913
rect 6020 909 6076 913
rect 6468 909 6524 913
rect 6916 909 6972 913
rect 7364 909 7420 913
rect 7812 909 7868 913
rect 8260 909 8316 913
rect 8708 909 8764 913
rect 99 882 137 883
rect 99 881 102 882
rect 54 851 102 881
rect 99 850 102 851
rect 134 881 137 882
rect 311 882 349 883
rect 311 881 314 882
rect 134 851 181 881
rect 267 851 314 881
rect 134 850 137 851
rect 99 849 137 850
rect 311 850 314 851
rect 346 881 349 882
rect 547 882 585 883
rect 547 881 550 882
rect 346 851 394 881
rect 502 851 550 881
rect 346 850 349 851
rect 311 849 349 850
rect 547 850 550 851
rect 582 881 585 882
rect 759 882 797 883
rect 759 881 762 882
rect 582 851 629 881
rect 715 851 762 881
rect 582 850 585 851
rect 547 849 585 850
rect 759 850 762 851
rect 794 881 797 882
rect 995 882 1033 883
rect 995 881 998 882
rect 794 851 842 881
rect 950 851 998 881
rect 794 850 797 851
rect 759 849 797 850
rect 995 850 998 851
rect 1030 881 1033 882
rect 1207 882 1245 883
rect 1207 881 1210 882
rect 1030 851 1077 881
rect 1163 851 1210 881
rect 1030 850 1033 851
rect 995 849 1033 850
rect 1207 850 1210 851
rect 1242 881 1245 882
rect 1443 882 1481 883
rect 1443 881 1446 882
rect 1242 851 1290 881
rect 1398 851 1446 881
rect 1242 850 1245 851
rect 1207 849 1245 850
rect 1443 850 1446 851
rect 1478 881 1481 882
rect 1655 882 1693 883
rect 1655 881 1658 882
rect 1478 851 1525 881
rect 1611 851 1658 881
rect 1478 850 1481 851
rect 1443 849 1481 850
rect 1655 850 1658 851
rect 1690 881 1693 882
rect 1891 882 1929 883
rect 1891 881 1894 882
rect 1690 851 1738 881
rect 1846 851 1894 881
rect 1690 850 1693 851
rect 1655 849 1693 850
rect 1891 850 1894 851
rect 1926 881 1929 882
rect 2103 882 2141 883
rect 2103 881 2106 882
rect 1926 851 1973 881
rect 2059 851 2106 881
rect 1926 850 1929 851
rect 1891 849 1929 850
rect 2103 850 2106 851
rect 2138 881 2141 882
rect 2339 882 2377 883
rect 2339 881 2342 882
rect 2138 851 2186 881
rect 2294 851 2342 881
rect 2138 850 2141 851
rect 2103 849 2141 850
rect 2339 850 2342 851
rect 2374 881 2377 882
rect 2551 882 2589 883
rect 2551 881 2554 882
rect 2374 851 2421 881
rect 2507 851 2554 881
rect 2374 850 2377 851
rect 2339 849 2377 850
rect 2551 850 2554 851
rect 2586 881 2589 882
rect 2787 882 2825 883
rect 2787 881 2790 882
rect 2586 851 2634 881
rect 2742 851 2790 881
rect 2586 850 2589 851
rect 2551 849 2589 850
rect 2787 850 2790 851
rect 2822 881 2825 882
rect 2999 882 3037 883
rect 2999 881 3002 882
rect 2822 851 2869 881
rect 2955 851 3002 881
rect 2822 850 2825 851
rect 2787 849 2825 850
rect 2999 850 3002 851
rect 3034 881 3037 882
rect 3235 882 3273 883
rect 3235 881 3238 882
rect 3034 851 3082 881
rect 3190 851 3238 881
rect 3034 850 3037 851
rect 2999 849 3037 850
rect 3235 850 3238 851
rect 3270 881 3273 882
rect 3447 882 3485 883
rect 3447 881 3450 882
rect 3270 851 3317 881
rect 3403 851 3450 881
rect 3270 850 3273 851
rect 3235 849 3273 850
rect 3447 850 3450 851
rect 3482 881 3485 882
rect 3683 882 3721 883
rect 3683 881 3686 882
rect 3482 851 3530 881
rect 3638 851 3686 881
rect 3482 850 3485 851
rect 3447 849 3485 850
rect 3683 850 3686 851
rect 3718 881 3721 882
rect 3895 882 3933 883
rect 3895 881 3898 882
rect 3718 851 3765 881
rect 3851 851 3898 881
rect 3718 850 3721 851
rect 3683 849 3721 850
rect 3895 850 3898 851
rect 3930 881 3933 882
rect 4131 882 4169 883
rect 4131 881 4134 882
rect 3930 851 3978 881
rect 4086 851 4134 881
rect 3930 850 3933 851
rect 3895 849 3933 850
rect 4131 850 4134 851
rect 4166 881 4169 882
rect 4343 882 4381 883
rect 4343 881 4346 882
rect 4166 851 4213 881
rect 4299 851 4346 881
rect 4166 850 4169 851
rect 4131 849 4169 850
rect 4343 850 4346 851
rect 4378 881 4381 882
rect 4579 882 4617 883
rect 4579 881 4582 882
rect 4378 851 4426 881
rect 4534 851 4582 881
rect 4378 850 4381 851
rect 4343 849 4381 850
rect 4579 850 4582 851
rect 4614 881 4617 882
rect 4791 882 4829 883
rect 4791 881 4794 882
rect 4614 851 4661 881
rect 4747 851 4794 881
rect 4614 850 4617 851
rect 4579 849 4617 850
rect 4791 850 4794 851
rect 4826 881 4829 882
rect 5027 882 5065 883
rect 5027 881 5030 882
rect 4826 851 4874 881
rect 4982 851 5030 881
rect 4826 850 4829 851
rect 4791 849 4829 850
rect 5027 850 5030 851
rect 5062 881 5065 882
rect 5239 882 5277 883
rect 5239 881 5242 882
rect 5062 851 5109 881
rect 5195 851 5242 881
rect 5062 850 5065 851
rect 5027 849 5065 850
rect 5239 850 5242 851
rect 5274 881 5277 882
rect 5475 882 5513 883
rect 5475 881 5478 882
rect 5274 851 5322 881
rect 5430 851 5478 881
rect 5274 850 5277 851
rect 5239 849 5277 850
rect 5475 850 5478 851
rect 5510 881 5513 882
rect 5687 882 5725 883
rect 5687 881 5690 882
rect 5510 851 5557 881
rect 5643 851 5690 881
rect 5510 850 5513 851
rect 5475 849 5513 850
rect 5687 850 5690 851
rect 5722 881 5725 882
rect 5923 882 5961 883
rect 5923 881 5926 882
rect 5722 851 5770 881
rect 5878 851 5926 881
rect 5722 850 5725 851
rect 5687 849 5725 850
rect 5923 850 5926 851
rect 5958 881 5961 882
rect 6135 882 6173 883
rect 6135 881 6138 882
rect 5958 851 6005 881
rect 6091 851 6138 881
rect 5958 850 5961 851
rect 5923 849 5961 850
rect 6135 850 6138 851
rect 6170 881 6173 882
rect 6371 882 6409 883
rect 6371 881 6374 882
rect 6170 851 6218 881
rect 6326 851 6374 881
rect 6170 850 6173 851
rect 6135 849 6173 850
rect 6371 850 6374 851
rect 6406 881 6409 882
rect 6583 882 6621 883
rect 6583 881 6586 882
rect 6406 851 6453 881
rect 6539 851 6586 881
rect 6406 850 6409 851
rect 6371 849 6409 850
rect 6583 850 6586 851
rect 6618 881 6621 882
rect 6819 882 6857 883
rect 6819 881 6822 882
rect 6618 851 6666 881
rect 6774 851 6822 881
rect 6618 850 6621 851
rect 6583 849 6621 850
rect 6819 850 6822 851
rect 6854 881 6857 882
rect 7031 882 7069 883
rect 7031 881 7034 882
rect 6854 851 6901 881
rect 6987 851 7034 881
rect 6854 850 6857 851
rect 6819 849 6857 850
rect 7031 850 7034 851
rect 7066 881 7069 882
rect 7267 882 7305 883
rect 7267 881 7270 882
rect 7066 851 7114 881
rect 7222 851 7270 881
rect 7066 850 7069 851
rect 7031 849 7069 850
rect 7267 850 7270 851
rect 7302 881 7305 882
rect 7479 882 7517 883
rect 7479 881 7482 882
rect 7302 851 7349 881
rect 7435 851 7482 881
rect 7302 850 7305 851
rect 7267 849 7305 850
rect 7479 850 7482 851
rect 7514 881 7517 882
rect 7715 882 7753 883
rect 7715 881 7718 882
rect 7514 851 7562 881
rect 7670 851 7718 881
rect 7514 850 7517 851
rect 7479 849 7517 850
rect 7715 850 7718 851
rect 7750 881 7753 882
rect 7927 882 7965 883
rect 7927 881 7930 882
rect 7750 851 7797 881
rect 7883 851 7930 881
rect 7750 850 7753 851
rect 7715 849 7753 850
rect 7927 850 7930 851
rect 7962 881 7965 882
rect 8163 882 8201 883
rect 8163 881 8166 882
rect 7962 851 8010 881
rect 8118 851 8166 881
rect 7962 850 7965 851
rect 7927 849 7965 850
rect 8163 850 8166 851
rect 8198 881 8201 882
rect 8375 882 8413 883
rect 8375 881 8378 882
rect 8198 851 8245 881
rect 8331 851 8378 881
rect 8198 850 8201 851
rect 8163 849 8201 850
rect 8375 850 8378 851
rect 8410 881 8413 882
rect 8611 882 8649 883
rect 8611 881 8614 882
rect 8410 851 8458 881
rect 8566 851 8614 881
rect 8410 850 8413 851
rect 8375 849 8413 850
rect 8611 850 8614 851
rect 8646 881 8649 882
rect 8823 882 8861 883
rect 8823 881 8826 882
rect 8646 851 8693 881
rect 8779 851 8826 881
rect 8646 850 8649 851
rect 8611 849 8649 850
rect 8823 850 8826 851
rect 8858 881 8861 882
rect 8858 851 8906 881
rect 8858 850 8861 851
rect 8823 849 8861 850
rect 196 820 252 823
rect 196 819 201 820
rect 35 789 201 819
rect 247 819 252 820
rect 644 820 700 823
rect 644 819 649 820
rect 247 789 413 819
rect 483 789 649 819
rect 695 819 700 820
rect 1092 820 1148 823
rect 1092 819 1097 820
rect 695 789 861 819
rect 931 789 1097 819
rect 1143 819 1148 820
rect 1540 820 1596 823
rect 1540 819 1545 820
rect 1143 789 1309 819
rect 1379 789 1545 819
rect 1591 819 1596 820
rect 1988 820 2044 823
rect 1988 819 1993 820
rect 1591 789 1757 819
rect 1827 789 1993 819
rect 2039 819 2044 820
rect 2436 820 2492 823
rect 2436 819 2441 820
rect 2039 789 2205 819
rect 2275 789 2441 819
rect 2487 819 2492 820
rect 2884 820 2940 823
rect 2884 819 2889 820
rect 2487 789 2653 819
rect 2723 789 2889 819
rect 2935 819 2940 820
rect 3332 820 3388 823
rect 3332 819 3337 820
rect 2935 789 3101 819
rect 3171 789 3337 819
rect 3383 819 3388 820
rect 3780 820 3836 823
rect 3780 819 3785 820
rect 3383 789 3549 819
rect 3619 789 3785 819
rect 3831 819 3836 820
rect 4228 820 4284 823
rect 4228 819 4233 820
rect 3831 789 3997 819
rect 4067 789 4233 819
rect 4279 819 4284 820
rect 4676 820 4732 823
rect 4676 819 4681 820
rect 4279 789 4445 819
rect 4515 789 4681 819
rect 4727 819 4732 820
rect 5124 820 5180 823
rect 5124 819 5129 820
rect 4727 789 4893 819
rect 4963 789 5129 819
rect 5175 819 5180 820
rect 5572 820 5628 823
rect 5572 819 5577 820
rect 5175 789 5341 819
rect 5411 789 5577 819
rect 5623 819 5628 820
rect 6020 820 6076 823
rect 6020 819 6025 820
rect 5623 789 5789 819
rect 5859 789 6025 819
rect 6071 819 6076 820
rect 6468 820 6524 823
rect 6468 819 6473 820
rect 6071 789 6237 819
rect 6307 789 6473 819
rect 6519 819 6524 820
rect 6916 820 6972 823
rect 6916 819 6921 820
rect 6519 789 6685 819
rect 6755 789 6921 819
rect 6967 819 6972 820
rect 7364 820 7420 823
rect 7364 819 7369 820
rect 6967 789 7133 819
rect 7203 789 7369 819
rect 7415 819 7420 820
rect 7812 820 7868 823
rect 7812 819 7817 820
rect 7415 789 7581 819
rect 7651 789 7817 819
rect 7863 819 7868 820
rect 8260 820 8316 823
rect 8260 819 8265 820
rect 7863 789 8029 819
rect 8099 789 8265 819
rect 8311 819 8316 820
rect 8708 820 8764 823
rect 8708 819 8713 820
rect 8311 789 8477 819
rect 8547 789 8713 819
rect 8759 819 8764 820
rect 8759 789 8925 819
rect 196 785 252 789
rect 644 785 700 789
rect 1092 785 1148 789
rect 1540 785 1596 789
rect 1988 785 2044 789
rect 2436 785 2492 789
rect 2884 785 2940 789
rect 3332 785 3388 789
rect 3780 785 3836 789
rect 4228 785 4284 789
rect 4676 785 4732 789
rect 5124 785 5180 789
rect 5572 785 5628 789
rect 6020 785 6076 789
rect 6468 785 6524 789
rect 6916 785 6972 789
rect 7364 785 7420 789
rect 7812 785 7868 789
rect 8260 785 8316 789
rect 8708 785 8764 789
rect 99 758 137 759
rect 99 757 102 758
rect 54 727 102 757
rect 99 726 102 727
rect 134 757 137 758
rect 311 758 349 759
rect 311 757 314 758
rect 134 727 181 757
rect 267 727 314 757
rect 134 726 137 727
rect 99 725 137 726
rect 311 726 314 727
rect 346 757 349 758
rect 547 758 585 759
rect 547 757 550 758
rect 346 727 394 757
rect 502 727 550 757
rect 346 726 349 727
rect 311 725 349 726
rect 547 726 550 727
rect 582 757 585 758
rect 759 758 797 759
rect 759 757 762 758
rect 582 727 629 757
rect 715 727 762 757
rect 582 726 585 727
rect 547 725 585 726
rect 759 726 762 727
rect 794 757 797 758
rect 995 758 1033 759
rect 995 757 998 758
rect 794 727 842 757
rect 950 727 998 757
rect 794 726 797 727
rect 759 725 797 726
rect 995 726 998 727
rect 1030 757 1033 758
rect 1207 758 1245 759
rect 1207 757 1210 758
rect 1030 727 1077 757
rect 1163 727 1210 757
rect 1030 726 1033 727
rect 995 725 1033 726
rect 1207 726 1210 727
rect 1242 757 1245 758
rect 1443 758 1481 759
rect 1443 757 1446 758
rect 1242 727 1290 757
rect 1398 727 1446 757
rect 1242 726 1245 727
rect 1207 725 1245 726
rect 1443 726 1446 727
rect 1478 757 1481 758
rect 1655 758 1693 759
rect 1655 757 1658 758
rect 1478 727 1525 757
rect 1611 727 1658 757
rect 1478 726 1481 727
rect 1443 725 1481 726
rect 1655 726 1658 727
rect 1690 757 1693 758
rect 1891 758 1929 759
rect 1891 757 1894 758
rect 1690 727 1738 757
rect 1846 727 1894 757
rect 1690 726 1693 727
rect 1655 725 1693 726
rect 1891 726 1894 727
rect 1926 757 1929 758
rect 2103 758 2141 759
rect 2103 757 2106 758
rect 1926 727 1973 757
rect 2059 727 2106 757
rect 1926 726 1929 727
rect 1891 725 1929 726
rect 2103 726 2106 727
rect 2138 757 2141 758
rect 2339 758 2377 759
rect 2339 757 2342 758
rect 2138 727 2186 757
rect 2294 727 2342 757
rect 2138 726 2141 727
rect 2103 725 2141 726
rect 2339 726 2342 727
rect 2374 757 2377 758
rect 2551 758 2589 759
rect 2551 757 2554 758
rect 2374 727 2421 757
rect 2507 727 2554 757
rect 2374 726 2377 727
rect 2339 725 2377 726
rect 2551 726 2554 727
rect 2586 757 2589 758
rect 2787 758 2825 759
rect 2787 757 2790 758
rect 2586 727 2634 757
rect 2742 727 2790 757
rect 2586 726 2589 727
rect 2551 725 2589 726
rect 2787 726 2790 727
rect 2822 757 2825 758
rect 2999 758 3037 759
rect 2999 757 3002 758
rect 2822 727 2869 757
rect 2955 727 3002 757
rect 2822 726 2825 727
rect 2787 725 2825 726
rect 2999 726 3002 727
rect 3034 757 3037 758
rect 3235 758 3273 759
rect 3235 757 3238 758
rect 3034 727 3082 757
rect 3190 727 3238 757
rect 3034 726 3037 727
rect 2999 725 3037 726
rect 3235 726 3238 727
rect 3270 757 3273 758
rect 3447 758 3485 759
rect 3447 757 3450 758
rect 3270 727 3317 757
rect 3403 727 3450 757
rect 3270 726 3273 727
rect 3235 725 3273 726
rect 3447 726 3450 727
rect 3482 757 3485 758
rect 3683 758 3721 759
rect 3683 757 3686 758
rect 3482 727 3530 757
rect 3638 727 3686 757
rect 3482 726 3485 727
rect 3447 725 3485 726
rect 3683 726 3686 727
rect 3718 757 3721 758
rect 3895 758 3933 759
rect 3895 757 3898 758
rect 3718 727 3765 757
rect 3851 727 3898 757
rect 3718 726 3721 727
rect 3683 725 3721 726
rect 3895 726 3898 727
rect 3930 757 3933 758
rect 4131 758 4169 759
rect 4131 757 4134 758
rect 3930 727 3978 757
rect 4086 727 4134 757
rect 3930 726 3933 727
rect 3895 725 3933 726
rect 4131 726 4134 727
rect 4166 757 4169 758
rect 4343 758 4381 759
rect 4343 757 4346 758
rect 4166 727 4213 757
rect 4299 727 4346 757
rect 4166 726 4169 727
rect 4131 725 4169 726
rect 4343 726 4346 727
rect 4378 757 4381 758
rect 4579 758 4617 759
rect 4579 757 4582 758
rect 4378 727 4426 757
rect 4534 727 4582 757
rect 4378 726 4381 727
rect 4343 725 4381 726
rect 4579 726 4582 727
rect 4614 757 4617 758
rect 4791 758 4829 759
rect 4791 757 4794 758
rect 4614 727 4661 757
rect 4747 727 4794 757
rect 4614 726 4617 727
rect 4579 725 4617 726
rect 4791 726 4794 727
rect 4826 757 4829 758
rect 5027 758 5065 759
rect 5027 757 5030 758
rect 4826 727 4874 757
rect 4982 727 5030 757
rect 4826 726 4829 727
rect 4791 725 4829 726
rect 5027 726 5030 727
rect 5062 757 5065 758
rect 5239 758 5277 759
rect 5239 757 5242 758
rect 5062 727 5109 757
rect 5195 727 5242 757
rect 5062 726 5065 727
rect 5027 725 5065 726
rect 5239 726 5242 727
rect 5274 757 5277 758
rect 5475 758 5513 759
rect 5475 757 5478 758
rect 5274 727 5322 757
rect 5430 727 5478 757
rect 5274 726 5277 727
rect 5239 725 5277 726
rect 5475 726 5478 727
rect 5510 757 5513 758
rect 5687 758 5725 759
rect 5687 757 5690 758
rect 5510 727 5557 757
rect 5643 727 5690 757
rect 5510 726 5513 727
rect 5475 725 5513 726
rect 5687 726 5690 727
rect 5722 757 5725 758
rect 5923 758 5961 759
rect 5923 757 5926 758
rect 5722 727 5770 757
rect 5878 727 5926 757
rect 5722 726 5725 727
rect 5687 725 5725 726
rect 5923 726 5926 727
rect 5958 757 5961 758
rect 6135 758 6173 759
rect 6135 757 6138 758
rect 5958 727 6005 757
rect 6091 727 6138 757
rect 5958 726 5961 727
rect 5923 725 5961 726
rect 6135 726 6138 727
rect 6170 757 6173 758
rect 6371 758 6409 759
rect 6371 757 6374 758
rect 6170 727 6218 757
rect 6326 727 6374 757
rect 6170 726 6173 727
rect 6135 725 6173 726
rect 6371 726 6374 727
rect 6406 757 6409 758
rect 6583 758 6621 759
rect 6583 757 6586 758
rect 6406 727 6453 757
rect 6539 727 6586 757
rect 6406 726 6409 727
rect 6371 725 6409 726
rect 6583 726 6586 727
rect 6618 757 6621 758
rect 6819 758 6857 759
rect 6819 757 6822 758
rect 6618 727 6666 757
rect 6774 727 6822 757
rect 6618 726 6621 727
rect 6583 725 6621 726
rect 6819 726 6822 727
rect 6854 757 6857 758
rect 7031 758 7069 759
rect 7031 757 7034 758
rect 6854 727 6901 757
rect 6987 727 7034 757
rect 6854 726 6857 727
rect 6819 725 6857 726
rect 7031 726 7034 727
rect 7066 757 7069 758
rect 7267 758 7305 759
rect 7267 757 7270 758
rect 7066 727 7114 757
rect 7222 727 7270 757
rect 7066 726 7069 727
rect 7031 725 7069 726
rect 7267 726 7270 727
rect 7302 757 7305 758
rect 7479 758 7517 759
rect 7479 757 7482 758
rect 7302 727 7349 757
rect 7435 727 7482 757
rect 7302 726 7305 727
rect 7267 725 7305 726
rect 7479 726 7482 727
rect 7514 757 7517 758
rect 7715 758 7753 759
rect 7715 757 7718 758
rect 7514 727 7562 757
rect 7670 727 7718 757
rect 7514 726 7517 727
rect 7479 725 7517 726
rect 7715 726 7718 727
rect 7750 757 7753 758
rect 7927 758 7965 759
rect 7927 757 7930 758
rect 7750 727 7797 757
rect 7883 727 7930 757
rect 7750 726 7753 727
rect 7715 725 7753 726
rect 7927 726 7930 727
rect 7962 757 7965 758
rect 8163 758 8201 759
rect 8163 757 8166 758
rect 7962 727 8010 757
rect 8118 727 8166 757
rect 7962 726 7965 727
rect 7927 725 7965 726
rect 8163 726 8166 727
rect 8198 757 8201 758
rect 8375 758 8413 759
rect 8375 757 8378 758
rect 8198 727 8245 757
rect 8331 727 8378 757
rect 8198 726 8201 727
rect 8163 725 8201 726
rect 8375 726 8378 727
rect 8410 757 8413 758
rect 8611 758 8649 759
rect 8611 757 8614 758
rect 8410 727 8458 757
rect 8566 727 8614 757
rect 8410 726 8413 727
rect 8375 725 8413 726
rect 8611 726 8614 727
rect 8646 757 8649 758
rect 8823 758 8861 759
rect 8823 757 8826 758
rect 8646 727 8693 757
rect 8779 727 8826 757
rect 8646 726 8649 727
rect 8611 725 8649 726
rect 8823 726 8826 727
rect 8858 757 8861 758
rect 8858 727 8906 757
rect 8858 726 8861 727
rect 8823 725 8861 726
rect 196 696 252 699
rect 196 695 201 696
rect 35 665 201 695
rect 247 695 252 696
rect 644 696 700 699
rect 644 695 649 696
rect 247 665 413 695
rect 483 665 649 695
rect 695 695 700 696
rect 1092 696 1148 699
rect 1092 695 1097 696
rect 695 665 861 695
rect 931 665 1097 695
rect 1143 695 1148 696
rect 1540 696 1596 699
rect 1540 695 1545 696
rect 1143 665 1309 695
rect 1379 665 1545 695
rect 1591 695 1596 696
rect 1988 696 2044 699
rect 1988 695 1993 696
rect 1591 665 1757 695
rect 1827 665 1993 695
rect 2039 695 2044 696
rect 2436 696 2492 699
rect 2436 695 2441 696
rect 2039 665 2205 695
rect 2275 665 2441 695
rect 2487 695 2492 696
rect 2884 696 2940 699
rect 2884 695 2889 696
rect 2487 665 2653 695
rect 2723 665 2889 695
rect 2935 695 2940 696
rect 3332 696 3388 699
rect 3332 695 3337 696
rect 2935 665 3101 695
rect 3171 665 3337 695
rect 3383 695 3388 696
rect 3780 696 3836 699
rect 3780 695 3785 696
rect 3383 665 3549 695
rect 3619 665 3785 695
rect 3831 695 3836 696
rect 4228 696 4284 699
rect 4228 695 4233 696
rect 3831 665 3997 695
rect 4067 665 4233 695
rect 4279 695 4284 696
rect 4676 696 4732 699
rect 4676 695 4681 696
rect 4279 665 4445 695
rect 4515 665 4681 695
rect 4727 695 4732 696
rect 5124 696 5180 699
rect 5124 695 5129 696
rect 4727 665 4893 695
rect 4963 665 5129 695
rect 5175 695 5180 696
rect 5572 696 5628 699
rect 5572 695 5577 696
rect 5175 665 5341 695
rect 5411 665 5577 695
rect 5623 695 5628 696
rect 6020 696 6076 699
rect 6020 695 6025 696
rect 5623 665 5789 695
rect 5859 665 6025 695
rect 6071 695 6076 696
rect 6468 696 6524 699
rect 6468 695 6473 696
rect 6071 665 6237 695
rect 6307 665 6473 695
rect 6519 695 6524 696
rect 6916 696 6972 699
rect 6916 695 6921 696
rect 6519 665 6685 695
rect 6755 665 6921 695
rect 6967 695 6972 696
rect 7364 696 7420 699
rect 7364 695 7369 696
rect 6967 665 7133 695
rect 7203 665 7369 695
rect 7415 695 7420 696
rect 7812 696 7868 699
rect 7812 695 7817 696
rect 7415 665 7581 695
rect 7651 665 7817 695
rect 7863 695 7868 696
rect 8260 696 8316 699
rect 8260 695 8265 696
rect 7863 665 8029 695
rect 8099 665 8265 695
rect 8311 695 8316 696
rect 8708 696 8764 699
rect 8708 695 8713 696
rect 8311 665 8477 695
rect 8547 665 8713 695
rect 8759 695 8764 696
rect 8759 665 8925 695
rect 196 661 252 665
rect 644 661 700 665
rect 1092 661 1148 665
rect 1540 661 1596 665
rect 1988 661 2044 665
rect 2436 661 2492 665
rect 2884 661 2940 665
rect 3332 661 3388 665
rect 3780 661 3836 665
rect 4228 661 4284 665
rect 4676 661 4732 665
rect 5124 661 5180 665
rect 5572 661 5628 665
rect 6020 661 6076 665
rect 6468 661 6524 665
rect 6916 661 6972 665
rect 7364 661 7420 665
rect 7812 661 7868 665
rect 8260 661 8316 665
rect 8708 661 8764 665
rect 196 574 252 577
rect 196 573 201 574
rect 35 543 201 573
rect 247 573 252 574
rect 644 574 700 577
rect 644 573 649 574
rect 247 543 413 573
rect 483 543 649 573
rect 695 573 700 574
rect 1092 574 1148 577
rect 1092 573 1097 574
rect 695 543 861 573
rect 931 543 1097 573
rect 1143 573 1148 574
rect 1540 574 1596 577
rect 1540 573 1545 574
rect 1143 543 1309 573
rect 1379 543 1545 573
rect 1591 573 1596 574
rect 1988 574 2044 577
rect 1988 573 1993 574
rect 1591 543 1757 573
rect 1827 543 1993 573
rect 2039 573 2044 574
rect 2436 574 2492 577
rect 2436 573 2441 574
rect 2039 543 2205 573
rect 2275 543 2441 573
rect 2487 573 2492 574
rect 2884 574 2940 577
rect 2884 573 2889 574
rect 2487 543 2653 573
rect 2723 543 2889 573
rect 2935 573 2940 574
rect 3332 574 3388 577
rect 3332 573 3337 574
rect 2935 543 3101 573
rect 3171 543 3337 573
rect 3383 573 3388 574
rect 3780 574 3836 577
rect 3780 573 3785 574
rect 3383 543 3549 573
rect 3619 543 3785 573
rect 3831 573 3836 574
rect 4228 574 4284 577
rect 4228 573 4233 574
rect 3831 543 3997 573
rect 4067 543 4233 573
rect 4279 573 4284 574
rect 4676 574 4732 577
rect 4676 573 4681 574
rect 4279 543 4445 573
rect 4515 543 4681 573
rect 4727 573 4732 574
rect 5124 574 5180 577
rect 5124 573 5129 574
rect 4727 543 4893 573
rect 4963 543 5129 573
rect 5175 573 5180 574
rect 5572 574 5628 577
rect 5572 573 5577 574
rect 5175 543 5341 573
rect 5411 543 5577 573
rect 5623 573 5628 574
rect 6020 574 6076 577
rect 6020 573 6025 574
rect 5623 543 5789 573
rect 5859 543 6025 573
rect 6071 573 6076 574
rect 6468 574 6524 577
rect 6468 573 6473 574
rect 6071 543 6237 573
rect 6307 543 6473 573
rect 6519 573 6524 574
rect 6916 574 6972 577
rect 6916 573 6921 574
rect 6519 543 6685 573
rect 6755 543 6921 573
rect 6967 573 6972 574
rect 7364 574 7420 577
rect 7364 573 7369 574
rect 6967 543 7133 573
rect 7203 543 7369 573
rect 7415 573 7420 574
rect 7812 574 7868 577
rect 7812 573 7817 574
rect 7415 543 7581 573
rect 7651 543 7817 573
rect 7863 573 7868 574
rect 8260 574 8316 577
rect 8260 573 8265 574
rect 7863 543 8029 573
rect 8099 543 8265 573
rect 8311 573 8316 574
rect 8708 574 8764 577
rect 8708 573 8713 574
rect 8311 543 8477 573
rect 8547 543 8713 573
rect 8759 573 8764 574
rect 8759 543 8925 573
rect 196 539 252 543
rect 644 539 700 543
rect 1092 539 1148 543
rect 1540 539 1596 543
rect 1988 539 2044 543
rect 2436 539 2492 543
rect 2884 539 2940 543
rect 3332 539 3388 543
rect 3780 539 3836 543
rect 4228 539 4284 543
rect 4676 539 4732 543
rect 5124 539 5180 543
rect 5572 539 5628 543
rect 6020 539 6076 543
rect 6468 539 6524 543
rect 6916 539 6972 543
rect 7364 539 7420 543
rect 7812 539 7868 543
rect 8260 539 8316 543
rect 8708 539 8764 543
rect 99 511 137 512
rect 99 510 102 511
rect 54 480 102 510
rect 99 479 102 480
rect 134 510 137 511
rect 311 511 349 512
rect 311 510 314 511
rect 134 480 181 510
rect 267 480 314 510
rect 134 479 137 480
rect 99 478 137 479
rect 311 479 314 480
rect 346 510 349 511
rect 547 511 585 512
rect 547 510 550 511
rect 346 480 394 510
rect 502 480 550 510
rect 346 479 349 480
rect 311 478 349 479
rect 547 479 550 480
rect 582 510 585 511
rect 759 511 797 512
rect 759 510 762 511
rect 582 480 629 510
rect 715 480 762 510
rect 582 479 585 480
rect 547 478 585 479
rect 759 479 762 480
rect 794 510 797 511
rect 995 511 1033 512
rect 995 510 998 511
rect 794 480 842 510
rect 950 480 998 510
rect 794 479 797 480
rect 759 478 797 479
rect 995 479 998 480
rect 1030 510 1033 511
rect 1207 511 1245 512
rect 1207 510 1210 511
rect 1030 480 1077 510
rect 1163 480 1210 510
rect 1030 479 1033 480
rect 995 478 1033 479
rect 1207 479 1210 480
rect 1242 510 1245 511
rect 1443 511 1481 512
rect 1443 510 1446 511
rect 1242 480 1290 510
rect 1398 480 1446 510
rect 1242 479 1245 480
rect 1207 478 1245 479
rect 1443 479 1446 480
rect 1478 510 1481 511
rect 1655 511 1693 512
rect 1655 510 1658 511
rect 1478 480 1525 510
rect 1611 480 1658 510
rect 1478 479 1481 480
rect 1443 478 1481 479
rect 1655 479 1658 480
rect 1690 510 1693 511
rect 1891 511 1929 512
rect 1891 510 1894 511
rect 1690 480 1738 510
rect 1846 480 1894 510
rect 1690 479 1693 480
rect 1655 478 1693 479
rect 1891 479 1894 480
rect 1926 510 1929 511
rect 2103 511 2141 512
rect 2103 510 2106 511
rect 1926 480 1973 510
rect 2059 480 2106 510
rect 1926 479 1929 480
rect 1891 478 1929 479
rect 2103 479 2106 480
rect 2138 510 2141 511
rect 2339 511 2377 512
rect 2339 510 2342 511
rect 2138 480 2186 510
rect 2294 480 2342 510
rect 2138 479 2141 480
rect 2103 478 2141 479
rect 2339 479 2342 480
rect 2374 510 2377 511
rect 2551 511 2589 512
rect 2551 510 2554 511
rect 2374 480 2421 510
rect 2507 480 2554 510
rect 2374 479 2377 480
rect 2339 478 2377 479
rect 2551 479 2554 480
rect 2586 510 2589 511
rect 2787 511 2825 512
rect 2787 510 2790 511
rect 2586 480 2634 510
rect 2742 480 2790 510
rect 2586 479 2589 480
rect 2551 478 2589 479
rect 2787 479 2790 480
rect 2822 510 2825 511
rect 2999 511 3037 512
rect 2999 510 3002 511
rect 2822 480 2869 510
rect 2955 480 3002 510
rect 2822 479 2825 480
rect 2787 478 2825 479
rect 2999 479 3002 480
rect 3034 510 3037 511
rect 3235 511 3273 512
rect 3235 510 3238 511
rect 3034 480 3082 510
rect 3190 480 3238 510
rect 3034 479 3037 480
rect 2999 478 3037 479
rect 3235 479 3238 480
rect 3270 510 3273 511
rect 3447 511 3485 512
rect 3447 510 3450 511
rect 3270 480 3317 510
rect 3403 480 3450 510
rect 3270 479 3273 480
rect 3235 478 3273 479
rect 3447 479 3450 480
rect 3482 510 3485 511
rect 3683 511 3721 512
rect 3683 510 3686 511
rect 3482 480 3530 510
rect 3638 480 3686 510
rect 3482 479 3485 480
rect 3447 478 3485 479
rect 3683 479 3686 480
rect 3718 510 3721 511
rect 3895 511 3933 512
rect 3895 510 3898 511
rect 3718 480 3765 510
rect 3851 480 3898 510
rect 3718 479 3721 480
rect 3683 478 3721 479
rect 3895 479 3898 480
rect 3930 510 3933 511
rect 4131 511 4169 512
rect 4131 510 4134 511
rect 3930 480 3978 510
rect 4086 480 4134 510
rect 3930 479 3933 480
rect 3895 478 3933 479
rect 4131 479 4134 480
rect 4166 510 4169 511
rect 4343 511 4381 512
rect 4343 510 4346 511
rect 4166 480 4213 510
rect 4299 480 4346 510
rect 4166 479 4169 480
rect 4131 478 4169 479
rect 4343 479 4346 480
rect 4378 510 4381 511
rect 4579 511 4617 512
rect 4579 510 4582 511
rect 4378 480 4426 510
rect 4534 480 4582 510
rect 4378 479 4381 480
rect 4343 478 4381 479
rect 4579 479 4582 480
rect 4614 510 4617 511
rect 4791 511 4829 512
rect 4791 510 4794 511
rect 4614 480 4661 510
rect 4747 480 4794 510
rect 4614 479 4617 480
rect 4579 478 4617 479
rect 4791 479 4794 480
rect 4826 510 4829 511
rect 5027 511 5065 512
rect 5027 510 5030 511
rect 4826 480 4874 510
rect 4982 480 5030 510
rect 4826 479 4829 480
rect 4791 478 4829 479
rect 5027 479 5030 480
rect 5062 510 5065 511
rect 5239 511 5277 512
rect 5239 510 5242 511
rect 5062 480 5109 510
rect 5195 480 5242 510
rect 5062 479 5065 480
rect 5027 478 5065 479
rect 5239 479 5242 480
rect 5274 510 5277 511
rect 5475 511 5513 512
rect 5475 510 5478 511
rect 5274 480 5322 510
rect 5430 480 5478 510
rect 5274 479 5277 480
rect 5239 478 5277 479
rect 5475 479 5478 480
rect 5510 510 5513 511
rect 5687 511 5725 512
rect 5687 510 5690 511
rect 5510 480 5557 510
rect 5643 480 5690 510
rect 5510 479 5513 480
rect 5475 478 5513 479
rect 5687 479 5690 480
rect 5722 510 5725 511
rect 5923 511 5961 512
rect 5923 510 5926 511
rect 5722 480 5770 510
rect 5878 480 5926 510
rect 5722 479 5725 480
rect 5687 478 5725 479
rect 5923 479 5926 480
rect 5958 510 5961 511
rect 6135 511 6173 512
rect 6135 510 6138 511
rect 5958 480 6005 510
rect 6091 480 6138 510
rect 5958 479 5961 480
rect 5923 478 5961 479
rect 6135 479 6138 480
rect 6170 510 6173 511
rect 6371 511 6409 512
rect 6371 510 6374 511
rect 6170 480 6218 510
rect 6326 480 6374 510
rect 6170 479 6173 480
rect 6135 478 6173 479
rect 6371 479 6374 480
rect 6406 510 6409 511
rect 6583 511 6621 512
rect 6583 510 6586 511
rect 6406 480 6453 510
rect 6539 480 6586 510
rect 6406 479 6409 480
rect 6371 478 6409 479
rect 6583 479 6586 480
rect 6618 510 6621 511
rect 6819 511 6857 512
rect 6819 510 6822 511
rect 6618 480 6666 510
rect 6774 480 6822 510
rect 6618 479 6621 480
rect 6583 478 6621 479
rect 6819 479 6822 480
rect 6854 510 6857 511
rect 7031 511 7069 512
rect 7031 510 7034 511
rect 6854 480 6901 510
rect 6987 480 7034 510
rect 6854 479 6857 480
rect 6819 478 6857 479
rect 7031 479 7034 480
rect 7066 510 7069 511
rect 7267 511 7305 512
rect 7267 510 7270 511
rect 7066 480 7114 510
rect 7222 480 7270 510
rect 7066 479 7069 480
rect 7031 478 7069 479
rect 7267 479 7270 480
rect 7302 510 7305 511
rect 7479 511 7517 512
rect 7479 510 7482 511
rect 7302 480 7349 510
rect 7435 480 7482 510
rect 7302 479 7305 480
rect 7267 478 7305 479
rect 7479 479 7482 480
rect 7514 510 7517 511
rect 7715 511 7753 512
rect 7715 510 7718 511
rect 7514 480 7562 510
rect 7670 480 7718 510
rect 7514 479 7517 480
rect 7479 478 7517 479
rect 7715 479 7718 480
rect 7750 510 7753 511
rect 7927 511 7965 512
rect 7927 510 7930 511
rect 7750 480 7797 510
rect 7883 480 7930 510
rect 7750 479 7753 480
rect 7715 478 7753 479
rect 7927 479 7930 480
rect 7962 510 7965 511
rect 8163 511 8201 512
rect 8163 510 8166 511
rect 7962 480 8010 510
rect 8118 480 8166 510
rect 7962 479 7965 480
rect 7927 478 7965 479
rect 8163 479 8166 480
rect 8198 510 8201 511
rect 8375 511 8413 512
rect 8375 510 8378 511
rect 8198 480 8245 510
rect 8331 480 8378 510
rect 8198 479 8201 480
rect 8163 478 8201 479
rect 8375 479 8378 480
rect 8410 510 8413 511
rect 8611 511 8649 512
rect 8611 510 8614 511
rect 8410 480 8458 510
rect 8566 480 8614 510
rect 8410 479 8413 480
rect 8375 478 8413 479
rect 8611 479 8614 480
rect 8646 510 8649 511
rect 8823 511 8861 512
rect 8823 510 8826 511
rect 8646 480 8693 510
rect 8779 480 8826 510
rect 8646 479 8649 480
rect 8611 478 8649 479
rect 8823 479 8826 480
rect 8858 510 8861 511
rect 8858 480 8906 510
rect 8858 479 8861 480
rect 8823 478 8861 479
rect 196 449 252 452
rect 196 448 201 449
rect 35 418 201 448
rect 247 448 252 449
rect 644 449 700 452
rect 644 448 649 449
rect 247 418 413 448
rect 483 418 649 448
rect 695 448 700 449
rect 1092 449 1148 452
rect 1092 448 1097 449
rect 695 418 861 448
rect 931 418 1097 448
rect 1143 448 1148 449
rect 1540 449 1596 452
rect 1540 448 1545 449
rect 1143 418 1309 448
rect 1379 418 1545 448
rect 1591 448 1596 449
rect 1988 449 2044 452
rect 1988 448 1993 449
rect 1591 418 1757 448
rect 1827 418 1993 448
rect 2039 448 2044 449
rect 2436 449 2492 452
rect 2436 448 2441 449
rect 2039 418 2205 448
rect 2275 418 2441 448
rect 2487 448 2492 449
rect 2884 449 2940 452
rect 2884 448 2889 449
rect 2487 418 2653 448
rect 2723 418 2889 448
rect 2935 448 2940 449
rect 3332 449 3388 452
rect 3332 448 3337 449
rect 2935 418 3101 448
rect 3171 418 3337 448
rect 3383 448 3388 449
rect 3780 449 3836 452
rect 3780 448 3785 449
rect 3383 418 3549 448
rect 3619 418 3785 448
rect 3831 448 3836 449
rect 4228 449 4284 452
rect 4228 448 4233 449
rect 3831 418 3997 448
rect 4067 418 4233 448
rect 4279 448 4284 449
rect 4676 449 4732 452
rect 4676 448 4681 449
rect 4279 418 4445 448
rect 4515 418 4681 448
rect 4727 448 4732 449
rect 5124 449 5180 452
rect 5124 448 5129 449
rect 4727 418 4893 448
rect 4963 418 5129 448
rect 5175 448 5180 449
rect 5572 449 5628 452
rect 5572 448 5577 449
rect 5175 418 5341 448
rect 5411 418 5577 448
rect 5623 448 5628 449
rect 6020 449 6076 452
rect 6020 448 6025 449
rect 5623 418 5789 448
rect 5859 418 6025 448
rect 6071 448 6076 449
rect 6468 449 6524 452
rect 6468 448 6473 449
rect 6071 418 6237 448
rect 6307 418 6473 448
rect 6519 448 6524 449
rect 6916 449 6972 452
rect 6916 448 6921 449
rect 6519 418 6685 448
rect 6755 418 6921 448
rect 6967 448 6972 449
rect 7364 449 7420 452
rect 7364 448 7369 449
rect 6967 418 7133 448
rect 7203 418 7369 448
rect 7415 448 7420 449
rect 7812 449 7868 452
rect 7812 448 7817 449
rect 7415 418 7581 448
rect 7651 418 7817 448
rect 7863 448 7868 449
rect 8260 449 8316 452
rect 8260 448 8265 449
rect 7863 418 8029 448
rect 8099 418 8265 448
rect 8311 448 8316 449
rect 8708 449 8764 452
rect 8708 448 8713 449
rect 8311 418 8477 448
rect 8547 418 8713 448
rect 8759 448 8764 449
rect 8759 418 8925 448
rect 196 414 252 418
rect 644 414 700 418
rect 1092 414 1148 418
rect 1540 414 1596 418
rect 1988 414 2044 418
rect 2436 414 2492 418
rect 2884 414 2940 418
rect 3332 414 3388 418
rect 3780 414 3836 418
rect 4228 414 4284 418
rect 4676 414 4732 418
rect 5124 414 5180 418
rect 5572 414 5628 418
rect 6020 414 6076 418
rect 6468 414 6524 418
rect 6916 414 6972 418
rect 7364 414 7420 418
rect 7812 414 7868 418
rect 8260 414 8316 418
rect 8708 414 8764 418
rect 99 387 137 388
rect 99 386 102 387
rect 54 356 102 386
rect 99 355 102 356
rect 134 386 137 387
rect 311 387 349 388
rect 311 386 314 387
rect 134 356 181 386
rect 267 356 314 386
rect 134 355 137 356
rect 99 354 137 355
rect 311 355 314 356
rect 346 386 349 387
rect 547 387 585 388
rect 547 386 550 387
rect 346 356 394 386
rect 502 356 550 386
rect 346 355 349 356
rect 311 354 349 355
rect 547 355 550 356
rect 582 386 585 387
rect 759 387 797 388
rect 759 386 762 387
rect 582 356 629 386
rect 715 356 762 386
rect 582 355 585 356
rect 547 354 585 355
rect 759 355 762 356
rect 794 386 797 387
rect 995 387 1033 388
rect 995 386 998 387
rect 794 356 842 386
rect 950 356 998 386
rect 794 355 797 356
rect 759 354 797 355
rect 995 355 998 356
rect 1030 386 1033 387
rect 1207 387 1245 388
rect 1207 386 1210 387
rect 1030 356 1077 386
rect 1163 356 1210 386
rect 1030 355 1033 356
rect 995 354 1033 355
rect 1207 355 1210 356
rect 1242 386 1245 387
rect 1443 387 1481 388
rect 1443 386 1446 387
rect 1242 356 1290 386
rect 1398 356 1446 386
rect 1242 355 1245 356
rect 1207 354 1245 355
rect 1443 355 1446 356
rect 1478 386 1481 387
rect 1655 387 1693 388
rect 1655 386 1658 387
rect 1478 356 1525 386
rect 1611 356 1658 386
rect 1478 355 1481 356
rect 1443 354 1481 355
rect 1655 355 1658 356
rect 1690 386 1693 387
rect 1891 387 1929 388
rect 1891 386 1894 387
rect 1690 356 1738 386
rect 1846 356 1894 386
rect 1690 355 1693 356
rect 1655 354 1693 355
rect 1891 355 1894 356
rect 1926 386 1929 387
rect 2103 387 2141 388
rect 2103 386 2106 387
rect 1926 356 1973 386
rect 2059 356 2106 386
rect 1926 355 1929 356
rect 1891 354 1929 355
rect 2103 355 2106 356
rect 2138 386 2141 387
rect 2339 387 2377 388
rect 2339 386 2342 387
rect 2138 356 2186 386
rect 2294 356 2342 386
rect 2138 355 2141 356
rect 2103 354 2141 355
rect 2339 355 2342 356
rect 2374 386 2377 387
rect 2551 387 2589 388
rect 2551 386 2554 387
rect 2374 356 2421 386
rect 2507 356 2554 386
rect 2374 355 2377 356
rect 2339 354 2377 355
rect 2551 355 2554 356
rect 2586 386 2589 387
rect 2787 387 2825 388
rect 2787 386 2790 387
rect 2586 356 2634 386
rect 2742 356 2790 386
rect 2586 355 2589 356
rect 2551 354 2589 355
rect 2787 355 2790 356
rect 2822 386 2825 387
rect 2999 387 3037 388
rect 2999 386 3002 387
rect 2822 356 2869 386
rect 2955 356 3002 386
rect 2822 355 2825 356
rect 2787 354 2825 355
rect 2999 355 3002 356
rect 3034 386 3037 387
rect 3235 387 3273 388
rect 3235 386 3238 387
rect 3034 356 3082 386
rect 3190 356 3238 386
rect 3034 355 3037 356
rect 2999 354 3037 355
rect 3235 355 3238 356
rect 3270 386 3273 387
rect 3447 387 3485 388
rect 3447 386 3450 387
rect 3270 356 3317 386
rect 3403 356 3450 386
rect 3270 355 3273 356
rect 3235 354 3273 355
rect 3447 355 3450 356
rect 3482 386 3485 387
rect 3683 387 3721 388
rect 3683 386 3686 387
rect 3482 356 3530 386
rect 3638 356 3686 386
rect 3482 355 3485 356
rect 3447 354 3485 355
rect 3683 355 3686 356
rect 3718 386 3721 387
rect 3895 387 3933 388
rect 3895 386 3898 387
rect 3718 356 3765 386
rect 3851 356 3898 386
rect 3718 355 3721 356
rect 3683 354 3721 355
rect 3895 355 3898 356
rect 3930 386 3933 387
rect 4131 387 4169 388
rect 4131 386 4134 387
rect 3930 356 3978 386
rect 4086 356 4134 386
rect 3930 355 3933 356
rect 3895 354 3933 355
rect 4131 355 4134 356
rect 4166 386 4169 387
rect 4343 387 4381 388
rect 4343 386 4346 387
rect 4166 356 4213 386
rect 4299 356 4346 386
rect 4166 355 4169 356
rect 4131 354 4169 355
rect 4343 355 4346 356
rect 4378 386 4381 387
rect 4579 387 4617 388
rect 4579 386 4582 387
rect 4378 356 4426 386
rect 4534 356 4582 386
rect 4378 355 4381 356
rect 4343 354 4381 355
rect 4579 355 4582 356
rect 4614 386 4617 387
rect 4791 387 4829 388
rect 4791 386 4794 387
rect 4614 356 4661 386
rect 4747 356 4794 386
rect 4614 355 4617 356
rect 4579 354 4617 355
rect 4791 355 4794 356
rect 4826 386 4829 387
rect 5027 387 5065 388
rect 5027 386 5030 387
rect 4826 356 4874 386
rect 4982 356 5030 386
rect 4826 355 4829 356
rect 4791 354 4829 355
rect 5027 355 5030 356
rect 5062 386 5065 387
rect 5239 387 5277 388
rect 5239 386 5242 387
rect 5062 356 5109 386
rect 5195 356 5242 386
rect 5062 355 5065 356
rect 5027 354 5065 355
rect 5239 355 5242 356
rect 5274 386 5277 387
rect 5475 387 5513 388
rect 5475 386 5478 387
rect 5274 356 5322 386
rect 5430 356 5478 386
rect 5274 355 5277 356
rect 5239 354 5277 355
rect 5475 355 5478 356
rect 5510 386 5513 387
rect 5687 387 5725 388
rect 5687 386 5690 387
rect 5510 356 5557 386
rect 5643 356 5690 386
rect 5510 355 5513 356
rect 5475 354 5513 355
rect 5687 355 5690 356
rect 5722 386 5725 387
rect 5923 387 5961 388
rect 5923 386 5926 387
rect 5722 356 5770 386
rect 5878 356 5926 386
rect 5722 355 5725 356
rect 5687 354 5725 355
rect 5923 355 5926 356
rect 5958 386 5961 387
rect 6135 387 6173 388
rect 6135 386 6138 387
rect 5958 356 6005 386
rect 6091 356 6138 386
rect 5958 355 5961 356
rect 5923 354 5961 355
rect 6135 355 6138 356
rect 6170 386 6173 387
rect 6371 387 6409 388
rect 6371 386 6374 387
rect 6170 356 6218 386
rect 6326 356 6374 386
rect 6170 355 6173 356
rect 6135 354 6173 355
rect 6371 355 6374 356
rect 6406 386 6409 387
rect 6583 387 6621 388
rect 6583 386 6586 387
rect 6406 356 6453 386
rect 6539 356 6586 386
rect 6406 355 6409 356
rect 6371 354 6409 355
rect 6583 355 6586 356
rect 6618 386 6621 387
rect 6819 387 6857 388
rect 6819 386 6822 387
rect 6618 356 6666 386
rect 6774 356 6822 386
rect 6618 355 6621 356
rect 6583 354 6621 355
rect 6819 355 6822 356
rect 6854 386 6857 387
rect 7031 387 7069 388
rect 7031 386 7034 387
rect 6854 356 6901 386
rect 6987 356 7034 386
rect 6854 355 6857 356
rect 6819 354 6857 355
rect 7031 355 7034 356
rect 7066 386 7069 387
rect 7267 387 7305 388
rect 7267 386 7270 387
rect 7066 356 7114 386
rect 7222 356 7270 386
rect 7066 355 7069 356
rect 7031 354 7069 355
rect 7267 355 7270 356
rect 7302 386 7305 387
rect 7479 387 7517 388
rect 7479 386 7482 387
rect 7302 356 7349 386
rect 7435 356 7482 386
rect 7302 355 7305 356
rect 7267 354 7305 355
rect 7479 355 7482 356
rect 7514 386 7517 387
rect 7715 387 7753 388
rect 7715 386 7718 387
rect 7514 356 7562 386
rect 7670 356 7718 386
rect 7514 355 7517 356
rect 7479 354 7517 355
rect 7715 355 7718 356
rect 7750 386 7753 387
rect 7927 387 7965 388
rect 7927 386 7930 387
rect 7750 356 7797 386
rect 7883 356 7930 386
rect 7750 355 7753 356
rect 7715 354 7753 355
rect 7927 355 7930 356
rect 7962 386 7965 387
rect 8163 387 8201 388
rect 8163 386 8166 387
rect 7962 356 8010 386
rect 8118 356 8166 386
rect 7962 355 7965 356
rect 7927 354 7965 355
rect 8163 355 8166 356
rect 8198 386 8201 387
rect 8375 387 8413 388
rect 8375 386 8378 387
rect 8198 356 8245 386
rect 8331 356 8378 386
rect 8198 355 8201 356
rect 8163 354 8201 355
rect 8375 355 8378 356
rect 8410 386 8413 387
rect 8611 387 8649 388
rect 8611 386 8614 387
rect 8410 356 8458 386
rect 8566 356 8614 386
rect 8410 355 8413 356
rect 8375 354 8413 355
rect 8611 355 8614 356
rect 8646 386 8649 387
rect 8823 387 8861 388
rect 8823 386 8826 387
rect 8646 356 8693 386
rect 8779 356 8826 386
rect 8646 355 8649 356
rect 8611 354 8649 355
rect 8823 355 8826 356
rect 8858 386 8861 387
rect 8858 356 8906 386
rect 8858 355 8861 356
rect 8823 354 8861 355
rect 196 325 252 328
rect 196 324 201 325
rect 35 294 201 324
rect 247 324 252 325
rect 644 325 700 328
rect 644 324 649 325
rect 247 294 413 324
rect 483 294 649 324
rect 695 324 700 325
rect 1092 325 1148 328
rect 1092 324 1097 325
rect 695 294 861 324
rect 931 294 1097 324
rect 1143 324 1148 325
rect 1540 325 1596 328
rect 1540 324 1545 325
rect 1143 294 1309 324
rect 1379 294 1545 324
rect 1591 324 1596 325
rect 1988 325 2044 328
rect 1988 324 1993 325
rect 1591 294 1757 324
rect 1827 294 1993 324
rect 2039 324 2044 325
rect 2436 325 2492 328
rect 2436 324 2441 325
rect 2039 294 2205 324
rect 2275 294 2441 324
rect 2487 324 2492 325
rect 2884 325 2940 328
rect 2884 324 2889 325
rect 2487 294 2653 324
rect 2723 294 2889 324
rect 2935 324 2940 325
rect 3332 325 3388 328
rect 3332 324 3337 325
rect 2935 294 3101 324
rect 3171 294 3337 324
rect 3383 324 3388 325
rect 3780 325 3836 328
rect 3780 324 3785 325
rect 3383 294 3549 324
rect 3619 294 3785 324
rect 3831 324 3836 325
rect 4228 325 4284 328
rect 4228 324 4233 325
rect 3831 294 3997 324
rect 4067 294 4233 324
rect 4279 324 4284 325
rect 4676 325 4732 328
rect 4676 324 4681 325
rect 4279 294 4445 324
rect 4515 294 4681 324
rect 4727 324 4732 325
rect 5124 325 5180 328
rect 5124 324 5129 325
rect 4727 294 4893 324
rect 4963 294 5129 324
rect 5175 324 5180 325
rect 5572 325 5628 328
rect 5572 324 5577 325
rect 5175 294 5341 324
rect 5411 294 5577 324
rect 5623 324 5628 325
rect 6020 325 6076 328
rect 6020 324 6025 325
rect 5623 294 5789 324
rect 5859 294 6025 324
rect 6071 324 6076 325
rect 6468 325 6524 328
rect 6468 324 6473 325
rect 6071 294 6237 324
rect 6307 294 6473 324
rect 6519 324 6524 325
rect 6916 325 6972 328
rect 6916 324 6921 325
rect 6519 294 6685 324
rect 6755 294 6921 324
rect 6967 324 6972 325
rect 7364 325 7420 328
rect 7364 324 7369 325
rect 6967 294 7133 324
rect 7203 294 7369 324
rect 7415 324 7420 325
rect 7812 325 7868 328
rect 7812 324 7817 325
rect 7415 294 7581 324
rect 7651 294 7817 324
rect 7863 324 7868 325
rect 8260 325 8316 328
rect 8260 324 8265 325
rect 7863 294 8029 324
rect 8099 294 8265 324
rect 8311 324 8316 325
rect 8708 325 8764 328
rect 8708 324 8713 325
rect 8311 294 8477 324
rect 8547 294 8713 324
rect 8759 324 8764 325
rect 8759 294 8925 324
rect 196 290 252 294
rect 644 290 700 294
rect 1092 290 1148 294
rect 1540 290 1596 294
rect 1988 290 2044 294
rect 2436 290 2492 294
rect 2884 290 2940 294
rect 3332 290 3388 294
rect 3780 290 3836 294
rect 4228 290 4284 294
rect 4676 290 4732 294
rect 5124 290 5180 294
rect 5572 290 5628 294
rect 6020 290 6076 294
rect 6468 290 6524 294
rect 6916 290 6972 294
rect 7364 290 7420 294
rect 7812 290 7868 294
rect 8260 290 8316 294
rect 8708 290 8764 294
rect 99 263 137 264
rect 99 262 102 263
rect 54 232 102 262
rect 99 231 102 232
rect 134 262 137 263
rect 311 263 349 264
rect 311 262 314 263
rect 134 232 181 262
rect 267 232 314 262
rect 134 231 137 232
rect 99 230 137 231
rect 311 231 314 232
rect 346 262 349 263
rect 547 263 585 264
rect 547 262 550 263
rect 346 232 394 262
rect 502 232 550 262
rect 346 231 349 232
rect 311 230 349 231
rect 547 231 550 232
rect 582 262 585 263
rect 759 263 797 264
rect 759 262 762 263
rect 582 232 629 262
rect 715 232 762 262
rect 582 231 585 232
rect 547 230 585 231
rect 759 231 762 232
rect 794 262 797 263
rect 995 263 1033 264
rect 995 262 998 263
rect 794 232 842 262
rect 950 232 998 262
rect 794 231 797 232
rect 759 230 797 231
rect 995 231 998 232
rect 1030 262 1033 263
rect 1207 263 1245 264
rect 1207 262 1210 263
rect 1030 232 1077 262
rect 1163 232 1210 262
rect 1030 231 1033 232
rect 995 230 1033 231
rect 1207 231 1210 232
rect 1242 262 1245 263
rect 1443 263 1481 264
rect 1443 262 1446 263
rect 1242 232 1290 262
rect 1398 232 1446 262
rect 1242 231 1245 232
rect 1207 230 1245 231
rect 1443 231 1446 232
rect 1478 262 1481 263
rect 1655 263 1693 264
rect 1655 262 1658 263
rect 1478 232 1525 262
rect 1611 232 1658 262
rect 1478 231 1481 232
rect 1443 230 1481 231
rect 1655 231 1658 232
rect 1690 262 1693 263
rect 1891 263 1929 264
rect 1891 262 1894 263
rect 1690 232 1738 262
rect 1846 232 1894 262
rect 1690 231 1693 232
rect 1655 230 1693 231
rect 1891 231 1894 232
rect 1926 262 1929 263
rect 2103 263 2141 264
rect 2103 262 2106 263
rect 1926 232 1973 262
rect 2059 232 2106 262
rect 1926 231 1929 232
rect 1891 230 1929 231
rect 2103 231 2106 232
rect 2138 262 2141 263
rect 2339 263 2377 264
rect 2339 262 2342 263
rect 2138 232 2186 262
rect 2294 232 2342 262
rect 2138 231 2141 232
rect 2103 230 2141 231
rect 2339 231 2342 232
rect 2374 262 2377 263
rect 2551 263 2589 264
rect 2551 262 2554 263
rect 2374 232 2421 262
rect 2507 232 2554 262
rect 2374 231 2377 232
rect 2339 230 2377 231
rect 2551 231 2554 232
rect 2586 262 2589 263
rect 2787 263 2825 264
rect 2787 262 2790 263
rect 2586 232 2634 262
rect 2742 232 2790 262
rect 2586 231 2589 232
rect 2551 230 2589 231
rect 2787 231 2790 232
rect 2822 262 2825 263
rect 2999 263 3037 264
rect 2999 262 3002 263
rect 2822 232 2869 262
rect 2955 232 3002 262
rect 2822 231 2825 232
rect 2787 230 2825 231
rect 2999 231 3002 232
rect 3034 262 3037 263
rect 3235 263 3273 264
rect 3235 262 3238 263
rect 3034 232 3082 262
rect 3190 232 3238 262
rect 3034 231 3037 232
rect 2999 230 3037 231
rect 3235 231 3238 232
rect 3270 262 3273 263
rect 3447 263 3485 264
rect 3447 262 3450 263
rect 3270 232 3317 262
rect 3403 232 3450 262
rect 3270 231 3273 232
rect 3235 230 3273 231
rect 3447 231 3450 232
rect 3482 262 3485 263
rect 3683 263 3721 264
rect 3683 262 3686 263
rect 3482 232 3530 262
rect 3638 232 3686 262
rect 3482 231 3485 232
rect 3447 230 3485 231
rect 3683 231 3686 232
rect 3718 262 3721 263
rect 3895 263 3933 264
rect 3895 262 3898 263
rect 3718 232 3765 262
rect 3851 232 3898 262
rect 3718 231 3721 232
rect 3683 230 3721 231
rect 3895 231 3898 232
rect 3930 262 3933 263
rect 4131 263 4169 264
rect 4131 262 4134 263
rect 3930 232 3978 262
rect 4086 232 4134 262
rect 3930 231 3933 232
rect 3895 230 3933 231
rect 4131 231 4134 232
rect 4166 262 4169 263
rect 4343 263 4381 264
rect 4343 262 4346 263
rect 4166 232 4213 262
rect 4299 232 4346 262
rect 4166 231 4169 232
rect 4131 230 4169 231
rect 4343 231 4346 232
rect 4378 262 4381 263
rect 4579 263 4617 264
rect 4579 262 4582 263
rect 4378 232 4426 262
rect 4534 232 4582 262
rect 4378 231 4381 232
rect 4343 230 4381 231
rect 4579 231 4582 232
rect 4614 262 4617 263
rect 4791 263 4829 264
rect 4791 262 4794 263
rect 4614 232 4661 262
rect 4747 232 4794 262
rect 4614 231 4617 232
rect 4579 230 4617 231
rect 4791 231 4794 232
rect 4826 262 4829 263
rect 5027 263 5065 264
rect 5027 262 5030 263
rect 4826 232 4874 262
rect 4982 232 5030 262
rect 4826 231 4829 232
rect 4791 230 4829 231
rect 5027 231 5030 232
rect 5062 262 5065 263
rect 5239 263 5277 264
rect 5239 262 5242 263
rect 5062 232 5109 262
rect 5195 232 5242 262
rect 5062 231 5065 232
rect 5027 230 5065 231
rect 5239 231 5242 232
rect 5274 262 5277 263
rect 5475 263 5513 264
rect 5475 262 5478 263
rect 5274 232 5322 262
rect 5430 232 5478 262
rect 5274 231 5277 232
rect 5239 230 5277 231
rect 5475 231 5478 232
rect 5510 262 5513 263
rect 5687 263 5725 264
rect 5687 262 5690 263
rect 5510 232 5557 262
rect 5643 232 5690 262
rect 5510 231 5513 232
rect 5475 230 5513 231
rect 5687 231 5690 232
rect 5722 262 5725 263
rect 5923 263 5961 264
rect 5923 262 5926 263
rect 5722 232 5770 262
rect 5878 232 5926 262
rect 5722 231 5725 232
rect 5687 230 5725 231
rect 5923 231 5926 232
rect 5958 262 5961 263
rect 6135 263 6173 264
rect 6135 262 6138 263
rect 5958 232 6005 262
rect 6091 232 6138 262
rect 5958 231 5961 232
rect 5923 230 5961 231
rect 6135 231 6138 232
rect 6170 262 6173 263
rect 6371 263 6409 264
rect 6371 262 6374 263
rect 6170 232 6218 262
rect 6326 232 6374 262
rect 6170 231 6173 232
rect 6135 230 6173 231
rect 6371 231 6374 232
rect 6406 262 6409 263
rect 6583 263 6621 264
rect 6583 262 6586 263
rect 6406 232 6453 262
rect 6539 232 6586 262
rect 6406 231 6409 232
rect 6371 230 6409 231
rect 6583 231 6586 232
rect 6618 262 6621 263
rect 6819 263 6857 264
rect 6819 262 6822 263
rect 6618 232 6666 262
rect 6774 232 6822 262
rect 6618 231 6621 232
rect 6583 230 6621 231
rect 6819 231 6822 232
rect 6854 262 6857 263
rect 7031 263 7069 264
rect 7031 262 7034 263
rect 6854 232 6901 262
rect 6987 232 7034 262
rect 6854 231 6857 232
rect 6819 230 6857 231
rect 7031 231 7034 232
rect 7066 262 7069 263
rect 7267 263 7305 264
rect 7267 262 7270 263
rect 7066 232 7114 262
rect 7222 232 7270 262
rect 7066 231 7069 232
rect 7031 230 7069 231
rect 7267 231 7270 232
rect 7302 262 7305 263
rect 7479 263 7517 264
rect 7479 262 7482 263
rect 7302 232 7349 262
rect 7435 232 7482 262
rect 7302 231 7305 232
rect 7267 230 7305 231
rect 7479 231 7482 232
rect 7514 262 7517 263
rect 7715 263 7753 264
rect 7715 262 7718 263
rect 7514 232 7562 262
rect 7670 232 7718 262
rect 7514 231 7517 232
rect 7479 230 7517 231
rect 7715 231 7718 232
rect 7750 262 7753 263
rect 7927 263 7965 264
rect 7927 262 7930 263
rect 7750 232 7797 262
rect 7883 232 7930 262
rect 7750 231 7753 232
rect 7715 230 7753 231
rect 7927 231 7930 232
rect 7962 262 7965 263
rect 8163 263 8201 264
rect 8163 262 8166 263
rect 7962 232 8010 262
rect 8118 232 8166 262
rect 7962 231 7965 232
rect 7927 230 7965 231
rect 8163 231 8166 232
rect 8198 262 8201 263
rect 8375 263 8413 264
rect 8375 262 8378 263
rect 8198 232 8245 262
rect 8331 232 8378 262
rect 8198 231 8201 232
rect 8163 230 8201 231
rect 8375 231 8378 232
rect 8410 262 8413 263
rect 8611 263 8649 264
rect 8611 262 8614 263
rect 8410 232 8458 262
rect 8566 232 8614 262
rect 8410 231 8413 232
rect 8375 230 8413 231
rect 8611 231 8614 232
rect 8646 262 8649 263
rect 8823 263 8861 264
rect 8823 262 8826 263
rect 8646 232 8693 262
rect 8779 232 8826 262
rect 8646 231 8649 232
rect 8611 230 8649 231
rect 8823 231 8826 232
rect 8858 262 8861 263
rect 8858 232 8906 262
rect 8858 231 8861 232
rect 8823 230 8861 231
rect 196 201 252 204
rect 196 200 201 201
rect 35 170 201 200
rect 247 200 252 201
rect 644 201 700 204
rect 644 200 649 201
rect 247 170 413 200
rect 483 170 649 200
rect 695 200 700 201
rect 1092 201 1148 204
rect 1092 200 1097 201
rect 695 170 861 200
rect 931 170 1097 200
rect 1143 200 1148 201
rect 1540 201 1596 204
rect 1540 200 1545 201
rect 1143 170 1309 200
rect 1379 170 1545 200
rect 1591 200 1596 201
rect 1988 201 2044 204
rect 1988 200 1993 201
rect 1591 170 1757 200
rect 1827 170 1993 200
rect 2039 200 2044 201
rect 2436 201 2492 204
rect 2436 200 2441 201
rect 2039 170 2205 200
rect 2275 170 2441 200
rect 2487 200 2492 201
rect 2884 201 2940 204
rect 2884 200 2889 201
rect 2487 170 2653 200
rect 2723 170 2889 200
rect 2935 200 2940 201
rect 3332 201 3388 204
rect 3332 200 3337 201
rect 2935 170 3101 200
rect 3171 170 3337 200
rect 3383 200 3388 201
rect 3780 201 3836 204
rect 3780 200 3785 201
rect 3383 170 3549 200
rect 3619 170 3785 200
rect 3831 200 3836 201
rect 4228 201 4284 204
rect 4228 200 4233 201
rect 3831 170 3997 200
rect 4067 170 4233 200
rect 4279 200 4284 201
rect 4676 201 4732 204
rect 4676 200 4681 201
rect 4279 170 4445 200
rect 4515 170 4681 200
rect 4727 200 4732 201
rect 5124 201 5180 204
rect 5124 200 5129 201
rect 4727 170 4893 200
rect 4963 170 5129 200
rect 5175 200 5180 201
rect 5572 201 5628 204
rect 5572 200 5577 201
rect 5175 170 5341 200
rect 5411 170 5577 200
rect 5623 200 5628 201
rect 6020 201 6076 204
rect 6020 200 6025 201
rect 5623 170 5789 200
rect 5859 170 6025 200
rect 6071 200 6076 201
rect 6468 201 6524 204
rect 6468 200 6473 201
rect 6071 170 6237 200
rect 6307 170 6473 200
rect 6519 200 6524 201
rect 6916 201 6972 204
rect 6916 200 6921 201
rect 6519 170 6685 200
rect 6755 170 6921 200
rect 6967 200 6972 201
rect 7364 201 7420 204
rect 7364 200 7369 201
rect 6967 170 7133 200
rect 7203 170 7369 200
rect 7415 200 7420 201
rect 7812 201 7868 204
rect 7812 200 7817 201
rect 7415 170 7581 200
rect 7651 170 7817 200
rect 7863 200 7868 201
rect 8260 201 8316 204
rect 8260 200 8265 201
rect 7863 170 8029 200
rect 8099 170 8265 200
rect 8311 200 8316 201
rect 8708 201 8764 204
rect 8708 200 8713 201
rect 8311 170 8477 200
rect 8547 170 8713 200
rect 8759 200 8764 201
rect 8759 170 8925 200
rect 196 166 252 170
rect 644 166 700 170
rect 1092 166 1148 170
rect 1540 166 1596 170
rect 1988 166 2044 170
rect 2436 166 2492 170
rect 2884 166 2940 170
rect 3332 166 3388 170
rect 3780 166 3836 170
rect 4228 166 4284 170
rect 4676 166 4732 170
rect 5124 166 5180 170
rect 5572 166 5628 170
rect 6020 166 6076 170
rect 6468 166 6524 170
rect 6916 166 6972 170
rect 7364 166 7420 170
rect 7812 166 7868 170
rect 8260 166 8316 170
rect 8708 166 8764 170
rect 99 139 137 140
rect 99 138 102 139
rect 54 108 102 138
rect 99 107 102 108
rect 134 138 137 139
rect 311 139 349 140
rect 311 138 314 139
rect 134 108 181 138
rect 267 108 314 138
rect 134 107 137 108
rect 99 106 137 107
rect 311 107 314 108
rect 346 138 349 139
rect 547 139 585 140
rect 547 138 550 139
rect 346 108 394 138
rect 502 108 550 138
rect 346 107 349 108
rect 311 106 349 107
rect 547 107 550 108
rect 582 138 585 139
rect 759 139 797 140
rect 759 138 762 139
rect 582 108 629 138
rect 715 108 762 138
rect 582 107 585 108
rect 547 106 585 107
rect 759 107 762 108
rect 794 138 797 139
rect 995 139 1033 140
rect 995 138 998 139
rect 794 108 842 138
rect 950 108 998 138
rect 794 107 797 108
rect 759 106 797 107
rect 995 107 998 108
rect 1030 138 1033 139
rect 1207 139 1245 140
rect 1207 138 1210 139
rect 1030 108 1077 138
rect 1163 108 1210 138
rect 1030 107 1033 108
rect 995 106 1033 107
rect 1207 107 1210 108
rect 1242 138 1245 139
rect 1443 139 1481 140
rect 1443 138 1446 139
rect 1242 108 1290 138
rect 1398 108 1446 138
rect 1242 107 1245 108
rect 1207 106 1245 107
rect 1443 107 1446 108
rect 1478 138 1481 139
rect 1655 139 1693 140
rect 1655 138 1658 139
rect 1478 108 1525 138
rect 1611 108 1658 138
rect 1478 107 1481 108
rect 1443 106 1481 107
rect 1655 107 1658 108
rect 1690 138 1693 139
rect 1891 139 1929 140
rect 1891 138 1894 139
rect 1690 108 1738 138
rect 1846 108 1894 138
rect 1690 107 1693 108
rect 1655 106 1693 107
rect 1891 107 1894 108
rect 1926 138 1929 139
rect 2103 139 2141 140
rect 2103 138 2106 139
rect 1926 108 1973 138
rect 2059 108 2106 138
rect 1926 107 1929 108
rect 1891 106 1929 107
rect 2103 107 2106 108
rect 2138 138 2141 139
rect 2339 139 2377 140
rect 2339 138 2342 139
rect 2138 108 2186 138
rect 2294 108 2342 138
rect 2138 107 2141 108
rect 2103 106 2141 107
rect 2339 107 2342 108
rect 2374 138 2377 139
rect 2551 139 2589 140
rect 2551 138 2554 139
rect 2374 108 2421 138
rect 2507 108 2554 138
rect 2374 107 2377 108
rect 2339 106 2377 107
rect 2551 107 2554 108
rect 2586 138 2589 139
rect 2787 139 2825 140
rect 2787 138 2790 139
rect 2586 108 2634 138
rect 2742 108 2790 138
rect 2586 107 2589 108
rect 2551 106 2589 107
rect 2787 107 2790 108
rect 2822 138 2825 139
rect 2999 139 3037 140
rect 2999 138 3002 139
rect 2822 108 2869 138
rect 2955 108 3002 138
rect 2822 107 2825 108
rect 2787 106 2825 107
rect 2999 107 3002 108
rect 3034 138 3037 139
rect 3235 139 3273 140
rect 3235 138 3238 139
rect 3034 108 3082 138
rect 3190 108 3238 138
rect 3034 107 3037 108
rect 2999 106 3037 107
rect 3235 107 3238 108
rect 3270 138 3273 139
rect 3447 139 3485 140
rect 3447 138 3450 139
rect 3270 108 3317 138
rect 3403 108 3450 138
rect 3270 107 3273 108
rect 3235 106 3273 107
rect 3447 107 3450 108
rect 3482 138 3485 139
rect 3683 139 3721 140
rect 3683 138 3686 139
rect 3482 108 3530 138
rect 3638 108 3686 138
rect 3482 107 3485 108
rect 3447 106 3485 107
rect 3683 107 3686 108
rect 3718 138 3721 139
rect 3895 139 3933 140
rect 3895 138 3898 139
rect 3718 108 3765 138
rect 3851 108 3898 138
rect 3718 107 3721 108
rect 3683 106 3721 107
rect 3895 107 3898 108
rect 3930 138 3933 139
rect 4131 139 4169 140
rect 4131 138 4134 139
rect 3930 108 3978 138
rect 4086 108 4134 138
rect 3930 107 3933 108
rect 3895 106 3933 107
rect 4131 107 4134 108
rect 4166 138 4169 139
rect 4343 139 4381 140
rect 4343 138 4346 139
rect 4166 108 4213 138
rect 4299 108 4346 138
rect 4166 107 4169 108
rect 4131 106 4169 107
rect 4343 107 4346 108
rect 4378 138 4381 139
rect 4579 139 4617 140
rect 4579 138 4582 139
rect 4378 108 4426 138
rect 4534 108 4582 138
rect 4378 107 4381 108
rect 4343 106 4381 107
rect 4579 107 4582 108
rect 4614 138 4617 139
rect 4791 139 4829 140
rect 4791 138 4794 139
rect 4614 108 4661 138
rect 4747 108 4794 138
rect 4614 107 4617 108
rect 4579 106 4617 107
rect 4791 107 4794 108
rect 4826 138 4829 139
rect 5027 139 5065 140
rect 5027 138 5030 139
rect 4826 108 4874 138
rect 4982 108 5030 138
rect 4826 107 4829 108
rect 4791 106 4829 107
rect 5027 107 5030 108
rect 5062 138 5065 139
rect 5239 139 5277 140
rect 5239 138 5242 139
rect 5062 108 5109 138
rect 5195 108 5242 138
rect 5062 107 5065 108
rect 5027 106 5065 107
rect 5239 107 5242 108
rect 5274 138 5277 139
rect 5475 139 5513 140
rect 5475 138 5478 139
rect 5274 108 5322 138
rect 5430 108 5478 138
rect 5274 107 5277 108
rect 5239 106 5277 107
rect 5475 107 5478 108
rect 5510 138 5513 139
rect 5687 139 5725 140
rect 5687 138 5690 139
rect 5510 108 5557 138
rect 5643 108 5690 138
rect 5510 107 5513 108
rect 5475 106 5513 107
rect 5687 107 5690 108
rect 5722 138 5725 139
rect 5923 139 5961 140
rect 5923 138 5926 139
rect 5722 108 5770 138
rect 5878 108 5926 138
rect 5722 107 5725 108
rect 5687 106 5725 107
rect 5923 107 5926 108
rect 5958 138 5961 139
rect 6135 139 6173 140
rect 6135 138 6138 139
rect 5958 108 6005 138
rect 6091 108 6138 138
rect 5958 107 5961 108
rect 5923 106 5961 107
rect 6135 107 6138 108
rect 6170 138 6173 139
rect 6371 139 6409 140
rect 6371 138 6374 139
rect 6170 108 6218 138
rect 6326 108 6374 138
rect 6170 107 6173 108
rect 6135 106 6173 107
rect 6371 107 6374 108
rect 6406 138 6409 139
rect 6583 139 6621 140
rect 6583 138 6586 139
rect 6406 108 6453 138
rect 6539 108 6586 138
rect 6406 107 6409 108
rect 6371 106 6409 107
rect 6583 107 6586 108
rect 6618 138 6621 139
rect 6819 139 6857 140
rect 6819 138 6822 139
rect 6618 108 6666 138
rect 6774 108 6822 138
rect 6618 107 6621 108
rect 6583 106 6621 107
rect 6819 107 6822 108
rect 6854 138 6857 139
rect 7031 139 7069 140
rect 7031 138 7034 139
rect 6854 108 6901 138
rect 6987 108 7034 138
rect 6854 107 6857 108
rect 6819 106 6857 107
rect 7031 107 7034 108
rect 7066 138 7069 139
rect 7267 139 7305 140
rect 7267 138 7270 139
rect 7066 108 7114 138
rect 7222 108 7270 138
rect 7066 107 7069 108
rect 7031 106 7069 107
rect 7267 107 7270 108
rect 7302 138 7305 139
rect 7479 139 7517 140
rect 7479 138 7482 139
rect 7302 108 7349 138
rect 7435 108 7482 138
rect 7302 107 7305 108
rect 7267 106 7305 107
rect 7479 107 7482 108
rect 7514 138 7517 139
rect 7715 139 7753 140
rect 7715 138 7718 139
rect 7514 108 7562 138
rect 7670 108 7718 138
rect 7514 107 7517 108
rect 7479 106 7517 107
rect 7715 107 7718 108
rect 7750 138 7753 139
rect 7927 139 7965 140
rect 7927 138 7930 139
rect 7750 108 7797 138
rect 7883 108 7930 138
rect 7750 107 7753 108
rect 7715 106 7753 107
rect 7927 107 7930 108
rect 7962 138 7965 139
rect 8163 139 8201 140
rect 8163 138 8166 139
rect 7962 108 8010 138
rect 8118 108 8166 138
rect 7962 107 7965 108
rect 7927 106 7965 107
rect 8163 107 8166 108
rect 8198 138 8201 139
rect 8375 139 8413 140
rect 8375 138 8378 139
rect 8198 108 8245 138
rect 8331 108 8378 138
rect 8198 107 8201 108
rect 8163 106 8201 107
rect 8375 107 8378 108
rect 8410 138 8413 139
rect 8611 139 8649 140
rect 8611 138 8614 139
rect 8410 108 8458 138
rect 8566 108 8614 138
rect 8410 107 8413 108
rect 8375 106 8413 107
rect 8611 107 8614 108
rect 8646 138 8649 139
rect 8823 139 8861 140
rect 8823 138 8826 139
rect 8646 108 8693 138
rect 8779 108 8826 138
rect 8646 107 8649 108
rect 8611 106 8649 107
rect 8823 107 8826 108
rect 8858 138 8861 139
rect 8858 108 8906 138
rect 8858 107 8861 108
rect 8823 106 8861 107
rect 196 77 252 80
rect 196 76 201 77
rect 35 46 201 76
rect 247 76 252 77
rect 644 77 700 80
rect 644 76 649 77
rect 247 46 413 76
rect 483 46 649 76
rect 695 76 700 77
rect 1092 77 1148 80
rect 1092 76 1097 77
rect 695 46 861 76
rect 931 46 1097 76
rect 1143 76 1148 77
rect 1540 77 1596 80
rect 1540 76 1545 77
rect 1143 46 1309 76
rect 1379 46 1545 76
rect 1591 76 1596 77
rect 1988 77 2044 80
rect 1988 76 1993 77
rect 1591 46 1757 76
rect 1827 46 1993 76
rect 2039 76 2044 77
rect 2436 77 2492 80
rect 2436 76 2441 77
rect 2039 46 2205 76
rect 2275 46 2441 76
rect 2487 76 2492 77
rect 2884 77 2940 80
rect 2884 76 2889 77
rect 2487 46 2653 76
rect 2723 46 2889 76
rect 2935 76 2940 77
rect 3332 77 3388 80
rect 3332 76 3337 77
rect 2935 46 3101 76
rect 3171 46 3337 76
rect 3383 76 3388 77
rect 3780 77 3836 80
rect 3780 76 3785 77
rect 3383 46 3549 76
rect 3619 46 3785 76
rect 3831 76 3836 77
rect 4228 77 4284 80
rect 4228 76 4233 77
rect 3831 46 3997 76
rect 4067 46 4233 76
rect 4279 76 4284 77
rect 4676 77 4732 80
rect 4676 76 4681 77
rect 4279 46 4445 76
rect 4515 46 4681 76
rect 4727 76 4732 77
rect 5124 77 5180 80
rect 5124 76 5129 77
rect 4727 46 4893 76
rect 4963 46 5129 76
rect 5175 76 5180 77
rect 5572 77 5628 80
rect 5572 76 5577 77
rect 5175 46 5341 76
rect 5411 46 5577 76
rect 5623 76 5628 77
rect 6020 77 6076 80
rect 6020 76 6025 77
rect 5623 46 5789 76
rect 5859 46 6025 76
rect 6071 76 6076 77
rect 6468 77 6524 80
rect 6468 76 6473 77
rect 6071 46 6237 76
rect 6307 46 6473 76
rect 6519 76 6524 77
rect 6916 77 6972 80
rect 6916 76 6921 77
rect 6519 46 6685 76
rect 6755 46 6921 76
rect 6967 76 6972 77
rect 7364 77 7420 80
rect 7364 76 7369 77
rect 6967 46 7133 76
rect 7203 46 7369 76
rect 7415 76 7420 77
rect 7812 77 7868 80
rect 7812 76 7817 77
rect 7415 46 7581 76
rect 7651 46 7817 76
rect 7863 76 7868 77
rect 8260 77 8316 80
rect 8260 76 8265 77
rect 7863 46 8029 76
rect 8099 46 8265 76
rect 8311 76 8316 77
rect 8708 77 8764 80
rect 8708 76 8713 77
rect 8311 46 8477 76
rect 8547 46 8713 76
rect 8759 76 8764 77
rect 8759 46 8925 76
rect 196 42 252 46
rect 644 42 700 46
rect 1092 42 1148 46
rect 1540 42 1596 46
rect 1988 42 2044 46
rect 2436 42 2492 46
rect 2884 42 2940 46
rect 3332 42 3388 46
rect 3780 42 3836 46
rect 4228 42 4284 46
rect 4676 42 4732 46
rect 5124 42 5180 46
rect 5572 42 5628 46
rect 6020 42 6076 46
rect 6468 42 6524 46
rect 6916 42 6972 46
rect 7364 42 7420 46
rect 7812 42 7868 46
rect 8260 42 8316 46
rect 8708 42 8764 46
<< via3 >>
rect 102 2336 134 2368
rect 314 2336 346 2368
rect 550 2336 582 2368
rect 762 2336 794 2368
rect 998 2336 1030 2368
rect 1210 2336 1242 2368
rect 1446 2336 1478 2368
rect 1658 2336 1690 2368
rect 1894 2336 1926 2368
rect 2106 2336 2138 2368
rect 2342 2336 2374 2368
rect 2554 2336 2586 2368
rect 2790 2336 2822 2368
rect 3002 2336 3034 2368
rect 3238 2336 3270 2368
rect 3450 2336 3482 2368
rect 3686 2336 3718 2368
rect 3898 2336 3930 2368
rect 4134 2336 4166 2368
rect 4346 2336 4378 2368
rect 4582 2336 4614 2368
rect 4794 2336 4826 2368
rect 5030 2336 5062 2368
rect 5242 2336 5274 2368
rect 5478 2336 5510 2368
rect 5690 2336 5722 2368
rect 5926 2336 5958 2368
rect 6138 2336 6170 2368
rect 6374 2336 6406 2368
rect 6586 2336 6618 2368
rect 6822 2336 6854 2368
rect 7034 2336 7066 2368
rect 7270 2336 7302 2368
rect 7482 2336 7514 2368
rect 7718 2336 7750 2368
rect 7930 2336 7962 2368
rect 8166 2336 8198 2368
rect 8378 2336 8410 2368
rect 8614 2336 8646 2368
rect 8826 2336 8858 2368
rect 102 2212 134 2244
rect 314 2212 346 2244
rect 550 2212 582 2244
rect 762 2212 794 2244
rect 998 2212 1030 2244
rect 1210 2212 1242 2244
rect 1446 2212 1478 2244
rect 1658 2212 1690 2244
rect 1894 2212 1926 2244
rect 2106 2212 2138 2244
rect 2342 2212 2374 2244
rect 2554 2212 2586 2244
rect 2790 2212 2822 2244
rect 3002 2212 3034 2244
rect 3238 2212 3270 2244
rect 3450 2212 3482 2244
rect 3686 2212 3718 2244
rect 3898 2212 3930 2244
rect 4134 2212 4166 2244
rect 4346 2212 4378 2244
rect 4582 2212 4614 2244
rect 4794 2212 4826 2244
rect 5030 2212 5062 2244
rect 5242 2212 5274 2244
rect 5478 2212 5510 2244
rect 5690 2212 5722 2244
rect 5926 2212 5958 2244
rect 6138 2212 6170 2244
rect 6374 2212 6406 2244
rect 6586 2212 6618 2244
rect 6822 2212 6854 2244
rect 7034 2212 7066 2244
rect 7270 2212 7302 2244
rect 7482 2212 7514 2244
rect 7718 2212 7750 2244
rect 7930 2212 7962 2244
rect 8166 2212 8198 2244
rect 8378 2212 8410 2244
rect 8614 2212 8646 2244
rect 8826 2212 8858 2244
rect 102 2088 134 2120
rect 314 2088 346 2120
rect 550 2088 582 2120
rect 762 2088 794 2120
rect 998 2088 1030 2120
rect 1210 2088 1242 2120
rect 1446 2088 1478 2120
rect 1658 2088 1690 2120
rect 1894 2088 1926 2120
rect 2106 2088 2138 2120
rect 2342 2088 2374 2120
rect 2554 2088 2586 2120
rect 2790 2088 2822 2120
rect 3002 2088 3034 2120
rect 3238 2088 3270 2120
rect 3450 2088 3482 2120
rect 3686 2088 3718 2120
rect 3898 2088 3930 2120
rect 4134 2088 4166 2120
rect 4346 2088 4378 2120
rect 4582 2088 4614 2120
rect 4794 2088 4826 2120
rect 5030 2088 5062 2120
rect 5242 2088 5274 2120
rect 5478 2088 5510 2120
rect 5690 2088 5722 2120
rect 5926 2088 5958 2120
rect 6138 2088 6170 2120
rect 6374 2088 6406 2120
rect 6586 2088 6618 2120
rect 6822 2088 6854 2120
rect 7034 2088 7066 2120
rect 7270 2088 7302 2120
rect 7482 2088 7514 2120
rect 7718 2088 7750 2120
rect 7930 2088 7962 2120
rect 8166 2088 8198 2120
rect 8378 2088 8410 2120
rect 8614 2088 8646 2120
rect 8826 2088 8858 2120
rect 102 1964 134 1996
rect 314 1964 346 1996
rect 550 1964 582 1996
rect 762 1964 794 1996
rect 998 1964 1030 1996
rect 1210 1964 1242 1996
rect 1446 1964 1478 1996
rect 1658 1964 1690 1996
rect 1894 1964 1926 1996
rect 2106 1964 2138 1996
rect 2342 1964 2374 1996
rect 2554 1964 2586 1996
rect 2790 1964 2822 1996
rect 3002 1964 3034 1996
rect 3238 1964 3270 1996
rect 3450 1964 3482 1996
rect 3686 1964 3718 1996
rect 3898 1964 3930 1996
rect 4134 1964 4166 1996
rect 4346 1964 4378 1996
rect 4582 1964 4614 1996
rect 4794 1964 4826 1996
rect 5030 1964 5062 1996
rect 5242 1964 5274 1996
rect 5478 1964 5510 1996
rect 5690 1964 5722 1996
rect 5926 1964 5958 1996
rect 6138 1964 6170 1996
rect 6374 1964 6406 1996
rect 6586 1964 6618 1996
rect 6822 1964 6854 1996
rect 7034 1964 7066 1996
rect 7270 1964 7302 1996
rect 7482 1964 7514 1996
rect 7718 1964 7750 1996
rect 7930 1964 7962 1996
rect 8166 1964 8198 1996
rect 8378 1964 8410 1996
rect 8614 1964 8646 1996
rect 8826 1964 8858 1996
rect 102 1717 134 1749
rect 314 1717 346 1749
rect 550 1717 582 1749
rect 762 1717 794 1749
rect 998 1717 1030 1749
rect 1210 1717 1242 1749
rect 1446 1717 1478 1749
rect 1658 1717 1690 1749
rect 1894 1717 1926 1749
rect 2106 1717 2138 1749
rect 2342 1717 2374 1749
rect 2554 1717 2586 1749
rect 2790 1717 2822 1749
rect 3002 1717 3034 1749
rect 3238 1717 3270 1749
rect 3450 1717 3482 1749
rect 3686 1717 3718 1749
rect 3898 1717 3930 1749
rect 4134 1717 4166 1749
rect 4346 1717 4378 1749
rect 4582 1717 4614 1749
rect 4794 1717 4826 1749
rect 5030 1717 5062 1749
rect 5242 1717 5274 1749
rect 5478 1717 5510 1749
rect 5690 1717 5722 1749
rect 5926 1717 5958 1749
rect 6138 1717 6170 1749
rect 6374 1717 6406 1749
rect 6586 1717 6618 1749
rect 6822 1717 6854 1749
rect 7034 1717 7066 1749
rect 7270 1717 7302 1749
rect 7482 1717 7514 1749
rect 7718 1717 7750 1749
rect 7930 1717 7962 1749
rect 8166 1717 8198 1749
rect 8378 1717 8410 1749
rect 8614 1717 8646 1749
rect 8826 1717 8858 1749
rect 102 1593 134 1625
rect 314 1593 346 1625
rect 550 1593 582 1625
rect 762 1593 794 1625
rect 998 1593 1030 1625
rect 1210 1593 1242 1625
rect 1446 1593 1478 1625
rect 1658 1593 1690 1625
rect 1894 1593 1926 1625
rect 2106 1593 2138 1625
rect 2342 1593 2374 1625
rect 2554 1593 2586 1625
rect 2790 1593 2822 1625
rect 3002 1593 3034 1625
rect 3238 1593 3270 1625
rect 3450 1593 3482 1625
rect 3686 1593 3718 1625
rect 3898 1593 3930 1625
rect 4134 1593 4166 1625
rect 4346 1593 4378 1625
rect 4582 1593 4614 1625
rect 4794 1593 4826 1625
rect 5030 1593 5062 1625
rect 5242 1593 5274 1625
rect 5478 1593 5510 1625
rect 5690 1593 5722 1625
rect 5926 1593 5958 1625
rect 6138 1593 6170 1625
rect 6374 1593 6406 1625
rect 6586 1593 6618 1625
rect 6822 1593 6854 1625
rect 7034 1593 7066 1625
rect 7270 1593 7302 1625
rect 7482 1593 7514 1625
rect 7718 1593 7750 1625
rect 7930 1593 7962 1625
rect 8166 1593 8198 1625
rect 8378 1593 8410 1625
rect 8614 1593 8646 1625
rect 8826 1593 8858 1625
rect 102 1469 134 1501
rect 314 1469 346 1501
rect 550 1469 582 1501
rect 762 1469 794 1501
rect 998 1469 1030 1501
rect 1210 1469 1242 1501
rect 1446 1469 1478 1501
rect 1658 1469 1690 1501
rect 1894 1469 1926 1501
rect 2106 1469 2138 1501
rect 2342 1469 2374 1501
rect 2554 1469 2586 1501
rect 2790 1469 2822 1501
rect 3002 1469 3034 1501
rect 3238 1469 3270 1501
rect 3450 1469 3482 1501
rect 3686 1469 3718 1501
rect 3898 1469 3930 1501
rect 4134 1469 4166 1501
rect 4346 1469 4378 1501
rect 4582 1469 4614 1501
rect 4794 1469 4826 1501
rect 5030 1469 5062 1501
rect 5242 1469 5274 1501
rect 5478 1469 5510 1501
rect 5690 1469 5722 1501
rect 5926 1469 5958 1501
rect 6138 1469 6170 1501
rect 6374 1469 6406 1501
rect 6586 1469 6618 1501
rect 6822 1469 6854 1501
rect 7034 1469 7066 1501
rect 7270 1469 7302 1501
rect 7482 1469 7514 1501
rect 7718 1469 7750 1501
rect 7930 1469 7962 1501
rect 8166 1469 8198 1501
rect 8378 1469 8410 1501
rect 8614 1469 8646 1501
rect 8826 1469 8858 1501
rect 102 1345 134 1377
rect 314 1345 346 1377
rect 550 1345 582 1377
rect 762 1345 794 1377
rect 998 1345 1030 1377
rect 1210 1345 1242 1377
rect 1446 1345 1478 1377
rect 1658 1345 1690 1377
rect 1894 1345 1926 1377
rect 2106 1345 2138 1377
rect 2342 1345 2374 1377
rect 2554 1345 2586 1377
rect 2790 1345 2822 1377
rect 3002 1345 3034 1377
rect 3238 1345 3270 1377
rect 3450 1345 3482 1377
rect 3686 1345 3718 1377
rect 3898 1345 3930 1377
rect 4134 1345 4166 1377
rect 4346 1345 4378 1377
rect 4582 1345 4614 1377
rect 4794 1345 4826 1377
rect 5030 1345 5062 1377
rect 5242 1345 5274 1377
rect 5478 1345 5510 1377
rect 5690 1345 5722 1377
rect 5926 1345 5958 1377
rect 6138 1345 6170 1377
rect 6374 1345 6406 1377
rect 6586 1345 6618 1377
rect 6822 1345 6854 1377
rect 7034 1345 7066 1377
rect 7270 1345 7302 1377
rect 7482 1345 7514 1377
rect 7718 1345 7750 1377
rect 7930 1345 7962 1377
rect 8166 1345 8198 1377
rect 8378 1345 8410 1377
rect 8614 1345 8646 1377
rect 8826 1345 8858 1377
rect 102 1098 134 1130
rect 314 1098 346 1130
rect 550 1098 582 1130
rect 762 1098 794 1130
rect 998 1098 1030 1130
rect 1210 1098 1242 1130
rect 1446 1098 1478 1130
rect 1658 1098 1690 1130
rect 1894 1098 1926 1130
rect 2106 1098 2138 1130
rect 2342 1098 2374 1130
rect 2554 1098 2586 1130
rect 2790 1098 2822 1130
rect 3002 1098 3034 1130
rect 3238 1098 3270 1130
rect 3450 1098 3482 1130
rect 3686 1098 3718 1130
rect 3898 1098 3930 1130
rect 4134 1098 4166 1130
rect 4346 1098 4378 1130
rect 4582 1098 4614 1130
rect 4794 1098 4826 1130
rect 5030 1098 5062 1130
rect 5242 1098 5274 1130
rect 5478 1098 5510 1130
rect 5690 1098 5722 1130
rect 5926 1098 5958 1130
rect 6138 1098 6170 1130
rect 6374 1098 6406 1130
rect 6586 1098 6618 1130
rect 6822 1098 6854 1130
rect 7034 1098 7066 1130
rect 7270 1098 7302 1130
rect 7482 1098 7514 1130
rect 7718 1098 7750 1130
rect 7930 1098 7962 1130
rect 8166 1098 8198 1130
rect 8378 1098 8410 1130
rect 8614 1098 8646 1130
rect 8826 1098 8858 1130
rect 102 974 134 1006
rect 314 974 346 1006
rect 550 974 582 1006
rect 762 974 794 1006
rect 998 974 1030 1006
rect 1210 974 1242 1006
rect 1446 974 1478 1006
rect 1658 974 1690 1006
rect 1894 974 1926 1006
rect 2106 974 2138 1006
rect 2342 974 2374 1006
rect 2554 974 2586 1006
rect 2790 974 2822 1006
rect 3002 974 3034 1006
rect 3238 974 3270 1006
rect 3450 974 3482 1006
rect 3686 974 3718 1006
rect 3898 974 3930 1006
rect 4134 974 4166 1006
rect 4346 974 4378 1006
rect 4582 974 4614 1006
rect 4794 974 4826 1006
rect 5030 974 5062 1006
rect 5242 974 5274 1006
rect 5478 974 5510 1006
rect 5690 974 5722 1006
rect 5926 974 5958 1006
rect 6138 974 6170 1006
rect 6374 974 6406 1006
rect 6586 974 6618 1006
rect 6822 974 6854 1006
rect 7034 974 7066 1006
rect 7270 974 7302 1006
rect 7482 974 7514 1006
rect 7718 974 7750 1006
rect 7930 974 7962 1006
rect 8166 974 8198 1006
rect 8378 974 8410 1006
rect 8614 974 8646 1006
rect 8826 974 8858 1006
rect 102 850 134 882
rect 314 850 346 882
rect 550 850 582 882
rect 762 850 794 882
rect 998 850 1030 882
rect 1210 850 1242 882
rect 1446 850 1478 882
rect 1658 850 1690 882
rect 1894 850 1926 882
rect 2106 850 2138 882
rect 2342 850 2374 882
rect 2554 850 2586 882
rect 2790 850 2822 882
rect 3002 850 3034 882
rect 3238 850 3270 882
rect 3450 850 3482 882
rect 3686 850 3718 882
rect 3898 850 3930 882
rect 4134 850 4166 882
rect 4346 850 4378 882
rect 4582 850 4614 882
rect 4794 850 4826 882
rect 5030 850 5062 882
rect 5242 850 5274 882
rect 5478 850 5510 882
rect 5690 850 5722 882
rect 5926 850 5958 882
rect 6138 850 6170 882
rect 6374 850 6406 882
rect 6586 850 6618 882
rect 6822 850 6854 882
rect 7034 850 7066 882
rect 7270 850 7302 882
rect 7482 850 7514 882
rect 7718 850 7750 882
rect 7930 850 7962 882
rect 8166 850 8198 882
rect 8378 850 8410 882
rect 8614 850 8646 882
rect 8826 850 8858 882
rect 102 726 134 758
rect 314 726 346 758
rect 550 726 582 758
rect 762 726 794 758
rect 998 726 1030 758
rect 1210 726 1242 758
rect 1446 726 1478 758
rect 1658 726 1690 758
rect 1894 726 1926 758
rect 2106 726 2138 758
rect 2342 726 2374 758
rect 2554 726 2586 758
rect 2790 726 2822 758
rect 3002 726 3034 758
rect 3238 726 3270 758
rect 3450 726 3482 758
rect 3686 726 3718 758
rect 3898 726 3930 758
rect 4134 726 4166 758
rect 4346 726 4378 758
rect 4582 726 4614 758
rect 4794 726 4826 758
rect 5030 726 5062 758
rect 5242 726 5274 758
rect 5478 726 5510 758
rect 5690 726 5722 758
rect 5926 726 5958 758
rect 6138 726 6170 758
rect 6374 726 6406 758
rect 6586 726 6618 758
rect 6822 726 6854 758
rect 7034 726 7066 758
rect 7270 726 7302 758
rect 7482 726 7514 758
rect 7718 726 7750 758
rect 7930 726 7962 758
rect 8166 726 8198 758
rect 8378 726 8410 758
rect 8614 726 8646 758
rect 8826 726 8858 758
rect 102 479 134 511
rect 314 479 346 511
rect 550 479 582 511
rect 762 479 794 511
rect 998 479 1030 511
rect 1210 479 1242 511
rect 1446 479 1478 511
rect 1658 479 1690 511
rect 1894 479 1926 511
rect 2106 479 2138 511
rect 2342 479 2374 511
rect 2554 479 2586 511
rect 2790 479 2822 511
rect 3002 479 3034 511
rect 3238 479 3270 511
rect 3450 479 3482 511
rect 3686 479 3718 511
rect 3898 479 3930 511
rect 4134 479 4166 511
rect 4346 479 4378 511
rect 4582 479 4614 511
rect 4794 479 4826 511
rect 5030 479 5062 511
rect 5242 479 5274 511
rect 5478 479 5510 511
rect 5690 479 5722 511
rect 5926 479 5958 511
rect 6138 479 6170 511
rect 6374 479 6406 511
rect 6586 479 6618 511
rect 6822 479 6854 511
rect 7034 479 7066 511
rect 7270 479 7302 511
rect 7482 479 7514 511
rect 7718 479 7750 511
rect 7930 479 7962 511
rect 8166 479 8198 511
rect 8378 479 8410 511
rect 8614 479 8646 511
rect 8826 479 8858 511
rect 102 355 134 387
rect 314 355 346 387
rect 550 355 582 387
rect 762 355 794 387
rect 998 355 1030 387
rect 1210 355 1242 387
rect 1446 355 1478 387
rect 1658 355 1690 387
rect 1894 355 1926 387
rect 2106 355 2138 387
rect 2342 355 2374 387
rect 2554 355 2586 387
rect 2790 355 2822 387
rect 3002 355 3034 387
rect 3238 355 3270 387
rect 3450 355 3482 387
rect 3686 355 3718 387
rect 3898 355 3930 387
rect 4134 355 4166 387
rect 4346 355 4378 387
rect 4582 355 4614 387
rect 4794 355 4826 387
rect 5030 355 5062 387
rect 5242 355 5274 387
rect 5478 355 5510 387
rect 5690 355 5722 387
rect 5926 355 5958 387
rect 6138 355 6170 387
rect 6374 355 6406 387
rect 6586 355 6618 387
rect 6822 355 6854 387
rect 7034 355 7066 387
rect 7270 355 7302 387
rect 7482 355 7514 387
rect 7718 355 7750 387
rect 7930 355 7962 387
rect 8166 355 8198 387
rect 8378 355 8410 387
rect 8614 355 8646 387
rect 8826 355 8858 387
rect 102 231 134 263
rect 314 231 346 263
rect 550 231 582 263
rect 762 231 794 263
rect 998 231 1030 263
rect 1210 231 1242 263
rect 1446 231 1478 263
rect 1658 231 1690 263
rect 1894 231 1926 263
rect 2106 231 2138 263
rect 2342 231 2374 263
rect 2554 231 2586 263
rect 2790 231 2822 263
rect 3002 231 3034 263
rect 3238 231 3270 263
rect 3450 231 3482 263
rect 3686 231 3718 263
rect 3898 231 3930 263
rect 4134 231 4166 263
rect 4346 231 4378 263
rect 4582 231 4614 263
rect 4794 231 4826 263
rect 5030 231 5062 263
rect 5242 231 5274 263
rect 5478 231 5510 263
rect 5690 231 5722 263
rect 5926 231 5958 263
rect 6138 231 6170 263
rect 6374 231 6406 263
rect 6586 231 6618 263
rect 6822 231 6854 263
rect 7034 231 7066 263
rect 7270 231 7302 263
rect 7482 231 7514 263
rect 7718 231 7750 263
rect 7930 231 7962 263
rect 8166 231 8198 263
rect 8378 231 8410 263
rect 8614 231 8646 263
rect 8826 231 8858 263
rect 102 107 134 139
rect 314 107 346 139
rect 550 107 582 139
rect 762 107 794 139
rect 998 107 1030 139
rect 1210 107 1242 139
rect 1446 107 1478 139
rect 1658 107 1690 139
rect 1894 107 1926 139
rect 2106 107 2138 139
rect 2342 107 2374 139
rect 2554 107 2586 139
rect 2790 107 2822 139
rect 3002 107 3034 139
rect 3238 107 3270 139
rect 3450 107 3482 139
rect 3686 107 3718 139
rect 3898 107 3930 139
rect 4134 107 4166 139
rect 4346 107 4378 139
rect 4582 107 4614 139
rect 4794 107 4826 139
rect 5030 107 5062 139
rect 5242 107 5274 139
rect 5478 107 5510 139
rect 5690 107 5722 139
rect 5926 107 5958 139
rect 6138 107 6170 139
rect 6374 107 6406 139
rect 6586 107 6618 139
rect 6822 107 6854 139
rect 7034 107 7066 139
rect 7270 107 7302 139
rect 7482 107 7514 139
rect 7718 107 7750 139
rect 7930 107 7962 139
rect 8166 107 8198 139
rect 8378 107 8410 139
rect 8614 107 8646 139
rect 8826 107 8858 139
<< metal4 >>
rect 0 2460 8960 2492
rect 101 2369 134 2460
rect 314 2369 347 2460
rect 549 2369 582 2460
rect 762 2369 795 2460
rect 997 2369 1030 2460
rect 1210 2369 1243 2460
rect 1445 2369 1478 2460
rect 1658 2369 1691 2460
rect 1893 2369 1926 2460
rect 2106 2369 2139 2460
rect 2341 2369 2374 2460
rect 2554 2369 2587 2460
rect 2789 2369 2822 2460
rect 3002 2369 3035 2460
rect 3237 2369 3270 2460
rect 3450 2369 3483 2460
rect 3685 2369 3718 2460
rect 3898 2369 3931 2460
rect 4133 2369 4166 2460
rect 4346 2369 4379 2460
rect 4581 2369 4614 2460
rect 4794 2369 4827 2460
rect 5029 2369 5062 2460
rect 5242 2369 5275 2460
rect 5477 2369 5510 2460
rect 5690 2369 5723 2460
rect 5925 2369 5958 2460
rect 6138 2369 6171 2460
rect 6373 2369 6406 2460
rect 6586 2369 6619 2460
rect 6821 2369 6854 2460
rect 7034 2369 7067 2460
rect 7269 2369 7302 2460
rect 7482 2369 7515 2460
rect 7717 2369 7750 2460
rect 7930 2369 7963 2460
rect 8165 2369 8198 2460
rect 8378 2369 8411 2460
rect 8613 2369 8646 2460
rect 8826 2369 8859 2460
rect 99 2368 137 2369
rect 99 2367 102 2368
rect 54 2337 102 2367
rect 99 2336 102 2337
rect 134 2367 137 2368
rect 311 2368 349 2369
rect 311 2367 314 2368
rect 134 2337 181 2367
rect 267 2337 314 2367
rect 134 2336 137 2337
rect 99 2335 137 2336
rect 311 2336 314 2337
rect 346 2367 349 2368
rect 547 2368 585 2369
rect 547 2367 550 2368
rect 346 2337 394 2367
rect 502 2337 550 2367
rect 346 2336 349 2337
rect 311 2335 349 2336
rect 547 2336 550 2337
rect 582 2367 585 2368
rect 759 2368 797 2369
rect 759 2367 762 2368
rect 582 2337 629 2367
rect 715 2337 762 2367
rect 582 2336 585 2337
rect 547 2335 585 2336
rect 759 2336 762 2337
rect 794 2367 797 2368
rect 995 2368 1033 2369
rect 995 2367 998 2368
rect 794 2337 842 2367
rect 950 2337 998 2367
rect 794 2336 797 2337
rect 759 2335 797 2336
rect 995 2336 998 2337
rect 1030 2367 1033 2368
rect 1207 2368 1245 2369
rect 1207 2367 1210 2368
rect 1030 2337 1077 2367
rect 1163 2337 1210 2367
rect 1030 2336 1033 2337
rect 995 2335 1033 2336
rect 1207 2336 1210 2337
rect 1242 2367 1245 2368
rect 1443 2368 1481 2369
rect 1443 2367 1446 2368
rect 1242 2337 1290 2367
rect 1398 2337 1446 2367
rect 1242 2336 1245 2337
rect 1207 2335 1245 2336
rect 1443 2336 1446 2337
rect 1478 2367 1481 2368
rect 1655 2368 1693 2369
rect 1655 2367 1658 2368
rect 1478 2337 1525 2367
rect 1611 2337 1658 2367
rect 1478 2336 1481 2337
rect 1443 2335 1481 2336
rect 1655 2336 1658 2337
rect 1690 2367 1693 2368
rect 1891 2368 1929 2369
rect 1891 2367 1894 2368
rect 1690 2337 1738 2367
rect 1846 2337 1894 2367
rect 1690 2336 1693 2337
rect 1655 2335 1693 2336
rect 1891 2336 1894 2337
rect 1926 2367 1929 2368
rect 2103 2368 2141 2369
rect 2103 2367 2106 2368
rect 1926 2337 1973 2367
rect 2059 2337 2106 2367
rect 1926 2336 1929 2337
rect 1891 2335 1929 2336
rect 2103 2336 2106 2337
rect 2138 2367 2141 2368
rect 2339 2368 2377 2369
rect 2339 2367 2342 2368
rect 2138 2337 2186 2367
rect 2294 2337 2342 2367
rect 2138 2336 2141 2337
rect 2103 2335 2141 2336
rect 2339 2336 2342 2337
rect 2374 2367 2377 2368
rect 2551 2368 2589 2369
rect 2551 2367 2554 2368
rect 2374 2337 2421 2367
rect 2507 2337 2554 2367
rect 2374 2336 2377 2337
rect 2339 2335 2377 2336
rect 2551 2336 2554 2337
rect 2586 2367 2589 2368
rect 2787 2368 2825 2369
rect 2787 2367 2790 2368
rect 2586 2337 2634 2367
rect 2742 2337 2790 2367
rect 2586 2336 2589 2337
rect 2551 2335 2589 2336
rect 2787 2336 2790 2337
rect 2822 2367 2825 2368
rect 2999 2368 3037 2369
rect 2999 2367 3002 2368
rect 2822 2337 2869 2367
rect 2955 2337 3002 2367
rect 2822 2336 2825 2337
rect 2787 2335 2825 2336
rect 2999 2336 3002 2337
rect 3034 2367 3037 2368
rect 3235 2368 3273 2369
rect 3235 2367 3238 2368
rect 3034 2337 3082 2367
rect 3190 2337 3238 2367
rect 3034 2336 3037 2337
rect 2999 2335 3037 2336
rect 3235 2336 3238 2337
rect 3270 2367 3273 2368
rect 3447 2368 3485 2369
rect 3447 2367 3450 2368
rect 3270 2337 3317 2367
rect 3403 2337 3450 2367
rect 3270 2336 3273 2337
rect 3235 2335 3273 2336
rect 3447 2336 3450 2337
rect 3482 2367 3485 2368
rect 3683 2368 3721 2369
rect 3683 2367 3686 2368
rect 3482 2337 3530 2367
rect 3638 2337 3686 2367
rect 3482 2336 3485 2337
rect 3447 2335 3485 2336
rect 3683 2336 3686 2337
rect 3718 2367 3721 2368
rect 3895 2368 3933 2369
rect 3895 2367 3898 2368
rect 3718 2337 3765 2367
rect 3851 2337 3898 2367
rect 3718 2336 3721 2337
rect 3683 2335 3721 2336
rect 3895 2336 3898 2337
rect 3930 2367 3933 2368
rect 4131 2368 4169 2369
rect 4131 2367 4134 2368
rect 3930 2337 3978 2367
rect 4086 2337 4134 2367
rect 3930 2336 3933 2337
rect 3895 2335 3933 2336
rect 4131 2336 4134 2337
rect 4166 2367 4169 2368
rect 4343 2368 4381 2369
rect 4343 2367 4346 2368
rect 4166 2337 4213 2367
rect 4299 2337 4346 2367
rect 4166 2336 4169 2337
rect 4131 2335 4169 2336
rect 4343 2336 4346 2337
rect 4378 2367 4381 2368
rect 4579 2368 4617 2369
rect 4579 2367 4582 2368
rect 4378 2337 4426 2367
rect 4534 2337 4582 2367
rect 4378 2336 4381 2337
rect 4343 2335 4381 2336
rect 4579 2336 4582 2337
rect 4614 2367 4617 2368
rect 4791 2368 4829 2369
rect 4791 2367 4794 2368
rect 4614 2337 4661 2367
rect 4747 2337 4794 2367
rect 4614 2336 4617 2337
rect 4579 2335 4617 2336
rect 4791 2336 4794 2337
rect 4826 2367 4829 2368
rect 5027 2368 5065 2369
rect 5027 2367 5030 2368
rect 4826 2337 4874 2367
rect 4982 2337 5030 2367
rect 4826 2336 4829 2337
rect 4791 2335 4829 2336
rect 5027 2336 5030 2337
rect 5062 2367 5065 2368
rect 5239 2368 5277 2369
rect 5239 2367 5242 2368
rect 5062 2337 5109 2367
rect 5195 2337 5242 2367
rect 5062 2336 5065 2337
rect 5027 2335 5065 2336
rect 5239 2336 5242 2337
rect 5274 2367 5277 2368
rect 5475 2368 5513 2369
rect 5475 2367 5478 2368
rect 5274 2337 5322 2367
rect 5430 2337 5478 2367
rect 5274 2336 5277 2337
rect 5239 2335 5277 2336
rect 5475 2336 5478 2337
rect 5510 2367 5513 2368
rect 5687 2368 5725 2369
rect 5687 2367 5690 2368
rect 5510 2337 5557 2367
rect 5643 2337 5690 2367
rect 5510 2336 5513 2337
rect 5475 2335 5513 2336
rect 5687 2336 5690 2337
rect 5722 2367 5725 2368
rect 5923 2368 5961 2369
rect 5923 2367 5926 2368
rect 5722 2337 5770 2367
rect 5878 2337 5926 2367
rect 5722 2336 5725 2337
rect 5687 2335 5725 2336
rect 5923 2336 5926 2337
rect 5958 2367 5961 2368
rect 6135 2368 6173 2369
rect 6135 2367 6138 2368
rect 5958 2337 6005 2367
rect 6091 2337 6138 2367
rect 5958 2336 5961 2337
rect 5923 2335 5961 2336
rect 6135 2336 6138 2337
rect 6170 2367 6173 2368
rect 6371 2368 6409 2369
rect 6371 2367 6374 2368
rect 6170 2337 6218 2367
rect 6326 2337 6374 2367
rect 6170 2336 6173 2337
rect 6135 2335 6173 2336
rect 6371 2336 6374 2337
rect 6406 2367 6409 2368
rect 6583 2368 6621 2369
rect 6583 2367 6586 2368
rect 6406 2337 6453 2367
rect 6539 2337 6586 2367
rect 6406 2336 6409 2337
rect 6371 2335 6409 2336
rect 6583 2336 6586 2337
rect 6618 2367 6621 2368
rect 6819 2368 6857 2369
rect 6819 2367 6822 2368
rect 6618 2337 6666 2367
rect 6774 2337 6822 2367
rect 6618 2336 6621 2337
rect 6583 2335 6621 2336
rect 6819 2336 6822 2337
rect 6854 2367 6857 2368
rect 7031 2368 7069 2369
rect 7031 2367 7034 2368
rect 6854 2337 6901 2367
rect 6987 2337 7034 2367
rect 6854 2336 6857 2337
rect 6819 2335 6857 2336
rect 7031 2336 7034 2337
rect 7066 2367 7069 2368
rect 7267 2368 7305 2369
rect 7267 2367 7270 2368
rect 7066 2337 7114 2367
rect 7222 2337 7270 2367
rect 7066 2336 7069 2337
rect 7031 2335 7069 2336
rect 7267 2336 7270 2337
rect 7302 2367 7305 2368
rect 7479 2368 7517 2369
rect 7479 2367 7482 2368
rect 7302 2337 7349 2367
rect 7435 2337 7482 2367
rect 7302 2336 7305 2337
rect 7267 2335 7305 2336
rect 7479 2336 7482 2337
rect 7514 2367 7517 2368
rect 7715 2368 7753 2369
rect 7715 2367 7718 2368
rect 7514 2337 7562 2367
rect 7670 2337 7718 2367
rect 7514 2336 7517 2337
rect 7479 2335 7517 2336
rect 7715 2336 7718 2337
rect 7750 2367 7753 2368
rect 7927 2368 7965 2369
rect 7927 2367 7930 2368
rect 7750 2337 7797 2367
rect 7883 2337 7930 2367
rect 7750 2336 7753 2337
rect 7715 2335 7753 2336
rect 7927 2336 7930 2337
rect 7962 2367 7965 2368
rect 8163 2368 8201 2369
rect 8163 2367 8166 2368
rect 7962 2337 8010 2367
rect 8118 2337 8166 2367
rect 7962 2336 7965 2337
rect 7927 2335 7965 2336
rect 8163 2336 8166 2337
rect 8198 2367 8201 2368
rect 8375 2368 8413 2369
rect 8375 2367 8378 2368
rect 8198 2337 8245 2367
rect 8331 2337 8378 2367
rect 8198 2336 8201 2337
rect 8163 2335 8201 2336
rect 8375 2336 8378 2337
rect 8410 2367 8413 2368
rect 8611 2368 8649 2369
rect 8611 2367 8614 2368
rect 8410 2337 8458 2367
rect 8566 2337 8614 2367
rect 8410 2336 8413 2337
rect 8375 2335 8413 2336
rect 8611 2336 8614 2337
rect 8646 2367 8649 2368
rect 8823 2368 8861 2369
rect 8823 2367 8826 2368
rect 8646 2337 8693 2367
rect 8779 2337 8826 2367
rect 8646 2336 8649 2337
rect 8611 2335 8649 2336
rect 8823 2336 8826 2337
rect 8858 2367 8861 2368
rect 8858 2337 8906 2367
rect 8858 2336 8861 2337
rect 8823 2335 8861 2336
rect 101 2245 134 2335
rect 314 2245 347 2335
rect 549 2245 582 2335
rect 762 2245 795 2335
rect 997 2245 1030 2335
rect 1210 2245 1243 2335
rect 1445 2245 1478 2335
rect 1658 2245 1691 2335
rect 1893 2245 1926 2335
rect 2106 2245 2139 2335
rect 2341 2245 2374 2335
rect 2554 2245 2587 2335
rect 2789 2245 2822 2335
rect 3002 2245 3035 2335
rect 3237 2245 3270 2335
rect 3450 2245 3483 2335
rect 3685 2245 3718 2335
rect 3898 2245 3931 2335
rect 4133 2245 4166 2335
rect 4346 2245 4379 2335
rect 4581 2245 4614 2335
rect 4794 2245 4827 2335
rect 5029 2245 5062 2335
rect 5242 2245 5275 2335
rect 5477 2245 5510 2335
rect 5690 2245 5723 2335
rect 5925 2245 5958 2335
rect 6138 2245 6171 2335
rect 6373 2245 6406 2335
rect 6586 2245 6619 2335
rect 6821 2245 6854 2335
rect 7034 2245 7067 2335
rect 7269 2245 7302 2335
rect 7482 2245 7515 2335
rect 7717 2245 7750 2335
rect 7930 2245 7963 2335
rect 8165 2245 8198 2335
rect 8378 2245 8411 2335
rect 8613 2245 8646 2335
rect 8826 2245 8859 2335
rect 99 2244 137 2245
rect 99 2243 102 2244
rect 54 2213 102 2243
rect 99 2212 102 2213
rect 134 2243 137 2244
rect 311 2244 349 2245
rect 311 2243 314 2244
rect 134 2213 181 2243
rect 267 2213 314 2243
rect 134 2212 137 2213
rect 99 2211 137 2212
rect 311 2212 314 2213
rect 346 2243 349 2244
rect 547 2244 585 2245
rect 547 2243 550 2244
rect 346 2213 394 2243
rect 502 2213 550 2243
rect 346 2212 349 2213
rect 311 2211 349 2212
rect 547 2212 550 2213
rect 582 2243 585 2244
rect 759 2244 797 2245
rect 759 2243 762 2244
rect 582 2213 629 2243
rect 715 2213 762 2243
rect 582 2212 585 2213
rect 547 2211 585 2212
rect 759 2212 762 2213
rect 794 2243 797 2244
rect 995 2244 1033 2245
rect 995 2243 998 2244
rect 794 2213 842 2243
rect 950 2213 998 2243
rect 794 2212 797 2213
rect 759 2211 797 2212
rect 995 2212 998 2213
rect 1030 2243 1033 2244
rect 1207 2244 1245 2245
rect 1207 2243 1210 2244
rect 1030 2213 1077 2243
rect 1163 2213 1210 2243
rect 1030 2212 1033 2213
rect 995 2211 1033 2212
rect 1207 2212 1210 2213
rect 1242 2243 1245 2244
rect 1443 2244 1481 2245
rect 1443 2243 1446 2244
rect 1242 2213 1290 2243
rect 1398 2213 1446 2243
rect 1242 2212 1245 2213
rect 1207 2211 1245 2212
rect 1443 2212 1446 2213
rect 1478 2243 1481 2244
rect 1655 2244 1693 2245
rect 1655 2243 1658 2244
rect 1478 2213 1525 2243
rect 1611 2213 1658 2243
rect 1478 2212 1481 2213
rect 1443 2211 1481 2212
rect 1655 2212 1658 2213
rect 1690 2243 1693 2244
rect 1891 2244 1929 2245
rect 1891 2243 1894 2244
rect 1690 2213 1738 2243
rect 1846 2213 1894 2243
rect 1690 2212 1693 2213
rect 1655 2211 1693 2212
rect 1891 2212 1894 2213
rect 1926 2243 1929 2244
rect 2103 2244 2141 2245
rect 2103 2243 2106 2244
rect 1926 2213 1973 2243
rect 2059 2213 2106 2243
rect 1926 2212 1929 2213
rect 1891 2211 1929 2212
rect 2103 2212 2106 2213
rect 2138 2243 2141 2244
rect 2339 2244 2377 2245
rect 2339 2243 2342 2244
rect 2138 2213 2186 2243
rect 2294 2213 2342 2243
rect 2138 2212 2141 2213
rect 2103 2211 2141 2212
rect 2339 2212 2342 2213
rect 2374 2243 2377 2244
rect 2551 2244 2589 2245
rect 2551 2243 2554 2244
rect 2374 2213 2421 2243
rect 2507 2213 2554 2243
rect 2374 2212 2377 2213
rect 2339 2211 2377 2212
rect 2551 2212 2554 2213
rect 2586 2243 2589 2244
rect 2787 2244 2825 2245
rect 2787 2243 2790 2244
rect 2586 2213 2634 2243
rect 2742 2213 2790 2243
rect 2586 2212 2589 2213
rect 2551 2211 2589 2212
rect 2787 2212 2790 2213
rect 2822 2243 2825 2244
rect 2999 2244 3037 2245
rect 2999 2243 3002 2244
rect 2822 2213 2869 2243
rect 2955 2213 3002 2243
rect 2822 2212 2825 2213
rect 2787 2211 2825 2212
rect 2999 2212 3002 2213
rect 3034 2243 3037 2244
rect 3235 2244 3273 2245
rect 3235 2243 3238 2244
rect 3034 2213 3082 2243
rect 3190 2213 3238 2243
rect 3034 2212 3037 2213
rect 2999 2211 3037 2212
rect 3235 2212 3238 2213
rect 3270 2243 3273 2244
rect 3447 2244 3485 2245
rect 3447 2243 3450 2244
rect 3270 2213 3317 2243
rect 3403 2213 3450 2243
rect 3270 2212 3273 2213
rect 3235 2211 3273 2212
rect 3447 2212 3450 2213
rect 3482 2243 3485 2244
rect 3683 2244 3721 2245
rect 3683 2243 3686 2244
rect 3482 2213 3530 2243
rect 3638 2213 3686 2243
rect 3482 2212 3485 2213
rect 3447 2211 3485 2212
rect 3683 2212 3686 2213
rect 3718 2243 3721 2244
rect 3895 2244 3933 2245
rect 3895 2243 3898 2244
rect 3718 2213 3765 2243
rect 3851 2213 3898 2243
rect 3718 2212 3721 2213
rect 3683 2211 3721 2212
rect 3895 2212 3898 2213
rect 3930 2243 3933 2244
rect 4131 2244 4169 2245
rect 4131 2243 4134 2244
rect 3930 2213 3978 2243
rect 4086 2213 4134 2243
rect 3930 2212 3933 2213
rect 3895 2211 3933 2212
rect 4131 2212 4134 2213
rect 4166 2243 4169 2244
rect 4343 2244 4381 2245
rect 4343 2243 4346 2244
rect 4166 2213 4213 2243
rect 4299 2213 4346 2243
rect 4166 2212 4169 2213
rect 4131 2211 4169 2212
rect 4343 2212 4346 2213
rect 4378 2243 4381 2244
rect 4579 2244 4617 2245
rect 4579 2243 4582 2244
rect 4378 2213 4426 2243
rect 4534 2213 4582 2243
rect 4378 2212 4381 2213
rect 4343 2211 4381 2212
rect 4579 2212 4582 2213
rect 4614 2243 4617 2244
rect 4791 2244 4829 2245
rect 4791 2243 4794 2244
rect 4614 2213 4661 2243
rect 4747 2213 4794 2243
rect 4614 2212 4617 2213
rect 4579 2211 4617 2212
rect 4791 2212 4794 2213
rect 4826 2243 4829 2244
rect 5027 2244 5065 2245
rect 5027 2243 5030 2244
rect 4826 2213 4874 2243
rect 4982 2213 5030 2243
rect 4826 2212 4829 2213
rect 4791 2211 4829 2212
rect 5027 2212 5030 2213
rect 5062 2243 5065 2244
rect 5239 2244 5277 2245
rect 5239 2243 5242 2244
rect 5062 2213 5109 2243
rect 5195 2213 5242 2243
rect 5062 2212 5065 2213
rect 5027 2211 5065 2212
rect 5239 2212 5242 2213
rect 5274 2243 5277 2244
rect 5475 2244 5513 2245
rect 5475 2243 5478 2244
rect 5274 2213 5322 2243
rect 5430 2213 5478 2243
rect 5274 2212 5277 2213
rect 5239 2211 5277 2212
rect 5475 2212 5478 2213
rect 5510 2243 5513 2244
rect 5687 2244 5725 2245
rect 5687 2243 5690 2244
rect 5510 2213 5557 2243
rect 5643 2213 5690 2243
rect 5510 2212 5513 2213
rect 5475 2211 5513 2212
rect 5687 2212 5690 2213
rect 5722 2243 5725 2244
rect 5923 2244 5961 2245
rect 5923 2243 5926 2244
rect 5722 2213 5770 2243
rect 5878 2213 5926 2243
rect 5722 2212 5725 2213
rect 5687 2211 5725 2212
rect 5923 2212 5926 2213
rect 5958 2243 5961 2244
rect 6135 2244 6173 2245
rect 6135 2243 6138 2244
rect 5958 2213 6005 2243
rect 6091 2213 6138 2243
rect 5958 2212 5961 2213
rect 5923 2211 5961 2212
rect 6135 2212 6138 2213
rect 6170 2243 6173 2244
rect 6371 2244 6409 2245
rect 6371 2243 6374 2244
rect 6170 2213 6218 2243
rect 6326 2213 6374 2243
rect 6170 2212 6173 2213
rect 6135 2211 6173 2212
rect 6371 2212 6374 2213
rect 6406 2243 6409 2244
rect 6583 2244 6621 2245
rect 6583 2243 6586 2244
rect 6406 2213 6453 2243
rect 6539 2213 6586 2243
rect 6406 2212 6409 2213
rect 6371 2211 6409 2212
rect 6583 2212 6586 2213
rect 6618 2243 6621 2244
rect 6819 2244 6857 2245
rect 6819 2243 6822 2244
rect 6618 2213 6666 2243
rect 6774 2213 6822 2243
rect 6618 2212 6621 2213
rect 6583 2211 6621 2212
rect 6819 2212 6822 2213
rect 6854 2243 6857 2244
rect 7031 2244 7069 2245
rect 7031 2243 7034 2244
rect 6854 2213 6901 2243
rect 6987 2213 7034 2243
rect 6854 2212 6857 2213
rect 6819 2211 6857 2212
rect 7031 2212 7034 2213
rect 7066 2243 7069 2244
rect 7267 2244 7305 2245
rect 7267 2243 7270 2244
rect 7066 2213 7114 2243
rect 7222 2213 7270 2243
rect 7066 2212 7069 2213
rect 7031 2211 7069 2212
rect 7267 2212 7270 2213
rect 7302 2243 7305 2244
rect 7479 2244 7517 2245
rect 7479 2243 7482 2244
rect 7302 2213 7349 2243
rect 7435 2213 7482 2243
rect 7302 2212 7305 2213
rect 7267 2211 7305 2212
rect 7479 2212 7482 2213
rect 7514 2243 7517 2244
rect 7715 2244 7753 2245
rect 7715 2243 7718 2244
rect 7514 2213 7562 2243
rect 7670 2213 7718 2243
rect 7514 2212 7517 2213
rect 7479 2211 7517 2212
rect 7715 2212 7718 2213
rect 7750 2243 7753 2244
rect 7927 2244 7965 2245
rect 7927 2243 7930 2244
rect 7750 2213 7797 2243
rect 7883 2213 7930 2243
rect 7750 2212 7753 2213
rect 7715 2211 7753 2212
rect 7927 2212 7930 2213
rect 7962 2243 7965 2244
rect 8163 2244 8201 2245
rect 8163 2243 8166 2244
rect 7962 2213 8010 2243
rect 8118 2213 8166 2243
rect 7962 2212 7965 2213
rect 7927 2211 7965 2212
rect 8163 2212 8166 2213
rect 8198 2243 8201 2244
rect 8375 2244 8413 2245
rect 8375 2243 8378 2244
rect 8198 2213 8245 2243
rect 8331 2213 8378 2243
rect 8198 2212 8201 2213
rect 8163 2211 8201 2212
rect 8375 2212 8378 2213
rect 8410 2243 8413 2244
rect 8611 2244 8649 2245
rect 8611 2243 8614 2244
rect 8410 2213 8458 2243
rect 8566 2213 8614 2243
rect 8410 2212 8413 2213
rect 8375 2211 8413 2212
rect 8611 2212 8614 2213
rect 8646 2243 8649 2244
rect 8823 2244 8861 2245
rect 8823 2243 8826 2244
rect 8646 2213 8693 2243
rect 8779 2213 8826 2243
rect 8646 2212 8649 2213
rect 8611 2211 8649 2212
rect 8823 2212 8826 2213
rect 8858 2243 8861 2244
rect 8858 2213 8906 2243
rect 8858 2212 8861 2213
rect 8823 2211 8861 2212
rect 101 2121 134 2211
rect 314 2121 347 2211
rect 549 2121 582 2211
rect 762 2121 795 2211
rect 997 2121 1030 2211
rect 1210 2121 1243 2211
rect 1445 2121 1478 2211
rect 1658 2121 1691 2211
rect 1893 2121 1926 2211
rect 2106 2121 2139 2211
rect 2341 2121 2374 2211
rect 2554 2121 2587 2211
rect 2789 2121 2822 2211
rect 3002 2121 3035 2211
rect 3237 2121 3270 2211
rect 3450 2121 3483 2211
rect 3685 2121 3718 2211
rect 3898 2121 3931 2211
rect 4133 2121 4166 2211
rect 4346 2121 4379 2211
rect 4581 2121 4614 2211
rect 4794 2121 4827 2211
rect 5029 2121 5062 2211
rect 5242 2121 5275 2211
rect 5477 2121 5510 2211
rect 5690 2121 5723 2211
rect 5925 2121 5958 2211
rect 6138 2121 6171 2211
rect 6373 2121 6406 2211
rect 6586 2121 6619 2211
rect 6821 2121 6854 2211
rect 7034 2121 7067 2211
rect 7269 2121 7302 2211
rect 7482 2121 7515 2211
rect 7717 2121 7750 2211
rect 7930 2121 7963 2211
rect 8165 2121 8198 2211
rect 8378 2121 8411 2211
rect 8613 2121 8646 2211
rect 8826 2121 8859 2211
rect 99 2120 137 2121
rect 99 2119 102 2120
rect 54 2089 102 2119
rect 99 2088 102 2089
rect 134 2119 137 2120
rect 311 2120 349 2121
rect 311 2119 314 2120
rect 134 2089 181 2119
rect 267 2089 314 2119
rect 134 2088 137 2089
rect 99 2087 137 2088
rect 311 2088 314 2089
rect 346 2119 349 2120
rect 547 2120 585 2121
rect 547 2119 550 2120
rect 346 2089 394 2119
rect 502 2089 550 2119
rect 346 2088 349 2089
rect 311 2087 349 2088
rect 547 2088 550 2089
rect 582 2119 585 2120
rect 759 2120 797 2121
rect 759 2119 762 2120
rect 582 2089 629 2119
rect 715 2089 762 2119
rect 582 2088 585 2089
rect 547 2087 585 2088
rect 759 2088 762 2089
rect 794 2119 797 2120
rect 995 2120 1033 2121
rect 995 2119 998 2120
rect 794 2089 842 2119
rect 950 2089 998 2119
rect 794 2088 797 2089
rect 759 2087 797 2088
rect 995 2088 998 2089
rect 1030 2119 1033 2120
rect 1207 2120 1245 2121
rect 1207 2119 1210 2120
rect 1030 2089 1077 2119
rect 1163 2089 1210 2119
rect 1030 2088 1033 2089
rect 995 2087 1033 2088
rect 1207 2088 1210 2089
rect 1242 2119 1245 2120
rect 1443 2120 1481 2121
rect 1443 2119 1446 2120
rect 1242 2089 1290 2119
rect 1398 2089 1446 2119
rect 1242 2088 1245 2089
rect 1207 2087 1245 2088
rect 1443 2088 1446 2089
rect 1478 2119 1481 2120
rect 1655 2120 1693 2121
rect 1655 2119 1658 2120
rect 1478 2089 1525 2119
rect 1611 2089 1658 2119
rect 1478 2088 1481 2089
rect 1443 2087 1481 2088
rect 1655 2088 1658 2089
rect 1690 2119 1693 2120
rect 1891 2120 1929 2121
rect 1891 2119 1894 2120
rect 1690 2089 1738 2119
rect 1846 2089 1894 2119
rect 1690 2088 1693 2089
rect 1655 2087 1693 2088
rect 1891 2088 1894 2089
rect 1926 2119 1929 2120
rect 2103 2120 2141 2121
rect 2103 2119 2106 2120
rect 1926 2089 1973 2119
rect 2059 2089 2106 2119
rect 1926 2088 1929 2089
rect 1891 2087 1929 2088
rect 2103 2088 2106 2089
rect 2138 2119 2141 2120
rect 2339 2120 2377 2121
rect 2339 2119 2342 2120
rect 2138 2089 2186 2119
rect 2294 2089 2342 2119
rect 2138 2088 2141 2089
rect 2103 2087 2141 2088
rect 2339 2088 2342 2089
rect 2374 2119 2377 2120
rect 2551 2120 2589 2121
rect 2551 2119 2554 2120
rect 2374 2089 2421 2119
rect 2507 2089 2554 2119
rect 2374 2088 2377 2089
rect 2339 2087 2377 2088
rect 2551 2088 2554 2089
rect 2586 2119 2589 2120
rect 2787 2120 2825 2121
rect 2787 2119 2790 2120
rect 2586 2089 2634 2119
rect 2742 2089 2790 2119
rect 2586 2088 2589 2089
rect 2551 2087 2589 2088
rect 2787 2088 2790 2089
rect 2822 2119 2825 2120
rect 2999 2120 3037 2121
rect 2999 2119 3002 2120
rect 2822 2089 2869 2119
rect 2955 2089 3002 2119
rect 2822 2088 2825 2089
rect 2787 2087 2825 2088
rect 2999 2088 3002 2089
rect 3034 2119 3037 2120
rect 3235 2120 3273 2121
rect 3235 2119 3238 2120
rect 3034 2089 3082 2119
rect 3190 2089 3238 2119
rect 3034 2088 3037 2089
rect 2999 2087 3037 2088
rect 3235 2088 3238 2089
rect 3270 2119 3273 2120
rect 3447 2120 3485 2121
rect 3447 2119 3450 2120
rect 3270 2089 3317 2119
rect 3403 2089 3450 2119
rect 3270 2088 3273 2089
rect 3235 2087 3273 2088
rect 3447 2088 3450 2089
rect 3482 2119 3485 2120
rect 3683 2120 3721 2121
rect 3683 2119 3686 2120
rect 3482 2089 3530 2119
rect 3638 2089 3686 2119
rect 3482 2088 3485 2089
rect 3447 2087 3485 2088
rect 3683 2088 3686 2089
rect 3718 2119 3721 2120
rect 3895 2120 3933 2121
rect 3895 2119 3898 2120
rect 3718 2089 3765 2119
rect 3851 2089 3898 2119
rect 3718 2088 3721 2089
rect 3683 2087 3721 2088
rect 3895 2088 3898 2089
rect 3930 2119 3933 2120
rect 4131 2120 4169 2121
rect 4131 2119 4134 2120
rect 3930 2089 3978 2119
rect 4086 2089 4134 2119
rect 3930 2088 3933 2089
rect 3895 2087 3933 2088
rect 4131 2088 4134 2089
rect 4166 2119 4169 2120
rect 4343 2120 4381 2121
rect 4343 2119 4346 2120
rect 4166 2089 4213 2119
rect 4299 2089 4346 2119
rect 4166 2088 4169 2089
rect 4131 2087 4169 2088
rect 4343 2088 4346 2089
rect 4378 2119 4381 2120
rect 4579 2120 4617 2121
rect 4579 2119 4582 2120
rect 4378 2089 4426 2119
rect 4534 2089 4582 2119
rect 4378 2088 4381 2089
rect 4343 2087 4381 2088
rect 4579 2088 4582 2089
rect 4614 2119 4617 2120
rect 4791 2120 4829 2121
rect 4791 2119 4794 2120
rect 4614 2089 4661 2119
rect 4747 2089 4794 2119
rect 4614 2088 4617 2089
rect 4579 2087 4617 2088
rect 4791 2088 4794 2089
rect 4826 2119 4829 2120
rect 5027 2120 5065 2121
rect 5027 2119 5030 2120
rect 4826 2089 4874 2119
rect 4982 2089 5030 2119
rect 4826 2088 4829 2089
rect 4791 2087 4829 2088
rect 5027 2088 5030 2089
rect 5062 2119 5065 2120
rect 5239 2120 5277 2121
rect 5239 2119 5242 2120
rect 5062 2089 5109 2119
rect 5195 2089 5242 2119
rect 5062 2088 5065 2089
rect 5027 2087 5065 2088
rect 5239 2088 5242 2089
rect 5274 2119 5277 2120
rect 5475 2120 5513 2121
rect 5475 2119 5478 2120
rect 5274 2089 5322 2119
rect 5430 2089 5478 2119
rect 5274 2088 5277 2089
rect 5239 2087 5277 2088
rect 5475 2088 5478 2089
rect 5510 2119 5513 2120
rect 5687 2120 5725 2121
rect 5687 2119 5690 2120
rect 5510 2089 5557 2119
rect 5643 2089 5690 2119
rect 5510 2088 5513 2089
rect 5475 2087 5513 2088
rect 5687 2088 5690 2089
rect 5722 2119 5725 2120
rect 5923 2120 5961 2121
rect 5923 2119 5926 2120
rect 5722 2089 5770 2119
rect 5878 2089 5926 2119
rect 5722 2088 5725 2089
rect 5687 2087 5725 2088
rect 5923 2088 5926 2089
rect 5958 2119 5961 2120
rect 6135 2120 6173 2121
rect 6135 2119 6138 2120
rect 5958 2089 6005 2119
rect 6091 2089 6138 2119
rect 5958 2088 5961 2089
rect 5923 2087 5961 2088
rect 6135 2088 6138 2089
rect 6170 2119 6173 2120
rect 6371 2120 6409 2121
rect 6371 2119 6374 2120
rect 6170 2089 6218 2119
rect 6326 2089 6374 2119
rect 6170 2088 6173 2089
rect 6135 2087 6173 2088
rect 6371 2088 6374 2089
rect 6406 2119 6409 2120
rect 6583 2120 6621 2121
rect 6583 2119 6586 2120
rect 6406 2089 6453 2119
rect 6539 2089 6586 2119
rect 6406 2088 6409 2089
rect 6371 2087 6409 2088
rect 6583 2088 6586 2089
rect 6618 2119 6621 2120
rect 6819 2120 6857 2121
rect 6819 2119 6822 2120
rect 6618 2089 6666 2119
rect 6774 2089 6822 2119
rect 6618 2088 6621 2089
rect 6583 2087 6621 2088
rect 6819 2088 6822 2089
rect 6854 2119 6857 2120
rect 7031 2120 7069 2121
rect 7031 2119 7034 2120
rect 6854 2089 6901 2119
rect 6987 2089 7034 2119
rect 6854 2088 6857 2089
rect 6819 2087 6857 2088
rect 7031 2088 7034 2089
rect 7066 2119 7069 2120
rect 7267 2120 7305 2121
rect 7267 2119 7270 2120
rect 7066 2089 7114 2119
rect 7222 2089 7270 2119
rect 7066 2088 7069 2089
rect 7031 2087 7069 2088
rect 7267 2088 7270 2089
rect 7302 2119 7305 2120
rect 7479 2120 7517 2121
rect 7479 2119 7482 2120
rect 7302 2089 7349 2119
rect 7435 2089 7482 2119
rect 7302 2088 7305 2089
rect 7267 2087 7305 2088
rect 7479 2088 7482 2089
rect 7514 2119 7517 2120
rect 7715 2120 7753 2121
rect 7715 2119 7718 2120
rect 7514 2089 7562 2119
rect 7670 2089 7718 2119
rect 7514 2088 7517 2089
rect 7479 2087 7517 2088
rect 7715 2088 7718 2089
rect 7750 2119 7753 2120
rect 7927 2120 7965 2121
rect 7927 2119 7930 2120
rect 7750 2089 7797 2119
rect 7883 2089 7930 2119
rect 7750 2088 7753 2089
rect 7715 2087 7753 2088
rect 7927 2088 7930 2089
rect 7962 2119 7965 2120
rect 8163 2120 8201 2121
rect 8163 2119 8166 2120
rect 7962 2089 8010 2119
rect 8118 2089 8166 2119
rect 7962 2088 7965 2089
rect 7927 2087 7965 2088
rect 8163 2088 8166 2089
rect 8198 2119 8201 2120
rect 8375 2120 8413 2121
rect 8375 2119 8378 2120
rect 8198 2089 8245 2119
rect 8331 2089 8378 2119
rect 8198 2088 8201 2089
rect 8163 2087 8201 2088
rect 8375 2088 8378 2089
rect 8410 2119 8413 2120
rect 8611 2120 8649 2121
rect 8611 2119 8614 2120
rect 8410 2089 8458 2119
rect 8566 2089 8614 2119
rect 8410 2088 8413 2089
rect 8375 2087 8413 2088
rect 8611 2088 8614 2089
rect 8646 2119 8649 2120
rect 8823 2120 8861 2121
rect 8823 2119 8826 2120
rect 8646 2089 8693 2119
rect 8779 2089 8826 2119
rect 8646 2088 8649 2089
rect 8611 2087 8649 2088
rect 8823 2088 8826 2089
rect 8858 2119 8861 2120
rect 8858 2089 8906 2119
rect 8858 2088 8861 2089
rect 8823 2087 8861 2088
rect 101 1997 134 2087
rect 314 1997 347 2087
rect 549 1997 582 2087
rect 762 1997 795 2087
rect 997 1997 1030 2087
rect 1210 1997 1243 2087
rect 1445 1997 1478 2087
rect 1658 1997 1691 2087
rect 1893 1997 1926 2087
rect 2106 1997 2139 2087
rect 2341 1997 2374 2087
rect 2554 1997 2587 2087
rect 2789 1997 2822 2087
rect 3002 1997 3035 2087
rect 3237 1997 3270 2087
rect 3450 1997 3483 2087
rect 3685 1997 3718 2087
rect 3898 1997 3931 2087
rect 4133 1997 4166 2087
rect 4346 1997 4379 2087
rect 4581 1997 4614 2087
rect 4794 1997 4827 2087
rect 5029 1997 5062 2087
rect 5242 1997 5275 2087
rect 5477 1997 5510 2087
rect 5690 1997 5723 2087
rect 5925 1997 5958 2087
rect 6138 1997 6171 2087
rect 6373 1997 6406 2087
rect 6586 1997 6619 2087
rect 6821 1997 6854 2087
rect 7034 1997 7067 2087
rect 7269 1997 7302 2087
rect 7482 1997 7515 2087
rect 7717 1997 7750 2087
rect 7930 1997 7963 2087
rect 8165 1997 8198 2087
rect 8378 1997 8411 2087
rect 8613 1997 8646 2087
rect 8826 1997 8859 2087
rect 99 1996 137 1997
rect 99 1995 102 1996
rect 54 1965 102 1995
rect 99 1964 102 1965
rect 134 1995 137 1996
rect 311 1996 349 1997
rect 311 1995 314 1996
rect 134 1965 181 1995
rect 267 1965 314 1995
rect 134 1964 137 1965
rect 99 1963 137 1964
rect 311 1964 314 1965
rect 346 1995 349 1996
rect 547 1996 585 1997
rect 547 1995 550 1996
rect 346 1965 394 1995
rect 502 1965 550 1995
rect 346 1964 349 1965
rect 311 1963 349 1964
rect 547 1964 550 1965
rect 582 1995 585 1996
rect 759 1996 797 1997
rect 759 1995 762 1996
rect 582 1965 629 1995
rect 715 1965 762 1995
rect 582 1964 585 1965
rect 547 1963 585 1964
rect 759 1964 762 1965
rect 794 1995 797 1996
rect 995 1996 1033 1997
rect 995 1995 998 1996
rect 794 1965 842 1995
rect 950 1965 998 1995
rect 794 1964 797 1965
rect 759 1963 797 1964
rect 995 1964 998 1965
rect 1030 1995 1033 1996
rect 1207 1996 1245 1997
rect 1207 1995 1210 1996
rect 1030 1965 1077 1995
rect 1163 1965 1210 1995
rect 1030 1964 1033 1965
rect 995 1963 1033 1964
rect 1207 1964 1210 1965
rect 1242 1995 1245 1996
rect 1443 1996 1481 1997
rect 1443 1995 1446 1996
rect 1242 1965 1290 1995
rect 1398 1965 1446 1995
rect 1242 1964 1245 1965
rect 1207 1963 1245 1964
rect 1443 1964 1446 1965
rect 1478 1995 1481 1996
rect 1655 1996 1693 1997
rect 1655 1995 1658 1996
rect 1478 1965 1525 1995
rect 1611 1965 1658 1995
rect 1478 1964 1481 1965
rect 1443 1963 1481 1964
rect 1655 1964 1658 1965
rect 1690 1995 1693 1996
rect 1891 1996 1929 1997
rect 1891 1995 1894 1996
rect 1690 1965 1738 1995
rect 1846 1965 1894 1995
rect 1690 1964 1693 1965
rect 1655 1963 1693 1964
rect 1891 1964 1894 1965
rect 1926 1995 1929 1996
rect 2103 1996 2141 1997
rect 2103 1995 2106 1996
rect 1926 1965 1973 1995
rect 2059 1965 2106 1995
rect 1926 1964 1929 1965
rect 1891 1963 1929 1964
rect 2103 1964 2106 1965
rect 2138 1995 2141 1996
rect 2339 1996 2377 1997
rect 2339 1995 2342 1996
rect 2138 1965 2186 1995
rect 2294 1965 2342 1995
rect 2138 1964 2141 1965
rect 2103 1963 2141 1964
rect 2339 1964 2342 1965
rect 2374 1995 2377 1996
rect 2551 1996 2589 1997
rect 2551 1995 2554 1996
rect 2374 1965 2421 1995
rect 2507 1965 2554 1995
rect 2374 1964 2377 1965
rect 2339 1963 2377 1964
rect 2551 1964 2554 1965
rect 2586 1995 2589 1996
rect 2787 1996 2825 1997
rect 2787 1995 2790 1996
rect 2586 1965 2634 1995
rect 2742 1965 2790 1995
rect 2586 1964 2589 1965
rect 2551 1963 2589 1964
rect 2787 1964 2790 1965
rect 2822 1995 2825 1996
rect 2999 1996 3037 1997
rect 2999 1995 3002 1996
rect 2822 1965 2869 1995
rect 2955 1965 3002 1995
rect 2822 1964 2825 1965
rect 2787 1963 2825 1964
rect 2999 1964 3002 1965
rect 3034 1995 3037 1996
rect 3235 1996 3273 1997
rect 3235 1995 3238 1996
rect 3034 1965 3082 1995
rect 3190 1965 3238 1995
rect 3034 1964 3037 1965
rect 2999 1963 3037 1964
rect 3235 1964 3238 1965
rect 3270 1995 3273 1996
rect 3447 1996 3485 1997
rect 3447 1995 3450 1996
rect 3270 1965 3317 1995
rect 3403 1965 3450 1995
rect 3270 1964 3273 1965
rect 3235 1963 3273 1964
rect 3447 1964 3450 1965
rect 3482 1995 3485 1996
rect 3683 1996 3721 1997
rect 3683 1995 3686 1996
rect 3482 1965 3530 1995
rect 3638 1965 3686 1995
rect 3482 1964 3485 1965
rect 3447 1963 3485 1964
rect 3683 1964 3686 1965
rect 3718 1995 3721 1996
rect 3895 1996 3933 1997
rect 3895 1995 3898 1996
rect 3718 1965 3765 1995
rect 3851 1965 3898 1995
rect 3718 1964 3721 1965
rect 3683 1963 3721 1964
rect 3895 1964 3898 1965
rect 3930 1995 3933 1996
rect 4131 1996 4169 1997
rect 4131 1995 4134 1996
rect 3930 1965 3978 1995
rect 4086 1965 4134 1995
rect 3930 1964 3933 1965
rect 3895 1963 3933 1964
rect 4131 1964 4134 1965
rect 4166 1995 4169 1996
rect 4343 1996 4381 1997
rect 4343 1995 4346 1996
rect 4166 1965 4213 1995
rect 4299 1965 4346 1995
rect 4166 1964 4169 1965
rect 4131 1963 4169 1964
rect 4343 1964 4346 1965
rect 4378 1995 4381 1996
rect 4579 1996 4617 1997
rect 4579 1995 4582 1996
rect 4378 1965 4426 1995
rect 4534 1965 4582 1995
rect 4378 1964 4381 1965
rect 4343 1963 4381 1964
rect 4579 1964 4582 1965
rect 4614 1995 4617 1996
rect 4791 1996 4829 1997
rect 4791 1995 4794 1996
rect 4614 1965 4661 1995
rect 4747 1965 4794 1995
rect 4614 1964 4617 1965
rect 4579 1963 4617 1964
rect 4791 1964 4794 1965
rect 4826 1995 4829 1996
rect 5027 1996 5065 1997
rect 5027 1995 5030 1996
rect 4826 1965 4874 1995
rect 4982 1965 5030 1995
rect 4826 1964 4829 1965
rect 4791 1963 4829 1964
rect 5027 1964 5030 1965
rect 5062 1995 5065 1996
rect 5239 1996 5277 1997
rect 5239 1995 5242 1996
rect 5062 1965 5109 1995
rect 5195 1965 5242 1995
rect 5062 1964 5065 1965
rect 5027 1963 5065 1964
rect 5239 1964 5242 1965
rect 5274 1995 5277 1996
rect 5475 1996 5513 1997
rect 5475 1995 5478 1996
rect 5274 1965 5322 1995
rect 5430 1965 5478 1995
rect 5274 1964 5277 1965
rect 5239 1963 5277 1964
rect 5475 1964 5478 1965
rect 5510 1995 5513 1996
rect 5687 1996 5725 1997
rect 5687 1995 5690 1996
rect 5510 1965 5557 1995
rect 5643 1965 5690 1995
rect 5510 1964 5513 1965
rect 5475 1963 5513 1964
rect 5687 1964 5690 1965
rect 5722 1995 5725 1996
rect 5923 1996 5961 1997
rect 5923 1995 5926 1996
rect 5722 1965 5770 1995
rect 5878 1965 5926 1995
rect 5722 1964 5725 1965
rect 5687 1963 5725 1964
rect 5923 1964 5926 1965
rect 5958 1995 5961 1996
rect 6135 1996 6173 1997
rect 6135 1995 6138 1996
rect 5958 1965 6005 1995
rect 6091 1965 6138 1995
rect 5958 1964 5961 1965
rect 5923 1963 5961 1964
rect 6135 1964 6138 1965
rect 6170 1995 6173 1996
rect 6371 1996 6409 1997
rect 6371 1995 6374 1996
rect 6170 1965 6218 1995
rect 6326 1965 6374 1995
rect 6170 1964 6173 1965
rect 6135 1963 6173 1964
rect 6371 1964 6374 1965
rect 6406 1995 6409 1996
rect 6583 1996 6621 1997
rect 6583 1995 6586 1996
rect 6406 1965 6453 1995
rect 6539 1965 6586 1995
rect 6406 1964 6409 1965
rect 6371 1963 6409 1964
rect 6583 1964 6586 1965
rect 6618 1995 6621 1996
rect 6819 1996 6857 1997
rect 6819 1995 6822 1996
rect 6618 1965 6666 1995
rect 6774 1965 6822 1995
rect 6618 1964 6621 1965
rect 6583 1963 6621 1964
rect 6819 1964 6822 1965
rect 6854 1995 6857 1996
rect 7031 1996 7069 1997
rect 7031 1995 7034 1996
rect 6854 1965 6901 1995
rect 6987 1965 7034 1995
rect 6854 1964 6857 1965
rect 6819 1963 6857 1964
rect 7031 1964 7034 1965
rect 7066 1995 7069 1996
rect 7267 1996 7305 1997
rect 7267 1995 7270 1996
rect 7066 1965 7114 1995
rect 7222 1965 7270 1995
rect 7066 1964 7069 1965
rect 7031 1963 7069 1964
rect 7267 1964 7270 1965
rect 7302 1995 7305 1996
rect 7479 1996 7517 1997
rect 7479 1995 7482 1996
rect 7302 1965 7349 1995
rect 7435 1965 7482 1995
rect 7302 1964 7305 1965
rect 7267 1963 7305 1964
rect 7479 1964 7482 1965
rect 7514 1995 7517 1996
rect 7715 1996 7753 1997
rect 7715 1995 7718 1996
rect 7514 1965 7562 1995
rect 7670 1965 7718 1995
rect 7514 1964 7517 1965
rect 7479 1963 7517 1964
rect 7715 1964 7718 1965
rect 7750 1995 7753 1996
rect 7927 1996 7965 1997
rect 7927 1995 7930 1996
rect 7750 1965 7797 1995
rect 7883 1965 7930 1995
rect 7750 1964 7753 1965
rect 7715 1963 7753 1964
rect 7927 1964 7930 1965
rect 7962 1995 7965 1996
rect 8163 1996 8201 1997
rect 8163 1995 8166 1996
rect 7962 1965 8010 1995
rect 8118 1965 8166 1995
rect 7962 1964 7965 1965
rect 7927 1963 7965 1964
rect 8163 1964 8166 1965
rect 8198 1995 8201 1996
rect 8375 1996 8413 1997
rect 8375 1995 8378 1996
rect 8198 1965 8245 1995
rect 8331 1965 8378 1995
rect 8198 1964 8201 1965
rect 8163 1963 8201 1964
rect 8375 1964 8378 1965
rect 8410 1995 8413 1996
rect 8611 1996 8649 1997
rect 8611 1995 8614 1996
rect 8410 1965 8458 1995
rect 8566 1965 8614 1995
rect 8410 1964 8413 1965
rect 8375 1963 8413 1964
rect 8611 1964 8614 1965
rect 8646 1995 8649 1996
rect 8823 1996 8861 1997
rect 8823 1995 8826 1996
rect 8646 1965 8693 1995
rect 8779 1965 8826 1995
rect 8646 1964 8649 1965
rect 8611 1963 8649 1964
rect 8823 1964 8826 1965
rect 8858 1995 8861 1996
rect 8858 1965 8906 1995
rect 8858 1964 8861 1965
rect 8823 1963 8861 1964
rect 101 1873 134 1963
rect 314 1873 347 1963
rect 549 1917 582 1963
rect 762 1917 795 1963
rect 997 1917 1030 1963
rect 1210 1917 1243 1963
rect 1445 1917 1478 1963
rect 1658 1917 1691 1963
rect 1893 1873 1926 1963
rect 2106 1873 2139 1963
rect 2341 1873 2374 1963
rect 2554 1873 2587 1963
rect 2789 1917 2822 1963
rect 3002 1917 3035 1963
rect 3237 1917 3270 1963
rect 3450 1917 3483 1963
rect 3685 1917 3718 1963
rect 3898 1917 3931 1963
rect 4133 1873 4166 1963
rect 4346 1873 4379 1963
rect 4581 1873 4614 1963
rect 4794 1873 4827 1963
rect 5029 1917 5062 1963
rect 5242 1917 5275 1963
rect 5477 1917 5510 1963
rect 5690 1917 5723 1963
rect 5925 1917 5958 1963
rect 6138 1917 6171 1963
rect 6373 1873 6406 1963
rect 6586 1873 6619 1963
rect 6821 1873 6854 1963
rect 7034 1873 7067 1963
rect 7269 1917 7302 1963
rect 7482 1917 7515 1963
rect 7717 1917 7750 1963
rect 7930 1917 7963 1963
rect 8165 1917 8198 1963
rect 8378 1917 8411 1963
rect 8613 1873 8646 1963
rect 8826 1873 8859 1963
rect 0 1841 448 1873
rect 549 1841 1691 1873
rect 1792 1841 2688 1873
rect 2789 1841 3931 1873
rect 4032 1841 4928 1873
rect 5029 1841 6171 1873
rect 6272 1841 7168 1873
rect 7269 1841 8411 1873
rect 8512 1841 8960 1873
rect 101 1750 134 1841
rect 314 1750 347 1841
rect 549 1750 582 1841
rect 762 1750 795 1841
rect 997 1750 1030 1841
rect 1210 1750 1243 1841
rect 1445 1750 1478 1841
rect 1658 1750 1691 1841
rect 1893 1750 1926 1841
rect 2106 1750 2139 1841
rect 2341 1750 2374 1841
rect 2554 1750 2587 1841
rect 2789 1750 2822 1841
rect 3002 1750 3035 1841
rect 3237 1750 3270 1841
rect 3450 1750 3483 1841
rect 3685 1750 3718 1841
rect 3898 1750 3931 1841
rect 4133 1750 4166 1841
rect 4346 1750 4379 1841
rect 4581 1750 4614 1841
rect 4794 1750 4827 1841
rect 5029 1750 5062 1841
rect 5242 1750 5275 1841
rect 5477 1750 5510 1841
rect 5690 1750 5723 1841
rect 5925 1750 5958 1841
rect 6138 1750 6171 1841
rect 6373 1750 6406 1841
rect 6586 1750 6619 1841
rect 6821 1750 6854 1841
rect 7034 1750 7067 1841
rect 7269 1750 7302 1841
rect 7482 1750 7515 1841
rect 7717 1750 7750 1841
rect 7930 1750 7963 1841
rect 8165 1750 8198 1841
rect 8378 1750 8411 1841
rect 8613 1750 8646 1841
rect 8826 1750 8859 1841
rect 99 1749 137 1750
rect 99 1748 102 1749
rect 54 1718 102 1748
rect 99 1717 102 1718
rect 134 1748 137 1749
rect 311 1749 349 1750
rect 311 1748 314 1749
rect 134 1718 181 1748
rect 267 1718 314 1748
rect 134 1717 137 1718
rect 99 1716 137 1717
rect 311 1717 314 1718
rect 346 1748 349 1749
rect 547 1749 585 1750
rect 547 1748 550 1749
rect 346 1718 394 1748
rect 502 1718 550 1748
rect 346 1717 349 1718
rect 311 1716 349 1717
rect 547 1717 550 1718
rect 582 1748 585 1749
rect 759 1749 797 1750
rect 759 1748 762 1749
rect 582 1718 629 1748
rect 715 1718 762 1748
rect 582 1717 585 1718
rect 547 1716 585 1717
rect 759 1717 762 1718
rect 794 1748 797 1749
rect 995 1749 1033 1750
rect 995 1748 998 1749
rect 794 1718 842 1748
rect 950 1718 998 1748
rect 794 1717 797 1718
rect 759 1716 797 1717
rect 995 1717 998 1718
rect 1030 1748 1033 1749
rect 1207 1749 1245 1750
rect 1207 1748 1210 1749
rect 1030 1718 1077 1748
rect 1163 1718 1210 1748
rect 1030 1717 1033 1718
rect 995 1716 1033 1717
rect 1207 1717 1210 1718
rect 1242 1748 1245 1749
rect 1443 1749 1481 1750
rect 1443 1748 1446 1749
rect 1242 1718 1290 1748
rect 1398 1718 1446 1748
rect 1242 1717 1245 1718
rect 1207 1716 1245 1717
rect 1443 1717 1446 1718
rect 1478 1748 1481 1749
rect 1655 1749 1693 1750
rect 1655 1748 1658 1749
rect 1478 1718 1525 1748
rect 1611 1718 1658 1748
rect 1478 1717 1481 1718
rect 1443 1716 1481 1717
rect 1655 1717 1658 1718
rect 1690 1748 1693 1749
rect 1891 1749 1929 1750
rect 1891 1748 1894 1749
rect 1690 1718 1738 1748
rect 1846 1718 1894 1748
rect 1690 1717 1693 1718
rect 1655 1716 1693 1717
rect 1891 1717 1894 1718
rect 1926 1748 1929 1749
rect 2103 1749 2141 1750
rect 2103 1748 2106 1749
rect 1926 1718 1973 1748
rect 2059 1718 2106 1748
rect 1926 1717 1929 1718
rect 1891 1716 1929 1717
rect 2103 1717 2106 1718
rect 2138 1748 2141 1749
rect 2339 1749 2377 1750
rect 2339 1748 2342 1749
rect 2138 1718 2186 1748
rect 2294 1718 2342 1748
rect 2138 1717 2141 1718
rect 2103 1716 2141 1717
rect 2339 1717 2342 1718
rect 2374 1748 2377 1749
rect 2551 1749 2589 1750
rect 2551 1748 2554 1749
rect 2374 1718 2421 1748
rect 2507 1718 2554 1748
rect 2374 1717 2377 1718
rect 2339 1716 2377 1717
rect 2551 1717 2554 1718
rect 2586 1748 2589 1749
rect 2787 1749 2825 1750
rect 2787 1748 2790 1749
rect 2586 1718 2634 1748
rect 2742 1718 2790 1748
rect 2586 1717 2589 1718
rect 2551 1716 2589 1717
rect 2787 1717 2790 1718
rect 2822 1748 2825 1749
rect 2999 1749 3037 1750
rect 2999 1748 3002 1749
rect 2822 1718 2869 1748
rect 2955 1718 3002 1748
rect 2822 1717 2825 1718
rect 2787 1716 2825 1717
rect 2999 1717 3002 1718
rect 3034 1748 3037 1749
rect 3235 1749 3273 1750
rect 3235 1748 3238 1749
rect 3034 1718 3082 1748
rect 3190 1718 3238 1748
rect 3034 1717 3037 1718
rect 2999 1716 3037 1717
rect 3235 1717 3238 1718
rect 3270 1748 3273 1749
rect 3447 1749 3485 1750
rect 3447 1748 3450 1749
rect 3270 1718 3317 1748
rect 3403 1718 3450 1748
rect 3270 1717 3273 1718
rect 3235 1716 3273 1717
rect 3447 1717 3450 1718
rect 3482 1748 3485 1749
rect 3683 1749 3721 1750
rect 3683 1748 3686 1749
rect 3482 1718 3530 1748
rect 3638 1718 3686 1748
rect 3482 1717 3485 1718
rect 3447 1716 3485 1717
rect 3683 1717 3686 1718
rect 3718 1748 3721 1749
rect 3895 1749 3933 1750
rect 3895 1748 3898 1749
rect 3718 1718 3765 1748
rect 3851 1718 3898 1748
rect 3718 1717 3721 1718
rect 3683 1716 3721 1717
rect 3895 1717 3898 1718
rect 3930 1748 3933 1749
rect 4131 1749 4169 1750
rect 4131 1748 4134 1749
rect 3930 1718 3978 1748
rect 4086 1718 4134 1748
rect 3930 1717 3933 1718
rect 3895 1716 3933 1717
rect 4131 1717 4134 1718
rect 4166 1748 4169 1749
rect 4343 1749 4381 1750
rect 4343 1748 4346 1749
rect 4166 1718 4213 1748
rect 4299 1718 4346 1748
rect 4166 1717 4169 1718
rect 4131 1716 4169 1717
rect 4343 1717 4346 1718
rect 4378 1748 4381 1749
rect 4579 1749 4617 1750
rect 4579 1748 4582 1749
rect 4378 1718 4426 1748
rect 4534 1718 4582 1748
rect 4378 1717 4381 1718
rect 4343 1716 4381 1717
rect 4579 1717 4582 1718
rect 4614 1748 4617 1749
rect 4791 1749 4829 1750
rect 4791 1748 4794 1749
rect 4614 1718 4661 1748
rect 4747 1718 4794 1748
rect 4614 1717 4617 1718
rect 4579 1716 4617 1717
rect 4791 1717 4794 1718
rect 4826 1748 4829 1749
rect 5027 1749 5065 1750
rect 5027 1748 5030 1749
rect 4826 1718 4874 1748
rect 4982 1718 5030 1748
rect 4826 1717 4829 1718
rect 4791 1716 4829 1717
rect 5027 1717 5030 1718
rect 5062 1748 5065 1749
rect 5239 1749 5277 1750
rect 5239 1748 5242 1749
rect 5062 1718 5109 1748
rect 5195 1718 5242 1748
rect 5062 1717 5065 1718
rect 5027 1716 5065 1717
rect 5239 1717 5242 1718
rect 5274 1748 5277 1749
rect 5475 1749 5513 1750
rect 5475 1748 5478 1749
rect 5274 1718 5322 1748
rect 5430 1718 5478 1748
rect 5274 1717 5277 1718
rect 5239 1716 5277 1717
rect 5475 1717 5478 1718
rect 5510 1748 5513 1749
rect 5687 1749 5725 1750
rect 5687 1748 5690 1749
rect 5510 1718 5557 1748
rect 5643 1718 5690 1748
rect 5510 1717 5513 1718
rect 5475 1716 5513 1717
rect 5687 1717 5690 1718
rect 5722 1748 5725 1749
rect 5923 1749 5961 1750
rect 5923 1748 5926 1749
rect 5722 1718 5770 1748
rect 5878 1718 5926 1748
rect 5722 1717 5725 1718
rect 5687 1716 5725 1717
rect 5923 1717 5926 1718
rect 5958 1748 5961 1749
rect 6135 1749 6173 1750
rect 6135 1748 6138 1749
rect 5958 1718 6005 1748
rect 6091 1718 6138 1748
rect 5958 1717 5961 1718
rect 5923 1716 5961 1717
rect 6135 1717 6138 1718
rect 6170 1748 6173 1749
rect 6371 1749 6409 1750
rect 6371 1748 6374 1749
rect 6170 1718 6218 1748
rect 6326 1718 6374 1748
rect 6170 1717 6173 1718
rect 6135 1716 6173 1717
rect 6371 1717 6374 1718
rect 6406 1748 6409 1749
rect 6583 1749 6621 1750
rect 6583 1748 6586 1749
rect 6406 1718 6453 1748
rect 6539 1718 6586 1748
rect 6406 1717 6409 1718
rect 6371 1716 6409 1717
rect 6583 1717 6586 1718
rect 6618 1748 6621 1749
rect 6819 1749 6857 1750
rect 6819 1748 6822 1749
rect 6618 1718 6666 1748
rect 6774 1718 6822 1748
rect 6618 1717 6621 1718
rect 6583 1716 6621 1717
rect 6819 1717 6822 1718
rect 6854 1748 6857 1749
rect 7031 1749 7069 1750
rect 7031 1748 7034 1749
rect 6854 1718 6901 1748
rect 6987 1718 7034 1748
rect 6854 1717 6857 1718
rect 6819 1716 6857 1717
rect 7031 1717 7034 1718
rect 7066 1748 7069 1749
rect 7267 1749 7305 1750
rect 7267 1748 7270 1749
rect 7066 1718 7114 1748
rect 7222 1718 7270 1748
rect 7066 1717 7069 1718
rect 7031 1716 7069 1717
rect 7267 1717 7270 1718
rect 7302 1748 7305 1749
rect 7479 1749 7517 1750
rect 7479 1748 7482 1749
rect 7302 1718 7349 1748
rect 7435 1718 7482 1748
rect 7302 1717 7305 1718
rect 7267 1716 7305 1717
rect 7479 1717 7482 1718
rect 7514 1748 7517 1749
rect 7715 1749 7753 1750
rect 7715 1748 7718 1749
rect 7514 1718 7562 1748
rect 7670 1718 7718 1748
rect 7514 1717 7517 1718
rect 7479 1716 7517 1717
rect 7715 1717 7718 1718
rect 7750 1748 7753 1749
rect 7927 1749 7965 1750
rect 7927 1748 7930 1749
rect 7750 1718 7797 1748
rect 7883 1718 7930 1748
rect 7750 1717 7753 1718
rect 7715 1716 7753 1717
rect 7927 1717 7930 1718
rect 7962 1748 7965 1749
rect 8163 1749 8201 1750
rect 8163 1748 8166 1749
rect 7962 1718 8010 1748
rect 8118 1718 8166 1748
rect 7962 1717 7965 1718
rect 7927 1716 7965 1717
rect 8163 1717 8166 1718
rect 8198 1748 8201 1749
rect 8375 1749 8413 1750
rect 8375 1748 8378 1749
rect 8198 1718 8245 1748
rect 8331 1718 8378 1748
rect 8198 1717 8201 1718
rect 8163 1716 8201 1717
rect 8375 1717 8378 1718
rect 8410 1748 8413 1749
rect 8611 1749 8649 1750
rect 8611 1748 8614 1749
rect 8410 1718 8458 1748
rect 8566 1718 8614 1748
rect 8410 1717 8413 1718
rect 8375 1716 8413 1717
rect 8611 1717 8614 1718
rect 8646 1748 8649 1749
rect 8823 1749 8861 1750
rect 8823 1748 8826 1749
rect 8646 1718 8693 1748
rect 8779 1718 8826 1748
rect 8646 1717 8649 1718
rect 8611 1716 8649 1717
rect 8823 1717 8826 1718
rect 8858 1748 8861 1749
rect 8858 1718 8906 1748
rect 8858 1717 8861 1718
rect 8823 1716 8861 1717
rect 101 1626 134 1716
rect 314 1626 347 1716
rect 549 1626 582 1716
rect 762 1626 795 1716
rect 997 1626 1030 1716
rect 1210 1626 1243 1716
rect 1445 1626 1478 1716
rect 1658 1626 1691 1716
rect 1893 1626 1926 1716
rect 2106 1626 2139 1716
rect 2341 1626 2374 1716
rect 2554 1626 2587 1716
rect 2789 1626 2822 1716
rect 3002 1626 3035 1716
rect 3237 1626 3270 1716
rect 3450 1626 3483 1716
rect 3685 1626 3718 1716
rect 3898 1626 3931 1716
rect 4133 1626 4166 1716
rect 4346 1626 4379 1716
rect 4581 1626 4614 1716
rect 4794 1626 4827 1716
rect 5029 1626 5062 1716
rect 5242 1626 5275 1716
rect 5477 1626 5510 1716
rect 5690 1626 5723 1716
rect 5925 1626 5958 1716
rect 6138 1626 6171 1716
rect 6373 1626 6406 1716
rect 6586 1626 6619 1716
rect 6821 1626 6854 1716
rect 7034 1626 7067 1716
rect 7269 1626 7302 1716
rect 7482 1626 7515 1716
rect 7717 1626 7750 1716
rect 7930 1626 7963 1716
rect 8165 1626 8198 1716
rect 8378 1626 8411 1716
rect 8613 1626 8646 1716
rect 8826 1626 8859 1716
rect 99 1625 137 1626
rect 99 1624 102 1625
rect 54 1594 102 1624
rect 99 1593 102 1594
rect 134 1624 137 1625
rect 311 1625 349 1626
rect 311 1624 314 1625
rect 134 1594 181 1624
rect 267 1594 314 1624
rect 134 1593 137 1594
rect 99 1592 137 1593
rect 311 1593 314 1594
rect 346 1624 349 1625
rect 547 1625 585 1626
rect 547 1624 550 1625
rect 346 1594 394 1624
rect 502 1594 550 1624
rect 346 1593 349 1594
rect 311 1592 349 1593
rect 547 1593 550 1594
rect 582 1624 585 1625
rect 759 1625 797 1626
rect 759 1624 762 1625
rect 582 1594 629 1624
rect 715 1594 762 1624
rect 582 1593 585 1594
rect 547 1592 585 1593
rect 759 1593 762 1594
rect 794 1624 797 1625
rect 995 1625 1033 1626
rect 995 1624 998 1625
rect 794 1594 842 1624
rect 950 1594 998 1624
rect 794 1593 797 1594
rect 759 1592 797 1593
rect 995 1593 998 1594
rect 1030 1624 1033 1625
rect 1207 1625 1245 1626
rect 1207 1624 1210 1625
rect 1030 1594 1077 1624
rect 1163 1594 1210 1624
rect 1030 1593 1033 1594
rect 995 1592 1033 1593
rect 1207 1593 1210 1594
rect 1242 1624 1245 1625
rect 1443 1625 1481 1626
rect 1443 1624 1446 1625
rect 1242 1594 1290 1624
rect 1398 1594 1446 1624
rect 1242 1593 1245 1594
rect 1207 1592 1245 1593
rect 1443 1593 1446 1594
rect 1478 1624 1481 1625
rect 1655 1625 1693 1626
rect 1655 1624 1658 1625
rect 1478 1594 1525 1624
rect 1611 1594 1658 1624
rect 1478 1593 1481 1594
rect 1443 1592 1481 1593
rect 1655 1593 1658 1594
rect 1690 1624 1693 1625
rect 1891 1625 1929 1626
rect 1891 1624 1894 1625
rect 1690 1594 1738 1624
rect 1846 1594 1894 1624
rect 1690 1593 1693 1594
rect 1655 1592 1693 1593
rect 1891 1593 1894 1594
rect 1926 1624 1929 1625
rect 2103 1625 2141 1626
rect 2103 1624 2106 1625
rect 1926 1594 1973 1624
rect 2059 1594 2106 1624
rect 1926 1593 1929 1594
rect 1891 1592 1929 1593
rect 2103 1593 2106 1594
rect 2138 1624 2141 1625
rect 2339 1625 2377 1626
rect 2339 1624 2342 1625
rect 2138 1594 2186 1624
rect 2294 1594 2342 1624
rect 2138 1593 2141 1594
rect 2103 1592 2141 1593
rect 2339 1593 2342 1594
rect 2374 1624 2377 1625
rect 2551 1625 2589 1626
rect 2551 1624 2554 1625
rect 2374 1594 2421 1624
rect 2507 1594 2554 1624
rect 2374 1593 2377 1594
rect 2339 1592 2377 1593
rect 2551 1593 2554 1594
rect 2586 1624 2589 1625
rect 2787 1625 2825 1626
rect 2787 1624 2790 1625
rect 2586 1594 2634 1624
rect 2742 1594 2790 1624
rect 2586 1593 2589 1594
rect 2551 1592 2589 1593
rect 2787 1593 2790 1594
rect 2822 1624 2825 1625
rect 2999 1625 3037 1626
rect 2999 1624 3002 1625
rect 2822 1594 2869 1624
rect 2955 1594 3002 1624
rect 2822 1593 2825 1594
rect 2787 1592 2825 1593
rect 2999 1593 3002 1594
rect 3034 1624 3037 1625
rect 3235 1625 3273 1626
rect 3235 1624 3238 1625
rect 3034 1594 3082 1624
rect 3190 1594 3238 1624
rect 3034 1593 3037 1594
rect 2999 1592 3037 1593
rect 3235 1593 3238 1594
rect 3270 1624 3273 1625
rect 3447 1625 3485 1626
rect 3447 1624 3450 1625
rect 3270 1594 3317 1624
rect 3403 1594 3450 1624
rect 3270 1593 3273 1594
rect 3235 1592 3273 1593
rect 3447 1593 3450 1594
rect 3482 1624 3485 1625
rect 3683 1625 3721 1626
rect 3683 1624 3686 1625
rect 3482 1594 3530 1624
rect 3638 1594 3686 1624
rect 3482 1593 3485 1594
rect 3447 1592 3485 1593
rect 3683 1593 3686 1594
rect 3718 1624 3721 1625
rect 3895 1625 3933 1626
rect 3895 1624 3898 1625
rect 3718 1594 3765 1624
rect 3851 1594 3898 1624
rect 3718 1593 3721 1594
rect 3683 1592 3721 1593
rect 3895 1593 3898 1594
rect 3930 1624 3933 1625
rect 4131 1625 4169 1626
rect 4131 1624 4134 1625
rect 3930 1594 3978 1624
rect 4086 1594 4134 1624
rect 3930 1593 3933 1594
rect 3895 1592 3933 1593
rect 4131 1593 4134 1594
rect 4166 1624 4169 1625
rect 4343 1625 4381 1626
rect 4343 1624 4346 1625
rect 4166 1594 4213 1624
rect 4299 1594 4346 1624
rect 4166 1593 4169 1594
rect 4131 1592 4169 1593
rect 4343 1593 4346 1594
rect 4378 1624 4381 1625
rect 4579 1625 4617 1626
rect 4579 1624 4582 1625
rect 4378 1594 4426 1624
rect 4534 1594 4582 1624
rect 4378 1593 4381 1594
rect 4343 1592 4381 1593
rect 4579 1593 4582 1594
rect 4614 1624 4617 1625
rect 4791 1625 4829 1626
rect 4791 1624 4794 1625
rect 4614 1594 4661 1624
rect 4747 1594 4794 1624
rect 4614 1593 4617 1594
rect 4579 1592 4617 1593
rect 4791 1593 4794 1594
rect 4826 1624 4829 1625
rect 5027 1625 5065 1626
rect 5027 1624 5030 1625
rect 4826 1594 4874 1624
rect 4982 1594 5030 1624
rect 4826 1593 4829 1594
rect 4791 1592 4829 1593
rect 5027 1593 5030 1594
rect 5062 1624 5065 1625
rect 5239 1625 5277 1626
rect 5239 1624 5242 1625
rect 5062 1594 5109 1624
rect 5195 1594 5242 1624
rect 5062 1593 5065 1594
rect 5027 1592 5065 1593
rect 5239 1593 5242 1594
rect 5274 1624 5277 1625
rect 5475 1625 5513 1626
rect 5475 1624 5478 1625
rect 5274 1594 5322 1624
rect 5430 1594 5478 1624
rect 5274 1593 5277 1594
rect 5239 1592 5277 1593
rect 5475 1593 5478 1594
rect 5510 1624 5513 1625
rect 5687 1625 5725 1626
rect 5687 1624 5690 1625
rect 5510 1594 5557 1624
rect 5643 1594 5690 1624
rect 5510 1593 5513 1594
rect 5475 1592 5513 1593
rect 5687 1593 5690 1594
rect 5722 1624 5725 1625
rect 5923 1625 5961 1626
rect 5923 1624 5926 1625
rect 5722 1594 5770 1624
rect 5878 1594 5926 1624
rect 5722 1593 5725 1594
rect 5687 1592 5725 1593
rect 5923 1593 5926 1594
rect 5958 1624 5961 1625
rect 6135 1625 6173 1626
rect 6135 1624 6138 1625
rect 5958 1594 6005 1624
rect 6091 1594 6138 1624
rect 5958 1593 5961 1594
rect 5923 1592 5961 1593
rect 6135 1593 6138 1594
rect 6170 1624 6173 1625
rect 6371 1625 6409 1626
rect 6371 1624 6374 1625
rect 6170 1594 6218 1624
rect 6326 1594 6374 1624
rect 6170 1593 6173 1594
rect 6135 1592 6173 1593
rect 6371 1593 6374 1594
rect 6406 1624 6409 1625
rect 6583 1625 6621 1626
rect 6583 1624 6586 1625
rect 6406 1594 6453 1624
rect 6539 1594 6586 1624
rect 6406 1593 6409 1594
rect 6371 1592 6409 1593
rect 6583 1593 6586 1594
rect 6618 1624 6621 1625
rect 6819 1625 6857 1626
rect 6819 1624 6822 1625
rect 6618 1594 6666 1624
rect 6774 1594 6822 1624
rect 6618 1593 6621 1594
rect 6583 1592 6621 1593
rect 6819 1593 6822 1594
rect 6854 1624 6857 1625
rect 7031 1625 7069 1626
rect 7031 1624 7034 1625
rect 6854 1594 6901 1624
rect 6987 1594 7034 1624
rect 6854 1593 6857 1594
rect 6819 1592 6857 1593
rect 7031 1593 7034 1594
rect 7066 1624 7069 1625
rect 7267 1625 7305 1626
rect 7267 1624 7270 1625
rect 7066 1594 7114 1624
rect 7222 1594 7270 1624
rect 7066 1593 7069 1594
rect 7031 1592 7069 1593
rect 7267 1593 7270 1594
rect 7302 1624 7305 1625
rect 7479 1625 7517 1626
rect 7479 1624 7482 1625
rect 7302 1594 7349 1624
rect 7435 1594 7482 1624
rect 7302 1593 7305 1594
rect 7267 1592 7305 1593
rect 7479 1593 7482 1594
rect 7514 1624 7517 1625
rect 7715 1625 7753 1626
rect 7715 1624 7718 1625
rect 7514 1594 7562 1624
rect 7670 1594 7718 1624
rect 7514 1593 7517 1594
rect 7479 1592 7517 1593
rect 7715 1593 7718 1594
rect 7750 1624 7753 1625
rect 7927 1625 7965 1626
rect 7927 1624 7930 1625
rect 7750 1594 7797 1624
rect 7883 1594 7930 1624
rect 7750 1593 7753 1594
rect 7715 1592 7753 1593
rect 7927 1593 7930 1594
rect 7962 1624 7965 1625
rect 8163 1625 8201 1626
rect 8163 1624 8166 1625
rect 7962 1594 8010 1624
rect 8118 1594 8166 1624
rect 7962 1593 7965 1594
rect 7927 1592 7965 1593
rect 8163 1593 8166 1594
rect 8198 1624 8201 1625
rect 8375 1625 8413 1626
rect 8375 1624 8378 1625
rect 8198 1594 8245 1624
rect 8331 1594 8378 1624
rect 8198 1593 8201 1594
rect 8163 1592 8201 1593
rect 8375 1593 8378 1594
rect 8410 1624 8413 1625
rect 8611 1625 8649 1626
rect 8611 1624 8614 1625
rect 8410 1594 8458 1624
rect 8566 1594 8614 1624
rect 8410 1593 8413 1594
rect 8375 1592 8413 1593
rect 8611 1593 8614 1594
rect 8646 1624 8649 1625
rect 8823 1625 8861 1626
rect 8823 1624 8826 1625
rect 8646 1594 8693 1624
rect 8779 1594 8826 1624
rect 8646 1593 8649 1594
rect 8611 1592 8649 1593
rect 8823 1593 8826 1594
rect 8858 1624 8861 1625
rect 8858 1594 8906 1624
rect 8858 1593 8861 1594
rect 8823 1592 8861 1593
rect 101 1502 134 1592
rect 314 1502 347 1592
rect 549 1502 582 1592
rect 762 1502 795 1592
rect 997 1502 1030 1592
rect 1210 1502 1243 1592
rect 1445 1502 1478 1592
rect 1658 1502 1691 1592
rect 1893 1502 1926 1592
rect 2106 1502 2139 1592
rect 2341 1502 2374 1592
rect 2554 1502 2587 1592
rect 2789 1502 2822 1592
rect 3002 1502 3035 1592
rect 3237 1502 3270 1592
rect 3450 1502 3483 1592
rect 3685 1502 3718 1592
rect 3898 1502 3931 1592
rect 4133 1502 4166 1592
rect 4346 1502 4379 1592
rect 4581 1502 4614 1592
rect 4794 1502 4827 1592
rect 5029 1502 5062 1592
rect 5242 1502 5275 1592
rect 5477 1502 5510 1592
rect 5690 1502 5723 1592
rect 5925 1502 5958 1592
rect 6138 1502 6171 1592
rect 6373 1502 6406 1592
rect 6586 1502 6619 1592
rect 6821 1502 6854 1592
rect 7034 1502 7067 1592
rect 7269 1502 7302 1592
rect 7482 1502 7515 1592
rect 7717 1502 7750 1592
rect 7930 1502 7963 1592
rect 8165 1502 8198 1592
rect 8378 1502 8411 1592
rect 8613 1502 8646 1592
rect 8826 1502 8859 1592
rect 99 1501 137 1502
rect 99 1500 102 1501
rect 54 1470 102 1500
rect 99 1469 102 1470
rect 134 1500 137 1501
rect 311 1501 349 1502
rect 311 1500 314 1501
rect 134 1470 181 1500
rect 267 1470 314 1500
rect 134 1469 137 1470
rect 99 1468 137 1469
rect 311 1469 314 1470
rect 346 1500 349 1501
rect 547 1501 585 1502
rect 547 1500 550 1501
rect 346 1470 394 1500
rect 502 1470 550 1500
rect 346 1469 349 1470
rect 311 1468 349 1469
rect 547 1469 550 1470
rect 582 1500 585 1501
rect 759 1501 797 1502
rect 759 1500 762 1501
rect 582 1470 629 1500
rect 715 1470 762 1500
rect 582 1469 585 1470
rect 547 1468 585 1469
rect 759 1469 762 1470
rect 794 1500 797 1501
rect 995 1501 1033 1502
rect 995 1500 998 1501
rect 794 1470 842 1500
rect 950 1470 998 1500
rect 794 1469 797 1470
rect 759 1468 797 1469
rect 995 1469 998 1470
rect 1030 1500 1033 1501
rect 1207 1501 1245 1502
rect 1207 1500 1210 1501
rect 1030 1470 1077 1500
rect 1163 1470 1210 1500
rect 1030 1469 1033 1470
rect 995 1468 1033 1469
rect 1207 1469 1210 1470
rect 1242 1500 1245 1501
rect 1443 1501 1481 1502
rect 1443 1500 1446 1501
rect 1242 1470 1290 1500
rect 1398 1470 1446 1500
rect 1242 1469 1245 1470
rect 1207 1468 1245 1469
rect 1443 1469 1446 1470
rect 1478 1500 1481 1501
rect 1655 1501 1693 1502
rect 1655 1500 1658 1501
rect 1478 1470 1525 1500
rect 1611 1470 1658 1500
rect 1478 1469 1481 1470
rect 1443 1468 1481 1469
rect 1655 1469 1658 1470
rect 1690 1500 1693 1501
rect 1891 1501 1929 1502
rect 1891 1500 1894 1501
rect 1690 1470 1738 1500
rect 1846 1470 1894 1500
rect 1690 1469 1693 1470
rect 1655 1468 1693 1469
rect 1891 1469 1894 1470
rect 1926 1500 1929 1501
rect 2103 1501 2141 1502
rect 2103 1500 2106 1501
rect 1926 1470 1973 1500
rect 2059 1470 2106 1500
rect 1926 1469 1929 1470
rect 1891 1468 1929 1469
rect 2103 1469 2106 1470
rect 2138 1500 2141 1501
rect 2339 1501 2377 1502
rect 2339 1500 2342 1501
rect 2138 1470 2186 1500
rect 2294 1470 2342 1500
rect 2138 1469 2141 1470
rect 2103 1468 2141 1469
rect 2339 1469 2342 1470
rect 2374 1500 2377 1501
rect 2551 1501 2589 1502
rect 2551 1500 2554 1501
rect 2374 1470 2421 1500
rect 2507 1470 2554 1500
rect 2374 1469 2377 1470
rect 2339 1468 2377 1469
rect 2551 1469 2554 1470
rect 2586 1500 2589 1501
rect 2787 1501 2825 1502
rect 2787 1500 2790 1501
rect 2586 1470 2634 1500
rect 2742 1470 2790 1500
rect 2586 1469 2589 1470
rect 2551 1468 2589 1469
rect 2787 1469 2790 1470
rect 2822 1500 2825 1501
rect 2999 1501 3037 1502
rect 2999 1500 3002 1501
rect 2822 1470 2869 1500
rect 2955 1470 3002 1500
rect 2822 1469 2825 1470
rect 2787 1468 2825 1469
rect 2999 1469 3002 1470
rect 3034 1500 3037 1501
rect 3235 1501 3273 1502
rect 3235 1500 3238 1501
rect 3034 1470 3082 1500
rect 3190 1470 3238 1500
rect 3034 1469 3037 1470
rect 2999 1468 3037 1469
rect 3235 1469 3238 1470
rect 3270 1500 3273 1501
rect 3447 1501 3485 1502
rect 3447 1500 3450 1501
rect 3270 1470 3317 1500
rect 3403 1470 3450 1500
rect 3270 1469 3273 1470
rect 3235 1468 3273 1469
rect 3447 1469 3450 1470
rect 3482 1500 3485 1501
rect 3683 1501 3721 1502
rect 3683 1500 3686 1501
rect 3482 1470 3530 1500
rect 3638 1470 3686 1500
rect 3482 1469 3485 1470
rect 3447 1468 3485 1469
rect 3683 1469 3686 1470
rect 3718 1500 3721 1501
rect 3895 1501 3933 1502
rect 3895 1500 3898 1501
rect 3718 1470 3765 1500
rect 3851 1470 3898 1500
rect 3718 1469 3721 1470
rect 3683 1468 3721 1469
rect 3895 1469 3898 1470
rect 3930 1500 3933 1501
rect 4131 1501 4169 1502
rect 4131 1500 4134 1501
rect 3930 1470 3978 1500
rect 4086 1470 4134 1500
rect 3930 1469 3933 1470
rect 3895 1468 3933 1469
rect 4131 1469 4134 1470
rect 4166 1500 4169 1501
rect 4343 1501 4381 1502
rect 4343 1500 4346 1501
rect 4166 1470 4213 1500
rect 4299 1470 4346 1500
rect 4166 1469 4169 1470
rect 4131 1468 4169 1469
rect 4343 1469 4346 1470
rect 4378 1500 4381 1501
rect 4579 1501 4617 1502
rect 4579 1500 4582 1501
rect 4378 1470 4426 1500
rect 4534 1470 4582 1500
rect 4378 1469 4381 1470
rect 4343 1468 4381 1469
rect 4579 1469 4582 1470
rect 4614 1500 4617 1501
rect 4791 1501 4829 1502
rect 4791 1500 4794 1501
rect 4614 1470 4661 1500
rect 4747 1470 4794 1500
rect 4614 1469 4617 1470
rect 4579 1468 4617 1469
rect 4791 1469 4794 1470
rect 4826 1500 4829 1501
rect 5027 1501 5065 1502
rect 5027 1500 5030 1501
rect 4826 1470 4874 1500
rect 4982 1470 5030 1500
rect 4826 1469 4829 1470
rect 4791 1468 4829 1469
rect 5027 1469 5030 1470
rect 5062 1500 5065 1501
rect 5239 1501 5277 1502
rect 5239 1500 5242 1501
rect 5062 1470 5109 1500
rect 5195 1470 5242 1500
rect 5062 1469 5065 1470
rect 5027 1468 5065 1469
rect 5239 1469 5242 1470
rect 5274 1500 5277 1501
rect 5475 1501 5513 1502
rect 5475 1500 5478 1501
rect 5274 1470 5322 1500
rect 5430 1470 5478 1500
rect 5274 1469 5277 1470
rect 5239 1468 5277 1469
rect 5475 1469 5478 1470
rect 5510 1500 5513 1501
rect 5687 1501 5725 1502
rect 5687 1500 5690 1501
rect 5510 1470 5557 1500
rect 5643 1470 5690 1500
rect 5510 1469 5513 1470
rect 5475 1468 5513 1469
rect 5687 1469 5690 1470
rect 5722 1500 5725 1501
rect 5923 1501 5961 1502
rect 5923 1500 5926 1501
rect 5722 1470 5770 1500
rect 5878 1470 5926 1500
rect 5722 1469 5725 1470
rect 5687 1468 5725 1469
rect 5923 1469 5926 1470
rect 5958 1500 5961 1501
rect 6135 1501 6173 1502
rect 6135 1500 6138 1501
rect 5958 1470 6005 1500
rect 6091 1470 6138 1500
rect 5958 1469 5961 1470
rect 5923 1468 5961 1469
rect 6135 1469 6138 1470
rect 6170 1500 6173 1501
rect 6371 1501 6409 1502
rect 6371 1500 6374 1501
rect 6170 1470 6218 1500
rect 6326 1470 6374 1500
rect 6170 1469 6173 1470
rect 6135 1468 6173 1469
rect 6371 1469 6374 1470
rect 6406 1500 6409 1501
rect 6583 1501 6621 1502
rect 6583 1500 6586 1501
rect 6406 1470 6453 1500
rect 6539 1470 6586 1500
rect 6406 1469 6409 1470
rect 6371 1468 6409 1469
rect 6583 1469 6586 1470
rect 6618 1500 6621 1501
rect 6819 1501 6857 1502
rect 6819 1500 6822 1501
rect 6618 1470 6666 1500
rect 6774 1470 6822 1500
rect 6618 1469 6621 1470
rect 6583 1468 6621 1469
rect 6819 1469 6822 1470
rect 6854 1500 6857 1501
rect 7031 1501 7069 1502
rect 7031 1500 7034 1501
rect 6854 1470 6901 1500
rect 6987 1470 7034 1500
rect 6854 1469 6857 1470
rect 6819 1468 6857 1469
rect 7031 1469 7034 1470
rect 7066 1500 7069 1501
rect 7267 1501 7305 1502
rect 7267 1500 7270 1501
rect 7066 1470 7114 1500
rect 7222 1470 7270 1500
rect 7066 1469 7069 1470
rect 7031 1468 7069 1469
rect 7267 1469 7270 1470
rect 7302 1500 7305 1501
rect 7479 1501 7517 1502
rect 7479 1500 7482 1501
rect 7302 1470 7349 1500
rect 7435 1470 7482 1500
rect 7302 1469 7305 1470
rect 7267 1468 7305 1469
rect 7479 1469 7482 1470
rect 7514 1500 7517 1501
rect 7715 1501 7753 1502
rect 7715 1500 7718 1501
rect 7514 1470 7562 1500
rect 7670 1470 7718 1500
rect 7514 1469 7517 1470
rect 7479 1468 7517 1469
rect 7715 1469 7718 1470
rect 7750 1500 7753 1501
rect 7927 1501 7965 1502
rect 7927 1500 7930 1501
rect 7750 1470 7797 1500
rect 7883 1470 7930 1500
rect 7750 1469 7753 1470
rect 7715 1468 7753 1469
rect 7927 1469 7930 1470
rect 7962 1500 7965 1501
rect 8163 1501 8201 1502
rect 8163 1500 8166 1501
rect 7962 1470 8010 1500
rect 8118 1470 8166 1500
rect 7962 1469 7965 1470
rect 7927 1468 7965 1469
rect 8163 1469 8166 1470
rect 8198 1500 8201 1501
rect 8375 1501 8413 1502
rect 8375 1500 8378 1501
rect 8198 1470 8245 1500
rect 8331 1470 8378 1500
rect 8198 1469 8201 1470
rect 8163 1468 8201 1469
rect 8375 1469 8378 1470
rect 8410 1500 8413 1501
rect 8611 1501 8649 1502
rect 8611 1500 8614 1501
rect 8410 1470 8458 1500
rect 8566 1470 8614 1500
rect 8410 1469 8413 1470
rect 8375 1468 8413 1469
rect 8611 1469 8614 1470
rect 8646 1500 8649 1501
rect 8823 1501 8861 1502
rect 8823 1500 8826 1501
rect 8646 1470 8693 1500
rect 8779 1470 8826 1500
rect 8646 1469 8649 1470
rect 8611 1468 8649 1469
rect 8823 1469 8826 1470
rect 8858 1500 8861 1501
rect 8858 1470 8906 1500
rect 8858 1469 8861 1470
rect 8823 1468 8861 1469
rect 101 1378 134 1468
rect 314 1378 347 1468
rect 549 1378 582 1468
rect 762 1378 795 1468
rect 997 1378 1030 1468
rect 1210 1378 1243 1468
rect 1445 1378 1478 1468
rect 1658 1378 1691 1468
rect 1893 1378 1926 1468
rect 2106 1378 2139 1468
rect 2341 1378 2374 1468
rect 2554 1378 2587 1468
rect 2789 1378 2822 1468
rect 3002 1378 3035 1468
rect 3237 1378 3270 1468
rect 3450 1378 3483 1468
rect 3685 1378 3718 1468
rect 3898 1378 3931 1468
rect 4133 1378 4166 1468
rect 4346 1378 4379 1468
rect 4581 1378 4614 1468
rect 4794 1378 4827 1468
rect 5029 1378 5062 1468
rect 5242 1378 5275 1468
rect 5477 1378 5510 1468
rect 5690 1378 5723 1468
rect 5925 1378 5958 1468
rect 6138 1378 6171 1468
rect 6373 1378 6406 1468
rect 6586 1378 6619 1468
rect 6821 1378 6854 1468
rect 7034 1378 7067 1468
rect 7269 1378 7302 1468
rect 7482 1378 7515 1468
rect 7717 1378 7750 1468
rect 7930 1378 7963 1468
rect 8165 1378 8198 1468
rect 8378 1378 8411 1468
rect 8613 1378 8646 1468
rect 8826 1378 8859 1468
rect 99 1377 137 1378
rect 99 1376 102 1377
rect 54 1346 102 1376
rect 99 1345 102 1346
rect 134 1376 137 1377
rect 311 1377 349 1378
rect 311 1376 314 1377
rect 134 1346 181 1376
rect 267 1346 314 1376
rect 134 1345 137 1346
rect 99 1344 137 1345
rect 311 1345 314 1346
rect 346 1376 349 1377
rect 547 1377 585 1378
rect 547 1376 550 1377
rect 346 1346 394 1376
rect 502 1346 550 1376
rect 346 1345 349 1346
rect 311 1344 349 1345
rect 547 1345 550 1346
rect 582 1376 585 1377
rect 759 1377 797 1378
rect 759 1376 762 1377
rect 582 1346 629 1376
rect 715 1346 762 1376
rect 582 1345 585 1346
rect 547 1344 585 1345
rect 759 1345 762 1346
rect 794 1376 797 1377
rect 995 1377 1033 1378
rect 995 1376 998 1377
rect 794 1346 842 1376
rect 950 1346 998 1376
rect 794 1345 797 1346
rect 759 1344 797 1345
rect 995 1345 998 1346
rect 1030 1376 1033 1377
rect 1207 1377 1245 1378
rect 1207 1376 1210 1377
rect 1030 1346 1077 1376
rect 1163 1346 1210 1376
rect 1030 1345 1033 1346
rect 995 1344 1033 1345
rect 1207 1345 1210 1346
rect 1242 1376 1245 1377
rect 1443 1377 1481 1378
rect 1443 1376 1446 1377
rect 1242 1346 1290 1376
rect 1398 1346 1446 1376
rect 1242 1345 1245 1346
rect 1207 1344 1245 1345
rect 1443 1345 1446 1346
rect 1478 1376 1481 1377
rect 1655 1377 1693 1378
rect 1655 1376 1658 1377
rect 1478 1346 1525 1376
rect 1611 1346 1658 1376
rect 1478 1345 1481 1346
rect 1443 1344 1481 1345
rect 1655 1345 1658 1346
rect 1690 1376 1693 1377
rect 1891 1377 1929 1378
rect 1891 1376 1894 1377
rect 1690 1346 1738 1376
rect 1846 1346 1894 1376
rect 1690 1345 1693 1346
rect 1655 1344 1693 1345
rect 1891 1345 1894 1346
rect 1926 1376 1929 1377
rect 2103 1377 2141 1378
rect 2103 1376 2106 1377
rect 1926 1346 1973 1376
rect 2059 1346 2106 1376
rect 1926 1345 1929 1346
rect 1891 1344 1929 1345
rect 2103 1345 2106 1346
rect 2138 1376 2141 1377
rect 2339 1377 2377 1378
rect 2339 1376 2342 1377
rect 2138 1346 2186 1376
rect 2294 1346 2342 1376
rect 2138 1345 2141 1346
rect 2103 1344 2141 1345
rect 2339 1345 2342 1346
rect 2374 1376 2377 1377
rect 2551 1377 2589 1378
rect 2551 1376 2554 1377
rect 2374 1346 2421 1376
rect 2507 1346 2554 1376
rect 2374 1345 2377 1346
rect 2339 1344 2377 1345
rect 2551 1345 2554 1346
rect 2586 1376 2589 1377
rect 2787 1377 2825 1378
rect 2787 1376 2790 1377
rect 2586 1346 2634 1376
rect 2742 1346 2790 1376
rect 2586 1345 2589 1346
rect 2551 1344 2589 1345
rect 2787 1345 2790 1346
rect 2822 1376 2825 1377
rect 2999 1377 3037 1378
rect 2999 1376 3002 1377
rect 2822 1346 2869 1376
rect 2955 1346 3002 1376
rect 2822 1345 2825 1346
rect 2787 1344 2825 1345
rect 2999 1345 3002 1346
rect 3034 1376 3037 1377
rect 3235 1377 3273 1378
rect 3235 1376 3238 1377
rect 3034 1346 3082 1376
rect 3190 1346 3238 1376
rect 3034 1345 3037 1346
rect 2999 1344 3037 1345
rect 3235 1345 3238 1346
rect 3270 1376 3273 1377
rect 3447 1377 3485 1378
rect 3447 1376 3450 1377
rect 3270 1346 3317 1376
rect 3403 1346 3450 1376
rect 3270 1345 3273 1346
rect 3235 1344 3273 1345
rect 3447 1345 3450 1346
rect 3482 1376 3485 1377
rect 3683 1377 3721 1378
rect 3683 1376 3686 1377
rect 3482 1346 3530 1376
rect 3638 1346 3686 1376
rect 3482 1345 3485 1346
rect 3447 1344 3485 1345
rect 3683 1345 3686 1346
rect 3718 1376 3721 1377
rect 3895 1377 3933 1378
rect 3895 1376 3898 1377
rect 3718 1346 3765 1376
rect 3851 1346 3898 1376
rect 3718 1345 3721 1346
rect 3683 1344 3721 1345
rect 3895 1345 3898 1346
rect 3930 1376 3933 1377
rect 4131 1377 4169 1378
rect 4131 1376 4134 1377
rect 3930 1346 3978 1376
rect 4086 1346 4134 1376
rect 3930 1345 3933 1346
rect 3895 1344 3933 1345
rect 4131 1345 4134 1346
rect 4166 1376 4169 1377
rect 4343 1377 4381 1378
rect 4343 1376 4346 1377
rect 4166 1346 4213 1376
rect 4299 1346 4346 1376
rect 4166 1345 4169 1346
rect 4131 1344 4169 1345
rect 4343 1345 4346 1346
rect 4378 1376 4381 1377
rect 4579 1377 4617 1378
rect 4579 1376 4582 1377
rect 4378 1346 4426 1376
rect 4534 1346 4582 1376
rect 4378 1345 4381 1346
rect 4343 1344 4381 1345
rect 4579 1345 4582 1346
rect 4614 1376 4617 1377
rect 4791 1377 4829 1378
rect 4791 1376 4794 1377
rect 4614 1346 4661 1376
rect 4747 1346 4794 1376
rect 4614 1345 4617 1346
rect 4579 1344 4617 1345
rect 4791 1345 4794 1346
rect 4826 1376 4829 1377
rect 5027 1377 5065 1378
rect 5027 1376 5030 1377
rect 4826 1346 4874 1376
rect 4982 1346 5030 1376
rect 4826 1345 4829 1346
rect 4791 1344 4829 1345
rect 5027 1345 5030 1346
rect 5062 1376 5065 1377
rect 5239 1377 5277 1378
rect 5239 1376 5242 1377
rect 5062 1346 5109 1376
rect 5195 1346 5242 1376
rect 5062 1345 5065 1346
rect 5027 1344 5065 1345
rect 5239 1345 5242 1346
rect 5274 1376 5277 1377
rect 5475 1377 5513 1378
rect 5475 1376 5478 1377
rect 5274 1346 5322 1376
rect 5430 1346 5478 1376
rect 5274 1345 5277 1346
rect 5239 1344 5277 1345
rect 5475 1345 5478 1346
rect 5510 1376 5513 1377
rect 5687 1377 5725 1378
rect 5687 1376 5690 1377
rect 5510 1346 5557 1376
rect 5643 1346 5690 1376
rect 5510 1345 5513 1346
rect 5475 1344 5513 1345
rect 5687 1345 5690 1346
rect 5722 1376 5725 1377
rect 5923 1377 5961 1378
rect 5923 1376 5926 1377
rect 5722 1346 5770 1376
rect 5878 1346 5926 1376
rect 5722 1345 5725 1346
rect 5687 1344 5725 1345
rect 5923 1345 5926 1346
rect 5958 1376 5961 1377
rect 6135 1377 6173 1378
rect 6135 1376 6138 1377
rect 5958 1346 6005 1376
rect 6091 1346 6138 1376
rect 5958 1345 5961 1346
rect 5923 1344 5961 1345
rect 6135 1345 6138 1346
rect 6170 1376 6173 1377
rect 6371 1377 6409 1378
rect 6371 1376 6374 1377
rect 6170 1346 6218 1376
rect 6326 1346 6374 1376
rect 6170 1345 6173 1346
rect 6135 1344 6173 1345
rect 6371 1345 6374 1346
rect 6406 1376 6409 1377
rect 6583 1377 6621 1378
rect 6583 1376 6586 1377
rect 6406 1346 6453 1376
rect 6539 1346 6586 1376
rect 6406 1345 6409 1346
rect 6371 1344 6409 1345
rect 6583 1345 6586 1346
rect 6618 1376 6621 1377
rect 6819 1377 6857 1378
rect 6819 1376 6822 1377
rect 6618 1346 6666 1376
rect 6774 1346 6822 1376
rect 6618 1345 6621 1346
rect 6583 1344 6621 1345
rect 6819 1345 6822 1346
rect 6854 1376 6857 1377
rect 7031 1377 7069 1378
rect 7031 1376 7034 1377
rect 6854 1346 6901 1376
rect 6987 1346 7034 1376
rect 6854 1345 6857 1346
rect 6819 1344 6857 1345
rect 7031 1345 7034 1346
rect 7066 1376 7069 1377
rect 7267 1377 7305 1378
rect 7267 1376 7270 1377
rect 7066 1346 7114 1376
rect 7222 1346 7270 1376
rect 7066 1345 7069 1346
rect 7031 1344 7069 1345
rect 7267 1345 7270 1346
rect 7302 1376 7305 1377
rect 7479 1377 7517 1378
rect 7479 1376 7482 1377
rect 7302 1346 7349 1376
rect 7435 1346 7482 1376
rect 7302 1345 7305 1346
rect 7267 1344 7305 1345
rect 7479 1345 7482 1346
rect 7514 1376 7517 1377
rect 7715 1377 7753 1378
rect 7715 1376 7718 1377
rect 7514 1346 7562 1376
rect 7670 1346 7718 1376
rect 7514 1345 7517 1346
rect 7479 1344 7517 1345
rect 7715 1345 7718 1346
rect 7750 1376 7753 1377
rect 7927 1377 7965 1378
rect 7927 1376 7930 1377
rect 7750 1346 7797 1376
rect 7883 1346 7930 1376
rect 7750 1345 7753 1346
rect 7715 1344 7753 1345
rect 7927 1345 7930 1346
rect 7962 1376 7965 1377
rect 8163 1377 8201 1378
rect 8163 1376 8166 1377
rect 7962 1346 8010 1376
rect 8118 1346 8166 1376
rect 7962 1345 7965 1346
rect 7927 1344 7965 1345
rect 8163 1345 8166 1346
rect 8198 1376 8201 1377
rect 8375 1377 8413 1378
rect 8375 1376 8378 1377
rect 8198 1346 8245 1376
rect 8331 1346 8378 1376
rect 8198 1345 8201 1346
rect 8163 1344 8201 1345
rect 8375 1345 8378 1346
rect 8410 1376 8413 1377
rect 8611 1377 8649 1378
rect 8611 1376 8614 1377
rect 8410 1346 8458 1376
rect 8566 1346 8614 1376
rect 8410 1345 8413 1346
rect 8375 1344 8413 1345
rect 8611 1345 8614 1346
rect 8646 1376 8649 1377
rect 8823 1377 8861 1378
rect 8823 1376 8826 1377
rect 8646 1346 8693 1376
rect 8779 1346 8826 1376
rect 8646 1345 8649 1346
rect 8611 1344 8649 1345
rect 8823 1345 8826 1346
rect 8858 1376 8861 1377
rect 8858 1346 8906 1376
rect 8858 1345 8861 1346
rect 8823 1344 8861 1345
rect 101 1254 134 1344
rect 314 1254 347 1344
rect 549 1254 582 1344
rect 762 1254 795 1344
rect 997 1254 1030 1344
rect 1210 1254 1243 1344
rect 1445 1254 1478 1344
rect 1658 1254 1691 1344
rect 1893 1254 1926 1344
rect 2106 1254 2139 1344
rect 2341 1254 2374 1344
rect 2554 1254 2587 1344
rect 2789 1254 2822 1344
rect 3002 1254 3035 1344
rect 3237 1254 3270 1344
rect 3450 1254 3483 1344
rect 3685 1254 3718 1344
rect 3898 1254 3931 1344
rect 4133 1254 4166 1344
rect 4346 1254 4379 1344
rect 4581 1254 4614 1344
rect 4794 1254 4827 1344
rect 5029 1254 5062 1344
rect 5242 1254 5275 1344
rect 5477 1254 5510 1344
rect 5690 1254 5723 1344
rect 5925 1254 5958 1344
rect 6138 1254 6171 1344
rect 6373 1254 6406 1344
rect 6586 1254 6619 1344
rect 6821 1254 6854 1344
rect 7034 1254 7067 1344
rect 7269 1254 7302 1344
rect 7482 1254 7515 1344
rect 7717 1254 7750 1344
rect 7930 1254 7963 1344
rect 8165 1254 8198 1344
rect 8378 1254 8411 1344
rect 8613 1254 8646 1344
rect 8826 1254 8859 1344
rect 0 1222 448 1254
rect 549 1222 1691 1254
rect 1792 1222 2688 1254
rect 2789 1222 3931 1254
rect 4032 1222 4928 1254
rect 5029 1222 6171 1254
rect 6272 1222 7168 1254
rect 7269 1222 8411 1254
rect 8512 1222 8960 1254
rect 101 1131 134 1222
rect 314 1131 347 1222
rect 549 1131 582 1222
rect 762 1131 795 1222
rect 997 1131 1030 1222
rect 1210 1131 1243 1222
rect 1445 1131 1478 1222
rect 1658 1131 1691 1222
rect 1893 1131 1926 1222
rect 2106 1131 2139 1222
rect 2341 1131 2374 1222
rect 2554 1131 2587 1222
rect 2789 1131 2822 1222
rect 3002 1131 3035 1222
rect 3237 1131 3270 1222
rect 3450 1131 3483 1222
rect 3685 1131 3718 1222
rect 3898 1131 3931 1222
rect 4133 1131 4166 1222
rect 4346 1131 4379 1222
rect 4581 1131 4614 1222
rect 4794 1131 4827 1222
rect 5029 1131 5062 1222
rect 5242 1131 5275 1222
rect 5477 1131 5510 1222
rect 5690 1131 5723 1222
rect 5925 1131 5958 1222
rect 6138 1131 6171 1222
rect 6373 1131 6406 1222
rect 6586 1131 6619 1222
rect 6821 1131 6854 1222
rect 7034 1131 7067 1222
rect 7269 1131 7302 1222
rect 7482 1131 7515 1222
rect 7717 1131 7750 1222
rect 7930 1131 7963 1222
rect 8165 1131 8198 1222
rect 8378 1131 8411 1222
rect 8613 1131 8646 1222
rect 8826 1131 8859 1222
rect 99 1130 137 1131
rect 99 1129 102 1130
rect 54 1099 102 1129
rect 99 1098 102 1099
rect 134 1129 137 1130
rect 311 1130 349 1131
rect 311 1129 314 1130
rect 134 1099 181 1129
rect 267 1099 314 1129
rect 134 1098 137 1099
rect 99 1097 137 1098
rect 311 1098 314 1099
rect 346 1129 349 1130
rect 547 1130 585 1131
rect 547 1129 550 1130
rect 346 1099 394 1129
rect 502 1099 550 1129
rect 346 1098 349 1099
rect 311 1097 349 1098
rect 547 1098 550 1099
rect 582 1129 585 1130
rect 759 1130 797 1131
rect 759 1129 762 1130
rect 582 1099 629 1129
rect 715 1099 762 1129
rect 582 1098 585 1099
rect 547 1097 585 1098
rect 759 1098 762 1099
rect 794 1129 797 1130
rect 995 1130 1033 1131
rect 995 1129 998 1130
rect 794 1099 842 1129
rect 950 1099 998 1129
rect 794 1098 797 1099
rect 759 1097 797 1098
rect 995 1098 998 1099
rect 1030 1129 1033 1130
rect 1207 1130 1245 1131
rect 1207 1129 1210 1130
rect 1030 1099 1077 1129
rect 1163 1099 1210 1129
rect 1030 1098 1033 1099
rect 995 1097 1033 1098
rect 1207 1098 1210 1099
rect 1242 1129 1245 1130
rect 1443 1130 1481 1131
rect 1443 1129 1446 1130
rect 1242 1099 1290 1129
rect 1398 1099 1446 1129
rect 1242 1098 1245 1099
rect 1207 1097 1245 1098
rect 1443 1098 1446 1099
rect 1478 1129 1481 1130
rect 1655 1130 1693 1131
rect 1655 1129 1658 1130
rect 1478 1099 1525 1129
rect 1611 1099 1658 1129
rect 1478 1098 1481 1099
rect 1443 1097 1481 1098
rect 1655 1098 1658 1099
rect 1690 1129 1693 1130
rect 1891 1130 1929 1131
rect 1891 1129 1894 1130
rect 1690 1099 1738 1129
rect 1846 1099 1894 1129
rect 1690 1098 1693 1099
rect 1655 1097 1693 1098
rect 1891 1098 1894 1099
rect 1926 1129 1929 1130
rect 2103 1130 2141 1131
rect 2103 1129 2106 1130
rect 1926 1099 1973 1129
rect 2059 1099 2106 1129
rect 1926 1098 1929 1099
rect 1891 1097 1929 1098
rect 2103 1098 2106 1099
rect 2138 1129 2141 1130
rect 2339 1130 2377 1131
rect 2339 1129 2342 1130
rect 2138 1099 2186 1129
rect 2294 1099 2342 1129
rect 2138 1098 2141 1099
rect 2103 1097 2141 1098
rect 2339 1098 2342 1099
rect 2374 1129 2377 1130
rect 2551 1130 2589 1131
rect 2551 1129 2554 1130
rect 2374 1099 2421 1129
rect 2507 1099 2554 1129
rect 2374 1098 2377 1099
rect 2339 1097 2377 1098
rect 2551 1098 2554 1099
rect 2586 1129 2589 1130
rect 2787 1130 2825 1131
rect 2787 1129 2790 1130
rect 2586 1099 2634 1129
rect 2742 1099 2790 1129
rect 2586 1098 2589 1099
rect 2551 1097 2589 1098
rect 2787 1098 2790 1099
rect 2822 1129 2825 1130
rect 2999 1130 3037 1131
rect 2999 1129 3002 1130
rect 2822 1099 2869 1129
rect 2955 1099 3002 1129
rect 2822 1098 2825 1099
rect 2787 1097 2825 1098
rect 2999 1098 3002 1099
rect 3034 1129 3037 1130
rect 3235 1130 3273 1131
rect 3235 1129 3238 1130
rect 3034 1099 3082 1129
rect 3190 1099 3238 1129
rect 3034 1098 3037 1099
rect 2999 1097 3037 1098
rect 3235 1098 3238 1099
rect 3270 1129 3273 1130
rect 3447 1130 3485 1131
rect 3447 1129 3450 1130
rect 3270 1099 3317 1129
rect 3403 1099 3450 1129
rect 3270 1098 3273 1099
rect 3235 1097 3273 1098
rect 3447 1098 3450 1099
rect 3482 1129 3485 1130
rect 3683 1130 3721 1131
rect 3683 1129 3686 1130
rect 3482 1099 3530 1129
rect 3638 1099 3686 1129
rect 3482 1098 3485 1099
rect 3447 1097 3485 1098
rect 3683 1098 3686 1099
rect 3718 1129 3721 1130
rect 3895 1130 3933 1131
rect 3895 1129 3898 1130
rect 3718 1099 3765 1129
rect 3851 1099 3898 1129
rect 3718 1098 3721 1099
rect 3683 1097 3721 1098
rect 3895 1098 3898 1099
rect 3930 1129 3933 1130
rect 4131 1130 4169 1131
rect 4131 1129 4134 1130
rect 3930 1099 3978 1129
rect 4086 1099 4134 1129
rect 3930 1098 3933 1099
rect 3895 1097 3933 1098
rect 4131 1098 4134 1099
rect 4166 1129 4169 1130
rect 4343 1130 4381 1131
rect 4343 1129 4346 1130
rect 4166 1099 4213 1129
rect 4299 1099 4346 1129
rect 4166 1098 4169 1099
rect 4131 1097 4169 1098
rect 4343 1098 4346 1099
rect 4378 1129 4381 1130
rect 4579 1130 4617 1131
rect 4579 1129 4582 1130
rect 4378 1099 4426 1129
rect 4534 1099 4582 1129
rect 4378 1098 4381 1099
rect 4343 1097 4381 1098
rect 4579 1098 4582 1099
rect 4614 1129 4617 1130
rect 4791 1130 4829 1131
rect 4791 1129 4794 1130
rect 4614 1099 4661 1129
rect 4747 1099 4794 1129
rect 4614 1098 4617 1099
rect 4579 1097 4617 1098
rect 4791 1098 4794 1099
rect 4826 1129 4829 1130
rect 5027 1130 5065 1131
rect 5027 1129 5030 1130
rect 4826 1099 4874 1129
rect 4982 1099 5030 1129
rect 4826 1098 4829 1099
rect 4791 1097 4829 1098
rect 5027 1098 5030 1099
rect 5062 1129 5065 1130
rect 5239 1130 5277 1131
rect 5239 1129 5242 1130
rect 5062 1099 5109 1129
rect 5195 1099 5242 1129
rect 5062 1098 5065 1099
rect 5027 1097 5065 1098
rect 5239 1098 5242 1099
rect 5274 1129 5277 1130
rect 5475 1130 5513 1131
rect 5475 1129 5478 1130
rect 5274 1099 5322 1129
rect 5430 1099 5478 1129
rect 5274 1098 5277 1099
rect 5239 1097 5277 1098
rect 5475 1098 5478 1099
rect 5510 1129 5513 1130
rect 5687 1130 5725 1131
rect 5687 1129 5690 1130
rect 5510 1099 5557 1129
rect 5643 1099 5690 1129
rect 5510 1098 5513 1099
rect 5475 1097 5513 1098
rect 5687 1098 5690 1099
rect 5722 1129 5725 1130
rect 5923 1130 5961 1131
rect 5923 1129 5926 1130
rect 5722 1099 5770 1129
rect 5878 1099 5926 1129
rect 5722 1098 5725 1099
rect 5687 1097 5725 1098
rect 5923 1098 5926 1099
rect 5958 1129 5961 1130
rect 6135 1130 6173 1131
rect 6135 1129 6138 1130
rect 5958 1099 6005 1129
rect 6091 1099 6138 1129
rect 5958 1098 5961 1099
rect 5923 1097 5961 1098
rect 6135 1098 6138 1099
rect 6170 1129 6173 1130
rect 6371 1130 6409 1131
rect 6371 1129 6374 1130
rect 6170 1099 6218 1129
rect 6326 1099 6374 1129
rect 6170 1098 6173 1099
rect 6135 1097 6173 1098
rect 6371 1098 6374 1099
rect 6406 1129 6409 1130
rect 6583 1130 6621 1131
rect 6583 1129 6586 1130
rect 6406 1099 6453 1129
rect 6539 1099 6586 1129
rect 6406 1098 6409 1099
rect 6371 1097 6409 1098
rect 6583 1098 6586 1099
rect 6618 1129 6621 1130
rect 6819 1130 6857 1131
rect 6819 1129 6822 1130
rect 6618 1099 6666 1129
rect 6774 1099 6822 1129
rect 6618 1098 6621 1099
rect 6583 1097 6621 1098
rect 6819 1098 6822 1099
rect 6854 1129 6857 1130
rect 7031 1130 7069 1131
rect 7031 1129 7034 1130
rect 6854 1099 6901 1129
rect 6987 1099 7034 1129
rect 6854 1098 6857 1099
rect 6819 1097 6857 1098
rect 7031 1098 7034 1099
rect 7066 1129 7069 1130
rect 7267 1130 7305 1131
rect 7267 1129 7270 1130
rect 7066 1099 7114 1129
rect 7222 1099 7270 1129
rect 7066 1098 7069 1099
rect 7031 1097 7069 1098
rect 7267 1098 7270 1099
rect 7302 1129 7305 1130
rect 7479 1130 7517 1131
rect 7479 1129 7482 1130
rect 7302 1099 7349 1129
rect 7435 1099 7482 1129
rect 7302 1098 7305 1099
rect 7267 1097 7305 1098
rect 7479 1098 7482 1099
rect 7514 1129 7517 1130
rect 7715 1130 7753 1131
rect 7715 1129 7718 1130
rect 7514 1099 7562 1129
rect 7670 1099 7718 1129
rect 7514 1098 7517 1099
rect 7479 1097 7517 1098
rect 7715 1098 7718 1099
rect 7750 1129 7753 1130
rect 7927 1130 7965 1131
rect 7927 1129 7930 1130
rect 7750 1099 7797 1129
rect 7883 1099 7930 1129
rect 7750 1098 7753 1099
rect 7715 1097 7753 1098
rect 7927 1098 7930 1099
rect 7962 1129 7965 1130
rect 8163 1130 8201 1131
rect 8163 1129 8166 1130
rect 7962 1099 8010 1129
rect 8118 1099 8166 1129
rect 7962 1098 7965 1099
rect 7927 1097 7965 1098
rect 8163 1098 8166 1099
rect 8198 1129 8201 1130
rect 8375 1130 8413 1131
rect 8375 1129 8378 1130
rect 8198 1099 8245 1129
rect 8331 1099 8378 1129
rect 8198 1098 8201 1099
rect 8163 1097 8201 1098
rect 8375 1098 8378 1099
rect 8410 1129 8413 1130
rect 8611 1130 8649 1131
rect 8611 1129 8614 1130
rect 8410 1099 8458 1129
rect 8566 1099 8614 1129
rect 8410 1098 8413 1099
rect 8375 1097 8413 1098
rect 8611 1098 8614 1099
rect 8646 1129 8649 1130
rect 8823 1130 8861 1131
rect 8823 1129 8826 1130
rect 8646 1099 8693 1129
rect 8779 1099 8826 1129
rect 8646 1098 8649 1099
rect 8611 1097 8649 1098
rect 8823 1098 8826 1099
rect 8858 1129 8861 1130
rect 8858 1099 8906 1129
rect 8858 1098 8861 1099
rect 8823 1097 8861 1098
rect 101 1007 134 1097
rect 314 1007 347 1097
rect 549 1007 582 1097
rect 762 1007 795 1097
rect 997 1007 1030 1097
rect 1210 1007 1243 1097
rect 1445 1007 1478 1097
rect 1658 1007 1691 1097
rect 1893 1007 1926 1097
rect 2106 1007 2139 1097
rect 2341 1007 2374 1097
rect 2554 1007 2587 1097
rect 2789 1007 2822 1097
rect 3002 1007 3035 1097
rect 3237 1007 3270 1097
rect 3450 1007 3483 1097
rect 3685 1007 3718 1097
rect 3898 1007 3931 1097
rect 4133 1007 4166 1097
rect 4346 1007 4379 1097
rect 4581 1007 4614 1097
rect 4794 1007 4827 1097
rect 5029 1007 5062 1097
rect 5242 1007 5275 1097
rect 5477 1007 5510 1097
rect 5690 1007 5723 1097
rect 5925 1007 5958 1097
rect 6138 1007 6171 1097
rect 6373 1007 6406 1097
rect 6586 1007 6619 1097
rect 6821 1007 6854 1097
rect 7034 1007 7067 1097
rect 7269 1007 7302 1097
rect 7482 1007 7515 1097
rect 7717 1007 7750 1097
rect 7930 1007 7963 1097
rect 8165 1007 8198 1097
rect 8378 1007 8411 1097
rect 8613 1007 8646 1097
rect 8826 1007 8859 1097
rect 99 1006 137 1007
rect 99 1005 102 1006
rect 54 975 102 1005
rect 99 974 102 975
rect 134 1005 137 1006
rect 311 1006 349 1007
rect 311 1005 314 1006
rect 134 975 181 1005
rect 267 975 314 1005
rect 134 974 137 975
rect 99 973 137 974
rect 311 974 314 975
rect 346 1005 349 1006
rect 547 1006 585 1007
rect 547 1005 550 1006
rect 346 975 394 1005
rect 502 975 550 1005
rect 346 974 349 975
rect 311 973 349 974
rect 547 974 550 975
rect 582 1005 585 1006
rect 759 1006 797 1007
rect 759 1005 762 1006
rect 582 975 629 1005
rect 715 975 762 1005
rect 582 974 585 975
rect 547 973 585 974
rect 759 974 762 975
rect 794 1005 797 1006
rect 995 1006 1033 1007
rect 995 1005 998 1006
rect 794 975 842 1005
rect 950 975 998 1005
rect 794 974 797 975
rect 759 973 797 974
rect 995 974 998 975
rect 1030 1005 1033 1006
rect 1207 1006 1245 1007
rect 1207 1005 1210 1006
rect 1030 975 1077 1005
rect 1163 975 1210 1005
rect 1030 974 1033 975
rect 995 973 1033 974
rect 1207 974 1210 975
rect 1242 1005 1245 1006
rect 1443 1006 1481 1007
rect 1443 1005 1446 1006
rect 1242 975 1290 1005
rect 1398 975 1446 1005
rect 1242 974 1245 975
rect 1207 973 1245 974
rect 1443 974 1446 975
rect 1478 1005 1481 1006
rect 1655 1006 1693 1007
rect 1655 1005 1658 1006
rect 1478 975 1525 1005
rect 1611 975 1658 1005
rect 1478 974 1481 975
rect 1443 973 1481 974
rect 1655 974 1658 975
rect 1690 1005 1693 1006
rect 1891 1006 1929 1007
rect 1891 1005 1894 1006
rect 1690 975 1738 1005
rect 1846 975 1894 1005
rect 1690 974 1693 975
rect 1655 973 1693 974
rect 1891 974 1894 975
rect 1926 1005 1929 1006
rect 2103 1006 2141 1007
rect 2103 1005 2106 1006
rect 1926 975 1973 1005
rect 2059 975 2106 1005
rect 1926 974 1929 975
rect 1891 973 1929 974
rect 2103 974 2106 975
rect 2138 1005 2141 1006
rect 2339 1006 2377 1007
rect 2339 1005 2342 1006
rect 2138 975 2186 1005
rect 2294 975 2342 1005
rect 2138 974 2141 975
rect 2103 973 2141 974
rect 2339 974 2342 975
rect 2374 1005 2377 1006
rect 2551 1006 2589 1007
rect 2551 1005 2554 1006
rect 2374 975 2421 1005
rect 2507 975 2554 1005
rect 2374 974 2377 975
rect 2339 973 2377 974
rect 2551 974 2554 975
rect 2586 1005 2589 1006
rect 2787 1006 2825 1007
rect 2787 1005 2790 1006
rect 2586 975 2634 1005
rect 2742 975 2790 1005
rect 2586 974 2589 975
rect 2551 973 2589 974
rect 2787 974 2790 975
rect 2822 1005 2825 1006
rect 2999 1006 3037 1007
rect 2999 1005 3002 1006
rect 2822 975 2869 1005
rect 2955 975 3002 1005
rect 2822 974 2825 975
rect 2787 973 2825 974
rect 2999 974 3002 975
rect 3034 1005 3037 1006
rect 3235 1006 3273 1007
rect 3235 1005 3238 1006
rect 3034 975 3082 1005
rect 3190 975 3238 1005
rect 3034 974 3037 975
rect 2999 973 3037 974
rect 3235 974 3238 975
rect 3270 1005 3273 1006
rect 3447 1006 3485 1007
rect 3447 1005 3450 1006
rect 3270 975 3317 1005
rect 3403 975 3450 1005
rect 3270 974 3273 975
rect 3235 973 3273 974
rect 3447 974 3450 975
rect 3482 1005 3485 1006
rect 3683 1006 3721 1007
rect 3683 1005 3686 1006
rect 3482 975 3530 1005
rect 3638 975 3686 1005
rect 3482 974 3485 975
rect 3447 973 3485 974
rect 3683 974 3686 975
rect 3718 1005 3721 1006
rect 3895 1006 3933 1007
rect 3895 1005 3898 1006
rect 3718 975 3765 1005
rect 3851 975 3898 1005
rect 3718 974 3721 975
rect 3683 973 3721 974
rect 3895 974 3898 975
rect 3930 1005 3933 1006
rect 4131 1006 4169 1007
rect 4131 1005 4134 1006
rect 3930 975 3978 1005
rect 4086 975 4134 1005
rect 3930 974 3933 975
rect 3895 973 3933 974
rect 4131 974 4134 975
rect 4166 1005 4169 1006
rect 4343 1006 4381 1007
rect 4343 1005 4346 1006
rect 4166 975 4213 1005
rect 4299 975 4346 1005
rect 4166 974 4169 975
rect 4131 973 4169 974
rect 4343 974 4346 975
rect 4378 1005 4381 1006
rect 4579 1006 4617 1007
rect 4579 1005 4582 1006
rect 4378 975 4426 1005
rect 4534 975 4582 1005
rect 4378 974 4381 975
rect 4343 973 4381 974
rect 4579 974 4582 975
rect 4614 1005 4617 1006
rect 4791 1006 4829 1007
rect 4791 1005 4794 1006
rect 4614 975 4661 1005
rect 4747 975 4794 1005
rect 4614 974 4617 975
rect 4579 973 4617 974
rect 4791 974 4794 975
rect 4826 1005 4829 1006
rect 5027 1006 5065 1007
rect 5027 1005 5030 1006
rect 4826 975 4874 1005
rect 4982 975 5030 1005
rect 4826 974 4829 975
rect 4791 973 4829 974
rect 5027 974 5030 975
rect 5062 1005 5065 1006
rect 5239 1006 5277 1007
rect 5239 1005 5242 1006
rect 5062 975 5109 1005
rect 5195 975 5242 1005
rect 5062 974 5065 975
rect 5027 973 5065 974
rect 5239 974 5242 975
rect 5274 1005 5277 1006
rect 5475 1006 5513 1007
rect 5475 1005 5478 1006
rect 5274 975 5322 1005
rect 5430 975 5478 1005
rect 5274 974 5277 975
rect 5239 973 5277 974
rect 5475 974 5478 975
rect 5510 1005 5513 1006
rect 5687 1006 5725 1007
rect 5687 1005 5690 1006
rect 5510 975 5557 1005
rect 5643 975 5690 1005
rect 5510 974 5513 975
rect 5475 973 5513 974
rect 5687 974 5690 975
rect 5722 1005 5725 1006
rect 5923 1006 5961 1007
rect 5923 1005 5926 1006
rect 5722 975 5770 1005
rect 5878 975 5926 1005
rect 5722 974 5725 975
rect 5687 973 5725 974
rect 5923 974 5926 975
rect 5958 1005 5961 1006
rect 6135 1006 6173 1007
rect 6135 1005 6138 1006
rect 5958 975 6005 1005
rect 6091 975 6138 1005
rect 5958 974 5961 975
rect 5923 973 5961 974
rect 6135 974 6138 975
rect 6170 1005 6173 1006
rect 6371 1006 6409 1007
rect 6371 1005 6374 1006
rect 6170 975 6218 1005
rect 6326 975 6374 1005
rect 6170 974 6173 975
rect 6135 973 6173 974
rect 6371 974 6374 975
rect 6406 1005 6409 1006
rect 6583 1006 6621 1007
rect 6583 1005 6586 1006
rect 6406 975 6453 1005
rect 6539 975 6586 1005
rect 6406 974 6409 975
rect 6371 973 6409 974
rect 6583 974 6586 975
rect 6618 1005 6621 1006
rect 6819 1006 6857 1007
rect 6819 1005 6822 1006
rect 6618 975 6666 1005
rect 6774 975 6822 1005
rect 6618 974 6621 975
rect 6583 973 6621 974
rect 6819 974 6822 975
rect 6854 1005 6857 1006
rect 7031 1006 7069 1007
rect 7031 1005 7034 1006
rect 6854 975 6901 1005
rect 6987 975 7034 1005
rect 6854 974 6857 975
rect 6819 973 6857 974
rect 7031 974 7034 975
rect 7066 1005 7069 1006
rect 7267 1006 7305 1007
rect 7267 1005 7270 1006
rect 7066 975 7114 1005
rect 7222 975 7270 1005
rect 7066 974 7069 975
rect 7031 973 7069 974
rect 7267 974 7270 975
rect 7302 1005 7305 1006
rect 7479 1006 7517 1007
rect 7479 1005 7482 1006
rect 7302 975 7349 1005
rect 7435 975 7482 1005
rect 7302 974 7305 975
rect 7267 973 7305 974
rect 7479 974 7482 975
rect 7514 1005 7517 1006
rect 7715 1006 7753 1007
rect 7715 1005 7718 1006
rect 7514 975 7562 1005
rect 7670 975 7718 1005
rect 7514 974 7517 975
rect 7479 973 7517 974
rect 7715 974 7718 975
rect 7750 1005 7753 1006
rect 7927 1006 7965 1007
rect 7927 1005 7930 1006
rect 7750 975 7797 1005
rect 7883 975 7930 1005
rect 7750 974 7753 975
rect 7715 973 7753 974
rect 7927 974 7930 975
rect 7962 1005 7965 1006
rect 8163 1006 8201 1007
rect 8163 1005 8166 1006
rect 7962 975 8010 1005
rect 8118 975 8166 1005
rect 7962 974 7965 975
rect 7927 973 7965 974
rect 8163 974 8166 975
rect 8198 1005 8201 1006
rect 8375 1006 8413 1007
rect 8375 1005 8378 1006
rect 8198 975 8245 1005
rect 8331 975 8378 1005
rect 8198 974 8201 975
rect 8163 973 8201 974
rect 8375 974 8378 975
rect 8410 1005 8413 1006
rect 8611 1006 8649 1007
rect 8611 1005 8614 1006
rect 8410 975 8458 1005
rect 8566 975 8614 1005
rect 8410 974 8413 975
rect 8375 973 8413 974
rect 8611 974 8614 975
rect 8646 1005 8649 1006
rect 8823 1006 8861 1007
rect 8823 1005 8826 1006
rect 8646 975 8693 1005
rect 8779 975 8826 1005
rect 8646 974 8649 975
rect 8611 973 8649 974
rect 8823 974 8826 975
rect 8858 1005 8861 1006
rect 8858 975 8906 1005
rect 8858 974 8861 975
rect 8823 973 8861 974
rect 101 883 134 973
rect 314 883 347 973
rect 549 883 582 973
rect 762 883 795 973
rect 997 883 1030 973
rect 1210 883 1243 973
rect 1445 883 1478 973
rect 1658 883 1691 973
rect 1893 883 1926 973
rect 2106 883 2139 973
rect 2341 883 2374 973
rect 2554 883 2587 973
rect 2789 883 2822 973
rect 3002 883 3035 973
rect 3237 883 3270 973
rect 3450 883 3483 973
rect 3685 883 3718 973
rect 3898 883 3931 973
rect 4133 883 4166 973
rect 4346 883 4379 973
rect 4581 883 4614 973
rect 4794 883 4827 973
rect 5029 883 5062 973
rect 5242 883 5275 973
rect 5477 883 5510 973
rect 5690 883 5723 973
rect 5925 883 5958 973
rect 6138 883 6171 973
rect 6373 883 6406 973
rect 6586 883 6619 973
rect 6821 883 6854 973
rect 7034 883 7067 973
rect 7269 883 7302 973
rect 7482 883 7515 973
rect 7717 883 7750 973
rect 7930 883 7963 973
rect 8165 883 8198 973
rect 8378 883 8411 973
rect 8613 883 8646 973
rect 8826 883 8859 973
rect 99 882 137 883
rect 99 881 102 882
rect 54 851 102 881
rect 99 850 102 851
rect 134 881 137 882
rect 311 882 349 883
rect 311 881 314 882
rect 134 851 181 881
rect 267 851 314 881
rect 134 850 137 851
rect 99 849 137 850
rect 311 850 314 851
rect 346 881 349 882
rect 547 882 585 883
rect 547 881 550 882
rect 346 851 394 881
rect 502 851 550 881
rect 346 850 349 851
rect 311 849 349 850
rect 547 850 550 851
rect 582 881 585 882
rect 759 882 797 883
rect 759 881 762 882
rect 582 851 629 881
rect 715 851 762 881
rect 582 850 585 851
rect 547 849 585 850
rect 759 850 762 851
rect 794 881 797 882
rect 995 882 1033 883
rect 995 881 998 882
rect 794 851 842 881
rect 950 851 998 881
rect 794 850 797 851
rect 759 849 797 850
rect 995 850 998 851
rect 1030 881 1033 882
rect 1207 882 1245 883
rect 1207 881 1210 882
rect 1030 851 1077 881
rect 1163 851 1210 881
rect 1030 850 1033 851
rect 995 849 1033 850
rect 1207 850 1210 851
rect 1242 881 1245 882
rect 1443 882 1481 883
rect 1443 881 1446 882
rect 1242 851 1290 881
rect 1398 851 1446 881
rect 1242 850 1245 851
rect 1207 849 1245 850
rect 1443 850 1446 851
rect 1478 881 1481 882
rect 1655 882 1693 883
rect 1655 881 1658 882
rect 1478 851 1525 881
rect 1611 851 1658 881
rect 1478 850 1481 851
rect 1443 849 1481 850
rect 1655 850 1658 851
rect 1690 881 1693 882
rect 1891 882 1929 883
rect 1891 881 1894 882
rect 1690 851 1738 881
rect 1846 851 1894 881
rect 1690 850 1693 851
rect 1655 849 1693 850
rect 1891 850 1894 851
rect 1926 881 1929 882
rect 2103 882 2141 883
rect 2103 881 2106 882
rect 1926 851 1973 881
rect 2059 851 2106 881
rect 1926 850 1929 851
rect 1891 849 1929 850
rect 2103 850 2106 851
rect 2138 881 2141 882
rect 2339 882 2377 883
rect 2339 881 2342 882
rect 2138 851 2186 881
rect 2294 851 2342 881
rect 2138 850 2141 851
rect 2103 849 2141 850
rect 2339 850 2342 851
rect 2374 881 2377 882
rect 2551 882 2589 883
rect 2551 881 2554 882
rect 2374 851 2421 881
rect 2507 851 2554 881
rect 2374 850 2377 851
rect 2339 849 2377 850
rect 2551 850 2554 851
rect 2586 881 2589 882
rect 2787 882 2825 883
rect 2787 881 2790 882
rect 2586 851 2634 881
rect 2742 851 2790 881
rect 2586 850 2589 851
rect 2551 849 2589 850
rect 2787 850 2790 851
rect 2822 881 2825 882
rect 2999 882 3037 883
rect 2999 881 3002 882
rect 2822 851 2869 881
rect 2955 851 3002 881
rect 2822 850 2825 851
rect 2787 849 2825 850
rect 2999 850 3002 851
rect 3034 881 3037 882
rect 3235 882 3273 883
rect 3235 881 3238 882
rect 3034 851 3082 881
rect 3190 851 3238 881
rect 3034 850 3037 851
rect 2999 849 3037 850
rect 3235 850 3238 851
rect 3270 881 3273 882
rect 3447 882 3485 883
rect 3447 881 3450 882
rect 3270 851 3317 881
rect 3403 851 3450 881
rect 3270 850 3273 851
rect 3235 849 3273 850
rect 3447 850 3450 851
rect 3482 881 3485 882
rect 3683 882 3721 883
rect 3683 881 3686 882
rect 3482 851 3530 881
rect 3638 851 3686 881
rect 3482 850 3485 851
rect 3447 849 3485 850
rect 3683 850 3686 851
rect 3718 881 3721 882
rect 3895 882 3933 883
rect 3895 881 3898 882
rect 3718 851 3765 881
rect 3851 851 3898 881
rect 3718 850 3721 851
rect 3683 849 3721 850
rect 3895 850 3898 851
rect 3930 881 3933 882
rect 4131 882 4169 883
rect 4131 881 4134 882
rect 3930 851 3978 881
rect 4086 851 4134 881
rect 3930 850 3933 851
rect 3895 849 3933 850
rect 4131 850 4134 851
rect 4166 881 4169 882
rect 4343 882 4381 883
rect 4343 881 4346 882
rect 4166 851 4213 881
rect 4299 851 4346 881
rect 4166 850 4169 851
rect 4131 849 4169 850
rect 4343 850 4346 851
rect 4378 881 4381 882
rect 4579 882 4617 883
rect 4579 881 4582 882
rect 4378 851 4426 881
rect 4534 851 4582 881
rect 4378 850 4381 851
rect 4343 849 4381 850
rect 4579 850 4582 851
rect 4614 881 4617 882
rect 4791 882 4829 883
rect 4791 881 4794 882
rect 4614 851 4661 881
rect 4747 851 4794 881
rect 4614 850 4617 851
rect 4579 849 4617 850
rect 4791 850 4794 851
rect 4826 881 4829 882
rect 5027 882 5065 883
rect 5027 881 5030 882
rect 4826 851 4874 881
rect 4982 851 5030 881
rect 4826 850 4829 851
rect 4791 849 4829 850
rect 5027 850 5030 851
rect 5062 881 5065 882
rect 5239 882 5277 883
rect 5239 881 5242 882
rect 5062 851 5109 881
rect 5195 851 5242 881
rect 5062 850 5065 851
rect 5027 849 5065 850
rect 5239 850 5242 851
rect 5274 881 5277 882
rect 5475 882 5513 883
rect 5475 881 5478 882
rect 5274 851 5322 881
rect 5430 851 5478 881
rect 5274 850 5277 851
rect 5239 849 5277 850
rect 5475 850 5478 851
rect 5510 881 5513 882
rect 5687 882 5725 883
rect 5687 881 5690 882
rect 5510 851 5557 881
rect 5643 851 5690 881
rect 5510 850 5513 851
rect 5475 849 5513 850
rect 5687 850 5690 851
rect 5722 881 5725 882
rect 5923 882 5961 883
rect 5923 881 5926 882
rect 5722 851 5770 881
rect 5878 851 5926 881
rect 5722 850 5725 851
rect 5687 849 5725 850
rect 5923 850 5926 851
rect 5958 881 5961 882
rect 6135 882 6173 883
rect 6135 881 6138 882
rect 5958 851 6005 881
rect 6091 851 6138 881
rect 5958 850 5961 851
rect 5923 849 5961 850
rect 6135 850 6138 851
rect 6170 881 6173 882
rect 6371 882 6409 883
rect 6371 881 6374 882
rect 6170 851 6218 881
rect 6326 851 6374 881
rect 6170 850 6173 851
rect 6135 849 6173 850
rect 6371 850 6374 851
rect 6406 881 6409 882
rect 6583 882 6621 883
rect 6583 881 6586 882
rect 6406 851 6453 881
rect 6539 851 6586 881
rect 6406 850 6409 851
rect 6371 849 6409 850
rect 6583 850 6586 851
rect 6618 881 6621 882
rect 6819 882 6857 883
rect 6819 881 6822 882
rect 6618 851 6666 881
rect 6774 851 6822 881
rect 6618 850 6621 851
rect 6583 849 6621 850
rect 6819 850 6822 851
rect 6854 881 6857 882
rect 7031 882 7069 883
rect 7031 881 7034 882
rect 6854 851 6901 881
rect 6987 851 7034 881
rect 6854 850 6857 851
rect 6819 849 6857 850
rect 7031 850 7034 851
rect 7066 881 7069 882
rect 7267 882 7305 883
rect 7267 881 7270 882
rect 7066 851 7114 881
rect 7222 851 7270 881
rect 7066 850 7069 851
rect 7031 849 7069 850
rect 7267 850 7270 851
rect 7302 881 7305 882
rect 7479 882 7517 883
rect 7479 881 7482 882
rect 7302 851 7349 881
rect 7435 851 7482 881
rect 7302 850 7305 851
rect 7267 849 7305 850
rect 7479 850 7482 851
rect 7514 881 7517 882
rect 7715 882 7753 883
rect 7715 881 7718 882
rect 7514 851 7562 881
rect 7670 851 7718 881
rect 7514 850 7517 851
rect 7479 849 7517 850
rect 7715 850 7718 851
rect 7750 881 7753 882
rect 7927 882 7965 883
rect 7927 881 7930 882
rect 7750 851 7797 881
rect 7883 851 7930 881
rect 7750 850 7753 851
rect 7715 849 7753 850
rect 7927 850 7930 851
rect 7962 881 7965 882
rect 8163 882 8201 883
rect 8163 881 8166 882
rect 7962 851 8010 881
rect 8118 851 8166 881
rect 7962 850 7965 851
rect 7927 849 7965 850
rect 8163 850 8166 851
rect 8198 881 8201 882
rect 8375 882 8413 883
rect 8375 881 8378 882
rect 8198 851 8245 881
rect 8331 851 8378 881
rect 8198 850 8201 851
rect 8163 849 8201 850
rect 8375 850 8378 851
rect 8410 881 8413 882
rect 8611 882 8649 883
rect 8611 881 8614 882
rect 8410 851 8458 881
rect 8566 851 8614 881
rect 8410 850 8413 851
rect 8375 849 8413 850
rect 8611 850 8614 851
rect 8646 881 8649 882
rect 8823 882 8861 883
rect 8823 881 8826 882
rect 8646 851 8693 881
rect 8779 851 8826 881
rect 8646 850 8649 851
rect 8611 849 8649 850
rect 8823 850 8826 851
rect 8858 881 8861 882
rect 8858 851 8906 881
rect 8858 850 8861 851
rect 8823 849 8861 850
rect 101 759 134 849
rect 314 759 347 849
rect 549 759 582 849
rect 762 759 795 849
rect 997 759 1030 849
rect 1210 759 1243 849
rect 1445 759 1478 849
rect 1658 759 1691 849
rect 1893 759 1926 849
rect 2106 759 2139 849
rect 2341 759 2374 849
rect 2554 759 2587 849
rect 2789 759 2822 849
rect 3002 759 3035 849
rect 3237 759 3270 849
rect 3450 759 3483 849
rect 3685 759 3718 849
rect 3898 759 3931 849
rect 4133 759 4166 849
rect 4346 759 4379 849
rect 4581 759 4614 849
rect 4794 759 4827 849
rect 5029 759 5062 849
rect 5242 759 5275 849
rect 5477 759 5510 849
rect 5690 759 5723 849
rect 5925 759 5958 849
rect 6138 759 6171 849
rect 6373 759 6406 849
rect 6586 759 6619 849
rect 6821 759 6854 849
rect 7034 759 7067 849
rect 7269 759 7302 849
rect 7482 759 7515 849
rect 7717 759 7750 849
rect 7930 759 7963 849
rect 8165 759 8198 849
rect 8378 759 8411 849
rect 8613 759 8646 849
rect 8826 759 8859 849
rect 99 758 137 759
rect 99 757 102 758
rect 54 727 102 757
rect 99 726 102 727
rect 134 757 137 758
rect 311 758 349 759
rect 311 757 314 758
rect 134 727 181 757
rect 267 727 314 757
rect 134 726 137 727
rect 99 725 137 726
rect 311 726 314 727
rect 346 757 349 758
rect 547 758 585 759
rect 547 757 550 758
rect 346 727 394 757
rect 502 727 550 757
rect 346 726 349 727
rect 311 725 349 726
rect 547 726 550 727
rect 582 757 585 758
rect 759 758 797 759
rect 759 757 762 758
rect 582 727 629 757
rect 715 727 762 757
rect 582 726 585 727
rect 547 725 585 726
rect 759 726 762 727
rect 794 757 797 758
rect 995 758 1033 759
rect 995 757 998 758
rect 794 727 842 757
rect 950 727 998 757
rect 794 726 797 727
rect 759 725 797 726
rect 995 726 998 727
rect 1030 757 1033 758
rect 1207 758 1245 759
rect 1207 757 1210 758
rect 1030 727 1077 757
rect 1163 727 1210 757
rect 1030 726 1033 727
rect 995 725 1033 726
rect 1207 726 1210 727
rect 1242 757 1245 758
rect 1443 758 1481 759
rect 1443 757 1446 758
rect 1242 727 1290 757
rect 1398 727 1446 757
rect 1242 726 1245 727
rect 1207 725 1245 726
rect 1443 726 1446 727
rect 1478 757 1481 758
rect 1655 758 1693 759
rect 1655 757 1658 758
rect 1478 727 1525 757
rect 1611 727 1658 757
rect 1478 726 1481 727
rect 1443 725 1481 726
rect 1655 726 1658 727
rect 1690 757 1693 758
rect 1891 758 1929 759
rect 1891 757 1894 758
rect 1690 727 1738 757
rect 1846 727 1894 757
rect 1690 726 1693 727
rect 1655 725 1693 726
rect 1891 726 1894 727
rect 1926 757 1929 758
rect 2103 758 2141 759
rect 2103 757 2106 758
rect 1926 727 1973 757
rect 2059 727 2106 757
rect 1926 726 1929 727
rect 1891 725 1929 726
rect 2103 726 2106 727
rect 2138 757 2141 758
rect 2339 758 2377 759
rect 2339 757 2342 758
rect 2138 727 2186 757
rect 2294 727 2342 757
rect 2138 726 2141 727
rect 2103 725 2141 726
rect 2339 726 2342 727
rect 2374 757 2377 758
rect 2551 758 2589 759
rect 2551 757 2554 758
rect 2374 727 2421 757
rect 2507 727 2554 757
rect 2374 726 2377 727
rect 2339 725 2377 726
rect 2551 726 2554 727
rect 2586 757 2589 758
rect 2787 758 2825 759
rect 2787 757 2790 758
rect 2586 727 2634 757
rect 2742 727 2790 757
rect 2586 726 2589 727
rect 2551 725 2589 726
rect 2787 726 2790 727
rect 2822 757 2825 758
rect 2999 758 3037 759
rect 2999 757 3002 758
rect 2822 727 2869 757
rect 2955 727 3002 757
rect 2822 726 2825 727
rect 2787 725 2825 726
rect 2999 726 3002 727
rect 3034 757 3037 758
rect 3235 758 3273 759
rect 3235 757 3238 758
rect 3034 727 3082 757
rect 3190 727 3238 757
rect 3034 726 3037 727
rect 2999 725 3037 726
rect 3235 726 3238 727
rect 3270 757 3273 758
rect 3447 758 3485 759
rect 3447 757 3450 758
rect 3270 727 3317 757
rect 3403 727 3450 757
rect 3270 726 3273 727
rect 3235 725 3273 726
rect 3447 726 3450 727
rect 3482 757 3485 758
rect 3683 758 3721 759
rect 3683 757 3686 758
rect 3482 727 3530 757
rect 3638 727 3686 757
rect 3482 726 3485 727
rect 3447 725 3485 726
rect 3683 726 3686 727
rect 3718 757 3721 758
rect 3895 758 3933 759
rect 3895 757 3898 758
rect 3718 727 3765 757
rect 3851 727 3898 757
rect 3718 726 3721 727
rect 3683 725 3721 726
rect 3895 726 3898 727
rect 3930 757 3933 758
rect 4131 758 4169 759
rect 4131 757 4134 758
rect 3930 727 3978 757
rect 4086 727 4134 757
rect 3930 726 3933 727
rect 3895 725 3933 726
rect 4131 726 4134 727
rect 4166 757 4169 758
rect 4343 758 4381 759
rect 4343 757 4346 758
rect 4166 727 4213 757
rect 4299 727 4346 757
rect 4166 726 4169 727
rect 4131 725 4169 726
rect 4343 726 4346 727
rect 4378 757 4381 758
rect 4579 758 4617 759
rect 4579 757 4582 758
rect 4378 727 4426 757
rect 4534 727 4582 757
rect 4378 726 4381 727
rect 4343 725 4381 726
rect 4579 726 4582 727
rect 4614 757 4617 758
rect 4791 758 4829 759
rect 4791 757 4794 758
rect 4614 727 4661 757
rect 4747 727 4794 757
rect 4614 726 4617 727
rect 4579 725 4617 726
rect 4791 726 4794 727
rect 4826 757 4829 758
rect 5027 758 5065 759
rect 5027 757 5030 758
rect 4826 727 4874 757
rect 4982 727 5030 757
rect 4826 726 4829 727
rect 4791 725 4829 726
rect 5027 726 5030 727
rect 5062 757 5065 758
rect 5239 758 5277 759
rect 5239 757 5242 758
rect 5062 727 5109 757
rect 5195 727 5242 757
rect 5062 726 5065 727
rect 5027 725 5065 726
rect 5239 726 5242 727
rect 5274 757 5277 758
rect 5475 758 5513 759
rect 5475 757 5478 758
rect 5274 727 5322 757
rect 5430 727 5478 757
rect 5274 726 5277 727
rect 5239 725 5277 726
rect 5475 726 5478 727
rect 5510 757 5513 758
rect 5687 758 5725 759
rect 5687 757 5690 758
rect 5510 727 5557 757
rect 5643 727 5690 757
rect 5510 726 5513 727
rect 5475 725 5513 726
rect 5687 726 5690 727
rect 5722 757 5725 758
rect 5923 758 5961 759
rect 5923 757 5926 758
rect 5722 727 5770 757
rect 5878 727 5926 757
rect 5722 726 5725 727
rect 5687 725 5725 726
rect 5923 726 5926 727
rect 5958 757 5961 758
rect 6135 758 6173 759
rect 6135 757 6138 758
rect 5958 727 6005 757
rect 6091 727 6138 757
rect 5958 726 5961 727
rect 5923 725 5961 726
rect 6135 726 6138 727
rect 6170 757 6173 758
rect 6371 758 6409 759
rect 6371 757 6374 758
rect 6170 727 6218 757
rect 6326 727 6374 757
rect 6170 726 6173 727
rect 6135 725 6173 726
rect 6371 726 6374 727
rect 6406 757 6409 758
rect 6583 758 6621 759
rect 6583 757 6586 758
rect 6406 727 6453 757
rect 6539 727 6586 757
rect 6406 726 6409 727
rect 6371 725 6409 726
rect 6583 726 6586 727
rect 6618 757 6621 758
rect 6819 758 6857 759
rect 6819 757 6822 758
rect 6618 727 6666 757
rect 6774 727 6822 757
rect 6618 726 6621 727
rect 6583 725 6621 726
rect 6819 726 6822 727
rect 6854 757 6857 758
rect 7031 758 7069 759
rect 7031 757 7034 758
rect 6854 727 6901 757
rect 6987 727 7034 757
rect 6854 726 6857 727
rect 6819 725 6857 726
rect 7031 726 7034 727
rect 7066 757 7069 758
rect 7267 758 7305 759
rect 7267 757 7270 758
rect 7066 727 7114 757
rect 7222 727 7270 757
rect 7066 726 7069 727
rect 7031 725 7069 726
rect 7267 726 7270 727
rect 7302 757 7305 758
rect 7479 758 7517 759
rect 7479 757 7482 758
rect 7302 727 7349 757
rect 7435 727 7482 757
rect 7302 726 7305 727
rect 7267 725 7305 726
rect 7479 726 7482 727
rect 7514 757 7517 758
rect 7715 758 7753 759
rect 7715 757 7718 758
rect 7514 727 7562 757
rect 7670 727 7718 757
rect 7514 726 7517 727
rect 7479 725 7517 726
rect 7715 726 7718 727
rect 7750 757 7753 758
rect 7927 758 7965 759
rect 7927 757 7930 758
rect 7750 727 7797 757
rect 7883 727 7930 757
rect 7750 726 7753 727
rect 7715 725 7753 726
rect 7927 726 7930 727
rect 7962 757 7965 758
rect 8163 758 8201 759
rect 8163 757 8166 758
rect 7962 727 8010 757
rect 8118 727 8166 757
rect 7962 726 7965 727
rect 7927 725 7965 726
rect 8163 726 8166 727
rect 8198 757 8201 758
rect 8375 758 8413 759
rect 8375 757 8378 758
rect 8198 727 8245 757
rect 8331 727 8378 757
rect 8198 726 8201 727
rect 8163 725 8201 726
rect 8375 726 8378 727
rect 8410 757 8413 758
rect 8611 758 8649 759
rect 8611 757 8614 758
rect 8410 727 8458 757
rect 8566 727 8614 757
rect 8410 726 8413 727
rect 8375 725 8413 726
rect 8611 726 8614 727
rect 8646 757 8649 758
rect 8823 758 8861 759
rect 8823 757 8826 758
rect 8646 727 8693 757
rect 8779 727 8826 757
rect 8646 726 8649 727
rect 8611 725 8649 726
rect 8823 726 8826 727
rect 8858 757 8861 758
rect 8858 727 8906 757
rect 8858 726 8861 727
rect 8823 725 8861 726
rect 101 635 134 725
rect 314 635 347 725
rect 549 635 582 725
rect 762 635 795 725
rect 997 635 1030 725
rect 1210 635 1243 725
rect 1445 635 1478 725
rect 1658 635 1691 725
rect 1893 635 1926 725
rect 2106 635 2139 725
rect 2341 635 2374 725
rect 2554 635 2587 725
rect 2789 635 2822 725
rect 3002 635 3035 725
rect 3237 635 3270 725
rect 3450 635 3483 725
rect 3685 635 3718 725
rect 3898 635 3931 725
rect 4133 635 4166 725
rect 4346 635 4379 725
rect 4581 635 4614 725
rect 4794 635 4827 725
rect 5029 635 5062 725
rect 5242 635 5275 725
rect 5477 635 5510 725
rect 5690 635 5723 725
rect 5925 635 5958 725
rect 6138 635 6171 725
rect 6373 635 6406 725
rect 6586 635 6619 725
rect 6821 635 6854 725
rect 7034 635 7067 725
rect 7269 635 7302 725
rect 7482 635 7515 725
rect 7717 635 7750 725
rect 7930 635 7963 725
rect 8165 635 8198 725
rect 8378 635 8411 725
rect 8613 635 8646 725
rect 8826 635 8859 725
rect 0 603 448 635
rect 549 603 1691 635
rect 1792 603 2688 635
rect 2789 603 3931 635
rect 4032 603 4928 635
rect 5029 603 6171 635
rect 6272 603 7168 635
rect 7269 603 8411 635
rect 8512 603 8960 635
rect 101 512 134 603
rect 314 512 347 603
rect 549 512 582 559
rect 762 512 795 559
rect 997 512 1030 559
rect 1210 512 1243 559
rect 1445 512 1478 559
rect 1658 512 1691 559
rect 1893 512 1926 603
rect 2106 512 2139 603
rect 2341 512 2374 603
rect 2554 512 2587 603
rect 2789 512 2822 559
rect 3002 512 3035 559
rect 3237 512 3270 603
rect 3450 512 3483 603
rect 3685 512 3718 559
rect 3898 512 3931 559
rect 4133 512 4166 603
rect 4346 512 4379 603
rect 4581 512 4614 603
rect 4794 512 4827 603
rect 5029 512 5062 559
rect 5242 512 5275 559
rect 5477 512 5510 603
rect 5690 512 5723 603
rect 5925 512 5958 559
rect 6138 512 6171 559
rect 6373 512 6406 603
rect 6586 512 6619 603
rect 6821 512 6854 603
rect 7034 512 7067 603
rect 7269 512 7302 559
rect 7482 512 7515 559
rect 7717 512 7750 603
rect 7930 512 7963 559
rect 8165 512 8198 559
rect 8378 512 8411 559
rect 8613 512 8646 603
rect 8826 512 8859 603
rect 99 511 137 512
rect 99 510 102 511
rect 54 480 102 510
rect 99 479 102 480
rect 134 510 137 511
rect 311 511 349 512
rect 311 510 314 511
rect 134 480 181 510
rect 267 480 314 510
rect 134 479 137 480
rect 99 478 137 479
rect 311 479 314 480
rect 346 510 349 511
rect 547 511 585 512
rect 547 510 550 511
rect 346 480 394 510
rect 502 480 550 510
rect 346 479 349 480
rect 311 478 349 479
rect 547 479 550 480
rect 582 510 585 511
rect 759 511 797 512
rect 759 510 762 511
rect 582 480 629 510
rect 715 480 762 510
rect 582 479 585 480
rect 547 478 585 479
rect 759 479 762 480
rect 794 510 797 511
rect 995 511 1033 512
rect 995 510 998 511
rect 794 480 842 510
rect 950 480 998 510
rect 794 479 797 480
rect 759 478 797 479
rect 995 479 998 480
rect 1030 510 1033 511
rect 1207 511 1245 512
rect 1207 510 1210 511
rect 1030 480 1077 510
rect 1163 480 1210 510
rect 1030 479 1033 480
rect 995 478 1033 479
rect 1207 479 1210 480
rect 1242 510 1245 511
rect 1443 511 1481 512
rect 1443 510 1446 511
rect 1242 480 1290 510
rect 1398 480 1446 510
rect 1242 479 1245 480
rect 1207 478 1245 479
rect 1443 479 1446 480
rect 1478 510 1481 511
rect 1655 511 1693 512
rect 1655 510 1658 511
rect 1478 480 1525 510
rect 1611 480 1658 510
rect 1478 479 1481 480
rect 1443 478 1481 479
rect 1655 479 1658 480
rect 1690 510 1693 511
rect 1891 511 1929 512
rect 1891 510 1894 511
rect 1690 480 1738 510
rect 1846 480 1894 510
rect 1690 479 1693 480
rect 1655 478 1693 479
rect 1891 479 1894 480
rect 1926 510 1929 511
rect 2103 511 2141 512
rect 2103 510 2106 511
rect 1926 480 1973 510
rect 2059 480 2106 510
rect 1926 479 1929 480
rect 1891 478 1929 479
rect 2103 479 2106 480
rect 2138 510 2141 511
rect 2339 511 2377 512
rect 2339 510 2342 511
rect 2138 480 2186 510
rect 2294 480 2342 510
rect 2138 479 2141 480
rect 2103 478 2141 479
rect 2339 479 2342 480
rect 2374 510 2377 511
rect 2551 511 2589 512
rect 2551 510 2554 511
rect 2374 480 2421 510
rect 2507 480 2554 510
rect 2374 479 2377 480
rect 2339 478 2377 479
rect 2551 479 2554 480
rect 2586 510 2589 511
rect 2787 511 2825 512
rect 2787 510 2790 511
rect 2586 480 2634 510
rect 2742 480 2790 510
rect 2586 479 2589 480
rect 2551 478 2589 479
rect 2787 479 2790 480
rect 2822 510 2825 511
rect 2999 511 3037 512
rect 2999 510 3002 511
rect 2822 480 2869 510
rect 2955 480 3002 510
rect 2822 479 2825 480
rect 2787 478 2825 479
rect 2999 479 3002 480
rect 3034 510 3037 511
rect 3235 511 3273 512
rect 3235 510 3238 511
rect 3034 480 3082 510
rect 3190 480 3238 510
rect 3034 479 3037 480
rect 2999 478 3037 479
rect 3235 479 3238 480
rect 3270 510 3273 511
rect 3447 511 3485 512
rect 3447 510 3450 511
rect 3270 480 3317 510
rect 3403 480 3450 510
rect 3270 479 3273 480
rect 3235 478 3273 479
rect 3447 479 3450 480
rect 3482 510 3485 511
rect 3683 511 3721 512
rect 3683 510 3686 511
rect 3482 480 3530 510
rect 3638 480 3686 510
rect 3482 479 3485 480
rect 3447 478 3485 479
rect 3683 479 3686 480
rect 3718 510 3721 511
rect 3895 511 3933 512
rect 3895 510 3898 511
rect 3718 480 3765 510
rect 3851 480 3898 510
rect 3718 479 3721 480
rect 3683 478 3721 479
rect 3895 479 3898 480
rect 3930 510 3933 511
rect 4131 511 4169 512
rect 4131 510 4134 511
rect 3930 480 3978 510
rect 4086 480 4134 510
rect 3930 479 3933 480
rect 3895 478 3933 479
rect 4131 479 4134 480
rect 4166 510 4169 511
rect 4343 511 4381 512
rect 4343 510 4346 511
rect 4166 480 4213 510
rect 4299 480 4346 510
rect 4166 479 4169 480
rect 4131 478 4169 479
rect 4343 479 4346 480
rect 4378 510 4381 511
rect 4579 511 4617 512
rect 4579 510 4582 511
rect 4378 480 4426 510
rect 4534 480 4582 510
rect 4378 479 4381 480
rect 4343 478 4381 479
rect 4579 479 4582 480
rect 4614 510 4617 511
rect 4791 511 4829 512
rect 4791 510 4794 511
rect 4614 480 4661 510
rect 4747 480 4794 510
rect 4614 479 4617 480
rect 4579 478 4617 479
rect 4791 479 4794 480
rect 4826 510 4829 511
rect 5027 511 5065 512
rect 5027 510 5030 511
rect 4826 480 4874 510
rect 4982 480 5030 510
rect 4826 479 4829 480
rect 4791 478 4829 479
rect 5027 479 5030 480
rect 5062 510 5065 511
rect 5239 511 5277 512
rect 5239 510 5242 511
rect 5062 480 5109 510
rect 5195 480 5242 510
rect 5062 479 5065 480
rect 5027 478 5065 479
rect 5239 479 5242 480
rect 5274 510 5277 511
rect 5475 511 5513 512
rect 5475 510 5478 511
rect 5274 480 5322 510
rect 5430 480 5478 510
rect 5274 479 5277 480
rect 5239 478 5277 479
rect 5475 479 5478 480
rect 5510 510 5513 511
rect 5687 511 5725 512
rect 5687 510 5690 511
rect 5510 480 5557 510
rect 5643 480 5690 510
rect 5510 479 5513 480
rect 5475 478 5513 479
rect 5687 479 5690 480
rect 5722 510 5725 511
rect 5923 511 5961 512
rect 5923 510 5926 511
rect 5722 480 5770 510
rect 5878 480 5926 510
rect 5722 479 5725 480
rect 5687 478 5725 479
rect 5923 479 5926 480
rect 5958 510 5961 511
rect 6135 511 6173 512
rect 6135 510 6138 511
rect 5958 480 6005 510
rect 6091 480 6138 510
rect 5958 479 5961 480
rect 5923 478 5961 479
rect 6135 479 6138 480
rect 6170 510 6173 511
rect 6371 511 6409 512
rect 6371 510 6374 511
rect 6170 480 6218 510
rect 6326 480 6374 510
rect 6170 479 6173 480
rect 6135 478 6173 479
rect 6371 479 6374 480
rect 6406 510 6409 511
rect 6583 511 6621 512
rect 6583 510 6586 511
rect 6406 480 6453 510
rect 6539 480 6586 510
rect 6406 479 6409 480
rect 6371 478 6409 479
rect 6583 479 6586 480
rect 6618 510 6621 511
rect 6819 511 6857 512
rect 6819 510 6822 511
rect 6618 480 6666 510
rect 6774 480 6822 510
rect 6618 479 6621 480
rect 6583 478 6621 479
rect 6819 479 6822 480
rect 6854 510 6857 511
rect 7031 511 7069 512
rect 7031 510 7034 511
rect 6854 480 6901 510
rect 6987 480 7034 510
rect 6854 479 6857 480
rect 6819 478 6857 479
rect 7031 479 7034 480
rect 7066 510 7069 511
rect 7267 511 7305 512
rect 7267 510 7270 511
rect 7066 480 7114 510
rect 7222 480 7270 510
rect 7066 479 7069 480
rect 7031 478 7069 479
rect 7267 479 7270 480
rect 7302 510 7305 511
rect 7479 511 7517 512
rect 7479 510 7482 511
rect 7302 480 7349 510
rect 7435 480 7482 510
rect 7302 479 7305 480
rect 7267 478 7305 479
rect 7479 479 7482 480
rect 7514 510 7517 511
rect 7715 511 7753 512
rect 7715 510 7718 511
rect 7514 480 7562 510
rect 7670 480 7718 510
rect 7514 479 7517 480
rect 7479 478 7517 479
rect 7715 479 7718 480
rect 7750 510 7753 511
rect 7927 511 7965 512
rect 7927 510 7930 511
rect 7750 480 7797 510
rect 7883 480 7930 510
rect 7750 479 7753 480
rect 7715 478 7753 479
rect 7927 479 7930 480
rect 7962 510 7965 511
rect 8163 511 8201 512
rect 8163 510 8166 511
rect 7962 480 8010 510
rect 8118 480 8166 510
rect 7962 479 7965 480
rect 7927 478 7965 479
rect 8163 479 8166 480
rect 8198 510 8201 511
rect 8375 511 8413 512
rect 8375 510 8378 511
rect 8198 480 8245 510
rect 8331 480 8378 510
rect 8198 479 8201 480
rect 8163 478 8201 479
rect 8375 479 8378 480
rect 8410 510 8413 511
rect 8611 511 8649 512
rect 8611 510 8614 511
rect 8410 480 8458 510
rect 8566 480 8614 510
rect 8410 479 8413 480
rect 8375 478 8413 479
rect 8611 479 8614 480
rect 8646 510 8649 511
rect 8823 511 8861 512
rect 8823 510 8826 511
rect 8646 480 8693 510
rect 8779 480 8826 510
rect 8646 479 8649 480
rect 8611 478 8649 479
rect 8823 479 8826 480
rect 8858 510 8861 511
rect 8858 480 8906 510
rect 8858 479 8861 480
rect 8823 478 8861 479
rect 101 388 134 478
rect 314 388 347 478
rect 549 388 582 478
rect 762 388 795 478
rect 997 388 1030 478
rect 1210 388 1243 478
rect 1445 388 1478 478
rect 1658 388 1691 478
rect 1893 388 1926 478
rect 2106 388 2139 478
rect 2341 388 2374 478
rect 2554 388 2587 478
rect 2789 388 2822 478
rect 3002 388 3035 478
rect 3237 388 3270 478
rect 3450 388 3483 478
rect 3685 388 3718 478
rect 3898 388 3931 478
rect 4133 388 4166 478
rect 4346 388 4379 478
rect 4581 388 4614 478
rect 4794 388 4827 478
rect 5029 388 5062 478
rect 5242 388 5275 478
rect 5477 433 5510 478
rect 5690 433 5723 478
rect 5925 388 5958 478
rect 6138 388 6171 478
rect 6373 388 6406 478
rect 6586 388 6619 478
rect 6821 388 6854 478
rect 7034 388 7067 478
rect 7269 388 7302 478
rect 7482 388 7515 478
rect 7717 432 7750 478
rect 7930 388 7963 478
rect 8165 388 8198 478
rect 8378 388 8411 478
rect 8613 388 8646 478
rect 8826 388 8859 478
rect 99 387 137 388
rect 99 386 102 387
rect 54 356 102 386
rect 99 355 102 356
rect 134 386 137 387
rect 311 387 349 388
rect 311 386 314 387
rect 134 356 181 386
rect 267 356 314 386
rect 134 355 137 356
rect 99 354 137 355
rect 311 355 314 356
rect 346 386 349 387
rect 547 387 585 388
rect 547 386 550 387
rect 346 356 394 386
rect 502 356 550 386
rect 346 355 349 356
rect 311 354 349 355
rect 547 355 550 356
rect 582 386 585 387
rect 759 387 797 388
rect 759 386 762 387
rect 582 356 629 386
rect 715 356 762 386
rect 582 355 585 356
rect 547 354 585 355
rect 759 355 762 356
rect 794 386 797 387
rect 995 387 1033 388
rect 995 386 998 387
rect 794 356 842 386
rect 950 356 998 386
rect 794 355 797 356
rect 759 354 797 355
rect 995 355 998 356
rect 1030 386 1033 387
rect 1207 387 1245 388
rect 1207 386 1210 387
rect 1030 356 1077 386
rect 1163 356 1210 386
rect 1030 355 1033 356
rect 995 354 1033 355
rect 1207 355 1210 356
rect 1242 386 1245 387
rect 1443 387 1481 388
rect 1443 386 1446 387
rect 1242 356 1290 386
rect 1398 356 1446 386
rect 1242 355 1245 356
rect 1207 354 1245 355
rect 1443 355 1446 356
rect 1478 386 1481 387
rect 1655 387 1693 388
rect 1655 386 1658 387
rect 1478 356 1525 386
rect 1611 356 1658 386
rect 1478 355 1481 356
rect 1443 354 1481 355
rect 1655 355 1658 356
rect 1690 386 1693 387
rect 1891 387 1929 388
rect 1891 386 1894 387
rect 1690 356 1738 386
rect 1846 356 1894 386
rect 1690 355 1693 356
rect 1655 354 1693 355
rect 1891 355 1894 356
rect 1926 386 1929 387
rect 2103 387 2141 388
rect 2103 386 2106 387
rect 1926 356 1973 386
rect 2059 356 2106 386
rect 1926 355 1929 356
rect 1891 354 1929 355
rect 2103 355 2106 356
rect 2138 386 2141 387
rect 2339 387 2377 388
rect 2339 386 2342 387
rect 2138 356 2186 386
rect 2294 356 2342 386
rect 2138 355 2141 356
rect 2103 354 2141 355
rect 2339 355 2342 356
rect 2374 386 2377 387
rect 2551 387 2589 388
rect 2551 386 2554 387
rect 2374 356 2421 386
rect 2507 356 2554 386
rect 2374 355 2377 356
rect 2339 354 2377 355
rect 2551 355 2554 356
rect 2586 386 2589 387
rect 2787 387 2825 388
rect 2787 386 2790 387
rect 2586 356 2634 386
rect 2742 356 2790 386
rect 2586 355 2589 356
rect 2551 354 2589 355
rect 2787 355 2790 356
rect 2822 386 2825 387
rect 2999 387 3037 388
rect 2999 386 3002 387
rect 2822 356 2869 386
rect 2955 356 3002 386
rect 2822 355 2825 356
rect 2787 354 2825 355
rect 2999 355 3002 356
rect 3034 386 3037 387
rect 3235 387 3273 388
rect 3235 386 3238 387
rect 3034 356 3082 386
rect 3190 356 3238 386
rect 3034 355 3037 356
rect 2999 354 3037 355
rect 3235 355 3238 356
rect 3270 386 3273 387
rect 3447 387 3485 388
rect 3447 386 3450 387
rect 3270 356 3317 386
rect 3403 356 3450 386
rect 3270 355 3273 356
rect 3235 354 3273 355
rect 3447 355 3450 356
rect 3482 386 3485 387
rect 3683 387 3721 388
rect 3683 386 3686 387
rect 3482 356 3530 386
rect 3638 356 3686 386
rect 3482 355 3485 356
rect 3447 354 3485 355
rect 3683 355 3686 356
rect 3718 386 3721 387
rect 3895 387 3933 388
rect 3895 386 3898 387
rect 3718 356 3765 386
rect 3851 356 3898 386
rect 3718 355 3721 356
rect 3683 354 3721 355
rect 3895 355 3898 356
rect 3930 386 3933 387
rect 4131 387 4169 388
rect 4131 386 4134 387
rect 3930 356 3978 386
rect 4086 356 4134 386
rect 3930 355 3933 356
rect 3895 354 3933 355
rect 4131 355 4134 356
rect 4166 386 4169 387
rect 4343 387 4381 388
rect 4343 386 4346 387
rect 4166 356 4213 386
rect 4299 356 4346 386
rect 4166 355 4169 356
rect 4131 354 4169 355
rect 4343 355 4346 356
rect 4378 386 4381 387
rect 4579 387 4617 388
rect 4579 386 4582 387
rect 4378 356 4426 386
rect 4534 356 4582 386
rect 4378 355 4381 356
rect 4343 354 4381 355
rect 4579 355 4582 356
rect 4614 386 4617 387
rect 4791 387 4829 388
rect 4791 386 4794 387
rect 4614 356 4661 386
rect 4747 356 4794 386
rect 4614 355 4617 356
rect 4579 354 4617 355
rect 4791 355 4794 356
rect 4826 386 4829 387
rect 5027 387 5065 388
rect 5027 386 5030 387
rect 4826 356 4874 386
rect 4982 356 5030 386
rect 4826 355 4829 356
rect 4791 354 4829 355
rect 5027 355 5030 356
rect 5062 386 5065 387
rect 5239 387 5277 388
rect 5239 386 5242 387
rect 5062 356 5109 386
rect 5195 356 5242 386
rect 5062 355 5065 356
rect 5027 354 5065 355
rect 5239 355 5242 356
rect 5274 386 5277 387
rect 5475 387 5513 388
rect 5475 386 5478 387
rect 5274 356 5322 386
rect 5430 356 5478 386
rect 5274 355 5277 356
rect 5239 354 5277 355
rect 5475 355 5478 356
rect 5510 386 5513 387
rect 5687 387 5725 388
rect 5687 386 5690 387
rect 5510 356 5557 386
rect 5643 356 5690 386
rect 5510 355 5513 356
rect 5475 354 5513 355
rect 5687 355 5690 356
rect 5722 386 5725 387
rect 5923 387 5961 388
rect 5923 386 5926 387
rect 5722 356 5770 386
rect 5878 356 5926 386
rect 5722 355 5725 356
rect 5687 354 5725 355
rect 5923 355 5926 356
rect 5958 386 5961 387
rect 6135 387 6173 388
rect 6135 386 6138 387
rect 5958 356 6005 386
rect 6091 356 6138 386
rect 5958 355 5961 356
rect 5923 354 5961 355
rect 6135 355 6138 356
rect 6170 386 6173 387
rect 6371 387 6409 388
rect 6371 386 6374 387
rect 6170 356 6218 386
rect 6326 356 6374 386
rect 6170 355 6173 356
rect 6135 354 6173 355
rect 6371 355 6374 356
rect 6406 386 6409 387
rect 6583 387 6621 388
rect 6583 386 6586 387
rect 6406 356 6453 386
rect 6539 356 6586 386
rect 6406 355 6409 356
rect 6371 354 6409 355
rect 6583 355 6586 356
rect 6618 386 6621 387
rect 6819 387 6857 388
rect 6819 386 6822 387
rect 6618 356 6666 386
rect 6774 356 6822 386
rect 6618 355 6621 356
rect 6583 354 6621 355
rect 6819 355 6822 356
rect 6854 386 6857 387
rect 7031 387 7069 388
rect 7031 386 7034 387
rect 6854 356 6901 386
rect 6987 356 7034 386
rect 6854 355 6857 356
rect 6819 354 6857 355
rect 7031 355 7034 356
rect 7066 386 7069 387
rect 7267 387 7305 388
rect 7267 386 7270 387
rect 7066 356 7114 386
rect 7222 356 7270 386
rect 7066 355 7069 356
rect 7031 354 7069 355
rect 7267 355 7270 356
rect 7302 386 7305 387
rect 7479 387 7517 388
rect 7479 386 7482 387
rect 7302 356 7349 386
rect 7435 356 7482 386
rect 7302 355 7305 356
rect 7267 354 7305 355
rect 7479 355 7482 356
rect 7514 386 7517 387
rect 7715 387 7753 388
rect 7715 386 7718 387
rect 7514 356 7562 386
rect 7670 356 7718 386
rect 7514 355 7517 356
rect 7479 354 7517 355
rect 7715 355 7718 356
rect 7750 386 7753 387
rect 7927 387 7965 388
rect 7927 386 7930 387
rect 7750 356 7797 386
rect 7883 356 7930 386
rect 7750 355 7753 356
rect 7715 354 7753 355
rect 7927 355 7930 356
rect 7962 386 7965 387
rect 8163 387 8201 388
rect 8163 386 8166 387
rect 7962 356 8010 386
rect 8118 356 8166 386
rect 7962 355 7965 356
rect 7927 354 7965 355
rect 8163 355 8166 356
rect 8198 386 8201 387
rect 8375 387 8413 388
rect 8375 386 8378 387
rect 8198 356 8245 386
rect 8331 356 8378 386
rect 8198 355 8201 356
rect 8163 354 8201 355
rect 8375 355 8378 356
rect 8410 386 8413 387
rect 8611 387 8649 388
rect 8611 386 8614 387
rect 8410 356 8458 386
rect 8566 356 8614 386
rect 8410 355 8413 356
rect 8375 354 8413 355
rect 8611 355 8614 356
rect 8646 386 8649 387
rect 8823 387 8861 388
rect 8823 386 8826 387
rect 8646 356 8693 386
rect 8779 356 8826 386
rect 8646 355 8649 356
rect 8611 354 8649 355
rect 8823 355 8826 356
rect 8858 386 8861 387
rect 8858 356 8906 386
rect 8858 355 8861 356
rect 8823 354 8861 355
rect 101 264 134 354
rect 314 264 347 354
rect 549 264 582 354
rect 762 264 795 354
rect 997 264 1030 354
rect 1210 264 1243 354
rect 1445 264 1478 354
rect 1658 264 1691 354
rect 1893 264 1926 354
rect 2106 264 2139 354
rect 2341 264 2374 354
rect 2554 264 2587 354
rect 2789 264 2822 354
rect 3002 264 3035 354
rect 3237 309 3270 354
rect 3450 309 3483 354
rect 3685 264 3718 354
rect 3898 264 3931 354
rect 4133 264 4166 354
rect 4346 264 4379 354
rect 4581 264 4614 354
rect 4794 264 4827 354
rect 5029 264 5062 354
rect 5242 264 5275 354
rect 5477 264 5510 354
rect 5690 264 5723 354
rect 5925 264 5958 354
rect 6138 264 6171 354
rect 6373 264 6406 354
rect 6586 264 6619 354
rect 6821 264 6854 354
rect 7034 264 7067 354
rect 7269 264 7302 354
rect 7482 264 7515 354
rect 7717 264 7750 354
rect 7930 264 7963 354
rect 8165 264 8198 354
rect 8378 264 8411 354
rect 8613 264 8646 354
rect 8826 264 8859 354
rect 99 263 137 264
rect 99 262 102 263
rect 54 232 102 262
rect 99 231 102 232
rect 134 262 137 263
rect 311 263 349 264
rect 311 262 314 263
rect 134 232 181 262
rect 267 232 314 262
rect 134 231 137 232
rect 99 230 137 231
rect 311 231 314 232
rect 346 262 349 263
rect 547 263 585 264
rect 547 262 550 263
rect 346 232 394 262
rect 502 232 550 262
rect 346 231 349 232
rect 311 230 349 231
rect 547 231 550 232
rect 582 262 585 263
rect 759 263 797 264
rect 759 262 762 263
rect 582 232 629 262
rect 715 232 762 262
rect 582 231 585 232
rect 547 230 585 231
rect 759 231 762 232
rect 794 262 797 263
rect 995 263 1033 264
rect 995 262 998 263
rect 794 232 842 262
rect 950 232 998 262
rect 794 231 797 232
rect 759 230 797 231
rect 995 231 998 232
rect 1030 262 1033 263
rect 1207 263 1245 264
rect 1207 262 1210 263
rect 1030 232 1077 262
rect 1163 232 1210 262
rect 1030 231 1033 232
rect 995 230 1033 231
rect 1207 231 1210 232
rect 1242 262 1245 263
rect 1443 263 1481 264
rect 1443 262 1446 263
rect 1242 232 1290 262
rect 1398 232 1446 262
rect 1242 231 1245 232
rect 1207 230 1245 231
rect 1443 231 1446 232
rect 1478 262 1481 263
rect 1655 263 1693 264
rect 1655 262 1658 263
rect 1478 232 1525 262
rect 1611 232 1658 262
rect 1478 231 1481 232
rect 1443 230 1481 231
rect 1655 231 1658 232
rect 1690 262 1693 263
rect 1891 263 1929 264
rect 1891 262 1894 263
rect 1690 232 1738 262
rect 1846 232 1894 262
rect 1690 231 1693 232
rect 1655 230 1693 231
rect 1891 231 1894 232
rect 1926 262 1929 263
rect 2103 263 2141 264
rect 2103 262 2106 263
rect 1926 232 1973 262
rect 2059 232 2106 262
rect 1926 231 1929 232
rect 1891 230 1929 231
rect 2103 231 2106 232
rect 2138 262 2141 263
rect 2339 263 2377 264
rect 2339 262 2342 263
rect 2138 232 2186 262
rect 2294 232 2342 262
rect 2138 231 2141 232
rect 2103 230 2141 231
rect 2339 231 2342 232
rect 2374 262 2377 263
rect 2551 263 2589 264
rect 2551 262 2554 263
rect 2374 232 2421 262
rect 2507 232 2554 262
rect 2374 231 2377 232
rect 2339 230 2377 231
rect 2551 231 2554 232
rect 2586 262 2589 263
rect 2787 263 2825 264
rect 2787 262 2790 263
rect 2586 232 2634 262
rect 2742 232 2790 262
rect 2586 231 2589 232
rect 2551 230 2589 231
rect 2787 231 2790 232
rect 2822 262 2825 263
rect 2999 263 3037 264
rect 2999 262 3002 263
rect 2822 232 2869 262
rect 2955 232 3002 262
rect 2822 231 2825 232
rect 2787 230 2825 231
rect 2999 231 3002 232
rect 3034 262 3037 263
rect 3235 263 3273 264
rect 3235 262 3238 263
rect 3034 232 3082 262
rect 3190 232 3238 262
rect 3034 231 3037 232
rect 2999 230 3037 231
rect 3235 231 3238 232
rect 3270 262 3273 263
rect 3447 263 3485 264
rect 3447 262 3450 263
rect 3270 232 3317 262
rect 3403 232 3450 262
rect 3270 231 3273 232
rect 3235 230 3273 231
rect 3447 231 3450 232
rect 3482 262 3485 263
rect 3683 263 3721 264
rect 3683 262 3686 263
rect 3482 232 3530 262
rect 3638 232 3686 262
rect 3482 231 3485 232
rect 3447 230 3485 231
rect 3683 231 3686 232
rect 3718 262 3721 263
rect 3895 263 3933 264
rect 3895 262 3898 263
rect 3718 232 3765 262
rect 3851 232 3898 262
rect 3718 231 3721 232
rect 3683 230 3721 231
rect 3895 231 3898 232
rect 3930 262 3933 263
rect 4131 263 4169 264
rect 4131 262 4134 263
rect 3930 232 3978 262
rect 4086 232 4134 262
rect 3930 231 3933 232
rect 3895 230 3933 231
rect 4131 231 4134 232
rect 4166 262 4169 263
rect 4343 263 4381 264
rect 4343 262 4346 263
rect 4166 232 4213 262
rect 4299 232 4346 262
rect 4166 231 4169 232
rect 4131 230 4169 231
rect 4343 231 4346 232
rect 4378 262 4381 263
rect 4579 263 4617 264
rect 4579 262 4582 263
rect 4378 232 4426 262
rect 4534 232 4582 262
rect 4378 231 4381 232
rect 4343 230 4381 231
rect 4579 231 4582 232
rect 4614 262 4617 263
rect 4791 263 4829 264
rect 4791 262 4794 263
rect 4614 232 4661 262
rect 4747 232 4794 262
rect 4614 231 4617 232
rect 4579 230 4617 231
rect 4791 231 4794 232
rect 4826 262 4829 263
rect 5027 263 5065 264
rect 5027 262 5030 263
rect 4826 232 4874 262
rect 4982 232 5030 262
rect 4826 231 4829 232
rect 4791 230 4829 231
rect 5027 231 5030 232
rect 5062 262 5065 263
rect 5239 263 5277 264
rect 5239 262 5242 263
rect 5062 232 5109 262
rect 5195 232 5242 262
rect 5062 231 5065 232
rect 5027 230 5065 231
rect 5239 231 5242 232
rect 5274 262 5277 263
rect 5475 263 5513 264
rect 5475 262 5478 263
rect 5274 232 5322 262
rect 5430 232 5478 262
rect 5274 231 5277 232
rect 5239 230 5277 231
rect 5475 231 5478 232
rect 5510 262 5513 263
rect 5687 263 5725 264
rect 5687 262 5690 263
rect 5510 232 5557 262
rect 5643 232 5690 262
rect 5510 231 5513 232
rect 5475 230 5513 231
rect 5687 231 5690 232
rect 5722 262 5725 263
rect 5923 263 5961 264
rect 5923 262 5926 263
rect 5722 232 5770 262
rect 5878 232 5926 262
rect 5722 231 5725 232
rect 5687 230 5725 231
rect 5923 231 5926 232
rect 5958 262 5961 263
rect 6135 263 6173 264
rect 6135 262 6138 263
rect 5958 232 6005 262
rect 6091 232 6138 262
rect 5958 231 5961 232
rect 5923 230 5961 231
rect 6135 231 6138 232
rect 6170 262 6173 263
rect 6371 263 6409 264
rect 6371 262 6374 263
rect 6170 232 6218 262
rect 6326 232 6374 262
rect 6170 231 6173 232
rect 6135 230 6173 231
rect 6371 231 6374 232
rect 6406 262 6409 263
rect 6583 263 6621 264
rect 6583 262 6586 263
rect 6406 232 6453 262
rect 6539 232 6586 262
rect 6406 231 6409 232
rect 6371 230 6409 231
rect 6583 231 6586 232
rect 6618 262 6621 263
rect 6819 263 6857 264
rect 6819 262 6822 263
rect 6618 232 6666 262
rect 6774 232 6822 262
rect 6618 231 6621 232
rect 6583 230 6621 231
rect 6819 231 6822 232
rect 6854 262 6857 263
rect 7031 263 7069 264
rect 7031 262 7034 263
rect 6854 232 6901 262
rect 6987 232 7034 262
rect 6854 231 6857 232
rect 6819 230 6857 231
rect 7031 231 7034 232
rect 7066 262 7069 263
rect 7267 263 7305 264
rect 7267 262 7270 263
rect 7066 232 7114 262
rect 7222 232 7270 262
rect 7066 231 7069 232
rect 7031 230 7069 231
rect 7267 231 7270 232
rect 7302 262 7305 263
rect 7479 263 7517 264
rect 7479 262 7482 263
rect 7302 232 7349 262
rect 7435 232 7482 262
rect 7302 231 7305 232
rect 7267 230 7305 231
rect 7479 231 7482 232
rect 7514 262 7517 263
rect 7715 263 7753 264
rect 7715 262 7718 263
rect 7514 232 7562 262
rect 7670 232 7718 262
rect 7514 231 7517 232
rect 7479 230 7517 231
rect 7715 231 7718 232
rect 7750 262 7753 263
rect 7927 263 7965 264
rect 7927 262 7930 263
rect 7750 232 7797 262
rect 7883 232 7930 262
rect 7750 231 7753 232
rect 7715 230 7753 231
rect 7927 231 7930 232
rect 7962 262 7965 263
rect 8163 263 8201 264
rect 8163 262 8166 263
rect 7962 232 8010 262
rect 8118 232 8166 262
rect 7962 231 7965 232
rect 7927 230 7965 231
rect 8163 231 8166 232
rect 8198 262 8201 263
rect 8375 263 8413 264
rect 8375 262 8378 263
rect 8198 232 8245 262
rect 8331 232 8378 262
rect 8198 231 8201 232
rect 8163 230 8201 231
rect 8375 231 8378 232
rect 8410 262 8413 263
rect 8611 263 8649 264
rect 8611 262 8614 263
rect 8410 232 8458 262
rect 8566 232 8614 262
rect 8410 231 8413 232
rect 8375 230 8413 231
rect 8611 231 8614 232
rect 8646 262 8649 263
rect 8823 263 8861 264
rect 8823 262 8826 263
rect 8646 232 8693 262
rect 8779 232 8826 262
rect 8646 231 8649 232
rect 8611 230 8649 231
rect 8823 231 8826 232
rect 8858 262 8861 263
rect 8858 232 8906 262
rect 8858 231 8861 232
rect 8823 230 8861 231
rect 101 140 134 230
rect 314 140 347 230
rect 549 140 582 230
rect 762 140 795 230
rect 997 140 1030 230
rect 1210 140 1243 230
rect 1445 140 1478 230
rect 1658 140 1691 230
rect 1893 140 1926 230
rect 2106 140 2139 230
rect 2341 140 2374 230
rect 2554 140 2587 230
rect 2789 140 2822 230
rect 3002 140 3035 230
rect 3237 140 3270 230
rect 3450 140 3483 230
rect 3685 140 3718 230
rect 3898 140 3931 230
rect 4133 140 4166 230
rect 4346 140 4379 230
rect 4581 140 4614 230
rect 4794 140 4827 230
rect 5029 140 5062 230
rect 5242 140 5275 230
rect 5477 140 5510 230
rect 5690 140 5723 230
rect 5925 140 5958 230
rect 6138 140 6171 230
rect 6373 140 6406 230
rect 6586 140 6619 230
rect 6821 140 6854 230
rect 7034 140 7067 230
rect 7269 140 7302 230
rect 7482 140 7515 230
rect 7717 140 7750 230
rect 7930 140 7963 230
rect 8165 140 8198 230
rect 8378 140 8411 230
rect 8613 140 8646 230
rect 8826 140 8859 230
rect 99 139 137 140
rect 99 138 102 139
rect 54 108 102 138
rect 99 107 102 108
rect 134 138 137 139
rect 311 139 349 140
rect 311 138 314 139
rect 134 108 181 138
rect 267 108 314 138
rect 134 107 137 108
rect 99 106 137 107
rect 311 107 314 108
rect 346 138 349 139
rect 547 139 585 140
rect 547 138 550 139
rect 346 108 394 138
rect 502 108 550 138
rect 346 107 349 108
rect 311 106 349 107
rect 547 107 550 108
rect 582 138 585 139
rect 759 139 797 140
rect 759 138 762 139
rect 582 108 629 138
rect 715 108 762 138
rect 582 107 585 108
rect 547 106 585 107
rect 759 107 762 108
rect 794 138 797 139
rect 995 139 1033 140
rect 995 138 998 139
rect 794 108 842 138
rect 950 108 998 138
rect 794 107 797 108
rect 759 106 797 107
rect 995 107 998 108
rect 1030 138 1033 139
rect 1207 139 1245 140
rect 1207 138 1210 139
rect 1030 108 1077 138
rect 1163 108 1210 138
rect 1030 107 1033 108
rect 995 106 1033 107
rect 1207 107 1210 108
rect 1242 138 1245 139
rect 1443 139 1481 140
rect 1443 138 1446 139
rect 1242 108 1290 138
rect 1398 108 1446 138
rect 1242 107 1245 108
rect 1207 106 1245 107
rect 1443 107 1446 108
rect 1478 138 1481 139
rect 1655 139 1693 140
rect 1655 138 1658 139
rect 1478 108 1525 138
rect 1611 108 1658 138
rect 1478 107 1481 108
rect 1443 106 1481 107
rect 1655 107 1658 108
rect 1690 138 1693 139
rect 1891 139 1929 140
rect 1891 138 1894 139
rect 1690 108 1738 138
rect 1846 108 1894 138
rect 1690 107 1693 108
rect 1655 106 1693 107
rect 1891 107 1894 108
rect 1926 138 1929 139
rect 2103 139 2141 140
rect 2103 138 2106 139
rect 1926 108 1973 138
rect 2059 108 2106 138
rect 1926 107 1929 108
rect 1891 106 1929 107
rect 2103 107 2106 108
rect 2138 138 2141 139
rect 2339 139 2377 140
rect 2339 138 2342 139
rect 2138 108 2186 138
rect 2294 108 2342 138
rect 2138 107 2141 108
rect 2103 106 2141 107
rect 2339 107 2342 108
rect 2374 138 2377 139
rect 2551 139 2589 140
rect 2551 138 2554 139
rect 2374 108 2421 138
rect 2507 108 2554 138
rect 2374 107 2377 108
rect 2339 106 2377 107
rect 2551 107 2554 108
rect 2586 138 2589 139
rect 2787 139 2825 140
rect 2787 138 2790 139
rect 2586 108 2634 138
rect 2742 108 2790 138
rect 2586 107 2589 108
rect 2551 106 2589 107
rect 2787 107 2790 108
rect 2822 138 2825 139
rect 2999 139 3037 140
rect 2999 138 3002 139
rect 2822 108 2869 138
rect 2955 108 3002 138
rect 2822 107 2825 108
rect 2787 106 2825 107
rect 2999 107 3002 108
rect 3034 138 3037 139
rect 3235 139 3273 140
rect 3235 138 3238 139
rect 3034 108 3082 138
rect 3190 108 3238 138
rect 3034 107 3037 108
rect 2999 106 3037 107
rect 3235 107 3238 108
rect 3270 138 3273 139
rect 3447 139 3485 140
rect 3447 138 3450 139
rect 3270 108 3317 138
rect 3403 108 3450 138
rect 3270 107 3273 108
rect 3235 106 3273 107
rect 3447 107 3450 108
rect 3482 138 3485 139
rect 3683 139 3721 140
rect 3683 138 3686 139
rect 3482 108 3530 138
rect 3638 108 3686 138
rect 3482 107 3485 108
rect 3447 106 3485 107
rect 3683 107 3686 108
rect 3718 138 3721 139
rect 3895 139 3933 140
rect 3895 138 3898 139
rect 3718 108 3765 138
rect 3851 108 3898 138
rect 3718 107 3721 108
rect 3683 106 3721 107
rect 3895 107 3898 108
rect 3930 138 3933 139
rect 4131 139 4169 140
rect 4131 138 4134 139
rect 3930 108 3978 138
rect 4086 108 4134 138
rect 3930 107 3933 108
rect 3895 106 3933 107
rect 4131 107 4134 108
rect 4166 138 4169 139
rect 4343 139 4381 140
rect 4343 138 4346 139
rect 4166 108 4213 138
rect 4299 108 4346 138
rect 4166 107 4169 108
rect 4131 106 4169 107
rect 4343 107 4346 108
rect 4378 138 4381 139
rect 4579 139 4617 140
rect 4579 138 4582 139
rect 4378 108 4426 138
rect 4534 108 4582 138
rect 4378 107 4381 108
rect 4343 106 4381 107
rect 4579 107 4582 108
rect 4614 138 4617 139
rect 4791 139 4829 140
rect 4791 138 4794 139
rect 4614 108 4661 138
rect 4747 108 4794 138
rect 4614 107 4617 108
rect 4579 106 4617 107
rect 4791 107 4794 108
rect 4826 138 4829 139
rect 5027 139 5065 140
rect 5027 138 5030 139
rect 4826 108 4874 138
rect 4982 108 5030 138
rect 4826 107 4829 108
rect 4791 106 4829 107
rect 5027 107 5030 108
rect 5062 138 5065 139
rect 5239 139 5277 140
rect 5239 138 5242 139
rect 5062 108 5109 138
rect 5195 108 5242 138
rect 5062 107 5065 108
rect 5027 106 5065 107
rect 5239 107 5242 108
rect 5274 138 5277 139
rect 5475 139 5513 140
rect 5475 138 5478 139
rect 5274 108 5322 138
rect 5430 108 5478 138
rect 5274 107 5277 108
rect 5239 106 5277 107
rect 5475 107 5478 108
rect 5510 138 5513 139
rect 5687 139 5725 140
rect 5687 138 5690 139
rect 5510 108 5557 138
rect 5643 108 5690 138
rect 5510 107 5513 108
rect 5475 106 5513 107
rect 5687 107 5690 108
rect 5722 138 5725 139
rect 5923 139 5961 140
rect 5923 138 5926 139
rect 5722 108 5770 138
rect 5878 108 5926 138
rect 5722 107 5725 108
rect 5687 106 5725 107
rect 5923 107 5926 108
rect 5958 138 5961 139
rect 6135 139 6173 140
rect 6135 138 6138 139
rect 5958 108 6005 138
rect 6091 108 6138 138
rect 5958 107 5961 108
rect 5923 106 5961 107
rect 6135 107 6138 108
rect 6170 138 6173 139
rect 6371 139 6409 140
rect 6371 138 6374 139
rect 6170 108 6218 138
rect 6326 108 6374 138
rect 6170 107 6173 108
rect 6135 106 6173 107
rect 6371 107 6374 108
rect 6406 138 6409 139
rect 6583 139 6621 140
rect 6583 138 6586 139
rect 6406 108 6453 138
rect 6539 108 6586 138
rect 6406 107 6409 108
rect 6371 106 6409 107
rect 6583 107 6586 108
rect 6618 138 6621 139
rect 6819 139 6857 140
rect 6819 138 6822 139
rect 6618 108 6666 138
rect 6774 108 6822 138
rect 6618 107 6621 108
rect 6583 106 6621 107
rect 6819 107 6822 108
rect 6854 138 6857 139
rect 7031 139 7069 140
rect 7031 138 7034 139
rect 6854 108 6901 138
rect 6987 108 7034 138
rect 6854 107 6857 108
rect 6819 106 6857 107
rect 7031 107 7034 108
rect 7066 138 7069 139
rect 7267 139 7305 140
rect 7267 138 7270 139
rect 7066 108 7114 138
rect 7222 108 7270 138
rect 7066 107 7069 108
rect 7031 106 7069 107
rect 7267 107 7270 108
rect 7302 138 7305 139
rect 7479 139 7517 140
rect 7479 138 7482 139
rect 7302 108 7349 138
rect 7435 108 7482 138
rect 7302 107 7305 108
rect 7267 106 7305 107
rect 7479 107 7482 108
rect 7514 138 7517 139
rect 7715 139 7753 140
rect 7715 138 7718 139
rect 7514 108 7562 138
rect 7670 108 7718 138
rect 7514 107 7517 108
rect 7479 106 7517 107
rect 7715 107 7718 108
rect 7750 138 7753 139
rect 7927 139 7965 140
rect 7927 138 7930 139
rect 7750 108 7797 138
rect 7883 108 7930 138
rect 7750 107 7753 108
rect 7715 106 7753 107
rect 7927 107 7930 108
rect 7962 138 7965 139
rect 8163 139 8201 140
rect 8163 138 8166 139
rect 7962 108 8010 138
rect 8118 108 8166 138
rect 7962 107 7965 108
rect 7927 106 7965 107
rect 8163 107 8166 108
rect 8198 138 8201 139
rect 8375 139 8413 140
rect 8375 138 8378 139
rect 8198 108 8245 138
rect 8331 108 8378 138
rect 8198 107 8201 108
rect 8163 106 8201 107
rect 8375 107 8378 108
rect 8410 138 8413 139
rect 8611 139 8649 140
rect 8611 138 8614 139
rect 8410 108 8458 138
rect 8566 108 8614 138
rect 8410 107 8413 108
rect 8375 106 8413 107
rect 8611 107 8614 108
rect 8646 138 8649 139
rect 8823 139 8861 140
rect 8823 138 8826 139
rect 8646 108 8693 138
rect 8779 108 8826 138
rect 8646 107 8649 108
rect 8611 106 8649 107
rect 8823 107 8826 108
rect 8858 138 8861 139
rect 8858 108 8906 138
rect 8858 107 8861 108
rect 8823 106 8861 107
rect 101 16 134 106
rect 314 16 347 106
rect 549 16 582 106
rect 762 16 795 106
rect 997 16 1030 106
rect 1210 16 1243 106
rect 1445 16 1478 106
rect 1658 16 1691 106
rect 1893 16 1926 106
rect 2106 16 2139 106
rect 2341 16 2374 106
rect 2554 16 2587 106
rect 2789 16 2822 106
rect 3002 16 3035 106
rect 3237 61 3270 106
rect 3450 61 3483 106
rect 3685 16 3718 106
rect 3898 16 3931 106
rect 4133 16 4166 106
rect 4346 16 4379 106
rect 4581 16 4614 106
rect 4794 16 4827 106
rect 5029 16 5062 106
rect 5242 16 5275 106
rect 5477 62 5510 106
rect 5690 62 5723 106
rect 5925 16 5958 106
rect 6138 16 6171 106
rect 6373 16 6406 106
rect 6586 16 6619 106
rect 6821 16 6854 106
rect 7034 16 7067 106
rect 7269 16 7302 106
rect 7482 16 7515 106
rect 7717 61 7750 106
rect 7930 61 7963 106
rect 8165 16 8198 106
rect 8378 16 8411 106
rect 8613 16 8646 106
rect 8826 16 8859 106
rect 0 -16 8960 16
<< labels >>
rlabel metal2 16 27 16 59 7 dummy_bot
rlabel metal4 0 -16 0 16 7 dummy-top
rlabel metal4 549 603 549 635 7 top_8
rlabel metal3 483 665 483 695 7 bot_8
rlabel metal4 2789 603 2789 633 7 top_4
rlabel metal3 2723 665 2723 695 7 bot_4
rlabel metal4 5029 603 5029 633 7 top_2
rlabel metal3 4963 665 4963 695 7 bot_2
rlabel metal4 7269 603 7269 633 7 top_1
rlabel metal3 7203 665 7203 695 7 bot_1
<< end >>
