* NGSPICE file created from adc_clkgen_with_edgedetect.ext - technology: sky130A

.subckt sky130_fd_sc_hd__inv_2 A Y VPWR VGND VNB VPB
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=5.2e+11p ps=5.04e+06u w=1e+06u l=150000u
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=3.38e+11p pd=3.64e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__decap_4 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=4.524e+11p pd=4.52e+06u as=0p ps=0u w=870000u l=1.05e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=2.86e+11p pd=3.24e+06u as=0p ps=0u w=550000u l=1.05e+06u
.ends

.subckt sky130_fd_sc_hd__mux2_1 VGND VPWR S A1 A0 X VNB VPB
X0 VPWR a_505_21# a_535_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=4.553e+11p pd=4.29e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X1 a_505_21# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X2 a_218_374# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X3 VGND a_505_21# a_439_47# VNB sky130_fd_pr__nfet_01v8 ad=5.155e+11p pd=4.31e+06u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4 a_76_199# A0 a_218_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X5 a_505_21# S VGND VNB sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X6 a_439_47# A0 a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X7 a_535_374# A1 a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_76_199# A1 a_218_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X9 a_218_47# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VPWR VPB VNB
D0 VNB DIODE sky130_fd_pr__diode_pw2nd_05v5 pj=2.64e+06u area=4.347e+11p
.ends

.subckt sky130_fd_sc_hd__decap_6 VPWR VGND VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=4.524e+11p pd=4.52e+06u as=0p ps=0u w=870000u l=1.97e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=2.86e+11p pd=3.24e+06u as=0p ps=0u w=550000u l=1.97e+06u
.ends

.subckt sky130_fd_sc_hd__or2_1 A X B VGND VPWR VNB VPB
X0 VGND A a_68_297# VNB sky130_fd_pr__nfet_01v8 ad=3.097e+11p pd=3.33e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X1 a_68_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 X a_68_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X3 VPWR A a_150_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=2.915e+11p pd=2.67e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X4 X a_68_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=3.4e+11p pd=2.68e+06u as=0p ps=0u w=1e+06u l=150000u
X5 a_150_297# B a_68_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__decap_3 VPWR VGND VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=4.524e+11p pd=4.52e+06u as=0p ps=0u w=870000u l=590000u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=2.86e+11p pd=3.24e+06u as=0p ps=0u w=550000u l=590000u
.ends

.subckt sky130_mm_sc_hd_dlyPoly5ns VPWR in out VGND VNB VPB
X0 a_851_95# in VGND VNB sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=1.0453e+12p ps=9.52e+06u w=420000u l=3.83e+06u
X1 a_1724_71# a_851_95# VGND VNB sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X2 VPWR out a_1724_71# VNB sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3 VGND out a_1783_329# VPB sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u
X4 a_1783_329# out VGND VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5 a_1724_71# out VPWR VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VGND a_851_95# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X7 a_1783_329# a_851_95# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.72e+11p ps=4.38e+06u w=800000u l=150000u
X8 out a_851_95# a_1783_329# VPB sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X9 a_851_95# in VPWR VPB sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X10 out a_851_95# a_1724_71# VNB sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
C0 VGND a_851_95# 1.77fF
C1 VGND VNB 1.45fF
C2 VPWR VNB 1.20fF
C3 in VNB 1.50fF
C4 VPB VNB 2.04fF
.ends

.subckt sky130_fd_sc_hd__and2_1 VPWR VGND X B A VNB VPB
X0 VPWR B a_59_75# VPB sky130_fd_pr__pfet_01v8_hvt ad=4.507e+11p pd=4.18e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X1 X a_59_75# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=4.75e+11p pd=2.95e+06u as=0p ps=0u w=1e+06u l=150000u
X2 VGND B a_145_75# VNB sky130_fd_pr__nfet_01v8 ad=2.236e+11p pd=2.08e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X3 a_59_75# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 X a_59_75# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X5 a_145_75# A a_59_75# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__decap_8 VPWR VGND VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=4.524e+11p pd=4.52e+06u as=0p ps=0u w=870000u l=2.89e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=2.86e+11p pd=3.24e+06u as=0p ps=0u w=550000u l=2.89e+06u
C0 VGND VPWR 1.26fF
C1 VPWR VNB 1.11fF
.ends

.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=4.524e+11p pd=4.52e+06u as=0p ps=0u w=870000u l=4.73e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=2.86e+11p pd=3.24e+06u as=0p ps=0u w=550000u l=4.73e+06u
C0 VGND VPWR 1.27fF
C1 VPWR VNB 1.62fF
C2 VGND VNB 1.45fF
C3 VPB VNB 1.14fF
.ends

.subckt sky130_fd_sc_hd__nor2b_1 B_N Y A VGND VPWR VNB VPB
X0 Y a_74_47# a_265_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X1 VPWR B_N a_74_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=3.146e+11p pd=2.78e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X2 a_265_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=3.695e+11p ps=3.79e+06u w=650000u l=150000u
X4 VGND B_N a_74_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X5 VGND a_74_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__and2b_1 X A_N B VGND VPWR VNB VPB
X0 VPWR B a_207_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=5.986e+11p pd=5e+06u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X1 X a_207_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X2 a_297_47# a_27_413# a_207_413# VNB sky130_fd_pr__nfet_01v8 ad=1.008e+11p pd=1.32e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X3 X a_207_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=3.118e+11p ps=3.34e+06u w=650000u l=150000u
X4 a_207_413# a_27_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VPWR A_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X6 VGND B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_27_413# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__buf_1 VGND VPWR X A VNB VPB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=2.291e+11p pd=2.16e+06u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X1 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=1.508e+11p ps=1.62e+06u w=520000u l=150000u
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X3 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
.ends

.subckt sky130_fd_sc_hd__buf_4 VPWR VGND X A VNB VPB
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=8e+11p pd=7.6e+06u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=5.2e+11p ps=5.5e+06u w=650000u l=150000u
X5 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X9 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
.ends

.subckt adc_clkgen_with_edgedetect VGND VPWR clk_comp_out clk_dig_out dlycontrol1_in[0]
+ dlycontrol1_in[1] dlycontrol1_in[2] dlycontrol1_in[3] dlycontrol1_in[4] dlycontrol2_in[0]
+ dlycontrol2_in[1] dlycontrol2_in[2] dlycontrol2_in[3] dlycontrol2_in[4] dlycontrol3_in[0]
+ dlycontrol3_in[1] dlycontrol3_in[2] dlycontrol3_in[3] dlycontrol3_in[4] dlycontrol4_in[0]
+ dlycontrol4_in[1] dlycontrol4_in[2] dlycontrol4_in[3] dlycontrol4_in[4] dlycontrol4_in[5]
+ ena_in enable_dlycontrol_in ndecision_finish_in nsample_n_in nsample_n_out nsample_p_in
+ nsample_p_out sample_n_in sample_n_out sample_p_in sample_p_out start_conv_in
Xclkgen.delay_155ns_2.genblk1\[0\].control_invert dlycontrol2_in[0] clkgen.delay_155ns_2.genblk1\[0\].bypass_enable/B
+ VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_12_32 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_2.genblk1\[0\].dly_binary.out_mux VGND VPWR clkgen.delay_155ns_2.genblk1\[0\].bypass_enable/X
+ outbuf_1/A clkgen.delay_155ns_2.genblk1\[0\].dly_binary.out_mux/A0 clkgen.delay_155ns_2.genblk1\[0\].dly_binary.out_mux/X
+ VGND VPWR sky130_fd_sc_hd__mux2_1
Xclkgen.delay_155ns_2.genblk1\[2\].dly_binary.out_mux VGND VPWR clkgen.delay_155ns_2.genblk1\[2\].bypass_enable/X
+ clkgen.delay_155ns_2.genblk1\[1\].dly_binary.out_mux/X clkgen.delay_155ns_2.genblk1\[2\].dly_binary.out_mux/A0
+ clkgen.delay_155ns_2.genblk1\[2\].dly_binary.out_mux/X VGND VPWR sky130_fd_sc_hd__mux2_1
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.out_mux VGND VPWR clkgen.delay_155ns_2.genblk1\[4\].bypass_enable/X
+ clkgen.delay_155ns_2.genblk1\[3\].dly_binary.out_mux/X clkgen.delay_155ns_2.genblk1\[4\].dly_binary.out_mux/A0
+ clkgen.nor1/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_9_11 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.delay_155ns_1.genblk1\[2\].control_invert_A dlycontrol1_in[2] VGND
+ VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_2_121 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xedgedetect.or1 edgedetect.or1/A clkgen.nor1/B_N inbuf_1/X VGND VPWR VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_20_32 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xclkgen.delay_155ns_3.genblk1\[0\].dly_binary.genblk1\[0\].delay_unit VPWR clkgen.delay_155ns_3.genblk1\[0\].dly_binary.and_bypass_switch/X
+ clkgen.delay_155ns_3.genblk1\[0\].dly_binary.out_mux/A0 VGND VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[1\].bypass_enable VPWR VGND edgedetect.dly_315ns_1.genblk1\[1\].bypass_enable/X
+ edgedetect.dly_315ns_1.genblk1\[1\].bypass_enable/B edgedetect.dly_315ns_1.enablebuffer/X
+ VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_3_271 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_315 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_164 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.delay_155ns_2.genblk1\[1\].control_invert_A dlycontrol2_in[1] VGND
+ VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit VPWR clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit/in
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_10_307 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.delay_155ns_2.genblk1\[1\].dly_binary.and_bypass_switch_A_N clkgen.delay_155ns_2.genblk1\[1\].bypass_enable/X
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_5_311 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
Xclkgen.delay_155ns_1.genblk1\[2\].bypass_enable VPWR VGND clkgen.delay_155ns_1.genblk1\[2\].bypass_enable/X
+ clkgen.delay_155ns_1.genblk1\[2\].bypass_enable/B clkgen.delay_155ns_1.enablebuffer/X
+ VGND VPWR sky130_fd_sc_hd__and2_1
Xclkgen.delay_155ns_2.genblk1\[3\].bypass_enable VPWR VGND clkgen.delay_155ns_2.genblk1\[3\].bypass_enable/X
+ clkgen.delay_155ns_2.genblk1\[3\].bypass_enable/B clkgen.delay_155ns_2.enablebuffer/X
+ VGND VPWR sky130_fd_sc_hd__and2_1
Xclkgen.delay_155ns_3.genblk1\[4\].bypass_enable VPWR VGND clkgen.delay_155ns_3.genblk1\[4\].bypass_enable/X
+ clkgen.delay_155ns_3.genblk1\[4\].bypass_enable/B clkgen.delay_155ns_3.enablebuffer/X
+ VGND VPWR sky130_fd_sc_hd__and2_1
XANTENNA_clkgen.delay_155ns_3.genblk1\[0\].control_invert_A dlycontrol3_in[0] VGND
+ VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[3\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[3\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[4\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_clkgen.delay_155ns_3.genblk1\[4\].bypass_enable_A clkgen.delay_155ns_3.enablebuffer/X
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_20_276 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_32 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_276 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_214 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit VPWR clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit/in
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[2\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[1\].control_invert dlycontrol4_in[1] edgedetect.dly_315ns_1.genblk1\[1\].bypass_enable/B
+ VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_16_121 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[8\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[8\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[9\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_outbuf_6_A nsample_n_in VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_7_9 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.delay_155ns_1.genblk1\[4\].dly_binary.and_bypass_switch_A_N clkgen.delay_155ns_1.genblk1\[4\].bypass_enable/X
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_2_304 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit VPWR clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit/in
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit VPWR clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit/in
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_14_274 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_3 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xedgedetect.nor1 inbuf_2/X edgedetect.or1/A edgedetect.nor1/A VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__nor2b_1
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[0\].delay_unit VPWR clkgen.delay_155ns_2.genblk1\[4\].dly_binary.and_bypass_switch/X
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_11_288 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[1\].control_invert dlycontrol3_in[1] clkgen.delay_155ns_3.genblk1\[1\].bypass_enable/B
+ VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_232 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_13_125 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit VPWR clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit/in
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_2_316 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit VPWR clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit/in
+ clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_5_154 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[10\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[9\].delay_unit/out
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[11\].delay_unit/in VGND
+ VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[10\].delay_unit VPWR clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit/out
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_edgedetect.dly_315ns_1.genblk1\[5\].bypass_enable_A edgedetect.dly_315ns_1.enablebuffer/X
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_19_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit/in VGND
+ VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit VPWR clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit/in
+ clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_0_244 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_3 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit VPWR clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit/in
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.and_bypass_switch_A_N edgedetect.dly_315ns_1.genblk1\[3\].bypass_enable/X
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[0\].delay_unit VPWR clkgen.delay_155ns_2.genblk1\[3\].dly_binary.and_bypass_switch/X
+ clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[15\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[15\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[16\].delay_unit/in VGND
+ VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit VPWR clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit/in
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.out_mux/A0 VGND VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.nor1 clkgen.nor1/B_N clkgen.nor1/Y clkgen.nor1/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2b_1
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit VPWR clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit/in
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit/out VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_1_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.delay_155ns_1.genblk1\[4\].dly_binary.and_bypass_switch_B clkgen.delay_155ns_1.genblk1\[3\].dly_binary.out_mux/X
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit VPWR clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit/in
+ clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_6_16 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_7 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[2\].dly_binary.genblk1\[1\].delay_unit VPWR clkgen.delay_155ns_3.genblk1\[2\].dly_binary.genblk1\[1\].delay_unit/in
+ clkgen.delay_155ns_3.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_1.genblk1\[2\].control_invert dlycontrol1_in[2] clkgen.delay_155ns_1.genblk1\[2\].bypass_enable/B
+ VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[22\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[22\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[23\].delay_unit/in VGND
+ VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_edgedetect.dly_315ns_1.enablebuffer_A enable_dlycontrol_in VGND VPWR VPWR
+ VGND sky130_fd_sc_hd__diode_2
XANTENNA_outbuf_4_A sample_n_in VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_20_214 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[27\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[27\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[28\].delay_unit/in VGND
+ VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_11_214 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA_inbuf_3_A ndecision_finish_in VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_clkgen.delay_155ns_1.genblk1\[1\].control_invert_A dlycontrol1_in[1] VGND
+ VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_clkgen.delay_155ns_2.enablebuffer_A enable_dlycontrol_in VGND VPWR VPWR VGND
+ sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit VPWR clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit/in
+ clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_1_3 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_284 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_317 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xclkgen.delay_155ns_2.genblk1\[2\].dly_binary.genblk1\[0\].delay_unit VPWR clkgen.delay_155ns_2.genblk1\[2\].dly_binary.and_bypass_switch/X
+ clkgen.delay_155ns_2.genblk1\[2\].dly_binary.genblk1\[1\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_20_9 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.clkdig_inverter clkgen.clkdig_inverter/A outbuf_1/A VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_3_243 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_313 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_0 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkgen.delay_155ns_2.genblk1\[0\].control_invert_A dlycontrol2_in[0] VGND
+ VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_13_117 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xedgedetect.dly_315ns_1.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.out_mux/A0 VGND VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_14_245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit VPWR clkgen.delay_155ns_3.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit/in
+ clkgen.delay_155ns_3.genblk1\[1\].dly_binary.out_mux/A0 VGND VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_9_260 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_182 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_315 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_277 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XANTENNA_clkgen.delay_155ns_1.genblk1\[4\].dly_binary.out_mux_S clkgen.delay_155ns_1.genblk1\[4\].bypass_enable/X
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xedgedetect.dly_315ns_1.genblk1\[0\].dly_binary.out_mux VGND VPWR edgedetect.dly_315ns_1.genblk1\[0\].bypass_enable/X
+ inbuf_2/X edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.out_mux/A0 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.out_mux/X
+ VGND VPWR sky130_fd_sc_hd__mux2_1
XPHY_1 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xedgedetect.dly_315ns_1.genblk1\[2\].dly_binary.out_mux VGND VPWR edgedetect.dly_315ns_1.genblk1\[2\].bypass_enable/X
+ edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.out_mux/X edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.out_mux/A0
+ edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.out_mux/X VGND VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_edgedetect.dly_315ns_1.genblk1\[0\].bypass_enable_A edgedetect.dly_315ns_1.enablebuffer/X
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xedgedetect.dly_315ns_1.genblk1\[0\].dly_binary.and_bypass_switch edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.and_bypass_switch/X
+ edgedetect.dly_315ns_1.genblk1\[0\].bypass_enable/X inbuf_2/X VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__and2b_1
XFILLER_7_83 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_195 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xinbuf_1 VGND VPWR inbuf_1/X ena_in VGND VPWR sky130_fd_sc_hd__buf_1
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.out_mux VGND VPWR edgedetect.dly_315ns_1.genblk1\[4\].bypass_enable/X
+ edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.out_mux/X edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.out_mux/A0
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.out_mux/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_12_17 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_276 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_243 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_2.genblk1\[1\].dly_binary.genblk1\[0\].delay_unit VPWR clkgen.delay_155ns_2.genblk1\[1\].dly_binary.and_bypass_switch/X
+ clkgen.delay_155ns_2.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_4_62 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_172 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_16 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[2\].bypass_enable VPWR VGND edgedetect.dly_315ns_1.genblk1\[2\].bypass_enable/X
+ edgedetect.dly_315ns_1.genblk1\[2\].bypass_enable/B edgedetect.dly_315ns_1.enablebuffer/X
+ VGND VPWR sky130_fd_sc_hd__and2_1
Xclkgen.delay_155ns_2.genblk1\[3\].control_invert dlycontrol2_in[3] clkgen.delay_155ns_2.genblk1\[3\].bypass_enable/B
+ VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_1_63 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[10\].delay_unit VPWR clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit/out
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_3_289 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XANTENNA_clkgen.delay_155ns_2.genblk1\[4\].dly_binary.and_bypass_switch_A_N clkgen.delay_155ns_2.genblk1\[4\].bypass_enable/X
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_0_226 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_259 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[3\].bypass_enable VPWR VGND clkgen.delay_155ns_1.genblk1\[3\].bypass_enable/X
+ clkgen.delay_155ns_1.genblk1\[3\].bypass_enable/B clkgen.delay_155ns_1.enablebuffer/X
+ VGND VPWR sky130_fd_sc_hd__and2_1
XPHY_2 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xclkgen.delay_155ns_2.genblk1\[4\].bypass_enable VPWR VGND clkgen.delay_155ns_2.genblk1\[4\].bypass_enable/X
+ clkgen.delay_155ns_2.genblk1\[4\].bypass_enable/B clkgen.delay_155ns_2.enablebuffer/X
+ VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_7_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xinbuf_2 VGND VPWR inbuf_2/X start_conv_in VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_12_163 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA_clkgen.delay_155ns_1.genblk1\[2\].dly_binary.out_mux_S clkgen.delay_155ns_1.genblk1\[2\].bypass_enable/X
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit VPWR clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit/in
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.out_mux/A0 VGND VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_1.genblk1\[0\].dly_binary.out_mux VGND VPWR clkgen.delay_155ns_1.genblk1\[0\].bypass_enable/X
+ inbuf_3/X clkgen.delay_155ns_1.genblk1\[0\].dly_binary.out_mux/A0 clkgen.delay_155ns_1.genblk1\[0\].dly_binary.out_mux/X
+ VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_9_295 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[2\].dly_binary.out_mux VGND VPWR clkgen.delay_155ns_1.genblk1\[2\].bypass_enable/X
+ clkgen.delay_155ns_1.genblk1\[1\].dly_binary.out_mux/X clkgen.delay_155ns_1.genblk1\[2\].dly_binary.out_mux/A0
+ clkgen.delay_155ns_1.genblk1\[2\].dly_binary.out_mux/X VGND VPWR sky130_fd_sc_hd__mux2_1
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.out_mux VGND VPWR clkgen.delay_155ns_1.genblk1\[4\].bypass_enable/X
+ clkgen.delay_155ns_1.genblk1\[3\].dly_binary.out_mux/X clkgen.delay_155ns_1.genblk1\[4\].dly_binary.out_mux/A0
+ clkgen.clkdig_inverter/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_1_31 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[1\].dly_binary.and_bypass_switch edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.and_bypass_switch/X
+ edgedetect.dly_315ns_1.genblk1\[1\].bypass_enable/X edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.out_mux/X
+ VGND VPWR VGND VPWR sky130_fd_sc_hd__and2b_1
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[4\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[4\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[5\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_inbuf_1_A ena_in VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_19_125 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_238 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[2\].delay_unit VPWR clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[2\].delay_unit/in
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_2.genblk1\[0\].dly_binary.genblk1\[0\].delay_unit VPWR clkgen.delay_155ns_2.genblk1\[0\].dly_binary.and_bypass_switch/X
+ clkgen.delay_155ns_2.genblk1\[0\].dly_binary.out_mux/A0 VGND VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
XPHY_3 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_74 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xinbuf_3 VGND VPWR inbuf_3/X ndecision_finish_in VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_8_124 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_edgedetect.dly_315ns_1.genblk1\[5\].control_invert_A dlycontrol4_in[5] VGND
+ VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xedgedetect.dly_315ns_1.genblk1\[4\].control_invert dlycontrol4_in[4] edgedetect.dly_315ns_1.genblk1\[4\].bypass_enable/B
+ VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_1_311 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkgen.delay_155ns_1.genblk1\[0\].dly_binary.out_mux_S clkgen.delay_155ns_1.genblk1\[0\].bypass_enable/X
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[9\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[9\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[9\].delay_unit/out VGND
+ VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_13_84 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkgen.delay_155ns_2.genblk1\[0\].dly_binary.and_bypass_switch_B outbuf_1/A
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit VPWR clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit/in
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit VPWR clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit/in
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_20_19 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.delay_155ns_1.genblk1\[2\].dly_binary.and_bypass_switch_A_N clkgen.delay_155ns_1.genblk1\[2\].bypass_enable/X
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit VPWR clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit/in
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[2\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_3_214 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[0\].bypass_enable VPWR VGND clkgen.delay_155ns_3.genblk1\[0\].bypass_enable/X
+ clkgen.delay_155ns_3.genblk1\[0\].bypass_enable/B clkgen.delay_155ns_3.enablebuffer/X
+ VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_2_280 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XANTENNA_clkgen.delay_155ns_3.genblk1\[2\].bypass_enable_A clkgen.delay_155ns_3.enablebuffer/X
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_3.genblk1\[1\].dly_binary.out_mux VGND VPWR clkgen.delay_155ns_3.genblk1\[1\].bypass_enable/X
+ clkgen.delay_155ns_3.genblk1\[0\].dly_binary.out_mux/X clkgen.delay_155ns_3.genblk1\[1\].dly_binary.out_mux/A0
+ clkgen.delay_155ns_3.genblk1\[1\].dly_binary.out_mux/X VGND VPWR sky130_fd_sc_hd__mux2_1
XPHY_4 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xclkgen.delay_155ns_3.genblk1\[3\].dly_binary.out_mux VGND VPWR clkgen.delay_155ns_3.genblk1\[3\].bypass_enable/X
+ clkgen.delay_155ns_3.genblk1\[2\].dly_binary.out_mux/X clkgen.delay_155ns_3.genblk1\[3\].dly_binary.out_mux/A0
+ clkgen.delay_155ns_3.genblk1\[3\].dly_binary.out_mux/X VGND VPWR sky130_fd_sc_hd__mux2_1
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_3.genblk1\[4\].control_invert dlycontrol3_in[4] clkgen.delay_155ns_3.genblk1\[4\].bypass_enable/B
+ VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_4_32 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_150 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_74 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit VPWR clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit/in
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[2\].dly_binary.and_bypass_switch edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.and_bypass_switch/X
+ edgedetect.dly_315ns_1.genblk1\[2\].bypass_enable/X edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.out_mux/X
+ VGND VPWR VGND VPWR sky130_fd_sc_hd__and2b_1
XFILLER_13_260 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.delay_155ns_2.genblk1\[4\].dly_binary.out_mux_S clkgen.delay_155ns_2.genblk1\[4\].bypass_enable/X
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit VPWR clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit/in
+ clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_clkgen.delay_155ns_1.genblk1\[0\].control_invert_A dlycontrol1_in[0] VGND
+ VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[0\].delay_unit VPWR clkgen.delay_155ns_1.genblk1\[4\].dly_binary.and_bypass_switch/X
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_3_259 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_292 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[11\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[11\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[12\].delay_unit/in VGND
+ VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_clkgen.delay_155ns_3.genblk1\[2\].bypass_enable_B clkgen.delay_155ns_3.genblk1\[2\].bypass_enable/B
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_8_307 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit VPWR clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit/in
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit/out VGND
+ VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
XPHY_5 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit VPWR clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit/in
+ clkgen.delay_155ns_3.genblk1\[3\].dly_binary.out_mux/A0 VGND VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit/in VGND
+ VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_17_214 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit VPWR clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit/in
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_4_173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit VPWR clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit/in
+ clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_13_272 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_254 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_143 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[16\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[16\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[17\].delay_unit/in VGND
+ VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.and_bypass_switch_A_N edgedetect.dly_315ns_1.genblk1\[1\].bypass_enable/X
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_5_290 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_63 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.delay_155ns_2.genblk1\[2\].dly_binary.out_mux_S clkgen.delay_155ns_2.genblk1\[2\].bypass_enable/X
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_18_183 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_260 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[0\].control_invert dlycontrol1_in[0] clkgen.delay_155ns_1.genblk1\[0\].bypass_enable/B
+ VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_208 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_15_175 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_6 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_22 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit VPWR clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit/in
+ clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_3.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit VPWR clkgen.delay_155ns_3.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit/in
+ clkgen.delay_155ns_3.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[3\].dly_binary.and_bypass_switch edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.and_bypass_switch/X
+ edgedetect.dly_315ns_1.genblk1\[3\].bypass_enable/X edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.out_mux/X
+ VGND VPWR VGND VPWR sky130_fd_sc_hd__and2b_1
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[23\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[23\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[24\].delay_unit/in VGND
+ VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_edgedetect.dly_315ns_1.genblk1\[3\].bypass_enable_A edgedetect.dly_315ns_1.enablebuffer/X
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[0\].delay_unit VPWR clkgen.delay_155ns_1.genblk1\[3\].dly_binary.and_bypass_switch/X
+ clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_13_240 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_247 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.out_mux_S edgedetect.dly_315ns_1.genblk1\[4\].bypass_enable/X
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_19_31 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_272 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[28\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[28\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[29\].delay_unit/in VGND
+ VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit VPWR clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit/in
+ clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[30\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[30\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[31\].delay_unit/in VGND
+ VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_15_143 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA_clkgen.delay_155ns_2.genblk1\[0\].dly_binary.out_mux_S clkgen.delay_155ns_2.genblk1\[0\].bypass_enable/X
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XPHY_7 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xclkgen.delay_155ns_2.genblk1\[2\].dly_binary.genblk1\[1\].delay_unit VPWR clkgen.delay_155ns_2.genblk1\[2\].dly_binary.genblk1\[1\].delay_unit/in
+ clkgen.delay_155ns_2.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_16_43 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_124 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_164 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_208 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.enablebuffer VPWR VGND edgedetect.dly_315ns_1.enablebuffer/X
+ enable_dlycontrol_in VGND VPWR sky130_fd_sc_hd__buf_4
Xclkgen.delay_155ns_1.genblk1\[2\].dly_binary.genblk1\[0\].delay_unit VPWR clkgen.delay_155ns_1.genblk1\[2\].dly_binary.and_bypass_switch/X
+ clkgen.delay_155ns_1.genblk1\[2\].dly_binary.genblk1\[1\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.and_bypass_switch edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.and_bypass_switch/X
+ edgedetect.dly_315ns_1.genblk1\[4\].bypass_enable/X edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.out_mux/X
+ VGND VPWR VGND VPWR sky130_fd_sc_hd__and2b_1
XFILLER_16_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_8 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_302 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XANTENNA_edgedetect.dly_315ns_1.genblk1\[4\].control_invert_A dlycontrol4_in[4] VGND
+ VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_4_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.enablebuffer VPWR VGND clkgen.delay_155ns_1.enablebuffer/X enable_dlycontrol_in
+ VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_13_56 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xedgedetect.dly_315ns_1.genblk1\[3\].bypass_enable VPWR VGND edgedetect.dly_315ns_1.genblk1\[3\].bypass_enable/X
+ edgedetect.dly_315ns_1.genblk1\[3\].bypass_enable/B edgedetect.dly_315ns_1.enablebuffer/X
+ VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_5_90 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xclkgen.delay_155ns_2.genblk1\[1\].control_invert dlycontrol2_in[1] clkgen.delay_155ns_2.genblk1\[1\].bypass_enable/B
+ VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
Xclkgen.delay_155ns_2.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit VPWR clkgen.delay_155ns_2.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit/in
+ clkgen.delay_155ns_2.genblk1\[1\].dly_binary.out_mux/A0 VGND VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_5_260 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_315 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[4\].bypass_enable VPWR VGND clkgen.delay_155ns_1.genblk1\[4\].bypass_enable/X
+ clkgen.delay_155ns_1.genblk1\[4\].bypass_enable/B clkgen.delay_155ns_1.enablebuffer/X
+ VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_2_230 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[0\].dly_binary.and_bypass_switch clkgen.delay_155ns_3.genblk1\[0\].dly_binary.and_bypass_switch/X
+ clkgen.delay_155ns_3.genblk1\[0\].bypass_enable/X clkgen.nor1/Y VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__and2b_1
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit VPWR clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit/in
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XPHY_9 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_56 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.delay_155ns_1.genblk1\[4\].dly_binary.out_mux_A0 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.out_mux/A0
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_4_314 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA_clkgen.delay_155ns_1.enablebuffer_A enable_dlycontrol_in VGND VPWR VPWR VGND
+ sky130_fd_sc_hd__diode_2
XFILLER_11_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.delay_155ns_2.genblk1\[2\].dly_binary.and_bypass_switch_A_N clkgen.delay_155ns_2.genblk1\[2\].bypass_enable/X
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[0\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.and_bypass_switch/X
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[1\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_13_254 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[1\].dly_binary.genblk1\[0\].delay_unit VPWR clkgen.delay_155ns_1.genblk1\[1\].dly_binary.and_bypass_switch/X
+ clkgen.delay_155ns_1.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_18_313 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_272 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.and_bypass_switch edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.and_bypass_switch/X
+ edgedetect.dly_315ns_1.genblk1\[5\].bypass_enable/X edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.out_mux/X
+ VGND VPWR VGND VPWR sky130_fd_sc_hd__and2b_1
XFILLER_15_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_242 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_90 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[5\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[5\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[6\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_clkgen.delay_155ns_1.genblk1\[4\].dly_binary.out_mux_A1 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.out_mux/X
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xedgedetect.dly_315ns_1.genblk1\[2\].control_invert dlycontrol4_in[2] edgedetect.dly_315ns_1.genblk1\[2\].bypass_enable/B
+ VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_1_307 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit VPWR clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit/in
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_16_285 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_16 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_266 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_218 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_2.genblk1\[0\].bypass_enable VPWR VGND clkgen.delay_155ns_2.genblk1\[0\].bypass_enable/X
+ clkgen.delay_155ns_2.genblk1\[0\].bypass_enable/B clkgen.delay_155ns_2.enablebuffer/X
+ VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_5_284 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[1\].bypass_enable VPWR VGND clkgen.delay_155ns_3.genblk1\[1\].bypass_enable/X
+ clkgen.delay_155ns_3.genblk1\[1\].bypass_enable/B clkgen.delay_155ns_3.enablebuffer/X
+ VGND VPWR sky130_fd_sc_hd__and2_1
Xclkgen.delay_155ns_3.genblk1\[1\].dly_binary.and_bypass_switch clkgen.delay_155ns_3.genblk1\[1\].dly_binary.and_bypass_switch/X
+ clkgen.delay_155ns_3.genblk1\[1\].bypass_enable/X clkgen.delay_155ns_3.genblk1\[0\].dly_binary.out_mux/X
+ VGND VPWR VGND VPWR sky130_fd_sc_hd__and2b_1
XFILLER_10_59 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_254 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit VPWR clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit/in
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_clkgen.delay_155ns_3.genblk1\[4\].control_invert_A dlycontrol3_in[4] VGND
+ VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit VPWR clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit/in
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_2.genblk1\[0\].dly_binary.and_bypass_switch clkgen.delay_155ns_2.genblk1\[0\].dly_binary.and_bypass_switch/X
+ clkgen.delay_155ns_2.genblk1\[0\].bypass_enable/X outbuf_1/A VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__and2b_1
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[0\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.and_bypass_switch/X
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[2\].delay_unit VPWR clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[2\].delay_unit/in
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_14_3 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xclkgen.delay_155ns_1.genblk1\[0\].dly_binary.genblk1\[0\].delay_unit VPWR clkgen.delay_155ns_1.genblk1\[0\].dly_binary.and_bypass_switch/X
+ clkgen.delay_155ns_1.genblk1\[0\].dly_binary.out_mux/A0 VGND VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_clkgen.delay_155ns_1.genblk1\[0\].dly_binary.and_bypass_switch_A_N clkgen.delay_155ns_1.genblk1\[0\].bypass_enable/X
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_3.genblk1\[2\].control_invert dlycontrol3_in[2] clkgen.delay_155ns_3.genblk1\[2\].bypass_enable/B
+ VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_13_278 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_204 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_208 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_5_241 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit VPWR clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit/in
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_10_16 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_200 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_266 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit VPWR clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit/in
+ clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_14_170 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit VPWR clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit/in
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[2\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_20_173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_155 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[12\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[12\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[13\].delay_unit/in VGND
+ VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_2.genblk1\[1\].dly_binary.out_mux VGND VPWR clkgen.delay_155ns_2.genblk1\[1\].bypass_enable/X
+ clkgen.delay_155ns_2.genblk1\[0\].dly_binary.out_mux/X clkgen.delay_155ns_2.genblk1\[1\].dly_binary.out_mux/A0
+ clkgen.delay_155ns_2.genblk1\[1\].dly_binary.out_mux/X VGND VPWR sky130_fd_sc_hd__mux2_1
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit VPWR clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit/in
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.and_bypass_switch_A_N edgedetect.dly_315ns_1.genblk1\[4\].bypass_enable/X
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_2.genblk1\[3\].dly_binary.out_mux VGND VPWR clkgen.delay_155ns_2.genblk1\[3\].bypass_enable/X
+ clkgen.delay_155ns_2.genblk1\[2\].dly_binary.out_mux/X clkgen.delay_155ns_2.genblk1\[3\].dly_binary.out_mux/A0
+ clkgen.delay_155ns_2.genblk1\[3\].dly_binary.out_mux/X VGND VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_clkgen.delay_155ns_3.genblk1\[0\].bypass_enable_A clkgen.delay_155ns_3.enablebuffer/X
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_13_224 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[2\].dly_binary.and_bypass_switch clkgen.delay_155ns_3.genblk1\[2\].dly_binary.and_bypass_switch/X
+ clkgen.delay_155ns_3.genblk1\[2\].bypass_enable/X clkgen.delay_155ns_3.genblk1\[1\].dly_binary.out_mux/X
+ VGND VPWR VGND VPWR sky130_fd_sc_hd__and2b_1
XFILLER_9_217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_194 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_183 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit/in VGND
+ VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_8_272 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xclkgen.delay_155ns_2.genblk1\[1\].dly_binary.and_bypass_switch clkgen.delay_155ns_2.genblk1\[1\].dly_binary.and_bypass_switch/X
+ clkgen.delay_155ns_2.genblk1\[1\].bypass_enable/X clkgen.delay_155ns_2.genblk1\[0\].dly_binary.out_mux/X
+ VGND VPWR VGND VPWR sky130_fd_sc_hd__and2b_1
Xedgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[0\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.and_bypass_switch/X
+ edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit VPWR clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit/in
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit VPWR clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit/in
+ clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_2_223 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_124 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[17\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[17\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[18\].delay_unit/in VGND
+ VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_1.genblk1\[0\].dly_binary.and_bypass_switch clkgen.delay_155ns_1.genblk1\[0\].dly_binary.and_bypass_switch/X
+ clkgen.delay_155ns_1.genblk1\[0\].bypass_enable/X inbuf_3/X VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__and2b_1
XFILLER_2_62 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_300 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_315 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_16 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_152 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_152 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_112 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_94 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_3_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit VPWR clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit/in
+ clkgen.delay_155ns_2.genblk1\[3\].dly_binary.out_mux/A0 VGND VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_edgedetect.dly_315ns_1.genblk1\[3\].control_invert_A dlycontrol4_in[3] VGND
+ VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_13_17 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[3\].control_invert dlycontrol1_in[3] clkgen.delay_155ns_1.genblk1\[3\].bypass_enable/B
+ VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
Xclkgen.delay_155ns_3.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit VPWR clkgen.delay_155ns_3.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit/in
+ clkgen.delay_155ns_3.genblk1\[2\].dly_binary.out_mux/A0 VGND VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[24\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[24\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[25\].delay_unit/in VGND
+ VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit VPWR clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit/in
+ clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_5_232 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_254 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_164 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[29\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[29\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[30\].delay_unit/in VGND
+ VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_3.genblk1\[3\].dly_binary.and_bypass_switch clkgen.delay_155ns_3.genblk1\[3\].dly_binary.and_bypass_switch/X
+ clkgen.delay_155ns_3.genblk1\[3\].bypass_enable/X clkgen.delay_155ns_3.genblk1\[2\].dly_binary.out_mux/X
+ VGND VPWR VGND VPWR sky130_fd_sc_hd__and2b_1
Xedgedetect.dly_315ns_1.genblk1\[2\].dly_binary.genblk1\[0\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.and_bypass_switch/X
+ edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.genblk1\[1\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_8_62 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit VPWR clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit/in
+ clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_17_71 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_212 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[31\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[31\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.out_mux/A0 VGND VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_0_311 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
Xclkgen.delay_155ns_2.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit VPWR clkgen.delay_155ns_2.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit/in
+ clkgen.delay_155ns_2.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_2.genblk1\[2\].dly_binary.and_bypass_switch clkgen.delay_155ns_2.genblk1\[2\].dly_binary.and_bypass_switch/X
+ clkgen.delay_155ns_2.genblk1\[2\].bypass_enable/X clkgen.delay_155ns_2.genblk1\[1\].dly_binary.out_mux/X
+ VGND VPWR VGND VPWR sky130_fd_sc_hd__and2b_1
XFILLER_12_270 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_307 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[1\].dly_binary.and_bypass_switch clkgen.delay_155ns_1.genblk1\[1\].dly_binary.and_bypass_switch/X
+ clkgen.delay_155ns_1.genblk1\[1\].bypass_enable/X clkgen.delay_155ns_1.genblk1\[0\].dly_binary.out_mux/X
+ VGND VPWR VGND VPWR sky130_fd_sc_hd__and2b_1
XFILLER_14_94 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_266 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_edgedetect.dly_315ns_1.genblk1\[1\].bypass_enable_A edgedetect.dly_315ns_1.enablebuffer/X
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_2_236 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_276 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_243 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[2\].dly_binary.genblk1\[1\].delay_unit VPWR clkgen.delay_155ns_1.genblk1\[2\].dly_binary.genblk1\[1\].delay_unit/in
+ clkgen.delay_155ns_1.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[4\].bypass_enable VPWR VGND edgedetect.dly_315ns_1.genblk1\[4\].bypass_enable/X
+ edgedetect.dly_315ns_1.genblk1\[4\].bypass_enable/B edgedetect.dly_315ns_1.enablebuffer/X
+ VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_5_31 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.delay_155ns_2.genblk1\[4\].control_invert_A dlycontrol2_in[4] VGND
+ VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_outbuf_5_A nsample_p_in VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_5_223 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_278 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_2.enablebuffer VPWR VGND clkgen.delay_155ns_2.enablebuffer/X enable_dlycontrol_in
+ VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_2_248 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_303 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xedgedetect.dly_315ns_1.genblk1\[1\].dly_binary.genblk1\[0\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.and_bypass_switch/X
+ edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_2_32 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.and_bypass_switch clkgen.delay_155ns_3.genblk1\[4\].dly_binary.and_bypass_switch/X
+ clkgen.delay_155ns_3.genblk1\[4\].bypass_enable/X clkgen.delay_155ns_3.genblk1\[3\].dly_binary.out_mux/X
+ VGND VPWR VGND VPWR sky130_fd_sc_hd__and2b_1
XANTENNA_clkgen.delay_155ns_3.genblk1\[3\].control_invert_A dlycontrol3_in[3] VGND
+ VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.out_mux_A0 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.out_mux/A0
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_14_163 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_3 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xclkgen.delay_155ns_2.genblk1\[4\].control_invert dlycontrol2_in[4] clkgen.delay_155ns_2.genblk1\[4\].bypass_enable/B
+ VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
Xclkgen.delay_155ns_2.genblk1\[3\].dly_binary.and_bypass_switch clkgen.delay_155ns_2.genblk1\[3\].dly_binary.and_bypass_switch/X
+ clkgen.delay_155ns_2.genblk1\[3\].bypass_enable/X clkgen.delay_155ns_2.genblk1\[2\].dly_binary.out_mux/X
+ VGND VPWR VGND VPWR sky130_fd_sc_hd__and2b_1
XFILLER_16_247 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_203 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[2\].dly_binary.and_bypass_switch clkgen.delay_155ns_1.genblk1\[2\].dly_binary.and_bypass_switch/X
+ clkgen.delay_155ns_1.genblk1\[2\].bypass_enable/X clkgen.delay_155ns_1.genblk1\[1\].dly_binary.out_mux/X
+ VGND VPWR VGND VPWR sky130_fd_sc_hd__and2b_1
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit VPWR clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit/in
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[1\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[1\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[2\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_4_290 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XANTENNA_clkgen.delay_155ns_2.genblk1\[0\].dly_binary.and_bypass_switch_A_N clkgen.delay_155ns_2.genblk1\[0\].bypass_enable/X
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XPHY_40 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_183 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_271 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xclkgen.delay_155ns_1.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit VPWR clkgen.delay_155ns_1.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit/in
+ clkgen.delay_155ns_1.genblk1\[1\].dly_binary.out_mux/A0 VGND VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_20_315 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_315 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.clkdig_inverter_A clkgen.clkdig_inverter/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_11_31 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_311 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_32 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[0\].control_invert dlycontrol4_in[0] edgedetect.dly_315ns_1.genblk1\[0\].bypass_enable/B
+ VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[6\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[6\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[7\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_3_152 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[0\].bypass_enable VPWR VGND clkgen.delay_155ns_1.genblk1\[0\].bypass_enable/X
+ clkgen.delay_155ns_1.genblk1\[0\].bypass_enable/B clkgen.delay_155ns_1.enablebuffer/X
+ VGND VPWR sky130_fd_sc_hd__and2_1
Xedgedetect.dly_315ns_1.genblk1\[0\].dly_binary.genblk1\[0\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.and_bypass_switch/X
+ edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.out_mux/A0 VGND VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_8_200 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_2.genblk1\[1\].bypass_enable VPWR VGND clkgen.delay_155ns_2.genblk1\[1\].bypass_enable/X
+ clkgen.delay_155ns_2.genblk1\[1\].bypass_enable/B clkgen.delay_155ns_2.enablebuffer/X
+ VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_12_284 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
Xclkgen.delay_155ns_3.genblk1\[2\].bypass_enable VPWR VGND clkgen.delay_155ns_3.genblk1\[2\].bypass_enable/X
+ clkgen.delay_155ns_3.genblk1\[2\].bypass_enable/B clkgen.delay_155ns_3.enablebuffer/X
+ VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_10_3 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_266 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit VPWR clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit/in
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[10\].delay_unit VPWR clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit/out
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_clkgen.delay_155ns_3.genblk1\[3\].bypass_enable_A clkgen.delay_155ns_3.enablebuffer/X
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xedgedetect.dly_315ns_1.genblk1\[5\].control_invert dlycontrol4_in[5] edgedetect.dly_315ns_1.genblk1\[5\].bypass_enable/B
+ VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XPHY_41 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_30 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_313 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_283 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.and_bypass_switch clkgen.delay_155ns_2.genblk1\[4\].dly_binary.and_bypass_switch/X
+ clkgen.delay_155ns_2.genblk1\[4\].bypass_enable/X clkgen.delay_155ns_2.genblk1\[3\].dly_binary.out_mux/X
+ VGND VPWR VGND VPWR sky130_fd_sc_hd__and2b_1
XANTENNA_clkgen.delay_155ns_1.genblk1\[3\].dly_binary.and_bypass_switch_A_N clkgen.delay_155ns_1.genblk1\[3\].bypass_enable/X
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_1.genblk1\[3\].dly_binary.and_bypass_switch clkgen.delay_155ns_1.genblk1\[3\].dly_binary.and_bypass_switch/X
+ clkgen.delay_155ns_1.genblk1\[3\].bypass_enable/X clkgen.delay_155ns_1.genblk1\[2\].dly_binary.out_mux/X
+ VGND VPWR VGND VPWR sky130_fd_sc_hd__and2b_1
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit VPWR clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit/in
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit/out VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_3_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit VPWR clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit/in
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.out_mux/A0 VGND VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_0_304 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[2\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_17_31 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[0\].control_invert dlycontrol3_in[0] clkgen.delay_155ns_3.genblk1\[0\].bypass_enable/B
+ VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit VPWR clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit/in
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_12_7 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_252 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_edgedetect.dly_315ns_1.genblk1\[2\].control_invert_A dlycontrol4_in[2] VGND
+ VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XPHY_31 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA_outbuf_3_A sample_p_in VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XPHY_20 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_152 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_295 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[1\].dly_binary.out_mux VGND VPWR edgedetect.dly_315ns_1.genblk1\[1\].bypass_enable/X
+ edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.out_mux/X edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.out_mux/A0
+ edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.out_mux/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_11_306 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_199 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit VPWR clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit/in
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[3\].dly_binary.out_mux VGND VPWR edgedetect.dly_315ns_1.genblk1\[3\].bypass_enable/X
+ edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.out_mux/X edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.out_mux/A0
+ edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.out_mux/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_19_214 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.out_mux VGND VPWR edgedetect.dly_315ns_1.genblk1\[5\].bypass_enable/X
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.out_mux/X edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.out_mux/A0
+ edgedetect.nor1/A VGND VPWR sky130_fd_sc_hd__mux2_1
Xclkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit VPWR clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit/in
+ clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_inbuf_2_A start_conv_in VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_0_3 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[2\].delay_unit VPWR clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[2\].delay_unit/in
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_clkgen.delay_155ns_1.genblk1\[3\].dly_binary.out_mux_S clkgen.delay_155ns_1.genblk1\[3\].bypass_enable/X
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[13\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[13\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[14\].delay_unit/in VGND
+ VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_12_264 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit VPWR clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit/in
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_14_88 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_32 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.and_bypass_switch clkgen.delay_155ns_1.genblk1\[4\].dly_binary.and_bypass_switch/X
+ clkgen.delay_155ns_1.genblk1\[4\].bypass_enable/X clkgen.delay_155ns_1.genblk1\[3\].dly_binary.out_mux/X
+ VGND VPWR VGND VPWR sky130_fd_sc_hd__and2b_1
XPHY_10 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit/in VGND
+ VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
Xoutbuf_1 VPWR VGND clk_dig_out outbuf_1/A VGND VPWR sky130_fd_sc_hd__buf_4
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit VPWR clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit/in
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_edgedetect.dly_315ns_1.genblk1\[4\].bypass_enable_A edgedetect.dly_315ns_1.enablebuffer/X
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit VPWR clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit/in
+ clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[18\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[18\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[19\].delay_unit/in VGND
+ VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_clkgen.delay_155ns_1.genblk1\[4\].control_invert_A dlycontrol1_in[4] VGND
+ VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_16_218 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[20\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[20\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[21\].delay_unit/in VGND
+ VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_1.genblk1\[1\].control_invert dlycontrol1_in[1] clkgen.delay_155ns_1.genblk1\[1\].bypass_enable/B
+ VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
Xclkgen.delay_155ns_1.genblk1\[1\].dly_binary.out_mux VGND VPWR clkgen.delay_155ns_1.genblk1\[1\].bypass_enable/X
+ clkgen.delay_155ns_1.genblk1\[0\].dly_binary.out_mux/X clkgen.delay_155ns_1.genblk1\[1\].dly_binary.out_mux/A0
+ clkgen.delay_155ns_1.genblk1\[1\].dly_binary.out_mux/X VGND VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_edgedetect.nor1_B_N inbuf_2/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_12_276 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xedgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_1.genblk1\[3\].dly_binary.out_mux VGND VPWR clkgen.delay_155ns_1.genblk1\[3\].bypass_enable/X
+ clkgen.delay_155ns_1.genblk1\[2\].dly_binary.out_mux/X clkgen.delay_155ns_1.genblk1\[3\].dly_binary.out_mux/A0
+ clkgen.delay_155ns_1.genblk1\[3\].dly_binary.out_mux/X VGND VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_clkgen.delay_155ns_1.genblk1\[1\].dly_binary.out_mux_S clkgen.delay_155ns_1.genblk1\[1\].bypass_enable/X
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_clkgen.delay_155ns_2.genblk1\[3\].control_invert_A dlycontrol2_in[3] VGND
+ VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XPHY_33 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_11 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[25\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[25\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[26\].delay_unit/in VGND
+ VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit VPWR clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit/in
+ clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
Xoutbuf_2 VPWR VGND clk_comp_out outbuf_2/A VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_14_124 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.delay_155ns_3.genblk1\[2\].control_invert_A dlycontrol3_in[2] VGND
+ VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_19_3 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_164 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_78 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_90 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_259 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[2\].dly_binary.genblk1\[1\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.genblk1\[1\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit VPWR clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit/in
+ clkgen.delay_155ns_1.genblk1\[3\].dly_binary.out_mux/A0 VGND VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_2.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit VPWR clkgen.delay_155ns_2.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit/in
+ clkgen.delay_155ns_2.genblk1\[2\].dly_binary.out_mux/A0 VGND VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_4_251 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_284 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_12 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_16 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xoutbuf_3 VPWR VGND sample_p_out sample_p_in VGND VPWR sky130_fd_sc_hd__buf_4
Xclkgen.delay_155ns_3.genblk1\[0\].dly_binary.out_mux VGND VPWR clkgen.delay_155ns_3.genblk1\[0\].bypass_enable/X
+ clkgen.nor1/Y clkgen.delay_155ns_3.genblk1\[0\].dly_binary.out_mux/A0 clkgen.delay_155ns_3.genblk1\[0\].dly_binary.out_mux/X
+ VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_6_313 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xclkgen.delay_155ns_3.genblk1\[2\].dly_binary.out_mux VGND VPWR clkgen.delay_155ns_3.genblk1\[2\].bypass_enable/X
+ clkgen.delay_155ns_3.genblk1\[1\].dly_binary.out_mux/X clkgen.delay_155ns_3.genblk1\[2\].dly_binary.out_mux/A0
+ clkgen.delay_155ns_3.genblk1\[2\].dly_binary.out_mux/X VGND VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_outbuf_1_A outbuf_1/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xedgedetect.dly_315ns_1.genblk1\[5\].bypass_enable VPWR VGND edgedetect.dly_315ns_1.genblk1\[5\].bypass_enable/X
+ edgedetect.dly_315ns_1.genblk1\[5\].bypass_enable/B edgedetect.dly_315ns_1.enablebuffer/X
+ VGND VPWR sky130_fd_sc_hd__and2_1
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.out_mux VGND VPWR clkgen.delay_155ns_3.genblk1\[4\].bypass_enable/X
+ clkgen.delay_155ns_3.genblk1\[3\].dly_binary.out_mux/X clkgen.delay_155ns_3.genblk1\[4\].dly_binary.out_mux/A0
+ outbuf_2/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_6_198 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit VPWR clkgen.delay_155ns_1.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit/in
+ clkgen.delay_155ns_1.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_17_315 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_263 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_35 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_307 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_24 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_13 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xoutbuf_4 VPWR VGND sample_n_out sample_n_in VGND VPWR sky130_fd_sc_hd__buf_4
Xclkgen.delay_155ns_3.enablebuffer VPWR VGND clkgen.delay_155ns_3.enablebuffer/X enable_dlycontrol_in
+ VGND VPWR sky130_fd_sc_hd__buf_4
XANTENNA_clkgen.delay_155ns_2.genblk1\[3\].dly_binary.out_mux_S clkgen.delay_155ns_2.genblk1\[3\].bypass_enable/X
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_2.genblk1\[2\].control_invert dlycontrol2_in[2] clkgen.delay_155ns_2.genblk1\[2\].bypass_enable/B
+ VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_3_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.out_mux/A0 VGND VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_8_16 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.delay_155ns_2.genblk1\[4\].dly_binary.out_mux_A0 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.out_mux/A0
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_15_276 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_243 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_191 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.delay_155ns_2.genblk1\[3\].dly_binary.and_bypass_switch_A_N clkgen.delay_155ns_2.genblk1\[3\].bypass_enable/X
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_14_59 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_edgedetect.dly_315ns_1.genblk1\[1\].control_invert_A dlycontrol4_in[1] VGND
+ VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit VPWR clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit/in
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_17_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_275 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_36 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xedgedetect.dly_315ns_1.genblk1\[0\].bypass_enable VPWR VGND edgedetect.dly_315ns_1.genblk1\[0\].bypass_enable/X
+ edgedetect.dly_315ns_1.genblk1\[0\].bypass_enable/B edgedetect.dly_315ns_1.enablebuffer/X
+ VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_9_301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xoutbuf_5 VPWR VGND nsample_p_out nsample_p_in VGND VPWR sky130_fd_sc_hd__buf_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[2\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[2\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[3\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.and_bypass_switch_B inbuf_2/X
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_18_274 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_174 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[0\].delay_unit VPWR clkgen.delay_155ns_3.genblk1\[4\].dly_binary.and_bypass_switch/X
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_1.genblk1\[1\].bypass_enable VPWR VGND clkgen.delay_155ns_1.genblk1\[1\].bypass_enable/X
+ clkgen.delay_155ns_1.genblk1\[1\].bypass_enable/B clkgen.delay_155ns_1.enablebuffer/X
+ VGND VPWR sky130_fd_sc_hd__and2_1
Xclkgen.delay_155ns_2.genblk1\[2\].bypass_enable VPWR VGND clkgen.delay_155ns_2.genblk1\[2\].bypass_enable/X
+ clkgen.delay_155ns_2.genblk1\[2\].bypass_enable/B clkgen.delay_155ns_2.enablebuffer/X
+ VGND VPWR sky130_fd_sc_hd__and2_1
XANTENNA_clkgen.delay_155ns_2.genblk1\[1\].dly_binary.out_mux_S clkgen.delay_155ns_2.genblk1\[1\].bypass_enable/X
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_17_3 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xclkgen.delay_155ns_3.genblk1\[3\].bypass_enable VPWR VGND clkgen.delay_155ns_3.genblk1\[3\].bypass_enable/X
+ clkgen.delay_155ns_3.genblk1\[3\].bypass_enable/B clkgen.delay_155ns_3.enablebuffer/X
+ VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_20_291 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_258 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[7\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[7\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[8\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_14_16 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[3\].control_invert dlycontrol4_in[3] edgedetect.dly_315ns_1.genblk1\[3\].bypass_enable/B
+ VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XPHY_37 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_94 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit VPWR clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit/in
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit VPWR clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit/in
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
Xoutbuf_6 VPWR VGND nsample_n_out nsample_n_in VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_13_194 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_187 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_124 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.out_mux_S edgedetect.dly_315ns_1.genblk1\[3\].bypass_enable/X
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_clkgen.delay_155ns_1.genblk1\[3\].control_invert_A dlycontrol1_in[3] VGND
+ VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_0_63 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_204 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.delay_155ns_1.genblk1\[1\].dly_binary.and_bypass_switch_A_N clkgen.delay_155ns_1.genblk1\[1\].bypass_enable/X
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_clkgen.delay_155ns_2.genblk1\[0\].dly_binary.out_mux_A1 outbuf_1/A VGND VPWR
+ VPWR VGND sky130_fd_sc_hd__diode_2
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[2\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[2\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XPHY_38 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit VPWR clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit/in
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XPHY_16 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkgen.delay_155ns_2.genblk1\[2\].control_invert_A dlycontrol2_in[2] VGND
+ VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_6_62 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[3\].control_invert dlycontrol3_in[3] clkgen.delay_155ns_3.genblk1\[3\].bypass_enable/B
+ VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
Xclkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[0\].delay_unit VPWR clkgen.delay_155ns_3.genblk1\[3\].dly_binary.and_bypass_switch/X
+ clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_1_214 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_280 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_313 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA_clkgen.delay_155ns_3.enablebuffer_A enable_dlycontrol_in VGND VPWR VPWR VGND
+ sky130_fd_sc_hd__diode_2
XFILLER_7_3 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_63 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.delay_155ns_3.genblk1\[1\].control_invert_A dlycontrol3_in[1] VGND
+ VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_clkgen.delay_155ns_3.genblk1\[1\].bypass_enable_A clkgen.delay_155ns_3.enablebuffer/X
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_12_94 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_121 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit VPWR clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit/in
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit/out VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_9_40 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.out_mux_S edgedetect.dly_315ns_1.genblk1\[1\].bypass_enable/X
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit VPWR clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit/in
+ clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_8_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[10\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit/out
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit/in VGND
+ VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_11_282 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit VPWR clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit/in
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_20_94 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_212 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_28 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_17 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_259 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[14\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[14\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[15\].delay_unit/in VGND
+ VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_9_315 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit VPWR clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit/in
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_0_292 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_178 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_31 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.out_mux/A0 VGND VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_12_62 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit VPWR clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit/in
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_15_214 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xclkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit VPWR clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit/in
+ clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_3.genblk1\[2\].dly_binary.genblk1\[0\].delay_unit VPWR clkgen.delay_155ns_3.genblk1\[2\].dly_binary.and_bypass_switch/X
+ clkgen.delay_155ns_3.genblk1\[2\].dly_binary.genblk1\[1\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_18_94 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[19\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[19\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[20\].delay_unit/in VGND
+ VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_11_294 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_243 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[21\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[21\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[22\].delay_unit/in VGND
+ VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_15_3 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA_edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.out_mux_A1 inbuf_2/X VGND
+ VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_7_276 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_202 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_117 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_29 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_18 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_227 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.out_mux/A0 VGND VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_0_271 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
Xclkgen.delay_155ns_1.genblk1\[4\].control_invert dlycontrol1_in[4] clkgen.delay_155ns_1.genblk1\[4\].bypass_enable/B
+ VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_16_194 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_153 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_167 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[26\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[26\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[27\].delay_unit/in VGND
+ VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_18_245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit VPWR clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit/in
+ clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_9_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_edgedetect.dly_315ns_1.genblk1\[2\].bypass_enable_A edgedetect.dly_315ns_1.enablebuffer/X
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_18_62 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_63 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA_edgedetect.dly_315ns_1.genblk1\[0\].control_invert_A dlycontrol4_in[0] VGND
+ VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_4_269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_32 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_19 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_239 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_17_107 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_63 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[1\].dly_binary.genblk1\[0\].delay_unit VPWR clkgen.delay_155ns_3.genblk1\[1\].dly_binary.and_bypass_switch/X
+ clkgen.delay_155ns_3.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_9_136 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_191 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_3 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_183 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_194 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_182 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_3 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_31 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_307 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xclkgen.delay_155ns_1.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit VPWR clkgen.delay_155ns_1.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit/in
+ clkgen.delay_155ns_1.genblk1\[2\].dly_binary.out_mux/A0 VGND VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
C0 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.out_mux/X VGND 1.60fF
C1 dlycontrol4_in[5] nsample_p_out 1.09fF
C2 VGND outbuf_1/A 5.38fF
C3 VPWR clkgen.delay_155ns_2.genblk1\[4\].dly_binary.out_mux/A0 5.54fF
C4 dlycontrol1_in[0] clkgen.delay_155ns_1.genblk1\[4\].bypass_enable/X 1.22fF
C5 VPWR clkgen.delay_155ns_2.genblk1\[2\].bypass_enable/B 1.11fF
C6 VGND clkgen.delay_155ns_2.genblk1\[2\].bypass_enable/X 9.03fF
C7 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[12\].delay_unit/in VPWR 1.03fF
C8 clkgen.delay_155ns_1.genblk1\[0\].bypass_enable/X VGND 4.11fF
C9 dlycontrol3_in[1] clkgen.delay_155ns_3.genblk1\[1\].bypass_enable/B 1.82fF
C10 clkgen.delay_155ns_3.genblk1\[4\].bypass_enable/X VPWR 2.16fF
C11 enable_dlycontrol_in VPWR 9.87fF
C12 dlycontrol1_in[0] dlycontrol1_in[1] 1.30fF
C13 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.out_mux/A0 VGND 1.06fF
C14 clkgen.delay_155ns_2.genblk1\[3\].bypass_enable/X clkgen.delay_155ns_2.genblk1\[1\].bypass_enable/X 1.95fF
C15 VPWR clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit/in 2.08fF
C16 dlycontrol3_in[2] VPWR 4.72fF
C17 clkgen.delay_155ns_3.genblk1\[0\].bypass_enable/B VPWR 1.96fF
C18 edgedetect.dly_315ns_1.enablebuffer/X edgedetect.dly_315ns_1.genblk1\[3\].bypass_enable/X 4.08fF
C19 clk_dig_out dlycontrol1_in[4] 1.15fF
C20 edgedetect.dly_315ns_1.genblk1\[2\].bypass_enable/X clkgen.delay_155ns_3.genblk1\[1\].bypass_enable/B 1.14fF
C21 VPWR edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit/out 2.04fF
C22 dlycontrol4_in[3] clkgen.delay_155ns_3.genblk1\[0\].bypass_enable/X 1.28fF
C23 dlycontrol4_in[3] edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.out_mux/X 1.61fF
C24 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.out_mux/A0 clkgen.delay_155ns_3.genblk1\[2\].bypass_enable/X 1.19fF
C25 edgedetect.dly_315ns_1.genblk1\[4\].bypass_enable/B nsample_p_in 2.06fF
C26 clkgen.delay_155ns_2.genblk1\[4\].bypass_enable/X VGND 4.26fF
C27 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.out_mux/X clkgen.delay_155ns_2.genblk1\[2\].bypass_enable/X 2.94fF
C28 dlycontrol3_in[0] VGND 3.53fF
C29 dlycontrol4_in[2] inbuf_2/X 1.69fF
C30 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.and_bypass_switch/X VPWR 1.42fF
C31 dlycontrol4_in[4] VPWR 3.22fF
C32 dlycontrol4_in[0] VPWR 4.45fF
C33 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.and_bypass_switch/X dlycontrol2_in[4] 1.50fF
C34 VPWR clkgen.delay_155ns_1.genblk1\[3\].dly_binary.out_mux/A0 1.33fF
C35 edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.and_bypass_switch/X VPWR 1.90fF
C36 edgedetect.dly_315ns_1.genblk1\[1\].bypass_enable/X clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit/in 1.42fF
C37 VPWR edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit/in 1.16fF
C38 sample_p_in VGND 3.15fF
C39 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.out_mux/X VPWR 1.45fF
C40 enable_dlycontrol_in dlycontrol1_in[0] 1.27fF
C41 enable_dlycontrol_in clkgen.delay_155ns_1.genblk1\[2\].bypass_enable/X 3.80fF
C42 VPWR outbuf_1/A 5.73fF
C43 edgedetect.or1/A inbuf_1/X 2.08fF
C44 dlycontrol4_in[0] clkgen.delay_155ns_3.enablebuffer/X 2.68fF
C45 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.out_mux/A0 clk_dig_out 1.31fF
C46 VPWR clkgen.delay_155ns_3.genblk1\[3\].dly_binary.and_bypass_switch/X 1.15fF
C47 dlycontrol3_in[0] dlycontrol2_in[3] 1.93fF
C48 inbuf_1/X ndecision_finish_in 1.70fF
C49 clkgen.delay_155ns_1.genblk1\[2\].bypass_enable/X clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit/in 1.68fF
C50 VPWR clkgen.delay_155ns_2.genblk1\[2\].bypass_enable/X 5.29fF
C51 dlycontrol3_in[2] clkgen.delay_155ns_1.genblk1\[2\].bypass_enable/X 1.40fF
C52 dlycontrol1_in[3] dlycontrol1_in[4] 1.19fF
C53 clkgen.delay_155ns_1.genblk1\[0\].bypass_enable/X VPWR 4.31fF
C54 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.out_mux/X VPWR 1.72fF
C55 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit/in VPWR 1.04fF
C56 dlycontrol2_in[4] VGND 1.69fF
C57 clkgen.delay_155ns_2.genblk1\[0\].bypass_enable/B clkgen.delay_155ns_2.genblk1\[3\].bypass_enable/X 1.60fF
C58 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.out_mux/X dlycontrol3_in[0] 2.12fF
C59 dlycontrol2_in[2] clkgen.delay_155ns_2.genblk1\[4\].dly_binary.out_mux/A0 5.05fF
C60 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.out_mux/A0 VGND 2.03fF
C61 clkgen.delay_155ns_3.genblk1\[3\].bypass_enable/X VPWR 1.81fF
C62 dlycontrol2_in[0] VGND 3.95fF
C63 clkgen.delay_155ns_1.genblk1\[2\].dly_binary.out_mux/A0 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.and_bypass_switch/X 1.79fF
C64 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit/in VPWR 1.06fF
C65 clkgen.delay_155ns_3.genblk1\[1\].bypass_enable/X VGND 1.85fF
C66 ena_in clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit/in 1.11fF
C67 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.out_mux/A0 VPWR 1.65fF
C68 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.and_bypass_switch/X clkgen.delay_155ns_2.genblk1\[3\].bypass_enable/X 1.45fF
C69 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.out_mux/A0 dlycontrol4_in[2] 6.26fF
C70 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit/in dlycontrol4_in[1] 1.01fF
C71 clkgen.delay_155ns_3.genblk1\[2\].bypass_enable/B VGND 1.74fF
C72 dlycontrol3_in[4] VGND 4.04fF
C73 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.out_mux/A0 clkgen.delay_155ns_2.genblk1\[0\].bypass_enable/X 2.08fF
C74 ena_in clkgen.delay_155ns_1.genblk1\[3\].bypass_enable/X 1.93fF
C75 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.and_bypass_switch/X clkgen.delay_155ns_3.genblk1\[1\].bypass_enable/B 3.28fF
C76 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.out_mux/A0 VGND 1.96fF
C77 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.out_mux/A0 start_conv_in 2.67fF
C78 VPWR clkgen.delay_155ns_1.genblk1\[1\].bypass_enable/B 1.31fF
C79 clkgen.delay_155ns_2.genblk1\[4\].bypass_enable/X VPWR 4.99fF
C80 VGND inbuf_2/X 6.36fF
C81 dlycontrol3_in[0] VPWR 5.05fF
C82 edgedetect.dly_315ns_1.genblk1\[1\].bypass_enable/X inbuf_2/X 2.29fF
C83 dlycontrol2_in[1] clkgen.delay_155ns_3.genblk1\[4\].bypass_enable/X 1.26fF
C84 VPWR clk_comp_out 1.36fF
C85 clkgen.clkdig_inverter/A VGND 7.11fF
C86 clkgen.delay_155ns_1.genblk1\[2\].dly_binary.out_mux/X clkgen.delay_155ns_3.genblk1\[2\].bypass_enable/B 5.54fF
C87 VPWR clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit/in 1.06fF
C88 clkgen.delay_155ns_2.genblk1\[3\].bypass_enable/X VGND 4.11fF
C89 dlycontrol1_in[0] clkgen.delay_155ns_1.genblk1\[1\].dly_binary.out_mux/A0 1.90fF
C90 dlycontrol2_in[3] clkgen.delay_155ns_3.genblk1\[2\].bypass_enable/B 1.42fF
C91 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit/in VPWR 1.02fF
C92 clkgen.delay_155ns_1.genblk1\[0\].bypass_enable/X clkgen.delay_155ns_1.genblk1\[2\].bypass_enable/X 1.19fF
C93 sample_p_in VPWR 2.12fF
C94 clkgen.delay_155ns_3.genblk1\[1\].bypass_enable/X dlycontrol4_in[1] 2.41fF
C95 VGND clk_dig_out 1.28fF
C96 clkgen.delay_155ns_3.genblk1\[2\].bypass_enable/B dlycontrol4_in[1] 1.25fF
C97 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[23\].delay_unit/in VPWR 1.04fF
C98 VGND edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[20\].delay_unit/in 1.83fF
C99 VPWR clkgen.delay_155ns_3.genblk1\[2\].dly_binary.out_mux/X 1.12fF
C100 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[30\].delay_unit/in VPWR 1.05fF
C101 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit/in VPWR 1.06fF
C102 clkgen.delay_155ns_3.genblk1\[4\].bypass_enable/B VPWR 1.01fF
C103 edgedetect.nor1/A VGND 2.11fF
C104 ena_in clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit/in 2.85fF
C105 dlycontrol4_in[0] edgedetect.dly_315ns_1.genblk1\[5\].bypass_enable/X 2.48fF
C106 inbuf_3/X VPWR 1.42fF
C107 dlycontrol2_in[4] VPWR 2.91fF
C108 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.out_mux/A0 VPWR 1.16fF
C109 dlycontrol1_in[2] VGND 1.54fF
C110 dlycontrol2_in[0] VPWR 3.65fF
C111 clkgen.nor1/A dlycontrol2_in[2] 1.22fF
C112 clkgen.delay_155ns_3.genblk1\[1\].bypass_enable/X VPWR 2.72fF
C113 clkgen.delay_155ns_2.genblk1\[0\].bypass_enable/X VGND 6.45fF
C114 clkgen.delay_155ns_3.genblk1\[2\].bypass_enable/B sample_n_in 2.44fF
C115 dlycontrol3_in[0] dlycontrol1_in[0] 1.72fF
C116 clkgen.delay_155ns_2.genblk1\[1\].bypass_enable/B VGND 1.35fF
C117 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.out_mux/A0 VGND 4.50fF
C118 clkgen.delay_155ns_3.genblk1\[2\].bypass_enable/B VPWR 2.87fF
C119 dlycontrol3_in[4] VPWR 3.86fF
C120 dlycontrol4_in[4] edgedetect.dly_315ns_1.genblk1\[3\].bypass_enable/X 6.74fF
C121 start_conv_in VGND 7.29fF
C122 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.out_mux/A0 dlycontrol1_in[4] 5.00fF
C123 VGND dlycontrol1_in[3] 3.01fF
C124 edgedetect.dly_315ns_1.genblk1\[0\].bypass_enable/X inbuf_2/X 3.48fF
C125 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.out_mux/A0 VPWR 1.76fF
C126 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.out_mux/A0 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.out_mux/X 1.95fF
C127 VPWR inbuf_2/X 7.11fF
C128 dlycontrol2_in[3] clkgen.delay_155ns_2.genblk1\[0\].bypass_enable/X 1.74fF
C129 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit/in VPWR 1.31fF
C130 clkgen.clkdig_inverter/A VPWR 1.33fF
C131 nsample_p_out edgedetect.dly_315ns_1.genblk1\[3\].bypass_enable/X 4.74fF
C132 VGND clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit/in 1.81fF
C133 VPWR clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit/in 1.14fF
C134 clkgen.delay_155ns_2.genblk1\[0\].dly_binary.out_mux/X edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.and_bypass_switch/X 1.05fF
C135 clkgen.delay_155ns_2.genblk1\[3\].bypass_enable/X VPWR 6.52fF
C136 edgedetect.dly_315ns_1.genblk1\[2\].bypass_enable/B nsample_p_out 1.92fF
C137 clkgen.delay_155ns_2.genblk1\[0\].dly_binary.and_bypass_switch/X clkgen.delay_155ns_1.genblk1\[4\].dly_binary.and_bypass_switch/X 1.46fF
C138 VPWR clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit/in 1.10fF
C139 clkgen.delay_155ns_2.genblk1\[2\].bypass_enable/X edgedetect.dly_315ns_1.genblk1\[3\].bypass_enable/X 2.09fF
C140 ena_in clkgen.delay_155ns_1.genblk1\[0\].bypass_enable/X 1.07fF
C141 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.out_mux/X clkgen.delay_155ns_2.genblk1\[0\].bypass_enable/X 4.04fF
C142 VPWR clk_dig_out 2.43fF
C143 dlycontrol2_in[3] dlycontrol1_in[3] 1.32fF
C144 clkgen.delay_155ns_3.enablebuffer/X inbuf_2/X 1.68fF
C145 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.out_mux/A0 dlycontrol4_in[1] 3.66fF
C146 edgedetect.nor1/A edgedetect.dly_315ns_1.genblk1\[0\].bypass_enable/X 3.21fF
C147 clkgen.clkdig_inverter/A nsample_n_in 1.11fF
C148 VPWR edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[20\].delay_unit/in 2.64fF
C149 VGND clkgen.delay_155ns_3.genblk1\[2\].bypass_enable/X 1.99fF
C150 edgedetect.nor1/A VPWR 3.51fF
C151 clkgen.delay_155ns_2.genblk1\[4\].bypass_enable/X ndecision_finish_in 6.88fF
C152 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.and_bypass_switch/X VPWR 1.10fF
C153 clkgen.delay_155ns_2.genblk1\[4\].bypass_enable/X clkgen.delay_155ns_3.genblk1\[0\].bypass_enable/X 1.10fF
C154 clkgen.delay_155ns_2.genblk1\[4\].bypass_enable/X dlycontrol2_in[1] 1.03fF
C155 dlycontrol1_in[2] VPWR 2.59fF
C156 VGND clkgen.delay_155ns_3.genblk1\[4\].dly_binary.out_mux/A0 2.74fF
C157 clkgen.delay_155ns_2.genblk1\[0\].bypass_enable/X VPWR 6.27fF
C158 clkgen.delay_155ns_2.genblk1\[1\].bypass_enable/X VGND 4.49fF
C159 clkgen.delay_155ns_2.genblk1\[1\].bypass_enable/B VPWR 1.60fF
C160 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.out_mux/A0 VPWR 6.53fF
C161 VPWR edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit/in 1.01fF
C162 VGND edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit/in 1.81fF
C163 VGND dlycontrol1_in[4] 2.60fF
C164 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.out_mux/A0 clkgen.delay_155ns_2.genblk1\[2\].bypass_enable/X 1.76fF
C165 clkgen.delay_155ns_1.genblk1\[3\].bypass_enable/X dlycontrol1_in[1] 1.78fF
C166 start_conv_in VPWR 7.70fF
C167 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit/in dlycontrol1_in[3] 1.11fF
C168 VPWR dlycontrol1_in[3] 4.84fF
C169 VPWR edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[21\].delay_unit/in 1.46fF
C170 clkgen.delay_155ns_3.genblk1\[2\].bypass_enable/X dlycontrol4_in[1] 1.12fF
C171 dlycontrol3_in[4] dlycontrol2_in[2] 2.03fF
C172 enable_dlycontrol_in clkgen.delay_155ns_1.genblk1\[4\].bypass_enable/X 3.03fF
C173 clkgen.delay_155ns_2.genblk1\[1\].dly_binary.out_mux/X VPWR 1.41fF
C174 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit/in clkgen.delay_155ns_2.genblk1\[1\].bypass_enable/X 1.03fF
C175 edgedetect.dly_315ns_1.genblk1\[3\].bypass_enable/B clkgen.delay_155ns_2.genblk1\[4\].dly_binary.out_mux/A0 2.20fF
C176 dlycontrol2_in[0] dlycontrol2_in[1] 3.42fF
C177 VPWR clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit/in 1.19fF
C178 clkgen.delay_155ns_3.genblk1\[1\].bypass_enable/X clkgen.delay_155ns_3.genblk1\[0\].bypass_enable/X 1.27fF
C179 dlycontrol4_in[2] VGND 3.67fF
C180 dlycontrol4_in[4] nsample_p_in 4.38fF
C181 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.out_mux/A0 VPWR 2.28fF
C182 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.out_mux/X edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.out_mux/A0 1.17fF
C183 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.out_mux/A0 VGND 2.44fF
C184 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit/in VPWR 1.35fF
C185 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.out_mux/X dlycontrol1_in[4] 2.23fF
C186 clkgen.delay_155ns_2.genblk1\[0\].dly_binary.out_mux/X clkgen.delay_155ns_2.genblk1\[1\].dly_binary.and_bypass_switch/X 1.17fF
C187 enable_dlycontrol_in dlycontrol1_in[1] 1.06fF
C188 dlycontrol1_in[0] clkgen.delay_155ns_2.genblk1\[0\].bypass_enable/X 1.08fF
C189 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.out_mux/A0 edgedetect.dly_315ns_1.genblk1\[5\].bypass_enable/X 1.13fF
C190 VPWR clkgen.delay_155ns_3.genblk1\[2\].bypass_enable/X 2.67fF
C191 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[27\].delay_unit/in VPWR 2.50fF
C192 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit/in clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit/in 1.01fF
C193 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.and_bypass_switch/X clkgen.delay_155ns_1.genblk1\[1\].dly_binary.out_mux/A0 1.81fF
C194 VPWR clkgen.delay_155ns_3.genblk1\[4\].dly_binary.out_mux/A0 2.26fF
C195 clkgen.delay_155ns_2.genblk1\[1\].bypass_enable/X sample_n_in 3.82fF
C196 ndecision_finish_in clkgen.delay_155ns_2.genblk1\[3\].bypass_enable/X 1.27fF
C197 VPWR clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit/in 1.08fF
C198 clkgen.delay_155ns_2.genblk1\[1\].bypass_enable/X VPWR 8.03fF
C199 clkgen.delay_155ns_1.genblk1\[4\].bypass_enable/X outbuf_1/A 1.43fF
C200 dlycontrol4_in[2] dlycontrol4_in[1] 2.82fF
C201 VPWR edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit/in 2.39fF
C202 VPWR dlycontrol1_in[4] 2.69fF
C203 edgedetect.dly_315ns_1.genblk1\[1\].bypass_enable/B VGND 1.43fF
C204 dlycontrol4_in[5] edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit/in 1.28fF
C205 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.out_mux/X clkgen.delay_155ns_1.genblk1\[4\].dly_binary.out_mux/A0 1.94fF
C206 ena_in clk_dig_out 2.14fF
C207 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[6\].delay_unit/in VPWR 1.21fF
C208 clkgen.delay_155ns_1.genblk1\[3\].bypass_enable/X clkgen.delay_155ns_1.genblk1\[3\].dly_binary.out_mux/A0 2.70fF
C209 dlycontrol4_in[5] VGND 1.88fF
C210 enable_dlycontrol_in dlycontrol3_in[2] 1.90fF
C211 dlycontrol3_in[0] clkgen.delay_155ns_1.genblk1\[4\].dly_binary.and_bypass_switch/X 3.39fF
C212 clkgen.delay_155ns_1.genblk1\[3\].bypass_enable/X outbuf_1/A 1.73fF
C213 dlycontrol4_in[2] VPWR 4.16fF
C214 edgedetect.dly_315ns_1.genblk1\[1\].bypass_enable/X VGND 5.55fF
C215 clkgen.delay_155ns_1.genblk1\[1\].bypass_enable/X VGND 2.45fF
C216 clkgen.delay_155ns_2.genblk1\[0\].dly_binary.and_bypass_switch/X clkgen.delay_155ns_2.genblk1\[2\].bypass_enable/X 1.28fF
C217 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.out_mux/A0 VPWR 3.69fF
C218 edgedetect.dly_315ns_1.genblk1\[4\].bypass_enable/X sample_p_in 2.62fF
C219 edgedetect.dly_315ns_1.genblk1\[5\].bypass_enable/B VPWR 1.32fF
C220 ena_in clkgen.delay_155ns_2.genblk1\[0\].bypass_enable/X 1.02fF
C221 dlycontrol2_in[1] start_conv_in 1.67fF
C222 clkgen.delay_155ns_1.genblk1\[0\].bypass_enable/X clkgen.delay_155ns_1.genblk1\[3\].bypass_enable/X 4.07fF
C223 dlycontrol2_in[1] dlycontrol1_in[3] 3.43fF
C224 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit/in VPWR 1.05fF
C225 dlycontrol2_in[3] VGND 2.48fF
C226 ena_in start_conv_in 2.09fF
C227 VPWR clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit/in 1.13fF
C228 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[29\].delay_unit/in VGND 1.30fF
C229 VGND clkgen.delay_155ns_3.genblk1\[0\].dly_binary.out_mux/X 1.19fF
C230 clkgen.delay_155ns_3.genblk1\[2\].bypass_enable/X dlycontrol2_in[2] 1.30fF
C231 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.out_mux/X VGND 3.31fF
C232 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.and_bypass_switch/X VPWR 2.80fF
C233 VGND dlycontrol4_in[1] 3.37fF
C234 dlycontrol4_in[4] edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit/out 1.18fF
C235 dlycontrol3_in[0] dlycontrol1_in[1] 1.47fF
C236 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.out_mux/A0 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit/in 1.71fF
C237 edgedetect.dly_315ns_1.genblk1\[4\].bypass_enable/X clkgen.delay_155ns_3.genblk1\[2\].bypass_enable/B 1.97fF
C238 dlycontrol3_in[0] clkgen.delay_155ns_2.genblk1\[0\].dly_binary.and_bypass_switch/X 2.52fF
C239 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit/in VPWR 2.16fF
C240 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.and_bypass_switch/X dlycontrol3_in[4] 1.37fF
C241 dlycontrol3_in[1] dlycontrol4_in[2] 1.77fF
C242 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.out_mux/X outbuf_1/A 1.29fF
C243 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit/in VGND 1.22fF
C244 edgedetect.dly_315ns_1.genblk1\[0\].bypass_enable/X VGND 2.17fF
C245 clkgen.delay_155ns_2.genblk1\[4\].bypass_enable/X clkgen.delay_155ns_2.genblk1\[4\].dly_binary.out_mux/A0 1.73fF
C246 VGND sample_n_in 2.93fF
C247 dlycontrol4_in[5] VPWR 3.73fF
C248 clkgen.delay_155ns_1.genblk1\[1\].bypass_enable/X sample_n_in 1.16fF
C249 dlycontrol2_in[0] clkgen.delay_155ns_1.genblk1\[4\].bypass_enable/X 1.94fF
C250 VGND VPWR 95.42fF
C251 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.out_mux/X VGND 2.58fF
C252 edgedetect.dly_315ns_1.genblk1\[1\].bypass_enable/X VPWR 7.52fF
C253 clkgen.delay_155ns_1.genblk1\[1\].bypass_enable/X VPWR 3.47fF
C254 dlycontrol4_in[3] inbuf_2/X 2.78fF
C255 dlycontrol2_in[0] inbuf_1/X 1.80fF
C256 VPWR clkgen.delay_155ns_3.genblk1\[1\].dly_binary.out_mux/X 1.04fF
C257 clkgen.delay_155ns_1.genblk1\[0\].bypass_enable/X clkgen.delay_155ns_1.genblk1\[3\].dly_binary.out_mux/A0 2.42fF
C258 clkgen.delay_155ns_3.enablebuffer/X VGND 5.01fF
C259 edgedetect.dly_315ns_1.genblk1\[1\].bypass_enable/X clkgen.delay_155ns_3.enablebuffer/X 1.16fF
C260 ena_in dlycontrol1_in[4] 3.02fF
C261 dlycontrol2_in[3] sample_n_in 2.45fF
C262 outbuf_1/A clkgen.delay_155ns_2.genblk1\[2\].bypass_enable/X 2.96fF
C263 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit/in VGND 1.29fF
C264 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit/in VPWR 1.09fF
C265 dlycontrol2_in[3] VPWR 3.28fF
C266 dlycontrol3_in[0] dlycontrol3_in[2] 1.16fF
C267 clkgen.delay_155ns_1.genblk1\[4\].bypass_enable/X clkgen.delay_155ns_2.genblk1\[3\].bypass_enable/X 2.15fF
C268 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit/in clkgen.delay_155ns_1.genblk1\[0\].dly_binary.and_bypass_switch/X 1.13fF
C269 dlycontrol2_in[4] clkgen.delay_155ns_2.genblk1\[4\].dly_binary.out_mux/A0 5.39fF
C270 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[29\].delay_unit/in VPWR 1.28fF
C271 VPWR clkgen.delay_155ns_3.genblk1\[0\].dly_binary.out_mux/X 1.01fF
C272 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.out_mux/A0 outbuf_1/A 1.21fF
C273 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.out_mux/X VPWR 4.72fF
C274 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit/in VPWR 1.11fF
C275 VPWR dlycontrol4_in[1] 4.60fF
C276 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit/in VPWR 1.02fF
C277 clkgen.clkdig_inverter/A dlycontrol1_in[1] 1.87fF
C278 dlycontrol1_in[0] VGND 3.62fF
C279 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[22\].delay_unit/in VPWR 1.53fF
C280 clkgen.delay_155ns_1.genblk1\[2\].bypass_enable/X VGND 3.38fF
C281 clkgen.delay_155ns_1.genblk1\[1\].bypass_enable/X clkgen.delay_155ns_1.genblk1\[2\].bypass_enable/X 3.19fF
C282 dlycontrol3_in[1] VGND 5.76fF
C283 dlycontrol4_in[5] edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit/in 1.63fF
C284 clkgen.delay_155ns_3.enablebuffer/X dlycontrol4_in[1] 1.21fF
C285 edgedetect.dly_315ns_1.genblk1\[0\].bypass_enable/X VPWR 3.07fF
C286 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit/in VGND 1.27fF
C287 clkgen.delay_155ns_1.genblk1\[2\].dly_binary.out_mux/A0 dlycontrol1_in[4] 2.00fF
C288 VPWR sample_n_in 2.28fF
C289 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit/in VPWR 1.16fF
C290 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.out_mux/X VPWR 4.00fF
C291 dlycontrol2_in[3] dlycontrol1_in[0] 1.47fF
C292 edgedetect.dly_315ns_1.genblk1\[2\].bypass_enable/X VGND 2.28fF
C293 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[24\].delay_unit/in VPWR 1.04fF
C294 dlycontrol3_in[0] clkgen.delay_155ns_2.genblk1\[2\].bypass_enable/X 3.60fF
C295 edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.out_mux/X edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit/in 5.34fF
C296 edgedetect.dly_315ns_1.genblk1\[4\].bypass_enable/X edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.out_mux/A0 1.43fF
C297 edgedetect.dly_315ns_1.genblk1\[0\].bypass_enable/X clkgen.delay_155ns_3.enablebuffer/X 1.98fF
C298 clkgen.delay_155ns_2.genblk1\[2\].bypass_enable/X clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit/in 1.38fF
C299 dlycontrol1_in[2] dlycontrol1_in[1] 5.54fF
C300 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.out_mux/X dlycontrol1_in[0] 1.68fF
C301 clkgen.delay_155ns_3.enablebuffer/X VPWR 5.52fF
C302 VGND dlycontrol2_in[2] 3.92fF
C303 VGND dlycontrol3_in[3] 3.32fF
C304 clkgen.delay_155ns_2.genblk1\[1\].dly_binary.and_bypass_switch/X VGND 1.19fF
C305 inbuf_1/X start_conv_in 1.48fF
C306 edgedetect.or1/A VGND 2.66fF
C307 clkgen.delay_155ns_3.genblk1\[1\].bypass_enable/X edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.and_bypass_switch/X 1.82fF
C308 edgedetect.dly_315ns_1.genblk1\[5\].bypass_enable/X VGND 1.61fF
C309 clkgen.delay_155ns_3.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit/in VPWR 1.10fF
C310 ndecision_finish_in VGND 3.67fF
C311 clkgen.nor1/A inbuf_3/X 1.21fF
C312 VGND clkgen.delay_155ns_3.genblk1\[0\].bypass_enable/X 3.22fF
C313 VPWR clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit/in 1.33fF
C314 dlycontrol2_in[0] outbuf_1/A 2.98fF
C315 dlycontrol2_in[1] VGND 2.90fF
C316 edgedetect.dly_315ns_1.genblk1\[1\].bypass_enable/X clkgen.delay_155ns_3.genblk1\[0\].bypass_enable/X 1.62fF
C317 edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.out_mux/X VGND 2.56fF
C318 clkgen.delay_155ns_1.genblk1\[3\].bypass_enable/X start_conv_in 2.07fF
C319 clkgen.delay_155ns_1.genblk1\[0\].bypass_enable/X inbuf_3/X 1.11fF
C320 dlycontrol1_in[0] VPWR 4.44fF
C321 clkgen.delay_155ns_1.genblk1\[2\].bypass_enable/X VPWR 6.03fF
C322 dlycontrol2_in[0] clkgen.delay_155ns_2.genblk1\[2\].bypass_enable/X 1.39fF
C323 ena_in VGND 2.46fF
C324 dlycontrol3_in[1] VPWR 7.34fF
C325 dlycontrol4_in[5] edgedetect.dly_315ns_1.genblk1\[2\].bypass_enable/B 2.62fF
C326 VGND edgedetect.dly_315ns_1.genblk1\[3\].bypass_enable/X 3.04fF
C327 clkgen.delay_155ns_2.genblk1\[1\].bypass_enable/X clkgen.delay_155ns_2.enablebuffer/X 1.04fF
C328 edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.out_mux/X edgedetect.dly_315ns_1.genblk1\[3\].bypass_enable/X 1.09fF
C329 dlycontrol4_in[5] edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.and_bypass_switch/X 1.13fF
C330 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit/in VPWR 1.15fF
C331 clkgen.delay_155ns_3.genblk1\[0\].dly_binary.out_mux/X dlycontrol3_in[3] 1.23fF
C332 edgedetect.dly_315ns_1.enablebuffer/X dlycontrol4_in[2] 1.13fF
C333 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit/in VPWR 3.48fF
C334 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.and_bypass_switch/X VGND 1.69fF
C335 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.and_bypass_switch/X VGND 1.51fF
C336 clkgen.delay_155ns_3.genblk1\[4\].bypass_enable/X dlycontrol1_in[3] 1.28fF
C337 clkgen.delay_155ns_1.genblk1\[4\].bypass_enable/X clkgen.delay_155ns_2.genblk1\[1\].bypass_enable/X 3.18fF
C338 edgedetect.dly_315ns_1.genblk1\[2\].bypass_enable/X VPWR 3.02fF
C339 edgedetect.dly_315ns_1.genblk1\[2\].bypass_enable/X edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.out_mux/X 1.93fF
C340 VPWR edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit/in 1.16fF
C341 edgedetect.dly_315ns_1.genblk1\[4\].bypass_enable/X dlycontrol4_in[2] 1.63fF
C342 dlycontrol1_in[0] clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit/in 2.33fF
C343 edgedetect.nor1/A edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.and_bypass_switch/X 1.51fF
C344 clkgen.delay_155ns_2.genblk1\[4\].bypass_enable/X clkgen.delay_155ns_3.genblk1\[3\].dly_binary.out_mux/A0 1.33fF
C345 edgedetect.dly_315ns_1.genblk1\[0\].bypass_enable/X dlycontrol3_in[3] 2.63fF
C346 VPWR dlycontrol2_in[2] 3.67fF
C347 outbuf_2/A clkgen.delay_155ns_3.genblk1\[4\].dly_binary.out_mux/A0 3.90fF
C348 clkgen.delay_155ns_1.genblk1\[2\].dly_binary.out_mux/A0 VGND 1.08fF
C349 VGND nsample_n_out 2.26fF
C350 VPWR dlycontrol3_in[3] 2.46fF
C351 dlycontrol4_in[3] edgedetect.dly_315ns_1.genblk1\[5\].bypass_enable/B 1.14fF
C352 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.out_mux/A0 VGND 1.79fF
C353 clkgen.delay_155ns_2.genblk1\[1\].dly_binary.and_bypass_switch/X VPWR 1.18fF
C354 clkgen.delay_155ns_2.genblk1\[4\].bypass_enable/X dlycontrol3_in[4] 2.48fF
C355 clkgen.delay_155ns_1.genblk1\[0\].bypass_enable/X clk_dig_out 1.30fF
C356 clkgen.delay_155ns_2.genblk1\[3\].bypass_enable/B VPWR 1.25fF
C357 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.out_mux/X dlycontrol1_in[3] 1.74fF
C358 edgedetect.dly_315ns_1.genblk1\[0\].bypass_enable/X clkgen.delay_155ns_3.genblk1\[0\].bypass_enable/X 1.98fF
C359 edgedetect.or1/A VPWR 2.54fF
C360 edgedetect.dly_315ns_1.genblk1\[5\].bypass_enable/X VPWR 3.88fF
C361 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[18\].delay_unit/in VPWR 1.14fF
C362 ndecision_finish_in VPWR 5.62fF
C363 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit/in VPWR 1.02fF
C364 VPWR clkgen.delay_155ns_3.genblk1\[0\].bypass_enable/X 2.23fF
C365 dlycontrol2_in[1] VPWR 4.87fF
C366 edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.out_mux/X VPWR 1.24fF
C367 clkgen.delay_155ns_3.enablebuffer/X dlycontrol3_in[3] 1.11fF
C368 clkgen.delay_155ns_2.genblk1\[4\].bypass_enable/X inbuf_2/X 1.35fF
C369 ena_in VPWR 3.46fF
C370 clkgen.delay_155ns_2.genblk1\[4\].bypass_enable/X clkgen.delay_155ns_2.genblk1\[3\].bypass_enable/X 1.31fF
C371 VPWR edgedetect.dly_315ns_1.genblk1\[3\].bypass_enable/X 3.67fF
C372 outbuf_1/A dlycontrol1_in[3] 1.32fF
C373 dlycontrol4_in[5] edgedetect.dly_315ns_1.enablebuffer/X 1.07fF
C374 edgedetect.dly_315ns_1.genblk1\[2\].bypass_enable/B VPWR 1.07fF
C375 clkgen.delay_155ns_3.enablebuffer/X edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.out_mux/X 1.19fF
C376 clkgen.delay_155ns_3.genblk1\[0\].bypass_enable/B clkgen.delay_155ns_3.genblk1\[2\].bypass_enable/X 1.02fF
C377 edgedetect.dly_315ns_1.enablebuffer/X VGND 5.84fF
C378 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.and_bypass_switch/X VPWR 3.61fF
C379 edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.out_mux/X edgedetect.dly_315ns_1.enablebuffer/X 1.21fF
C380 enable_dlycontrol_in clkgen.delay_155ns_2.genblk1\[1\].bypass_enable/X 4.61fF
C381 clkgen.delay_155ns_1.genblk1\[0\].bypass_enable/X start_conv_in 1.59fF
C382 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.out_mux/A0 clkgen.delay_155ns_1.genblk1\[3\].bypass_enable/X 1.23fF
C383 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.and_bypass_switch/X VPWR 2.36fF
C384 dlycontrol4_in[5] nsample_p_in 2.09fF
C385 edgedetect.dly_315ns_1.genblk1\[4\].bypass_enable/X VGND 4.42fF
C386 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit/in VPWR 2.32fF
C387 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.and_bypass_switch/X VGND 1.86fF
C388 dlycontrol3_in[1] edgedetect.dly_315ns_1.genblk1\[5\].bypass_enable/X 1.02fF
C389 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[27\].delay_unit/in dlycontrol4_in[4] 1.33fF
C390 dlycontrol4_in[3] VGND 4.64fF
C391 edgedetect.dly_315ns_1.genblk1\[1\].bypass_enable/X dlycontrol4_in[3] 1.94fF
C392 VGND clkgen.delay_155ns_2.enablebuffer/X 1.38fF
C393 clkgen.delay_155ns_2.genblk1\[3\].bypass_enable/X dlycontrol2_in[4] 1.15fF
C394 clkgen.delay_155ns_1.genblk1\[2\].dly_binary.out_mux/A0 VPWR 1.03fF
C395 clkgen.delay_155ns_1.genblk1\[2\].bypass_enable/B clkgen.delay_155ns_1.genblk1\[3\].bypass_enable/X 1.10fF
C396 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.out_mux/A0 VPWR 2.36fF
C397 ena_in dlycontrol1_in[0] 1.24fF
C398 edgedetect.dly_315ns_1.enablebuffer/X clkgen.delay_155ns_3.genblk1\[0\].dly_binary.out_mux/X 1.84fF
C399 dlycontrol2_in[0] clkgen.delay_155ns_2.genblk1\[3\].bypass_enable/X 2.81fF
C400 clkgen.delay_155ns_1.genblk1\[0\].bypass_enable/X clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit/in 1.13fF
C401 edgedetect.dly_315ns_1.enablebuffer/X dlycontrol4_in[1] 2.41fF
C402 clkgen.delay_155ns_1.genblk1\[4\].bypass_enable/X VGND 6.02fF
C403 clkgen.delay_155ns_3.genblk1\[1\].bypass_enable/B VGND 1.81fF
C404 edgedetect.dly_315ns_1.genblk1\[2\].bypass_enable/X edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.out_mux/X 2.59fF
C405 clkgen.delay_155ns_3.genblk1\[0\].bypass_enable/B dlycontrol4_in[2] 3.75fF
C406 nsample_n_in nsample_n_out 1.63fF
C407 inbuf_1/X VGND 1.93fF
C408 dlycontrol3_in[1] edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.and_bypass_switch/X 1.22fF
C409 VGND dlycontrol1_in[1] 1.24fF
C410 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit/in VPWR 1.13fF
C411 ndecision_finish_in dlycontrol2_in[2] 1.04fF
C412 clkgen.delay_155ns_2.genblk1\[1\].bypass_enable/X clkgen.delay_155ns_2.genblk1\[2\].bypass_enable/X 1.02fF
C413 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[15\].delay_unit/in VPWR 1.16fF
C414 edgedetect.dly_315ns_1.genblk1\[3\].bypass_enable/X edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit/in 5.35fF
C415 clkgen.delay_155ns_2.genblk1\[0\].dly_binary.and_bypass_switch/X VGND 1.39fF
C416 VGND outbuf_2/A 2.93fF
C417 edgedetect.dly_315ns_1.genblk1\[3\].bypass_enable/B VGND 1.21fF
C418 edgedetect.dly_315ns_1.enablebuffer/X VPWR 8.29fF
C419 clkgen.delay_155ns_1.enablebuffer/X VGND 1.20fF
C420 clkgen.delay_155ns_1.genblk1\[0\].bypass_enable/X dlycontrol1_in[4] 1.30fF
C421 clkgen.delay_155ns_1.genblk1\[3\].bypass_enable/X VGND 3.34fF
C422 edgedetect.or1/A dlycontrol2_in[1] 1.68fF
C423 edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.out_mux/X edgedetect.dly_315ns_1.genblk1\[5\].bypass_enable/X 1.14fF
C424 clkgen.delay_155ns_3.genblk1\[1\].bypass_enable/X edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.out_mux/A0 3.01fF
C425 dlycontrol1_in[2] clkgen.delay_155ns_3.genblk1\[2\].bypass_enable/B 3.46fF
C426 ndecision_finish_in dlycontrol2_in[1] 1.90fF
C427 clkgen.delay_155ns_1.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit/in VPWR 1.20fF
C428 clkgen.delay_155ns_3.genblk1\[0\].dly_binary.and_bypass_switch/X VPWR 1.30fF
C429 edgedetect.nor1/A inbuf_2/X 1.07fF
C430 edgedetect.dly_315ns_1.genblk1\[4\].bypass_enable/X VPWR 9.19fF
C431 edgedetect.dly_315ns_1.genblk1\[4\].bypass_enable/X edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.out_mux/X 1.61fF
C432 VGND clkgen.delay_155ns_2.genblk1\[4\].dly_binary.out_mux/A0 5.61fF
C433 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.and_bypass_switch/X VPWR 2.68fF
C434 dlycontrol2_in[0] start_conv_in 1.02fF
C435 VPWR nsample_p_in 1.17fF
C436 dlycontrol2_in[0] dlycontrol1_in[3] 2.69fF
C437 dlycontrol4_in[3] VPWR 6.06fF
C438 VGND clkgen.delay_155ns_2.genblk1\[2\].bypass_enable/B 1.29fF
C439 VPWR clkgen.delay_155ns_2.enablebuffer/X 1.22fF
C440 dlycontrol1_in[2] clkgen.clkdig_inverter/A 3.79fF
C441 clkgen.delay_155ns_3.genblk1\[4\].bypass_enable/X VGND 1.19fF
C442 clkgen.delay_155ns_1.genblk1\[2\].bypass_enable/B clkgen.delay_155ns_1.genblk1\[3\].bypass_enable/B 1.15fF
C443 enable_dlycontrol_in VGND 5.10fF
C444 enable_dlycontrol_in clkgen.delay_155ns_1.genblk1\[1\].bypass_enable/X 1.04fF
C445 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.out_mux/X clkgen.delay_155ns_2.genblk1\[0\].dly_binary.and_bypass_switch/X 2.42fF
C446 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.and_bypass_switch/X edgedetect.dly_315ns_1.genblk1\[5\].bypass_enable/X 1.64fF
C447 clkgen.delay_155ns_1.genblk1\[4\].bypass_enable/X VPWR 5.52fF
C448 VGND clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit/in 1.37fF
C449 dlycontrol3_in[2] VGND 3.82fF
C450 dlycontrol3_in[2] clkgen.delay_155ns_1.genblk1\[1\].bypass_enable/X 7.93fF
C451 clkgen.delay_155ns_3.genblk1\[0\].bypass_enable/B VGND 2.44fF
C452 clkgen.delay_155ns_3.genblk1\[1\].bypass_enable/B VPWR 2.46fF
C453 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit/in VPWR 1.15fF
C454 clkgen.delay_155ns_2.genblk1\[3\].bypass_enable/X start_conv_in 1.51fF
C455 dlycontrol1_in[1] sample_n_in 3.53fF
C456 VPWR edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit/in 1.21fF
C457 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.out_mux/X VGND 1.25fF
C458 clkgen.delay_155ns_1.genblk1\[2\].dly_binary.and_bypass_switch/X VPWR 1.42fF
C459 inbuf_1/X VPWR 3.42fF
C460 start_conv_in clk_dig_out 4.55fF
C461 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit/in VPWR 1.02fF
C462 VPWR dlycontrol1_in[1] 2.74fF
C463 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.out_mux/A0 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.out_mux/A0 2.58fF
C464 dlycontrol4_in[5] dlycontrol4_in[4] 7.83fF
C465 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.and_bypass_switch/X dlycontrol1_in[0] 2.31fF
C466 clkgen.clkdig_inverter/A clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit/in 1.19fF
C467 clkgen.delay_155ns_1.genblk1\[3\].bypass_enable/X sample_n_in 1.25fF
C468 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.and_bypass_switch/X VGND 1.82fF
C469 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit/in VPWR 1.09fF
C470 clkgen.delay_155ns_2.genblk1\[0\].dly_binary.and_bypass_switch/X VPWR 2.96fF
C471 VPWR outbuf_2/A 3.48fF
C472 dlycontrol4_in[4] VGND 1.06fF
C473 dlycontrol4_in[0] VGND 3.41fF
C474 edgedetect.dly_315ns_1.genblk1\[3\].bypass_enable/B VPWR 1.84fF
C475 clkgen.delay_155ns_1.enablebuffer/X VPWR 1.77fF
C476 clkgen.delay_155ns_1.genblk1\[3\].bypass_enable/B VGND 2.83fF
C477 edgedetect.dly_315ns_1.genblk1\[1\].bypass_enable/X dlycontrol4_in[0] 9.40fF
C478 clkgen.delay_155ns_1.genblk1\[3\].bypass_enable/X VPWR 3.47fF
C479 clkgen.delay_155ns_1.genblk1\[3\].bypass_enable/B clkgen.delay_155ns_1.genblk1\[1\].bypass_enable/X 1.24fF
C480 VGND clkgen.delay_155ns_1.genblk1\[3\].dly_binary.out_mux/A0 1.85fF
C481 edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.and_bypass_switch/X VGND 2.33fF
C482 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit/in 0 1.32fF
C483 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit/in 0 1.12fF
C484 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit/in 0 1.22fF
C485 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit/in 0 1.04fF
C486 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit/in 0 1.37fF
C487 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit/out 0 1.08fF
C488 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit/in 0 1.28fF
C489 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit/in 0 1.00fF
C490 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit/in 0 1.03fF
C491 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit/in 0 1.07fF
C492 edgedetect.dly_315ns_1.genblk1\[3\].bypass_enable/X 0 1.85fF
C493 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit/in 0 1.05fF
C494 nsample_p_in 0 1.04fF
C495 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.out_mux/A0 0 3.87fF
C496 edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit/in 0 1.02fF
C497 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[26\].delay_unit/in 0 1.13fF
C498 dlycontrol1_in[1] 0 1.08fF
C499 VPWR 0 571.41fF
C500 VGND 0 54.47fF
C501 start_conv_in 0 1.80fF
C502 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.and_bypass_switch/X 0 1.23fF
C503 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.out_mux/A0 0 2.11fF
C504 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit/in 0 1.36fF
C505 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit/in 0 1.19fF
C506 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit/in 0 1.08fF
C507 edgedetect.dly_315ns_1.enablebuffer/X 0 -2.35fF
C508 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit/in 0 1.01fF
C509 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit/in 0 1.09fF
C510 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit/in 0 1.35fF
C511 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit/in 0 1.15fF
C512 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit/in 0 1.08fF
C513 clkgen.delay_155ns_1.genblk1\[2\].dly_binary.out_mux/X 0 1.48fF
C514 ena_in 0 1.08fF
C515 edgedetect.dly_315ns_1.genblk1\[0\].bypass_enable/X 0 1.06fF
C516 dlycontrol2_in[0] 0 1.76fF
C517 clkgen.clkdig_inverter/A 0 1.33fF
C518 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit/in 0 1.01fF
C519 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[27\].delay_unit/in 0 1.14fF
C520 dlycontrol1_in[2] 0 1.03fF
C521 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit/in 0 1.25fF
C522 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit/in 0 1.41fF
C523 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit/in 0 1.23fF
.ends

