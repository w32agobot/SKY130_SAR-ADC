magic
tech sky130A
timestamp 1664895328
<< nwell >>
rect 0 253 502 440
<< nmos >>
rect 116 126 131 168
rect 164 126 179 168
rect 308 127 323 169
rect 356 127 371 169
<< pmos >>
rect 116 271 131 351
rect 164 271 179 351
rect 308 272 323 352
rect 356 272 371 352
<< ndiff >>
rect 85 162 116 168
rect 85 132 91 162
rect 108 132 116 162
rect 85 126 116 132
rect 131 162 164 168
rect 131 132 139 162
rect 156 132 164 162
rect 131 126 164 132
rect 179 162 210 168
rect 179 132 187 162
rect 204 132 210 162
rect 179 126 210 132
rect 277 163 308 169
rect 277 133 283 163
rect 300 133 308 163
rect 277 127 308 133
rect 323 163 356 169
rect 323 133 331 163
rect 348 133 356 163
rect 323 127 356 133
rect 371 163 402 169
rect 371 133 379 163
rect 396 133 402 163
rect 371 127 402 133
<< pdiff >>
rect 85 345 116 351
rect 85 277 91 345
rect 108 277 116 345
rect 85 271 116 277
rect 131 345 164 351
rect 131 277 139 345
rect 156 277 164 345
rect 131 271 164 277
rect 179 345 210 351
rect 179 277 187 345
rect 204 277 210 345
rect 179 271 210 277
rect 277 346 308 352
rect 277 278 283 346
rect 300 278 308 346
rect 277 272 308 278
rect 323 346 356 352
rect 323 278 331 346
rect 348 278 356 346
rect 323 272 356 278
rect 371 346 402 352
rect 371 278 379 346
rect 396 278 402 346
rect 371 272 402 278
<< ndiffc >>
rect 91 132 108 162
rect 139 132 156 162
rect 187 132 204 162
rect 283 133 300 163
rect 331 133 348 163
rect 379 133 396 163
<< pdiffc >>
rect 91 277 108 345
rect 139 277 156 345
rect 187 277 204 345
rect 283 278 300 346
rect 331 278 348 346
rect 379 278 396 346
<< psubdiff >>
rect 91 74 115 91
rect 132 74 163 91
rect 180 74 215 91
rect 232 74 267 91
rect 284 74 314 91
rect 331 74 363 91
rect 380 74 396 91
<< nsubdiff >>
rect 151 419 403 422
rect 151 402 163 419
rect 180 402 215 419
rect 232 402 267 419
rect 284 402 315 419
rect 332 402 362 419
rect 379 402 403 419
rect 151 399 403 402
<< psubdiffcont >>
rect 115 74 132 91
rect 163 74 180 91
rect 215 74 232 91
rect 267 74 284 91
rect 314 74 331 91
rect 363 74 380 91
<< nsubdiffcont >>
rect 163 402 180 419
rect 215 402 232 419
rect 267 402 284 419
rect 315 402 332 419
rect 362 402 379 419
<< poly >>
rect 106 409 140 414
rect 106 391 114 409
rect 132 391 140 409
rect 106 374 140 391
rect 106 359 179 374
rect 116 351 131 359
rect 164 351 179 359
rect 308 352 323 365
rect 356 352 371 365
rect 116 168 131 271
rect 164 168 179 271
rect 308 215 323 272
rect 205 214 323 215
rect 356 214 371 272
rect 205 209 371 214
rect 205 192 213 209
rect 230 200 371 209
rect 230 192 249 200
rect 205 187 249 192
rect 308 187 371 200
rect 308 169 323 187
rect 356 169 371 187
rect 116 113 131 126
rect 164 113 179 126
rect 308 114 323 127
rect 356 114 371 127
rect 417 110 444 118
rect 417 93 422 110
rect 439 93 444 110
rect 417 85 444 93
<< polycont >>
rect 114 391 132 409
rect 213 192 230 209
rect 422 93 439 110
<< locali >>
rect 17 461 74 502
rect 427 474 485 502
rect 17 444 24 461
rect 68 444 74 461
rect 17 353 74 444
rect 420 461 485 474
rect 420 444 428 461
rect 477 444 485 461
rect 151 419 403 422
rect 114 409 132 417
rect 151 402 163 419
rect 180 402 215 419
rect 232 402 267 419
rect 284 402 315 419
rect 332 402 362 419
rect 379 402 403 419
rect 151 399 403 402
rect 114 386 132 391
rect 114 369 115 386
rect 17 336 23 353
rect 64 336 74 353
rect 17 304 74 336
rect 17 287 23 304
rect 64 287 74 304
rect 17 133 74 287
rect 91 345 108 353
rect 91 269 108 277
rect 139 345 156 353
rect 17 116 57 133
rect 17 51 74 116
rect 91 162 108 170
rect 91 91 108 132
rect 139 164 156 277
rect 187 345 204 399
rect 187 269 204 277
rect 283 346 300 399
rect 283 270 300 278
rect 331 346 348 354
rect 178 209 238 210
rect 178 204 213 209
rect 197 192 213 204
rect 230 192 238 209
rect 197 187 238 192
rect 139 124 156 132
rect 187 162 204 170
rect 187 91 204 132
rect 283 163 300 171
rect 283 91 300 133
rect 331 163 348 278
rect 379 346 396 399
rect 379 270 396 278
rect 420 353 485 444
rect 420 336 429 353
rect 478 336 485 353
rect 420 304 485 336
rect 420 287 429 304
rect 478 287 485 304
rect 331 125 348 133
rect 379 163 396 171
rect 379 91 396 133
rect 91 74 115 91
rect 132 74 163 91
rect 180 74 215 91
rect 232 74 267 91
rect 284 74 314 91
rect 331 74 363 91
rect 380 74 396 91
rect 420 170 485 287
rect 420 141 429 170
rect 478 141 485 170
rect 420 110 485 141
rect 420 93 422 110
rect 439 93 485 110
rect 17 34 23 51
rect 68 34 74 51
rect 17 0 74 34
rect 420 51 485 93
rect 420 34 429 51
rect 478 34 485 51
rect 420 30 485 34
rect 427 0 485 30
<< viali >>
rect 24 444 68 461
rect 428 444 477 461
rect 163 402 180 419
rect 215 402 232 419
rect 267 402 284 419
rect 315 402 332 419
rect 362 402 379 419
rect 115 369 132 386
rect 23 336 64 353
rect 23 287 64 304
rect 91 298 108 321
rect 57 116 74 133
rect 187 300 204 323
rect 331 300 348 335
rect 178 187 197 204
rect 139 162 156 164
rect 139 144 156 162
rect 429 336 478 353
rect 429 287 478 304
rect 115 74 132 91
rect 163 74 180 91
rect 215 74 232 91
rect 267 74 284 91
rect 314 74 331 91
rect 363 74 380 91
rect 429 141 478 170
rect 23 34 68 51
rect 429 34 478 51
<< metal1 >>
rect 17 461 74 502
rect 427 474 485 502
rect 17 444 24 461
rect 68 444 74 461
rect 17 441 74 444
rect 420 461 485 474
rect 420 444 428 461
rect 477 444 485 461
rect 420 441 485 444
rect 0 419 502 427
rect 0 403 163 419
rect 0 399 98 403
rect 149 402 163 403
rect 180 402 215 419
rect 232 402 267 419
rect 284 402 315 419
rect 332 402 362 419
rect 379 402 502 419
rect 149 399 502 402
rect 109 386 138 389
rect 109 385 115 386
rect 0 370 115 385
rect 109 369 115 370
rect 132 369 138 386
rect 109 366 138 369
rect 331 370 502 385
rect 17 353 70 356
rect 17 336 23 353
rect 64 336 70 353
rect 331 342 348 370
rect 420 353 485 356
rect 17 304 70 336
rect 327 335 351 342
rect 17 287 23 304
rect 64 287 70 304
rect 85 323 210 327
rect 85 321 187 323
rect 85 298 91 321
rect 108 300 187 321
rect 204 300 210 323
rect 108 298 210 300
rect 85 295 210 298
rect 327 300 331 335
rect 348 300 351 335
rect 327 287 351 300
rect 420 336 429 353
rect 478 336 485 353
rect 420 304 485 336
rect 420 287 429 304
rect 478 287 485 304
rect 17 284 70 287
rect 420 284 485 287
rect 0 256 502 270
rect 78 229 421 242
rect 0 228 502 229
rect 0 215 97 228
rect 404 215 502 228
rect 172 204 203 208
rect 172 201 178 204
rect 0 187 178 201
rect 197 187 203 204
rect 172 182 203 187
rect 244 187 502 201
rect 135 164 159 172
rect 54 142 83 145
rect 54 124 57 142
rect 135 144 139 164
rect 156 156 159 164
rect 244 156 259 187
rect 156 144 259 156
rect 135 140 259 144
rect 420 170 485 173
rect 420 141 429 170
rect 478 141 485 170
rect 135 138 159 140
rect 420 138 485 141
rect 0 116 57 124
rect 83 116 502 124
rect 0 110 502 116
rect 0 91 502 96
rect 0 74 115 91
rect 132 74 163 91
rect 180 74 215 91
rect 232 74 267 91
rect 284 74 314 91
rect 331 74 363 91
rect 380 74 502 91
rect 0 68 502 74
rect 17 51 74 54
rect 17 34 23 51
rect 68 34 74 51
rect 17 0 74 34
rect 420 51 485 54
rect 420 34 429 51
rect 478 34 485 51
rect 420 30 485 34
rect 427 0 485 30
<< via1 >>
rect 57 133 83 142
rect 57 116 74 133
rect 74 116 83 133
<< metal2 >>
rect 16 481 486 486
rect 16 453 21 481
rect 49 453 69 481
rect 97 453 117 481
rect 145 453 165 481
rect 193 453 213 481
rect 241 453 261 481
rect 289 453 309 481
rect 337 453 357 481
rect 385 453 405 481
rect 433 453 453 481
rect 481 453 486 481
rect 16 433 486 453
rect 16 405 21 433
rect 49 405 165 433
rect 193 405 309 433
rect 337 405 453 433
rect 481 405 486 433
rect 16 385 486 405
rect 16 357 21 385
rect 49 357 165 385
rect 193 357 309 385
rect 337 357 453 385
rect 481 357 486 385
rect 16 337 486 357
rect 16 309 21 337
rect 49 309 69 337
rect 97 309 117 337
rect 145 309 165 337
rect 193 309 213 337
rect 241 309 261 337
rect 289 309 309 337
rect 337 309 357 337
rect 385 309 405 337
rect 433 309 453 337
rect 481 309 486 337
rect 16 304 486 309
rect 16 289 198 304
rect 16 261 21 289
rect 49 261 165 289
rect 193 261 198 289
rect 304 289 486 304
rect 16 241 198 261
rect 16 213 21 241
rect 49 213 165 241
rect 193 213 198 241
rect 230 230 272 272
rect 304 261 309 289
rect 337 261 453 289
rect 481 261 486 289
rect 304 241 486 261
rect 16 198 198 213
rect 304 213 309 241
rect 337 213 453 241
rect 481 213 486 241
rect 304 198 486 213
rect 16 193 486 198
rect 16 165 21 193
rect 49 165 69 193
rect 97 165 117 193
rect 145 165 165 193
rect 193 165 213 193
rect 241 165 261 193
rect 289 165 309 193
rect 337 165 357 193
rect 385 165 405 193
rect 433 165 453 193
rect 481 165 486 193
rect 16 145 486 165
rect 16 117 21 145
rect 49 142 165 145
rect 49 117 57 142
rect 16 116 57 117
rect 83 117 165 142
rect 193 117 309 145
rect 337 117 453 145
rect 481 117 486 145
rect 83 116 486 117
rect 16 97 486 116
rect 16 69 21 97
rect 49 69 165 97
rect 193 69 309 97
rect 337 69 453 97
rect 481 69 486 97
rect 16 49 486 69
rect 16 21 21 49
rect 49 21 69 49
rect 97 21 117 49
rect 145 21 165 49
rect 193 21 213 49
rect 241 21 261 49
rect 289 21 309 49
rect 337 21 357 49
rect 385 21 405 49
rect 433 21 453 49
rect 481 21 486 49
rect 16 16 486 21
<< via2 >>
rect 21 453 49 481
rect 69 453 97 481
rect 117 453 145 481
rect 165 453 193 481
rect 213 453 241 481
rect 261 453 289 481
rect 309 453 337 481
rect 357 453 385 481
rect 405 453 433 481
rect 453 453 481 481
rect 21 405 49 433
rect 165 405 193 433
rect 309 405 337 433
rect 453 405 481 433
rect 21 357 49 385
rect 165 357 193 385
rect 309 357 337 385
rect 453 357 481 385
rect 21 309 49 337
rect 69 309 97 337
rect 117 309 145 337
rect 165 309 193 337
rect 213 309 241 337
rect 261 309 289 337
rect 309 309 337 337
rect 357 309 385 337
rect 405 309 433 337
rect 453 309 481 337
rect 21 261 49 289
rect 165 261 193 289
rect 21 213 49 241
rect 165 213 193 241
rect 309 261 337 289
rect 453 261 481 289
rect 309 213 337 241
rect 453 213 481 241
rect 21 165 49 193
rect 69 165 97 193
rect 117 165 145 193
rect 165 165 193 193
rect 213 165 241 193
rect 261 165 289 193
rect 309 165 337 193
rect 357 165 385 193
rect 405 165 433 193
rect 453 165 481 193
rect 21 117 49 145
rect 165 117 193 145
rect 309 117 337 145
rect 453 117 481 145
rect 21 69 49 97
rect 165 69 193 97
rect 309 69 337 97
rect 453 69 481 97
rect 21 21 49 49
rect 69 21 97 49
rect 117 21 145 49
rect 165 21 193 49
rect 213 21 241 49
rect 261 21 289 49
rect 309 21 337 49
rect 357 21 385 49
rect 405 21 433 49
rect 453 21 481 49
<< metal3 >>
rect 18 481 484 484
rect 18 453 21 481
rect 49 453 69 481
rect 97 453 117 481
rect 145 453 165 481
rect 193 453 213 481
rect 241 453 261 481
rect 289 453 309 481
rect 337 453 357 481
rect 385 453 405 481
rect 433 453 453 481
rect 481 453 484 481
rect 18 450 484 453
rect 18 433 52 450
rect 18 405 21 433
rect 49 405 52 433
rect 162 433 196 450
rect 18 385 52 405
rect 18 357 21 385
rect 49 357 52 385
rect 82 412 132 420
rect 82 378 90 412
rect 124 378 132 412
rect 82 370 132 378
rect 162 405 165 433
rect 193 405 196 433
rect 306 433 340 450
rect 162 385 196 405
rect 18 340 52 357
rect 162 357 165 385
rect 193 357 196 385
rect 226 412 276 420
rect 226 378 234 412
rect 268 378 276 412
rect 226 370 276 378
rect 306 405 309 433
rect 337 405 340 433
rect 450 433 484 450
rect 306 385 340 405
rect 162 340 196 357
rect 306 357 309 385
rect 337 357 340 385
rect 370 412 420 420
rect 370 378 378 412
rect 412 378 420 412
rect 370 370 420 378
rect 450 405 453 433
rect 481 405 484 433
rect 450 385 484 405
rect 306 340 340 357
rect 450 357 453 385
rect 481 357 484 385
rect 450 340 484 357
rect 18 337 484 340
rect 18 309 21 337
rect 49 309 69 337
rect 97 309 117 337
rect 145 309 165 337
rect 193 309 213 337
rect 241 309 261 337
rect 289 309 309 337
rect 337 309 357 337
rect 385 309 405 337
rect 433 309 453 337
rect 481 309 484 337
rect 18 306 484 309
rect 18 289 52 306
rect 18 261 21 289
rect 49 261 52 289
rect 162 289 196 306
rect 18 241 52 261
rect 18 213 21 241
rect 49 213 52 241
rect 82 268 132 276
rect 82 234 90 268
rect 124 234 132 268
rect 82 226 132 234
rect 162 261 165 289
rect 193 261 196 289
rect 162 241 196 261
rect 18 196 52 213
rect 162 213 165 241
rect 193 213 196 241
rect 162 196 196 213
rect 306 289 340 306
rect 306 261 309 289
rect 337 261 340 289
rect 450 289 484 306
rect 306 241 340 261
rect 306 213 309 241
rect 337 213 340 241
rect 370 268 420 276
rect 370 234 378 268
rect 412 234 420 268
rect 370 226 420 234
rect 450 261 453 289
rect 481 261 484 289
rect 450 241 484 261
rect 306 196 340 213
rect 450 213 453 241
rect 481 213 484 241
rect 450 196 484 213
rect 18 193 484 196
rect 18 165 21 193
rect 49 165 69 193
rect 97 165 117 193
rect 145 165 165 193
rect 193 165 213 193
rect 241 165 261 193
rect 289 165 309 193
rect 337 165 357 193
rect 385 165 405 193
rect 433 165 453 193
rect 481 165 484 193
rect 18 162 484 165
rect 18 145 52 162
rect 18 117 21 145
rect 49 117 52 145
rect 162 145 196 162
rect 18 97 52 117
rect 18 69 21 97
rect 49 69 52 97
rect 82 124 132 132
rect 82 90 90 124
rect 124 90 132 124
rect 82 82 132 90
rect 162 117 165 145
rect 193 117 196 145
rect 306 145 340 162
rect 162 97 196 117
rect 18 52 52 69
rect 162 69 165 97
rect 193 69 196 97
rect 226 124 276 132
rect 226 90 234 124
rect 268 90 276 124
rect 226 82 276 90
rect 306 117 309 145
rect 337 117 340 145
rect 450 145 484 162
rect 306 97 340 117
rect 162 52 196 69
rect 306 69 309 97
rect 337 69 340 97
rect 370 124 420 132
rect 370 90 378 124
rect 412 90 420 124
rect 370 82 420 90
rect 450 117 453 145
rect 481 117 484 145
rect 450 97 484 117
rect 306 52 340 69
rect 450 69 453 97
rect 481 69 484 97
rect 450 52 484 69
rect 18 49 484 52
rect 18 21 21 49
rect 49 21 69 49
rect 97 21 117 49
rect 145 21 165 49
rect 193 21 213 49
rect 241 21 261 49
rect 289 21 309 49
rect 337 21 357 49
rect 385 21 405 49
rect 433 21 453 49
rect 481 21 484 49
rect 18 18 484 21
<< via3 >>
rect 90 378 124 412
rect 234 378 268 412
rect 378 378 412 412
rect 90 234 124 268
rect 378 234 412 268
rect 90 90 124 124
rect 234 90 268 124
rect 378 90 412 124
<< metal4 >>
rect 92 420 122 467
rect 236 420 266 467
rect 380 420 410 467
rect 82 412 132 420
rect 82 410 90 412
rect 35 380 90 410
rect 82 378 90 380
rect 124 410 132 412
rect 226 412 276 420
rect 226 410 234 412
rect 124 380 234 410
rect 124 378 132 380
rect 82 370 132 378
rect 226 378 234 380
rect 268 410 276 412
rect 370 412 420 420
rect 370 410 378 412
rect 268 380 378 410
rect 268 378 276 380
rect 226 370 276 378
rect 370 378 378 380
rect 412 410 420 412
rect 412 380 467 410
rect 412 378 420 380
rect 370 370 420 378
rect 92 276 122 370
rect 236 323 266 370
rect 380 276 410 370
rect 82 268 132 276
rect 82 266 90 268
rect 35 236 90 266
rect 82 234 90 236
rect 124 266 132 268
rect 370 268 420 276
rect 370 266 378 268
rect 124 236 179 266
rect 323 236 378 266
rect 124 234 132 236
rect 82 226 132 234
rect 370 234 378 236
rect 412 266 420 268
rect 412 236 467 266
rect 412 234 420 236
rect 370 226 420 234
rect 92 132 122 226
rect 236 132 266 179
rect 380 132 410 226
rect 82 124 132 132
rect 82 122 90 124
rect 35 92 90 122
rect 82 90 90 92
rect 124 122 132 124
rect 226 124 276 132
rect 226 122 234 124
rect 124 92 234 122
rect 124 90 132 92
rect 82 82 132 90
rect 226 90 234 92
rect 268 122 276 124
rect 370 124 420 132
rect 370 122 378 124
rect 268 92 378 122
rect 268 90 276 92
rect 226 82 276 90
rect 370 90 378 92
rect 412 122 420 124
rect 412 92 467 122
rect 412 90 420 92
rect 370 82 420 90
rect 92 35 122 82
rect 236 35 266 82
rect 380 35 410 82
<< comment >>
rect 0 486 16 502
rect 486 486 502 502
rect 69 375 154 399
rect 215 378 281 402
rect 69 130 97 375
rect 156 345 184 375
rect 179 214 203 344
rect 215 281 239 378
rect 282 358 303 381
rect 299 304 316 358
rect 288 302 316 304
rect 279 301 316 302
rect 279 288 304 301
rect 272 281 300 288
rect 215 279 300 281
rect 215 272 288 279
rect 215 257 279 272
rect 215 230 239 257
rect 280 239 301 261
rect 280 238 318 239
rect 214 214 239 230
rect 179 198 214 214
rect 150 130 178 159
rect 179 157 203 198
rect 69 129 178 130
rect 69 106 153 129
rect 215 103 239 214
rect 301 99 318 238
rect 335 99 358 401
rect 0 0 16 16
rect 486 0 502 16
<< labels >>
rlabel metal1 0 399 0 427 7 VDD
port 2 w
rlabel metal1 0 256 0 270 7 colon_n
port 3 w
rlabel metal1 0 215 0 229 7 col_n
port 4 w
rlabel metal1 0 110 0 124 7 vcom
port 5 w
rlabel metal1 0 68 0 96 7 VSS
port 6 w
rlabel locali 427 0 485 0 5 row_n
port 7 s
rlabel metal4 92 467 122 467 1 ctop
port 1 n
rlabel metal1 0 187 0 201 7 sample_i
port 12 w
rlabel metal1 0 370 0 385 7 sample_n_i
port 13 w
rlabel metal1 502 370 502 385 3 sample_n_o
port 14 e
rlabel metal1 502 187 502 201 3 sample_o
port 15 e
<< end >>
