* NGSPICE file created from adc_array_circuit.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_01v8_J7MSU8 a_n111_n68# a_n81_n42# a_15_n42# a_n15_n68#
+ a_n173_n42# a_81_n68# a_111_n42# VSUBS
X0 a_15_n42# a_n15_n68# a_n81_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1 a_111_n42# a_81_n68# a_15_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X2 a_n81_n42# a_n111_n68# a_n173_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_MJPTSJ a_63_n42# a_n125_n42# a_n63_n68# a_33_n68#
+ a_n33_n42# VSUBS
X0 a_63_n42# a_33_n68# a_n33_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=1.302e+11p pd=1.46e+06u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1 a_n33_n42# a_n63_n68# a_n125_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_5CE3MA a_111_n80# a_81_n106# a_n15_n106# a_n111_n106#
+ a_n81_n80# a_15_n80# w_n209_n116# a_n173_n80#
X0 a_n81_n80# a_n111_n106# a_n173_n80# w_n209_n116# sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=2.48e+11p ps=2.22e+06u w=800000u l=150000u
X1 a_111_n80# a_81_n106# a_15_n80# w_n209_n116# sky130_fd_pr__pfet_01v8 ad=2.48e+11p pd=2.22e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2 a_15_n80# a_n15_n106# a_n81_n80# w_n209_n116# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_5CSGFE w_n161_n116# a_33_n106# a_63_n80# a_n125_n80#
+ a_n63_n106# a_n33_n80#
X0 a_n33_n80# a_n63_n106# a_n125_n80# w_n161_n116# sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=2.48e+11p ps=2.22e+06u w=800000u l=150000u
X1 a_63_n80# a_33_n106# a_n33_n80# w_n161_n116# sky130_fd_pr__pfet_01v8 ad=2.48e+11p pd=2.22e+06u as=0p ps=0u w=800000u l=150000u
.ends

.subckt adc_array_circuit
Xsky130_fd_pr__nfet_01v8_J7MSU8_0 colon_n li_722_732# VSS col_n li_322_734# row_n
+ li_722_732# VSS sky130_fd_pr__nfet_01v8_J7MSU8
Xsky130_fd_pr__nfet_01v8_MJPTSJ_0 vcom li_322_734# sample_n sample li_418_782# VSS
+ sky130_fd_pr__nfet_01v8_MJPTSJ
Xsky130_fd_pr__pfet_01v8_5CE3MA_0 li_322_734# col_n row_n colon_n VDD vint1 VDD li_322_734#
+ sky130_fd_pr__pfet_01v8_5CE3MA
Xsky130_fd_pr__pfet_01v8_5CSGFE_0 VDD sample li_322_734# vcom sample_n li_418_782#
+ sky130_fd_pr__pfet_01v8_5CSGFE
.ends

