magic
tech sky130A
timestamp 1659006126
<< metal2 >>
rect 14 513 518 518
rect 14 485 19 513
rect 47 485 67 513
rect 95 485 115 513
rect 143 485 156 513
rect 184 485 204 513
rect 232 485 252 513
rect 280 485 300 513
rect 328 485 348 513
rect 376 485 389 513
rect 417 485 437 513
rect 465 485 485 513
rect 513 485 518 513
rect 14 465 518 485
rect 14 437 19 465
rect 47 437 252 465
rect 280 437 485 465
rect 513 437 518 465
rect 14 417 518 437
rect 14 389 19 417
rect 47 389 252 417
rect 280 389 485 417
rect 513 389 518 417
rect 14 376 518 389
rect 14 348 19 376
rect 47 348 252 376
rect 280 348 485 376
rect 513 348 518 376
rect 14 328 518 348
rect 14 300 19 328
rect 47 300 252 328
rect 280 300 485 328
rect 513 300 518 328
rect 14 280 518 300
rect 14 252 19 280
rect 47 252 67 280
rect 95 252 115 280
rect 143 252 156 280
rect 184 252 204 280
rect 232 252 252 280
rect 280 252 300 280
rect 328 252 348 280
rect 376 252 389 280
rect 417 252 437 280
rect 465 252 485 280
rect 513 252 518 280
rect 14 232 518 252
rect 14 204 19 232
rect 47 204 252 232
rect 280 204 485 232
rect 513 204 518 232
rect 14 184 518 204
rect 14 156 19 184
rect 47 156 252 184
rect 280 156 485 184
rect 513 156 518 184
rect 14 143 518 156
rect 14 115 19 143
rect 47 115 252 143
rect 280 115 485 143
rect 513 115 518 143
rect 14 95 518 115
rect 14 67 19 95
rect 47 67 252 95
rect 280 67 485 95
rect 513 67 518 95
rect 14 47 518 67
rect 14 19 19 47
rect 47 19 67 47
rect 95 19 115 47
rect 143 19 156 47
rect 184 19 204 47
rect 232 19 252 47
rect 280 19 300 47
rect 328 19 348 47
rect 376 19 389 47
rect 417 19 437 47
rect 465 19 485 47
rect 513 19 518 47
rect 14 14 518 19
<< via2 >>
rect 19 485 47 513
rect 67 485 95 513
rect 115 485 143 513
rect 156 485 184 513
rect 204 485 232 513
rect 252 485 280 513
rect 300 485 328 513
rect 348 485 376 513
rect 389 485 417 513
rect 437 485 465 513
rect 485 485 513 513
rect 19 437 47 465
rect 252 437 280 465
rect 485 437 513 465
rect 19 389 47 417
rect 252 389 280 417
rect 485 389 513 417
rect 19 348 47 376
rect 252 348 280 376
rect 485 348 513 376
rect 19 300 47 328
rect 252 300 280 328
rect 485 300 513 328
rect 19 252 47 280
rect 67 252 95 280
rect 115 252 143 280
rect 156 252 184 280
rect 204 252 232 280
rect 252 252 280 280
rect 300 252 328 280
rect 348 252 376 280
rect 389 252 417 280
rect 437 252 465 280
rect 485 252 513 280
rect 19 204 47 232
rect 252 204 280 232
rect 485 204 513 232
rect 19 156 47 184
rect 252 156 280 184
rect 485 156 513 184
rect 19 115 47 143
rect 252 115 280 143
rect 485 115 513 143
rect 19 67 47 95
rect 252 67 280 95
rect 485 67 513 95
rect 19 19 47 47
rect 67 19 95 47
rect 115 19 143 47
rect 156 19 184 47
rect 204 19 232 47
rect 252 19 280 47
rect 300 19 328 47
rect 348 19 376 47
rect 389 19 417 47
rect 437 19 465 47
rect 485 19 513 47
<< metal3 >>
rect 16 513 516 516
rect 16 485 19 513
rect 47 485 67 513
rect 95 485 115 513
rect 143 485 156 513
rect 184 485 204 513
rect 232 485 252 513
rect 280 485 300 513
rect 328 485 348 513
rect 376 485 389 513
rect 417 485 437 513
rect 465 485 485 513
rect 513 485 516 513
rect 16 482 516 485
rect 16 465 50 482
rect 16 437 19 465
rect 47 437 50 465
rect 249 465 283 482
rect 16 417 50 437
rect 16 389 19 417
rect 47 389 50 417
rect 80 444 130 452
rect 80 410 88 444
rect 122 410 130 444
rect 80 402 130 410
rect 169 444 219 452
rect 169 410 177 444
rect 211 410 219 444
rect 169 402 219 410
rect 249 437 252 465
rect 280 437 283 465
rect 482 465 516 482
rect 249 417 283 437
rect 16 376 50 389
rect 16 348 19 376
rect 47 348 50 376
rect 249 389 252 417
rect 280 389 283 417
rect 313 444 363 452
rect 313 410 321 444
rect 355 410 363 444
rect 313 402 363 410
rect 402 444 452 452
rect 402 410 410 444
rect 444 410 452 444
rect 402 402 452 410
rect 482 437 485 465
rect 513 437 516 465
rect 482 417 516 437
rect 249 376 283 389
rect 16 328 50 348
rect 16 300 19 328
rect 47 300 50 328
rect 80 355 130 363
rect 80 321 88 355
rect 122 321 130 355
rect 80 313 130 321
rect 169 355 219 363
rect 169 321 177 355
rect 211 321 219 355
rect 169 313 219 321
rect 249 348 252 376
rect 280 348 283 376
rect 482 389 485 417
rect 513 389 516 417
rect 482 376 516 389
rect 249 328 283 348
rect 16 283 50 300
rect 249 300 252 328
rect 280 300 283 328
rect 313 355 363 363
rect 313 321 321 355
rect 355 321 363 355
rect 313 313 363 321
rect 402 355 452 363
rect 402 321 410 355
rect 444 321 452 355
rect 402 313 452 321
rect 482 348 485 376
rect 513 348 516 376
rect 482 328 516 348
rect 249 283 283 300
rect 482 300 485 328
rect 513 300 516 328
rect 482 283 516 300
rect 16 280 516 283
rect 16 252 19 280
rect 47 252 67 280
rect 95 252 115 280
rect 143 252 156 280
rect 184 252 204 280
rect 232 252 252 280
rect 280 252 300 280
rect 328 252 348 280
rect 376 252 389 280
rect 417 252 437 280
rect 465 252 485 280
rect 513 252 516 280
rect 16 249 516 252
rect 16 232 50 249
rect 16 204 19 232
rect 47 204 50 232
rect 249 232 283 249
rect 16 184 50 204
rect 16 156 19 184
rect 47 156 50 184
rect 80 211 130 219
rect 80 177 88 211
rect 122 177 130 211
rect 80 169 130 177
rect 169 211 219 219
rect 169 177 177 211
rect 211 177 219 211
rect 169 169 219 177
rect 249 204 252 232
rect 280 204 283 232
rect 482 232 516 249
rect 249 184 283 204
rect 16 143 50 156
rect 16 115 19 143
rect 47 115 50 143
rect 249 156 252 184
rect 280 156 283 184
rect 313 211 363 219
rect 313 177 321 211
rect 355 177 363 211
rect 313 169 363 177
rect 402 211 452 219
rect 402 177 410 211
rect 444 177 452 211
rect 402 169 452 177
rect 482 204 485 232
rect 513 204 516 232
rect 482 184 516 204
rect 249 143 283 156
rect 16 95 50 115
rect 16 67 19 95
rect 47 67 50 95
rect 80 122 130 130
rect 80 88 88 122
rect 122 88 130 122
rect 80 80 130 88
rect 169 122 219 130
rect 169 88 177 122
rect 211 88 219 122
rect 169 80 219 88
rect 249 115 252 143
rect 280 115 283 143
rect 482 156 485 184
rect 513 156 516 184
rect 482 143 516 156
rect 249 95 283 115
rect 16 50 50 67
rect 249 67 252 95
rect 280 67 283 95
rect 313 122 363 130
rect 313 88 321 122
rect 355 88 363 122
rect 313 80 363 88
rect 402 122 452 130
rect 402 88 410 122
rect 444 88 452 122
rect 402 80 452 88
rect 482 115 485 143
rect 513 115 516 143
rect 482 95 516 115
rect 249 50 283 67
rect 482 67 485 95
rect 513 67 516 95
rect 482 50 516 67
rect 16 47 516 50
rect 16 19 19 47
rect 47 19 67 47
rect 95 19 115 47
rect 143 19 156 47
rect 184 19 204 47
rect 232 19 252 47
rect 280 19 300 47
rect 328 19 348 47
rect 376 19 389 47
rect 417 19 437 47
rect 465 19 485 47
rect 513 19 516 47
rect 16 16 516 19
<< via3 >>
rect 88 410 122 444
rect 177 410 211 444
rect 321 410 355 444
rect 410 410 444 444
rect 88 321 122 355
rect 177 321 211 355
rect 321 321 355 355
rect 410 321 444 355
rect 88 177 122 211
rect 177 177 211 211
rect 321 177 355 211
rect 410 177 444 211
rect 88 88 122 122
rect 177 88 211 122
rect 321 88 355 122
rect 410 88 444 122
<< metal4 >>
rect 90 452 120 532
rect 179 452 209 532
rect 323 452 353 532
rect 412 452 442 532
rect 80 444 130 452
rect 80 442 88 444
rect 0 412 88 442
rect 80 410 88 412
rect 122 442 130 444
rect 169 444 219 452
rect 169 442 177 444
rect 122 412 177 442
rect 122 410 130 412
rect 80 402 130 410
rect 169 410 177 412
rect 211 442 219 444
rect 313 444 363 452
rect 313 442 321 444
rect 211 412 321 442
rect 211 410 219 412
rect 169 402 219 410
rect 313 410 321 412
rect 355 442 363 444
rect 402 444 452 452
rect 402 442 410 444
rect 355 412 410 442
rect 355 410 363 412
rect 313 402 363 410
rect 402 410 410 412
rect 444 442 452 444
rect 444 412 532 442
rect 444 410 452 412
rect 402 402 452 410
rect 90 363 120 402
rect 179 363 209 402
rect 323 363 353 402
rect 412 363 442 402
rect 80 355 130 363
rect 80 353 88 355
rect 0 323 88 353
rect 80 321 88 323
rect 122 353 130 355
rect 169 355 219 363
rect 169 353 177 355
rect 122 323 177 353
rect 122 321 130 323
rect 80 313 130 321
rect 169 321 177 323
rect 211 353 219 355
rect 313 355 363 363
rect 313 353 321 355
rect 211 323 321 353
rect 211 321 219 323
rect 169 313 219 321
rect 313 321 321 323
rect 355 353 363 355
rect 402 355 452 363
rect 402 353 410 355
rect 355 323 410 353
rect 355 321 363 323
rect 313 313 363 321
rect 402 321 410 323
rect 444 353 452 355
rect 444 323 532 353
rect 444 321 452 323
rect 402 313 452 321
rect 90 266 120 313
rect 179 266 209 313
rect 323 266 353 313
rect 412 266 442 313
rect 80 211 130 219
rect 80 209 88 211
rect 0 179 88 209
rect 80 177 88 179
rect 122 209 130 211
rect 169 211 219 219
rect 169 209 177 211
rect 122 179 177 209
rect 122 177 130 179
rect 80 169 130 177
rect 169 177 177 179
rect 211 209 219 211
rect 313 211 363 219
rect 313 209 321 211
rect 211 179 321 209
rect 211 177 219 179
rect 169 169 219 177
rect 313 177 321 179
rect 355 209 363 211
rect 402 211 452 219
rect 402 209 410 211
rect 355 179 410 209
rect 355 177 363 179
rect 313 169 363 177
rect 402 177 410 179
rect 444 209 452 211
rect 444 179 532 209
rect 444 177 452 179
rect 402 169 452 177
rect 90 130 120 169
rect 179 130 209 169
rect 323 130 353 169
rect 412 130 442 169
rect 80 122 130 130
rect 80 120 88 122
rect 0 90 88 120
rect 80 88 88 90
rect 122 120 130 122
rect 169 122 219 130
rect 169 120 177 122
rect 122 90 177 120
rect 122 88 130 90
rect 80 80 130 88
rect 169 88 177 90
rect 211 120 219 122
rect 313 122 363 130
rect 313 120 321 122
rect 211 90 321 120
rect 211 88 219 90
rect 169 80 219 88
rect 313 88 321 90
rect 355 120 363 122
rect 402 122 452 130
rect 402 120 410 122
rect 355 90 410 120
rect 355 88 363 90
rect 313 80 363 88
rect 402 88 410 90
rect 444 120 452 122
rect 444 90 532 120
rect 444 88 452 90
rect 402 80 452 88
rect 90 0 120 80
rect 179 0 209 80
rect 323 0 353 80
rect 412 0 442 80
<< comment >>
rect 0 518 14 532
rect 518 518 532 532
rect 0 0 14 14
rect 518 1 532 15
<< labels >>
rlabel metal2 14 54 14 54 7 cbot
port 2 w
rlabel metal4 0 104 0 105 3 cfloating
rlabel metal4 104 532 104 532 5 ctop
port 3 s
<< end >>
