* NGSPICE file created from delay_macrocell.ext - technology: sky130A

.subckt delay_macrocell in VPWR out VGND VNB VPB
X0 VGND cap_top a_968_80# VNB sky130_fd_pr__nfet_01v8 ad=2.604e+11p pd=2.92e+06u as=5.292e+11p ps=5.88e+06u w=420000u l=150000u
X1 cap_top VGND sky130_fd_pr__cap_mim_m3_1 l=1.93e+06u w=3.68e+06u
X2 cap_top in VGND VNB sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=4e+06u
X3 out cap_top a_968_80# VNB sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4 a_968_80# cap_top VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 cap_top VGND sky130_fd_pr__cap_mim_m3_1 l=1.93e+06u w=3.26e+06u
X6 a_968_80# cap_top out VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 cap_top in VPWR VPB sky130_fd_pr__pfet_01v8 ad=2.32e+11p pd=2.18e+06u as=4.96e+11p ps=4.44e+06u w=800000u l=4e+06u
X8 VPWR out a_968_80# VNB sky130_fd_pr__nfet_01v8 ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X9 VGND out a_968_308# VPB sky130_fd_pr__pfet_01v8 ad=3.52e+11p pd=2.48e+06u as=1.008e+12p ps=8.92e+06u w=800000u l=150000u
X10 VPWR cap_top a_968_308# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11 out cap_top a_968_308# VPB sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12 a_968_308# cap_top VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X13 a_968_308# cap_top out VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
.ends

