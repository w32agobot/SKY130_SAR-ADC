VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO adc_comp_latch
  CLASS BLOCK ;
  FOREIGN adc_comp_latch ;
  ORIGIN 0.000 0.000 ;
  SIZE 42.000 BY 129.000 ;
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 28.380 68.020 36.290 68.040 ;
        RECT 16.590 66.000 36.290 68.020 ;
        RECT 16.590 65.910 28.050 66.000 ;
        RECT 19.220 65.900 20.430 65.910 ;
        RECT 22.260 64.160 28.050 65.910 ;
        RECT 31.240 65.760 36.290 66.000 ;
        RECT 14.230 62.070 16.440 64.060 ;
        RECT 32.040 62.300 34.610 62.560 ;
        RECT 28.560 60.280 34.610 62.300 ;
      LAYER li1 ;
        RECT 28.390 67.650 31.130 68.140 ;
        RECT 31.680 67.690 35.910 67.860 ;
        RECT 15.700 67.190 21.060 67.430 ;
        RECT 23.280 67.240 26.900 67.480 ;
        RECT 15.700 64.060 16.130 67.190 ;
        RECT 16.840 67.100 20.850 67.190 ;
        RECT 16.840 66.390 17.010 67.100 ;
        RECT 17.800 66.390 17.970 67.100 ;
        RECT 18.760 66.390 18.930 67.100 ;
        RECT 19.720 66.390 19.890 67.100 ;
        RECT 20.680 66.390 20.850 67.100 ;
        RECT 24.960 67.070 25.410 67.240 ;
        RECT 24.110 66.900 26.200 67.070 ;
        RECT 24.110 64.640 24.280 66.900 ;
        RECT 25.070 64.640 25.240 66.900 ;
        RECT 26.030 64.640 26.200 66.900 ;
        RECT 29.280 66.290 29.450 67.650 ;
        RECT 30.240 66.290 30.410 67.650 ;
        RECT 14.100 63.860 16.130 64.060 ;
        RECT 14.100 62.940 14.280 63.860 ;
        RECT 14.540 63.700 14.960 63.860 ;
        RECT 15.230 62.940 15.450 63.860 ;
        RECT 15.710 63.700 16.130 63.860 ;
        RECT 14.100 62.750 14.980 62.940 ;
        RECT 15.230 62.750 16.150 62.940 ;
        RECT 29.280 60.650 29.450 62.010 ;
        RECT 30.240 60.650 30.410 62.010 ;
        RECT 30.850 60.650 31.130 67.650 ;
        RECT 32.440 66.250 32.610 67.690 ;
        RECT 34.920 66.250 35.090 67.690 ;
        RECT 28.400 60.630 31.130 60.650 ;
        RECT 33.240 60.630 33.410 62.070 ;
        RECT 28.400 60.460 34.230 60.630 ;
      LAYER mcon ;
        RECT 28.860 67.860 29.040 68.040 ;
        RECT 29.240 67.860 29.420 68.040 ;
        RECT 29.620 67.860 29.800 68.040 ;
        RECT 30.000 67.860 30.180 68.040 ;
        RECT 30.380 67.860 30.560 68.040 ;
        RECT 30.760 67.860 30.940 68.040 ;
        RECT 15.760 67.220 15.930 67.400 ;
        RECT 16.150 67.220 16.320 67.400 ;
        RECT 16.510 67.220 16.680 67.400 ;
        RECT 16.930 67.220 17.100 67.390 ;
        RECT 17.350 67.220 17.520 67.390 ;
        RECT 17.770 67.220 17.940 67.390 ;
        RECT 18.190 67.220 18.360 67.390 ;
        RECT 18.610 67.220 18.780 67.390 ;
        RECT 19.030 67.220 19.200 67.390 ;
        RECT 19.450 67.220 19.620 67.390 ;
        RECT 19.870 67.220 20.040 67.390 ;
        RECT 20.290 67.220 20.460 67.390 ;
        RECT 20.740 67.220 20.910 67.390 ;
        RECT 23.470 67.270 23.640 67.440 ;
        RECT 23.890 67.270 24.060 67.440 ;
        RECT 24.310 67.270 24.480 67.440 ;
        RECT 24.730 67.270 24.900 67.440 ;
        RECT 25.150 67.270 25.320 67.440 ;
        RECT 25.570 67.270 25.740 67.440 ;
        RECT 25.990 67.270 26.160 67.440 ;
        RECT 26.410 67.270 26.580 67.440 ;
        RECT 14.660 63.890 14.840 64.060 ;
        RECT 15.830 63.890 16.010 64.060 ;
      LAYER met1 ;
        RECT 10.000 67.700 39.920 68.850 ;
        RECT 15.700 67.190 21.060 67.700 ;
        RECT 23.280 67.240 26.900 67.700 ;
        RECT 14.500 63.860 14.990 64.090 ;
        RECT 15.670 63.860 16.160 64.090 ;
      LAYER via ;
        RECT 10.320 67.790 11.120 68.740 ;
        RECT 39.020 67.790 39.820 68.740 ;
      LAYER met2 ;
        RECT 10.230 67.700 11.230 68.850 ;
        RECT 38.920 67.700 39.920 68.850 ;
      LAYER via2 ;
        RECT 10.320 67.790 11.120 68.740 ;
        RECT 39.020 67.790 39.820 68.740 ;
      LAYER met3 ;
        RECT 10.230 67.700 11.230 68.850 ;
        RECT 38.920 67.700 39.920 68.850 ;
      LAYER via3 ;
        RECT 10.320 67.790 11.120 68.740 ;
        RECT 39.020 67.790 39.820 68.740 ;
      LAYER met4 ;
        RECT 10.230 50.000 11.230 77.980 ;
        RECT 38.920 50.000 39.920 77.980 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 17.320 75.990 19.720 76.890 ;
        RECT 30.220 75.990 32.620 76.890 ;
        RECT 15.020 75.590 21.270 75.990 ;
        RECT 24.520 75.590 25.420 75.990 ;
        RECT 28.670 75.590 34.920 75.990 ;
        RECT 15.020 70.290 34.920 75.590 ;
        RECT 15.020 69.890 21.270 70.290 ;
        RECT 24.520 69.890 25.420 70.290 ;
        RECT 28.670 69.890 34.920 70.290 ;
        RECT 17.320 68.990 19.720 69.890 ;
        RECT 30.220 68.990 32.620 69.890 ;
        RECT 17.320 58.040 19.720 58.940 ;
        RECT 30.220 58.040 32.620 58.940 ;
        RECT 15.020 57.640 21.270 58.040 ;
        RECT 24.520 57.640 25.420 58.040 ;
        RECT 28.670 57.640 34.920 58.040 ;
        RECT 15.020 52.340 34.920 57.640 ;
        RECT 15.020 51.940 21.270 52.340 ;
        RECT 24.520 51.940 25.420 52.340 ;
        RECT 28.670 51.940 34.920 52.340 ;
        RECT 17.320 51.040 19.720 51.940 ;
        RECT 30.220 51.040 32.620 51.940 ;
      LAYER li1 ;
        RECT 12.940 76.990 37.330 77.980 ;
        RECT 12.940 74.540 14.120 76.990 ;
        RECT 17.370 76.490 19.670 76.990 ;
        RECT 30.270 76.490 32.570 76.990 ;
        RECT 14.520 76.090 35.420 76.490 ;
        RECT 12.940 50.990 13.930 74.540 ;
        RECT 14.520 69.790 14.920 76.090 ;
        RECT 17.370 76.040 19.670 76.090 ;
        RECT 30.270 76.040 32.570 76.090 ;
        RECT 15.720 74.890 34.220 75.490 ;
        RECT 18.320 74.290 18.670 74.890 ;
        RECT 16.070 74.090 18.670 74.290 ;
        RECT 18.320 73.490 18.670 74.090 ;
        RECT 16.070 73.290 18.670 73.490 ;
        RECT 19.270 73.390 19.470 74.890 ;
        RECT 20.070 73.390 20.270 74.890 ;
        RECT 20.870 73.390 21.070 74.890 ;
        RECT 21.670 73.390 21.870 74.890 ;
        RECT 22.470 73.390 22.670 74.890 ;
        RECT 23.270 73.390 23.470 74.890 ;
        RECT 24.070 73.390 24.270 74.890 ;
        RECT 24.870 73.390 25.070 74.890 ;
        RECT 25.670 73.390 25.870 74.890 ;
        RECT 26.470 73.390 26.670 74.890 ;
        RECT 27.270 73.390 27.470 74.890 ;
        RECT 28.070 73.390 28.270 74.890 ;
        RECT 28.870 73.390 29.070 74.890 ;
        RECT 29.670 73.390 29.870 74.890 ;
        RECT 30.470 73.390 30.670 74.890 ;
        RECT 31.270 74.290 31.620 74.890 ;
        RECT 31.270 74.090 33.870 74.290 ;
        RECT 31.270 73.490 31.620 74.090 ;
        RECT 31.270 73.290 33.820 73.490 ;
        RECT 16.070 72.390 18.670 72.590 ;
        RECT 18.320 71.790 18.670 72.390 ;
        RECT 16.070 71.590 18.670 71.790 ;
        RECT 18.320 70.990 18.670 71.590 ;
        RECT 19.270 70.990 19.470 72.490 ;
        RECT 20.070 70.990 20.270 72.490 ;
        RECT 20.870 70.990 21.070 72.490 ;
        RECT 21.670 70.990 21.870 72.490 ;
        RECT 22.470 70.990 22.670 72.490 ;
        RECT 23.270 70.990 23.470 72.490 ;
        RECT 24.070 70.990 24.270 72.490 ;
        RECT 24.870 70.990 25.070 72.490 ;
        RECT 25.670 70.990 25.870 72.490 ;
        RECT 26.470 70.990 26.670 72.490 ;
        RECT 27.270 70.990 27.470 72.490 ;
        RECT 28.070 70.990 28.270 72.490 ;
        RECT 28.870 70.990 29.070 72.490 ;
        RECT 29.670 70.990 29.870 72.490 ;
        RECT 30.470 70.990 30.670 72.490 ;
        RECT 31.270 72.390 33.820 72.590 ;
        RECT 31.270 71.790 31.620 72.390 ;
        RECT 31.270 71.590 33.870 71.790 ;
        RECT 31.270 70.990 31.620 71.590 ;
        RECT 15.720 70.390 34.220 70.990 ;
        RECT 17.370 69.790 19.670 69.840 ;
        RECT 30.270 69.790 32.570 69.840 ;
        RECT 35.020 69.790 35.420 76.090 ;
        RECT 14.520 69.390 35.420 69.790 ;
        RECT 17.370 68.990 19.670 69.390 ;
        RECT 30.270 68.990 32.570 69.390 ;
        RECT 29.280 64.410 29.450 65.200 ;
        RECT 30.240 64.410 30.410 65.200 ;
        RECT 31.960 64.740 32.130 65.440 ;
        RECT 34.440 64.740 34.610 65.440 ;
        RECT 36.340 64.740 37.330 76.990 ;
        RECT 31.830 64.480 37.330 64.740 ;
        RECT 28.740 64.320 30.520 64.410 ;
        RECT 28.060 63.980 30.520 64.320 ;
        RECT 14.520 61.060 14.980 61.230 ;
        RECT 15.690 61.060 16.150 61.230 ;
        RECT 14.540 60.530 14.960 61.060 ;
        RECT 15.710 60.530 16.130 61.060 ;
        RECT 17.320 60.310 17.490 61.570 ;
        RECT 18.280 60.310 18.450 61.560 ;
        RECT 19.240 60.310 19.410 61.560 ;
        RECT 20.200 60.310 20.370 61.560 ;
        RECT 24.110 60.450 24.280 63.030 ;
        RECT 25.070 60.450 25.240 63.030 ;
        RECT 26.030 60.450 26.200 63.030 ;
        RECT 28.060 62.350 28.400 63.980 ;
        RECT 28.740 63.890 30.520 63.980 ;
        RECT 29.280 63.100 29.450 63.890 ;
        RECT 30.240 63.100 30.410 63.890 ;
        RECT 32.640 63.590 33.070 64.480 ;
        RECT 32.760 62.880 32.930 63.590 ;
        RECT 27.710 62.010 28.400 62.350 ;
        RECT 17.320 60.240 20.370 60.310 ;
        RECT 24.080 60.260 26.340 60.450 ;
        RECT 27.710 60.260 28.110 62.010 ;
        RECT 16.750 60.030 20.840 60.240 ;
        RECT 17.370 58.540 19.670 60.030 ;
        RECT 27.710 59.910 32.570 60.260 ;
        RECT 30.270 58.540 32.570 59.910 ;
        RECT 14.520 58.140 35.420 58.540 ;
        RECT 14.520 51.840 14.920 58.140 ;
        RECT 17.370 58.090 19.670 58.140 ;
        RECT 30.270 58.090 32.570 58.140 ;
        RECT 15.720 56.940 34.220 57.540 ;
        RECT 18.320 56.340 18.670 56.940 ;
        RECT 16.070 56.140 18.670 56.340 ;
        RECT 18.320 55.540 18.670 56.140 ;
        RECT 16.070 55.340 18.670 55.540 ;
        RECT 19.270 55.440 19.470 56.940 ;
        RECT 20.070 55.440 20.270 56.940 ;
        RECT 20.870 55.440 21.070 56.940 ;
        RECT 21.670 55.440 21.870 56.940 ;
        RECT 22.470 55.440 22.670 56.940 ;
        RECT 23.270 55.440 23.470 56.940 ;
        RECT 24.070 55.440 24.270 56.940 ;
        RECT 24.870 55.440 25.070 56.940 ;
        RECT 25.670 55.440 25.870 56.940 ;
        RECT 26.470 55.440 26.670 56.940 ;
        RECT 27.270 55.440 27.470 56.940 ;
        RECT 28.070 55.440 28.270 56.940 ;
        RECT 28.870 55.440 29.070 56.940 ;
        RECT 29.670 55.440 29.870 56.940 ;
        RECT 30.470 55.440 30.670 56.940 ;
        RECT 31.270 56.340 31.620 56.940 ;
        RECT 31.270 56.140 33.870 56.340 ;
        RECT 31.270 55.540 31.620 56.140 ;
        RECT 31.270 55.340 33.820 55.540 ;
        RECT 16.070 54.440 18.670 54.640 ;
        RECT 18.320 53.840 18.670 54.440 ;
        RECT 16.070 53.640 18.670 53.840 ;
        RECT 18.320 53.040 18.670 53.640 ;
        RECT 19.270 53.040 19.470 54.540 ;
        RECT 20.070 53.040 20.270 54.540 ;
        RECT 20.870 53.040 21.070 54.540 ;
        RECT 21.670 53.040 21.870 54.540 ;
        RECT 22.470 53.040 22.670 54.540 ;
        RECT 23.270 53.040 23.470 54.540 ;
        RECT 24.070 53.040 24.270 54.540 ;
        RECT 24.870 53.040 25.070 54.540 ;
        RECT 25.670 53.040 25.870 54.540 ;
        RECT 26.470 53.040 26.670 54.540 ;
        RECT 27.270 53.040 27.470 54.540 ;
        RECT 28.070 53.040 28.270 54.540 ;
        RECT 28.870 53.040 29.070 54.540 ;
        RECT 29.670 53.040 29.870 54.540 ;
        RECT 30.470 53.040 30.670 54.540 ;
        RECT 31.270 54.440 33.820 54.640 ;
        RECT 31.270 53.840 31.620 54.440 ;
        RECT 31.270 53.640 33.870 53.840 ;
        RECT 31.270 53.040 31.620 53.640 ;
        RECT 15.720 52.440 34.220 53.040 ;
        RECT 17.370 51.840 19.670 51.890 ;
        RECT 30.270 51.840 32.570 51.890 ;
        RECT 35.020 51.840 35.420 58.140 ;
        RECT 14.520 51.440 35.420 51.840 ;
        RECT 17.370 50.990 19.670 51.440 ;
        RECT 30.270 50.990 32.570 51.440 ;
        RECT 36.340 50.990 37.330 64.480 ;
        RECT 12.940 50.000 37.330 50.990 ;
      LAYER mcon ;
        RECT 13.120 74.740 13.770 76.740 ;
        RECT 13.040 71.840 13.720 74.040 ;
        RECT 13.040 69.090 13.820 71.240 ;
        RECT 15.820 74.990 16.420 75.490 ;
        RECT 16.620 74.990 17.220 75.490 ;
        RECT 17.420 74.990 18.020 75.490 ;
        RECT 18.220 74.990 18.820 75.490 ;
        RECT 31.120 74.990 31.720 75.490 ;
        RECT 31.920 74.990 32.520 75.490 ;
        RECT 32.720 74.990 33.320 75.490 ;
        RECT 33.520 74.990 34.120 75.490 ;
        RECT 15.820 70.390 16.420 70.890 ;
        RECT 16.620 70.390 17.220 70.890 ;
        RECT 17.420 70.390 18.020 70.890 ;
        RECT 18.220 70.390 18.820 70.890 ;
        RECT 31.120 70.390 31.720 70.890 ;
        RECT 31.920 70.390 32.520 70.890 ;
        RECT 32.720 70.390 33.320 70.890 ;
        RECT 33.520 70.390 34.120 70.890 ;
        RECT 13.020 60.610 13.190 60.780 ;
        RECT 13.380 60.610 13.550 60.780 ;
        RECT 13.740 60.610 13.910 60.780 ;
        RECT 14.660 60.560 14.840 60.730 ;
        RECT 15.830 60.560 16.010 60.730 ;
        RECT 13.020 60.250 13.190 60.420 ;
        RECT 13.380 60.250 13.550 60.420 ;
        RECT 13.740 60.250 13.910 60.420 ;
        RECT 24.200 60.270 24.380 60.450 ;
        RECT 24.660 60.270 24.840 60.450 ;
        RECT 25.120 60.270 25.300 60.450 ;
        RECT 25.580 60.270 25.760 60.450 ;
        RECT 26.040 60.270 26.220 60.450 ;
        RECT 36.410 60.610 36.580 60.780 ;
        RECT 36.770 60.610 36.940 60.780 ;
        RECT 37.130 60.610 37.300 60.780 ;
        RECT 13.020 59.890 13.190 60.060 ;
        RECT 13.380 59.890 13.550 60.060 ;
        RECT 13.740 59.890 13.910 60.060 ;
        RECT 16.870 60.050 17.050 60.230 ;
        RECT 17.460 60.050 17.640 60.230 ;
        RECT 18.050 60.050 18.230 60.230 ;
        RECT 18.640 60.050 18.820 60.230 ;
        RECT 19.230 60.050 19.410 60.230 ;
        RECT 19.820 60.050 20.000 60.230 ;
        RECT 20.410 60.050 20.590 60.230 ;
        RECT 13.020 59.530 13.190 59.700 ;
        RECT 13.380 59.530 13.550 59.700 ;
        RECT 13.740 59.530 13.910 59.700 ;
        RECT 13.010 59.170 13.180 59.340 ;
        RECT 13.370 59.170 13.540 59.340 ;
        RECT 13.730 59.170 13.900 59.340 ;
        RECT 13.030 56.690 13.820 58.840 ;
        RECT 27.750 59.980 27.930 60.160 ;
        RECT 28.120 59.990 28.300 60.170 ;
        RECT 28.520 59.990 28.700 60.170 ;
        RECT 28.920 59.990 29.100 60.170 ;
        RECT 29.320 59.990 29.500 60.170 ;
        RECT 36.410 60.250 36.580 60.420 ;
        RECT 36.770 60.250 36.940 60.420 ;
        RECT 37.130 60.250 37.300 60.420 ;
        RECT 36.410 59.890 36.580 60.060 ;
        RECT 36.770 59.890 36.940 60.060 ;
        RECT 37.130 59.890 37.300 60.060 ;
        RECT 36.410 59.530 36.580 59.700 ;
        RECT 36.770 59.530 36.940 59.700 ;
        RECT 37.130 59.530 37.300 59.700 ;
        RECT 36.410 59.170 36.580 59.340 ;
        RECT 36.770 59.170 36.940 59.340 ;
        RECT 37.130 59.170 37.300 59.340 ;
        RECT 13.070 53.890 13.720 56.090 ;
        RECT 13.070 51.190 13.870 53.240 ;
        RECT 15.820 57.040 16.420 57.540 ;
        RECT 16.620 57.040 17.220 57.540 ;
        RECT 17.420 57.040 18.020 57.540 ;
        RECT 18.220 57.040 18.820 57.540 ;
        RECT 31.120 57.040 31.720 57.540 ;
        RECT 31.920 57.040 32.520 57.540 ;
        RECT 32.720 57.040 33.320 57.540 ;
        RECT 33.520 57.040 34.120 57.540 ;
        RECT 15.820 52.440 16.420 52.940 ;
        RECT 16.620 52.440 17.220 52.940 ;
        RECT 17.420 52.440 18.020 52.940 ;
        RECT 18.220 52.440 18.820 52.940 ;
        RECT 31.120 52.440 31.720 52.940 ;
        RECT 31.920 52.440 32.520 52.940 ;
        RECT 32.720 52.440 33.320 52.940 ;
        RECT 33.520 52.440 34.120 52.940 ;
      LAYER met1 ;
        RECT 12.940 75.690 17.320 76.890 ;
        RECT 32.620 75.690 35.820 76.890 ;
        RECT 12.940 75.540 16.420 75.690 ;
        RECT 33.520 75.540 35.820 75.690 ;
        RECT 12.940 75.390 24.520 75.540 ;
        RECT 25.420 75.390 35.820 75.540 ;
        RECT 12.940 74.940 18.920 75.390 ;
        RECT 31.020 74.940 35.820 75.390 ;
        RECT 12.940 74.540 15.320 74.940 ;
        RECT 15.770 74.890 24.520 74.940 ;
        RECT 12.940 71.740 13.820 74.140 ;
        RECT 14.120 74.040 15.320 74.540 ;
        RECT 15.920 73.540 16.070 74.890 ;
        RECT 16.520 73.540 16.670 74.890 ;
        RECT 17.120 73.540 17.270 74.890 ;
        RECT 17.720 73.540 17.870 74.890 ;
        RECT 18.320 74.790 24.520 74.890 ;
        RECT 25.420 74.890 34.170 74.940 ;
        RECT 25.420 74.790 31.620 74.890 ;
        RECT 18.320 74.340 18.920 74.790 ;
        RECT 31.020 74.340 31.620 74.790 ;
        RECT 18.320 74.190 24.520 74.340 ;
        RECT 25.420 74.190 31.620 74.340 ;
        RECT 18.320 73.740 18.920 74.190 ;
        RECT 31.020 73.740 31.620 74.190 ;
        RECT 18.320 73.590 24.520 73.740 ;
        RECT 25.420 73.590 31.620 73.740 ;
        RECT 18.320 73.390 18.920 73.590 ;
        RECT 31.020 73.390 31.620 73.590 ;
        RECT 32.070 73.540 32.220 74.890 ;
        RECT 32.670 73.540 32.820 74.890 ;
        RECT 33.270 73.540 33.420 74.890 ;
        RECT 33.870 73.540 34.020 74.890 ;
        RECT 34.620 74.040 35.820 74.940 ;
        RECT 14.120 71.340 15.320 71.840 ;
        RECT 12.940 70.940 15.320 71.340 ;
        RECT 15.920 70.990 16.070 72.290 ;
        RECT 16.520 70.990 16.670 72.290 ;
        RECT 17.120 70.990 17.270 72.290 ;
        RECT 17.720 70.990 17.870 72.290 ;
        RECT 18.320 72.140 24.520 72.290 ;
        RECT 25.420 72.140 31.620 72.290 ;
        RECT 18.320 71.690 18.920 72.140 ;
        RECT 31.020 71.690 31.620 72.140 ;
        RECT 18.320 71.540 24.520 71.690 ;
        RECT 25.420 71.540 31.620 71.690 ;
        RECT 18.320 71.090 18.920 71.540 ;
        RECT 31.020 71.090 31.620 71.540 ;
        RECT 18.320 70.990 24.520 71.090 ;
        RECT 15.770 70.940 24.520 70.990 ;
        RECT 25.420 70.990 31.620 71.090 ;
        RECT 32.070 70.990 32.220 72.290 ;
        RECT 32.670 70.990 32.820 72.290 ;
        RECT 33.270 70.990 33.420 72.290 ;
        RECT 33.870 70.990 34.020 72.290 ;
        RECT 25.420 70.940 34.170 70.990 ;
        RECT 34.620 70.940 35.820 71.840 ;
        RECT 12.940 70.490 18.920 70.940 ;
        RECT 31.020 70.490 35.820 70.940 ;
        RECT 12.940 70.340 24.520 70.490 ;
        RECT 25.420 70.340 35.820 70.490 ;
        RECT 12.940 70.190 16.420 70.340 ;
        RECT 33.520 70.190 35.820 70.340 ;
        RECT 12.940 68.990 17.320 70.190 ;
        RECT 32.620 68.990 35.820 70.190 ;
        RECT 12.940 60.780 13.940 60.880 ;
        RECT 12.940 60.260 16.210 60.780 ;
        RECT 24.080 60.260 26.340 60.480 ;
        RECT 36.340 60.260 37.330 60.880 ;
        RECT 10.000 59.100 38.570 60.260 ;
        RECT 12.930 57.740 17.320 58.940 ;
        RECT 32.620 57.740 35.820 58.940 ;
        RECT 12.930 57.590 16.420 57.740 ;
        RECT 33.520 57.590 35.820 57.740 ;
        RECT 12.930 57.440 24.520 57.590 ;
        RECT 25.420 57.440 35.820 57.590 ;
        RECT 12.930 56.990 18.920 57.440 ;
        RECT 31.020 56.990 35.820 57.440 ;
        RECT 12.930 56.590 15.320 56.990 ;
        RECT 15.770 56.940 24.520 56.990 ;
        RECT 12.940 53.790 13.820 56.190 ;
        RECT 14.120 56.090 15.320 56.590 ;
        RECT 15.920 55.590 16.070 56.940 ;
        RECT 16.520 55.590 16.670 56.940 ;
        RECT 17.120 55.590 17.270 56.940 ;
        RECT 17.720 55.590 17.870 56.940 ;
        RECT 18.320 56.840 24.520 56.940 ;
        RECT 25.420 56.940 34.170 56.990 ;
        RECT 25.420 56.840 31.620 56.940 ;
        RECT 18.320 56.390 18.920 56.840 ;
        RECT 31.020 56.390 31.620 56.840 ;
        RECT 18.320 56.240 24.520 56.390 ;
        RECT 25.420 56.240 31.620 56.390 ;
        RECT 18.320 55.790 18.920 56.240 ;
        RECT 31.020 55.790 31.620 56.240 ;
        RECT 18.320 55.640 24.520 55.790 ;
        RECT 25.420 55.640 31.620 55.790 ;
        RECT 18.320 55.440 18.920 55.640 ;
        RECT 31.020 55.440 31.620 55.640 ;
        RECT 32.070 55.590 32.220 56.940 ;
        RECT 32.670 55.590 32.820 56.940 ;
        RECT 33.270 55.590 33.420 56.940 ;
        RECT 33.870 55.590 34.020 56.940 ;
        RECT 34.620 56.090 35.820 56.990 ;
        RECT 14.120 53.390 15.320 53.890 ;
        RECT 12.940 52.990 15.320 53.390 ;
        RECT 15.920 53.040 16.070 54.340 ;
        RECT 16.520 53.040 16.670 54.340 ;
        RECT 17.120 53.040 17.270 54.340 ;
        RECT 17.720 53.040 17.870 54.340 ;
        RECT 18.320 54.190 24.520 54.340 ;
        RECT 25.420 54.190 31.620 54.340 ;
        RECT 18.320 53.740 18.920 54.190 ;
        RECT 31.020 53.740 31.620 54.190 ;
        RECT 18.320 53.590 24.520 53.740 ;
        RECT 25.420 53.590 31.620 53.740 ;
        RECT 18.320 53.140 18.920 53.590 ;
        RECT 31.020 53.140 31.620 53.590 ;
        RECT 18.320 53.040 24.520 53.140 ;
        RECT 15.770 52.990 24.520 53.040 ;
        RECT 25.420 53.040 31.620 53.140 ;
        RECT 32.070 53.040 32.220 54.340 ;
        RECT 32.670 53.040 32.820 54.340 ;
        RECT 33.270 53.040 33.420 54.340 ;
        RECT 33.870 53.040 34.020 54.340 ;
        RECT 25.420 52.990 34.170 53.040 ;
        RECT 34.620 52.990 35.820 53.890 ;
        RECT 12.940 52.540 18.920 52.990 ;
        RECT 31.020 52.540 35.820 52.990 ;
        RECT 12.940 52.390 24.520 52.540 ;
        RECT 25.420 52.390 35.820 52.540 ;
        RECT 12.940 52.240 16.420 52.390 ;
        RECT 33.520 52.240 35.820 52.390 ;
        RECT 12.940 51.040 17.320 52.240 ;
        RECT 32.620 51.040 35.820 52.240 ;
      LAYER via ;
        RECT 13.120 74.740 13.770 76.740 ;
        RECT 14.220 75.790 15.220 76.790 ;
        RECT 16.220 75.790 17.220 76.790 ;
        RECT 32.720 75.790 33.720 76.790 ;
        RECT 34.720 75.790 35.720 76.790 ;
        RECT 14.220 74.190 15.220 75.190 ;
        RECT 13.040 71.840 13.720 74.040 ;
        RECT 34.720 74.190 35.720 75.190 ;
        RECT 14.220 70.690 15.220 71.690 ;
        RECT 34.720 70.690 35.720 71.690 ;
        RECT 14.220 69.090 15.220 70.090 ;
        RECT 16.220 69.090 17.220 70.090 ;
        RECT 32.720 69.090 33.720 70.090 ;
        RECT 34.720 69.090 35.720 70.090 ;
        RECT 11.720 59.190 12.520 60.140 ;
        RECT 14.220 59.290 17.000 60.120 ;
        RECT 37.670 59.190 38.470 60.140 ;
        RECT 14.220 57.840 15.220 58.840 ;
        RECT 16.220 57.840 17.220 58.840 ;
        RECT 32.720 57.840 33.720 58.840 ;
        RECT 34.720 57.840 35.720 58.840 ;
        RECT 14.220 56.240 15.220 57.240 ;
        RECT 13.070 53.890 13.720 56.090 ;
        RECT 34.720 56.240 35.720 57.240 ;
        RECT 13.070 51.190 13.730 53.240 ;
        RECT 14.220 52.740 15.220 53.740 ;
        RECT 34.720 52.740 35.720 53.740 ;
        RECT 14.220 51.140 15.220 52.140 ;
        RECT 16.220 51.140 17.220 52.140 ;
        RECT 32.720 51.140 33.720 52.140 ;
        RECT 34.720 51.140 35.720 52.140 ;
      LAYER met2 ;
        RECT 12.940 75.690 17.320 76.890 ;
        RECT 32.620 75.690 35.820 76.890 ;
        RECT 12.940 74.740 16.070 75.690 ;
        RECT 33.870 74.740 35.820 75.690 ;
        RECT 12.940 74.590 18.070 74.740 ;
        RECT 12.940 74.540 16.070 74.590 ;
        RECT 14.120 74.140 16.070 74.540 ;
        RECT 12.940 71.740 13.820 74.140 ;
        RECT 14.120 74.040 18.070 74.140 ;
        RECT 15.520 73.990 18.070 74.040 ;
        RECT 15.520 73.390 16.070 73.990 ;
        RECT 15.520 73.090 18.070 73.390 ;
        RECT 18.670 73.090 18.820 74.740 ;
        RECT 19.270 73.090 19.420 74.740 ;
        RECT 19.870 73.090 20.020 74.740 ;
        RECT 20.470 73.090 20.620 74.740 ;
        RECT 21.070 73.090 21.220 74.740 ;
        RECT 21.670 73.090 21.820 74.740 ;
        RECT 22.270 73.090 22.420 74.740 ;
        RECT 22.870 73.090 23.020 74.740 ;
        RECT 23.470 73.090 23.620 74.740 ;
        RECT 24.070 73.090 24.220 74.740 ;
        RECT 24.670 73.090 25.270 74.740 ;
        RECT 25.720 73.090 25.870 74.740 ;
        RECT 26.320 73.090 26.470 74.740 ;
        RECT 26.920 73.090 27.070 74.740 ;
        RECT 27.520 73.090 27.670 74.740 ;
        RECT 28.120 73.090 28.270 74.740 ;
        RECT 28.720 73.090 28.870 74.740 ;
        RECT 29.320 73.090 29.470 74.740 ;
        RECT 29.920 73.090 30.070 74.740 ;
        RECT 30.520 73.090 30.670 74.740 ;
        RECT 31.120 73.090 31.270 74.740 ;
        RECT 31.870 74.590 35.820 74.740 ;
        RECT 33.870 74.140 35.820 74.590 ;
        RECT 31.870 74.040 35.820 74.140 ;
        RECT 31.870 73.990 34.420 74.040 ;
        RECT 33.870 73.390 34.420 73.990 ;
        RECT 31.870 73.090 34.420 73.390 ;
        RECT 15.520 72.790 34.420 73.090 ;
        RECT 15.520 72.340 18.070 72.790 ;
        RECT 15.520 71.890 16.070 72.340 ;
        RECT 15.520 71.840 18.070 71.890 ;
        RECT 14.120 71.740 18.070 71.840 ;
        RECT 14.120 71.290 16.070 71.740 ;
        RECT 14.120 71.140 18.070 71.290 ;
        RECT 18.670 71.140 18.820 72.790 ;
        RECT 19.270 71.140 19.420 72.790 ;
        RECT 19.870 71.140 20.020 72.790 ;
        RECT 20.470 71.140 20.620 72.790 ;
        RECT 21.070 71.140 21.220 72.790 ;
        RECT 21.670 71.140 21.820 72.790 ;
        RECT 22.270 71.140 22.420 72.790 ;
        RECT 22.870 71.140 23.020 72.790 ;
        RECT 23.470 71.140 23.620 72.790 ;
        RECT 24.070 71.140 24.220 72.790 ;
        RECT 24.670 71.140 25.270 72.790 ;
        RECT 25.720 71.140 25.870 72.790 ;
        RECT 26.320 71.140 26.470 72.790 ;
        RECT 26.920 71.140 27.070 72.790 ;
        RECT 27.520 71.140 27.670 72.790 ;
        RECT 28.120 71.140 28.270 72.790 ;
        RECT 28.720 71.140 28.870 72.790 ;
        RECT 29.320 71.140 29.470 72.790 ;
        RECT 29.920 71.140 30.070 72.790 ;
        RECT 30.520 71.140 30.670 72.790 ;
        RECT 31.120 71.140 31.270 72.790 ;
        RECT 31.870 72.340 34.420 72.790 ;
        RECT 33.870 71.890 34.420 72.340 ;
        RECT 31.870 71.840 34.420 71.890 ;
        RECT 31.870 71.740 35.820 71.840 ;
        RECT 33.870 71.290 35.820 71.740 ;
        RECT 31.870 71.140 35.820 71.290 ;
        RECT 14.120 70.190 16.070 71.140 ;
        RECT 33.870 70.190 35.820 71.140 ;
        RECT 14.120 68.990 17.320 70.190 ;
        RECT 32.620 68.990 35.820 70.190 ;
        RECT 11.610 59.100 12.610 60.260 ;
        RECT 14.080 59.260 17.230 60.260 ;
        RECT 14.120 58.940 17.270 59.260 ;
        RECT 37.570 59.100 38.570 60.260 ;
        RECT 14.120 57.740 17.320 58.940 ;
        RECT 32.620 57.740 35.820 58.940 ;
        RECT 14.120 56.790 16.070 57.740 ;
        RECT 33.870 56.790 35.820 57.740 ;
        RECT 14.120 56.640 18.070 56.790 ;
        RECT 14.120 56.190 16.070 56.640 ;
        RECT 12.940 53.790 13.820 56.190 ;
        RECT 14.120 56.090 18.070 56.190 ;
        RECT 15.520 56.040 18.070 56.090 ;
        RECT 15.520 55.440 16.070 56.040 ;
        RECT 15.520 55.140 18.070 55.440 ;
        RECT 18.670 55.140 18.820 56.790 ;
        RECT 19.270 55.140 19.420 56.790 ;
        RECT 19.870 55.140 20.020 56.790 ;
        RECT 20.470 55.140 20.620 56.790 ;
        RECT 21.070 55.140 21.220 56.790 ;
        RECT 21.670 55.140 21.820 56.790 ;
        RECT 22.270 55.140 22.420 56.790 ;
        RECT 22.870 55.140 23.020 56.790 ;
        RECT 23.470 55.140 23.620 56.790 ;
        RECT 24.070 55.140 24.220 56.790 ;
        RECT 24.670 55.140 25.270 56.790 ;
        RECT 25.720 55.140 25.870 56.790 ;
        RECT 26.320 55.140 26.470 56.790 ;
        RECT 26.920 55.140 27.070 56.790 ;
        RECT 27.520 55.140 27.670 56.790 ;
        RECT 28.120 55.140 28.270 56.790 ;
        RECT 28.720 55.140 28.870 56.790 ;
        RECT 29.320 55.140 29.470 56.790 ;
        RECT 29.920 55.140 30.070 56.790 ;
        RECT 30.520 55.140 30.670 56.790 ;
        RECT 31.120 55.140 31.270 56.790 ;
        RECT 31.870 56.640 35.820 56.790 ;
        RECT 33.870 56.190 35.820 56.640 ;
        RECT 31.870 56.090 35.820 56.190 ;
        RECT 31.870 56.040 34.420 56.090 ;
        RECT 33.870 55.440 34.420 56.040 ;
        RECT 31.870 55.140 34.420 55.440 ;
        RECT 15.520 54.840 34.420 55.140 ;
        RECT 15.520 54.390 18.070 54.840 ;
        RECT 15.520 53.940 16.070 54.390 ;
        RECT 15.520 53.890 18.070 53.940 ;
        RECT 14.120 53.790 18.070 53.890 ;
        RECT 14.120 53.390 16.070 53.790 ;
        RECT 12.940 53.340 16.070 53.390 ;
        RECT 12.940 53.190 18.070 53.340 ;
        RECT 18.670 53.190 18.820 54.840 ;
        RECT 19.270 53.190 19.420 54.840 ;
        RECT 19.870 53.190 20.020 54.840 ;
        RECT 20.470 53.190 20.620 54.840 ;
        RECT 21.070 53.190 21.220 54.840 ;
        RECT 21.670 53.190 21.820 54.840 ;
        RECT 22.270 53.190 22.420 54.840 ;
        RECT 22.870 53.190 23.020 54.840 ;
        RECT 23.470 53.190 23.620 54.840 ;
        RECT 24.070 53.190 24.220 54.840 ;
        RECT 24.670 53.190 25.270 54.840 ;
        RECT 25.720 53.190 25.870 54.840 ;
        RECT 26.320 53.190 26.470 54.840 ;
        RECT 26.920 53.190 27.070 54.840 ;
        RECT 27.520 53.190 27.670 54.840 ;
        RECT 28.120 53.190 28.270 54.840 ;
        RECT 28.720 53.190 28.870 54.840 ;
        RECT 29.320 53.190 29.470 54.840 ;
        RECT 29.920 53.190 30.070 54.840 ;
        RECT 30.520 53.190 30.670 54.840 ;
        RECT 31.120 53.190 31.270 54.840 ;
        RECT 31.870 54.390 34.420 54.840 ;
        RECT 33.870 53.940 34.420 54.390 ;
        RECT 31.870 53.890 34.420 53.940 ;
        RECT 31.870 53.790 35.820 53.890 ;
        RECT 33.870 53.340 35.820 53.790 ;
        RECT 31.870 53.190 35.820 53.340 ;
        RECT 12.940 52.240 16.070 53.190 ;
        RECT 33.870 52.240 35.820 53.190 ;
        RECT 12.940 51.040 17.320 52.240 ;
        RECT 32.620 51.040 35.820 52.240 ;
      LAYER via2 ;
        RECT 13.120 74.740 13.770 76.740 ;
        RECT 13.040 71.840 13.720 74.040 ;
        RECT 11.720 59.190 12.520 60.140 ;
        RECT 14.220 59.290 17.000 60.120 ;
        RECT 37.670 59.190 38.470 60.140 ;
        RECT 13.070 53.890 13.720 56.090 ;
        RECT 13.070 51.190 13.730 53.240 ;
      LAYER met3 ;
        RECT 12.940 74.540 13.810 76.890 ;
        RECT 14.120 75.640 17.320 76.890 ;
        RECT 19.720 76.040 30.220 76.890 ;
        RECT 32.620 75.640 35.820 76.890 ;
        RECT 14.120 74.490 35.820 75.640 ;
        RECT 12.940 71.740 13.820 74.140 ;
        RECT 14.120 71.740 14.970 74.140 ;
        RECT 15.370 71.390 34.570 74.490 ;
        RECT 34.970 71.740 35.820 74.140 ;
        RECT 14.120 70.240 35.820 71.390 ;
        RECT 14.120 68.990 17.320 70.240 ;
        RECT 19.720 68.990 30.220 69.840 ;
        RECT 32.620 68.990 35.820 70.240 ;
        RECT 11.610 59.100 12.610 60.260 ;
        RECT 14.080 59.260 17.230 60.260 ;
        RECT 37.570 59.100 38.570 60.260 ;
        RECT 14.120 57.690 17.320 58.940 ;
        RECT 19.720 58.090 30.220 58.940 ;
        RECT 32.620 57.690 35.820 58.940 ;
        RECT 14.120 56.540 35.820 57.690 ;
        RECT 12.940 53.790 13.820 56.190 ;
        RECT 14.120 53.790 14.970 56.190 ;
        RECT 15.370 53.440 34.570 56.540 ;
        RECT 34.970 53.790 35.820 56.190 ;
        RECT 12.940 51.040 13.800 53.390 ;
        RECT 14.120 52.290 35.820 53.440 ;
        RECT 14.120 51.040 17.320 52.290 ;
        RECT 19.720 51.040 30.220 51.890 ;
        RECT 32.620 51.040 35.820 52.290 ;
      LAYER via3 ;
        RECT 13.120 74.740 13.770 76.740 ;
        RECT 14.220 75.940 15.070 76.790 ;
        RECT 16.320 75.940 17.170 76.790 ;
        RECT 19.820 76.140 20.470 76.790 ;
        RECT 20.620 76.140 21.270 76.790 ;
        RECT 28.670 76.140 29.320 76.790 ;
        RECT 29.470 76.140 30.120 76.790 ;
        RECT 32.770 75.940 33.620 76.790 ;
        RECT 34.870 75.940 35.720 76.790 ;
        RECT 14.220 74.640 15.070 75.490 ;
        RECT 34.870 74.640 35.720 75.490 ;
        RECT 13.040 71.840 13.720 74.040 ;
        RECT 14.220 73.040 14.870 74.040 ;
        RECT 14.220 71.840 14.870 72.840 ;
        RECT 35.070 73.040 35.720 74.040 ;
        RECT 35.070 71.840 35.720 72.840 ;
        RECT 14.220 70.390 15.070 71.240 ;
        RECT 34.870 70.390 35.720 71.240 ;
        RECT 14.220 69.090 15.070 69.940 ;
        RECT 16.320 69.090 17.170 69.940 ;
        RECT 19.820 69.090 20.470 69.740 ;
        RECT 20.620 69.090 21.270 69.740 ;
        RECT 28.670 69.090 29.320 69.740 ;
        RECT 29.470 69.090 30.120 69.740 ;
        RECT 32.770 69.090 33.620 69.940 ;
        RECT 34.870 69.090 35.720 69.940 ;
        RECT 11.720 59.190 12.520 60.140 ;
        RECT 37.670 59.190 38.470 60.140 ;
        RECT 14.220 57.990 15.070 58.840 ;
        RECT 16.320 57.990 17.170 58.840 ;
        RECT 19.820 58.190 20.470 58.840 ;
        RECT 20.620 58.190 21.270 58.840 ;
        RECT 28.670 58.190 29.320 58.840 ;
        RECT 29.470 58.190 30.120 58.840 ;
        RECT 32.770 57.990 33.620 58.840 ;
        RECT 34.870 57.990 35.720 58.840 ;
        RECT 14.220 56.690 15.070 57.540 ;
        RECT 34.870 56.690 35.720 57.540 ;
        RECT 13.070 53.890 13.720 56.090 ;
        RECT 14.220 55.090 14.870 56.090 ;
        RECT 14.220 53.890 14.870 54.890 ;
        RECT 35.070 55.090 35.720 56.090 ;
        RECT 35.070 53.890 35.720 54.890 ;
        RECT 13.070 51.190 13.730 53.240 ;
        RECT 14.220 52.440 15.070 53.290 ;
        RECT 34.870 52.440 35.720 53.290 ;
        RECT 14.220 51.140 15.070 51.990 ;
        RECT 16.320 51.140 17.170 51.990 ;
        RECT 19.820 51.140 20.470 51.790 ;
        RECT 20.620 51.140 21.270 51.790 ;
        RECT 28.670 51.140 29.320 51.790 ;
        RECT 29.470 51.140 30.120 51.790 ;
        RECT 32.770 51.140 33.620 51.990 ;
        RECT 34.870 51.140 35.720 51.990 ;
      LAYER met4 ;
        RECT 11.610 50.000 12.610 77.980 ;
        RECT 12.940 75.840 17.270 76.890 ;
        RECT 12.940 74.540 15.170 75.840 ;
        RECT 19.720 75.440 30.220 76.890 ;
        RECT 32.670 75.840 35.820 76.890 ;
        RECT 15.570 74.140 34.370 75.440 ;
        RECT 34.770 74.540 35.820 75.840 ;
        RECT 12.940 71.740 35.820 74.140 ;
        RECT 14.120 70.040 15.170 71.340 ;
        RECT 15.570 70.440 34.370 71.740 ;
        RECT 14.120 68.990 17.270 70.040 ;
        RECT 19.720 68.990 30.220 70.440 ;
        RECT 34.770 70.040 35.820 71.340 ;
        RECT 32.670 68.990 35.820 70.040 ;
        RECT 14.120 57.890 17.270 58.940 ;
        RECT 14.120 56.590 15.170 57.890 ;
        RECT 19.720 57.490 30.220 58.940 ;
        RECT 32.670 57.890 35.820 58.940 ;
        RECT 15.570 56.190 34.370 57.490 ;
        RECT 34.770 56.590 35.820 57.890 ;
        RECT 12.940 53.790 35.820 56.190 ;
        RECT 12.940 52.090 15.170 53.390 ;
        RECT 15.570 52.490 34.370 53.790 ;
        RECT 12.940 51.040 17.270 52.090 ;
        RECT 19.720 51.040 30.220 52.490 ;
        RECT 34.770 52.090 35.820 53.390 ;
        RECT 32.670 51.040 35.820 52.090 ;
        RECT 37.570 50.000 38.570 77.980 ;
    END
  END VGND
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.189000 ;
    PORT
      LAYER li1 ;
        RECT 14.100 61.790 14.370 62.120 ;
      LAYER mcon ;
        RECT 14.180 61.870 14.350 62.040 ;
      LAYER met1 ;
        RECT 14.070 62.030 14.380 62.120 ;
        RECT 10.000 61.890 14.380 62.030 ;
        RECT 14.070 61.790 14.380 61.890 ;
    END
  END clk
  PIN inp
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.200000 ;
    PORT
      LAYER li1 ;
        RECT 19.630 65.220 19.990 65.520 ;
      LAYER mcon ;
        RECT 19.710 65.270 19.910 65.470 ;
      LAYER met1 ;
        RECT 10.000 65.410 19.990 65.550 ;
        RECT 19.630 65.220 19.990 65.410 ;
    END
  END inp
  PIN inn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.200000 ;
    PORT
      LAYER li1 ;
        RECT 17.670 64.970 18.030 65.270 ;
      LAYER mcon ;
        RECT 17.750 65.020 17.950 65.220 ;
      LAYER met1 ;
        RECT 10.000 65.130 18.030 65.270 ;
        RECT 17.670 64.970 18.030 65.130 ;
    END
  END inn
  PIN comp_trig
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.756400 ;
    PORT
      LAYER li1 ;
        RECT 32.280 61.230 32.450 63.340 ;
        RECT 33.240 62.880 33.510 63.340 ;
        RECT 33.340 62.780 33.510 62.880 ;
        RECT 33.340 62.590 35.370 62.780 ;
        RECT 34.200 61.230 34.370 62.590 ;
        RECT 34.690 62.540 35.370 62.590 ;
      LAYER mcon ;
        RECT 32.280 62.960 32.450 63.260 ;
        RECT 33.240 62.960 33.410 63.260 ;
        RECT 34.750 62.570 34.930 62.750 ;
        RECT 35.130 62.570 35.310 62.750 ;
      LAYER met1 ;
        RECT 32.250 63.180 32.480 63.320 ;
        RECT 33.210 63.180 33.440 63.320 ;
        RECT 32.250 63.040 33.440 63.180 ;
        RECT 32.250 62.900 32.480 63.040 ;
        RECT 33.210 62.900 33.440 63.040 ;
        RECT 34.690 62.730 35.370 62.780 ;
        RECT 34.690 62.590 40.050 62.730 ;
        RECT 34.690 62.540 35.370 62.590 ;
    END
  END comp_trig
  PIN latch_qn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.303000 ;
    ANTENNADIFFAREA 0.756400 ;
    PORT
      LAYER li1 ;
        RECT 32.060 65.810 32.390 66.070 ;
        RECT 33.960 64.980 34.130 67.090 ;
        RECT 35.880 65.730 36.050 67.090 ;
        RECT 35.020 65.540 36.170 65.730 ;
        RECT 35.020 65.440 35.190 65.540 ;
        RECT 35.500 65.490 36.170 65.540 ;
        RECT 34.920 64.980 35.190 65.440 ;
      LAYER mcon ;
        RECT 32.140 65.860 32.310 66.030 ;
        RECT 35.560 65.520 35.740 65.700 ;
        RECT 35.930 65.520 36.110 65.700 ;
        RECT 33.960 65.060 34.130 65.360 ;
        RECT 34.920 65.060 35.090 65.360 ;
      LAYER met1 ;
        RECT 32.060 66.050 32.390 66.070 ;
        RECT 31.400 65.870 33.190 66.050 ;
        RECT 32.060 65.810 32.390 65.870 ;
        RECT 33.010 65.310 33.190 65.870 ;
        RECT 35.500 65.680 36.170 65.730 ;
        RECT 35.500 65.540 40.050 65.680 ;
        RECT 35.500 65.490 36.170 65.540 ;
        RECT 33.930 65.310 34.160 65.420 ;
        RECT 33.010 65.280 34.160 65.310 ;
        RECT 34.890 65.280 35.120 65.420 ;
        RECT 33.010 65.140 35.120 65.280 ;
        RECT 33.010 65.130 34.160 65.140 ;
        RECT 33.930 65.000 34.160 65.130 ;
        RECT 34.890 65.000 35.120 65.140 ;
    END
  END latch_qn
  PIN latch_q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.303000 ;
    ANTENNADIFFAREA 0.756400 ;
    PORT
      LAYER li1 ;
        RECT 31.480 64.980 31.650 67.090 ;
        RECT 33.400 65.780 33.570 67.090 ;
        RECT 34.540 65.810 34.870 66.070 ;
        RECT 33.400 65.730 33.640 65.780 ;
        RECT 32.540 65.540 33.640 65.730 ;
        RECT 32.540 65.440 32.710 65.540 ;
        RECT 32.440 64.980 32.710 65.440 ;
      LAYER mcon ;
        RECT 34.620 65.860 34.790 66.030 ;
        RECT 33.440 65.580 33.610 65.750 ;
        RECT 31.480 65.060 31.650 65.360 ;
        RECT 32.440 65.060 32.610 65.360 ;
      LAYER met1 ;
        RECT 34.540 66.060 34.870 66.070 ;
        RECT 34.480 66.050 36.070 66.060 ;
        RECT 33.460 66.020 36.070 66.050 ;
        RECT 33.460 65.880 40.050 66.020 ;
        RECT 33.460 65.870 34.870 65.880 ;
        RECT 33.460 65.810 33.640 65.870 ;
        RECT 34.540 65.810 34.870 65.870 ;
        RECT 33.400 65.520 33.640 65.810 ;
        RECT 31.450 65.280 31.680 65.420 ;
        RECT 32.410 65.280 32.640 65.420 ;
        RECT 31.450 65.140 32.640 65.280 ;
        RECT 31.450 65.000 31.680 65.140 ;
        RECT 32.410 65.000 32.640 65.140 ;
    END
  END latch_q
  OBS
      LAYER li1 ;
        RECT 15.320 74.490 18.120 74.690 ;
        RECT 15.320 73.890 15.870 74.490 ;
        RECT 15.320 73.690 18.120 73.890 ;
        RECT 15.320 73.090 15.870 73.690 ;
        RECT 18.870 73.140 19.070 74.690 ;
        RECT 19.670 73.140 19.870 74.690 ;
        RECT 20.470 73.140 20.670 74.690 ;
        RECT 21.270 73.140 21.470 74.690 ;
        RECT 22.070 73.140 22.270 74.690 ;
        RECT 22.870 73.140 23.070 74.690 ;
        RECT 23.670 73.140 23.870 74.690 ;
        RECT 24.470 73.140 24.670 74.690 ;
        RECT 25.270 73.140 25.470 74.690 ;
        RECT 26.070 73.140 26.270 74.690 ;
        RECT 26.870 73.140 27.070 74.690 ;
        RECT 27.670 73.140 27.870 74.690 ;
        RECT 28.470 73.140 28.670 74.690 ;
        RECT 29.270 73.140 29.470 74.690 ;
        RECT 30.070 73.140 30.270 74.690 ;
        RECT 30.870 73.140 31.070 74.690 ;
        RECT 31.820 74.490 34.620 74.690 ;
        RECT 34.070 73.890 34.620 74.490 ;
        RECT 31.820 73.690 34.620 73.890 ;
        RECT 18.870 73.090 31.070 73.140 ;
        RECT 34.070 73.090 34.620 73.690 ;
        RECT 15.320 72.790 34.620 73.090 ;
        RECT 15.320 72.190 15.870 72.790 ;
        RECT 18.870 72.740 31.070 72.790 ;
        RECT 15.320 71.990 18.120 72.190 ;
        RECT 15.320 71.390 15.870 71.990 ;
        RECT 15.320 71.190 18.120 71.390 ;
        RECT 18.870 71.190 19.070 72.740 ;
        RECT 19.670 71.190 19.870 72.740 ;
        RECT 20.470 71.190 20.670 72.740 ;
        RECT 21.270 71.190 21.470 72.740 ;
        RECT 22.070 71.190 22.270 72.740 ;
        RECT 22.870 71.190 23.070 72.740 ;
        RECT 23.670 71.190 23.870 72.740 ;
        RECT 24.470 71.240 24.670 72.740 ;
        RECT 25.270 71.240 25.470 72.740 ;
        RECT 26.070 71.190 26.270 72.740 ;
        RECT 26.870 71.190 27.070 72.740 ;
        RECT 27.670 71.190 27.870 72.740 ;
        RECT 28.470 71.190 28.670 72.740 ;
        RECT 29.270 71.190 29.470 72.740 ;
        RECT 30.070 71.190 30.270 72.740 ;
        RECT 30.870 71.190 31.070 72.740 ;
        RECT 34.070 72.190 34.620 72.790 ;
        RECT 31.820 71.990 34.620 72.190 ;
        RECT 34.070 71.390 34.620 71.990 ;
        RECT 31.820 71.190 34.620 71.390 ;
        RECT 17.320 66.090 17.490 66.930 ;
        RECT 18.280 66.090 18.450 66.930 ;
        RECT 17.320 65.920 18.450 66.090 ;
        RECT 19.240 66.090 19.410 66.930 ;
        RECT 20.200 66.090 20.370 66.930 ;
        RECT 21.320 66.290 22.270 67.240 ;
        RECT 22.500 66.850 23.630 67.020 ;
        RECT 19.240 65.920 20.370 66.090 ;
        RECT 16.300 65.620 16.630 65.910 ;
        RECT 14.540 63.400 14.960 63.430 ;
        RECT 15.710 63.400 16.130 63.430 ;
        RECT 14.520 63.210 14.980 63.400 ;
        RECT 15.690 63.210 16.150 63.400 ;
        RECT 14.520 62.310 14.980 62.480 ;
        RECT 15.690 62.310 16.150 62.480 ;
        RECT 14.540 62.070 14.960 62.310 ;
        RECT 15.270 62.070 15.540 62.120 ;
        RECT 14.540 61.840 15.540 62.070 ;
        RECT 14.540 61.670 14.960 61.840 ;
        RECT 15.270 61.790 15.540 61.840 ;
        RECT 15.710 62.070 16.130 62.310 ;
        RECT 16.400 62.070 16.630 65.620 ;
        RECT 17.320 64.800 17.490 65.920 ;
        RECT 18.210 64.800 18.450 65.100 ;
        RECT 17.320 64.630 18.450 64.800 ;
        RECT 15.710 61.920 16.630 62.070 ;
        RECT 16.840 62.150 17.010 64.360 ;
        RECT 17.320 62.320 17.490 64.630 ;
        RECT 17.800 62.150 17.970 64.360 ;
        RECT 18.280 62.320 18.450 64.630 ;
        RECT 19.240 64.810 19.410 65.920 ;
        RECT 19.240 64.640 21.620 64.810 ;
        RECT 18.760 62.150 18.930 64.360 ;
        RECT 19.240 62.320 19.410 64.640 ;
        RECT 19.720 62.150 19.890 64.360 ;
        RECT 20.200 62.320 20.370 64.640 ;
        RECT 20.680 62.150 20.850 64.360 ;
        RECT 21.240 64.190 21.620 64.640 ;
        RECT 21.850 64.360 22.230 66.290 ;
        RECT 21.240 63.130 22.230 64.190 ;
        RECT 22.500 64.050 22.670 66.850 ;
        RECT 22.980 64.390 23.150 66.680 ;
        RECT 23.460 64.640 23.630 66.850 ;
        RECT 26.680 66.850 27.810 67.020 ;
        RECT 24.590 64.390 24.760 66.680 ;
        RECT 22.980 64.220 24.760 64.390 ;
        RECT 25.550 64.390 25.720 66.680 ;
        RECT 26.680 64.640 26.850 66.850 ;
        RECT 27.160 64.390 27.330 66.680 ;
        RECT 25.550 64.220 27.330 64.390 ;
        RECT 27.640 65.950 27.810 66.850 ;
        RECT 27.640 65.260 28.630 65.950 ;
        RECT 28.800 65.900 28.970 67.330 ;
        RECT 28.800 65.560 29.590 65.900 ;
        RECT 29.760 65.720 29.930 67.330 ;
        RECT 31.480 67.260 31.810 67.520 ;
        RECT 33.960 67.260 34.290 67.520 ;
        RECT 31.960 66.250 32.130 67.090 ;
        RECT 32.920 66.250 33.090 67.090 ;
        RECT 34.440 66.250 34.610 67.090 ;
        RECT 35.400 66.250 35.570 67.090 ;
        RECT 30.300 65.720 30.600 65.770 ;
        RECT 27.640 64.050 27.810 65.260 ;
        RECT 28.800 64.660 28.970 65.560 ;
        RECT 29.760 65.530 30.670 65.720 ;
        RECT 29.760 64.660 29.930 65.530 ;
        RECT 30.300 65.470 30.600 65.530 ;
        RECT 22.420 63.880 24.480 64.050 ;
        RECT 24.660 63.880 27.870 64.050 ;
        RECT 24.310 63.710 24.480 63.880 ;
        RECT 24.310 63.540 25.660 63.710 ;
        RECT 16.840 61.970 20.850 62.150 ;
        RECT 15.710 61.840 16.670 61.920 ;
        RECT 15.710 61.670 16.130 61.840 ;
        RECT 14.520 61.500 14.980 61.670 ;
        RECT 15.690 61.500 16.150 61.670 ;
        RECT 16.340 61.650 16.670 61.840 ;
        RECT 14.540 61.470 14.960 61.500 ;
        RECT 15.710 61.470 16.130 61.500 ;
        RECT 16.840 61.020 17.010 61.970 ;
        RECT 17.800 61.020 17.970 61.970 ;
        RECT 18.760 61.020 18.930 61.970 ;
        RECT 19.720 61.020 19.890 61.970 ;
        RECT 20.680 61.020 20.850 61.970 ;
        RECT 21.850 61.840 22.230 63.130 ;
        RECT 21.820 60.890 22.770 61.840 ;
        RECT 24.590 60.990 24.760 63.540 ;
        RECT 25.880 63.370 26.050 63.880 ;
        RECT 25.550 63.200 26.050 63.370 ;
        RECT 26.930 63.210 27.540 63.550 ;
        RECT 25.550 60.990 25.720 63.200 ;
        RECT 28.800 62.740 28.970 63.640 ;
        RECT 29.760 62.770 29.930 63.640 ;
        RECT 30.320 62.770 30.620 62.820 ;
        RECT 28.800 62.400 29.590 62.740 ;
        RECT 29.760 62.580 30.680 62.770 ;
        RECT 28.800 60.970 28.970 62.400 ;
        RECT 29.760 60.970 29.930 62.580 ;
        RECT 30.320 62.520 30.620 62.580 ;
        RECT 31.300 61.060 31.540 64.730 ;
        RECT 31.710 62.280 31.950 64.260 ;
        RECT 32.860 62.250 33.190 62.510 ;
        RECT 32.760 61.230 32.930 62.070 ;
        RECT 33.720 61.230 33.890 62.070 ;
        RECT 31.300 60.800 32.610 61.060 ;
        RECT 23.180 60.400 23.900 60.670 ;
        RECT 15.320 56.540 18.120 56.740 ;
        RECT 15.320 55.940 15.870 56.540 ;
        RECT 15.320 55.740 18.120 55.940 ;
        RECT 15.320 55.140 15.870 55.740 ;
        RECT 18.870 55.190 19.070 56.740 ;
        RECT 19.670 55.190 19.870 56.740 ;
        RECT 20.470 55.190 20.670 56.740 ;
        RECT 21.270 55.190 21.470 56.740 ;
        RECT 22.070 55.190 22.270 56.740 ;
        RECT 22.870 55.190 23.070 56.740 ;
        RECT 23.670 55.190 23.870 56.740 ;
        RECT 24.470 55.190 24.670 56.740 ;
        RECT 25.270 55.190 25.470 56.740 ;
        RECT 26.070 55.190 26.270 56.740 ;
        RECT 26.870 55.190 27.070 56.740 ;
        RECT 27.670 55.190 27.870 56.740 ;
        RECT 28.470 55.190 28.670 56.740 ;
        RECT 29.270 55.190 29.470 56.740 ;
        RECT 30.070 55.190 30.270 56.740 ;
        RECT 30.870 55.190 31.070 56.740 ;
        RECT 31.820 56.540 34.620 56.740 ;
        RECT 34.070 55.940 34.620 56.540 ;
        RECT 31.820 55.740 34.620 55.940 ;
        RECT 18.870 55.140 31.070 55.190 ;
        RECT 34.070 55.140 34.620 55.740 ;
        RECT 15.320 54.840 34.620 55.140 ;
        RECT 15.320 54.240 15.870 54.840 ;
        RECT 18.870 54.790 31.070 54.840 ;
        RECT 15.320 54.040 18.120 54.240 ;
        RECT 15.320 53.440 15.870 54.040 ;
        RECT 15.320 53.240 18.120 53.440 ;
        RECT 18.870 53.240 19.070 54.790 ;
        RECT 19.670 53.240 19.870 54.790 ;
        RECT 20.470 53.240 20.670 54.790 ;
        RECT 21.270 53.240 21.470 54.790 ;
        RECT 22.070 53.240 22.270 54.790 ;
        RECT 22.870 53.240 23.070 54.790 ;
        RECT 23.670 53.240 23.870 54.790 ;
        RECT 24.470 53.290 24.670 54.790 ;
        RECT 25.270 53.290 25.470 54.790 ;
        RECT 26.070 53.240 26.270 54.790 ;
        RECT 26.870 53.240 27.070 54.790 ;
        RECT 27.670 53.240 27.870 54.790 ;
        RECT 28.470 53.240 28.670 54.790 ;
        RECT 29.270 53.240 29.470 54.790 ;
        RECT 30.070 53.240 30.270 54.790 ;
        RECT 30.870 53.240 31.070 54.790 ;
        RECT 34.070 54.240 34.620 54.840 ;
        RECT 31.820 54.040 34.620 54.240 ;
        RECT 34.070 53.440 34.620 54.040 ;
        RECT 31.820 53.240 34.620 53.440 ;
      LAYER mcon ;
        RECT 15.420 73.540 15.670 73.790 ;
        RECT 15.420 73.090 15.670 73.340 ;
        RECT 34.270 73.490 34.520 73.740 ;
        RECT 34.270 73.040 34.520 73.290 ;
        RECT 15.420 72.590 15.670 72.840 ;
        RECT 15.420 72.140 15.670 72.390 ;
        RECT 34.270 72.540 34.520 72.790 ;
        RECT 34.270 72.090 34.520 72.340 ;
        RECT 21.420 66.390 22.170 67.140 ;
        RECT 14.600 63.220 14.900 63.390 ;
        RECT 15.770 63.220 16.070 63.390 ;
        RECT 14.600 62.310 14.900 62.480 ;
        RECT 15.770 62.310 16.070 62.480 ;
        RECT 15.350 61.870 15.520 62.040 ;
        RECT 18.240 64.890 18.420 65.070 ;
        RECT 21.950 65.240 22.130 65.420 ;
        RECT 21.950 64.870 22.130 65.050 ;
        RECT 21.950 64.500 22.130 64.680 ;
        RECT 21.950 63.950 22.130 64.130 ;
        RECT 28.420 65.700 28.600 65.870 ;
        RECT 28.420 65.340 28.600 65.510 ;
        RECT 34.040 67.320 34.210 67.490 ;
        RECT 30.330 65.530 30.510 65.710 ;
        RECT 21.950 63.570 22.130 63.750 ;
        RECT 21.950 63.200 22.130 63.380 ;
        RECT 21.920 60.990 22.670 61.740 ;
        RECT 26.960 63.290 27.140 63.470 ;
        RECT 27.330 63.290 27.510 63.470 ;
        RECT 30.360 62.580 30.530 62.760 ;
        RECT 31.330 62.640 31.510 62.820 ;
        RECT 31.740 64.020 31.920 64.200 ;
        RECT 31.740 62.340 31.920 62.520 ;
        RECT 32.940 62.290 33.110 62.460 ;
        RECT 23.260 60.450 23.430 60.620 ;
        RECT 23.650 60.450 23.820 60.620 ;
        RECT 15.420 55.590 15.670 55.840 ;
        RECT 15.420 55.140 15.670 55.390 ;
        RECT 34.270 55.540 34.520 55.790 ;
        RECT 34.270 55.090 34.520 55.340 ;
        RECT 15.420 54.640 15.670 54.890 ;
        RECT 15.420 54.190 15.670 54.440 ;
        RECT 34.270 54.590 34.520 54.840 ;
        RECT 34.270 54.140 34.520 54.390 ;
      LAYER met1 ;
        RECT 19.720 75.690 30.220 76.890 ;
        RECT 24.670 75.240 25.270 75.690 ;
        RECT 19.070 75.090 30.870 75.240 ;
        RECT 14.120 73.240 15.770 73.890 ;
        RECT 16.220 73.240 16.370 74.740 ;
        RECT 16.820 73.240 16.970 74.740 ;
        RECT 17.420 73.240 17.570 74.740 ;
        RECT 18.020 73.240 18.170 74.740 ;
        RECT 24.670 74.640 25.270 75.090 ;
        RECT 19.070 74.490 30.870 74.640 ;
        RECT 24.670 74.040 25.270 74.490 ;
        RECT 19.070 73.890 30.870 74.040 ;
        RECT 24.670 73.440 25.270 73.890 ;
        RECT 19.070 73.290 30.870 73.440 ;
        RECT 14.120 73.140 18.170 73.240 ;
        RECT 24.670 73.140 25.270 73.290 ;
        RECT 31.770 73.240 31.920 74.740 ;
        RECT 32.370 73.240 32.520 74.740 ;
        RECT 32.970 73.240 33.120 74.740 ;
        RECT 33.570 73.240 33.720 74.740 ;
        RECT 34.170 73.240 35.820 73.840 ;
        RECT 31.770 73.140 35.820 73.240 ;
        RECT 14.120 72.440 35.820 73.140 ;
        RECT 14.120 72.040 15.770 72.440 ;
        RECT 16.220 71.140 16.370 72.440 ;
        RECT 16.820 71.140 16.970 72.440 ;
        RECT 17.420 71.140 17.570 72.440 ;
        RECT 18.020 71.140 18.170 72.440 ;
        RECT 24.670 71.990 25.270 72.440 ;
        RECT 19.070 71.840 30.870 71.990 ;
        RECT 24.670 71.390 25.270 71.840 ;
        RECT 19.070 71.240 30.870 71.390 ;
        RECT 24.670 70.790 25.270 71.240 ;
        RECT 31.770 71.140 31.920 72.440 ;
        RECT 32.370 71.140 32.520 72.440 ;
        RECT 32.970 71.140 33.120 72.440 ;
        RECT 33.570 71.140 33.720 72.440 ;
        RECT 34.170 71.990 35.820 72.440 ;
        RECT 19.070 70.640 30.870 70.790 ;
        RECT 24.670 70.190 25.270 70.640 ;
        RECT 19.720 68.990 30.220 70.190 ;
        RECT 30.600 67.520 31.820 67.550 ;
        RECT 30.600 67.380 34.270 67.520 ;
        RECT 21.320 66.290 22.270 67.240 ;
        RECT 18.180 65.080 18.450 65.100 ;
        RECT 21.890 65.080 22.190 65.470 ;
        RECT 28.350 65.250 28.630 65.950 ;
        RECT 30.600 65.770 30.780 67.380 ;
        RECT 33.960 67.290 34.270 67.380 ;
        RECT 30.300 65.470 30.780 65.770 ;
        RECT 18.180 65.010 22.190 65.080 ;
        RECT 18.170 64.820 22.190 65.010 ;
        RECT 21.890 64.470 22.190 64.820 ;
        RECT 30.600 64.260 30.780 65.470 ;
        RECT 14.560 62.250 14.950 63.460 ;
        RECT 15.730 62.250 16.120 63.460 ;
        RECT 21.890 63.390 22.190 64.160 ;
        RECT 30.600 64.070 31.950 64.260 ;
        RECT 31.710 63.960 31.950 64.070 ;
        RECT 26.910 63.390 27.560 63.550 ;
        RECT 21.890 63.210 27.560 63.390 ;
        RECT 21.890 63.170 22.190 63.210 ;
        RECT 30.320 62.770 30.620 62.820 ;
        RECT 31.300 62.770 31.540 62.880 ;
        RECT 30.320 62.580 31.540 62.770 ;
        RECT 30.320 62.520 30.620 62.580 ;
        RECT 31.710 62.450 31.950 62.580 ;
        RECT 32.860 62.450 33.190 62.510 ;
        RECT 31.710 62.270 33.190 62.450 ;
        RECT 31.710 62.260 32.200 62.270 ;
        RECT 32.860 62.250 33.190 62.270 ;
        RECT 15.270 61.950 15.550 62.120 ;
        RECT 15.270 61.790 16.570 61.950 ;
        RECT 16.360 60.670 16.570 61.790 ;
        RECT 21.820 60.890 22.770 61.840 ;
        RECT 16.360 60.400 23.900 60.670 ;
        RECT 19.720 57.740 30.220 58.940 ;
        RECT 24.670 57.290 25.270 57.740 ;
        RECT 19.070 57.140 30.870 57.290 ;
        RECT 14.120 55.290 15.770 55.940 ;
        RECT 16.220 55.290 16.370 56.790 ;
        RECT 16.820 55.290 16.970 56.790 ;
        RECT 17.420 55.290 17.570 56.790 ;
        RECT 18.020 55.290 18.170 56.790 ;
        RECT 24.670 56.690 25.270 57.140 ;
        RECT 19.070 56.540 30.870 56.690 ;
        RECT 24.670 56.090 25.270 56.540 ;
        RECT 19.070 55.940 30.870 56.090 ;
        RECT 24.670 55.490 25.270 55.940 ;
        RECT 19.070 55.340 30.870 55.490 ;
        RECT 14.120 55.190 18.170 55.290 ;
        RECT 24.670 55.190 25.270 55.340 ;
        RECT 31.770 55.290 31.920 56.790 ;
        RECT 32.370 55.290 32.520 56.790 ;
        RECT 32.970 55.290 33.120 56.790 ;
        RECT 33.570 55.290 33.720 56.790 ;
        RECT 34.170 55.290 35.820 55.890 ;
        RECT 31.770 55.190 35.820 55.290 ;
        RECT 14.120 54.490 35.820 55.190 ;
        RECT 14.120 54.090 15.770 54.490 ;
        RECT 16.220 53.190 16.370 54.490 ;
        RECT 16.820 53.190 16.970 54.490 ;
        RECT 17.420 53.190 17.570 54.490 ;
        RECT 18.020 53.190 18.170 54.490 ;
        RECT 24.670 54.040 25.270 54.490 ;
        RECT 19.070 53.890 30.870 54.040 ;
        RECT 24.670 53.440 25.270 53.890 ;
        RECT 19.070 53.290 30.870 53.440 ;
        RECT 24.670 52.840 25.270 53.290 ;
        RECT 31.770 53.190 31.920 54.490 ;
        RECT 32.370 53.190 32.520 54.490 ;
        RECT 32.970 53.190 33.120 54.490 ;
        RECT 33.570 53.190 33.720 54.490 ;
        RECT 34.170 54.040 35.820 54.490 ;
        RECT 19.070 52.690 30.870 52.840 ;
        RECT 24.670 52.240 25.270 52.690 ;
        RECT 19.720 51.040 30.220 52.240 ;
      LAYER via ;
        RECT 19.820 75.790 20.820 76.790 ;
        RECT 20.920 75.790 21.920 76.790 ;
        RECT 24.520 75.790 25.420 76.790 ;
        RECT 28.020 75.790 29.020 76.790 ;
        RECT 29.120 75.790 30.120 76.790 ;
        RECT 14.220 73.190 15.220 73.740 ;
        RECT 34.720 73.190 35.720 73.740 ;
        RECT 14.220 72.140 15.220 72.690 ;
        RECT 34.720 72.140 35.720 72.690 ;
        RECT 19.820 69.090 20.820 70.090 ;
        RECT 20.920 69.090 21.920 70.090 ;
        RECT 24.520 69.090 25.420 70.090 ;
        RECT 28.020 69.090 29.020 70.090 ;
        RECT 29.120 69.090 30.120 70.090 ;
        RECT 21.420 66.390 22.170 67.140 ;
        RECT 21.920 60.990 22.670 61.740 ;
        RECT 19.820 57.840 20.820 58.840 ;
        RECT 20.920 57.840 21.920 58.840 ;
        RECT 24.520 57.840 25.420 58.840 ;
        RECT 28.020 57.840 29.020 58.840 ;
        RECT 29.120 57.840 30.120 58.840 ;
        RECT 14.220 55.240 15.220 55.790 ;
        RECT 34.720 55.240 35.720 55.790 ;
        RECT 14.220 54.190 15.220 54.740 ;
        RECT 34.720 54.190 35.720 54.740 ;
        RECT 19.820 51.140 20.820 52.140 ;
        RECT 20.920 51.140 21.920 52.140 ;
        RECT 24.520 51.140 25.420 52.140 ;
        RECT 28.020 51.140 29.020 52.140 ;
        RECT 29.120 51.140 30.120 52.140 ;
      LAYER met2 ;
        RECT 19.720 75.490 30.220 76.890 ;
        RECT 16.220 74.890 33.720 75.490 ;
        RECT 18.220 74.440 18.520 74.890 ;
        RECT 16.220 74.290 18.520 74.440 ;
        RECT 18.220 73.840 18.520 74.290 ;
        RECT 14.120 72.040 15.320 73.840 ;
        RECT 16.220 73.690 18.520 73.840 ;
        RECT 18.220 73.240 18.520 73.690 ;
        RECT 18.970 73.240 19.120 74.890 ;
        RECT 19.570 73.240 19.720 74.890 ;
        RECT 20.170 73.240 20.320 74.890 ;
        RECT 20.770 73.240 20.920 74.890 ;
        RECT 21.370 73.240 21.520 74.890 ;
        RECT 21.970 73.240 22.120 74.890 ;
        RECT 22.570 73.240 22.720 74.890 ;
        RECT 23.170 73.240 23.320 74.890 ;
        RECT 23.770 73.240 23.920 74.890 ;
        RECT 24.370 73.240 24.520 74.890 ;
        RECT 25.420 73.240 25.570 74.890 ;
        RECT 26.020 73.240 26.170 74.890 ;
        RECT 26.620 73.240 26.770 74.890 ;
        RECT 27.220 73.240 27.370 74.890 ;
        RECT 27.820 73.240 27.970 74.890 ;
        RECT 28.420 73.240 28.570 74.890 ;
        RECT 29.020 73.240 29.170 74.890 ;
        RECT 29.620 73.240 29.770 74.890 ;
        RECT 30.220 73.240 30.370 74.890 ;
        RECT 30.820 73.240 30.970 74.890 ;
        RECT 31.420 74.440 31.720 74.890 ;
        RECT 31.420 74.290 33.720 74.440 ;
        RECT 31.420 73.840 31.720 74.290 ;
        RECT 31.420 73.690 33.720 73.840 ;
        RECT 31.420 73.240 31.720 73.690 ;
        RECT 18.220 72.190 18.520 72.640 ;
        RECT 16.220 72.040 18.520 72.190 ;
        RECT 18.220 71.590 18.520 72.040 ;
        RECT 16.220 71.440 18.520 71.590 ;
        RECT 18.220 70.990 18.520 71.440 ;
        RECT 18.970 70.990 19.120 72.640 ;
        RECT 19.570 70.990 19.720 72.640 ;
        RECT 20.170 70.990 20.320 72.640 ;
        RECT 20.770 70.990 20.920 72.640 ;
        RECT 21.370 70.990 21.520 72.640 ;
        RECT 21.970 70.990 22.120 72.640 ;
        RECT 22.570 70.990 22.720 72.640 ;
        RECT 23.170 70.990 23.320 72.640 ;
        RECT 23.770 70.990 23.920 72.640 ;
        RECT 24.370 70.990 24.520 72.640 ;
        RECT 25.420 70.990 25.570 72.640 ;
        RECT 26.020 70.990 26.170 72.640 ;
        RECT 26.620 70.990 26.770 72.640 ;
        RECT 27.220 70.990 27.370 72.640 ;
        RECT 27.820 70.990 27.970 72.640 ;
        RECT 28.420 70.990 28.570 72.640 ;
        RECT 29.020 70.990 29.170 72.640 ;
        RECT 29.620 70.990 29.770 72.640 ;
        RECT 30.220 70.990 30.370 72.640 ;
        RECT 30.820 70.990 30.970 72.640 ;
        RECT 31.420 72.190 31.720 72.640 ;
        RECT 31.420 72.040 33.720 72.190 ;
        RECT 34.620 72.040 35.820 73.840 ;
        RECT 31.420 71.590 31.720 72.040 ;
        RECT 31.420 71.440 33.720 71.590 ;
        RECT 31.420 70.990 31.720 71.440 ;
        RECT 16.220 70.390 33.720 70.990 ;
        RECT 19.720 68.990 30.220 70.390 ;
        RECT 21.320 66.290 22.270 68.990 ;
        RECT 21.820 58.940 22.770 61.840 ;
        RECT 19.720 57.540 30.220 58.940 ;
        RECT 16.220 56.940 33.720 57.540 ;
        RECT 18.220 56.490 18.520 56.940 ;
        RECT 16.220 56.340 18.520 56.490 ;
        RECT 18.220 55.890 18.520 56.340 ;
        RECT 14.120 54.090 15.320 55.890 ;
        RECT 16.220 55.740 18.520 55.890 ;
        RECT 18.220 55.290 18.520 55.740 ;
        RECT 18.970 55.290 19.120 56.940 ;
        RECT 19.570 55.290 19.720 56.940 ;
        RECT 20.170 55.290 20.320 56.940 ;
        RECT 20.770 55.290 20.920 56.940 ;
        RECT 21.370 55.290 21.520 56.940 ;
        RECT 21.970 55.290 22.120 56.940 ;
        RECT 22.570 55.290 22.720 56.940 ;
        RECT 23.170 55.290 23.320 56.940 ;
        RECT 23.770 55.290 23.920 56.940 ;
        RECT 24.370 55.290 24.520 56.940 ;
        RECT 25.420 55.290 25.570 56.940 ;
        RECT 26.020 55.290 26.170 56.940 ;
        RECT 26.620 55.290 26.770 56.940 ;
        RECT 27.220 55.290 27.370 56.940 ;
        RECT 27.820 55.290 27.970 56.940 ;
        RECT 28.420 55.290 28.570 56.940 ;
        RECT 29.020 55.290 29.170 56.940 ;
        RECT 29.620 55.290 29.770 56.940 ;
        RECT 30.220 55.290 30.370 56.940 ;
        RECT 30.820 55.290 30.970 56.940 ;
        RECT 31.420 56.490 31.720 56.940 ;
        RECT 31.420 56.340 33.720 56.490 ;
        RECT 31.420 55.890 31.720 56.340 ;
        RECT 31.420 55.740 33.720 55.890 ;
        RECT 31.420 55.290 31.720 55.740 ;
        RECT 18.220 54.240 18.520 54.690 ;
        RECT 16.220 54.090 18.520 54.240 ;
        RECT 18.220 53.640 18.520 54.090 ;
        RECT 16.220 53.490 18.520 53.640 ;
        RECT 18.220 53.040 18.520 53.490 ;
        RECT 18.970 53.040 19.120 54.690 ;
        RECT 19.570 53.040 19.720 54.690 ;
        RECT 20.170 53.040 20.320 54.690 ;
        RECT 20.770 53.040 20.920 54.690 ;
        RECT 21.370 53.040 21.520 54.690 ;
        RECT 21.970 53.040 22.120 54.690 ;
        RECT 22.570 53.040 22.720 54.690 ;
        RECT 23.170 53.040 23.320 54.690 ;
        RECT 23.770 53.040 23.920 54.690 ;
        RECT 24.370 53.040 24.520 54.690 ;
        RECT 25.420 53.040 25.570 54.690 ;
        RECT 26.020 53.040 26.170 54.690 ;
        RECT 26.620 53.040 26.770 54.690 ;
        RECT 27.220 53.040 27.370 54.690 ;
        RECT 27.820 53.040 27.970 54.690 ;
        RECT 28.420 53.040 28.570 54.690 ;
        RECT 29.020 53.040 29.170 54.690 ;
        RECT 29.620 53.040 29.770 54.690 ;
        RECT 30.220 53.040 30.370 54.690 ;
        RECT 30.820 53.040 30.970 54.690 ;
        RECT 31.420 54.240 31.720 54.690 ;
        RECT 31.420 54.090 33.720 54.240 ;
        RECT 34.620 54.090 35.820 55.890 ;
        RECT 31.420 53.640 31.720 54.090 ;
        RECT 31.420 53.490 33.720 53.640 ;
        RECT 31.420 53.040 31.720 53.490 ;
        RECT 16.220 52.440 33.720 53.040 ;
        RECT 19.720 51.040 30.220 52.440 ;
  END
END adc_comp_latch
END LIBRARY

