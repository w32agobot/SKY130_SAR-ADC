magic
tech sky130A
timestamp 1659617841
<< metal2 >>
rect -416 1916 -384 1970
rect 1885 1916 1917 1953
rect 2094 1916 2126 1970
rect 4395 1916 4427 1953
rect 4604 1916 4636 1970
rect 6905 1916 6937 1953
rect 7114 1916 7146 1970
rect 9415 1916 9447 1953
rect -502 1886 9478 1916
rect -416 1885 1917 1886
rect -502 1817 -433 1847
rect -416 122 -384 1885
rect 476 1161 529 1194
rect 979 1168 1032 1201
rect 303 987 331 1037
rect 804 981 832 1031
rect 1328 984 1356 1034
rect 472 673 525 706
rect 971 675 1024 708
rect 804 510 846 554
rect 469 301 579 331
rect 958 300 1068 330
rect 1885 122 1917 1885
rect 2094 1885 4427 1886
rect 2008 1817 2077 1847
rect 2094 122 2126 1885
rect 2938 1172 3778 1195
rect 2816 983 2837 1041
rect 3184 683 3204 1054
rect 3688 977 3709 1035
rect 2930 660 3770 683
rect 3184 463 3204 660
rect 4395 122 4427 1885
rect 4604 1885 6937 1886
rect 4518 1817 4587 1847
rect 4604 122 4636 1885
rect 5480 1165 5568 1197
rect 5977 1165 6065 1197
rect 5324 977 5345 1035
rect 5681 972 5702 1030
rect 6195 970 6216 1028
rect 5486 662 5551 681
rect 5981 675 6069 707
rect 5686 538 5707 548
rect 5679 473 5707 538
rect 6905 122 6937 1885
rect 7114 1885 9447 1886
rect 7028 1817 7097 1847
rect 7114 122 7146 1885
rect 7990 1185 8078 1217
rect 8500 1167 8588 1199
rect 8200 966 8226 1052
rect 8701 972 8727 1058
rect 7999 668 8087 700
rect 8500 677 8588 709
rect 8194 461 8220 547
rect 9415 122 9447 1885
rect -416 93 414 122
rect 1142 93 1970 122
rect 2094 93 2924 122
rect 3652 93 4480 122
rect 4604 93 5434 122
rect 6162 93 6990 122
rect 7114 93 7944 122
rect 8672 93 9500 122
rect -416 68 -384 93
rect 1885 51 1917 93
rect 2094 68 2126 93
rect 4395 51 4427 93
rect 4604 68 4636 93
rect 6905 51 6937 93
rect 7114 68 7146 93
rect 9415 51 9447 93
<< metal4 >>
rect -411 1917 -381 1973
rect -502 1916 -381 1917
rect 1885 1916 1917 1953
rect 2099 1917 2129 1973
rect 2008 1916 2129 1917
rect 4395 1916 4427 1953
rect 4609 1917 4639 1973
rect 4518 1916 4639 1917
rect 6905 1916 6937 1953
rect 7119 1917 7149 1973
rect 7028 1916 7149 1917
rect 9415 1916 9447 1953
rect -502 1886 9496 1916
rect -411 56 -381 1886
rect 92 1471 122 1506
rect 380 1471 410 1506
rect 594 1471 624 1506
rect 882 1471 912 1506
rect 1096 1471 1126 1506
rect 1384 1471 1414 1506
rect 0 1384 71 1414
rect 466 1384 537 1414
rect 968 1384 1039 1414
rect 1435 1384 1506 1414
rect 0 1096 71 1126
rect 466 1096 537 1126
rect 968 1096 1039 1126
rect 1435 1096 1506 1126
rect 92 969 122 1039
rect 380 969 410 1039
rect 594 969 624 1039
rect 882 969 912 1039
rect 1096 969 1126 1039
rect 1384 969 1414 1039
rect 0 882 71 912
rect 466 882 537 912
rect 968 882 1039 912
rect 1435 882 1506 912
rect 0 594 71 624
rect 466 594 537 624
rect 969 594 1040 624
rect 1435 594 1506 624
rect 92 502 122 537
rect 380 502 410 537
rect 594 500 624 537
rect 882 500 912 537
rect 1096 502 1126 537
rect 1384 502 1414 537
rect 462 380 572 410
rect 950 380 1062 410
rect -158 92 155 122
rect 1313 121 1765 122
rect 1296 92 1765 121
rect 1885 51 1917 1886
rect 2099 56 2129 1886
rect 2602 1471 2632 1506
rect 2890 1471 2920 1506
rect 3104 1471 3134 1506
rect 3392 1471 3422 1506
rect 3606 1471 3636 1506
rect 3894 1471 3924 1506
rect 2510 1384 2581 1414
rect 2976 1384 3047 1414
rect 3478 1384 3549 1414
rect 3945 1384 4016 1414
rect 2510 1096 2581 1126
rect 2976 1096 3047 1126
rect 3478 1096 3549 1126
rect 3945 1096 4016 1126
rect 2602 969 2632 1039
rect 2890 969 2920 1039
rect 3104 969 3134 1039
rect 3392 969 3422 1039
rect 3606 969 3636 1039
rect 3894 969 3924 1039
rect 2510 882 2581 912
rect 2976 882 3047 912
rect 3478 882 3549 912
rect 3945 882 4016 912
rect 2510 594 2581 624
rect 2976 594 3047 624
rect 3479 594 3550 624
rect 3945 594 4016 624
rect 2602 502 2632 537
rect 2890 502 2920 537
rect 3104 467 3134 537
rect 3392 467 3422 537
rect 3606 502 3636 537
rect 3894 502 3924 537
rect 3012 380 3047 410
rect 3479 380 3514 410
rect 2352 92 2665 122
rect 3823 121 4275 122
rect 3806 92 4275 121
rect 3248 9 3278 73
rect 4395 51 4427 1886
rect 4609 56 4639 1886
rect 5112 1471 5142 1506
rect 5400 1471 5430 1506
rect 5614 1471 5644 1506
rect 5902 1471 5932 1506
rect 6116 1471 6146 1506
rect 6404 1471 6434 1506
rect 5020 1384 5091 1414
rect 5486 1384 5557 1414
rect 5988 1384 6059 1414
rect 6455 1384 6526 1414
rect 5020 1096 5091 1126
rect 5486 1096 5557 1126
rect 5988 1096 6059 1126
rect 6455 1096 6526 1126
rect 5112 969 5142 1039
rect 5400 969 5430 1039
rect 5614 969 5644 1039
rect 5902 969 5932 1039
rect 6116 969 6146 1039
rect 6404 969 6434 1039
rect 5020 882 5091 912
rect 5486 882 5557 912
rect 5988 882 6059 912
rect 6455 882 6526 912
rect 5020 594 5091 624
rect 5486 594 5557 624
rect 5989 594 6060 624
rect 6455 594 6526 624
rect 5112 502 5142 537
rect 5400 502 5430 537
rect 5614 467 5644 537
rect 5902 502 5932 537
rect 6116 502 6146 537
rect 6404 502 6434 537
rect 5522 380 5557 410
rect 4862 92 5175 122
rect 6333 121 6785 122
rect 6316 92 6785 121
rect 6905 51 6937 1886
rect 7119 56 7149 1886
rect 7622 1471 7652 1506
rect 7910 1471 7940 1506
rect 8124 1471 8154 1506
rect 8412 1471 8442 1506
rect 8626 1471 8656 1506
rect 8914 1471 8944 1506
rect 7530 1384 7601 1414
rect 7996 1384 8067 1414
rect 8498 1384 8569 1414
rect 8965 1384 9036 1414
rect 7530 1096 7601 1126
rect 7996 1096 8067 1126
rect 8498 1096 8569 1126
rect 8965 1096 9036 1126
rect 7622 969 7652 1039
rect 7910 969 7940 1039
rect 8124 969 8154 1039
rect 8412 969 8442 1039
rect 8626 969 8656 1039
rect 8914 969 8944 1039
rect 7530 882 7601 912
rect 7996 882 8067 912
rect 8498 882 8569 912
rect 8965 882 9036 912
rect 7530 594 7601 624
rect 7996 594 8067 624
rect 8499 594 8570 624
rect 8965 594 9036 624
rect 7622 502 7652 537
rect 7910 502 7940 537
rect 8124 467 8154 537
rect 8412 502 8442 537
rect 8626 502 8656 537
rect 8914 502 8944 537
rect 7372 92 7685 122
rect 8843 121 9295 122
rect 8826 92 9295 121
rect 9415 51 9447 1886
rect 5757 4 5788 49
rect 8268 -2 8298 51
use adc_array_wafflecap_8(1)_25um2  adc_array_wafflecap_8(1)_25um2_0
timestamp 1659612718
transform 1 0 8032 0 1 0
box 0 0 502 502
use adc_array_wafflecap_8(2)_25um2  adc_array_wafflecap_8(2)_25um2_0
timestamp 1659612673
transform 1 0 5522 0 1 0
box 0 0 502 502
use adc_array_wafflecap_8(4)_25um2  adc_array_wafflecap_8(4)_25um2_0
timestamp 1659612633
transform 1 0 3012 0 1 0
box 0 0 502 502
use adc_array_wafflecap_8(8)_25um2  adc_array_wafflecap_8(8)_25um2_0
array 0 3 2510 0 0 2008
timestamp 1659615172
transform 1 0 0 0 1 0
box 0 0 502 502
use adc_array_wafflecap_8(8)_25um2  adc_array_wafflecap_8(8)_25um2_1
array 0 3 2510 0 0 2008
timestamp 1659615172
transform 1 0 0 0 1 502
box 0 0 502 502
use adc_array_wafflecap_8(8)_25um2  adc_array_wafflecap_8(8)_25um2_2
array 0 3 2510 0 0 2008
timestamp 1659615172
transform 1 0 0 0 1 1004
box 0 0 502 502
use adc_array_wafflecap_8(8)_25um2  adc_array_wafflecap_8(8)_25um2_3
array 0 3 2510 0 0 2008
timestamp 1659615172
transform 1 0 502 0 1 1004
box 0 0 502 502
use adc_array_wafflecap_8(8)_25um2  adc_array_wafflecap_8(8)_25um2_4
array 0 3 2510 0 0 2008
timestamp 1659615172
transform 1 0 502 0 1 502
box 0 0 502 502
use adc_array_wafflecap_8(8)_25um2  adc_array_wafflecap_8(8)_25um2_5
array 0 3 2510 0 0 2008
timestamp 1659615172
transform 1 0 1004 0 1 1004
box 0 0 502 502
use adc_array_wafflecap_8(8)_25um2  adc_array_wafflecap_8(8)_25um2_6
array 0 3 2510 0 0 2008
timestamp 1659615172
transform 1 0 1004 0 1 502
box 0 0 502 502
use adc_array_wafflecap_8(8)_25um2  adc_array_wafflecap_8(8)_25um2_7
array 0 3 2510 0 0 2008
timestamp 1659615172
transform 1 0 1004 0 1 0
box 0 0 502 502
use adc_array_wafflecap_8(8)_25um2  adc_array_wafflecap_8(8)_25um2_8
array 0 3 2510 0 0 2008
timestamp 1659615172
transform 1 0 -502 0 1 0
box 0 0 502 502
use adc_array_wafflecap_8(8)_25um2  adc_array_wafflecap_8(8)_25um2_9
array 0 3 2510 0 0 2008
timestamp 1659615172
transform 1 0 -502 0 1 502
box 0 0 502 502
use adc_array_wafflecap_8(8)_25um2  adc_array_wafflecap_8(8)_25um2_10
array 0 3 2510 0 0 2008
timestamp 1659615172
transform 1 0 -502 0 1 1004
box 0 0 502 502
use adc_array_wafflecap_8(8)_25um2  adc_array_wafflecap_8(8)_25um2_11
array 0 3 2510 0 0 2008
timestamp 1659615172
transform 1 0 -502 0 1 1506
box 0 0 502 502
use adc_array_wafflecap_8(8)_25um2  adc_array_wafflecap_8(8)_25um2_12
array 0 3 2510 0 0 2008
timestamp 1659615172
transform 1 0 0 0 1 1506
box 0 0 502 502
use adc_array_wafflecap_8(8)_25um2  adc_array_wafflecap_8(8)_25um2_13
array 0 3 2510 0 0 2008
timestamp 1659615172
transform 1 0 502 0 1 1506
box 0 0 502 502
use adc_array_wafflecap_8(8)_25um2  adc_array_wafflecap_8(8)_25um2_14
array 0 3 2510 0 0 2008
timestamp 1659615172
transform 1 0 1004 0 1 1506
box 0 0 502 502
use adc_array_wafflecap_8(8)_25um2  adc_array_wafflecap_8(8)_25um2_15
array 0 3 2510 0 0 2008
timestamp 1659615172
transform 1 0 1506 0 1 1506
box 0 0 502 502
use adc_array_wafflecap_8(8)_25um2  adc_array_wafflecap_8(8)_25um2_16
array 0 3 2510 0 0 2008
timestamp 1659615172
transform 1 0 1506 0 1 1004
box 0 0 502 502
use adc_array_wafflecap_8(8)_25um2  adc_array_wafflecap_8(8)_25um2_17
array 0 3 2510 0 0 2008
timestamp 1659615172
transform 1 0 1506 0 1 502
box 0 0 502 502
use adc_array_wafflecap_8(8)_25um2  adc_array_wafflecap_8(8)_25um2_18
array 0 3 2510 0 0 2008
timestamp 1659615172
transform 1 0 1506 0 1 0
box 0 0 502 502
use adc_array_wafflecap_8(8)_25um2  adc_array_wafflecap_8(8)_25um2_19
timestamp 1659615172
transform 1 0 502 0 1 0
box 0 0 502 502
<< labels >>
rlabel metal4 -502 1886 -502 1917 7 ctop_dummy
rlabel metal2 -502 1817 -502 1847 7 cbot_dummy
rlabel metal4 3134 495 3134 515 3 ctop_4
rlabel metal4 5644 490 5644 510 3 ctop_2
rlabel metal4 8154 491 8154 511 3 ctop_1
rlabel metal2 8220 494 8220 514 3 cbot_1
rlabel metal2 5707 493 5707 513 3 cbot_2
rlabel metal2 3204 494 3204 514 3 cbot_4
rlabel metal4 3248 9 3278 9 5 floatingmetal4
rlabel metal4 5757 4 5788 4 5 floatingmetal2
rlabel metal4 8268 -2 8298 -2 5 floatingmetal1
rlabel metal4 594 500 624 500 5 ctop_8
rlabel metal2 804 510 846 510 5 cbot_8
<< end >>
