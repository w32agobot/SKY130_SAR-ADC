* NGSPICE file created from adc_vcm_gen.ext - technology: sky130A

.subckt sky130_fd_sc_hd__inv_1 A VGND VPWR Y VNB VPB
X0 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_K25L97 a_n29_0# a_129_0# a_n129_n26# w_n224_n36# a_n187_0#
+ a_29_n26#
X0 a_129_0# a_29_n26# a_n29_0# w_n224_n36# sky130_fd_pr__pfet_01v8 ad=1.45e+11p pd=1.58e+06u as=1.45e+11p ps=1.58e+06u w=500000u l=500000u
X1 a_n29_0# a_n129_n26# a_n187_0# w_n224_n36# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.45e+11p ps=1.58e+06u w=500000u l=500000u
.ends

.subckt sky130_fd_sc_hd__buf_4 A VGND VPWR X VNB VPB
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=8e+11p pd=7.6e+06u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=5.2e+11p ps=5.5e+06u w=650000u l=150000u
X5 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X9 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__dlymetal6s6s_1 A VGND VPWR X VNB VPB
X0 X a_629_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=5.82e+11p ps=5.85e+06u w=650000u l=150000u
X1 a_523_47# a_346_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X2 VGND a_240_47# a_346_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X3 a_240_47# a_63_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X4 VPWR a_240_47# a_346_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=8.445e+11p pd=7.95e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X5 VGND A a_63_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X6 VPWR A a_63_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X7 VPWR a_523_47# a_629_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X8 VGND a_523_47# a_629_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X9 a_523_47# a_346_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X10 a_240_47# a_63_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X11 X a_629_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_8PFHMD a_n129_n76# a_n29_n50# a_n187_n50# a_29_n76#
+ a_129_n50# VSUBS
X0 a_129_n50# a_29_n76# a_n29_n50# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45e+11p pd=1.58e+06u as=1.45e+11p ps=1.58e+06u w=500000u l=500000u
X1 a_n29_n50# a_n129_n76# a_n187_n50# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.45e+11p ps=1.58e+06u w=500000u l=500000u
.ends

.subckt adc_noise_decoup_cell1 nmoscap_top nmoscap_bot mimcap_top mimcap_bot pwell
X0 mimcap_top mimcap_bot sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X1 nmoscap_bot nmoscap_top nmoscap_bot pwell sky130_fd_pr__nfet_01v8 ad=2.296e+13p pd=6.84e+07u as=0p ps=0u w=1.64e+07u l=1.6e+07u
.ends

.subckt sky130_fd_sc_hd__nand2_1 A B VGND VPWR Y VNB VPB
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=5.2e+11p pd=5.04e+06u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1 Y A a_113_47# VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X2 a_113_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X3 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt adc_vcm_generator VDD VSS clk vcm
Xsky130_fd_sc_hd__inv_1_4 clk VSS VDD sky130_fd_sc_hd__inv_1_4/Y VSS VDD sky130_fd_sc_hd__inv_1
Xsky130_fd_pr__pfet_01v8_K25L97_0 mimtop2 vcm phi1_n VDD vcm phi1_n sky130_fd_pr__pfet_01v8_K25L97
Xsky130_fd_pr__pfet_01v8_K25L97_1 mimtop1 vcm phi1_n VDD vcm phi1_n sky130_fd_pr__pfet_01v8_K25L97
Xsky130_fd_pr__pfet_01v8_K25L97_2 mimtop2 adc_noise_decoup_cell1_3[6|5]/mimcap_bot
+ phi2_n VDD adc_noise_decoup_cell1_3[6|5]/mimcap_bot phi2_n sky130_fd_pr__pfet_01v8_K25L97
Xsky130_fd_pr__pfet_01v8_K25L97_3 VDD mimtop1 phi2_n VDD mimtop1 phi2_n sky130_fd_pr__pfet_01v8_K25L97
Xsky130_fd_pr__pfet_01v8_K25L97_4 adc_noise_decoup_cell1_3[6|5]/mimcap_bot VSS phi1_n
+ VDD VSS phi1_n sky130_fd_pr__pfet_01v8_K25L97
Xsky130_fd_sc_hd__buf_4_0 sky130_fd_sc_hd__inv_1_2/A VSS VDD phi1 VSS VDD sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_1 sky130_fd_sc_hd__inv_1_2/Y VSS VDD phi1_n VSS VDD sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_2 sky130_fd_sc_hd__inv_1_3/A VSS VDD phi2 VSS VDD sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_3 sky130_fd_sc_hd__inv_1_3/Y VSS VDD phi2_n VSS VDD sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__dlymetal6s6s_1_0 sky130_fd_sc_hd__nand2_1_0/Y VSS VDD sky130_fd_sc_hd__dlymetal6s6s_1_2/A
+ VSS VDD sky130_fd_sc_hd__dlymetal6s6s_1
Xsky130_fd_sc_hd__dlymetal6s6s_1_1 sky130_fd_sc_hd__nand2_1_1/Y VSS VDD sky130_fd_sc_hd__dlymetal6s6s_1_4/A
+ VSS VDD sky130_fd_sc_hd__dlymetal6s6s_1
Xsky130_fd_sc_hd__dlymetal6s6s_1_2 sky130_fd_sc_hd__dlymetal6s6s_1_2/A VSS VDD sky130_fd_sc_hd__dlymetal6s6s_1_3/A
+ VSS VDD sky130_fd_sc_hd__dlymetal6s6s_1
Xsky130_fd_sc_hd__dlymetal6s6s_1_3 sky130_fd_sc_hd__dlymetal6s6s_1_3/A VSS VDD sky130_fd_sc_hd__inv_1_0/A
+ VSS VDD sky130_fd_sc_hd__dlymetal6s6s_1
Xsky130_fd_pr__nfet_01v8_8PFHMD_0 phi1 mimtop2 vcm phi1 vcm VSS sky130_fd_pr__nfet_01v8_8PFHMD
Xsky130_fd_sc_hd__dlymetal6s6s_1_4 sky130_fd_sc_hd__dlymetal6s6s_1_4/A VSS VDD sky130_fd_sc_hd__dlymetal6s6s_1_5/A
+ VSS VDD sky130_fd_sc_hd__dlymetal6s6s_1
Xsky130_fd_sc_hd__dlymetal6s6s_1_5 sky130_fd_sc_hd__dlymetal6s6s_1_5/A VSS VDD sky130_fd_sc_hd__inv_1_1/A
+ VSS VDD sky130_fd_sc_hd__dlymetal6s6s_1
Xsky130_fd_pr__nfet_01v8_8PFHMD_1 phi1 mimtop1 vcm phi1 vcm VSS sky130_fd_pr__nfet_01v8_8PFHMD
Xadc_noise_decoup_cell1_0[0] VDD VSS VDD VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_0[1] VDD VSS VDD VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_0[2] VDD VSS VDD VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_0[3] VDD VSS VDD VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[0|0] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[1|0] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[2|0] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[3|0] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[4|0] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[5|0] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[6|0] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[0|1] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[1|1] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[2|1] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[3|1] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[4|1] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[5|1] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[6|1] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[0|2] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[1|2] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[2|2] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[3|2] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[4|2] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[5|2] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[6|2] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[0|3] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[1|3] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[2|3] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[3|3] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[4|3] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[5|3] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[6|3] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[0|4] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[1|4] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[2|4] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[3|4] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[4|4] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[5|4] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[6|4] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[0|5] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[1|5] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[2|5] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[3|5] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[4|5] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[5|5] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[6|5] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xsky130_fd_pr__nfet_01v8_8PFHMD_2 phi2 mimtop2 adc_noise_decoup_cell1_3[6|5]/mimcap_bot
+ phi2 adc_noise_decoup_cell1_3[6|5]/mimcap_bot VSS sky130_fd_pr__nfet_01v8_8PFHMD
Xadc_noise_decoup_cell1_3[0|0] vcm VSS mimtop1 adc_noise_decoup_cell1_3[6|5]/mimcap_bot
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[1|0] vcm VSS mimtop1 adc_noise_decoup_cell1_3[6|5]/mimcap_bot
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[2|0] vcm VSS mimtop1 adc_noise_decoup_cell1_3[6|5]/mimcap_bot
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[3|0] vcm VSS mimtop1 adc_noise_decoup_cell1_3[6|5]/mimcap_bot
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[4|0] vcm VSS mimtop1 adc_noise_decoup_cell1_3[6|5]/mimcap_bot
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[5|0] vcm VSS mimtop1 adc_noise_decoup_cell1_3[6|5]/mimcap_bot
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[6|0] vcm VSS mimtop1 adc_noise_decoup_cell1_3[6|5]/mimcap_bot
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[0|1] vcm VSS mimtop1 adc_noise_decoup_cell1_3[6|5]/mimcap_bot
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[1|1] vcm VSS mimtop1 adc_noise_decoup_cell1_3[6|5]/mimcap_bot
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[2|1] vcm VSS mimtop1 adc_noise_decoup_cell1_3[6|5]/mimcap_bot
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[3|1] vcm VSS mimtop1 adc_noise_decoup_cell1_3[6|5]/mimcap_bot
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[4|1] vcm VSS mimtop1 adc_noise_decoup_cell1_3[6|5]/mimcap_bot
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[5|1] vcm VSS mimtop1 adc_noise_decoup_cell1_3[6|5]/mimcap_bot
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[6|1] vcm VSS mimtop1 adc_noise_decoup_cell1_3[6|5]/mimcap_bot
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[0|2] vcm VSS mimtop1 adc_noise_decoup_cell1_3[6|5]/mimcap_bot
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[1|2] vcm VSS mimtop1 adc_noise_decoup_cell1_3[6|5]/mimcap_bot
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[2|2] vcm VSS mimtop1 adc_noise_decoup_cell1_3[6|5]/mimcap_bot
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[3|2] vcm VSS mimtop1 adc_noise_decoup_cell1_3[6|5]/mimcap_bot
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[4|2] vcm VSS mimtop1 adc_noise_decoup_cell1_3[6|5]/mimcap_bot
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[5|2] vcm VSS mimtop1 adc_noise_decoup_cell1_3[6|5]/mimcap_bot
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[6|2] vcm VSS mimtop1 adc_noise_decoup_cell1_3[6|5]/mimcap_bot
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[0|3] vcm VSS mimtop1 adc_noise_decoup_cell1_3[6|5]/mimcap_bot
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[1|3] vcm VSS mimtop1 adc_noise_decoup_cell1_3[6|5]/mimcap_bot
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[2|3] vcm VSS mimtop1 adc_noise_decoup_cell1_3[6|5]/mimcap_bot
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[3|3] vcm VSS mimtop1 adc_noise_decoup_cell1_3[6|5]/mimcap_bot
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[4|3] vcm VSS mimtop1 adc_noise_decoup_cell1_3[6|5]/mimcap_bot
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[5|3] vcm VSS mimtop1 adc_noise_decoup_cell1_3[6|5]/mimcap_bot
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[6|3] vcm VSS mimtop1 adc_noise_decoup_cell1_3[6|5]/mimcap_bot
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[0|4] vcm VSS mimtop1 adc_noise_decoup_cell1_3[6|5]/mimcap_bot
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[1|4] vcm VSS mimtop1 adc_noise_decoup_cell1_3[6|5]/mimcap_bot
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[2|4] vcm VSS mimtop1 adc_noise_decoup_cell1_3[6|5]/mimcap_bot
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[3|4] vcm VSS mimtop1 adc_noise_decoup_cell1_3[6|5]/mimcap_bot
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[4|4] vcm VSS mimtop1 adc_noise_decoup_cell1_3[6|5]/mimcap_bot
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[5|4] vcm VSS mimtop1 adc_noise_decoup_cell1_3[6|5]/mimcap_bot
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[6|4] vcm VSS mimtop1 adc_noise_decoup_cell1_3[6|5]/mimcap_bot
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[0|5] vcm VSS mimtop1 adc_noise_decoup_cell1_3[6|5]/mimcap_bot
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[1|5] vcm VSS mimtop1 adc_noise_decoup_cell1_3[6|5]/mimcap_bot
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[2|5] vcm VSS mimtop1 adc_noise_decoup_cell1_3[6|5]/mimcap_bot
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[3|5] vcm VSS mimtop1 adc_noise_decoup_cell1_3[6|5]/mimcap_bot
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[4|5] vcm VSS mimtop1 adc_noise_decoup_cell1_3[6|5]/mimcap_bot
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[5|5] vcm VSS mimtop1 adc_noise_decoup_cell1_3[6|5]/mimcap_bot
+ VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[6|5] vcm VSS mimtop1 adc_noise_decoup_cell1_3[6|5]/mimcap_bot
+ VSS adc_noise_decoup_cell1
Xsky130_fd_pr__nfet_01v8_8PFHMD_3 phi2 VDD mimtop1 phi2 mimtop1 VSS sky130_fd_pr__nfet_01v8_8PFHMD
Xsky130_fd_pr__nfet_01v8_8PFHMD_4 phi1 adc_noise_decoup_cell1_3[6|5]/mimcap_bot VSS
+ phi1 VSS VSS sky130_fd_pr__nfet_01v8_8PFHMD
Xsky130_fd_sc_hd__nand2_1_0 clk sky130_fd_sc_hd__inv_1_3/Y VSS VDD sky130_fd_sc_hd__nand2_1_0/Y
+ VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_1 sky130_fd_sc_hd__inv_1_2/Y sky130_fd_sc_hd__inv_1_4/Y
+ VSS VDD sky130_fd_sc_hd__nand2_1_1/Y VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__inv_1_0 sky130_fd_sc_hd__inv_1_0/A VSS VDD sky130_fd_sc_hd__inv_1_2/A
+ VSS VDD sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_1 sky130_fd_sc_hd__inv_1_1/A VSS VDD sky130_fd_sc_hd__inv_1_3/A
+ VSS VDD sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_2 sky130_fd_sc_hd__inv_1_2/A VSS VDD sky130_fd_sc_hd__inv_1_2/Y
+ VSS VDD sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_3 sky130_fd_sc_hd__inv_1_3/A VSS VDD sky130_fd_sc_hd__inv_1_3/Y
+ VSS VDD sky130_fd_sc_hd__inv_1
.ends

