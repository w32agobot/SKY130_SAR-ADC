* SPICE3 file created from Extract.ext - technology: sky130A

C0 cbot_dummy ctop_2 1.88fF
C1 cbot_dummy ctop_8 1.96fF
C2 ctop_dummy cbot_1 1.80fF
C3 cbot_2 floatingmetal2 3.31fF
C4 cbot_dummy ctop_dummy 247.72fF
C5 floatingmetal4 cbot_4 2.21fF
C6 ctop_4 ctop_dummy 2.67fF
C7 cbot_dummy cbot_2 16.01fF
C8 cbot_1 floatingmetal1 3.88fF
C9 cbot_dummy cbot_8 14.65fF
C10 ctop_dummy ctop_2 2.51fF
C11 ctop_1 cbot_1 29.29fF
C12 ctop_dummy ctop_8 2.62fF
C13 cbot_2 ctop_2 29.86fF
C14 cbot_dummy ctop_1 1.83fF
C15 cbot_dummy cbot_4 16.03fF
C16 ctop_8 cbot_8 28.51fF
C17 ctop_4 cbot_4 30.99fF
C18 ctop_dummy cbot_2 1.82fF
C19 ctop_dummy cbot_8 1.57fF
C20 cbot_dummy cbot_1 15.99fF
C21 ctop_1 ctop_dummy 2.47fF
C22 ctop_dummy cbot_4 1.83fF
C23 cbot_dummy ctop_4 1.98fF
C24 cbot_1 VSUBS 3.89fF
C25 cbot_2 VSUBS 3.90fF
C26 cbot_dummy VSUBS 43.58fF
C27 cbot_8 VSUBS 3.02fF
C28 ctop_dummy VSUBS 1.54fF
C29 cbot_4 VSUBS 3.90fF
