magic
tech sky130A
timestamp 1661509002
<< nwell >>
rect 144 2605 349 2759
<< poly >>
rect 1039 2460 1078 2465
rect 1039 2443 1047 2460
rect 1064 2443 1078 2460
rect 1039 2438 1078 2443
<< polycont >>
rect 1047 2443 1064 2460
<< locali >>
rect 291 3138 399 3141
rect 291 3120 297 3138
rect 314 3120 336 3138
rect 353 3120 372 3138
rect 389 3120 399 3138
rect 291 3117 399 3120
rect 291 2759 334 3117
rect 175 2739 334 2759
rect 248 2602 275 2610
rect 248 2585 256 2602
rect 273 2585 275 2602
rect 248 2582 275 2585
rect 248 2577 273 2582
rect 1039 2460 1078 2465
rect 1039 2443 1047 2460
rect 1064 2443 1078 2460
rect 1039 2438 1078 2443
<< viali >>
rect 297 3120 314 3138
rect 336 3120 353 3138
rect 372 3120 389 3138
rect 256 2585 273 2602
rect 1047 2443 1064 2460
rect 1086 2443 1103 2460
<< metal1 >>
rect 291 3138 399 3168
rect 291 3120 297 3138
rect 314 3120 336 3138
rect 353 3120 372 3138
rect 389 3120 399 3138
rect 291 3117 399 3120
rect 128 2601 158 2610
rect -61 2587 158 2601
rect 128 2577 158 2587
rect 248 2602 276 2610
rect 248 2585 256 2602
rect 273 2593 276 2602
rect 273 2585 378 2593
rect 248 2577 378 2585
rect 355 2563 378 2577
rect 114 2423 342 2476
rect 357 2465 378 2563
rect 357 2460 1111 2465
rect 357 2443 1047 2460
rect 1064 2443 1086 2460
rect 1103 2443 1111 2460
rect 357 2438 1111 2443
use adc_comp_circuit  adc_comp_circuit_0 ../adc_comp_circuit
timestamp 1661508802
transform 1 0 358 0 1 3087
box -419 -3013 2031 2339
use inverter  inverter_0 ../inverter
timestamp 1661503936
transform 1 0 144 0 1 2516
box -13 -65 104 246
use inverter  inverter_1
timestamp 1661503936
transform 1 0 261 0 1 2516
box -13 -65 104 246
<< labels >>
rlabel metal1 -61 2587 -61 2601 7 clk
port 1 w
rlabel locali 1039 2438 1039 2465 7 nclk
port 10 w
<< end >>
