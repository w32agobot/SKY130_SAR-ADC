magic
tech sky130A
magscale 1 2
timestamp 1661174129
<< error_s >>
rect 94 677 152 683
rect 286 677 344 683
rect 478 677 536 683
rect 670 677 728 683
rect 94 643 106 677
rect 286 643 298 677
rect 478 643 490 677
rect 670 643 682 677
rect 94 637 152 643
rect 286 637 344 643
rect 478 637 536 643
rect 670 637 728 643
rect 0 455 812 474
rect -2 434 812 455
rect -2 409 716 434
rect 0 396 716 409
<< nwell >>
rect 238 -316 560 220
<< nmos >>
rect 48 -910 78 -510
rect 144 -910 174 -510
rect 240 -910 270 -510
rect 336 -910 366 -510
rect 432 -910 462 -510
rect 528 -910 558 -510
rect 624 -910 654 -510
rect 720 -910 750 -510
rect 330 -1516 360 -1116
rect 426 -1516 456 -1116
<< pmos >>
rect 336 -280 366 120
rect 432 -280 462 120
<< ndiff >>
rect -14 -522 48 -510
rect -14 -898 -2 -522
rect 32 -898 48 -522
rect -14 -910 48 -898
rect 78 -522 144 -510
rect 78 -898 94 -522
rect 128 -898 144 -522
rect 78 -910 144 -898
rect 174 -522 240 -510
rect 174 -898 190 -522
rect 224 -898 240 -522
rect 174 -910 240 -898
rect 270 -522 336 -510
rect 270 -898 286 -522
rect 320 -898 336 -522
rect 270 -910 336 -898
rect 366 -522 432 -510
rect 366 -898 382 -522
rect 416 -898 432 -522
rect 366 -910 432 -898
rect 462 -522 528 -510
rect 462 -898 478 -522
rect 512 -898 528 -522
rect 462 -910 528 -898
rect 558 -522 624 -510
rect 558 -898 574 -522
rect 608 -898 624 -522
rect 558 -910 624 -898
rect 654 -522 720 -510
rect 654 -898 670 -522
rect 704 -898 720 -522
rect 654 -910 720 -898
rect 750 -522 812 -510
rect 750 -898 766 -522
rect 800 -898 812 -522
rect 750 -910 812 -898
rect 268 -1128 330 -1116
rect 268 -1504 280 -1128
rect 314 -1504 330 -1128
rect 268 -1516 330 -1504
rect 360 -1128 426 -1116
rect 360 -1504 376 -1128
rect 410 -1504 426 -1128
rect 360 -1516 426 -1504
rect 456 -1128 518 -1116
rect 456 -1504 472 -1128
rect 506 -1504 518 -1128
rect 456 -1516 518 -1504
<< pdiff >>
rect 274 108 336 120
rect 274 -268 286 108
rect 320 -268 336 108
rect 274 -280 336 -268
rect 366 108 432 120
rect 366 -268 382 108
rect 416 -268 432 108
rect 366 -280 432 -268
rect 462 108 524 120
rect 462 -268 478 108
rect 512 -268 524 108
rect 462 -280 524 -268
<< ndiffc >>
rect -2 -898 32 -522
rect 94 -898 128 -522
rect 190 -898 224 -522
rect 286 -898 320 -522
rect 382 -898 416 -522
rect 478 -898 512 -522
rect 574 -898 608 -522
rect 670 -898 704 -522
rect 766 -898 800 -522
rect 280 -1504 314 -1128
rect 376 -1504 410 -1128
rect 472 -1504 506 -1128
<< pdiffc >>
rect 286 -268 320 108
rect 382 -268 416 108
rect 478 -268 512 108
<< poly >>
rect 336 120 366 146
rect 432 120 462 146
rect 336 -316 366 -280
rect 432 -316 462 -280
rect 336 -346 462 -316
rect 48 -510 78 -484
rect 144 -510 174 -484
rect 240 -510 270 -484
rect 336 -510 366 -484
rect 432 -510 462 -484
rect 528 -510 558 -484
rect 624 -510 654 -484
rect 720 -510 750 -484
rect 48 -938 78 -910
rect 144 -938 174 -910
rect 240 -938 270 -910
rect 336 -938 366 -910
rect 48 -968 366 -938
rect 432 -938 462 -910
rect 528 -938 558 -910
rect 624 -938 654 -910
rect 720 -938 750 -910
rect 432 -968 750 -938
rect 330 -1116 360 -1090
rect 426 -1116 456 -1090
rect 330 -1542 360 -1516
rect 426 -1542 456 -1516
<< locali >>
rect 286 108 320 124
rect 286 -438 320 -268
rect 382 108 416 206
rect 382 -284 416 -268
rect 478 108 512 124
rect 94 -472 320 -438
rect -2 -522 32 -506
rect -2 -972 32 -898
rect 94 -522 128 -472
rect 94 -938 128 -898
rect 190 -522 224 -506
rect 190 -972 224 -898
rect 286 -522 320 -472
rect 478 -438 512 -268
rect 478 -472 704 -438
rect 286 -938 320 -898
rect 382 -522 416 -506
rect 382 -972 416 -898
rect 478 -522 512 -472
rect 478 -938 512 -898
rect 574 -522 608 -506
rect 574 -972 608 -898
rect 670 -522 704 -472
rect 670 -938 704 -898
rect 766 -522 800 -506
rect 766 -972 800 -898
rect -2 -1006 800 -972
rect 280 -1128 314 -1112
rect 280 -1520 314 -1504
rect 376 -1128 410 -1112
rect 376 -1520 410 -1504
rect 472 -1128 506 -1112
rect 472 -1520 506 -1504
<< viali >>
rect 286 -268 320 108
rect 382 -268 416 108
rect 478 -268 512 108
rect -2 -898 32 -522
rect 94 -898 128 -522
rect 190 -898 224 -522
rect 286 -898 320 -522
rect 382 -898 416 -522
rect 478 -898 512 -522
rect 574 -898 608 -522
rect 670 -898 704 -522
rect 766 -898 800 -522
rect 280 -1504 314 -1128
rect 376 -1504 410 -1128
rect 472 -1504 506 -1128
<< metal1 >>
rect 280 108 326 120
rect 280 -268 286 108
rect 320 -268 326 108
rect 280 -280 326 -268
rect 376 108 422 120
rect 376 -268 382 108
rect 416 -268 422 108
rect 376 -280 422 -268
rect 472 108 518 120
rect 472 -268 478 108
rect 512 -268 518 108
rect 472 -280 518 -268
rect -8 -522 38 -510
rect -8 -898 -2 -522
rect 32 -898 38 -522
rect -8 -910 38 -898
rect 88 -522 134 -510
rect 88 -898 94 -522
rect 128 -898 134 -522
rect 88 -910 134 -898
rect 184 -522 230 -510
rect 184 -898 190 -522
rect 224 -898 230 -522
rect 184 -910 230 -898
rect 280 -522 326 -510
rect 280 -898 286 -522
rect 320 -898 326 -522
rect 280 -910 326 -898
rect 376 -522 422 -510
rect 376 -898 382 -522
rect 416 -898 422 -522
rect 376 -910 422 -898
rect 472 -522 518 -510
rect 472 -898 478 -522
rect 512 -898 518 -522
rect 472 -910 518 -898
rect 568 -522 614 -510
rect 568 -898 574 -522
rect 608 -898 614 -522
rect 568 -910 614 -898
rect 664 -522 710 -510
rect 664 -898 670 -522
rect 704 -898 710 -522
rect 664 -910 710 -898
rect 760 -522 806 -510
rect 760 -898 766 -522
rect 800 -898 806 -522
rect 760 -910 806 -898
rect 274 -1128 320 -1116
rect 274 -1504 280 -1128
rect 314 -1504 320 -1128
rect 274 -1516 320 -1504
rect 370 -1128 416 -1116
rect 370 -1504 376 -1128
rect 410 -1504 416 -1128
rect 370 -1516 416 -1504
rect 466 -1128 512 -1116
rect 466 -1504 472 -1128
rect 506 -1504 512 -1128
rect 466 -1516 512 -1504
use sky130_fd_pr__pfet_01v8_52F6HE  sky130_fd_pr__pfet_01v8_52F6HE_0
timestamp 1661174129
transform 1 0 363 0 1 546
box -449 -150 449 150
<< end >>
