magic
tech sky130A
magscale 1 2
timestamp 1673705348
<< nwell >>
rect -10 48 408 452
<< nmos >>
rect 88 -216 118 -116
rect 184 -216 214 -116
rect 280 -216 310 -116
<< pmos >>
rect 88 110 118 310
rect 184 110 214 310
rect 280 110 310 310
<< ndiff >>
rect 26 -134 88 -116
rect 26 -204 38 -134
rect 72 -204 88 -134
rect 26 -216 88 -204
rect 118 -128 184 -116
rect 118 -204 134 -128
rect 168 -204 184 -128
rect 118 -216 184 -204
rect 214 -128 280 -116
rect 214 -204 230 -128
rect 264 -204 280 -128
rect 214 -216 280 -204
rect 310 -128 372 -116
rect 310 -204 326 -128
rect 360 -204 372 -128
rect 310 -216 372 -204
<< pdiff >>
rect 26 298 88 310
rect 26 122 38 298
rect 72 122 88 298
rect 26 110 88 122
rect 118 298 184 310
rect 118 122 134 298
rect 168 122 184 298
rect 118 110 184 122
rect 214 298 280 310
rect 214 122 230 298
rect 264 122 280 298
rect 214 110 280 122
rect 310 298 372 310
rect 310 122 326 298
rect 360 122 372 298
rect 310 110 372 122
<< ndiffc >>
rect 38 -204 72 -134
rect 134 -204 168 -128
rect 230 -204 264 -128
rect 326 -204 360 -128
<< pdiffc >>
rect 38 122 72 298
rect 134 122 168 298
rect 230 122 264 298
rect 326 122 360 298
<< psubdiff >>
rect -42 -304 -16 -270
rect 18 -304 52 -270
rect 86 -304 120 -270
rect 154 -304 188 -270
rect 222 -304 256 -270
rect 290 -304 324 -270
rect 358 -304 382 -270
rect -42 -306 382 -304
<< nsubdiff >>
rect 26 378 50 416
rect 88 378 126 416
rect 164 378 202 416
rect 240 378 278 416
rect 316 378 372 416
<< psubdiffcont >>
rect -16 -304 18 -270
rect 52 -304 86 -270
rect 120 -304 154 -270
rect 188 -304 222 -270
rect 256 -304 290 -270
rect 324 -304 358 -270
<< nsubdiffcont >>
rect 50 378 88 416
rect 126 378 164 416
rect 202 378 240 416
rect 278 378 316 416
<< poly >>
rect 88 310 118 336
rect 184 310 214 336
rect 280 310 310 336
rect 88 28 118 110
rect 184 84 214 110
rect 280 84 310 110
rect 184 48 310 84
rect 68 11 128 28
rect 68 -23 78 11
rect 112 -23 128 11
rect 68 -40 128 -23
rect 216 11 274 48
rect 216 -23 226 11
rect 260 -23 274 11
rect 88 -116 118 -40
rect 216 -70 274 -23
rect 184 -100 310 -70
rect 184 -116 214 -100
rect 280 -116 310 -100
rect 88 -242 118 -216
rect 184 -242 214 -216
rect 280 -242 310 -216
<< polycont >>
rect 78 -23 112 11
rect 226 -23 260 11
<< locali >>
rect -42 378 50 416
rect 88 378 126 416
rect 164 378 202 416
rect 240 378 278 416
rect 316 378 408 416
rect 38 298 72 314
rect 38 106 72 122
rect 134 298 168 378
rect 134 106 168 122
rect 230 298 264 314
rect 230 106 264 122
rect 326 298 360 378
rect 326 106 360 122
rect 68 12 128 28
rect 68 -24 78 12
rect 112 -24 128 12
rect 68 -40 128 -24
rect 216 12 262 28
rect 216 -24 226 12
rect 260 -24 262 12
rect 216 -40 262 -24
rect 38 -134 72 -112
rect 38 -220 72 -204
rect 134 -128 168 -112
rect 134 -270 168 -204
rect 230 -128 264 -112
rect 230 -220 264 -204
rect 326 -128 360 -112
rect 326 -270 360 -204
rect -42 -304 -16 -270
rect 18 -304 52 -270
rect 86 -304 120 -270
rect 154 -304 188 -270
rect 222 -304 256 -270
rect 290 -304 324 -270
rect 358 -304 382 -270
rect -42 -306 382 -304
<< viali >>
rect 38 122 72 186
rect 230 160 264 198
rect 78 11 112 12
rect 78 -23 112 11
rect 78 -24 112 -23
rect 226 11 260 12
rect 226 -23 260 11
rect 226 -24 260 -23
rect 38 -186 72 -134
rect 230 -188 264 -148
<< metal1 >>
rect 224 198 360 218
rect 32 186 78 198
rect 32 122 38 186
rect 72 122 78 186
rect 224 160 230 198
rect 264 160 360 198
rect 224 142 360 160
rect 32 116 78 122
rect 38 84 72 116
rect 38 56 272 84
rect 68 12 128 28
rect 68 8 78 12
rect -16 -20 78 8
rect 68 -24 78 -20
rect 112 -24 128 12
rect 68 -40 128 -24
rect 214 12 272 56
rect 214 -24 226 12
rect 260 -24 272 12
rect 214 -68 272 -24
rect 38 -96 272 -68
rect 326 8 360 142
rect 326 -20 408 8
rect 38 -124 72 -96
rect 32 -134 78 -124
rect 326 -128 360 -20
rect 32 -186 38 -134
rect 72 -186 78 -134
rect 32 -198 78 -186
rect 224 -148 360 -128
rect 224 -188 230 -148
rect 264 -188 360 -148
rect 224 -204 360 -188
<< labels >>
flabel metal1 356 -20 408 8 0 FreeSans 160 0 0 0 out
port 8 nsew
flabel metal1 -16 -20 34 8 0 FreeSans 160 0 0 0 in
port 12 nsew
flabel locali -42 -306 382 -270 0 FreeSans 160 0 0 0 VSS
port 13 nsew
flabel locali -42 378 408 416 0 FreeSans 160 0 0 0 VDD
port 14 nsew
<< end >>
