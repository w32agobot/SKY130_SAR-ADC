* SPICE3 file created from adc_array_wafflecap_8(4)x557aF_25um2.ext - technology: sky130A

.subckt adc_array_wafflecap_8(4)x557aF_25um2 cbot ctop
C0 ctop cbot 2.25fF
C1 nc cbot 2.16fF
C2 cbot VSUBS 2.01fF
.ends
