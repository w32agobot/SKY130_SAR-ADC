* SPICE3 file created from adc_array_fingercap_8(1)x360aF_topB_22um2.ext - technology: sky130A

C0 VSS floatingmetal 0.79fF
C1 cbot floatingmetal 2.36fF
C2 cbot VSS 3.09fF
C3 floatingmetal ctop 0.30fF
C4 VSS ctop 0.25fF
C5 cbot ctop 0.39fF
C6 floatingmetal VSUBS 0.71fF
C7 ctop VSUBS 0.25fF
C8 cbot VSUBS 0.43fF
C9 VSS VSUBS 1.80fF
