magic
tech sky130A
magscale 1 2
timestamp 1665667482
<< nwell >>
rect 0 873 141 880
rect 151 873 705 886
rect 859 873 1004 880
rect 0 506 1004 873
rect 141 499 859 506
<< locali >>
rect 34 924 148 1004
rect 34 888 46 924
rect 136 888 148 924
rect 34 706 148 888
rect 34 670 46 706
rect 136 670 148 706
rect 34 610 148 670
rect 34 574 46 610
rect 136 574 148 610
rect 34 266 148 574
rect 34 232 114 266
rect 34 102 148 232
rect 34 66 46 102
rect 136 66 148 102
rect 34 0 148 66
rect 854 924 970 1004
rect 854 888 866 924
rect 958 888 970 924
rect 854 706 970 888
rect 854 670 866 706
rect 958 670 970 706
rect 854 610 970 670
rect 854 574 866 610
rect 958 574 970 610
rect 854 340 970 574
rect 854 282 866 340
rect 958 282 970 340
rect 854 102 970 282
rect 854 66 866 102
rect 958 66 970 102
rect 854 0 970 66
<< viali >>
rect 46 888 136 924
rect 46 670 136 706
rect 46 574 136 610
rect 114 232 148 266
rect 46 66 136 102
rect 866 888 958 924
rect 866 670 958 706
rect 866 574 958 610
rect 866 282 958 340
rect 866 66 958 102
<< metal1 >>
rect 34 924 148 1004
rect 34 888 46 924
rect 136 888 148 924
rect 34 882 148 888
rect 854 924 970 1004
rect 854 888 866 924
rect 958 888 970 924
rect 854 882 970 888
rect 0 798 1004 854
rect 0 740 1004 770
rect 34 706 148 712
rect 34 670 46 706
rect 136 670 148 706
rect 34 610 148 670
rect 34 574 46 610
rect 136 574 148 610
rect 34 568 148 574
rect 854 706 970 712
rect 854 670 866 706
rect 958 670 970 706
rect 854 610 970 670
rect 854 574 866 610
rect 958 574 970 610
rect 854 568 970 574
rect 0 512 1004 540
rect 0 430 1004 458
rect 0 374 1004 402
rect 854 340 970 346
rect 854 282 866 340
rect 958 282 970 340
rect 108 266 154 278
rect 854 276 970 282
rect 108 248 114 266
rect 0 232 114 248
rect 148 248 154 266
rect 148 232 1004 248
rect 0 220 1004 232
rect 0 136 1004 192
rect 34 102 148 108
rect 34 66 46 102
rect 136 66 148 102
rect 34 0 148 66
rect 854 102 970 108
rect 854 66 866 102
rect 958 66 970 102
rect 854 0 970 66
<< metal2 >>
rect 32 962 972 972
rect 32 906 42 962
rect 98 906 138 962
rect 194 906 234 962
rect 290 906 330 962
rect 386 906 426 962
rect 482 906 522 962
rect 578 906 618 962
rect 674 906 714 962
rect 770 906 810 962
rect 866 906 906 962
rect 962 906 972 962
rect 32 866 972 906
rect 32 810 42 866
rect 98 810 330 866
rect 386 810 618 866
rect 674 810 906 866
rect 962 810 972 866
rect 32 776 972 810
rect 32 770 396 776
rect 32 714 42 770
rect 98 714 330 770
rect 386 714 396 770
rect 32 674 396 714
rect 608 770 972 776
rect 608 714 618 770
rect 674 714 906 770
rect 962 714 972 770
rect 32 618 42 674
rect 98 618 138 674
rect 194 618 234 674
rect 290 618 330 674
rect 386 618 396 674
rect 32 578 396 618
rect 474 691 530 700
rect 474 610 530 627
rect 608 674 972 714
rect 608 618 618 674
rect 674 618 714 674
rect 770 618 810 674
rect 866 618 906 674
rect 962 618 972 674
rect 32 522 42 578
rect 98 522 396 578
rect 32 512 396 522
rect 608 578 972 618
rect 608 522 906 578
rect 962 522 972 578
rect 608 512 972 522
rect 32 482 972 512
rect 32 426 42 482
rect 98 426 906 482
rect 962 426 972 482
rect 32 386 972 426
rect 32 330 42 386
rect 98 330 138 386
rect 194 330 234 386
rect 290 330 714 386
rect 770 330 810 386
rect 866 330 906 386
rect 962 330 972 386
rect 32 290 972 330
rect 32 234 42 290
rect 98 234 906 290
rect 962 234 972 290
rect 32 194 972 234
rect 32 138 42 194
rect 98 138 906 194
rect 962 138 972 194
rect 32 98 972 138
rect 32 42 42 98
rect 98 42 138 98
rect 194 42 234 98
rect 290 49 714 98
rect 290 42 330 49
rect 32 32 330 42
rect 650 42 714 49
rect 770 42 810 98
rect 866 42 906 98
rect 962 42 972 98
rect 650 32 972 42
<< via2 >>
rect 42 906 98 962
rect 138 906 194 962
rect 234 906 290 962
rect 330 906 386 962
rect 426 906 482 962
rect 522 906 578 962
rect 618 906 674 962
rect 714 906 770 962
rect 810 906 866 962
rect 906 906 962 962
rect 42 810 98 866
rect 330 810 386 866
rect 618 810 674 866
rect 906 810 962 866
rect 42 714 98 770
rect 330 714 386 770
rect 618 714 674 770
rect 906 714 962 770
rect 42 618 98 674
rect 138 618 194 674
rect 234 618 290 674
rect 330 618 386 674
rect 474 627 530 691
rect 618 618 674 674
rect 714 618 770 674
rect 810 618 866 674
rect 906 618 962 674
rect 42 522 98 578
rect 906 522 962 578
rect 42 426 98 482
rect 906 426 962 482
rect 42 330 98 386
rect 138 330 194 386
rect 234 330 290 386
rect 714 330 770 386
rect 810 330 866 386
rect 906 330 962 386
rect 42 234 98 290
rect 906 234 962 290
rect 42 138 98 194
rect 906 138 962 194
rect 42 42 98 98
rect 138 42 194 98
rect 234 42 290 98
rect 714 42 770 98
rect 810 42 866 98
rect 906 42 962 98
<< metal3 >>
rect 36 962 968 968
rect 36 906 42 962
rect 98 906 138 962
rect 194 906 234 962
rect 290 906 330 962
rect 386 906 426 962
rect 482 906 522 962
rect 578 906 618 962
rect 674 906 714 962
rect 770 906 810 962
rect 866 906 906 962
rect 962 906 968 962
rect 36 900 968 906
rect 36 866 104 900
rect 36 810 42 866
rect 98 810 104 866
rect 324 866 392 900
rect 36 770 104 810
rect 36 714 42 770
rect 98 714 104 770
rect 164 824 264 840
rect 164 756 180 824
rect 248 756 264 824
rect 164 740 264 756
rect 324 810 330 866
rect 386 810 392 866
rect 324 770 392 810
rect 36 680 104 714
rect 324 714 330 770
rect 386 714 392 770
rect 612 866 680 900
rect 612 810 618 866
rect 674 810 680 866
rect 900 866 968 900
rect 612 770 680 810
rect 324 680 392 714
rect 36 674 392 680
rect 36 618 42 674
rect 98 618 138 674
rect 194 618 234 674
rect 290 618 330 674
rect 386 618 392 674
rect 36 612 392 618
rect 468 691 536 732
rect 468 627 470 691
rect 534 627 536 691
rect 36 578 104 612
rect 468 582 536 627
rect 612 714 618 770
rect 674 714 680 770
rect 740 824 840 840
rect 740 756 756 824
rect 824 756 840 824
rect 740 740 840 756
rect 900 810 906 866
rect 962 810 968 866
rect 900 770 968 810
rect 612 680 680 714
rect 900 714 906 770
rect 962 714 968 770
rect 900 680 968 714
rect 612 674 968 680
rect 612 618 618 674
rect 674 618 714 674
rect 770 618 810 674
rect 866 618 906 674
rect 962 618 968 674
rect 612 612 968 618
rect 36 522 42 578
rect 98 522 104 578
rect 900 578 968 612
rect 36 482 104 522
rect 36 426 42 482
rect 98 426 104 482
rect 164 536 264 552
rect 164 468 180 536
rect 248 468 264 536
rect 164 452 264 468
rect 740 536 840 552
rect 740 468 756 536
rect 824 468 840 536
rect 740 452 840 468
rect 900 522 906 578
rect 962 522 968 578
rect 900 482 968 522
rect 36 392 104 426
rect 900 426 906 482
rect 962 426 968 482
rect 900 392 968 426
rect 36 386 324 392
rect 36 330 42 386
rect 98 330 138 386
rect 194 330 234 386
rect 290 330 324 386
rect 36 324 324 330
rect 692 386 968 392
rect 692 330 714 386
rect 770 330 810 386
rect 866 330 906 386
rect 962 330 968 386
rect 692 324 968 330
rect 36 290 104 324
rect 36 234 42 290
rect 98 234 104 290
rect 900 290 968 324
rect 36 194 104 234
rect 36 138 42 194
rect 98 138 104 194
rect 164 248 264 264
rect 164 180 180 248
rect 248 180 264 248
rect 164 164 264 180
rect 740 248 840 264
rect 740 180 756 248
rect 824 180 840 248
rect 740 164 840 180
rect 900 234 906 290
rect 962 234 968 290
rect 900 194 968 234
rect 36 104 104 138
rect 900 138 906 194
rect 962 138 968 194
rect 900 104 968 138
rect 36 98 324 104
rect 36 42 42 98
rect 98 42 138 98
rect 194 42 234 98
rect 290 42 324 98
rect 36 36 324 42
rect 692 98 968 104
rect 692 42 714 98
rect 770 42 810 98
rect 866 42 906 98
rect 962 42 968 98
rect 692 36 968 42
<< via3 >>
rect 180 756 248 824
rect 470 627 474 691
rect 474 627 530 691
rect 530 627 534 691
rect 756 756 824 824
rect 180 468 248 536
rect 756 468 824 536
rect 180 180 248 248
rect 756 180 824 248
<< metal4 >>
rect 184 840 244 934
rect 164 824 264 840
rect 164 820 180 824
rect 70 760 180 820
rect 164 756 180 760
rect 248 820 264 824
rect 248 760 360 820
rect 248 756 264 760
rect 164 740 264 756
rect 184 552 244 740
rect 472 732 532 934
rect 760 840 820 934
rect 740 824 840 840
rect 740 820 756 824
rect 646 760 756 820
rect 740 756 756 760
rect 824 820 840 824
rect 824 760 934 820
rect 824 756 840 760
rect 740 740 840 756
rect 470 698 534 732
rect 468 691 536 698
rect 468 627 470 691
rect 534 627 536 691
rect 468 612 536 627
rect 470 582 534 612
rect 164 536 264 552
rect 164 532 180 536
rect 70 472 180 532
rect 164 468 180 472
rect 248 468 264 536
rect 164 452 264 468
rect 184 264 244 452
rect 164 248 264 264
rect 164 244 180 248
rect 70 184 180 244
rect 164 180 180 184
rect 248 180 264 248
rect 164 164 264 180
rect 184 70 244 164
rect 472 49 532 582
rect 760 552 820 740
rect 740 536 840 552
rect 740 468 756 536
rect 824 532 840 536
rect 824 472 934 532
rect 824 468 840 472
rect 740 452 840 468
rect 760 264 820 452
rect 740 248 840 264
rect 740 180 756 248
rect 824 244 840 248
rect 824 184 934 244
rect 824 180 840 184
rect 740 164 840 180
rect 760 70 820 164
<< comment >>
rect 0 972 32 1004
rect 972 972 1004 1004
rect 0 0 32 32
rect 972 0 1004 32
use sky130_fd_pr__nfet_01v8_AVE2UL  sky130_fd_pr__nfet_01v8_AVE2UL_0
timestamp 1665667482
transform 1 0 504 0 1 231
box -323 -226 323 226
use sky130_fd_pr__pfet_01v8_KZGJBR  sky130_fd_pr__pfet_01v8_KZGJBR_0
timestamp 1665667482
transform 1 0 500 0 1 768
box -360 -238 359 237
<< labels >>
rlabel metal1 0 740 0 770 7 sample_n
port 2 w
rlabel metal1 0 512 0 540 7 colon_n
port 3 w
rlabel metal1 0 430 0 458 7 col_n
port 4 w
rlabel metal1 0 374 0 402 7 sample
port 5 w
rlabel metal1 0 220 0 248 7 vcom
port 6 w
rlabel metal1 0 136 0 192 7 VSS
port 7 w
rlabel locali 854 0 970 0 5 row_n
port 8 s
rlabel metal1 0 798 0 854 7 VDD
port 13 w
<< end >>
