magic
tech sky130A
magscale 1 2
timestamp 1673698727
<< nwell >>
rect -8 69 506 390
<< nmos >>
rect 186 -126 216 -42
rect 282 -126 312 -42
<< pmos >>
rect 90 106 120 266
rect 186 106 216 266
rect 282 106 312 266
rect 378 106 408 266
<< ndiff >>
rect 124 -54 186 -42
rect 124 -114 136 -54
rect 170 -114 186 -54
rect 124 -126 186 -114
rect 216 -54 282 -42
rect 216 -114 232 -54
rect 266 -114 282 -54
rect 216 -126 282 -114
rect 312 -54 374 -42
rect 312 -114 328 -54
rect 362 -114 374 -54
rect 312 -126 374 -114
<< pdiff >>
rect 28 254 90 266
rect 28 118 40 254
rect 74 118 90 254
rect 28 106 90 118
rect 120 254 186 266
rect 120 118 136 254
rect 170 118 186 254
rect 120 106 186 118
rect 216 254 282 266
rect 216 118 232 254
rect 266 118 282 254
rect 216 106 282 118
rect 312 254 378 266
rect 312 118 328 254
rect 362 118 378 254
rect 312 106 378 118
rect 408 254 470 266
rect 408 118 424 254
rect 458 118 470 254
rect 408 106 470 118
<< ndiffc >>
rect 136 -114 170 -54
rect 232 -114 266 -54
rect 328 -114 362 -54
<< pdiffc >>
rect 40 118 74 254
rect 136 118 170 254
rect 232 118 266 254
rect 328 118 362 254
rect 424 118 458 254
<< psubdiff >>
rect 62 -214 96 -180
rect 130 -214 164 -180
rect 198 -214 232 -180
rect 266 -214 300 -180
rect 334 -214 368 -180
rect 402 -214 436 -180
<< nsubdiff >>
rect 40 320 96 354
rect 130 320 164 354
rect 198 320 232 354
rect 266 320 300 354
rect 334 320 368 354
rect 402 320 458 354
<< psubdiffcont >>
rect 96 -214 130 -180
rect 164 -214 198 -180
rect 232 -214 266 -180
rect 300 -214 334 -180
rect 368 -214 402 -180
<< nsubdiffcont >>
rect 96 320 130 354
rect 164 320 198 354
rect 232 320 266 354
rect 300 320 334 354
rect 368 320 402 354
<< poly >>
rect 90 266 120 293
rect 186 266 216 292
rect 282 266 312 293
rect 378 266 408 292
rect 90 60 120 106
rect 186 66 216 106
rect 52 44 120 60
rect 52 10 70 44
rect 104 10 120 44
rect 52 0 120 10
rect 162 56 222 66
rect 282 60 312 106
rect 378 66 408 106
rect 162 22 178 56
rect 212 22 222 56
rect 162 6 222 22
rect 276 45 336 60
rect 276 11 286 45
rect 320 11 336 45
rect 186 -42 216 6
rect 276 1 336 11
rect 378 56 446 66
rect 378 22 396 56
rect 430 22 446 56
rect 378 6 446 22
rect 282 -42 312 1
rect 186 -152 216 -126
rect 282 -152 312 -126
<< polycont >>
rect 70 10 104 44
rect 178 22 212 56
rect 286 11 320 45
rect 396 22 430 56
<< locali >>
rect 40 320 96 354
rect 130 320 164 354
rect 198 320 232 354
rect 266 320 300 354
rect 334 320 368 354
rect 402 320 458 354
rect 40 254 74 320
rect 40 102 74 118
rect 136 254 170 270
rect 136 102 170 118
rect 232 254 266 270
rect 232 102 266 118
rect 328 254 362 270
rect 328 102 362 118
rect 424 254 458 320
rect 424 102 458 118
rect 52 44 120 60
rect 52 10 70 44
rect 104 10 120 44
rect 52 0 120 10
rect 162 56 230 66
rect 162 22 178 56
rect 212 22 230 56
rect 162 6 230 22
rect 268 45 336 60
rect 268 10 286 45
rect 320 10 336 45
rect 268 1 336 10
rect 378 56 446 66
rect 378 22 396 56
rect 430 22 446 56
rect 378 6 446 22
rect 136 -54 170 -38
rect 136 -180 170 -114
rect 232 -54 266 -38
rect 232 -130 266 -122
rect 328 -54 362 -38
rect 328 -180 362 -114
rect 62 -214 96 -180
rect 130 -214 164 -180
rect 198 -214 232 -180
rect 266 -214 300 -180
rect 334 -214 368 -180
rect 402 -214 436 -180
<< viali >>
rect 232 155 266 189
rect 70 10 104 44
rect 178 22 212 56
rect 286 11 320 44
rect 286 10 320 11
rect 396 22 430 56
rect 232 -114 266 -88
rect 232 -122 266 -114
<< metal1 >>
rect 223 198 275 204
rect 223 140 275 146
rect 22 84 476 112
rect 168 56 220 84
rect 386 56 438 84
rect 61 44 113 56
rect 61 10 70 44
rect 104 10 113 44
rect 168 22 178 56
rect 212 22 220 56
rect 168 10 220 22
rect 276 44 336 56
rect 276 10 286 44
rect 320 10 336 44
rect 386 22 396 56
rect 430 22 438 56
rect 386 10 438 22
rect 61 -19 113 10
rect 276 -19 336 10
rect 22 -47 476 -19
rect 223 -84 275 -76
rect 223 -147 275 -140
<< via1 >>
rect 223 189 275 198
rect 223 155 232 189
rect 232 155 266 189
rect 266 155 275 189
rect 223 146 275 155
rect 223 -88 275 -84
rect 223 -122 232 -88
rect 232 -122 266 -88
rect 266 -122 275 -88
rect 223 -140 275 -122
<< metal2 >>
rect 221 198 277 209
rect 221 146 223 198
rect 275 146 277 198
rect 221 135 277 146
rect 223 -84 275 135
rect 22 -140 223 -119
rect 275 -140 476 -119
rect 22 -147 476 -140
<< labels >>
flabel metal2 22 -147 476 -119 0 FreeSans 160 0 0 0 q
port 5 nsew
flabel metal1 22 84 476 112 0 FreeSans 160 0 0 0 a
port 6 nsew
flabel metal1 22 -47 476 -19 0 FreeSans 160 0 0 0 b
port 7 nsew
flabel locali 62 -214 436 -180 0 FreeSans 160 0 0 0 VSS
port 8 nsew
flabel locali 40 320 458 354 0 FreeSans 160 0 0 0 VDD
port 10 nsew
<< end >>
