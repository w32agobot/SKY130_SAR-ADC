magic
tech sky130A
magscale 1 2
timestamp 1661427359
<< nwell >>
rect -52 -178 2590 226
rect -52 -196 2336 -178
rect 474 -198 716 -196
rect 1178 -546 2336 -196
<< nmos >>
rect 48 -910 78 -510
rect 144 -910 174 -510
rect 240 -910 270 -510
rect 336 -910 366 -510
rect 432 -910 462 -510
rect 528 -910 558 -510
rect 624 -910 654 -510
rect 720 -910 750 -510
rect 48 -1170 78 -1070
rect 144 -1170 174 -1070
rect 240 -1170 270 -1070
rect 336 -1170 366 -1070
rect 432 -1170 462 -1070
rect 528 -1170 558 -1070
rect 624 -1170 654 -1070
rect 720 -1170 750 -1070
rect 1598 -1176 1628 -776
rect 1694 -1176 1724 -776
rect 1790 -1176 1820 -776
rect 1886 -1176 1916 -776
<< pmos >>
rect 48 -96 78 4
rect 144 -96 174 4
rect 240 -96 270 4
rect 336 -96 366 4
rect 432 -96 462 4
rect 528 -96 558 4
rect 624 -96 654 4
rect 720 -96 750 4
rect 1276 -446 1306 -46
rect 1372 -446 1402 -46
rect 1598 -446 1628 -46
rect 1694 -446 1724 -46
rect 1790 -446 1820 -46
rect 1886 -446 1916 -46
rect 2112 -446 2142 -46
rect 2208 -446 2238 -46
<< ndiff >>
rect -14 -522 48 -510
rect -14 -898 -2 -522
rect 32 -898 48 -522
rect -14 -910 48 -898
rect 78 -522 144 -510
rect 78 -898 94 -522
rect 128 -898 144 -522
rect 78 -910 144 -898
rect 174 -522 240 -510
rect 174 -898 190 -522
rect 224 -898 240 -522
rect 174 -910 240 -898
rect 270 -522 336 -510
rect 270 -898 286 -522
rect 320 -898 336 -522
rect 270 -910 336 -898
rect 366 -522 432 -510
rect 366 -898 382 -522
rect 416 -898 432 -522
rect 366 -910 432 -898
rect 462 -522 528 -510
rect 462 -898 478 -522
rect 512 -898 528 -522
rect 462 -910 528 -898
rect 558 -522 624 -510
rect 558 -898 574 -522
rect 608 -898 624 -522
rect 558 -910 624 -898
rect 654 -522 720 -510
rect 654 -898 670 -522
rect 704 -898 720 -522
rect 654 -910 720 -898
rect 750 -522 812 -510
rect 750 -898 766 -522
rect 800 -898 812 -522
rect 750 -910 812 -898
rect 1536 -788 1598 -776
rect -14 -1082 48 -1070
rect -14 -1158 -2 -1082
rect 32 -1158 48 -1082
rect -14 -1170 48 -1158
rect 78 -1082 144 -1070
rect 78 -1158 94 -1082
rect 128 -1158 144 -1082
rect 78 -1170 144 -1158
rect 174 -1082 240 -1070
rect 174 -1158 190 -1082
rect 224 -1158 240 -1082
rect 174 -1170 240 -1158
rect 270 -1082 336 -1070
rect 270 -1158 286 -1082
rect 320 -1158 336 -1082
rect 270 -1170 336 -1158
rect 366 -1082 432 -1070
rect 366 -1158 382 -1082
rect 416 -1158 432 -1082
rect 366 -1170 432 -1158
rect 462 -1082 528 -1070
rect 462 -1158 478 -1082
rect 512 -1158 528 -1082
rect 462 -1170 528 -1158
rect 558 -1082 624 -1070
rect 558 -1158 574 -1082
rect 608 -1158 624 -1082
rect 558 -1170 624 -1158
rect 654 -1082 720 -1070
rect 654 -1158 670 -1082
rect 704 -1158 720 -1082
rect 654 -1170 720 -1158
rect 750 -1082 812 -1070
rect 750 -1158 766 -1082
rect 800 -1158 812 -1082
rect 750 -1170 812 -1158
rect 1536 -1164 1548 -788
rect 1582 -1164 1598 -788
rect 1536 -1176 1598 -1164
rect 1628 -788 1694 -776
rect 1628 -1164 1644 -788
rect 1678 -1164 1694 -788
rect 1628 -1176 1694 -1164
rect 1724 -788 1790 -776
rect 1724 -1164 1740 -788
rect 1774 -1164 1790 -788
rect 1724 -1176 1790 -1164
rect 1820 -788 1886 -776
rect 1820 -1164 1836 -788
rect 1870 -1164 1886 -788
rect 1820 -1176 1886 -1164
rect 1916 -788 1978 -776
rect 1916 -1164 1932 -788
rect 1966 -1164 1978 -788
rect 1916 -1176 1978 -1164
<< pdiff >>
rect -14 -8 48 4
rect -14 -84 -2 -8
rect 32 -84 48 -8
rect -14 -96 48 -84
rect 78 -8 144 4
rect 78 -84 94 -8
rect 128 -84 144 -8
rect 78 -96 144 -84
rect 174 -8 240 4
rect 174 -84 190 -8
rect 224 -84 240 -8
rect 174 -96 240 -84
rect 270 -8 336 4
rect 270 -84 286 -8
rect 320 -84 336 -8
rect 270 -96 336 -84
rect 366 -8 432 4
rect 366 -84 382 -8
rect 416 -84 432 -8
rect 366 -96 432 -84
rect 462 -8 528 4
rect 462 -84 478 -8
rect 512 -84 528 -8
rect 462 -96 528 -84
rect 558 -8 624 4
rect 558 -84 574 -8
rect 608 -84 624 -8
rect 558 -96 624 -84
rect 654 -8 720 4
rect 654 -84 670 -8
rect 704 -84 720 -8
rect 654 -96 720 -84
rect 750 -8 812 4
rect 750 -84 766 -8
rect 800 -84 812 -8
rect 750 -96 812 -84
rect 1214 -58 1276 -46
rect 1214 -434 1226 -58
rect 1260 -434 1276 -58
rect 1214 -446 1276 -434
rect 1306 -58 1372 -46
rect 1306 -434 1322 -58
rect 1356 -434 1372 -58
rect 1306 -446 1372 -434
rect 1402 -58 1464 -46
rect 1402 -434 1418 -58
rect 1452 -434 1464 -58
rect 1402 -446 1464 -434
rect 1536 -58 1598 -46
rect 1536 -434 1548 -58
rect 1582 -434 1598 -58
rect 1536 -446 1598 -434
rect 1628 -58 1694 -46
rect 1628 -434 1644 -58
rect 1678 -434 1694 -58
rect 1628 -446 1694 -434
rect 1724 -58 1790 -46
rect 1724 -434 1740 -58
rect 1774 -434 1790 -58
rect 1724 -446 1790 -434
rect 1820 -58 1886 -46
rect 1820 -434 1836 -58
rect 1870 -434 1886 -58
rect 1820 -446 1886 -434
rect 1916 -58 1978 -46
rect 1916 -434 1932 -58
rect 1966 -434 1978 -58
rect 1916 -446 1978 -434
rect 2050 -58 2112 -46
rect 2050 -434 2062 -58
rect 2096 -434 2112 -58
rect 2050 -446 2112 -434
rect 2142 -58 2208 -46
rect 2142 -434 2158 -58
rect 2192 -434 2208 -58
rect 2142 -446 2208 -434
rect 2238 -58 2300 -46
rect 2238 -434 2254 -58
rect 2288 -434 2300 -58
rect 2238 -446 2300 -434
<< ndiffc >>
rect -2 -898 32 -522
rect 94 -898 128 -522
rect 190 -898 224 -522
rect 286 -898 320 -522
rect 382 -898 416 -522
rect 478 -898 512 -522
rect 574 -898 608 -522
rect 670 -898 704 -522
rect 766 -898 800 -522
rect -2 -1158 32 -1082
rect 94 -1158 128 -1082
rect 190 -1158 224 -1082
rect 286 -1158 320 -1082
rect 382 -1158 416 -1082
rect 478 -1158 512 -1082
rect 574 -1158 608 -1082
rect 670 -1158 704 -1082
rect 766 -1158 800 -1082
rect 1548 -1164 1582 -788
rect 1644 -1164 1678 -788
rect 1740 -1164 1774 -788
rect 1836 -1164 1870 -788
rect 1932 -1164 1966 -788
<< pdiffc >>
rect -2 -84 32 -8
rect 94 -84 128 -8
rect 190 -84 224 -8
rect 286 -84 320 -8
rect 382 -84 416 -8
rect 478 -84 512 -8
rect 574 -84 608 -8
rect 670 -84 704 -8
rect 766 -84 800 -8
rect 1226 -434 1260 -58
rect 1322 -434 1356 -58
rect 1418 -434 1452 -58
rect 1548 -434 1582 -58
rect 1644 -434 1678 -58
rect 1740 -434 1774 -58
rect 1836 -434 1870 -58
rect 1932 -434 1966 -58
rect 2062 -434 2096 -58
rect 2158 -434 2192 -58
rect 2254 -434 2288 -58
<< psubdiff >>
rect -286 4574 -164 4600
rect -286 4500 -262 4574
rect -188 4500 -164 4574
rect -286 4476 -164 4500
rect 262 4574 384 4600
rect 262 4500 286 4574
rect 360 4500 384 4574
rect 262 4476 384 4500
rect 810 4574 932 4600
rect 810 4500 834 4574
rect 908 4500 932 4574
rect 810 4476 932 4500
rect 1358 4574 1480 4600
rect 1358 4500 1382 4574
rect 1456 4500 1480 4574
rect 1358 4476 1480 4500
rect 1906 4574 2028 4600
rect 1906 4500 1930 4574
rect 2004 4500 2028 4574
rect 1906 4476 2028 4500
rect 2454 4574 2576 4600
rect 2454 4500 2478 4574
rect 2552 4500 2576 4574
rect 2454 4476 2576 4500
rect 3002 4574 3124 4600
rect 3002 4500 3026 4574
rect 3100 4500 3124 4574
rect 3002 4476 3124 4500
rect 3550 4574 3672 4600
rect 3550 4500 3574 4574
rect 3648 4500 3672 4574
rect 3550 4476 3672 4500
rect -512 4250 -390 4276
rect -512 4176 -488 4250
rect -414 4176 -390 4250
rect -512 4152 -390 4176
rect 3690 4182 3812 4208
rect 3690 4108 3714 4182
rect 3788 4108 3812 4182
rect 3690 4084 3812 4108
rect -512 3776 -390 3802
rect -512 3702 -488 3776
rect -414 3702 -390 3776
rect -512 3678 -390 3702
rect 3690 3708 3812 3734
rect 3690 3634 3714 3708
rect 3788 3634 3812 3708
rect 3690 3610 3812 3634
rect -512 3302 -390 3328
rect -512 3228 -488 3302
rect -414 3228 -390 3302
rect -512 3204 -390 3228
rect 3690 3234 3812 3260
rect 3690 3160 3714 3234
rect 3788 3160 3812 3234
rect 3690 3136 3812 3160
rect -512 2828 -390 2854
rect -512 2754 -488 2828
rect -414 2754 -390 2828
rect -512 2730 -390 2754
rect 3690 2760 3812 2786
rect 3690 2686 3714 2760
rect 3788 2686 3812 2760
rect 3690 2662 3812 2686
rect -512 2354 -390 2380
rect -512 2280 -488 2354
rect -414 2280 -390 2354
rect -512 2256 -390 2280
rect 3690 2286 3812 2312
rect 3690 2212 3714 2286
rect 3788 2212 3812 2286
rect 3690 2188 3812 2212
rect -512 1880 -390 1906
rect -512 1806 -488 1880
rect -414 1806 -390 1880
rect -512 1782 -390 1806
rect 3690 1810 3812 1836
rect 3690 1736 3714 1810
rect 3788 1736 3812 1810
rect 3690 1712 3812 1736
rect -512 1406 -390 1432
rect -512 1332 -488 1406
rect -414 1332 -390 1406
rect -512 1308 -390 1332
rect 3690 1334 3812 1360
rect 3690 1260 3714 1334
rect 3788 1260 3812 1334
rect 3690 1236 3812 1260
rect -512 932 -390 958
rect -512 858 -488 932
rect -414 858 -390 932
rect -512 834 -390 858
rect 3690 860 3812 886
rect 3690 786 3714 860
rect 3788 786 3812 860
rect 3690 762 3812 786
rect -512 458 -390 484
rect -512 384 -488 458
rect -414 384 -390 458
rect -512 360 -390 384
rect 3688 386 3810 412
rect 3688 312 3712 386
rect 3786 312 3810 386
rect 3688 288 3810 312
rect -512 -88 -390 -62
rect -512 -162 -488 -88
rect -414 -162 -390 -88
rect -512 -186 -390 -162
rect 3688 -86 3810 -60
rect 3688 -160 3712 -86
rect 3786 -160 3810 -86
rect 3688 -184 3810 -160
rect -434 -614 -312 -588
rect -434 -688 -410 -614
rect -336 -688 -312 -614
rect -434 -712 -312 -688
rect 3688 -560 3810 -534
rect 3688 -634 3712 -560
rect 3786 -634 3810 -560
rect 3688 -658 3810 -634
rect -434 -1088 -312 -1062
rect -434 -1162 -410 -1088
rect -336 -1162 -312 -1088
rect -434 -1186 -312 -1162
rect 3688 -1034 3810 -1008
rect 3688 -1108 3712 -1034
rect 3786 -1108 3810 -1034
rect 3688 -1132 3810 -1108
rect -26 -1228 830 -1226
rect -26 -1264 4 -1228
rect 40 -1264 122 -1228
rect 158 -1264 240 -1228
rect 276 -1264 358 -1228
rect 394 -1264 476 -1228
rect 512 -1264 594 -1228
rect 630 -1264 712 -1228
rect 748 -1264 830 -1228
rect -26 -1268 830 -1264
rect 1542 -1324 1566 -1288
rect 1602 -1324 1658 -1288
rect 1694 -1324 1750 -1288
rect 1786 -1324 1842 -1288
rect 1878 -1324 1934 -1288
rect 1970 -1324 1994 -1288
rect 1542 -1326 1994 -1324
rect -506 -1954 -384 -1928
rect -506 -2028 -482 -1954
rect -408 -2028 -384 -1954
rect -506 -2052 -384 -2028
rect 3688 -1984 3810 -1958
rect 3688 -2058 3712 -1984
rect 3786 -2058 3810 -1984
rect 3688 -2082 3810 -2058
rect -506 -2428 -384 -2402
rect -506 -2502 -482 -2428
rect -408 -2502 -384 -2428
rect -506 -2526 -384 -2502
rect 3688 -2458 3810 -2432
rect 3688 -2532 3712 -2458
rect 3786 -2532 3810 -2458
rect 3688 -2556 3810 -2532
rect -506 -2902 -384 -2876
rect -506 -2976 -482 -2902
rect -408 -2976 -384 -2902
rect -506 -3000 -384 -2976
rect 3688 -2932 3810 -2906
rect 3688 -3006 3712 -2932
rect 3786 -3006 3810 -2932
rect 3688 -3030 3810 -3006
rect -506 -3378 -384 -3352
rect -506 -3452 -482 -3378
rect -408 -3452 -384 -3378
rect -506 -3476 -384 -3452
rect 3688 -3406 3810 -3380
rect 3688 -3480 3712 -3406
rect 3786 -3480 3810 -3406
rect 3688 -3504 3810 -3480
rect -506 -3852 -384 -3826
rect -506 -3926 -482 -3852
rect -408 -3926 -384 -3852
rect -506 -3950 -384 -3926
rect 3688 -3880 3810 -3854
rect 3688 -3954 3712 -3880
rect 3786 -3954 3810 -3880
rect 3688 -3978 3810 -3954
rect -506 -4326 -384 -4300
rect -506 -4400 -482 -4326
rect -408 -4400 -384 -4326
rect -506 -4424 -384 -4400
rect 3688 -4354 3810 -4328
rect 3688 -4428 3712 -4354
rect 3786 -4428 3810 -4354
rect 3688 -4452 3810 -4428
rect -506 -4800 -384 -4774
rect -506 -4874 -482 -4800
rect -408 -4874 -384 -4800
rect -506 -4898 -384 -4874
rect 3690 -4828 3812 -4802
rect 3690 -4902 3714 -4828
rect 3788 -4902 3812 -4828
rect 3690 -4926 3812 -4902
rect -506 -5272 -384 -5246
rect -506 -5346 -482 -5272
rect -408 -5346 -384 -5272
rect -506 -5370 -384 -5346
rect 3690 -5302 3812 -5276
rect 3690 -5376 3714 -5302
rect 3788 -5376 3812 -5302
rect 3690 -5400 3812 -5376
rect -506 -5746 -384 -5720
rect -506 -5820 -482 -5746
rect -408 -5820 -384 -5746
rect -506 -5844 -384 -5820
rect 3690 -5776 3812 -5750
rect 3690 -5850 3714 -5776
rect 3788 -5850 3812 -5776
rect 3690 -5874 3812 -5850
rect -116 -6110 6 -6084
rect -116 -6184 -92 -6110
rect -18 -6184 6 -6110
rect -116 -6208 6 -6184
rect 432 -6110 554 -6084
rect 432 -6184 456 -6110
rect 530 -6184 554 -6110
rect 432 -6208 554 -6184
rect 980 -6110 1102 -6084
rect 980 -6184 1004 -6110
rect 1078 -6184 1102 -6110
rect 980 -6208 1102 -6184
rect 1528 -6110 1650 -6084
rect 1528 -6184 1552 -6110
rect 1626 -6184 1650 -6110
rect 1528 -6208 1650 -6184
rect 2076 -6110 2198 -6084
rect 2076 -6184 2100 -6110
rect 2174 -6184 2198 -6110
rect 2076 -6208 2198 -6184
rect 2624 -6110 2746 -6084
rect 2624 -6184 2648 -6110
rect 2722 -6184 2746 -6110
rect 2624 -6208 2746 -6184
rect 3174 -6110 3296 -6084
rect 3174 -6184 3198 -6110
rect 3272 -6184 3296 -6110
rect 3174 -6208 3296 -6184
<< nsubdiff >>
rect 1382 110 2106 118
rect -14 100 958 108
rect -14 66 16 100
rect 50 66 100 100
rect 134 66 184 100
rect 218 66 268 100
rect 302 66 352 100
rect 386 66 436 100
rect 470 66 520 100
rect 554 66 604 100
rect 638 66 688 100
rect 722 66 778 100
rect 812 66 868 100
rect 902 66 958 100
rect 1382 76 1420 110
rect 1454 76 1504 110
rect 1538 76 1588 110
rect 1622 76 1672 110
rect 1706 76 1756 110
rect 1790 76 1840 110
rect 1874 76 1924 110
rect 1958 76 2008 110
rect 2042 76 2106 110
rect 1382 70 2106 76
rect -14 60 958 66
<< psubdiffcont >>
rect -262 4500 -188 4574
rect 286 4500 360 4574
rect 834 4500 908 4574
rect 1382 4500 1456 4574
rect 1930 4500 2004 4574
rect 2478 4500 2552 4574
rect 3026 4500 3100 4574
rect 3574 4500 3648 4574
rect -488 4176 -414 4250
rect 3714 4108 3788 4182
rect -488 3702 -414 3776
rect 3714 3634 3788 3708
rect -488 3228 -414 3302
rect 3714 3160 3788 3234
rect -488 2754 -414 2828
rect 3714 2686 3788 2760
rect -488 2280 -414 2354
rect 3714 2212 3788 2286
rect -488 1806 -414 1880
rect 3714 1736 3788 1810
rect -488 1332 -414 1406
rect 3714 1260 3788 1334
rect -488 858 -414 932
rect 3714 786 3788 860
rect -488 384 -414 458
rect 3712 312 3786 386
rect -488 -162 -414 -88
rect 3712 -160 3786 -86
rect -410 -688 -336 -614
rect 3712 -634 3786 -560
rect -410 -1162 -336 -1088
rect 3712 -1108 3786 -1034
rect 4 -1264 40 -1228
rect 122 -1264 158 -1228
rect 240 -1264 276 -1228
rect 358 -1264 394 -1228
rect 476 -1264 512 -1228
rect 594 -1264 630 -1228
rect 712 -1264 748 -1228
rect 1566 -1324 1602 -1288
rect 1658 -1324 1694 -1288
rect 1750 -1324 1786 -1288
rect 1842 -1324 1878 -1288
rect 1934 -1324 1970 -1288
rect -482 -2028 -408 -1954
rect 3712 -2058 3786 -1984
rect -482 -2502 -408 -2428
rect 3712 -2532 3786 -2458
rect -482 -2976 -408 -2902
rect 3712 -3006 3786 -2932
rect -482 -3452 -408 -3378
rect 3712 -3480 3786 -3406
rect -482 -3926 -408 -3852
rect 3712 -3954 3786 -3880
rect -482 -4400 -408 -4326
rect 3712 -4428 3786 -4354
rect -482 -4874 -408 -4800
rect 3714 -4902 3788 -4828
rect -482 -5346 -408 -5272
rect 3714 -5376 3788 -5302
rect -482 -5820 -408 -5746
rect 3714 -5850 3788 -5776
rect -92 -6184 -18 -6110
rect 456 -6184 530 -6110
rect 1004 -6184 1078 -6110
rect 1552 -6184 1626 -6110
rect 2100 -6184 2174 -6110
rect 2648 -6184 2722 -6110
rect 3198 -6184 3272 -6110
<< nsubdiffcont >>
rect 16 66 50 100
rect 100 66 134 100
rect 184 66 218 100
rect 268 66 302 100
rect 352 66 386 100
rect 436 66 470 100
rect 520 66 554 100
rect 604 66 638 100
rect 688 66 722 100
rect 778 66 812 100
rect 868 66 902 100
rect 1420 76 1454 110
rect 1504 76 1538 110
rect 1588 76 1622 110
rect 1672 76 1706 110
rect 1756 76 1790 110
rect 1840 76 1874 110
rect 1924 76 1958 110
rect 2008 76 2042 110
<< poly >>
rect 48 4 78 30
rect 144 4 174 30
rect 240 4 270 30
rect 336 4 366 30
rect 432 4 462 30
rect 528 4 558 30
rect 624 4 654 30
rect 720 4 750 30
rect 1276 -46 1306 -20
rect 1372 -46 1402 -20
rect 1598 -46 1628 -20
rect 1694 -46 1724 -20
rect 1790 -46 1820 -20
rect 1886 -46 1916 -20
rect 2112 -46 2142 -20
rect 2208 -46 2238 -20
rect 48 -122 78 -96
rect 144 -122 174 -96
rect 240 -122 270 -96
rect 336 -122 366 -96
rect 432 -122 462 -96
rect 528 -122 558 -96
rect 624 -122 654 -96
rect 720 -122 750 -96
rect 48 -154 750 -122
rect 370 -238 428 -154
rect 370 -248 1068 -238
rect 370 -274 1018 -248
rect 1002 -282 1018 -274
rect 1052 -282 1068 -248
rect 1002 -292 1068 -282
rect 164 -334 236 -324
rect 164 -374 180 -334
rect 220 -374 236 -334
rect 164 -384 236 -374
rect 556 -332 628 -322
rect 556 -372 572 -332
rect 612 -372 628 -332
rect 556 -382 628 -372
rect 188 -454 226 -384
rect 572 -454 610 -382
rect 48 -484 366 -454
rect 48 -510 78 -484
rect 144 -510 174 -484
rect 240 -510 270 -484
rect 336 -510 366 -484
rect 432 -484 750 -454
rect 432 -510 462 -484
rect 528 -510 558 -484
rect 624 -510 654 -484
rect 720 -510 750 -484
rect 1276 -462 1306 -446
rect 1372 -462 1402 -446
rect 1276 -492 1402 -462
rect 1598 -462 1628 -446
rect 1694 -462 1724 -446
rect 1598 -492 1724 -462
rect 1276 -626 1306 -492
rect 1690 -558 1724 -492
rect 1658 -568 1724 -558
rect 1658 -602 1674 -568
rect 1708 -602 1724 -568
rect 1658 -612 1724 -602
rect 1276 -636 1342 -626
rect 1276 -670 1292 -636
rect 1326 -670 1342 -636
rect 1276 -680 1342 -670
rect 1598 -776 1628 -750
rect 1694 -776 1724 -612
rect 1790 -462 1820 -446
rect 1886 -462 1916 -446
rect 1790 -492 1916 -462
rect 2112 -462 2142 -446
rect 2208 -462 2238 -446
rect 2112 -492 2238 -462
rect 1790 -626 1824 -492
rect 2204 -626 2238 -492
rect 1790 -636 2082 -626
rect 1790 -670 1808 -636
rect 1842 -670 2082 -636
rect 1790 -680 2082 -670
rect 2172 -636 2238 -626
rect 2172 -670 2188 -636
rect 2222 -670 2238 -636
rect 2172 -680 2238 -670
rect 1790 -776 1820 -680
rect 1886 -776 1916 -750
rect 2026 -752 2082 -680
rect 2026 -762 2372 -752
rect 48 -938 78 -910
rect 144 -938 174 -910
rect 240 -938 270 -910
rect 336 -938 366 -910
rect 432 -938 462 -910
rect 528 -938 558 -910
rect 624 -938 654 -910
rect 720 -938 750 -910
rect 1002 -1000 1068 -990
rect 1002 -1014 1018 -1000
rect 48 -1034 1018 -1014
rect 1052 -1034 1068 -1000
rect 48 -1044 1068 -1034
rect 48 -1070 78 -1044
rect 144 -1070 174 -1044
rect 240 -1070 270 -1044
rect 336 -1070 366 -1044
rect 432 -1070 462 -1044
rect 528 -1070 558 -1044
rect 624 -1070 654 -1044
rect 720 -1070 750 -1044
rect 48 -1196 78 -1170
rect 144 -1196 174 -1170
rect 240 -1196 270 -1170
rect 336 -1196 366 -1170
rect 432 -1196 462 -1170
rect 528 -1196 558 -1170
rect 624 -1196 654 -1170
rect 720 -1196 750 -1170
rect 2026 -796 2322 -762
rect 2356 -796 2372 -762
rect 2026 -808 2372 -796
rect 2306 -832 2372 -808
rect 2306 -866 2322 -832
rect 2356 -866 2372 -832
rect 2306 -876 2372 -866
rect 1598 -1244 1628 -1176
rect 1694 -1202 1724 -1176
rect 1790 -1202 1820 -1176
rect 1886 -1244 1916 -1176
rect 1440 -1254 1916 -1244
rect 1440 -1288 1456 -1254
rect 1490 -1274 1916 -1254
rect 1490 -1288 1506 -1274
rect 1440 -1298 1506 -1288
<< polycont >>
rect 1018 -282 1052 -248
rect 180 -374 220 -334
rect 572 -372 612 -332
rect 1674 -602 1708 -568
rect 1292 -670 1326 -636
rect 1808 -670 1842 -636
rect 2188 -670 2222 -636
rect 1018 -1034 1052 -1000
rect 2322 -796 2356 -762
rect 2322 -866 2356 -832
rect 1456 -1288 1490 -1254
<< locali >>
rect -546 4574 3852 4630
rect -546 4500 -262 4574
rect -188 4500 286 4574
rect 360 4500 834 4574
rect 908 4500 1382 4574
rect 1456 4500 1930 4574
rect 2004 4500 2478 4574
rect 2552 4500 3026 4574
rect 3100 4500 3574 4574
rect 3648 4500 3852 4574
rect -546 4432 3852 4500
rect -546 4250 -348 4432
rect -546 4176 -488 4250
rect -414 4176 -348 4250
rect -546 3776 -348 4176
rect -546 3702 -488 3776
rect -414 3702 -348 3776
rect -546 3302 -348 3702
rect -546 3228 -488 3302
rect -414 3228 -348 3302
rect -546 2828 -348 3228
rect -546 2754 -488 2828
rect -414 2754 -348 2828
rect -546 2354 -348 2754
rect -546 2280 -488 2354
rect -414 2280 -348 2354
rect -546 1880 -348 2280
rect -546 1806 -488 1880
rect -414 1806 -348 1880
rect -546 1406 -348 1806
rect -546 1332 -488 1406
rect -414 1332 -348 1406
rect -546 932 -348 1332
rect -546 858 -488 932
rect -414 858 -348 932
rect -546 464 -348 858
rect 3654 4182 3852 4432
rect 3654 4108 3714 4182
rect 3788 4108 3852 4182
rect 3654 3708 3852 4108
rect 3654 3634 3714 3708
rect 3788 3634 3852 3708
rect 3654 3234 3852 3634
rect 3654 3160 3714 3234
rect 3788 3160 3852 3234
rect 3654 2760 3852 3160
rect 3654 2686 3714 2760
rect 3788 2686 3852 2760
rect 3654 2286 3852 2686
rect 3654 2212 3714 2286
rect 3788 2212 3852 2286
rect 3654 1810 3852 2212
rect 3654 1736 3714 1810
rect 3788 1736 3852 1810
rect 3654 1334 3852 1736
rect 3654 1260 3714 1334
rect 3788 1260 3852 1334
rect 3654 860 3852 1260
rect 3654 786 3714 860
rect 3788 786 3852 860
rect 3654 464 3852 786
rect -546 458 1276 464
rect -546 384 -488 458
rect -414 424 1276 458
rect -414 384 -322 424
rect -546 358 -322 384
rect -258 358 -214 424
rect -150 358 -106 424
rect -42 358 2 424
rect 66 358 110 424
rect 174 358 218 424
rect 282 358 326 424
rect 390 358 434 424
rect 498 358 542 424
rect 606 358 650 424
rect 714 358 758 424
rect 822 358 866 424
rect 930 358 978 424
rect 1042 358 1086 424
rect 1150 358 1194 424
rect 1258 358 1276 424
rect -546 336 1276 358
rect 2028 426 3852 464
rect 2028 424 2270 426
rect 2028 358 2054 424
rect 2118 358 2162 424
rect 2226 360 2270 424
rect 2334 424 3852 426
rect 2334 360 2376 424
rect 2226 358 2376 360
rect 2440 358 2486 424
rect 2550 358 2594 424
rect 2658 358 2700 424
rect 2764 358 2810 424
rect 2874 358 2918 424
rect 2982 358 3026 424
rect 3090 358 3134 424
rect 3198 358 3242 424
rect 3306 358 3354 424
rect 3418 358 3462 424
rect 3526 358 3570 424
rect 3634 386 3852 424
rect 3634 358 3712 386
rect -546 -88 -348 336
rect 2028 334 3712 358
rect 3654 312 3712 334
rect 3786 312 3852 386
rect 2558 152 2650 190
rect 2688 152 2726 190
rect 2764 152 2802 190
rect 2840 152 2878 190
rect 2916 152 3008 190
rect 2558 146 3008 152
rect -14 100 958 108
rect -14 66 16 100
rect 50 66 100 100
rect 134 66 184 100
rect 218 66 268 100
rect 302 66 352 100
rect 386 66 436 100
rect 470 66 520 100
rect 554 66 604 100
rect 638 66 688 100
rect 722 66 778 100
rect 812 66 868 100
rect 902 66 958 100
rect -14 60 958 66
rect 1138 100 1324 112
rect 1138 86 1246 100
rect -546 -162 -488 -88
rect -414 -162 -348 -88
rect -2 42 800 60
rect -2 -8 32 42
rect -2 -100 32 -84
rect 94 -8 128 8
rect -546 -458 -348 -162
rect 94 -160 128 -84
rect 190 -8 224 42
rect 190 -100 224 -84
rect 286 -8 320 8
rect 286 -160 320 -84
rect 382 -8 416 42
rect 382 -100 416 -84
rect 478 -8 512 8
rect 94 -194 320 -160
rect 164 -334 236 -324
rect 164 -374 180 -334
rect 220 -374 236 -334
rect 164 -384 236 -374
rect 286 -418 320 -194
rect -134 -452 320 -418
rect -546 -614 -198 -458
rect -546 -688 -410 -614
rect -336 -688 -198 -614
rect -546 -1088 -198 -688
rect -546 -1162 -410 -1088
rect -336 -1162 -198 -1088
rect -546 -1222 -198 -1162
rect -134 -1172 -74 -452
rect -2 -522 32 -506
rect -2 -948 32 -898
rect 94 -522 128 -452
rect 94 -914 128 -898
rect 190 -522 224 -506
rect 190 -948 224 -898
rect 286 -522 320 -452
rect 478 -160 512 -84
rect 574 -8 608 42
rect 574 -100 608 -84
rect 670 -8 704 8
rect 670 -160 704 -84
rect 766 -8 800 42
rect 1138 52 1174 86
rect 1208 52 1246 86
rect 1138 36 1246 52
rect 1310 36 1324 100
rect 1382 110 2106 118
rect 1382 76 1420 110
rect 1454 76 1504 110
rect 1538 76 1588 110
rect 1622 76 1672 110
rect 1706 76 1756 110
rect 1790 76 1840 110
rect 1874 76 1924 110
rect 1958 76 2008 110
rect 2042 76 2106 110
rect 1382 70 2106 76
rect 2198 100 2384 112
rect 2198 86 2304 100
rect 1718 36 1808 70
rect 2198 52 2232 86
rect 2266 52 2304 86
rect 2198 36 2304 52
rect 2368 36 2384 100
rect 1138 26 1324 36
rect 1138 -8 1452 26
rect 766 -100 800 -84
rect 1226 -58 1260 -8
rect 478 -194 704 -160
rect 478 -416 512 -194
rect 1002 -248 1068 -238
rect 1002 -282 1018 -248
rect 1052 -282 1068 -248
rect 556 -332 628 -322
rect 556 -372 572 -332
rect 612 -372 628 -332
rect 556 -382 628 -372
rect 478 -450 926 -416
rect 286 -914 320 -898
rect 382 -522 416 -506
rect 382 -948 416 -898
rect 478 -522 512 -450
rect 478 -914 512 -898
rect 574 -522 608 -506
rect 574 -948 608 -898
rect 670 -522 704 -450
rect 670 -914 704 -898
rect 766 -522 800 -506
rect 766 -948 800 -898
rect -2 -984 800 -948
rect -2 -1082 32 -984
rect -546 -1256 -530 -1222
rect -496 -1256 -458 -1222
rect -424 -1256 -386 -1222
rect -352 -1256 -314 -1222
rect -280 -1256 -242 -1222
rect -208 -1256 -198 -1222
rect -546 -1294 -198 -1256
rect -546 -1328 -530 -1294
rect -496 -1328 -458 -1294
rect -424 -1328 -386 -1294
rect -352 -1328 -314 -1294
rect -280 -1328 -242 -1294
rect -208 -1328 -198 -1294
rect -546 -1366 -198 -1328
rect -546 -1400 -530 -1366
rect -496 -1400 -458 -1366
rect -424 -1400 -386 -1366
rect -352 -1400 -314 -1366
rect -280 -1400 -242 -1366
rect -208 -1400 -198 -1366
rect -546 -1438 -198 -1400
rect -546 -1472 -530 -1438
rect -496 -1472 -458 -1438
rect -424 -1472 -386 -1438
rect -352 -1472 -314 -1438
rect -280 -1472 -242 -1438
rect -208 -1472 -198 -1438
rect -546 -1486 -198 -1472
rect -546 -1914 -348 -1486
rect -122 -1512 -88 -1172
rect -2 -1174 32 -1158
rect 94 -1082 128 -1064
rect 94 -1212 128 -1158
rect 190 -1082 224 -984
rect 190 -1174 224 -1158
rect 286 -1082 320 -1066
rect 286 -1212 320 -1158
rect 382 -1082 416 -984
rect 382 -1174 416 -1158
rect 478 -1082 512 -1066
rect 478 -1212 512 -1158
rect 574 -1082 608 -984
rect 574 -1174 608 -1158
rect 670 -1082 704 -1066
rect 670 -1212 704 -1158
rect 766 -1082 800 -984
rect 766 -1174 800 -1158
rect 94 -1226 704 -1212
rect -26 -1228 830 -1226
rect -26 -1264 4 -1228
rect 40 -1264 122 -1228
rect 158 -1264 240 -1228
rect 276 -1264 358 -1228
rect 394 -1264 476 -1228
rect 512 -1264 594 -1228
rect 630 -1264 712 -1228
rect 748 -1264 830 -1228
rect -26 -1268 830 -1264
rect 866 -1278 926 -450
rect 1002 -1000 1068 -282
rect 1226 -568 1260 -434
rect 1322 -58 1356 -42
rect 1322 -500 1356 -434
rect 1418 -58 1452 -8
rect 1418 -450 1452 -434
rect 1548 2 1966 36
rect 2198 26 2384 36
rect 1548 -58 1582 2
rect 1548 -450 1582 -434
rect 1644 -58 1678 -42
rect 1644 -500 1678 -434
rect 1740 -58 1774 2
rect 1740 -450 1774 -434
rect 1836 -58 1870 -42
rect 1322 -534 1678 -500
rect 1836 -500 1870 -434
rect 1932 -58 1966 2
rect 1932 -450 1966 -434
rect 2062 -8 2384 26
rect 2062 -58 2096 -8
rect 2062 -450 2096 -434
rect 2158 -58 2192 -42
rect 2158 -500 2192 -434
rect 1836 -534 2192 -500
rect 2254 -58 2288 -8
rect 3654 -86 3852 312
rect 3654 -160 3712 -86
rect 3786 -160 3852 -86
rect 2288 -326 2558 -192
rect 3176 -234 3306 -230
rect 3008 -236 3306 -234
rect 3008 -270 3188 -236
rect 3222 -270 3260 -236
rect 3294 -270 3306 -236
rect 3008 -272 3306 -270
rect 3176 -276 3306 -272
rect 2254 -568 2288 -434
rect 3654 -560 3852 -160
rect 1210 -602 1624 -568
rect 1658 -602 1674 -568
rect 1708 -602 2300 -568
rect 1002 -1034 1018 -1000
rect 1052 -1034 1068 -1000
rect 1002 -1278 1068 -1034
rect 1274 -670 1292 -636
rect 1326 -670 1342 -636
rect 1274 -1278 1342 -670
rect 1392 -946 1478 -602
rect 1590 -636 1624 -602
rect 1590 -670 1808 -636
rect 1842 -670 1858 -636
rect 1392 -980 1418 -946
rect 1452 -980 1478 -946
rect 1392 -1018 1478 -980
rect 1392 -1082 1402 -1018
rect 1466 -1082 1478 -1018
rect 1392 -1094 1478 -1082
rect 1548 -788 1582 -772
rect -122 -1518 8 -1512
rect -122 -1552 -110 -1518
rect -76 -1552 -38 -1518
rect -4 -1552 8 -1518
rect -122 -1558 8 -1552
rect 882 -1586 916 -1278
rect 784 -1592 916 -1586
rect 784 -1626 796 -1592
rect 830 -1626 868 -1592
rect 902 -1626 916 -1592
rect 784 -1632 916 -1626
rect 1018 -1660 1052 -1278
rect 1290 -1512 1324 -1278
rect 1440 -1288 1456 -1254
rect 1490 -1288 1506 -1254
rect 1548 -1288 1582 -1164
rect 1644 -788 1678 -670
rect 1902 -704 1936 -602
rect 1836 -738 1936 -704
rect 1644 -1180 1678 -1164
rect 1740 -788 1774 -772
rect 1740 -1288 1774 -1164
rect 1836 -788 1870 -738
rect 1836 -1180 1870 -1164
rect 1932 -788 1966 -772
rect 2016 -946 2102 -602
rect 2016 -980 2042 -946
rect 2076 -980 2102 -946
rect 2016 -1018 2102 -980
rect 2016 -1082 2026 -1018
rect 2090 -1082 2102 -1018
rect 2016 -1094 2102 -1082
rect 2136 -670 2188 -636
rect 2222 -670 2238 -636
rect 3654 -634 3712 -560
rect 3786 -634 3852 -560
rect 2136 -680 2238 -670
rect 1932 -1288 1966 -1164
rect 1244 -1518 1374 -1512
rect 1244 -1552 1256 -1518
rect 1290 -1552 1328 -1518
rect 1362 -1552 1374 -1518
rect 1244 -1558 1374 -1552
rect 936 -1666 1068 -1660
rect 936 -1700 948 -1666
rect 982 -1700 1020 -1666
rect 1054 -1700 1068 -1666
rect 936 -1706 1068 -1700
rect 1440 -1734 1506 -1288
rect 1542 -1324 1566 -1288
rect 1602 -1324 1658 -1288
rect 1694 -1324 1750 -1288
rect 1786 -1324 1842 -1288
rect 1878 -1324 1934 -1288
rect 1970 -1324 1994 -1288
rect 2136 -1314 2212 -680
rect 2306 -762 2372 -752
rect 2306 -796 2322 -762
rect 2356 -796 2372 -762
rect 2306 -832 2372 -796
rect 2306 -866 2322 -832
rect 2356 -866 2372 -832
rect 2306 -1004 2372 -866
rect 2306 -1140 2560 -1004
rect 3654 -1034 3852 -634
rect 3176 -1046 3306 -1042
rect 3008 -1048 3306 -1046
rect 3008 -1082 3188 -1048
rect 3222 -1082 3260 -1048
rect 3294 -1082 3306 -1048
rect 3008 -1084 3306 -1082
rect 3176 -1088 3306 -1084
rect 3654 -1108 3712 -1034
rect 3786 -1108 3852 -1034
rect 3654 -1222 3852 -1108
rect 3654 -1256 3668 -1222
rect 3702 -1256 3740 -1222
rect 3774 -1256 3812 -1222
rect 3846 -1256 3852 -1222
rect 3654 -1294 3852 -1256
rect 1542 -1326 1994 -1324
rect 2154 -1586 2188 -1314
rect 3654 -1328 3668 -1294
rect 3702 -1328 3740 -1294
rect 3774 -1328 3812 -1294
rect 3846 -1328 3852 -1294
rect 3654 -1366 3852 -1328
rect 3654 -1400 3668 -1366
rect 3702 -1400 3740 -1366
rect 3774 -1400 3812 -1366
rect 3846 -1400 3852 -1366
rect 3654 -1438 3852 -1400
rect 3654 -1472 3668 -1438
rect 3702 -1472 3740 -1438
rect 3774 -1472 3812 -1438
rect 3846 -1472 3852 -1438
rect 3654 -1510 3852 -1472
rect 3654 -1544 3668 -1510
rect 3702 -1544 3740 -1510
rect 3774 -1544 3812 -1510
rect 3846 -1544 3852 -1510
rect 2102 -1592 2232 -1586
rect 2102 -1626 2114 -1592
rect 2148 -1626 2186 -1592
rect 2220 -1626 2232 -1592
rect 2102 -1632 2232 -1626
rect 1440 -1740 1572 -1734
rect 1440 -1774 1452 -1740
rect 1486 -1774 1524 -1740
rect 1558 -1774 1572 -1740
rect 1440 -1780 1572 -1774
rect 3654 -1912 3852 -1544
rect -546 -1954 1346 -1914
rect -546 -2028 -482 -1954
rect -408 -2020 -252 -1954
rect -188 -2020 -144 -1954
rect -80 -2020 -36 -1954
rect 28 -2020 72 -1954
rect 136 -2020 180 -1954
rect 244 -2020 288 -1954
rect 352 -2020 396 -1954
rect 460 -2020 504 -1954
rect 568 -2020 612 -1954
rect 676 -2020 720 -1954
rect 784 -2020 828 -1954
rect 892 -2020 936 -1954
rect 1000 -2020 1048 -1954
rect 1112 -2020 1156 -1954
rect 1220 -2020 1264 -1954
rect 1328 -2020 1346 -1954
rect -408 -2028 1346 -2020
rect -546 -2042 1346 -2028
rect 2028 -1952 3852 -1912
rect 2028 -2018 2056 -1952
rect 2120 -2018 2164 -1952
rect 2228 -2018 2272 -1952
rect 2336 -2018 2380 -1952
rect 2444 -2018 2488 -1952
rect 2552 -2018 2596 -1952
rect 2660 -2018 2704 -1952
rect 2768 -2018 2812 -1952
rect 2876 -2018 2920 -1952
rect 2984 -2018 3028 -1952
rect 3092 -2018 3136 -1952
rect 3200 -2018 3244 -1952
rect 3308 -2018 3356 -1952
rect 3420 -2018 3464 -1952
rect 3528 -2018 3572 -1952
rect 3636 -1984 3852 -1952
rect 3636 -2018 3712 -1984
rect 2028 -2040 3712 -2018
rect -546 -2428 -348 -2042
rect -546 -2502 -482 -2428
rect -408 -2502 -348 -2428
rect -546 -2902 -348 -2502
rect -546 -2976 -482 -2902
rect -408 -2976 -348 -2902
rect -546 -3378 -348 -2976
rect -546 -3452 -482 -3378
rect -408 -3452 -348 -3378
rect -546 -3852 -348 -3452
rect -546 -3926 -482 -3852
rect -408 -3926 -348 -3852
rect -546 -4326 -348 -3926
rect -546 -4400 -482 -4326
rect -408 -4400 -348 -4326
rect -546 -4800 -348 -4400
rect -546 -4874 -482 -4800
rect -408 -4874 -348 -4800
rect -546 -5272 -348 -4874
rect -546 -5346 -482 -5272
rect -408 -5346 -348 -5272
rect -546 -5746 -348 -5346
rect -546 -5820 -482 -5746
rect -408 -5820 -348 -5746
rect -546 -6042 -348 -5820
rect 3654 -2058 3712 -2040
rect 3786 -2058 3852 -1984
rect 3654 -2458 3852 -2058
rect 3654 -2532 3712 -2458
rect 3786 -2532 3852 -2458
rect 3654 -2932 3852 -2532
rect 3654 -3006 3712 -2932
rect 3786 -3006 3852 -2932
rect 3654 -3406 3852 -3006
rect 3654 -3480 3712 -3406
rect 3786 -3480 3852 -3406
rect 3654 -3880 3852 -3480
rect 3654 -3954 3712 -3880
rect 3786 -3954 3852 -3880
rect 3654 -4354 3852 -3954
rect 3654 -4428 3712 -4354
rect 3786 -4428 3852 -4354
rect 3654 -4828 3852 -4428
rect 3654 -4902 3714 -4828
rect 3788 -4902 3852 -4828
rect 3654 -5302 3852 -4902
rect 3654 -5376 3714 -5302
rect 3788 -5376 3852 -5302
rect 3654 -5776 3852 -5376
rect 3654 -5850 3714 -5776
rect 3788 -5850 3852 -5776
rect 3654 -6042 3852 -5850
rect -546 -6110 3852 -6042
rect -546 -6184 -92 -6110
rect -18 -6184 456 -6110
rect 530 -6184 1004 -6110
rect 1078 -6184 1552 -6110
rect 1626 -6184 2100 -6110
rect 2174 -6184 2648 -6110
rect 2722 -6184 3198 -6110
rect 3272 -6184 3852 -6110
rect -546 -6240 3852 -6184
<< viali >>
rect -322 358 -258 424
rect -214 358 -150 424
rect -106 358 -42 424
rect 2 358 66 424
rect 110 358 174 424
rect 218 358 282 424
rect 326 358 390 424
rect 434 358 498 424
rect 542 358 606 424
rect 650 358 714 424
rect 758 358 822 424
rect 866 358 930 424
rect 978 358 1042 424
rect 1086 358 1150 424
rect 1194 358 1258 424
rect 2054 358 2118 424
rect 2162 358 2226 424
rect 2270 360 2334 426
rect 2376 358 2440 424
rect 2486 358 2550 424
rect 2594 358 2658 424
rect 2700 358 2764 424
rect 2810 358 2874 424
rect 2918 358 2982 424
rect 3026 358 3090 424
rect 3134 358 3198 424
rect 3242 358 3306 424
rect 3354 358 3418 424
rect 3462 358 3526 424
rect 3570 358 3634 424
rect 2650 152 2688 190
rect 2726 152 2764 190
rect 2802 152 2840 190
rect 2878 152 2916 190
rect 16 66 50 100
rect 100 66 134 100
rect 184 66 218 100
rect 268 66 302 100
rect 352 66 386 100
rect 436 66 470 100
rect 520 66 554 100
rect 604 66 638 100
rect 688 66 722 100
rect 778 66 812 100
rect 868 66 902 100
rect 180 -374 220 -334
rect 1174 52 1208 86
rect 1246 36 1310 100
rect 1420 76 1454 110
rect 1504 76 1538 110
rect 1588 76 1622 110
rect 1672 76 1706 110
rect 1756 76 1790 110
rect 1840 76 1874 110
rect 1924 76 1958 110
rect 2008 76 2042 110
rect 2232 52 2266 86
rect 2304 36 2368 100
rect 572 -372 612 -332
rect -530 -1256 -496 -1222
rect -458 -1256 -424 -1222
rect -386 -1256 -352 -1222
rect -314 -1256 -280 -1222
rect -242 -1256 -208 -1222
rect -530 -1328 -496 -1294
rect -458 -1328 -424 -1294
rect -386 -1328 -352 -1294
rect -314 -1328 -280 -1294
rect -242 -1328 -208 -1294
rect -530 -1400 -496 -1366
rect -458 -1400 -424 -1366
rect -386 -1400 -352 -1366
rect -314 -1400 -280 -1366
rect -242 -1400 -208 -1366
rect -530 -1472 -496 -1438
rect -458 -1472 -424 -1438
rect -386 -1472 -352 -1438
rect -314 -1472 -280 -1438
rect -242 -1472 -208 -1438
rect 4 -1264 40 -1228
rect 122 -1264 158 -1228
rect 240 -1264 276 -1228
rect 358 -1264 394 -1228
rect 476 -1264 512 -1228
rect 594 -1264 630 -1228
rect 712 -1264 748 -1228
rect 3188 -270 3222 -236
rect 3260 -270 3294 -236
rect 2642 -548 2676 -514
rect 2714 -548 2748 -514
rect 2794 -548 2828 -514
rect 2868 -548 2902 -514
rect 1418 -980 1452 -946
rect 1402 -1082 1466 -1018
rect -110 -1552 -76 -1518
rect -38 -1552 -4 -1518
rect 796 -1626 830 -1592
rect 868 -1626 902 -1592
rect 2042 -980 2076 -946
rect 2026 -1082 2090 -1018
rect 2650 -656 2688 -622
rect 2726 -656 2764 -622
rect 2802 -656 2840 -622
rect 2878 -656 2916 -622
rect 1256 -1552 1290 -1518
rect 1328 -1552 1362 -1518
rect 948 -1700 982 -1666
rect 1020 -1700 1054 -1666
rect 1566 -1324 1602 -1288
rect 1658 -1324 1694 -1288
rect 1750 -1324 1786 -1288
rect 1842 -1324 1878 -1288
rect 1934 -1324 1970 -1288
rect 3188 -1082 3222 -1048
rect 3260 -1082 3294 -1048
rect 3668 -1256 3702 -1222
rect 3740 -1256 3774 -1222
rect 3812 -1256 3846 -1222
rect 3668 -1328 3702 -1294
rect 3740 -1328 3774 -1294
rect 3812 -1328 3846 -1294
rect 2642 -1366 2676 -1332
rect 2714 -1368 2748 -1334
rect 2794 -1370 2828 -1336
rect 2870 -1366 2904 -1332
rect 3668 -1400 3702 -1366
rect 3740 -1400 3774 -1366
rect 3812 -1400 3846 -1366
rect 3668 -1472 3702 -1438
rect 3740 -1472 3774 -1438
rect 3812 -1472 3846 -1438
rect 3668 -1544 3702 -1510
rect 3740 -1544 3774 -1510
rect 3812 -1544 3846 -1510
rect 2114 -1626 2148 -1592
rect 2186 -1626 2220 -1592
rect 1452 -1774 1486 -1740
rect 1524 -1774 1558 -1740
rect -252 -2020 -188 -1954
rect -144 -2020 -80 -1954
rect -36 -2020 28 -1954
rect 72 -2020 136 -1954
rect 180 -2020 244 -1954
rect 288 -2020 352 -1954
rect 396 -2020 460 -1954
rect 504 -2020 568 -1954
rect 612 -2020 676 -1954
rect 720 -2020 784 -1954
rect 828 -2020 892 -1954
rect 936 -2020 1000 -1954
rect 1048 -2020 1112 -1954
rect 1156 -2020 1220 -1954
rect 1264 -2020 1328 -1954
rect 2056 -2018 2120 -1952
rect 2164 -2018 2228 -1952
rect 2272 -2018 2336 -1952
rect 2380 -2018 2444 -1952
rect 2488 -2018 2552 -1952
rect 2596 -2018 2660 -1952
rect 2704 -2018 2768 -1952
rect 2812 -2018 2876 -1952
rect 2920 -2018 2984 -1952
rect 3028 -2018 3092 -1952
rect 3136 -2018 3200 -1952
rect 3244 -2018 3308 -1952
rect 3356 -2018 3420 -1952
rect 3464 -2018 3528 -1952
rect 3572 -2018 3636 -1952
<< metal1 >>
rect -348 424 1276 464
rect -348 358 -322 424
rect -258 358 -214 424
rect -150 358 -106 424
rect -42 358 2 424
rect 66 358 110 424
rect 174 358 218 424
rect 282 358 326 424
rect 390 358 434 424
rect 498 358 542 424
rect 606 358 650 424
rect 718 358 758 424
rect 826 358 866 424
rect 934 358 978 424
rect 1042 358 1086 424
rect 1150 358 1194 424
rect 1258 358 1276 424
rect -348 336 1276 358
rect 2028 426 3652 464
rect 2028 424 2270 426
rect 2334 424 3652 426
rect 2028 358 2054 424
rect 2118 358 2162 424
rect 2226 358 2270 424
rect 2334 358 2376 424
rect 2442 358 2486 424
rect 2550 358 2594 424
rect 2658 358 2700 424
rect 2766 358 2810 424
rect 2874 358 2918 424
rect 2982 358 3026 424
rect 3094 358 3134 424
rect 3202 358 3242 424
rect 3310 358 3354 424
rect 3418 358 3462 424
rect 3526 358 3570 424
rect 3634 358 3652 424
rect 2028 336 3652 358
rect -714 190 3920 300
rect -714 162 2650 190
rect -14 100 958 162
rect -14 66 16 100
rect 50 66 100 100
rect 134 66 184 100
rect 218 66 268 100
rect 302 66 352 100
rect 386 66 436 100
rect 470 66 520 100
rect 554 66 604 100
rect 638 66 688 100
rect 722 66 778 100
rect 812 66 868 100
rect 902 66 958 100
rect -14 60 958 66
rect 1138 100 1324 112
rect 1138 36 1150 100
rect 1214 36 1246 100
rect 1310 36 1324 100
rect 1382 110 2106 162
rect 2556 152 2650 162
rect 2688 152 2726 190
rect 2764 152 2802 190
rect 2840 152 2878 190
rect 2916 162 3920 190
rect 2916 152 3090 162
rect 2556 146 3090 152
rect 1382 76 1420 110
rect 1454 76 1504 110
rect 1538 76 1588 110
rect 1622 76 1672 110
rect 1706 76 1756 110
rect 1790 76 1840 110
rect 1874 76 1924 110
rect 1958 76 2008 110
rect 2042 76 2106 110
rect 1382 70 2106 76
rect 2198 100 2384 112
rect 1138 26 1324 36
rect 2198 36 2208 100
rect 2272 36 2304 100
rect 2368 36 2384 100
rect 2198 26 2384 36
rect -714 -272 296 -244
rect 268 -322 296 -272
rect -714 -334 236 -324
rect -714 -352 180 -334
rect 164 -374 180 -352
rect 220 -374 236 -334
rect 268 -332 628 -322
rect 268 -352 572 -332
rect 164 -384 236 -374
rect 556 -372 572 -352
rect 612 -372 628 -332
rect 556 -382 628 -372
rect 2428 -514 2966 -506
rect 2428 -548 2642 -514
rect 2676 -548 2714 -514
rect 2748 -548 2794 -514
rect 2828 -548 2868 -514
rect 2902 -548 2966 -514
rect 2428 -560 2966 -548
rect 1392 -922 1478 -912
rect 1392 -986 1402 -922
rect 1466 -986 1478 -922
rect 1392 -1018 1478 -986
rect 1392 -1082 1402 -1018
rect 1466 -1082 1478 -1018
rect 1392 -1094 1478 -1082
rect 2016 -922 2102 -912
rect 2016 -986 2026 -922
rect 2090 -986 2102 -922
rect 2016 -1018 2102 -986
rect 2016 -1082 2026 -1018
rect 2090 -1082 2102 -1018
rect 2016 -1094 2102 -1082
rect -546 -1222 -198 -1202
rect -546 -1256 -530 -1222
rect -496 -1256 -458 -1222
rect -424 -1256 -386 -1222
rect -352 -1256 -314 -1222
rect -280 -1256 -242 -1222
rect -208 -1256 -198 -1222
rect -546 -1294 -198 -1256
rect -546 -1326 -530 -1294
rect -714 -1328 -530 -1326
rect -496 -1328 -458 -1294
rect -424 -1328 -386 -1294
rect -352 -1328 -314 -1294
rect -280 -1328 -242 -1294
rect -208 -1326 -198 -1294
rect -48 -1228 832 -1222
rect -48 -1264 4 -1228
rect 40 -1264 122 -1228
rect 158 -1264 240 -1228
rect 276 -1264 358 -1228
rect 394 -1264 476 -1228
rect 512 -1264 594 -1228
rect 630 -1264 712 -1228
rect 748 -1264 832 -1228
rect -48 -1326 832 -1264
rect 1542 -1288 1994 -1282
rect 1542 -1324 1566 -1288
rect 1602 -1324 1658 -1288
rect 1694 -1324 1750 -1288
rect 1786 -1324 1842 -1288
rect 1878 -1324 1934 -1288
rect 1970 -1324 1994 -1288
rect 1542 -1326 1994 -1324
rect 2428 -1326 2510 -560
rect 3008 -608 3090 146
rect 3176 -236 3920 -230
rect 3176 -270 3188 -236
rect 3222 -270 3260 -236
rect 3294 -270 3920 -236
rect 3176 -276 3920 -270
rect 2558 -622 3090 -608
rect 2558 -656 2650 -622
rect 2688 -656 2726 -622
rect 2764 -656 2802 -622
rect 2840 -656 2878 -622
rect 2916 -656 3090 -622
rect 2558 -662 3090 -656
rect 3176 -1048 3920 -1042
rect 3176 -1082 3188 -1048
rect 3222 -1082 3260 -1048
rect 3294 -1082 3920 -1048
rect 3176 -1088 3920 -1082
rect 3654 -1222 3852 -1202
rect 3654 -1256 3668 -1222
rect 3702 -1256 3740 -1222
rect 3774 -1256 3812 -1222
rect 3846 -1256 3852 -1222
rect 3654 -1294 3852 -1256
rect 3654 -1326 3668 -1294
rect -208 -1328 3668 -1326
rect 3702 -1328 3740 -1294
rect 3774 -1328 3812 -1294
rect 3846 -1326 3852 -1294
rect 3846 -1328 3920 -1326
rect -714 -1332 3920 -1328
rect -714 -1366 2642 -1332
rect 2676 -1334 2870 -1332
rect 2676 -1366 2714 -1334
rect -714 -1400 -530 -1366
rect -496 -1400 -458 -1366
rect -424 -1400 -386 -1366
rect -352 -1400 -314 -1366
rect -280 -1400 -242 -1366
rect -208 -1368 2714 -1366
rect 2748 -1336 2870 -1334
rect 2748 -1368 2794 -1336
rect -208 -1370 2794 -1368
rect 2828 -1366 2870 -1336
rect 2904 -1366 3920 -1332
rect 2828 -1370 3668 -1366
rect -208 -1400 3668 -1370
rect 3702 -1400 3740 -1366
rect 3774 -1400 3812 -1366
rect 3846 -1400 3920 -1366
rect -714 -1438 3920 -1400
rect -714 -1472 -530 -1438
rect -496 -1472 -458 -1438
rect -424 -1472 -386 -1438
rect -352 -1472 -314 -1438
rect -280 -1472 -242 -1438
rect -208 -1472 3668 -1438
rect 3702 -1472 3740 -1438
rect 3774 -1472 3812 -1438
rect 3846 -1472 3920 -1438
rect -714 -1484 3920 -1472
rect 3654 -1510 3852 -1484
rect -122 -1518 1374 -1512
rect -122 -1552 -110 -1518
rect -76 -1552 -38 -1518
rect -4 -1552 1256 -1518
rect 1290 -1552 1328 -1518
rect 1362 -1552 1374 -1518
rect -122 -1558 1374 -1552
rect 3654 -1544 3668 -1510
rect 3702 -1544 3740 -1510
rect 3774 -1544 3812 -1510
rect 3846 -1544 3852 -1510
rect 3654 -1556 3852 -1544
rect 784 -1592 2232 -1586
rect 784 -1626 796 -1592
rect 830 -1626 868 -1592
rect 902 -1626 2114 -1592
rect 2148 -1626 2186 -1592
rect 2220 -1626 2232 -1592
rect 784 -1632 2232 -1626
rect -716 -1666 3920 -1660
rect -716 -1700 948 -1666
rect 982 -1700 1020 -1666
rect 1054 -1700 3920 -1666
rect -716 -1706 3920 -1700
rect -716 -1740 3920 -1734
rect -716 -1774 1452 -1740
rect 1486 -1774 1524 -1740
rect 1558 -1774 3920 -1740
rect -716 -1780 3920 -1774
rect -278 -1954 1346 -1914
rect -278 -2020 -252 -1954
rect -188 -2020 -144 -1954
rect -80 -2020 -36 -1954
rect 28 -2020 72 -1954
rect 136 -2020 180 -1954
rect 244 -2020 288 -1954
rect 352 -2020 396 -1954
rect 460 -2020 504 -1954
rect 568 -2020 612 -1954
rect 676 -2020 720 -1954
rect 788 -2020 828 -1954
rect 896 -2020 936 -1954
rect 1004 -2020 1048 -1954
rect 1112 -2020 1156 -1954
rect 1220 -2020 1264 -1954
rect 1328 -2020 1346 -1954
rect -278 -2042 1346 -2020
rect 2030 -1952 3654 -1912
rect 2030 -2018 2056 -1952
rect 2120 -2018 2164 -1952
rect 2228 -2018 2272 -1952
rect 2336 -2018 2380 -1952
rect 2444 -2018 2488 -1952
rect 2552 -2018 2596 -1952
rect 2660 -2018 2704 -1952
rect 2768 -2018 2812 -1952
rect 2876 -2018 2920 -1952
rect 2984 -2018 3028 -1952
rect 3096 -2018 3136 -1952
rect 3204 -2018 3244 -1952
rect 3312 -2018 3356 -1952
rect 3420 -2018 3464 -1952
rect 3528 -2018 3572 -1952
rect 3636 -2018 3654 -1952
rect 2030 -2040 3654 -2018
<< via1 >>
rect -322 358 -258 424
rect -214 358 -150 424
rect -106 358 -42 424
rect 2 358 66 424
rect 110 358 174 424
rect 218 358 282 424
rect 326 358 390 424
rect 434 358 498 424
rect 542 358 606 424
rect 650 358 714 424
rect 714 358 718 424
rect 758 358 822 424
rect 822 358 826 424
rect 866 358 930 424
rect 930 358 934 424
rect 978 358 1042 424
rect 1086 358 1150 424
rect 1194 358 1258 424
rect 2054 358 2118 424
rect 2162 358 2226 424
rect 2270 360 2334 424
rect 2270 358 2334 360
rect 2378 358 2440 424
rect 2440 358 2442 424
rect 2486 358 2550 424
rect 2594 358 2658 424
rect 2702 358 2764 424
rect 2764 358 2766 424
rect 2810 358 2874 424
rect 2918 358 2982 424
rect 3026 358 3090 424
rect 3090 358 3094 424
rect 3134 358 3198 424
rect 3198 358 3202 424
rect 3242 358 3306 424
rect 3306 358 3310 424
rect 3354 358 3418 424
rect 3462 358 3526 424
rect 3570 358 3634 424
rect 1150 86 1214 100
rect 1150 52 1174 86
rect 1174 52 1208 86
rect 1208 52 1214 86
rect 1150 36 1214 52
rect 1246 36 1310 100
rect 2208 86 2272 100
rect 2208 52 2232 86
rect 2232 52 2266 86
rect 2266 52 2272 86
rect 2208 36 2272 52
rect 2304 36 2368 100
rect 1402 -946 1466 -922
rect 1402 -980 1418 -946
rect 1418 -980 1452 -946
rect 1452 -980 1466 -946
rect 1402 -986 1466 -980
rect 1402 -1082 1466 -1018
rect 2026 -946 2090 -922
rect 2026 -980 2042 -946
rect 2042 -980 2076 -946
rect 2076 -980 2090 -946
rect 2026 -986 2090 -980
rect 2026 -1082 2090 -1018
rect -252 -2020 -188 -1954
rect -144 -2020 -80 -1954
rect -36 -2020 28 -1954
rect 72 -2020 136 -1954
rect 180 -2020 244 -1954
rect 288 -2020 352 -1954
rect 396 -2020 460 -1954
rect 504 -2020 568 -1954
rect 612 -2020 676 -1954
rect 720 -2020 784 -1954
rect 784 -2020 788 -1954
rect 828 -2020 892 -1954
rect 892 -2020 896 -1954
rect 936 -2020 1000 -1954
rect 1000 -2020 1004 -1954
rect 1048 -2020 1112 -1954
rect 1156 -2020 1220 -1954
rect 1264 -2020 1328 -1954
rect 2056 -2018 2120 -1952
rect 2164 -2018 2228 -1952
rect 2272 -2018 2336 -1952
rect 2380 -2018 2444 -1952
rect 2488 -2018 2552 -1952
rect 2596 -2018 2660 -1952
rect 2704 -2018 2768 -1952
rect 2812 -2018 2876 -1952
rect 2920 -2018 2984 -1952
rect 3028 -2018 3092 -1952
rect 3092 -2018 3096 -1952
rect 3136 -2018 3200 -1952
rect 3200 -2018 3204 -1952
rect 3244 -2018 3308 -1952
rect 3308 -2018 3312 -1952
rect 3356 -2018 3420 -1952
rect 3464 -2018 3528 -1952
rect 3572 -2018 3636 -1952
<< metal2 >>
rect -348 424 1276 464
rect -348 358 -322 424
rect -258 358 -214 424
rect -150 358 -106 424
rect -42 358 2 424
rect 66 358 110 424
rect 174 358 218 424
rect 282 358 326 424
rect 390 358 434 424
rect 498 358 542 424
rect 606 358 650 424
rect 718 358 758 424
rect 826 358 866 424
rect 934 358 978 424
rect 1042 358 1086 424
rect 1150 358 1194 424
rect 1258 358 1276 424
rect -348 336 1276 358
rect 2028 424 3652 464
rect 2028 358 2054 424
rect 2118 358 2162 424
rect 2226 358 2270 424
rect 2334 358 2378 424
rect 2442 358 2486 424
rect 2550 358 2594 424
rect 2658 358 2702 424
rect 2766 358 2810 424
rect 2874 358 2918 424
rect 2982 358 3026 424
rect 3094 358 3134 424
rect 3202 358 3242 424
rect 3310 358 3354 424
rect 3418 358 3462 424
rect 3526 358 3570 424
rect 3634 358 3652 424
rect 2028 336 3652 358
rect 1138 100 1324 112
rect 1138 36 1150 100
rect 1214 36 1246 100
rect 1310 36 1324 100
rect 1138 26 1324 36
rect 2198 100 2384 112
rect 2198 36 2208 100
rect 2272 36 2304 100
rect 2368 36 2384 100
rect 2198 26 2384 36
rect 1392 -922 1478 -912
rect 1392 -986 1402 -922
rect 1466 -986 1478 -922
rect 1392 -1018 1478 -986
rect 1392 -1082 1402 -1018
rect 1466 -1082 1478 -1018
rect 1392 -1094 1478 -1082
rect 2016 -922 2102 -912
rect 2016 -986 2026 -922
rect 2090 -986 2102 -922
rect 2016 -1018 2102 -986
rect 2016 -1082 2026 -1018
rect 2090 -1082 2102 -1018
rect 2016 -1094 2102 -1082
rect -278 -1954 1346 -1914
rect -278 -2020 -252 -1954
rect -188 -2020 -144 -1954
rect -80 -2020 -36 -1954
rect 28 -2020 72 -1954
rect 136 -2020 180 -1954
rect 244 -2020 288 -1954
rect 352 -2020 396 -1954
rect 460 -2020 504 -1954
rect 568 -2020 612 -1954
rect 676 -2020 720 -1954
rect 788 -2020 828 -1954
rect 896 -2020 936 -1954
rect 1004 -2020 1048 -1954
rect 1112 -2020 1156 -1954
rect 1220 -2020 1264 -1954
rect 1328 -2020 1346 -1954
rect -278 -2042 1346 -2020
rect 2030 -1952 3654 -1912
rect 2030 -2018 2056 -1952
rect 2120 -2018 2164 -1952
rect 2228 -2018 2272 -1952
rect 2336 -2018 2380 -1952
rect 2444 -2018 2488 -1952
rect 2552 -2018 2596 -1952
rect 2660 -2018 2704 -1952
rect 2768 -2018 2812 -1952
rect 2876 -2018 2920 -1952
rect 2984 -2018 3028 -1952
rect 3096 -2018 3136 -1952
rect 3204 -2018 3244 -1952
rect 3312 -2018 3356 -1952
rect 3420 -2018 3464 -1952
rect 3528 -2018 3572 -1952
rect 3636 -2018 3654 -1952
rect 2030 -2040 3654 -2018
<< via2 >>
rect -322 358 -258 424
rect -214 358 -150 424
rect -106 358 -42 424
rect 2 358 66 424
rect 110 358 174 424
rect 218 358 282 424
rect 326 358 390 424
rect 434 358 498 424
rect 542 358 606 424
rect 650 358 718 424
rect 758 358 826 424
rect 866 358 934 424
rect 978 358 1042 424
rect 1086 358 1150 424
rect 1194 358 1258 424
rect 2054 358 2118 424
rect 2162 358 2226 424
rect 2270 358 2334 424
rect 2378 358 2442 424
rect 2486 358 2550 424
rect 2594 358 2658 424
rect 2702 358 2766 424
rect 2810 358 2874 424
rect 2918 358 2982 424
rect 3026 358 3094 424
rect 3134 358 3202 424
rect 3242 358 3310 424
rect 3354 358 3418 424
rect 3462 358 3526 424
rect 3570 358 3634 424
rect 1150 36 1214 100
rect 1246 36 1310 100
rect 2208 36 2272 100
rect 2304 36 2368 100
rect 1402 -986 1466 -922
rect 1402 -1082 1466 -1018
rect 2026 -986 2090 -922
rect 2026 -1082 2090 -1018
rect -252 -2020 -188 -1954
rect -144 -2020 -80 -1954
rect -36 -2020 28 -1954
rect 72 -2020 136 -1954
rect 180 -2020 244 -1954
rect 288 -2020 352 -1954
rect 396 -2020 460 -1954
rect 504 -2020 568 -1954
rect 612 -2020 676 -1954
rect 720 -2020 788 -1954
rect 828 -2020 896 -1954
rect 936 -2020 1004 -1954
rect 1048 -2020 1112 -1954
rect 1156 -2020 1220 -1954
rect 1264 -2020 1328 -1954
rect 2056 -2018 2120 -1952
rect 2164 -2018 2228 -1952
rect 2272 -2018 2336 -1952
rect 2380 -2018 2444 -1952
rect 2488 -2018 2552 -1952
rect 2596 -2018 2660 -1952
rect 2704 -2018 2768 -1952
rect 2812 -2018 2876 -1952
rect 2920 -2018 2984 -1952
rect 3028 -2018 3096 -1952
rect 3136 -2018 3204 -1952
rect 3244 -2018 3312 -1952
rect 3356 -2018 3420 -1952
rect 3464 -2018 3528 -1952
rect 3572 -2018 3636 -1952
<< metal3 >>
rect -279 3464 1620 4364
rect 1704 3464 3603 4364
rect 566 3364 672 3464
rect 2652 3364 2758 3464
rect -279 2464 1620 3364
rect 1704 2464 3603 3364
rect 568 2364 674 2464
rect 2650 2364 2756 2464
rect -279 1464 1620 2364
rect 1704 1464 3603 2364
rect 566 1364 672 1464
rect 2652 1364 2758 1464
rect -279 464 1620 1364
rect 1704 464 3603 1364
rect -348 424 1276 464
rect -348 358 -322 424
rect -258 358 -214 424
rect -150 358 -106 424
rect -42 358 2 424
rect 66 358 110 424
rect 174 358 218 424
rect 282 358 326 424
rect 390 358 434 424
rect 498 358 542 424
rect 606 358 650 424
rect 718 358 758 424
rect 826 358 866 424
rect 934 358 978 424
rect 1042 358 1086 424
rect 1150 358 1194 424
rect 1258 358 1276 424
rect -348 334 1276 358
rect 2028 424 3652 464
rect 2028 358 2054 424
rect 2118 358 2162 424
rect 2226 358 2270 424
rect 2334 358 2378 424
rect 2442 358 2486 424
rect 2550 358 2594 424
rect 2658 358 2702 424
rect 2766 358 2810 424
rect 2874 358 2918 424
rect 2982 358 3026 424
rect 3094 358 3134 424
rect 3202 358 3242 424
rect 3310 358 3354 424
rect 3418 358 3462 424
rect 3526 358 3570 424
rect 3634 358 3652 424
rect 2028 334 3652 358
rect 1138 100 1324 112
rect 1138 36 1150 100
rect 1310 36 1324 100
rect 1138 26 1324 36
rect 2198 100 2384 112
rect 2198 36 2208 100
rect 2368 36 2384 100
rect 2198 26 2384 36
rect 1392 -922 1478 -912
rect 1392 -986 1402 -922
rect 1466 -986 1478 -922
rect 1392 -1018 1478 -986
rect 1392 -1082 1402 -1018
rect 1466 -1082 1478 -1018
rect 1392 -1094 1478 -1082
rect 2016 -922 2102 -912
rect 2016 -986 2026 -922
rect 2090 -986 2102 -922
rect 2016 -1018 2102 -986
rect 2016 -1082 2026 -1018
rect 2090 -1082 2102 -1018
rect 2016 -1094 2102 -1082
rect -278 -1954 1346 -1914
rect -278 -2020 -252 -1954
rect -188 -2020 -144 -1954
rect -80 -2020 -36 -1954
rect 28 -2020 72 -1954
rect 136 -2020 180 -1954
rect 244 -2020 288 -1954
rect 352 -2020 396 -1954
rect 460 -2020 504 -1954
rect 568 -2020 612 -1954
rect 676 -2020 720 -1954
rect 788 -2020 828 -1954
rect 896 -2020 936 -1954
rect 1004 -2020 1048 -1954
rect 1112 -2020 1156 -1954
rect 1220 -2020 1264 -1954
rect 1328 -2020 1346 -1954
rect -278 -2042 1346 -2020
rect 2030 -1952 3654 -1912
rect 2030 -2018 2056 -1952
rect 2120 -2018 2164 -1952
rect 2228 -2018 2272 -1952
rect 2336 -2018 2380 -1952
rect 2444 -2018 2488 -1952
rect 2552 -2018 2596 -1952
rect 2660 -2018 2704 -1952
rect 2768 -2018 2812 -1952
rect 2876 -2018 2920 -1952
rect 2984 -2018 3028 -1952
rect 3096 -2018 3136 -1952
rect 3204 -2018 3244 -1952
rect 3312 -2018 3356 -1952
rect 3420 -2018 3464 -1952
rect 3528 -2018 3572 -1952
rect 3636 -2018 3654 -1952
rect 2030 -2040 3654 -2018
rect 2029 -2042 3654 -2040
rect -279 -2942 1620 -2042
rect 1704 -2942 3603 -2042
rect 566 -3042 672 -2942
rect 2652 -3042 2758 -2942
rect -279 -3942 1620 -3042
rect 1704 -3942 3603 -3042
rect 568 -4042 674 -3942
rect 2650 -4042 2756 -3942
rect -279 -4942 1620 -4042
rect 1704 -4942 3603 -4042
rect 566 -5042 672 -4942
rect 2652 -5042 2758 -4942
rect -279 -5942 1620 -5042
rect 1704 -5942 3603 -5042
<< via3 >>
rect 1150 36 1214 100
rect 1214 36 1246 100
rect 1246 36 1310 100
rect 2208 36 2272 100
rect 2272 36 2304 100
rect 2304 36 2368 100
rect 1402 -986 1466 -922
rect 1402 -1082 1466 -1018
rect 2026 -986 2090 -922
rect 2026 -1082 2090 -1018
<< mimcap >>
rect -179 4224 1421 4264
rect -179 3604 -139 4224
rect 1381 3604 1421 4224
rect -179 3564 1421 3604
rect 1903 4224 3503 4264
rect 1903 3604 1943 4224
rect 3463 3604 3503 4224
rect 1903 3564 3503 3604
rect -179 3224 1421 3264
rect -179 2604 -139 3224
rect 1381 2604 1421 3224
rect -179 2564 1421 2604
rect 1903 3224 3503 3264
rect 1903 2604 1943 3224
rect 3463 2604 3503 3224
rect 1903 2564 3503 2604
rect -179 2224 1421 2264
rect -179 1604 -139 2224
rect 1381 1604 1421 2224
rect -179 1564 1421 1604
rect 1903 2224 3503 2264
rect 1903 1604 1943 2224
rect 3463 1604 3503 2224
rect 1903 1564 3503 1604
rect -179 1224 1421 1264
rect -179 604 -139 1224
rect 1381 604 1421 1224
rect -179 564 1421 604
rect 1903 1224 3503 1264
rect 1903 604 1943 1224
rect 3463 604 3503 1224
rect 1903 564 3503 604
rect -179 -2182 1421 -2142
rect -179 -2802 -139 -2182
rect 1381 -2802 1421 -2182
rect -179 -2842 1421 -2802
rect 1903 -2182 3503 -2142
rect 1903 -2802 1943 -2182
rect 3463 -2802 3503 -2182
rect 1903 -2842 3503 -2802
rect -179 -3182 1421 -3142
rect -179 -3802 -139 -3182
rect 1381 -3802 1421 -3182
rect -179 -3842 1421 -3802
rect 1903 -3182 3503 -3142
rect 1903 -3802 1943 -3182
rect 3463 -3802 3503 -3182
rect 1903 -3842 3503 -3802
rect -179 -4182 1421 -4142
rect -179 -4802 -139 -4182
rect 1381 -4802 1421 -4182
rect -179 -4842 1421 -4802
rect 1903 -4182 3503 -4142
rect 1903 -4802 1943 -4182
rect 3463 -4802 3503 -4182
rect 1903 -4842 3503 -4802
rect -179 -5182 1421 -5142
rect -179 -5802 -139 -5182
rect 1381 -5802 1421 -5182
rect -179 -5842 1421 -5802
rect 1903 -5182 3503 -5142
rect 1903 -5802 1943 -5182
rect 3463 -5802 3503 -5182
rect 1903 -5842 3503 -5802
<< mimcapcontact >>
rect -139 3604 1381 4224
rect 1943 3604 3463 4224
rect -139 2604 1381 3224
rect 1943 2604 3463 3224
rect -139 1604 1381 2224
rect 1943 1604 3463 2224
rect -139 604 1381 1224
rect 1943 604 3463 1224
rect -139 -2802 1381 -2182
rect 1943 -2802 3463 -2182
rect -139 -3802 1381 -3182
rect 1943 -3802 3463 -3182
rect -139 -4802 1381 -4182
rect 1943 -4802 3463 -4182
rect -139 -5802 1381 -5182
rect 1943 -5802 3463 -5182
<< metal4 >>
rect 569 4225 673 4414
rect 2651 4225 2755 4414
rect -140 4224 1382 4225
rect -140 3604 -139 4224
rect 1381 3604 1382 4224
rect -140 3603 1382 3604
rect 1942 4224 3464 4225
rect 1942 3604 1943 4224
rect 3463 3604 3464 4224
rect 1942 3603 3464 3604
rect 569 3225 673 3603
rect 2651 3225 2755 3603
rect -140 3224 1382 3225
rect -140 2604 -139 3224
rect 1381 2604 1382 3224
rect -140 2603 1382 2604
rect 1942 3224 3464 3225
rect 1942 2604 1943 3224
rect 3463 2604 3464 3224
rect 1942 2603 3464 2604
rect 569 2225 673 2603
rect 2651 2225 2755 2603
rect -140 2224 1382 2225
rect -140 1604 -139 2224
rect 1381 1604 1382 2224
rect -140 1603 1382 1604
rect 1942 2224 3464 2225
rect 1942 1604 1943 2224
rect 3463 1604 3464 2224
rect 1942 1603 3464 1604
rect 569 1225 673 1603
rect 2651 1225 2755 1603
rect -140 1224 1382 1225
rect -140 604 -139 1224
rect 1381 604 1382 1224
rect -140 603 1382 604
rect 1942 1224 3464 1225
rect 1942 604 1943 1224
rect 3463 604 3464 1224
rect 1942 603 3464 604
rect 569 464 673 603
rect 2651 466 2755 603
rect 568 336 1324 464
rect 1138 100 1324 336
rect 1138 36 1150 100
rect 1310 36 1324 100
rect 1138 24 1324 36
rect 2198 414 2755 466
rect 2198 334 2754 414
rect 2198 100 2384 334
rect 2198 36 2208 100
rect 2368 36 2384 100
rect 2198 26 2384 36
rect 1392 -922 1478 -912
rect 1392 -986 1402 -922
rect 1466 -986 1478 -922
rect 1392 -1018 1478 -986
rect 1392 -1082 1402 -1018
rect 1466 -1082 1478 -1018
rect 1392 -1810 1478 -1082
rect 568 -1894 1478 -1810
rect 2016 -922 2102 -912
rect 2016 -986 2026 -922
rect 2090 -986 2102 -922
rect 2016 -1018 2102 -986
rect 2016 -1082 2026 -1018
rect 2090 -1082 2102 -1018
rect 2016 -1810 2102 -1082
rect 2016 -1894 2756 -1810
rect 568 -2008 674 -1894
rect 568 -2010 673 -2008
rect 569 -2181 673 -2010
rect 2650 -2181 2756 -1894
rect -140 -2182 1382 -2181
rect -140 -2802 -139 -2182
rect 1381 -2802 1382 -2182
rect -140 -2803 1382 -2802
rect 1942 -2182 3464 -2181
rect 1942 -2802 1943 -2182
rect 3463 -2802 3464 -2182
rect 1942 -2803 3464 -2802
rect 569 -3181 673 -2803
rect 2651 -3181 2755 -2803
rect -140 -3182 1382 -3181
rect -140 -3802 -139 -3182
rect 1381 -3802 1382 -3182
rect -140 -3803 1382 -3802
rect 1942 -3182 3464 -3181
rect 1942 -3802 1943 -3182
rect 3463 -3802 3464 -3182
rect 1942 -3803 3464 -3802
rect 569 -4181 673 -3803
rect 2651 -4181 2755 -3803
rect -140 -4182 1382 -4181
rect -140 -4802 -139 -4182
rect 1381 -4802 1382 -4182
rect -140 -4803 1382 -4802
rect 1942 -4182 3464 -4181
rect 1942 -4802 1943 -4182
rect 3463 -4802 3464 -4182
rect 1942 -4803 3464 -4802
rect 569 -5181 673 -4803
rect 2651 -5181 2755 -4803
rect -140 -5182 1382 -5181
rect -140 -5802 -139 -5182
rect 1381 -5802 1382 -5182
rect -140 -5803 1382 -5802
rect 1942 -5182 3464 -5181
rect 1942 -5802 1943 -5182
rect 3463 -5802 3464 -5182
rect 1942 -5803 3464 -5802
rect 569 -5992 673 -5803
rect 2651 -5992 2755 -5803
<< comment >>
rect -2 -58 30 -16
rect 194 -62 226 -20
rect 384 -64 416 -22
rect 576 -64 608 -22
rect 768 -62 800 -20
rect 1332 -350 1350 -146
rect 1554 -338 1574 -118
rect 1748 -366 1768 -146
rect 1942 -308 1962 -88
rect 2168 -350 2186 -146
rect 4 -752 36 -710
rect 192 -738 224 -696
rect 380 -736 412 -694
rect 584 -732 616 -690
rect 772 -724 804 -682
rect 1548 -1056 1576 -888
rect 1742 -1058 1770 -890
rect 1934 -1072 1962 -904
rect 96 -1140 128 -1098
rect 294 -1142 326 -1100
rect 482 -1140 514 -1098
rect 670 -1140 702 -1098
use adc_comp_buffer  adc_comp_buffer_0 ../adc_comp_buffer
timestamp 1661416858
transform 1 0 2600 0 1 -226
box -42 -326 408 452
use adc_comp_buffer  adc_comp_buffer_1
timestamp 1661416858
transform 1 0 2600 0 1 -1038
box -42 -326 408 452
<< labels >>
rlabel metal1 -714 -352 -714 -324 7 inn
port 6 w
rlabel metal1 -714 -272 -714 -244 7 inp
port 5 w
rlabel metal1 -714 162 -714 300 7 VDD
port 1 w
rlabel metal1 -714 -1484 -714 -1326 7 VSS
port 2 w
rlabel metal1 -716 -1706 -716 -1660 7 clk
port 3 w
rlabel metal1 -122 -1558 -122 -1512 7 op
rlabel metal1 784 -1632 784 -1586 7 on
rlabel locali 1210 -602 1210 -568 7 bn
rlabel locali 2300 -602 2300 -568 3 bp
rlabel metal1 3920 -276 3920 -230 3 outp
port 7 e
rlabel metal1 3920 -1088 3920 -1042 3 outn
port 8 e
rlabel metal1 -716 -1780 -716 -1734 7 nclk
port 4 w
<< end >>
