magic
tech sky130A
magscale 1 2
timestamp 1671363782
<< nwell >>
rect 111 880 1004 1004
rect 0 506 1004 880
rect 141 499 859 506
<< nmos >>
rect 227 51 271 431
rect 329 51 373 431
rect 431 51 475 431
rect 533 51 577 431
rect 635 51 679 431
rect 737 51 781 431
<< pmos >>
rect 223 588 267 968
rect 325 588 369 968
rect 427 588 471 968
rect 529 588 573 968
rect 631 588 675 968
rect 733 588 777 968
<< ndiff >>
rect 169 419 227 431
rect 169 100 181 419
rect 215 100 227 419
rect 169 51 227 100
rect 271 338 329 431
rect 271 63 283 338
rect 317 63 329 338
rect 271 51 329 63
rect 373 419 431 431
rect 373 63 385 419
rect 419 63 431 419
rect 373 51 431 63
rect 475 345 533 431
rect 475 63 487 345
rect 521 63 533 345
rect 475 51 533 63
rect 577 419 635 431
rect 577 63 589 419
rect 623 63 635 419
rect 577 51 635 63
rect 679 419 737 431
rect 679 63 691 419
rect 725 63 737 419
rect 679 51 737 63
rect 781 419 840 431
rect 781 103 793 419
rect 827 103 840 419
rect 781 51 840 103
<< pdiff >>
rect 170 928 223 968
rect 170 600 178 928
rect 212 600 223 928
rect 170 588 223 600
rect 267 956 325 968
rect 267 600 279 956
rect 313 600 325 956
rect 267 588 325 600
rect 369 956 427 968
rect 369 600 381 956
rect 415 600 427 956
rect 369 588 427 600
rect 471 956 529 968
rect 471 677 483 956
rect 517 677 529 956
rect 471 588 529 677
rect 573 956 631 968
rect 573 600 585 956
rect 619 600 631 956
rect 573 588 631 600
rect 675 956 733 968
rect 675 677 687 956
rect 721 677 733 956
rect 675 588 733 677
rect 777 930 835 968
rect 777 600 789 930
rect 823 600 835 930
rect 777 588 835 600
<< ndiffc >>
rect 181 100 215 419
rect 283 63 317 338
rect 385 63 419 419
rect 487 63 521 345
rect 589 63 623 419
rect 691 63 725 419
rect 793 103 827 419
<< pdiffc >>
rect 178 600 212 928
rect 279 600 313 956
rect 381 600 415 956
rect 483 677 517 956
rect 585 600 619 956
rect 687 677 721 956
rect 789 600 823 930
<< psubdiff >>
rect 895 192 970 216
rect 895 136 903 192
rect 963 136 970 192
rect 895 112 970 136
<< nsubdiff >>
rect 898 832 967 876
rect 898 776 907 832
rect 958 776 967 832
rect 898 720 967 776
<< psubdiffcont >>
rect 903 136 963 192
<< nsubdiffcont >>
rect 907 776 958 832
<< poly >>
rect 223 968 267 994
rect 325 968 369 994
rect 427 968 471 994
rect 529 968 573 994
rect 631 968 675 994
rect 733 968 777 994
rect 223 572 267 588
rect 325 572 369 588
rect 223 538 369 572
rect 223 486 269 538
rect 334 486 369 538
rect 427 573 471 588
rect 529 573 573 588
rect 631 573 675 588
rect 733 573 777 588
rect 427 569 777 573
rect 427 530 781 569
rect 427 518 668 530
rect 223 476 369 486
rect 635 478 668 518
rect 733 478 781 530
rect 223 450 577 476
rect 227 446 577 450
rect 227 431 271 446
rect 329 431 373 446
rect 431 431 475 446
rect 533 431 577 446
rect 635 446 781 478
rect 635 431 679 446
rect 737 431 781 446
rect 227 25 271 51
rect 329 25 373 51
rect 431 25 475 51
rect 533 25 577 51
rect 635 25 679 51
rect 737 25 781 51
<< polycont >>
rect 269 486 334 538
rect 668 478 733 530
<< locali >>
rect 34 970 148 1004
rect 34 924 142 970
rect 279 956 313 972
rect 34 888 46 924
rect 136 888 142 924
rect 34 102 142 888
rect 178 928 212 953
rect 212 600 279 627
rect 381 956 415 972
rect 313 600 381 627
rect 483 956 517 972
rect 483 661 517 677
rect 585 956 619 972
rect 415 600 585 627
rect 687 956 721 972
rect 856 970 970 1004
rect 687 661 721 677
rect 789 930 823 946
rect 619 600 789 627
rect 857 924 970 970
rect 857 888 868 924
rect 958 888 970 924
rect 857 882 970 888
rect 907 847 958 848
rect 907 760 958 776
rect 178 584 823 600
rect 857 667 970 715
rect 857 631 879 667
rect 958 631 970 667
rect 252 486 269 538
rect 334 486 350 538
rect 457 525 541 584
rect 857 531 970 631
rect 457 485 477 525
rect 523 485 541 525
rect 457 437 541 485
rect 652 525 668 530
rect 652 488 665 525
rect 652 478 668 488
rect 733 478 749 530
rect 34 66 46 102
rect 136 66 142 102
rect 177 419 827 437
rect 177 100 181 419
rect 215 396 385 419
rect 177 76 215 100
rect 283 338 317 362
rect 34 34 142 66
rect 283 47 317 56
rect 419 395 589 419
rect 385 47 419 63
rect 487 345 521 361
rect 487 47 521 56
rect 623 395 691 419
rect 589 47 623 63
rect 725 395 793 419
rect 792 103 793 395
rect 862 332 970 531
rect 862 292 878 332
rect 958 292 970 332
rect 862 230 970 292
rect 887 136 903 192
rect 963 136 979 192
rect 792 86 827 103
rect 691 47 725 63
rect 34 0 148 34
rect 854 0 970 51
<< viali >>
rect 46 888 136 924
rect 483 889 517 927
rect 687 888 721 926
rect 868 888 958 924
rect 907 832 958 847
rect 907 804 958 832
rect 879 631 958 667
rect 269 487 334 524
rect 477 485 523 525
rect 665 488 668 525
rect 668 488 708 525
rect 46 66 136 102
rect 283 63 317 98
rect 283 56 317 63
rect 487 63 521 98
rect 487 56 521 63
rect 878 292 958 332
rect 903 143 963 185
<< metal1 >>
rect 34 924 148 1004
rect 856 963 970 1004
rect 34 888 46 924
rect 136 888 148 924
rect 34 882 148 888
rect 266 882 272 934
rect 324 927 733 934
rect 324 889 483 927
rect 517 926 733 927
rect 517 889 687 926
rect 324 888 687 889
rect 721 888 733 926
rect 324 882 733 888
rect 856 924 879 963
rect 856 888 868 924
rect 961 888 970 963
rect 856 882 970 888
rect 0 847 1004 854
rect 0 804 907 847
rect 958 804 1004 847
rect 0 798 1004 804
rect 0 740 1004 770
rect 865 707 970 712
rect 48 673 837 701
rect 48 596 77 673
rect 0 568 77 596
rect 808 596 837 673
rect 865 632 876 707
rect 865 631 879 632
rect 958 631 970 707
rect 865 625 970 631
rect 105 559 780 588
rect 808 568 1004 596
rect 105 540 134 559
rect 0 512 134 540
rect 751 540 780 559
rect 257 524 352 531
rect 257 487 269 524
rect 334 487 352 524
rect 257 479 352 487
rect 404 479 410 531
rect 465 479 474 531
rect 526 479 535 531
rect 653 479 665 531
rect 717 479 723 531
rect 751 512 1004 540
rect 0 451 128 458
rect 748 451 1004 458
rect 0 430 1004 451
rect 99 423 776 430
rect 0 374 71 402
rect 42 342 71 374
rect 804 374 1004 402
rect 804 342 833 374
rect 42 314 833 342
rect 866 286 872 338
rect 964 286 970 338
rect 0 220 1004 258
rect 0 185 1004 192
rect 0 143 903 185
rect 963 143 1004 185
rect 0 136 1004 143
rect 34 102 148 108
rect 34 66 46 102
rect 136 66 148 102
rect 34 0 148 66
rect 258 56 272 108
rect 324 104 330 108
rect 854 107 970 108
rect 324 98 533 104
rect 324 56 487 98
rect 521 56 533 98
rect 258 47 533 56
rect 854 55 866 107
rect 958 55 970 107
rect 277 0 317 47
rect 854 0 970 55
<< via1 >>
rect 272 882 324 934
rect 879 924 961 963
rect 879 888 958 924
rect 958 888 961 924
rect 876 667 958 707
rect 876 632 879 667
rect 879 632 958 667
rect 352 479 404 531
rect 474 525 526 531
rect 474 485 477 525
rect 477 485 523 525
rect 523 485 526 525
rect 474 479 526 485
rect 665 525 717 531
rect 665 488 708 525
rect 708 488 717 525
rect 665 479 717 488
rect 872 332 964 338
rect 872 292 878 332
rect 878 292 958 332
rect 958 292 964 332
rect 872 286 964 292
rect 272 98 324 108
rect 272 56 283 98
rect 283 56 317 98
rect 317 56 324 98
rect 866 55 958 107
<< metal2 >>
rect 32 962 244 972
rect 32 906 42 962
rect 98 906 138 962
rect 194 906 244 962
rect 352 962 832 972
rect 32 866 244 906
rect 32 810 42 866
rect 98 810 244 866
rect 32 770 244 810
rect 32 714 42 770
rect 98 714 244 770
rect 32 674 244 714
rect 32 618 42 674
rect 98 618 138 674
rect 194 618 244 674
rect 32 578 244 618
rect 32 522 42 578
rect 98 522 244 578
rect 32 482 244 522
rect 32 426 42 482
rect 98 426 244 482
rect 32 386 244 426
rect 32 330 42 386
rect 98 330 138 386
rect 194 330 244 386
rect 32 290 244 330
rect 32 234 42 290
rect 98 234 244 290
rect 32 194 244 234
rect 32 138 42 194
rect 98 138 244 194
rect 32 98 244 138
rect 32 42 42 98
rect 98 42 138 98
rect 194 42 244 98
rect 272 934 324 940
rect 272 108 324 882
rect 352 906 426 962
rect 482 906 522 962
rect 578 906 618 962
rect 674 906 714 962
rect 770 906 832 962
rect 352 866 832 906
rect 352 810 618 866
rect 674 810 832 866
rect 352 578 832 810
rect 463 540 538 549
rect 272 50 324 56
rect 352 531 404 537
rect 352 472 404 479
rect 463 476 470 540
rect 534 476 538 540
rect 32 32 244 42
rect 352 0 391 472
rect 463 467 538 476
rect 567 431 628 578
rect 656 531 765 536
rect 656 479 665 531
rect 717 479 765 531
rect 656 472 765 479
rect 434 49 698 431
rect 726 0 765 472
rect 803 513 832 578
rect 865 963 972 972
rect 865 888 879 963
rect 961 888 972 963
rect 865 707 972 888
rect 865 632 876 707
rect 958 632 972 707
rect 865 552 972 632
rect 803 512 833 513
rect 803 482 972 512
rect 803 426 906 482
rect 962 426 972 482
rect 803 416 972 426
rect 861 338 972 359
rect 861 286 872 338
rect 964 286 972 338
rect 861 107 972 286
rect 861 55 866 107
rect 958 55 972 107
rect 861 32 972 55
<< via2 >>
rect 42 906 98 962
rect 138 906 194 962
rect 42 810 98 866
rect 42 714 98 770
rect 42 618 98 674
rect 138 618 194 674
rect 42 522 98 578
rect 42 426 98 482
rect 42 330 98 386
rect 138 330 194 386
rect 42 234 98 290
rect 42 138 98 194
rect 42 42 98 98
rect 138 42 194 98
rect 426 906 482 962
rect 522 906 578 962
rect 618 906 674 962
rect 714 906 770 962
rect 618 810 674 866
rect 470 531 534 540
rect 470 479 474 531
rect 474 479 526 531
rect 526 479 534 531
rect 470 476 534 479
rect 906 426 962 482
<< metal3 >>
rect 36 962 968 968
rect 36 906 42 962
rect 98 906 138 962
rect 194 906 426 962
rect 482 906 522 962
rect 578 906 618 962
rect 674 906 714 962
rect 770 906 968 962
rect 36 900 968 906
rect 36 866 104 900
rect 36 810 42 866
rect 98 810 104 866
rect 36 770 104 810
rect 36 714 42 770
rect 98 714 104 770
rect 164 824 264 840
rect 164 756 180 824
rect 248 756 264 824
rect 164 740 264 756
rect 36 680 104 714
rect 324 680 392 900
rect 36 674 392 680
rect 36 618 42 674
rect 98 618 138 674
rect 194 618 392 674
rect 36 612 392 618
rect 612 866 680 900
rect 612 810 618 866
rect 674 810 680 866
rect 612 680 680 810
rect 740 824 840 840
rect 740 756 756 824
rect 824 756 840 824
rect 740 740 840 756
rect 900 680 968 900
rect 612 612 968 680
rect 36 578 104 612
rect 36 522 42 578
rect 98 522 104 578
rect 36 482 104 522
rect 36 426 42 482
rect 98 426 104 482
rect 164 536 264 552
rect 164 468 180 536
rect 248 468 264 536
rect 164 452 264 468
rect 459 540 541 572
rect 459 476 470 540
rect 534 476 541 540
rect 459 450 541 476
rect 740 536 840 552
rect 740 468 756 536
rect 824 468 840 536
rect 740 452 840 468
rect 900 482 968 612
rect 36 392 104 426
rect 900 426 906 482
rect 962 426 968 482
rect 900 392 968 426
rect 36 386 324 392
rect 36 330 42 386
rect 98 330 138 386
rect 194 330 324 386
rect 36 324 324 330
rect 681 324 968 392
rect 36 290 104 324
rect 36 234 42 290
rect 98 234 104 290
rect 36 194 104 234
rect 36 138 42 194
rect 98 138 104 194
rect 164 248 264 264
rect 164 180 180 248
rect 248 180 264 248
rect 164 164 264 180
rect 740 248 840 264
rect 740 180 756 248
rect 824 180 840 248
rect 740 164 840 180
rect 36 104 104 138
rect 900 104 968 324
rect 36 98 324 104
rect 36 42 42 98
rect 98 42 138 98
rect 194 42 324 98
rect 36 36 324 42
rect 692 36 968 104
<< via3 >>
rect 180 756 248 824
rect 756 756 824 824
rect 180 468 248 536
rect 470 476 534 540
rect 756 468 824 536
rect 180 180 248 248
rect 756 180 824 248
<< metal4 >>
rect 184 840 244 934
rect 164 824 264 840
rect 164 820 180 824
rect 70 760 180 820
rect 164 756 180 760
rect 248 820 264 824
rect 248 760 360 820
rect 248 756 264 760
rect 164 740 264 756
rect 184 552 244 740
rect 164 536 264 552
rect 472 542 532 934
rect 760 840 820 934
rect 740 824 840 840
rect 740 820 756 824
rect 646 760 756 820
rect 740 756 756 760
rect 824 820 840 824
rect 824 760 934 820
rect 824 756 840 760
rect 740 740 840 756
rect 760 552 820 740
rect 164 532 180 536
rect 70 472 180 532
rect 164 468 180 472
rect 248 468 264 536
rect 468 540 536 542
rect 468 476 470 540
rect 534 476 536 540
rect 468 473 536 476
rect 740 536 840 552
rect 164 452 264 468
rect 184 264 244 452
rect 164 248 264 264
rect 164 244 180 248
rect 70 184 180 244
rect 164 180 180 184
rect 248 180 264 248
rect 164 164 264 180
rect 184 70 244 164
rect 472 48 532 473
rect 740 468 756 536
rect 824 532 840 536
rect 824 472 934 532
rect 824 468 840 472
rect 740 452 840 468
rect 760 264 820 452
rect 740 248 840 264
rect 740 180 756 248
rect 824 244 840 248
rect 824 184 934 244
rect 824 180 840 184
rect 740 164 840 180
rect 760 70 820 164
<< comment >>
rect 0 972 32 1004
rect 972 972 1004 1004
rect 0 0 32 32
rect 972 0 1004 32
<< labels >>
rlabel metal1 0 740 0 770 7 sample_n
port 2 w
rlabel metal1 0 512 0 540 7 rowon_n
port 3 w
rlabel metal1 0 430 0 458 7 row_n
port 4 w
rlabel metal1 0 220 0 248 7 vcom
port 6 w
rlabel metal1 0 136 0 192 7 VSS
port 7 w
rlabel locali 854 0 970 0 5 col_n
port 8 s
rlabel metal1 0 798 0 854 7 VDD
port 13 w
rlabel space 0 366 0 394 7 sample
port 5 w
flabel metal1 277 0 317 22 0 FreeSans 64 0 0 0 analog_in
port 16 nsew
flabel metal2 726 0 765 23 0 FreeSans 80 0 0 0 sw_n
port 19 nsew
flabel metal2 352 0 391 23 0 FreeSans 80 0 0 0 sw
port 17 nsew
<< end >>
