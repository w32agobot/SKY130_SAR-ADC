magic
tech sky130A
magscale 1 2
timestamp 1679566582
<< nwell >>
rect 0 464 1004 880
<< nmos >>
rect 321 236 351 356
rect 519 236 549 356
rect 717 236 747 356
<< pmos >>
rect 321 502 351 742
rect 519 502 549 742
rect 717 502 747 742
<< ndiff >>
rect 264 348 321 356
rect 264 244 276 348
rect 310 244 321 348
rect 264 236 321 244
rect 351 282 408 356
rect 351 244 362 282
rect 396 244 408 282
rect 351 236 408 244
rect 462 348 519 356
rect 462 244 474 348
rect 508 244 519 348
rect 462 236 519 244
rect 549 282 606 356
rect 549 244 560 282
rect 594 244 606 282
rect 549 236 606 244
rect 660 348 717 356
rect 660 244 672 348
rect 706 244 717 348
rect 660 236 717 244
rect 747 282 804 356
rect 747 244 758 282
rect 792 244 804 282
rect 747 236 804 244
<< pdiff >>
rect 264 734 321 742
rect 264 518 276 734
rect 310 518 321 734
rect 264 502 321 518
rect 351 734 408 742
rect 351 586 362 734
rect 396 586 408 734
rect 351 502 408 586
rect 462 734 519 742
rect 462 518 474 734
rect 508 518 519 734
rect 462 502 519 518
rect 549 734 606 742
rect 549 586 560 734
rect 594 586 606 734
rect 549 502 606 586
rect 660 734 717 742
rect 660 518 672 734
rect 706 518 717 734
rect 660 502 717 518
rect 747 734 804 742
rect 747 586 758 734
rect 792 586 804 734
rect 747 502 804 586
<< ndiffc >>
rect 276 244 310 348
rect 362 244 396 282
rect 474 244 508 348
rect 560 244 594 282
rect 672 244 706 348
rect 758 244 792 282
<< pdiffc >>
rect 276 518 310 734
rect 362 586 396 734
rect 474 518 508 734
rect 560 586 594 734
rect 672 518 706 734
rect 758 586 792 734
<< psubdiff >>
rect 182 148 230 182
rect 264 148 326 182
rect 360 148 430 182
rect 464 148 534 182
rect 568 148 628 182
rect 662 148 726 182
rect 760 148 792 182
<< nsubdiff >>
rect 198 838 806 844
rect 198 804 222 838
rect 256 804 326 838
rect 360 804 430 838
rect 464 804 534 838
rect 568 804 630 838
rect 664 804 724 838
rect 758 804 806 838
rect 198 798 806 804
<< psubdiffcont >>
rect 230 148 264 182
rect 326 148 360 182
rect 430 148 464 182
rect 534 148 568 182
rect 628 148 662 182
rect 726 148 760 182
<< nsubdiffcont >>
rect 222 804 256 838
rect 326 804 360 838
rect 430 804 464 838
rect 534 804 568 838
rect 630 804 664 838
rect 724 804 758 838
<< poly >>
rect 321 742 351 770
rect 519 742 549 770
rect 717 742 747 770
rect 321 466 351 502
rect 519 466 549 502
rect 717 466 747 502
rect 277 450 351 466
rect 277 416 287 450
rect 321 416 351 450
rect 277 400 351 416
rect 475 450 549 466
rect 475 416 485 450
rect 519 416 549 450
rect 475 400 549 416
rect 673 450 747 466
rect 673 416 683 450
rect 717 416 747 450
rect 673 400 747 416
rect 321 356 351 400
rect 519 356 549 400
rect 717 356 747 400
rect 321 210 351 236
rect 519 210 549 236
rect 717 210 747 236
<< polycont >>
rect 287 416 321 450
rect 485 416 519 450
rect 683 416 717 450
<< locali >>
rect 34 922 182 1004
rect 34 888 48 922
rect 136 888 182 922
rect 34 882 182 888
rect 910 922 970 1004
rect 910 888 922 922
rect 956 888 970 922
rect 910 882 970 888
rect 34 706 148 882
rect 182 838 820 844
rect 182 804 222 838
rect 256 804 326 838
rect 360 804 430 838
rect 464 804 534 838
rect 568 804 630 838
rect 664 804 724 838
rect 758 804 820 838
rect 182 798 820 804
rect 34 630 48 706
rect 130 630 148 706
rect 34 340 148 630
rect 276 734 310 750
rect 362 734 396 798
rect 362 570 396 586
rect 474 734 508 750
rect 310 518 389 536
rect 276 502 389 518
rect 560 734 594 798
rect 642 734 706 750
rect 642 733 672 734
rect 642 692 656 733
rect 642 672 672 692
rect 560 570 594 586
rect 508 518 587 536
rect 474 502 587 518
rect 758 734 792 798
rect 758 570 792 586
rect 706 518 785 536
rect 672 502 785 518
rect 355 466 389 502
rect 553 466 587 502
rect 186 450 321 466
rect 186 416 287 450
rect 186 400 321 416
rect 355 450 519 466
rect 355 416 485 450
rect 355 400 519 416
rect 553 450 717 466
rect 553 416 683 450
rect 553 400 717 416
rect 186 396 232 400
rect 186 362 192 396
rect 226 362 232 396
rect 355 366 389 400
rect 553 396 638 400
rect 553 366 585 396
rect 186 350 232 362
rect 34 292 48 340
rect 132 292 148 340
rect 34 106 148 292
rect 276 348 389 366
rect 310 332 389 348
rect 474 362 585 366
rect 619 362 638 396
rect 751 366 785 502
rect 474 348 638 362
rect 276 228 310 244
rect 362 282 396 298
rect 362 182 396 244
rect 508 332 638 348
rect 672 348 785 366
rect 474 228 508 244
rect 560 282 594 298
rect 560 182 594 244
rect 706 332 785 348
rect 854 340 970 882
rect 672 228 706 244
rect 758 282 792 298
rect 758 182 792 244
rect 182 148 230 182
rect 264 148 326 182
rect 360 148 430 182
rect 464 148 534 182
rect 568 148 628 182
rect 662 148 726 182
rect 760 148 792 182
rect 854 292 868 340
rect 956 292 970 340
rect 854 108 970 292
rect 34 102 182 106
rect 34 68 46 102
rect 136 68 182 102
rect 34 0 182 68
rect 910 102 970 108
rect 910 68 922 102
rect 958 68 970 102
rect 910 0 970 68
<< viali >>
rect 48 888 136 922
rect 922 888 956 922
rect 222 804 256 838
rect 326 804 360 838
rect 430 804 464 838
rect 534 804 568 838
rect 630 804 664 838
rect 724 804 758 838
rect 48 630 130 706
rect 656 692 672 733
rect 672 692 693 733
rect 192 362 226 396
rect 48 292 132 340
rect 585 362 619 396
rect 230 148 264 182
rect 326 148 360 182
rect 430 148 464 182
rect 534 148 568 182
rect 628 148 662 182
rect 726 148 760 182
rect 868 292 956 340
rect 46 68 136 102
rect 922 68 958 102
<< metal1 >>
rect 34 922 182 1004
rect 34 888 48 922
rect 136 888 182 922
rect 34 882 182 888
rect 910 922 970 1004
rect 910 888 922 922
rect 956 888 970 922
rect 910 882 970 888
rect 0 838 1004 854
rect 0 804 222 838
rect 256 804 326 838
rect 360 804 430 838
rect 464 804 534 838
rect 568 804 630 838
rect 664 804 724 838
rect 758 804 1004 838
rect 0 798 1004 804
rect 0 740 158 770
rect 642 740 1004 770
rect 642 738 816 740
rect 642 733 706 738
rect 34 706 142 712
rect 34 630 48 706
rect 130 630 142 706
rect 642 692 656 733
rect 693 692 706 733
rect 642 672 706 692
rect 34 624 142 630
rect 0 568 1004 596
rect 0 512 1004 540
rect 0 430 1004 458
rect 0 396 238 402
rect 0 374 192 396
rect 180 362 192 374
rect 226 362 238 396
rect 180 356 238 362
rect 573 396 1004 402
rect 573 362 585 396
rect 619 374 1004 396
rect 619 362 631 374
rect 573 356 631 362
rect 34 340 144 346
rect 34 292 48 340
rect 132 292 144 340
rect 34 286 144 292
rect 854 340 970 346
rect 854 292 868 340
rect 956 292 970 340
rect 854 286 970 292
rect 0 220 1004 258
rect 0 182 1004 192
rect 0 148 230 182
rect 264 148 326 182
rect 360 148 430 182
rect 464 148 534 182
rect 568 148 628 182
rect 662 148 726 182
rect 760 148 1004 182
rect 0 136 1004 148
rect 34 102 182 108
rect 34 68 46 102
rect 136 68 182 102
rect 34 0 182 68
rect 910 102 970 108
rect 910 68 922 102
rect 958 68 970 102
rect 910 0 970 68
<< metal2 >>
rect 32 962 972 972
rect 32 906 42 962
rect 98 906 138 962
rect 194 906 234 962
rect 290 906 330 962
rect 386 906 426 962
rect 482 906 522 962
rect 578 906 618 962
rect 674 906 714 962
rect 770 906 810 962
rect 866 906 906 962
rect 962 906 972 962
rect 32 866 972 906
rect 32 810 42 866
rect 98 810 330 866
rect 386 810 618 866
rect 674 810 906 866
rect 962 810 972 866
rect 32 770 972 810
rect 32 714 42 770
rect 98 714 330 770
rect 386 714 618 770
rect 674 714 906 770
rect 962 714 972 770
rect 32 674 972 714
rect 32 618 42 674
rect 98 618 138 674
rect 194 618 234 674
rect 290 618 330 674
rect 386 618 426 674
rect 482 618 522 674
rect 578 618 618 674
rect 674 618 714 674
rect 770 618 810 674
rect 866 618 906 674
rect 962 618 972 674
rect 32 608 972 618
rect 32 578 396 608
rect 32 522 42 578
rect 98 522 330 578
rect 386 522 396 578
rect 608 578 972 608
rect 32 482 396 522
rect 32 426 42 482
rect 98 426 330 482
rect 386 426 396 482
rect 460 460 544 544
rect 608 522 618 578
rect 674 522 906 578
rect 962 522 972 578
rect 608 482 972 522
rect 32 396 396 426
rect 608 426 618 482
rect 674 426 906 482
rect 962 426 972 482
rect 608 396 972 426
rect 32 386 972 396
rect 32 330 42 386
rect 98 330 138 386
rect 194 330 234 386
rect 290 330 330 386
rect 386 330 426 386
rect 482 330 522 386
rect 578 330 618 386
rect 674 330 714 386
rect 770 330 810 386
rect 866 330 906 386
rect 962 330 972 386
rect 32 290 972 330
rect 32 234 42 290
rect 98 234 330 290
rect 386 234 618 290
rect 674 234 906 290
rect 962 234 972 290
rect 32 194 972 234
rect 32 138 42 194
rect 98 138 330 194
rect 386 138 618 194
rect 674 138 906 194
rect 962 138 972 194
rect 32 98 972 138
rect 32 42 42 98
rect 98 42 138 98
rect 194 42 234 98
rect 290 42 330 98
rect 386 42 426 98
rect 482 42 522 98
rect 578 42 618 98
rect 674 42 714 98
rect 770 42 810 98
rect 866 42 906 98
rect 962 42 972 98
rect 32 32 972 42
<< via2 >>
rect 42 906 98 962
rect 138 906 194 962
rect 234 906 290 962
rect 330 906 386 962
rect 426 906 482 962
rect 522 906 578 962
rect 618 906 674 962
rect 714 906 770 962
rect 810 906 866 962
rect 906 906 962 962
rect 42 810 98 866
rect 330 810 386 866
rect 618 810 674 866
rect 906 810 962 866
rect 42 714 98 770
rect 330 714 386 770
rect 618 714 674 770
rect 906 714 962 770
rect 42 618 98 674
rect 138 618 194 674
rect 234 618 290 674
rect 330 618 386 674
rect 426 618 482 674
rect 522 618 578 674
rect 618 618 674 674
rect 714 618 770 674
rect 810 618 866 674
rect 906 618 962 674
rect 42 522 98 578
rect 330 522 386 578
rect 42 426 98 482
rect 330 426 386 482
rect 618 522 674 578
rect 906 522 962 578
rect 618 426 674 482
rect 906 426 962 482
rect 42 330 98 386
rect 138 330 194 386
rect 234 330 290 386
rect 330 330 386 386
rect 426 330 482 386
rect 522 330 578 386
rect 618 330 674 386
rect 714 330 770 386
rect 810 330 866 386
rect 906 330 962 386
rect 42 234 98 290
rect 330 234 386 290
rect 618 234 674 290
rect 906 234 962 290
rect 42 138 98 194
rect 330 138 386 194
rect 618 138 674 194
rect 906 138 962 194
rect 42 42 98 98
rect 138 42 194 98
rect 234 42 290 98
rect 330 42 386 98
rect 426 42 482 98
rect 522 42 578 98
rect 618 42 674 98
rect 714 42 770 98
rect 810 42 866 98
rect 906 42 962 98
<< metal3 >>
rect 36 962 968 968
rect 36 906 42 962
rect 98 906 138 962
rect 194 906 234 962
rect 290 906 330 962
rect 386 906 426 962
rect 482 906 522 962
rect 578 906 618 962
rect 674 906 714 962
rect 770 906 810 962
rect 866 906 906 962
rect 962 906 968 962
rect 36 900 968 906
rect 36 866 104 900
rect 36 810 42 866
rect 98 810 104 866
rect 324 866 392 900
rect 36 770 104 810
rect 36 714 42 770
rect 98 714 104 770
rect 164 824 264 840
rect 164 756 180 824
rect 248 756 264 824
rect 164 740 264 756
rect 324 810 330 866
rect 386 810 392 866
rect 612 866 680 900
rect 324 770 392 810
rect 36 680 104 714
rect 324 714 330 770
rect 386 714 392 770
rect 452 824 552 840
rect 452 756 468 824
rect 536 756 552 824
rect 452 740 552 756
rect 612 810 618 866
rect 674 810 680 866
rect 900 866 968 900
rect 612 770 680 810
rect 324 680 392 714
rect 612 714 618 770
rect 674 714 680 770
rect 740 824 840 840
rect 740 756 756 824
rect 824 756 840 824
rect 740 740 840 756
rect 900 810 906 866
rect 962 810 968 866
rect 900 770 968 810
rect 612 680 680 714
rect 900 714 906 770
rect 962 714 968 770
rect 900 680 968 714
rect 36 674 968 680
rect 36 618 42 674
rect 98 618 138 674
rect 194 618 234 674
rect 290 618 330 674
rect 386 618 426 674
rect 482 618 522 674
rect 578 618 618 674
rect 674 618 714 674
rect 770 618 810 674
rect 866 618 906 674
rect 962 618 968 674
rect 36 612 968 618
rect 36 578 104 612
rect 36 522 42 578
rect 98 522 104 578
rect 324 578 392 612
rect 36 482 104 522
rect 36 426 42 482
rect 98 426 104 482
rect 164 536 264 552
rect 164 468 180 536
rect 248 468 264 536
rect 164 452 264 468
rect 324 522 330 578
rect 386 522 392 578
rect 324 482 392 522
rect 36 392 104 426
rect 324 426 330 482
rect 386 426 392 482
rect 324 392 392 426
rect 612 578 680 612
rect 612 522 618 578
rect 674 522 680 578
rect 900 578 968 612
rect 612 482 680 522
rect 612 426 618 482
rect 674 426 680 482
rect 740 536 840 552
rect 740 468 756 536
rect 824 468 840 536
rect 740 452 840 468
rect 900 522 906 578
rect 962 522 968 578
rect 900 482 968 522
rect 612 392 680 426
rect 900 426 906 482
rect 962 426 968 482
rect 900 392 968 426
rect 36 386 968 392
rect 36 330 42 386
rect 98 330 138 386
rect 194 330 234 386
rect 290 330 330 386
rect 386 330 426 386
rect 482 330 522 386
rect 578 330 618 386
rect 674 330 714 386
rect 770 330 810 386
rect 866 330 906 386
rect 962 330 968 386
rect 36 324 968 330
rect 36 290 104 324
rect 36 234 42 290
rect 98 234 104 290
rect 324 290 392 324
rect 36 194 104 234
rect 36 138 42 194
rect 98 138 104 194
rect 164 248 264 264
rect 164 180 180 248
rect 248 180 264 248
rect 164 164 264 180
rect 324 234 330 290
rect 386 234 392 290
rect 612 290 680 324
rect 324 194 392 234
rect 36 104 104 138
rect 324 138 330 194
rect 386 138 392 194
rect 452 248 552 264
rect 452 180 468 248
rect 536 180 552 248
rect 452 164 552 180
rect 612 234 618 290
rect 674 234 680 290
rect 900 290 968 324
rect 612 194 680 234
rect 324 104 392 138
rect 612 138 618 194
rect 674 138 680 194
rect 740 248 840 264
rect 740 180 756 248
rect 824 180 840 248
rect 740 164 840 180
rect 900 234 906 290
rect 962 234 968 290
rect 900 194 968 234
rect 612 104 680 138
rect 900 138 906 194
rect 962 138 968 194
rect 900 104 968 138
rect 36 98 968 104
rect 36 42 42 98
rect 98 42 138 98
rect 194 42 234 98
rect 290 42 330 98
rect 386 42 426 98
rect 482 42 522 98
rect 578 42 618 98
rect 674 42 714 98
rect 770 42 810 98
rect 866 42 906 98
rect 962 42 968 98
rect 36 36 968 42
<< via3 >>
rect 180 756 248 824
rect 468 756 536 824
rect 756 756 824 824
rect 180 468 248 536
rect 756 468 824 536
rect 180 180 248 248
rect 468 180 536 248
rect 756 180 824 248
<< metal4 >>
rect 184 840 244 934
rect 472 840 532 934
rect 760 840 820 934
rect 164 824 264 840
rect 164 820 180 824
rect 70 760 180 820
rect 164 756 180 760
rect 248 820 264 824
rect 452 824 552 840
rect 452 820 468 824
rect 248 760 468 820
rect 248 756 264 760
rect 164 740 264 756
rect 452 756 468 760
rect 536 820 552 824
rect 740 824 840 840
rect 740 820 756 824
rect 536 760 756 820
rect 536 756 552 760
rect 452 740 552 756
rect 740 756 756 760
rect 824 820 840 824
rect 824 760 934 820
rect 824 756 840 760
rect 740 740 840 756
rect 184 552 244 740
rect 472 646 532 740
rect 760 552 820 740
rect 164 536 264 552
rect 164 532 180 536
rect 70 472 180 532
rect 164 468 180 472
rect 248 532 264 536
rect 740 536 840 552
rect 740 532 756 536
rect 248 472 358 532
rect 646 472 756 532
rect 248 468 264 472
rect 164 452 264 468
rect 740 468 756 472
rect 824 532 840 536
rect 824 472 934 532
rect 824 468 840 472
rect 740 452 840 468
rect 184 264 244 452
rect 472 264 532 358
rect 760 264 820 452
rect 164 248 264 264
rect 164 244 180 248
rect 70 184 180 244
rect 164 180 180 184
rect 248 244 264 248
rect 452 248 552 264
rect 452 244 468 248
rect 248 184 468 244
rect 248 180 264 184
rect 164 164 264 180
rect 452 180 468 184
rect 536 244 552 248
rect 740 248 840 264
rect 740 244 756 248
rect 536 184 756 244
rect 536 180 552 184
rect 452 164 552 180
rect 740 180 756 184
rect 824 244 840 248
rect 824 184 934 244
rect 824 180 840 184
rect 740 164 840 180
rect 184 70 244 164
rect 472 70 532 164
rect 760 70 820 164
<< comment >>
rect 0 972 32 1004
rect 972 972 1004 1004
rect 138 750 308 798
rect 430 756 562 804
rect 138 260 194 750
rect 312 690 368 750
rect 358 428 406 688
rect 430 562 478 756
rect 564 716 606 762
rect 598 608 632 716
rect 576 604 632 608
rect 558 602 632 604
rect 558 576 608 602
rect 544 562 600 576
rect 430 558 600 562
rect 430 544 576 558
rect 430 514 558 544
rect 430 460 478 514
rect 560 478 602 522
rect 560 476 636 478
rect 428 428 478 460
rect 358 396 428 428
rect 300 260 356 318
rect 358 314 406 396
rect 138 258 356 260
rect 138 212 306 258
rect 430 206 478 428
rect 602 198 636 476
rect 670 198 716 802
rect 0 0 32 32
rect 972 0 1004 32
<< labels >>
flabel metal1 837 798 1004 854 0 FreeSans 160 0 0 0 VDD
port 1 e power bidirectional
flabel metal1 0 136 1004 192 0 FreeSans 320 0 0 0 VSS
port 2 nsew ground bidirectional
flabel metal4 472 874 532 934 1 FreeSans 160 0 0 0 ctop
port 4 n
flabel metal1 34 0 182 108 5 FreeSans 320 0 0 0 col
port 5 s
flabel metal1 34 882 182 1004 1 FreeSans 320 0 0 0 col
port 5 n
flabel space 910 882 970 1004 1 FreeSans 320 0 0 0 col_n
port 6 n
flabel metal1 846 430 1004 458 0 FreeSans 160 0 0 0 row_n
port 7 e
flabel metal1 0 512 155 540 0 FreeSans 160 0 0 0 rowon_n
port 8 w
flabel metal1 849 512 1004 540 0 FreeSans 160 0 0 0 rowon_n
port 8 e
flabel metal1 846 374 1004 402 0 FreeSans 160 0 0 0 sample_o
port 10 e
flabel metal1 846 740 1004 770 0 FreeSans 160 0 0 0 sample_n_o
port 12 nsew
flabel metal1 0 568 156 596 7 FreeSans 160 0 0 0 off_n
port 13 w
flabel metal1 848 568 1004 596 3 FreeSans 160 0 0 0 off_n
port 13 e
rlabel metal2 500 972 500 972 1 cbot
flabel space 910 0 970 108 1 FreeSans 320 0 0 0 col_n
port 6 s
flabel metal1 0 798 167 854 0 FreeSans 160 0 0 0 VDD
port 1 w power bidirectional
flabel metal1 0 740 158 770 0 FreeSans 160 0 0 0 sample_n_i
port 11 nsew
flabel metal1 0 374 158 402 0 FreeSans 160 0 0 0 sample_i
port 9 w
flabel metal1 0 430 158 458 0 FreeSans 160 0 0 0 row_n
port 7 w
flabel metal1 0 220 1004 258 0 FreeSans 320 0 0 0 vcom
port 3 nsew
<< end >>
