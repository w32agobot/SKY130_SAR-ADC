* NGSPICE file created from adc_array_matrix_12bit.ext - technology: sky130A

.subckt adc_array_matrix_12bit_ext VDD VSS vcm sample sample_n row_n[0] row_n[1] row_n[2] row_n[3]
+ row_n[4] row_n[5] row_n[6] row_n[7] row_n[8] row_n[9] row_n[10] row_n[11] row_n[12] row_n[13] row_n[14]
+ row_n[15] rowon_n[0] rowon_n[1] rowon_n[2] rowon_n[3] rowon_n[4] rowon_n[5] rowon_n[6] rowon_n[7] rowon_n[8]
+ rowon_n[9] rowon_n[10] rowon_n[11] rowon_n[12] rowon_n[13] rowon_n[14] rowon_n[15] col_n[0] col_n[1] col_n[2]
+ col_n[3] col_n[4] col_n[5] col_n[6] col_n[7] col_n[8] col_n[9] col_n[10] col_n[11] col_n[12] col_n[13]
+ col_n[14] col_n[15] col_n[16] col_n[17] col_n[18] col_n[19] col_n[20] col_n[21] col_n[22] col_n[23] col_n[24]
+ col_n[25] col_n[26] col_n[27] col_n[28] col_n[29] col_n[30] col_n[31] en_bit_n[0] en_bit_n[1] en_bit_n[2] en_C0_n sw sw_n analog_in ctop rowoff_n[0] rowoff_n[1] rowoff_n[2]
+ rowoff_n[3] rowoff_n[4] rowoff_n[5] rowoff_n[6] rowoff_n[7] rowoff_n[8] rowoff_n[9] rowoff_n[10] rowoff_n[11]
+ rowoff_n[12] rowoff_n[13] rowoff_n[14] rowoff_n[15] col[0] col[1] col[2] col[3] col[4] col[5] col[6] col[7] col[8] col[9]
+ col[10] col[11] col[12] col[13] col[14] col[15] col[16] col[17] col[18] col[19] col[20] col[21] col[22]
+ col[23] col[24] col[25] col[26] col[27] col[28] col[29] col[30] col[31] 
X0 a_3970_15182# a_2346_15224# a_3878_15182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1 a_3878_9158# a_1962_9198# a_3970_9158# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2 VDD rowon_n[5] a_18938_7150# VDD sky130_fd_pr__pfet_01v8 ad=1.74408e+14p pd=1.50002e+09u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3 a_30986_7150# row_n[5] a_31478_7512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4 vcm a_1962_18234# a_32082_18194# VSS sky130_fd_pr__nfet_01v8 ad=7.72086e+13p pd=8.6578e+08u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5 a_12002_2130# a_2346_2172# a_11910_2130# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6 a_5374_4500# col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7 a_14410_15544# col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8 a_10906_12170# row_n[10] a_11398_12532# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X9 a_35398_9198# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=4.35964e+14p ps=2.02062e+09u w=420000u l=150000u
X10 VSS sample a_2346_8196# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X11 a_17422_7512# col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X12 a_18026_7150# a_2346_7192# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=1.47064e+14p ps=1.31646e+09u w=800000u l=150000u
X13 VSS row_n[4] a_9294_6186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X14 a_4370_15544# col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15 a_23046_11166# a_2346_11208# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X16 a_22346_10202# rowon_n[8] a_21950_10162# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X17 a_14922_11166# row_n[9] a_15414_11528# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X18 a_15414_2492# col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X19 a_4882_11166# row_n[9] a_5374_11528# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X20 a_34394_2170# col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X21 a_27062_12170# a_2346_12212# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X22 VSS row_n[6] a_26362_8194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X23 a_34090_3134# a_2346_3176# a_33998_3134# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X24 a_26058_18194# a_2346_18236# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X25 a_21342_2170# rowon_n[0] a_20946_2130# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X26 a_35002_9158# row_n[7] a_35494_9520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X27 a_23350_18234# VDD a_22954_18194# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X28 VSS row_n[13] a_20338_15222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X29 a_26970_14178# a_1962_14218# a_27062_14178# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X30 a_11302_8194# rowon_n[6] a_10906_8154# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X31 a_29982_4138# a_1962_4178# a_30074_4138# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X32 a_12306_4178# rowon_n[2] a_11910_4138# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X33 vcm a_1962_2170# a_13006_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X34 VDD rowon_n[3] a_22954_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X35 VSS row_n[12] a_24354_14218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X36 a_21342_11206# col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X37 a_34394_10202# col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X38 a_24962_17190# a_1962_17230# a_25054_17190# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X39 VDD sample a_2346_15224# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X40 a_18938_7150# a_1962_7190# a_19030_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X41 a_4274_13214# rowon_n[11] a_3878_13174# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X42 a_14314_13214# rowon_n[11] a_13918_13174# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X43 VSS row_n[8] a_11302_10202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X44 a_20034_7150# a_2346_7192# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X45 a_21038_3134# a_2346_3176# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X46 a_19430_18556# col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X47 a_19030_14178# a_2346_14220# a_18938_14178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X48 VDD sample_n a_1962_11206# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X49 a_11910_11166# a_1962_11206# a_12002_11166# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X50 VDD rowon_n[14] a_22954_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X51 a_28978_14178# row_n[12] a_29470_14540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X52 a_20434_13536# col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X53 a_33486_12532# col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X54 vcm a_1962_10202# a_29070_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X55 a_20338_6186# col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X56 a_15926_12170# a_1962_12210# a_16018_12170# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X57 a_3270_7190# rowon_n[5] a_2874_7150# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X58 VSS row_n[4] a_30378_6186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X59 a_4274_3174# rowon_n[1] a_3878_3134# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X60 VDD rowon_n[2] a_11910_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X61 a_5886_12170# a_1962_12210# a_5978_12170# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X62 VDD rowon_n[10] a_9902_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X63 a_16322_6186# rowon_n[4] a_15926_6146# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X64 vcm a_1962_6186# a_24050_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X65 a_35398_18234# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X66 VDD rowon_n[9] a_3878_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X67 VDD rowon_n[9] a_13918_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X68 VDD rowon_n[4] a_5886_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X69 VSS VDD a_12306_18234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X70 a_30074_17190# a_2346_17232# a_29982_17190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X71 a_16018_7150# a_2346_7192# a_15926_7150# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X72 a_26058_1126# a_2346_1168# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X73 a_25054_5142# a_2346_5184# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X74 a_13310_14218# col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X75 VDD en_C0_n a_3878_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X76 a_30986_17190# row_n[15] a_31478_17552# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X77 a_12002_16186# a_2346_16228# a_11910_16186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X78 a_34090_16186# a_2346_16228# a_33998_16186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X79 a_3270_14218# col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X80 vcm a_1962_13214# a_31078_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X81 a_25358_4178# col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X82 a_35002_16186# row_n[14] a_35494_16548# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X83 a_10906_8154# row_n[6] a_11398_8516# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X84 VSS row_n[6] a_34394_8194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X85 a_8290_5182# rowon_n[3] a_7894_5142# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X86 a_9294_1166# VSS a_8898_1126# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X87 a_2346_3176# sample VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X88 VSS row_n[2] a_35398_4178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X89 a_9994_9158# a_2346_9200# a_9902_9158# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X90 a_12402_16548# col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X91 a_19334_16226# rowon_n[14] a_18938_16186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X92 a_20338_11206# rowon_n[9] a_19942_11166# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X93 vcm a_1962_8194# a_28066_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X94 vcm a_1962_4178# a_29070_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X95 a_1962_10202# sample_n VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X96 a_25358_7190# rowon_n[5] a_24962_7150# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X97 a_25054_13174# a_2346_13216# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X98 a_13310_7190# col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X99 a_29070_7150# a_2346_7192# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X100 a_14314_3174# col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X101 a_16018_12170# a_2346_12212# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X102 a_33998_9158# a_1962_9198# a_34090_9158# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X103 VDD rowon_n[1] a_7894_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X104 a_24962_4138# row_n[2] a_25454_4500# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X105 a_5978_12170# a_2346_12212# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X106 a_2874_7150# row_n[5] a_3366_7512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X107 vcm a_1962_7190# a_17022_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X108 a_35494_4500# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X109 a_19942_11166# a_1962_11206# a_20034_11166# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X110 a_32994_10162# a_1962_10202# a_33086_10162# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X111 a_15926_6146# row_n[4] a_16418_6508# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X112 a_34394_18234# VDD a_33998_18194# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X113 a_27366_17230# col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X114 VSS row_n[13] a_31382_15222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X115 a_13918_1126# VDD a_14410_1488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X116 VSS row_n[12] a_35398_14218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X117 a_32386_11206# col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X118 a_6282_2170# col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X119 a_22954_18194# a_1962_18234# a_23046_18194# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X120 a_12306_14218# rowon_n[12] a_11910_14178# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X121 a_18330_5182# col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X122 a_19334_1166# en_bit_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X123 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X124 VDD rowon_n[15] a_29982_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X125 a_26058_15182# a_2346_15224# a_25966_15182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X126 VSS en_bit_n[0] a_20338_1166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X127 vcm a_1962_11206# a_27062_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X128 a_7894_5142# row_n[3] a_8386_5504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X129 a_30378_1166# VSS a_29982_1126# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X130 VDD rowon_n[14] a_33998_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X131 a_26970_15182# row_n[13] a_27462_15544# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X132 a_31478_13536# col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X133 a_3878_13174# a_1962_13214# a_3970_13174# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X134 a_13918_13174# a_1962_13214# a_14010_13174# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X135 a_23046_5142# a_2346_5184# a_22954_5142# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X136 VDD rowon_n[6] a_30986_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X137 a_17934_3134# row_n[1] a_18426_3496# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X138 a_29374_9198# col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X139 a_29982_12170# row_n[10] a_30474_12532# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X140 VSS row_n[1] a_24354_3174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X141 a_10394_7512# col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X142 a_33390_7190# rowon_n[5] a_32994_7150# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X143 a_34394_3174# rowon_n[1] a_33998_3134# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X144 a_18330_11206# rowon_n[9] a_17934_11166# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X145 a_10998_7150# a_2346_7192# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X146 VSS row_n[7] a_14314_9198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X147 a_27062_7150# a_2346_7192# a_26970_7150# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X148 a_28066_3134# a_2346_3176# a_27974_3134# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X149 vcm a_1962_9198# a_32082_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X150 a_18938_18194# VDD a_19430_18556# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X151 vcm a_1962_14218# a_8990_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X152 vcm a_1962_14218# a_19030_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X153 a_4974_9158# a_2346_9200# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X154 a_28978_9158# row_n[7] a_29470_9520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X155 a_8898_18194# VDD a_9390_18556# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X156 a_22954_8154# a_1962_8194# a_23046_8154# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X157 a_24450_1488# col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X158 a_19030_2130# a_2346_2172# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X159 VSS row_n[0] a_13310_2170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X160 a_23958_4138# a_1962_4178# a_24050_4138# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X161 a_33086_8154# a_2346_8196# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X162 a_23046_14178# a_2346_14220# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X163 VSS VDD a_29374_1166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X164 a_14410_9520# col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X165 a_15414_5504# col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X166 VSS row_n[13] a_29374_15222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X167 a_33390_13214# rowon_n[11] a_32994_13174# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X168 a_26362_12210# col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X169 VSS row_n[8] a_30378_10202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X170 a_16018_5142# a_2346_5184# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X171 VSS row_n[2] a_7286_4178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X172 a_30986_11166# a_1962_11206# a_31078_11166# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X173 a_2346_9200# sample VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X174 a_11910_7150# a_1962_7190# a_12002_7150# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X175 VDD rowon_n[15] a_27974_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X176 a_25454_14540# col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X177 a_35002_12170# a_1962_12210# a_35094_12170# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X178 a_25054_10162# a_2346_10204# a_24962_10162# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X179 a_27974_6146# a_1962_6186# a_28066_6146# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X180 a_32082_1126# a_2346_1168# a_31990_1126# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X181 a_5886_9158# a_1962_9198# a_5978_9158# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X182 a_33998_18194# a_1962_18234# a_34090_18194# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X183 a_29470_13536# col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X184 VDD rowon_n[9] a_32994_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X185 a_25966_10162# row_n[8] a_26458_10524# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X186 a_32994_7150# row_n[5] a_33486_7512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X187 a_7382_4500# col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X188 a_14010_2130# a_2346_2172# a_13918_2130# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X189 a_30986_2130# row_n[0] a_31478_2492# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X190 VDD rowon_n[0] a_18938_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X191 a_11910_14178# a_1962_14218# a_12002_14178# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X192 VDD rowon_n[10] a_8898_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X193 VDD sample_n a_1962_14218# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X194 a_16930_5142# a_1962_5182# a_17022_5142# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X195 a_17422_2492# col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X196 vcm a_1962_15222# a_23046_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X197 VSS row_n[6] a_28370_8194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X198 a_17022_17190# a_2346_17232# a_16930_17190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X199 a_8290_15222# col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X200 a_18330_15222# col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X201 a_6982_17190# a_2346_17232# a_6890_17190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X202 a_9902_17190# a_1962_17230# a_9994_17190# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X203 a_23350_2170# rowon_n[0] a_22954_2130# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X204 vcm a_1962_10202# a_14010_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X205 a_2966_9158# a_2346_9200# a_2874_9158# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X206 a_7382_17552# col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X207 a_17422_17552# col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X208 a_3878_14178# row_n[12] a_4370_14540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X209 a_13918_14178# row_n[12] a_14410_14540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X210 a_25358_12210# rowon_n[10] a_24962_12170# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X211 vcm a_1962_10202# a_3970_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X212 a_13310_8194# rowon_n[6] a_12914_8154# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X213 vcm a_1962_8194# a_21038_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X214 vcm a_1962_4178# a_22042_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X215 a_14314_4178# rowon_n[2] a_13918_4138# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X216 a_2346_16228# sample VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X217 a_17934_13174# row_n[11] a_18426_13536# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X218 a_29374_11206# rowon_n[9] a_28978_11166# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X219 a_31078_8154# a_2346_8196# a_30986_8154# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X220 vcm a_1962_2170# a_15014_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X221 a_7894_13174# row_n[11] a_8386_13536# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X222 VDD rowon_n[6] a_2874_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X223 VDD sample a_2346_1168# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X224 a_23046_3134# a_2346_3176# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X225 a_22042_7150# a_2346_7192# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X226 VDD sample a_2346_10204# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X227 VDD rowon_n[8] a_24962_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X228 VDD rowon_n[2] a_13918_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X229 vcm a_1962_18234# a_4974_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X230 vcm a_1962_18234# a_15014_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X231 VSS row_n[15] a_23350_17230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X232 VSS row_n[4] a_32386_6186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X233 a_6282_3174# rowon_n[1] a_5886_3134# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X234 vcm a_1962_6186# a_26058_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X235 VSS row_n[14] a_27366_16226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X236 a_31382_14218# rowon_n[12] a_30986_14178# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X237 a_24354_13214# col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X238 vcm a_1962_9198# a_3970_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X239 VDD rowon_n[4] a_7894_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X240 a_32082_17190# a_2346_17232# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X241 a_17326_15222# rowon_n[13] a_16930_15182# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X242 a_11302_5182# col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X243 a_12306_1166# col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X244 a_28066_1126# a_2346_1168# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X245 a_7286_15222# rowon_n[13] a_6890_15182# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X246 a_19942_14178# a_1962_14218# a_20034_14178# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X247 a_32994_13174# a_1962_13214# a_33086_13174# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X248 a_18026_7150# a_2346_7192# a_17934_7150# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X249 a_27062_5142# a_2346_5184# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X250 VDD VDD a_25966_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X251 a_3970_16186# a_2346_16228# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X252 a_14010_16186# a_2346_16228# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X253 a_23446_15544# col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X254 VSS row_n[9] a_8290_11206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X255 VSS row_n[9] a_18330_11206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X256 a_23046_11166# a_2346_11208# a_22954_11166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X257 VDD VSS a_5886_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X258 a_23958_11166# row_n[9] a_24450_11528# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X259 a_12914_8154# row_n[6] a_13406_8516# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X260 VDD rowon_n[6] a_24962_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X261 VDD rowon_n[11] a_6890_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X262 VDD rowon_n[11] a_16930_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X263 a_10906_3134# row_n[1] a_11398_3496# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X264 a_12306_17230# col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X265 a_22346_9198# col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X266 a_27366_7190# rowon_n[5] a_26970_7150# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X267 a_16322_3174# col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X268 vcm a_1962_4178# a_30074_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X269 a_16322_16226# col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X270 vcm a_1962_16226# a_21038_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X271 a_15318_7190# col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X272 a_15014_18194# a_2346_18236# a_14922_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X273 a_6282_16226# col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X274 vcm a_1962_15222# a_34090_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X275 a_4882_7150# row_n[5] a_5374_7512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X276 a_4974_18194# a_2346_18236# a_4882_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X277 vcm a_1962_7190# a_19030_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X278 a_17934_6146# row_n[4] a_18426_6508# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X279 a_21038_3134# a_2346_3176# a_20946_3134# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X280 a_15414_18556# col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X281 a_11910_15182# row_n[13] a_12402_15544# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X282 vcm a_1962_11206# a_12002_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X283 a_20034_7150# a_2346_7192# a_19942_7150# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X284 a_2874_2130# row_n[0] a_3366_2492# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X285 a_5374_18556# col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X286 a_21950_9158# row_n[7] a_22442_9520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X287 a_15926_1126# VDD a_16418_1488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X288 a_8290_2170# col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X289 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.64e+07u l=1.6e+07u
X290 a_28066_15182# a_2346_15224# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X291 a_9902_2130# a_1962_2170# a_9994_2130# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X292 VSS row_n[10] a_22346_12210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X293 VSS VDD a_22346_1166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X294 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.64e+07u l=1.6e+07u
X295 a_32386_1166# VSS a_31990_1126# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X296 a_31382_5182# rowon_n[3] a_30986_5142# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X297 a_26058_1126# a_2346_1168# a_25966_1126# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X298 VSS VDD a_21342_18234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X299 a_25054_5142# a_2346_5184# a_24962_5142# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X300 VDD rowon_n[12] a_20946_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X301 a_22346_14218# col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X302 a_16322_10202# rowon_n[8] a_15926_10162# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X303 VDD rowon_n[6] a_32994_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X304 a_26970_7150# row_n[5] a_27462_7512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X305 a_6282_10202# rowon_n[8] a_5886_10162# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X306 a_30074_18194# a_2346_18236# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X307 a_22442_10524# col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X308 a_20946_6146# a_1962_6186# a_21038_6146# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X309 a_5278_16226# rowon_n[14] a_4882_16186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X310 a_15318_16226# rowon_n[14] a_14922_16186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X311 a_31078_6146# a_2346_6188# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X312 VDD rowon_n[1] a_30986_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X313 a_20338_17230# col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X314 a_21438_16548# col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X315 a_30986_14178# a_1962_14218# a_31078_14178# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X316 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.64e+07u l=1.6e+07u
X317 a_18330_9198# rowon_n[7] a_17934_9158# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X318 a_30378_9198# col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X319 a_12402_7512# col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X320 a_13006_7150# a_2346_7192# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X321 VSS row_n[4] a_4274_6186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X322 a_6890_15182# a_1962_15222# a_6982_15182# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X323 a_16930_15182# a_1962_15222# a_17022_15182# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X324 vcm a_1962_9198# a_34090_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X325 a_29070_7150# a_2346_7192# a_28978_7150# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X326 a_10394_2492# col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X327 VSS row_n[13] a_4274_15222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X328 VSS row_n[13] a_14314_15222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X329 a_11302_12210# col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X330 a_19942_15182# row_n[13] a_20434_15544# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X331 a_15318_11206# col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X332 vcm a_1962_11206# a_20034_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X333 a_6982_9158# a_2346_9200# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X334 VSS row_n[6] a_21342_8194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X335 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X336 a_32994_14178# row_n[12] a_33486_14540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X337 a_14010_13174# a_2346_13216# a_13918_13174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X338 a_5278_11206# col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X339 vcm a_1962_10202# a_33086_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X340 a_24962_8154# a_1962_8194# a_25054_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X341 VSS row_n[0] a_15318_2170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X342 a_25966_4138# a_1962_4178# a_26058_4138# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X343 a_3970_13174# a_2346_13216# a_3878_13174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X344 VDD rowon_n[7] a_17934_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X345 a_29982_9158# row_n[7] a_30474_9520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X346 a_35094_8154# a_2346_8196# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X347 VDD rowon_n[3] a_18938_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X348 a_30986_5142# row_n[3] a_31478_5504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X349 VDD rowon_n[15] a_2874_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X350 VDD rowon_n[15] a_12914_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X351 vcm a_1962_16226# a_32082_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X352 a_10394_14540# col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X353 a_5978_2130# a_2346_2172# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X354 a_14410_13536# col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X355 a_10906_10162# row_n[8] a_11398_10524# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X356 VSS sample a_2346_6188# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X357 a_17422_5504# col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X358 a_18026_5142# a_2346_5184# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X359 VSS row_n[2] a_9294_4178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X360 a_4370_13536# col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X361 a_13918_7150# a_1962_7190# a_14010_7150# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X362 VSS row_n[4] a_26362_6186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X363 a_26058_16186# a_2346_16228# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X364 a_7894_9158# a_1962_9198# a_7986_9158# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X365 a_35002_7150# row_n[5] a_35494_7512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X366 a_9390_4500# col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X367 VSS VDD a_19334_18234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X368 a_23350_16226# rowon_n[14] a_22954_16186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X369 VSS row_n[11] a_20338_13214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X370 a_11302_6186# rowon_n[4] a_10906_6146# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X371 VSS row_n[10] a_33390_12210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X372 a_32994_2130# row_n[0] a_33486_2492# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X373 a_6890_2130# a_1962_2170# a_6982_2130# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X374 a_10298_12210# rowon_n[10] a_9902_12170# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X375 a_24962_15182# a_1962_15222# a_25054_15182# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X376 VDD sample a_2346_13216# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X377 a_18938_5142# a_1962_5182# a_19030_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X378 a_28066_12170# a_2346_12212# a_27974_12170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X379 a_4274_11206# rowon_n[9] a_3878_11166# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X380 a_14314_11206# rowon_n[9] a_13918_11166# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X381 a_10998_7150# a_2346_7192# a_10906_7150# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X382 a_21038_1126# a_2346_1168# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X383 a_20034_5142# a_2346_5184# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X384 a_8990_17190# a_2346_17232# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X385 a_19430_16548# col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X386 VDD rowon_n[12] a_31990_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X387 a_28978_12170# row_n[10] a_29470_12532# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X388 a_20434_11528# col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X389 a_33486_10524# col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X390 a_20338_4178# col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X391 a_3270_5182# rowon_n[3] a_2874_5142# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X392 a_4274_1166# en_C0_n a_3878_1126# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X393 VSS row_n[2] a_30378_4178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X394 a_31382_17230# col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X395 VDD rowon_n[8] a_9902_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X396 a_4974_9158# a_2346_9200# a_4882_9158# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X397 a_19030_2130# a_2346_2172# a_18938_2130# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X398 a_16322_4178# rowon_n[2] a_15926_4138# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X399 vcm a_1962_8194# a_23046_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X400 vcm a_1962_4178# a_24050_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X401 a_35398_16226# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X402 a_33086_8154# a_2346_8196# a_32994_8154# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X403 VSS row_n[14] a_12306_16226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X404 a_20338_7190# rowon_n[5] a_19942_7150# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X405 vcm a_1962_17230# a_26058_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X406 a_30074_15182# a_2346_15224# a_29982_15182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X407 a_24050_7150# a_2346_7192# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X408 a_16018_5142# a_2346_5184# a_15926_5142# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X409 a_25054_3134# a_2346_3176# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X410 a_34090_14178# a_2346_14220# a_33998_14178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X411 VDD rowon_n[1] a_2874_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X412 a_19942_4138# row_n[2] a_20434_4500# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X413 a_34490_18556# col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X414 a_30986_15182# row_n[13] a_31478_15544# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X415 a_12002_14178# a_2346_14220# a_11910_14178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X416 vcm a_1962_11206# a_31078_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X417 vcm a_1962_7190# a_12002_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X418 a_1962_2170# sample_n VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X419 a_30474_4500# col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X420 VDD VDD a_10906_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X421 vcm a_1962_12210# a_17022_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X422 a_10906_6146# row_n[4] a_11398_6508# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X423 VSS row_n[4] a_34394_6186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X424 a_2346_1168# sample VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X425 a_8290_3174# rowon_n[1] a_7894_3134# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X426 VDD rowon_n[2] a_15926_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X427 vcm a_1962_12210# a_6982_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X428 a_19334_14218# rowon_n[12] a_18938_14178# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X429 vcm a_1962_6186# a_28066_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X430 vcm a_1962_9198# a_5978_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X431 a_21038_12170# a_2346_12212# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X432 a_25358_5182# rowon_n[3] a_24962_5142# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X433 a_13310_5182# col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X434 a_14314_1166# col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X435 a_29070_5142# a_2346_5184# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X436 VDD VSS a_7894_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X437 VDD rowon_n[6] a_26970_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X438 a_2874_5142# row_n[3] a_3366_5504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X439 vcm a_1962_5182# a_17022_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X440 a_30378_17230# rowon_n[15] a_29982_17190# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X441 a_14922_8154# row_n[6] a_15414_8516# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X442 a_3970_11166# a_2346_11208# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X443 a_14010_11166# a_2346_11208# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X444 a_34394_16226# rowon_n[14] a_33998_16186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X445 a_27366_15222# col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X446 VSS row_n[11] a_31382_13214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X447 VDD rowon_n[1] a_24962_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X448 a_12914_3134# row_n[1] a_13406_3496# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X449 a_24354_9198# col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X450 VSS row_n[5] a_19334_7190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X451 a_29374_7190# rowon_n[5] a_28978_7150# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X452 a_22954_16186# a_1962_16226# a_23046_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X453 a_18330_3174# col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X454 a_6982_18194# a_2346_18236# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X455 a_17022_18194# a_2346_18236# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X456 a_26458_17552# col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X457 VDD rowon_n[13] a_29982_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X458 a_26058_13174# a_2346_13216# a_25966_13174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X459 a_30378_12210# col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X460 a_26970_13174# row_n[11] a_27462_13536# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X461 a_31478_11528# col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X462 a_22042_7150# a_2346_7192# a_21950_7150# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X463 a_23046_3134# a_2346_3176# a_22954_3134# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X464 VDD rowon_n[4] a_30986_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X465 a_4882_2130# row_n[0] a_5374_2492# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X466 vcm a_1962_12210# a_25054_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X467 a_23958_9158# row_n[7] a_24450_9520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X468 a_17934_1126# en_bit_n[1] a_18426_1488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X469 a_19334_18234# col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X470 vcm a_1962_18234# a_24050_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X471 a_29982_10162# row_n[8] a_30474_10524# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X472 a_9294_18234# col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X473 VSS VDD a_24354_1166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X474 a_9390_14540# col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X475 a_10394_5504# col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X476 a_33390_5182# rowon_n[3] a_32994_5142# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X477 a_28066_10162# a_2346_10204# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X478 a_10998_5142# a_2346_5184# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X479 a_28066_1126# a_2346_1168# a_27974_1126# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X480 a_27062_5142# a_2346_5184# a_26970_5142# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X481 a_19030_12170# a_2346_12212# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X482 a_18938_16186# row_n[14] a_19430_16548# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X483 a_28978_7150# row_n[5] a_29470_7512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X484 a_8898_16186# row_n[14] a_9390_16548# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X485 a_22954_6146# a_1962_6186# a_23046_6146# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X486 a_33086_6146# a_2346_6188# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X487 a_26970_2130# row_n[0] a_27462_2492# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X488 VDD rowon_n[1] a_32994_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X489 a_28370_17230# rowon_n[15] a_27974_17190# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X490 a_14410_7512# col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X491 VSS sample a_2346_18236# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X492 VSS row_n[11] a_29374_13214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X493 a_33390_11206# rowon_n[9] a_32994_11166# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X494 a_26362_10202# col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X495 a_15014_7150# a_2346_7192# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X496 a_16018_3134# a_2346_3176# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X497 a_2346_7192# sample VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X498 a_11910_5142# a_1962_5182# a_12002_5142# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X499 a_12402_2492# col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X500 a_9294_12210# rowon_n[10] a_8898_12170# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X501 a_16930_10162# a_1962_10202# a_17022_10162# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X502 a_8990_9158# a_2346_9200# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X503 VSS row_n[6] a_23350_8194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X504 a_31382_2170# col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X505 a_19334_2170# rowon_n[0] a_18938_2130# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X506 VDD rowon_n[13] a_27974_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X507 a_25454_12532# col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X508 a_6890_10162# a_1962_10202# a_6982_10162# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X509 VSS row_n[0] a_17326_2170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X510 a_27974_4138# a_1962_4178# a_28066_4138# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X511 a_33998_16186# a_1962_16226# a_34090_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X512 a_29470_11528# col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X513 a_32994_5142# row_n[3] a_33486_5504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X514 a_7986_2130# a_2346_2172# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X515 VDD rowon_n[8] a_8898_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X516 vcm a_1962_2170# a_9994_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X517 VSS row_n[15] a_7286_17230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X518 VSS row_n[15] a_17326_17230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X519 a_22042_17190# a_2346_17232# a_21950_17190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X520 a_15926_7150# a_1962_7190# a_16018_7150# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X521 a_16930_3134# a_1962_3174# a_17022_3134# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X522 a_18330_13214# col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X523 vcm a_1962_13214# a_23046_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X524 VSS row_n[4] a_28370_6186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X525 a_22954_17190# row_n[15] a_23446_17552# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X526 a_17022_15182# a_2346_15224# a_16930_15182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X527 a_8290_13214# col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X528 VSS row_n[7] a_6282_9198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X529 a_6982_15182# a_2346_15224# a_6890_15182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X530 a_9902_15182# a_1962_15222# a_9994_15182# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X531 a_17422_15544# col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X532 a_7382_15544# col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X533 a_3878_12170# row_n[10] a_4370_12532# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X534 a_13918_12170# row_n[10] a_14410_12532# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X535 a_26058_11166# a_2346_11208# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X536 a_25358_10202# rowon_n[8] a_24962_10162# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X537 a_13310_6186# rowon_n[4] a_12914_6146# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X538 vcm a_1962_6186# a_21038_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X539 a_17934_11166# row_n[9] a_18426_11528# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X540 a_31078_6146# a_2346_6188# a_30986_6146# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X541 a_35002_2130# row_n[0] a_35494_2492# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X542 a_8898_2130# a_1962_2170# a_8990_2130# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X543 a_7894_11166# row_n[9] a_8386_11528# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X544 VDD rowon_n[4] a_2874_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X545 a_6378_9520# col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X546 a_23046_1126# a_2346_1168# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X547 a_13006_7150# a_2346_7192# a_12914_7150# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X548 a_22042_5142# a_2346_5184# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X549 vcm a_1962_17230# a_10998_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X550 a_24962_10162# a_1962_10202# a_25054_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X551 VDD rowon_n[6] a_19942_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X552 a_26362_18234# VDD a_25966_18194# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X553 vcm a_1962_16226# a_4974_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X554 vcm a_1962_16226# a_15014_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X555 VSS row_n[13] a_23350_15222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X556 a_6982_9158# a_2346_9200# a_6890_9158# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X557 a_6282_1166# VSS a_5886_1126# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X558 VSS row_n[2] a_32386_4178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X559 vcm a_1962_8194# a_25054_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X560 vcm a_1962_4178# a_26058_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X561 VSS row_n[12] a_27366_14218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X562 a_24354_11206# col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X563 a_35094_8154# a_2346_8196# a_35002_8154# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X564 a_27974_17190# a_1962_17230# a_28066_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X565 a_5978_2130# a_2346_2172# a_5886_2130# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X566 VDD rowon_n[15] a_21950_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X567 a_32082_15182# a_2346_15224# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X568 a_17326_13214# rowon_n[11] a_16930_13174# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X569 a_22346_7190# rowon_n[5] a_21950_7150# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X570 a_11302_3174# col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X571 a_7286_13214# rowon_n[11] a_6890_13174# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X572 a_30986_9158# a_1962_9198# a_31078_9158# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X573 a_10298_7190# col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X574 a_18026_5142# a_2346_5184# a_17934_5142# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X575 a_27062_3134# a_2346_3176# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X576 VDD rowon_n[14] a_25966_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X577 a_3970_14178# a_2346_14220# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X578 a_14010_14178# a_2346_14220# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X579 a_23446_13536# col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X580 a_32482_4500# col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X581 a_18938_12170# a_1962_12210# a_19030_12170# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X582 vcm a_1962_7190# a_14010_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X583 a_12914_6146# row_n[4] a_13406_6508# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X584 VDD rowon_n[4] a_24962_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X585 a_8898_12170# a_1962_12210# a_8990_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X586 VDD rowon_n[9] a_6890_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X587 VDD rowon_n[9] a_16930_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X588 a_10906_1126# VDD a_11398_1488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X589 VSS VDD a_15318_18234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X590 a_20034_18194# a_2346_18236# a_19942_18194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X591 a_12306_15222# col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X592 vcm a_1962_9198# a_7986_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X593 a_3270_2170# col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X594 VSS VDD a_5278_18234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X595 a_10998_17190# a_2346_17232# a_10906_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X596 a_33086_17190# a_2346_17232# a_32994_17190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X597 a_16322_1166# col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X598 a_27366_5182# rowon_n[3] a_26970_5142# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X599 a_20946_18194# VDD a_21438_18556# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X600 a_16322_14218# col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X601 vcm a_1962_14218# a_21038_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X602 a_5278_8194# rowon_n[6] a_4882_8154# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X603 a_15318_5182# col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X604 a_33998_17190# row_n[15] a_34490_17552# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X605 a_15014_16186# a_2346_16228# a_14922_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X606 a_6282_14218# col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X607 vcm a_1962_13214# a_34090_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X608 a_19430_8516# col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X609 a_4882_5142# row_n[3] a_5374_5504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X610 vcm a_1962_2170# a_6982_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X611 a_11398_17552# col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X612 a_4974_16186# a_2346_16228# a_4882_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X613 VDD rowon_n[6] a_28978_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X614 vcm a_1962_5182# a_19030_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X615 a_21038_1126# a_2346_1168# a_20946_1126# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X616 a_20034_5142# a_2346_5184# a_19942_5142# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X617 a_15414_16548# col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X618 a_11910_13174# row_n[11] a_12402_13536# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X619 VDD rowon_n[1] a_26970_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X620 a_5374_16548# col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X621 a_21950_7150# row_n[5] a_22442_7512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X622 a_14922_3134# row_n[1] a_15414_3496# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X623 a_28066_13174# a_2346_13216# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X624 vcm a_1962_12210# a_9994_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X625 a_26362_9198# col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X626 VSS row_n[8] a_22346_10202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X627 a_22954_11166# a_1962_11206# a_23046_11166# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X628 a_31382_3174# rowon_n[1] a_30986_3134# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X629 a_25054_3134# a_2346_3176# a_24962_3134# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X630 VSS row_n[14] a_21342_16226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X631 a_24050_7150# a_2346_7192# a_23958_7150# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X632 VDD rowon_n[10] a_20946_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X633 a_25966_9158# row_n[7] a_26458_9520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X634 VDD rowon_n[4] a_32994_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X635 a_26970_5142# row_n[3] a_27462_5504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X636 a_1962_9198# sample_n VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X637 a_25966_18194# a_1962_18234# a_26058_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X638 a_30074_16186# a_2346_16228# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X639 a_19942_8154# a_1962_8194# a_20034_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X640 VDD VSS a_30986_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X641 VSS row_n[0] a_10298_2170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X642 a_31078_4138# a_2346_4180# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X643 a_20946_4138# a_1962_4178# a_21038_4138# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X644 VDD VDD a_19942_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X645 a_5278_14218# rowon_n[12] a_4882_14178# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X646 a_15318_14218# rowon_n[12] a_14922_14178# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X647 a_30074_8154# a_2346_8196# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X648 a_20338_15222# col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X649 a_12402_5504# col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X650 a_13006_5142# a_2346_5184# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X651 VSS row_n[2] a_4274_4178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X652 a_13310_17230# rowon_n[15] a_12914_17190# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X653 a_6890_13174# a_1962_13214# a_6982_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X654 a_16930_13174# a_1962_13214# a_17022_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X655 a_7286_7190# col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X656 a_3270_17230# rowon_n[15] a_2874_17190# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X657 a_29070_5142# a_2346_5184# a_28978_5142# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X658 VSS row_n[11] a_4274_13214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X659 VSS row_n[11] a_14314_13214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X660 a_32082_12170# a_2346_12212# a_31990_12170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X661 a_11302_10202# col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X662 a_19942_13174# row_n[11] a_20434_13536# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X663 VSS row_n[4] a_21342_6186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X664 a_32994_12170# row_n[10] a_33486_12532# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X665 a_14010_11166# a_2346_11208# a_13918_11166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X666 a_24962_6146# a_1962_6186# a_25054_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X667 a_31078_18194# a_2346_18236# a_30986_18194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X668 a_3970_11166# a_2346_11208# a_3878_11166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X669 a_2874_9158# a_1962_9198# a_2966_9158# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X670 VDD rowon_n[5] a_17934_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X671 a_29982_7150# row_n[5] a_30474_7512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X672 a_35094_6146# a_2346_6188# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X673 a_28978_2130# row_n[0] a_29470_2492# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X674 a_31990_18194# VDD a_32482_18556# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X675 VDD rowon_n[13] a_2874_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X676 VDD rowon_n[13] a_12914_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X677 vcm a_1962_14218# a_32082_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X678 a_10394_12532# col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X679 a_4370_4500# col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X680 a_14410_11528# col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X681 a_18026_3134# a_2346_3176# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X682 a_4370_11528# col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X683 a_17022_7150# a_2346_7192# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X684 VDD sample_n a_1962_2170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X685 vcm a_1962_17230# a_30074_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X686 a_13918_5142# a_1962_5182# a_14010_5142# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X687 a_33390_2170# col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X688 a_14410_2492# col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X689 VSS row_n[6] a_25358_8194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X690 VSS row_n[2] a_26362_4178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X691 a_35398_8194# rowon_n[6] a_35002_8154# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X692 a_26058_14178# a_2346_14220# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X693 a_35002_5142# row_n[3] a_35494_5504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X694 a_9994_2130# a_2346_2172# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X695 VSS row_n[14] a_19334_16226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X696 a_23350_14218# rowon_n[12] a_22954_14178# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X697 a_29374_12210# col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X698 VSS row_n[9] a_20338_11206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X699 VSS row_n[8] a_33390_10202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X700 a_11302_4178# rowon_n[2] a_10906_4138# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X701 a_24050_17190# a_2346_17232# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X702 a_33998_11166# a_1962_11206# a_34090_11166# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X703 a_10298_10202# rowon_n[8] a_9902_10162# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X704 a_26458_4500# col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X705 a_24962_13174# a_1962_13214# a_25054_13174# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X706 a_17934_7150# a_1962_7190# a_18026_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X707 a_18938_3134# a_1962_3174# a_19030_3134# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X708 VDD VDD a_17934_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X709 a_28466_14540# col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X710 VDD rowon_n[10] a_31990_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X711 a_28066_10162# a_2346_10204# a_27974_10162# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X712 a_10998_5142# a_2346_5184# a_10906_5142# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X713 a_20034_3134# a_2346_3176# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X714 a_8990_15182# a_2346_15224# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X715 VSS row_n[7] a_8290_9198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X716 a_28978_10162# row_n[8] a_29470_10524# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X717 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X718 a_3270_3174# rowon_n[1] a_2874_3134# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X719 VDD rowon_n[2] a_10906_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X720 VSS VDD a_34394_18234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X721 a_31382_15222# col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X722 a_9902_10162# a_1962_10202# a_9994_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X723 vcm a_1962_6186# a_23046_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X724 a_11302_18234# VDD a_10906_18194# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X725 a_35398_14218# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X726 a_33086_6146# a_2346_6188# a_32994_6146# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X727 a_29070_18194# a_2346_18236# a_28978_18194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X728 VSS row_n[12] a_12306_14218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X729 a_20338_5182# rowon_n[3] a_19942_5142# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X730 a_30474_17552# col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X731 vcm a_1962_15222# a_26058_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X732 a_30074_13174# a_2346_13216# a_29982_13174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X733 a_8386_9520# col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X734 a_15014_7150# a_2346_7192# a_14922_7150# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X735 a_25054_1126# a_2346_1168# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X736 a_16018_3134# a_2346_3176# a_15926_3134# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X737 a_24050_5142# a_2346_5184# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X738 a_2874_17190# a_1962_17230# a_2966_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X739 a_9994_17190# a_2346_17232# a_9902_17190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X740 a_12914_17190# a_1962_17230# a_13006_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X741 VDD VSS a_2874_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X742 a_34490_16548# col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X743 a_30986_13174# row_n[11] a_31478_13536# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X744 VDD rowon_n[6] a_21950_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X745 vcm a_1962_5182# a_12002_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X746 VDD rowon_n[14] a_10906_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X747 vcm a_1962_10202# a_17022_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X748 a_9902_8154# row_n[6] a_10394_8516# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X749 a_8290_1166# VSS a_7894_1126# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X750 VSS row_n[2] a_34394_4178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X751 a_6890_14178# row_n[12] a_7382_14540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X752 a_16930_14178# row_n[12] a_17422_14540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X753 vcm a_1962_10202# a_6982_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X754 a_8990_9158# a_2346_9200# a_8898_9158# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X755 VDD rowon_n[1] a_19942_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X756 vcm a_1962_4178# a_28066_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X757 a_24354_7190# rowon_n[5] a_23958_7150# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X758 a_7986_2130# a_2346_2172# a_7894_2130# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X759 a_25358_3174# rowon_n[1] a_24962_3134# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X760 a_29070_3134# a_2346_3176# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X761 a_13310_3174# col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X762 a_15318_9198# rowon_n[7] a_14922_9158# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X763 a_32994_9158# a_1962_9198# a_33086_9158# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X764 a_32082_10162# a_2346_10204# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X765 VDD rowon_n[4] a_26970_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X766 vcm a_1962_3174# a_17022_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X767 a_34490_4500# col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X768 vcm a_1962_18234# a_7986_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X769 vcm a_1962_18234# a_18026_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X770 VSS row_n[15] a_26362_17230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X771 a_30378_15222# rowon_n[13] a_29982_15182# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X772 vcm a_1962_7190# a_16018_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X773 a_14922_6146# row_n[4] a_15414_6508# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X774 a_31990_2130# a_1962_2170# a_32082_2130# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X775 a_34394_14218# rowon_n[12] a_33998_14178# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X776 a_27366_13214# col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X777 VSS row_n[9] a_31382_11206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X778 VDD VSS a_24962_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X779 a_22042_18194# a_2346_18236# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X780 a_12914_1126# VDD a_13406_1488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X781 VSS row_n[3] a_19334_5182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X782 a_13006_17190# a_2346_17232# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X783 a_35094_17190# a_2346_17232# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X784 a_5278_2170# col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X785 a_29374_5182# rowon_n[3] a_28978_5142# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X786 a_2966_17190# a_2346_17232# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X787 a_22954_14178# a_1962_14218# a_23046_14178# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X788 VDD rowon_n[7] a_14922_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X789 a_7286_8194# rowon_n[6] a_6890_8154# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X790 a_18330_1166# en_bit_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X791 VDD VDD a_28978_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X792 a_6982_16186# a_2346_16228# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X793 a_17022_16186# a_2346_16228# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X794 a_26458_15544# col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X795 VDD rowon_n[11] a_29982_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X796 a_26058_11166# a_2346_11208# a_25966_11166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X797 vcm a_1962_2170# a_8990_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X798 a_30378_10202# col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X799 a_26970_11166# row_n[9] a_27462_11528# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X800 a_23046_1126# a_2346_1168# a_22954_1126# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X801 a_19430_3496# col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X802 a_22042_5142# a_2346_5184# a_21950_5142# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X803 VDD rowon_n[1] a_28978_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X804 a_24962_14178# row_n[12] a_25454_14540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X805 vcm a_1962_10202# a_25054_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X806 a_23958_7150# row_n[5] a_24450_7512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X807 a_8990_12170# a_2346_12212# a_8898_12170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X808 a_28370_9198# col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X809 a_19334_16226# col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X810 vcm a_1962_16226# a_24050_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X811 a_21950_2130# row_n[0] a_22442_2492# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X812 a_10906_18194# a_1962_18234# a_10998_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X813 a_18026_18194# a_2346_18236# a_17934_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X814 a_9294_16226# col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X815 VSS sample_n a_1962_7190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X816 a_7986_18194# a_2346_18236# a_7894_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X817 a_9390_12532# col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X818 a_27366_2170# col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X819 a_33390_3174# rowon_n[1] a_32994_3134# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X820 a_10998_3134# a_2346_3176# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X821 a_18426_18556# col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X822 a_27062_3134# a_2346_3176# a_26970_3134# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X823 a_8386_18556# col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X824 vcm a_1962_9198# a_31078_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X825 a_17326_8194# col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X826 a_3970_9158# a_2346_9200# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X827 a_27974_9158# row_n[7] a_28466_9520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X828 a_28978_5142# row_n[3] a_29470_5504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X829 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.64e+07u l=1.6e+07u
X830 a_6890_8154# row_n[6] a_7382_8516# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X831 VSS row_n[0] a_12306_2170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X832 a_22954_4138# a_1962_4178# a_23046_4138# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X833 a_32082_8154# a_2346_8196# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X834 VDD VSS a_32994_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X835 a_33086_4138# a_2346_4180# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X836 a_28370_15222# rowon_n[13] a_27974_15182# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X837 VSS row_n[10] a_25358_12210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X838 a_30074_11166# a_2346_11208# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X839 a_14410_5504# col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X840 a_2966_2130# a_2346_2172# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X841 VSS sample a_2346_16228# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X842 VSS row_n[9] a_29374_11206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X843 a_2346_5184# sample VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X844 a_15014_5142# a_2346_5184# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X845 a_16018_1126# a_2346_1168# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X846 a_9294_7190# col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X847 VDD rowon_n[12] a_23958_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X848 a_12002_12170# a_2346_12212# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X849 a_34090_12170# a_2346_12212# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X850 a_10906_7150# a_1962_7190# a_10998_7150# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X851 a_11910_3134# a_1962_3174# a_12002_3134# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X852 a_1962_12210# sample_n VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X853 a_9294_10202# rowon_n[8] a_8898_10162# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X854 VSS row_n[4] a_23350_6186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X855 a_33086_18194# a_2346_18236# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X856 VDD rowon_n[11] a_27974_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X857 a_25454_10524# col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X858 a_10998_18194# a_2346_18236# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X859 a_23350_17230# col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X860 a_33998_14178# a_1962_14218# a_34090_14178# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X861 a_4882_9158# a_1962_9198# a_4974_9158# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X862 VDD rowon_n[0] a_17934_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X863 a_29982_2130# row_n[0] a_30474_2492# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X864 a_3878_2130# a_1962_2170# a_3970_2130# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X865 VSS row_n[13] a_7286_15222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X866 VSS row_n[13] a_17326_15222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X867 a_22042_15182# a_2346_15224# a_21950_15182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X868 a_4274_12210# col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X869 a_14314_12210# col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X870 a_15926_5142# a_1962_5182# a_16018_5142# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X871 a_16930_1126# a_1962_1166# a_17022_1126# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X872 a_18330_11206# col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X873 vcm a_1962_11206# a_23046_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X874 a_35398_2170# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X875 VSS row_n[2] a_28370_4178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X876 a_22954_15182# row_n[13] a_23446_15544# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X877 a_17022_13174# a_2346_13216# a_16930_13174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X878 a_8290_11206# col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X879 VSS row_n[6] a_27366_8194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X880 a_6982_13174# a_2346_13216# a_6890_13174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X881 a_9902_13174# a_1962_13214# a_9994_13174# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X882 VDD rowon_n[15] a_5886_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X883 VDD rowon_n[15] a_15926_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X884 a_3366_14540# col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X885 a_13406_14540# col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X886 a_17422_13536# col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X887 a_13918_10162# row_n[8] a_14410_10524# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X888 a_7382_13536# col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X889 a_3878_10162# row_n[8] a_4370_10524# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X890 vcm a_1962_8194# a_20034_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X891 vcm a_1962_4178# a_21038_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X892 a_13310_4178# rowon_n[2] a_12914_4138# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X893 a_26970_9158# a_1962_9198# a_27062_9158# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X894 a_30074_8154# a_2346_8196# a_29982_8154# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X895 VSS row_n[5] a_16322_7190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X896 a_31078_4138# a_2346_4180# a_30986_4138# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X897 a_28466_4500# col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X898 a_6378_7512# col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X899 a_13006_5142# a_2346_5184# a_12914_5142# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X900 a_22042_3134# a_2346_3176# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X901 a_22346_17230# rowon_n[15] a_21950_17190# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X902 vcm a_1962_15222# a_10998_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X903 VDD rowon_n[4] a_19942_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X904 a_4882_18194# VDD a_5374_18556# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X905 a_14922_18194# VDD a_15414_18556# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X906 a_26362_16226# rowon_n[14] a_25966_16186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X907 vcm a_1962_14218# a_4974_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X908 vcm a_1962_14218# a_15014_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X909 VSS row_n[11] a_23350_13214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X910 a_8990_10162# a_2346_10204# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X911 VDD rowon_n[2] a_12914_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X912 vcm a_1962_6186# a_25054_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X913 a_35094_6146# a_2346_6188# a_35002_6146# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X914 a_27974_15182# a_1962_15222# a_28066_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X915 a_32082_13174# a_2346_13216# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X916 vcm a_1962_9198# a_2966_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X917 VDD rowon_n[13] a_21950_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X918 a_17326_11206# rowon_n[9] a_16930_11166# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X919 a_11302_1166# col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X920 a_22346_5182# rowon_n[3] a_21950_5142# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X921 VDD rowon_n[12] a_35002_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X922 a_7286_11206# rowon_n[9] a_6890_11166# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X923 a_17022_7150# a_2346_7192# a_16930_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X924 a_10298_5182# col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X925 a_27062_1126# a_2346_1168# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X926 a_18026_3134# a_2346_3176# a_17934_3134# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X927 a_23446_11528# col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X928 a_21342_18234# col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X929 VDD rowon_n[6] a_23958_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X930 vcm a_1962_5182# a_14010_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X931 a_34394_17230# col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X932 VDD rowon_n[1] a_21950_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X933 VSS row_n[15] a_11302_17230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X934 a_9902_3134# row_n[1] a_10394_3496# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X935 a_29982_18194# a_1962_18234# a_30074_18194# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X936 VSS row_n[14] a_15318_16226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X937 a_20034_16186# a_2346_16228# a_19942_16186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X938 a_12306_13214# col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X939 vcm a_1962_17230# a_29070_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X940 VSS row_n[14] a_5278_16226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X941 a_10998_15182# a_2346_15224# a_10906_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X942 a_33086_15182# a_2346_15224# a_32994_15182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X943 a_21342_9198# col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X944 VSS row_n[7] a_31382_9198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X945 a_26362_7190# rowon_n[5] a_25966_7150# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X946 a_9994_2130# a_2346_2172# a_9902_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X947 a_27366_3174# rowon_n[1] a_26970_3134# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X948 a_15318_3174# col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X949 a_20946_16186# row_n[14] a_21438_16548# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X950 a_5278_6186# rowon_n[4] a_4882_6146# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X951 a_33998_15182# row_n[13] a_34490_15544# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X952 a_15014_14178# a_2346_14220# a_14922_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X953 vcm a_1962_11206# a_34090_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X954 a_17326_9198# rowon_n[7] a_16930_9158# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X955 a_35002_9158# a_1962_9198# a_35094_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X956 a_19430_6508# col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X957 VDD VDD a_13918_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X958 a_11398_15544# col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X959 a_4974_14178# a_2346_14220# a_4882_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X960 vcm a_1962_7190# a_18026_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X961 VDD rowon_n[4] a_28978_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X962 vcm a_1962_3174# a_19030_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X963 VDD VDD a_3878_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X964 a_20034_3134# a_2346_3176# a_19942_3134# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X965 a_11910_11166# row_n[9] a_12402_11528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X966 a_33998_2130# a_1962_2170# a_34090_2130# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X967 VDD VSS a_26970_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X968 a_20946_9158# row_n[7] a_21438_9520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X969 a_26058_8154# a_2346_8196# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X970 a_14922_1126# VDD a_15414_1488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X971 a_21950_5142# row_n[3] a_22442_5504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X972 a_31478_9520# col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X973 a_9902_14178# row_n[12] a_10394_14540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X974 vcm a_1962_10202# a_9994_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X975 a_21342_12210# rowon_n[10] a_20946_12170# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X976 VDD rowon_n[7] a_16930_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X977 a_9294_8194# rowon_n[6] a_8898_8154# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X978 a_20338_18234# VDD a_19942_18194# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X979 a_1962_17230# sample_n VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X980 a_31382_1166# VSS a_30986_1126# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X981 a_17022_11166# a_2346_11208# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X982 a_25054_1126# a_2346_1168# a_24962_1126# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X983 VSS row_n[12] a_21342_14218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X984 a_6982_11166# a_2346_11208# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X985 a_24050_5142# a_2346_5184# a_23958_5142# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X986 a_2346_18236# sample VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X987 a_21950_17190# a_1962_17230# a_22042_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X988 VDD rowon_n[8] a_20946_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X989 a_25966_7150# row_n[5] a_26458_7512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X990 a_25966_16186# a_1962_16226# a_26058_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X991 a_30074_14178# a_2346_14220# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X992 a_19942_6146# a_1962_6186# a_20034_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X993 a_9994_18194# a_2346_18236# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X994 VDD rowon_n[14] a_19942_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X995 a_30074_6146# a_2346_6188# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X996 a_23958_2130# row_n[0] a_24450_2492# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X997 a_20338_13214# col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X998 a_33390_12210# col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X999 a_12002_7150# a_2346_7192# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1000 a_29374_2170# col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1001 a_13006_3134# a_2346_3176# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1002 a_3270_15222# rowon_n[13] a_2874_15182# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1003 a_13310_15222# rowon_n[13] a_12914_15182# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1004 VSS row_n[10] a_10298_12210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1005 a_7286_5182# col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1006 a_32386_18234# col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1007 a_19334_8194# col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1008 a_29070_3134# a_2346_3176# a_28978_3134# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1009 a_32482_14540# col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1010 vcm a_1962_12210# a_28066_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1011 VSS row_n[9] a_4274_11206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1012 VSS row_n[9] a_14314_11206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1013 a_32082_10162# a_2346_10204# a_31990_10162# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1014 vcm a_1962_9198# a_33086_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1015 a_19942_11166# row_n[9] a_20434_11528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1016 a_8898_8154# row_n[6] a_9390_8516# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1017 VSS row_n[6] a_20338_8194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1018 VSS row_n[2] a_21342_4178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1019 vcm a_1962_18234# a_27062_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1020 a_31078_16186# a_2346_16228# a_30986_16186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1021 a_32994_10162# row_n[8] a_33486_10524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1022 a_30378_8194# rowon_n[6] a_29982_8154# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1023 VSS row_n[0] a_14314_2170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1024 a_24962_4138# a_1962_4178# a_25054_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1025 a_34090_8154# a_2346_8196# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1026 VDD rowon_n[3] a_17934_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1027 vcm a_1962_2170# a_32082_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1028 a_35094_4138# a_2346_4180# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1029 a_29982_5142# row_n[3] a_30474_5504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1030 a_31990_16186# row_n[14] a_32482_16548# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1031 VDD rowon_n[11] a_2874_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1032 VDD rowon_n[11] a_12914_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1033 a_10394_10524# col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1034 a_4974_2130# a_2346_2172# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1035 a_6890_3134# row_n[1] a_7382_3496# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1036 a_17022_5142# a_2346_5184# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1037 a_18026_1126# a_2346_1168# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1038 a_13918_3134# a_1962_3174# a_14010_3134# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1039 a_21438_4500# col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1040 vcm a_1962_15222# a_30074_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1041 a_12914_7150# a_1962_7190# a_13006_7150# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1042 VSS row_n[4] a_25358_6186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1043 VSS row_n[7] a_3270_9198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1044 a_35398_6186# rowon_n[4] a_35002_6146# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1045 a_18330_18234# VDD a_17934_18194# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1046 a_32386_12210# rowon_n[10] a_31990_12170# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1047 VSS row_n[12] a_19334_14218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1048 a_29374_10202# col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1049 ctop sw ctop VDD sky130_fd_pr__pfet_01v8 ad=2.7075e+12p pd=2.185e+07u as=0p ps=0u w=1.9e+06u l=220000u
X1050 a_24050_15182# a_2346_15224# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1051 a_20946_12170# a_1962_12210# a_21038_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1052 a_5886_2130# a_1962_2170# a_5978_2130# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1053 a_18938_1126# a_1962_1166# a_19030_1126# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1054 a_17934_5142# a_1962_5182# a_18026_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1055 VDD rowon_n[14] a_17934_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1056 a_28466_12532# col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1057 VDD rowon_n[8] a_31990_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1058 a_3366_9520# col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1059 VSS row_n[6] a_29374_8194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1060 a_20034_1126# a_2346_1168# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1061 a_10998_3134# a_2346_3176# a_10906_3134# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1062 a_8990_13174# a_2346_13216# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1063 a_16418_8516# col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1064 VSS row_n[15] a_30378_17230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1065 a_3270_1166# VSS a_2874_1126# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1066 VSS row_n[14] a_34394_16226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1067 a_31382_13214# col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1068 a_3970_9158# a_2346_9200# a_3878_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1069 a_32386_7190# col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1070 a_11302_16226# rowon_n[14] a_10906_16186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1071 vcm a_1962_4178# a_23046_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1072 a_25054_17190# a_2346_17232# a_24962_17190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1073 a_28978_9158# a_1962_9198# a_29070_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1074 a_32082_8154# a_2346_8196# a_31990_8154# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1075 VSS row_n[5] a_18330_7190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1076 a_33086_4138# a_2346_4180# a_32994_4138# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1077 a_29070_16186# a_2346_16228# a_28978_16186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1078 vcm a_1962_13214# a_26058_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1079 a_2966_2130# a_2346_2172# a_2874_2130# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1080 a_20338_3174# rowon_n[1] a_19942_3134# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1081 VDD VDD a_32994_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1082 a_25966_17190# row_n[15] a_26458_17552# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1083 a_30474_15544# col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1084 a_30074_11166# a_2346_11208# a_29982_11166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1085 a_8386_7512# col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1086 a_15014_5142# a_2346_5184# a_14922_5142# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1087 a_16018_1126# a_2346_1168# a_15926_1126# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1088 a_24050_3134# a_2346_3176# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1089 a_2874_15182# a_1962_15222# a_2966_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1090 a_9994_15182# a_2346_15224# a_9902_15182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1091 a_12914_15182# a_1962_15222# a_13006_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1092 a_10298_9198# rowon_n[7] a_9902_9158# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1093 a_30986_11166# row_n[9] a_31478_11528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1094 VDD rowon_n[4] a_21950_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1095 a_6378_2492# col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1096 vcm a_1962_3174# a_12002_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1097 vcm a_1962_7190# a_10998_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1098 a_9902_6146# row_n[4] a_10394_6508# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1099 a_6890_12170# row_n[10] a_7382_12532# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1100 a_16930_12170# row_n[10] a_17422_12532# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1101 VDD en_bit_n[0] a_19942_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1102 vcm a_1962_9198# a_4974_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1103 a_25358_1166# VSS a_24962_1126# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1104 a_24354_5182# rowon_n[3] a_23958_5142# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1105 VDD rowon_n[7] a_9902_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1106 a_13310_1166# col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1107 a_29070_1126# a_2346_1168# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1108 vcm a_1962_17230# a_14010_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1109 a_27974_10162# a_1962_10202# a_28066_10162# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1110 vcm a_1962_2170# a_3970_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1111 vcm a_1962_17230# a_3970_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1112 VDD rowon_n[6] a_25966_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1113 vcm a_1962_1166# a_17022_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1114 a_29374_18234# VDD a_28978_18194# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1115 vcm a_1962_16226# a_7986_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1116 vcm a_1962_16226# a_18026_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1117 VSS row_n[13] a_26362_15222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1118 a_30378_13214# rowon_n[11] a_29982_13174# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1119 vcm a_1962_5182# a_16018_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1120 VDD sample a_2346_8196# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1121 a_27366_11206# col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1122 VDD rowon_n[1] a_23958_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1123 a_22042_16186# a_2346_16228# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1124 VSS row_n[1] a_19334_3174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1125 VDD rowon_n[15] a_24962_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1126 a_13006_15182# a_2346_15224# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1127 a_35094_15182# a_2346_15224# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1128 a_31990_12170# a_1962_12210# a_32082_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1129 a_23350_9198# col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1130 a_28370_7190# rowon_n[5] a_27974_7150# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1131 a_29374_3174# rowon_n[1] a_28978_3134# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1132 a_2966_15182# a_2346_15224# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1133 VSS row_n[7] a_33390_9198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1134 VDD rowon_n[5] a_14922_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1135 a_7286_6186# rowon_n[4] a_6890_6146# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1136 VDD rowon_n[14] a_28978_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1137 a_6982_14178# a_2346_14220# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1138 a_17022_14178# a_2346_14220# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1139 a_26458_13536# col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1140 VDD rowon_n[9] a_29982_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1141 vcm a_1962_9198# a_27062_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1142 a_22346_2170# col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1143 a_24050_12170# a_2346_12212# a_23958_12170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1144 a_19430_1488# en_bit_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1145 a_22042_3134# a_2346_3176# a_21950_3134# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1146 VSS row_n[10] a_9294_12210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1147 a_12306_8194# col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1148 a_28066_8154# a_2346_8196# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1149 VDD VSS a_28978_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1150 VSS VDD a_18330_18234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1151 a_23046_18194# a_2346_18236# a_22954_18194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1152 a_24962_12170# row_n[10] a_25454_12532# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1153 a_22954_9158# row_n[7] a_23446_9520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1154 a_23958_5142# row_n[3] a_24450_5504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1155 VSS VDD a_8290_18234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1156 a_8990_10162# a_2346_10204# a_8898_10162# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1157 a_33486_9520# col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1158 a_23958_18194# VDD a_24450_18556# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1159 a_19334_14218# col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1160 vcm a_1962_14218# a_24050_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1161 a_10906_16186# a_1962_16226# a_10998_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1162 a_18026_16186# a_2346_16228# a_17934_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1163 VDD rowon_n[12] a_7894_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1164 a_9294_14218# col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1165 VSS sample_n a_1962_5182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1166 a_7986_16186# a_2346_16228# a_7894_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1167 a_9390_10524# col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1168 a_33390_1166# VSS a_32994_1126# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1169 a_10998_1126# a_2346_1168# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1170 a_18426_16548# col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1171 a_4274_7190# col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1172 a_27062_1126# a_2346_1168# a_26970_1126# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1173 a_8386_16548# col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1174 a_17326_6186# col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1175 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X1176 a_27974_7150# row_n[5] a_28466_7512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1177 vcm a_1962_12210# a_13006_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1178 a_6890_6146# row_n[4] a_7382_6508# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1179 vcm a_1962_12210# a_2966_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1180 a_32082_6146# a_2346_6188# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1181 a_25966_2130# row_n[0] a_26458_2492# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1182 a_28370_13214# rowon_n[11] a_27974_13174# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1183 VSS row_n[8] a_25358_10202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1184 vcm a_1962_18234# a_12002_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1185 a_25966_11166# a_1962_11206# a_26058_11166# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1186 a_14010_7150# a_2346_7192# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1187 a_15014_3134# a_2346_3176# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1188 a_2346_3176# sample VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1189 a_9294_5182# col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1190 VSS sample_n a_1962_12210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1191 VDD rowon_n[10] a_23958_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1192 vcm a_1962_9198# a_35094_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1193 a_10906_5142# a_1962_5182# a_10998_5142# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1194 a_11910_1126# a_1962_1166# a_12002_1126# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1195 a_30378_2170# col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1196 a_18330_2170# rowon_n[0] a_17934_2130# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1197 VSS row_n[2] a_23350_4178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1198 a_28978_18194# a_1962_18234# a_29070_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1199 a_33086_16186# a_2346_16228# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1200 VDD rowon_n[9] a_27974_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1201 VSS row_n[6] a_22346_8194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1202 a_32386_8194# rowon_n[6] a_31990_8154# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1203 a_10998_16186# a_2346_16228# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1204 vcm a_1962_2170# a_34090_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1205 a_23350_15222# col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1206 a_26058_8154# a_2346_8196# a_25966_8154# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1207 a_8898_3134# row_n[1] a_9390_3496# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1208 a_6982_2130# a_2346_2172# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1209 a_16322_17230# rowon_n[15] a_15926_17190# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1210 a_6282_17230# rowon_n[15] a_5886_17190# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1211 a_21950_9158# a_1962_9198# a_22042_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1212 VSS row_n[5] a_11302_7190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1213 a_22442_17552# col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1214 VSS row_n[11] a_7286_13214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1215 VSS row_n[11] a_17326_13214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1216 a_22042_13174# a_2346_13216# a_21950_13174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1217 a_35094_12170# a_2346_12212# a_35002_12170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1218 a_4274_10202# col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1219 a_14314_10202# col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1220 a_14922_7150# a_1962_7190# a_15014_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1221 a_15926_3134# a_1962_3174# a_16018_3134# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1222 a_23446_4500# col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1223 a_2966_12170# a_2346_12212# a_2874_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1224 a_13006_12170# a_2346_12212# a_12914_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1225 a_22954_13174# row_n[11] a_23446_13536# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1226 a_17022_11166# a_2346_11208# a_16930_11166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1227 VSS row_n[4] a_27366_6186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1228 a_6982_11166# a_2346_11208# a_6890_11166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1229 VSS row_n[7] a_5278_9198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1230 VDD rowon_n[13] a_5886_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1231 VDD rowon_n[13] a_15926_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1232 a_3366_12532# col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1233 a_13406_12532# col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1234 a_17422_11528# col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1235 a_7382_11528# col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1236 vcm a_1962_6186# a_20034_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1237 a_15318_18234# col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1238 vcm a_1962_18234# a_20034_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1239 a_30074_6146# a_2346_6188# a_29982_6146# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1240 VSS row_n[3] a_16322_5182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1241 a_7894_2130# a_1962_2170# a_7986_2130# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1242 a_5278_18234# col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1243 vcm a_1962_17230# a_33086_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1244 a_5374_9520# col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1245 a_31990_8154# row_n[6] a_32482_8516# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1246 a_6378_5504# col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1247 a_24050_10162# a_2346_10204# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1248 a_18426_8516# col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1249 a_12002_7150# a_2346_7192# a_11910_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1250 a_22042_1126# a_2346_1168# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1251 a_13006_3134# a_2346_3176# a_12914_3134# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1252 a_10906_17190# row_n[15] a_11398_17552# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1253 a_22346_15222# rowon_n[13] a_21950_15182# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1254 vcm a_1962_13214# a_10998_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1255 a_4882_16186# row_n[14] a_5374_16548# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1256 a_14922_16186# row_n[14] a_15414_16548# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1257 a_26362_14218# rowon_n[12] a_25966_14178# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1258 VSS row_n[9] a_23350_11206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1259 a_16418_3496# col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1260 a_34394_7190# col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1261 vcm a_1962_4178# a_25054_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1262 a_27062_17190# a_2346_17232# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1263 a_34090_8154# a_2346_8196# a_33998_8154# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1264 a_35094_4138# a_2346_4180# a_35002_4138# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1265 a_27974_13174# a_1962_13214# a_28066_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1266 VDD rowon_n[11] a_21950_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1267 a_21342_7190# rowon_n[5] a_20946_7150# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1268 a_4974_2130# a_2346_2172# a_4882_2130# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1269 a_22346_3174# rowon_n[1] a_21950_3134# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1270 a_10298_3174# col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1271 VDD rowon_n[10] a_35002_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1272 a_17022_5142# a_2346_5184# a_16930_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1273 a_18026_1126# a_2346_1168# a_17934_1126# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1274 a_12306_9198# rowon_n[7] a_11910_9158# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1275 a_29982_9158# a_1962_9198# a_30074_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1276 a_21342_16226# col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1277 vcm a_1962_7190# a_13006_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1278 VDD rowon_n[4] a_23958_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1279 a_8386_2492# col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1280 vcm a_1962_3174# a_14010_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1281 a_34394_15222# col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1282 a_12914_10162# a_1962_10202# a_13006_10162# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1283 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X1284 a_2874_10162# a_1962_10202# a_2966_10162# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1285 VDD VSS a_21950_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1286 a_4274_18234# VDD a_3878_18194# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1287 a_14314_18234# VDD a_13918_18194# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1288 VSS row_n[13] a_11302_15222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1289 a_21038_8154# a_2346_8196# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1290 a_9902_1126# VDD a_10394_1488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1291 a_20434_18556# col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1292 a_29982_16186# a_1962_16226# a_30074_16186# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1293 VSS row_n[12] a_15318_14218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1294 a_20034_14178# a_2346_14220# a_19942_14178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1295 a_12306_11206# col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1296 a_33486_17552# col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1297 vcm a_1962_15222# a_29070_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1298 VSS row_n[12] a_5278_14218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1299 a_10998_13174# a_2346_13216# a_10906_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1300 a_33086_13174# a_2346_13216# a_32994_13174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1301 a_15318_1166# col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1302 a_27366_1166# VSS a_26970_1126# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1303 a_26362_5182# rowon_n[3] a_25966_5142# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1304 a_5886_17190# a_1962_17230# a_5978_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1305 a_15926_17190# a_1962_17230# a_16018_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1306 VDD rowon_n[7] a_11910_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1307 a_4274_8194# rowon_n[6] a_3878_8154# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1308 a_5278_4178# rowon_n[2] a_4882_4138# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1309 VDD rowon_n[15] a_9902_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1310 a_33998_13174# row_n[11] a_34490_13536# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1311 vcm a_1962_2170# a_5978_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1312 VDD rowon_n[14] a_13918_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1313 a_11398_13536# col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1314 VDD rowon_n[6] a_27974_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1315 vcm a_1962_5182# a_18026_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1316 vcm a_1962_1166# a_19030_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1317 VDD rowon_n[14] a_3878_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1318 a_20034_1126# a_2346_1168# a_19942_1126# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1319 a_20946_7150# row_n[5] a_21438_7512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1320 a_26058_6146# a_2346_6188# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1321 VDD rowon_n[1] a_25966_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1322 vcm a_1962_18234# a_31078_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1323 a_31478_7512# col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1324 VDD rowon_n[2] a_4882_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1325 a_9902_12170# row_n[10] a_10394_12532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1326 a_21342_10202# rowon_n[8] a_20946_10162# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1327 a_25358_9198# col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1328 a_22042_11166# a_2346_11208# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1329 VSS row_n[7] a_35398_9198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1330 a_2346_8196# sample VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1331 VDD rowon_n[5] a_16930_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1332 a_9294_6186# rowon_n[4] a_8898_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1333 a_13006_10162# a_2346_10204# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1334 a_35094_10162# a_2346_10204# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1335 vcm a_1962_9198# a_29070_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1336 a_20338_16226# rowon_n[14] a_19942_16186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1337 a_1962_15222# sample_n VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1338 a_2966_10162# a_2346_10204# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1339 a_24354_2170# col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1340 VDD rowon_n[0] a_14922_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1341 a_14314_8194# col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1342 a_24050_3134# a_2346_3176# a_23958_3134# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1343 a_25054_18194# a_2346_18236# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1344 a_2346_16228# sample VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1345 a_21950_15182# a_1962_15222# a_22042_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1346 a_24962_9158# row_n[7] a_25454_9520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1347 a_25966_5142# row_n[3] a_26458_5504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1348 a_16018_17190# a_2346_17232# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1349 a_35494_9520# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1350 a_3878_8154# row_n[6] a_4370_8516# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1351 a_5978_17190# a_2346_17232# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1352 a_25966_14178# a_1962_14218# a_26058_14178# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1353 a_19942_4138# a_1962_4178# a_20034_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1354 a_9994_16186# a_2346_16228# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1355 a_30074_4138# a_2346_4180# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1356 a_20338_11206# col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1357 a_33390_10202# col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1358 a_12002_5142# a_2346_5184# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1359 a_13006_1126# a_2346_1168# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1360 a_3270_13214# rowon_n[11] a_2874_13174# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1361 a_13310_13214# rowon_n[11] a_12914_13174# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1362 VSS row_n[8] a_10298_10202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1363 a_6282_7190# col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1364 a_7286_3174# col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1365 a_32386_16226# col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1366 a_10906_11166# a_1962_11206# a_10998_11166# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1367 a_19334_6186# col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1368 a_29070_1126# a_2346_1168# a_28978_1126# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1369 a_27974_14178# row_n[12] a_28466_14540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1370 a_32482_12532# col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1371 vcm a_1962_10202# a_28066_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1372 a_14922_12170# a_1962_12210# a_15014_12170# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1373 a_8898_6146# row_n[4] a_9390_6508# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1374 VSS row_n[4] a_20338_6186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1375 vcm a_1962_16226# a_27062_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1376 a_31078_14178# a_2346_14220# a_30986_14178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1377 a_4882_12170# a_1962_12210# a_4974_12170# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1378 a_30378_6186# rowon_n[4] a_29982_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1379 a_13918_18194# a_1962_18234# a_14010_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1380 a_31478_18556# col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1381 a_34090_6146# a_2346_6188# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1382 a_27974_2130# row_n[0] a_28466_2492# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1383 a_3878_18194# a_1962_18234# a_3970_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1384 VDD rowon_n[9] a_2874_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1385 VDD rowon_n[9] a_12914_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1386 a_6890_1126# VDD a_7382_1488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1387 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.64e+07u l=1.6e+07u
X1388 a_17022_3134# a_2346_3176# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1389 a_13918_1126# a_1962_1166# a_14010_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1390 a_29982_17190# row_n[15] a_30474_17552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1391 vcm a_1962_13214# a_30074_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1392 a_12914_5142# a_1962_5182# a_13006_5142# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1393 VSS row_n[6] a_24354_8194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1394 VSS row_n[2] a_25358_4178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1395 a_11398_8516# col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1396 a_34394_8194# rowon_n[6] a_33998_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1397 a_35398_4178# rowon_n[2] a_35002_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1398 a_18330_16226# rowon_n[14] a_17934_16186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1399 VSS row_n[10] a_28370_12210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1400 a_33086_11166# a_2346_11208# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1401 a_32386_10202# rowon_n[8] a_31990_10162# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1402 a_28066_8154# a_2346_8196# a_27974_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1403 a_8990_2130# a_2346_2172# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1404 a_10998_11166# a_2346_11208# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1405 a_24050_13174# a_2346_13216# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1406 a_19030_7150# a_2346_7192# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1407 VDD rowon_n[12] a_26970_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1408 a_15014_12170# a_2346_12212# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1409 a_23958_9158# a_1962_9198# a_24050_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1410 VSS row_n[5] a_13310_7190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1411 a_4974_12170# a_2346_12212# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1412 a_17934_3134# a_1962_3174# a_18026_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1413 VDD rowon_n[2] a_35002_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1414 a_25454_4500# col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1415 a_28466_10524# col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1416 a_3366_7512# col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1417 VSS row_n[4] a_29374_6186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1418 a_10998_1126# a_2346_1168# a_10906_1126# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1419 VSS row_n[7] a_7286_9198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1420 a_16418_6508# col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1421 a_33390_18234# VDD a_32994_18194# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1422 a_26362_17230# col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1423 VSS row_n[13] a_30378_15222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1424 VSS row_n[12] a_34394_14218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1425 a_31382_11206# col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1426 VSS row_n[0] a_6282_2170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1427 a_32386_5182# col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1428 a_35002_17190# a_1962_17230# a_35094_17190# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1429 a_11302_14218# rowon_n[12] a_10906_14178# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1430 a_25054_15182# a_2346_15224# a_24962_15182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1431 a_7286_12210# col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1432 a_17326_12210# col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1433 vcm a_1962_12210# a_22042_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1434 a_32082_6146# a_2346_6188# a_31990_6146# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1435 VSS row_n[3] a_18330_5182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1436 a_29070_14178# a_2346_14220# a_28978_14178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1437 vcm a_1962_11206# a_26058_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1438 a_33998_8154# row_n[6] a_34490_8516# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1439 a_20338_1166# en_bit_n[0] a_19942_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1440 a_29470_18556# col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1441 VDD rowon_n[14] a_32994_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1442 a_25966_15182# row_n[13] a_26458_15544# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1443 a_30474_13536# col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1444 a_7382_9520# col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1445 a_8386_5504# col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1446 a_24050_1126# a_2346_1168# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1447 a_15014_3134# a_2346_3176# a_14922_3134# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1448 a_2874_13174# a_1962_13214# a_2966_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1449 a_9994_13174# a_2346_13216# a_9902_13174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1450 a_12914_13174# a_1962_13214# a_13006_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1451 a_14010_7150# a_2346_7192# a_13918_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1452 VDD rowon_n[15] a_8898_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1453 a_6378_14540# col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1454 a_16418_14540# col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1455 VDD rowon_n[6] a_20946_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1456 vcm a_1962_1166# a_12002_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1457 a_31990_3134# row_n[1] a_32482_3496# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1458 vcm a_1962_5182# a_10998_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1459 a_18426_3496# col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1460 a_6890_10162# row_n[8] a_7382_10524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1461 a_16930_10162# row_n[8] a_17422_10524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1462 a_23350_7190# rowon_n[5] a_22954_7150# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1463 a_6982_2130# a_2346_2172# a_6890_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1464 a_24354_3174# rowon_n[1] a_23958_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1465 VDD rowon_n[5] a_9902_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1466 a_25358_17230# rowon_n[15] a_24962_17190# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1467 vcm a_1962_15222# a_14010_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1468 vcm a_1962_15222# a_3970_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1469 a_14314_9198# rowon_n[7] a_13918_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1470 vcm a_1962_9198# a_22042_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1471 VDD rowon_n[4] a_25966_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1472 a_17934_18194# VDD a_18426_18556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1473 a_29374_16226# rowon_n[14] a_28978_16186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1474 vcm a_1962_14218# a_7986_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1475 vcm a_1962_14218# a_18026_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1476 VSS row_n[11] a_26362_13214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1477 a_30378_11206# rowon_n[9] a_29982_11166# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1478 vcm a_1962_7190# a_15014_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1479 vcm a_1962_3174# a_16018_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1480 a_7894_18194# VDD a_8386_18556# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1481 VDD sample a_2346_6188# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1482 a_30986_2130# a_1962_2170# a_31078_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1483 a_23046_8154# a_2346_8196# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1484 VDD VSS a_23958_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1485 a_22042_14178# a_2346_14220# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1486 VSS en_bit_n[2] a_19334_1166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1487 VDD rowon_n[13] a_24962_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1488 a_13006_13174# a_2346_13216# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1489 a_35094_13174# a_2346_13216# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1490 a_29374_1166# VSS a_28978_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1491 a_28370_5182# rowon_n[3] a_27974_5142# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1492 a_2966_13174# a_2346_13216# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1493 a_25358_12210# col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1494 VDD rowon_n[7] a_13918_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1495 VDD rowon_n[3] a_14922_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1496 a_7286_4178# rowon_n[2] a_6890_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1497 a_26458_11528# col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1498 a_29982_11166# a_1962_11206# a_30074_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1499 a_6282_8194# rowon_n[6] a_5886_8154# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1500 vcm a_1962_2170# a_7986_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1501 a_24354_18234# col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1502 a_24450_14540# col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1503 a_24050_10162# a_2346_10204# a_23958_10162# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1504 a_22042_1126# a_2346_1168# a_21950_1126# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1505 VSS row_n[8] a_9294_10202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1506 a_12306_6186# col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1507 a_28066_6146# a_2346_6188# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1508 VDD rowon_n[1] a_27974_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1509 a_32994_18194# a_1962_18234# a_33086_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1510 VSS row_n[14] a_18330_16226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1511 a_23046_16186# a_2346_16228# a_22954_16186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1512 a_24962_10162# row_n[8] a_25454_10524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1513 a_22954_7150# row_n[5] a_23446_7512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1514 VSS row_n[14] a_8290_16226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1515 a_33486_7512# col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1516 VDD rowon_n[2] a_6890_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1517 a_23958_16186# row_n[14] a_24450_16548# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1518 a_20946_2130# row_n[0] a_21438_2492# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1519 a_10906_14178# a_1962_14218# a_10998_14178# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1520 a_18026_14178# a_2346_14220# a_17934_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1521 VDD rowon_n[10] a_7894_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1522 a_31478_2492# col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1523 VSS sample_n a_1962_3174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1524 VDD VDD a_16930_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1525 a_7986_14178# a_2346_14220# a_7894_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1526 VDD VDD a_6890_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1527 a_26362_2170# col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1528 VDD rowon_n[0] a_16930_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1529 a_4274_5182# col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1530 vcm a_1962_9198# a_30074_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1531 a_16322_8194# col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1532 a_17326_4178# col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1533 a_27974_5142# row_n[3] a_28466_5504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1534 vcm a_1962_10202# a_13006_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1535 a_5886_8154# row_n[6] a_6378_8516# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1536 a_2874_14178# row_n[12] a_3366_14540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1537 a_12914_14178# row_n[12] a_13406_14540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1538 a_24354_12210# rowon_n[10] a_23958_12170# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1539 a_2346_11208# sample VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1540 vcm a_1962_10202# a_2966_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1541 a_21950_10162# a_1962_10202# a_22042_10162# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1542 a_32082_4138# a_2346_4180# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1543 a_28370_11206# rowon_n[9] a_27974_11166# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1544 a_21038_8154# a_2346_8196# a_20946_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1545 a_3878_3134# row_n[1] a_4370_3496# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1546 vcm a_1962_16226# a_12002_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1547 a_1962_2170# sample_n VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1548 a_14010_5142# a_2346_5184# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1549 a_2346_1168# sample VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1550 a_15014_1126# a_2346_1168# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1551 a_16930_4138# row_n[2] a_17422_4500# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1552 a_9994_11166# a_2346_11208# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1553 a_8290_7190# col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1554 a_9294_3174# col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1555 VSS sample_n a_1962_10202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1556 VDD rowon_n[8] a_23958_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1557 a_9902_7150# a_1962_7190# a_9994_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1558 a_10906_3134# a_1962_3174# a_10998_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1559 VSS row_n[15] a_22346_17230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1560 a_28978_16186# a_1962_16226# a_29070_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1561 a_33086_14178# a_2346_14220# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1562 VSS row_n[4] a_22346_6186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1563 a_32386_6186# rowon_n[4] a_31990_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1564 a_10998_14178# a_2346_14220# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1565 a_23350_13214# col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1566 a_26058_6146# a_2346_6188# a_25966_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1567 a_8898_1126# VDD a_9390_1488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1568 a_16322_15222# rowon_n[13] a_15926_15182# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1569 VSS row_n[10] a_13310_12210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1570 a_6282_15222# rowon_n[13] a_5886_15182# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1571 VSS row_n[10] a_3270_12210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1572 VSS row_n[3] a_11302_5182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1573 a_2874_2130# a_1962_2170# a_2966_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1574 a_22442_15544# col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1575 a_35494_14540# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1576 VSS row_n[9] a_7286_11206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1577 VSS row_n[9] a_17326_11206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1578 a_22042_11166# a_2346_11208# a_21950_11166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1579 a_35094_10162# a_2346_10204# a_35002_10162# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1580 a_14922_5142# a_1962_5182# a_15014_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1581 a_15926_1126# a_1962_1166# a_16018_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1582 a_22954_11166# row_n[9] a_23446_11528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1583 a_2966_10162# a_2346_10204# a_2874_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1584 a_13006_10162# a_2346_10204# a_12914_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1585 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X1586 VSS row_n[2] a_27366_4178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1587 VDD rowon_n[12] a_11910_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1588 a_13406_8516# col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1589 VDD rowon_n[11] a_5886_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1590 VDD rowon_n[11] a_15926_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1591 a_3366_10524# col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1592 a_13406_10524# col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1593 a_11302_17230# col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1594 a_11398_3496# col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1595 vcm a_1962_4178# a_20034_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1596 a_15318_16226# col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1597 vcm a_1962_16226# a_20034_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1598 a_25966_9158# a_1962_9198# a_26058_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1599 VSS row_n[5] a_15318_7190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1600 VSS row_n[1] a_16322_3174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1601 a_30074_4138# a_2346_4180# a_29982_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1602 a_14010_18194# a_2346_18236# a_13918_18194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1603 a_5278_16226# col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1604 vcm a_1962_15222# a_33086_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1605 a_27462_4500# col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1606 a_3970_18194# a_2346_18236# a_3878_18194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1607 a_5374_7512# col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1608 a_31990_6146# row_n[4] a_32482_6508# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1609 a_5978_7150# a_2346_7192# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1610 a_18426_6508# col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1611 a_12002_5142# a_2346_5184# a_11910_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1612 a_13006_1126# a_2346_1168# a_12914_1126# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1613 a_14410_18556# col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1614 a_10906_15182# row_n[13] a_11398_15544# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1615 a_22346_13214# rowon_n[11] a_21950_13174# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1616 vcm a_1962_11206# a_10998_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1617 VSS row_n[7] a_9294_9198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1618 a_4370_18556# col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1619 a_35398_12210# rowon_n[10] a_35002_12170# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1620 a_3366_2492# col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1621 a_16418_1488# col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1622 a_27062_15182# a_2346_15224# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1623 a_23958_12170# a_1962_12210# a_24050_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1624 VSS row_n[0] a_8290_2170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1625 a_34394_5182# col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1626 a_34090_6146# a_2346_6188# a_33998_6146# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1627 VDD rowon_n[9] a_21950_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1628 a_9390_9520# col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1629 a_10298_1166# col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1630 a_22346_1166# VSS a_21950_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1631 a_21342_5182# rowon_n[3] a_20946_5142# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1632 VDD rowon_n[8] a_35002_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1633 a_17022_3134# a_2346_3176# a_16930_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1634 VSS VDD a_20338_18234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1635 VSS row_n[15] a_33390_17230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1636 a_33998_3134# row_n[1] a_34490_3496# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1637 a_21342_14218# col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1638 VDD rowon_n[6] a_22954_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1639 a_6890_7150# a_1962_7190# a_6982_7150# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1640 vcm a_1962_5182# a_13006_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1641 vcm a_1962_1166# a_14010_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1642 a_10298_17230# rowon_n[15] a_9902_17190# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1643 a_34394_13214# col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1644 VDD sample a_2346_18236# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1645 a_28066_17190# a_2346_17232# a_27974_17190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1646 a_4274_16226# rowon_n[14] a_3878_16186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1647 a_14314_16226# rowon_n[14] a_13918_16186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1648 VSS row_n[11] a_11302_13214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1649 a_21038_6146# a_2346_6188# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1650 VDD rowon_n[1] a_20946_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1651 a_20434_16548# col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1652 a_29982_14178# a_1962_14218# a_30074_14178# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1653 a_28978_17190# row_n[15] a_29470_17552# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1654 a_33486_15544# col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1655 vcm a_1962_13214# a_29070_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1656 a_10998_11166# a_2346_11208# a_10906_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1657 a_33086_11166# a_2346_11208# a_32994_11166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1658 a_20338_9198# col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1659 a_8990_2130# a_2346_2172# a_8898_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1660 a_26362_3174# rowon_n[1] a_25966_3134# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1661 a_5886_15182# a_1962_15222# a_5978_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1662 a_15926_15182# a_1962_15222# a_16018_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1663 VSS row_n[7] a_30378_9198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1664 VDD rowon_n[5] a_11910_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1665 a_4274_6186# rowon_n[4] a_3878_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1666 VDD rowon_n[13] a_9902_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1667 a_33998_11166# row_n[9] a_34490_11528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1668 a_16322_9198# rowon_n[7] a_15926_9158# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1669 vcm a_1962_9198# a_24050_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1670 a_19030_7150# a_2346_7192# a_18938_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1671 a_10298_12210# col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1672 a_11398_11528# col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1673 VDD rowon_n[4] a_27974_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1674 VDD rowon_n[0] a_9902_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1675 vcm a_1962_3174# a_18026_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1676 VDD VSS a_25966_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1677 a_32994_2130# a_1962_2170# a_33086_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1678 a_15318_2170# rowon_n[0] a_14922_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1679 a_26058_4138# a_2346_4180# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1680 a_19942_9158# row_n[7] a_20434_9520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1681 a_25054_8154# a_2346_8196# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1682 a_20946_5142# row_n[3] a_21438_5504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1683 vcm a_1962_16226# a_31078_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1684 a_30474_9520# col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1685 a_1962_7190# sample_n VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1686 a_31478_5504# col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1687 a_9902_10162# row_n[8] a_10394_10524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1688 vcm a_1962_17230# a_17022_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1689 VDD rowon_n[7] a_15926_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1690 a_8290_8194# rowon_n[6] a_7894_8154# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1691 a_2346_6188# sample VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1692 VDD rowon_n[3] a_16930_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1693 a_9294_4178# rowon_n[2] a_8898_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1694 vcm a_1962_17230# a_6982_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1695 a_20338_14218# rowon_n[12] a_19942_14178# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1696 a_1962_13214# sample_n VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1697 a_21038_17190# a_2346_17232# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1698 a_14314_6186# col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1699 a_24050_1126# a_2346_1168# a_23958_1126# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1700 a_25054_16186# a_2346_16228# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1701 a_21950_13174# a_1962_13214# a_22042_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1702 a_24962_7150# row_n[5] a_25454_7512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1703 a_16018_15182# a_2346_15224# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1704 a_35494_7512# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1705 a_3878_6146# row_n[4] a_4370_6508# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1706 a_5978_15182# a_2346_15224# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1707 VDD rowon_n[2] a_8898_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1708 a_9994_14178# a_2346_14220# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1709 VSS row_n[10] a_32386_12210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1710 a_22954_2130# row_n[0] a_23446_2492# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1711 a_33486_2492# col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1712 VSS VDD a_31382_18234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1713 a_28370_2170# col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1714 a_12002_3134# a_2346_3176# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1715 VDD rowon_n[12] a_30986_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1716 a_27062_12170# a_2346_12212# a_26970_12170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1717 a_3270_11206# rowon_n[9] a_2874_11166# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1718 a_13310_11206# rowon_n[9] a_12914_11166# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1719 a_6282_5182# col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1720 a_7286_1166# col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1721 a_32386_14218# col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1722 a_19334_4178# col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1723 a_26058_18194# a_2346_18236# a_25966_18194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1724 a_27974_12170# row_n[10] a_28466_12532# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1725 a_32482_10524# col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1726 a_18330_8194# col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1727 VSS row_n[2] a_20338_4178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1728 a_26970_18194# VDD a_27462_18556# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1729 a_30378_17230# col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1730 vcm a_1962_14218# a_27062_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1731 a_7894_8154# row_n[6] a_8386_8516# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1732 a_30378_4178# rowon_n[2] a_29982_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1733 a_13918_16186# a_1962_16226# a_14010_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1734 a_31478_16548# col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1735 vcm a_1962_2170# a_31078_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1736 a_34090_4138# a_2346_4180# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1737 a_3878_16186# a_1962_16226# a_3970_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1738 a_23046_8154# a_2346_8196# a_22954_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1739 a_3970_2130# a_2346_2172# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1740 a_5886_3134# row_n[1] a_6378_3496# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1741 a_17022_1126# a_2346_1168# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1742 vcm a_1962_17230# a_25054_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1743 a_18938_4138# row_n[2] a_19430_4500# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1744 vcm a_1962_11206# a_30074_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1745 a_20434_4500# col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1746 a_29982_15182# row_n[13] a_30474_15544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1747 a_12914_3134# a_1962_3174# a_13006_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1748 VDD rowon_n[2] a_29982_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1749 vcm a_1962_12210# a_16018_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1750 VSS row_n[4] a_24354_6186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1751 vcm a_1962_12210# a_5978_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1752 a_11398_6508# col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1753 a_34394_6186# rowon_n[4] a_33998_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1754 a_18330_14218# rowon_n[12] a_17934_14178# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1755 VSS row_n[8] a_28370_10202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1756 a_19030_17190# a_2346_17232# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1757 a_28978_11166# a_1962_11206# a_29070_11166# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1758 a_28066_6146# a_2346_6188# a_27974_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1759 a_20034_12170# a_2346_12212# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1760 a_19030_5142# a_2346_5184# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1761 VDD rowon_n[10] a_26970_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1762 VSS row_n[3] a_13310_5182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1763 a_4882_2130# a_1962_2170# a_4974_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1764 a_17934_1126# a_1962_1166# a_18026_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1765 a_3366_5504# col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1766 VSS row_n[2] a_29374_4178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1767 a_15414_8516# col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1768 a_16018_8154# a_2346_8196# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1769 VSS VDD a_29374_18234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1770 a_33390_16226# rowon_n[14] a_32994_16186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1771 a_26362_15222# col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1772 VSS row_n[11] a_30378_13214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1773 a_13406_3496# col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1774 a_19334_7190# rowon_n[5] a_18938_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1775 a_31382_7190# col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1776 a_32386_3174# col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1777 a_9294_17230# rowon_n[15] a_8898_17190# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1778 a_35002_15182# a_1962_15222# a_35094_15182# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1779 a_25454_17552# col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1780 a_21950_14178# row_n[12] a_22442_14540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1781 a_25054_13174# a_2346_13216# a_24962_13174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1782 a_7286_10202# col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1783 a_17326_10202# col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1784 vcm a_1962_10202# a_22042_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1785 a_27974_9158# a_1962_9198# a_28066_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1786 VSS row_n[5] a_17326_7190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1787 VSS row_n[1] a_18330_3174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1788 a_32082_4138# a_2346_4180# a_31990_4138# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1789 a_5978_12170# a_2346_12212# a_5886_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1790 a_16018_12170# a_2346_12212# a_15926_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1791 a_33998_6146# row_n[4] a_34490_6508# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1792 a_29470_4500# col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1793 a_29470_16548# col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1794 a_25966_13174# row_n[11] a_26458_13536# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1795 a_30474_11528# col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1796 a_7382_7512# col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1797 a_7986_7150# a_2346_7192# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1798 a_14010_5142# a_2346_5184# a_13918_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1799 a_15014_1126# a_2346_1168# a_14922_1126# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1800 a_9994_11166# a_2346_11208# a_9902_11166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1801 a_26970_2130# a_1962_2170# a_27062_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1802 VDD rowon_n[13] a_8898_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1803 a_6378_12532# col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1804 a_16418_12532# col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1805 VDD rowon_n[4] a_20946_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1806 a_31990_1126# VDD a_32482_1488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1807 a_5374_2492# col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1808 vcm a_1962_3174# a_10998_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1809 vcm a_1962_7190# a_9994_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1810 a_18426_1488# en_bit_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1811 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.64e+07u l=1.6e+07u
X1812 a_16930_8154# a_1962_8194# a_17022_8154# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1813 a_18330_18234# col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1814 vcm a_1962_18234# a_23046_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1815 a_8290_18234# col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1816 a_24354_1166# VSS a_23958_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1817 a_23350_5182# rowon_n[3] a_22954_5142# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1818 a_27062_10162# a_2346_10204# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1819 VDD rowon_n[3] a_9902_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1820 a_13918_17190# row_n[15] a_14410_17552# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1821 a_25358_15222# rowon_n[13] a_24962_15182# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1822 vcm a_1962_13214# a_14010_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1823 vcm a_1962_2170# a_2966_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1824 a_3878_17190# row_n[15] a_4370_17552# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1825 vcm a_1962_13214# a_3970_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1826 vcm a_1962_1166# a_16018_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1827 a_17934_16186# row_n[14] a_18426_16548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1828 a_29374_14218# rowon_n[12] a_28978_14178# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1829 VSS row_n[9] a_26362_11206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1830 a_8898_7150# a_1962_7190# a_8990_7150# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1831 vcm a_1962_5182# a_15014_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1832 a_7894_16186# row_n[14] a_8386_16548# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1833 a_31078_12170# a_2346_12212# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1834 a_23046_6146# a_2346_6188# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1835 VDD rowon_n[1] a_22954_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1836 VDD rowon_n[11] a_24962_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1837 a_28370_3174# rowon_n[1] a_27974_3134# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1838 a_25358_10202# col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1839 VSS row_n[7] a_32386_9198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1840 VDD rowon_n[5] a_13918_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1841 a_6282_6186# rowon_n[4] a_5886_6146# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1842 a_24354_16226# col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1843 vcm a_1962_9198# a_26058_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1844 a_8290_12210# rowon_n[10] a_7894_12170# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1845 a_15926_10162# a_1962_10202# a_16018_10162# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1846 VSS row_n[0] a_31382_2170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1847 a_21342_2170# col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1848 VDD rowon_n[0] a_11910_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1849 a_24450_12532# col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1850 a_5886_10162# a_1962_10202# a_5978_10162# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1851 a_5978_7150# a_2346_7192# a_5886_7150# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1852 a_7286_18234# VDD a_6890_18194# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1853 a_17326_18234# VDD a_16930_18194# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1854 a_11302_8194# col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1855 a_27062_8154# a_2346_8196# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1856 a_35002_2130# a_1962_2170# a_35094_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1857 VDD VSS a_27974_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1858 a_17326_2170# rowon_n[0] a_16930_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1859 a_28066_4138# a_2346_4180# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1860 a_12306_4178# col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1861 a_23446_18556# col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1862 a_32994_16186# a_1962_16226# a_33086_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1863 VSS row_n[12] a_18330_14218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1864 a_23046_14178# a_2346_14220# a_22954_14178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1865 a_22954_5142# row_n[3] a_23446_5504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1866 VSS row_n[12] a_8290_14218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1867 a_32482_9520# col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1868 a_33486_5504# col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1869 a_18938_17190# a_1962_17230# a_19030_17190# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1870 a_8898_17190# a_1962_17230# a_8990_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1871 VDD rowon_n[8] a_7894_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1872 VSS sample_n a_1962_1166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1873 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X1874 VDD rowon_n[14] a_16930_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1875 VDD rowon_n[14] a_6890_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1876 a_11910_4138# row_n[2] a_12402_4500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1877 vcm a_1962_12210# a_35094_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1878 a_3270_7190# col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1879 a_4274_3174# col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1880 a_16322_6186# col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1881 vcm a_1962_18234# a_34090_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1882 vcm a_1962_7190# a_6982_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1883 a_12914_12170# row_n[10] a_13406_12532# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1884 a_5886_6146# row_n[4] a_6378_6508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1885 a_2874_12170# row_n[10] a_3366_12532# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1886 a_25054_11166# a_2346_11208# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1887 a_24354_10202# rowon_n[8] a_23958_10162# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1888 a_16018_10162# a_2346_10204# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1889 a_21038_6146# a_2346_6188# a_20946_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1890 a_35494_2492# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1891 a_3878_1126# en_C0_n a_4370_1488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1892 a_24962_2130# row_n[0] a_25454_2492# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1893 a_11910_18194# VDD a_12402_18556# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1894 vcm a_1962_14218# a_12002_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1895 a_5978_10162# a_2346_10204# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1896 VDD rowon_n[12] a_18938_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1897 a_29070_12170# a_2346_12212# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1898 a_14010_3134# a_2346_3176# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1899 a_8290_5182# col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1900 a_9294_1166# col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1901 a_28066_18194# a_2346_18236# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1902 vcm a_1962_17230# a_9994_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1903 a_9902_5142# a_1962_5182# a_9994_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1904 a_10906_1126# a_1962_1166# a_10998_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1905 VSS row_n[2] a_22346_4178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1906 VSS row_n[13] a_22346_15222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1907 a_28978_14178# a_1962_14218# a_29070_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1908 a_32386_4178# rowon_n[2] a_31990_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1909 a_31382_8194# rowon_n[6] a_30986_8154# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1910 vcm a_1962_2170# a_33086_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1911 a_23350_11206# col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1912 a_25054_8154# a_2346_8196# a_24962_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1913 a_26058_4138# a_2346_4180# a_25966_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1914 a_7894_3134# row_n[1] a_8386_3496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1915 VDD rowon_n[15] a_20946_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1916 a_16322_13214# rowon_n[11] a_15926_13174# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1917 VSS row_n[8] a_13310_10202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1918 a_6282_13214# rowon_n[11] a_5886_13174# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1919 a_3878_11166# a_1962_11206# a_3970_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1920 a_13918_11166# a_1962_11206# a_14010_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1921 VSS row_n[8] a_3270_10202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1922 a_20946_9158# a_1962_9198# a_21038_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1923 VSS row_n[5] a_10298_7190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1924 VSS row_n[1] a_11302_3174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1925 a_22442_13536# col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1926 a_35494_12532# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1927 a_31078_9158# a_2346_9200# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1928 a_14922_3134# a_1962_3174# a_15014_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1929 a_22442_4500# col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1930 a_17934_12170# a_1962_12210# a_18026_12170# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1931 VDD rowon_n[2] a_31990_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1932 a_7894_12170# a_1962_12210# a_7986_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1933 VDD rowon_n[10] a_11910_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1934 a_13406_6508# col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1935 VSS row_n[7] a_4274_9198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1936 a_6890_18194# a_1962_18234# a_6982_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1937 a_16930_18194# a_1962_18234# a_17022_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1938 VDD rowon_n[9] a_5886_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1939 VDD rowon_n[9] a_15926_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1940 VSS VDD a_14314_18234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1941 a_11302_15222# col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1942 a_11398_1488# col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1943 VSS VDD a_4274_18234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1944 a_32082_17190# a_2346_17232# a_31990_17190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1945 VSS row_n[0] a_3270_2170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1946 a_19942_18194# VDD a_20434_18556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1947 a_15318_14218# col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1948 vcm a_1962_14218# a_20034_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1949 VSS row_n[3] a_15318_5182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1950 VSS VDD a_16322_1166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1951 a_32994_17190# row_n[15] a_33486_17552# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1952 a_14010_16186# a_2346_16228# a_13918_16186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1953 a_5278_14218# col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1954 vcm a_1962_13214# a_33086_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1955 a_10394_17552# col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1956 a_3970_16186# a_2346_16228# a_3878_16186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1957 a_4370_9520# col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1958 VDD rowon_n[6] a_18938_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1959 a_30986_8154# row_n[6] a_31478_8516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1960 a_5374_5504# col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1961 a_17422_8516# col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1962 a_5978_5142# a_2346_5184# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1963 a_12002_3134# a_2346_3176# a_11910_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1964 a_14410_16548# col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1965 a_10906_13174# row_n[11] a_11398_13536# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1966 a_22346_11206# rowon_n[9] a_21950_11166# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1967 a_18026_8154# a_2346_8196# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1968 analog_in sw ctop VSS sky130_fd_pr__nfet_01v8 ad=1.102e+12p pd=8.76e+06u as=2.7645e+12p ps=2.191e+07u w=1.9e+06u l=220000u
X1969 a_4370_16548# col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1970 a_35398_10202# rowon_n[8] a_35002_10162# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1971 VDD sample_n a_1962_7190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1972 a_15414_3496# col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1973 a_27062_13174# a_2346_13216# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1974 VSS row_n[7] a_26362_9198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1975 a_33390_7190# col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1976 a_34394_3174# col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1977 a_18026_12170# a_2346_12212# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1978 a_34090_4138# a_2346_4180# a_33998_4138# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1979 a_7986_12170# a_2346_12212# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1980 a_9390_7512# col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1981 a_3970_2130# a_2346_2172# a_3878_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1982 a_21342_3174# rowon_n[1] a_20946_3134# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1983 a_35002_10162# a_1962_10202# a_35094_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1984 a_9994_7150# a_2346_7192# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1985 a_17022_1126# a_2346_1168# a_16930_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1986 a_29374_17230# col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1987 VSS row_n[14] a_20338_16226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1988 VSS row_n[13] a_33390_15222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1989 a_11302_9198# rowon_n[7] a_10906_9158# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1990 a_28978_2130# a_1962_2170# a_29070_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1991 VDD rowon_n[4] a_22954_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1992 a_6890_5142# a_1962_5182# a_6982_5142# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1993 a_7382_2492# col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1994 vcm a_1962_3174# a_13006_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1995 a_10298_15222# rowon_n[13] a_9902_15182# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1996 a_34394_11206# col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1997 a_26458_9520# col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1998 a_18938_8154# a_1962_8194# a_19030_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1999 a_24962_18194# a_1962_18234# a_25054_18194# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2000 VDD sample a_2346_16228# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2001 VDD VSS a_20946_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2002 a_10298_2170# rowon_n[0] a_9902_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2003 a_21038_4138# a_2346_4180# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2004 VDD rowon_n[15] a_31990_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2005 a_28066_15182# a_2346_15224# a_27974_15182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2006 a_4274_14218# rowon_n[12] a_3878_14178# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2007 a_14314_14218# rowon_n[12] a_13918_14178# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2008 VSS row_n[9] a_11302_11206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2009 a_20034_8154# a_2346_8196# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2010 a_28978_15182# row_n[13] a_29470_15544# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2011 a_33486_13536# col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2012 vcm a_1962_11206# a_29070_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2013 VDD rowon_n[3] a_11910_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2014 a_26362_1166# VSS a_25966_1126# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2015 a_5886_13174# a_1962_13214# a_5978_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2016 a_15926_13174# a_1962_13214# a_16018_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2017 VDD rowon_n[7] a_10906_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2018 a_3270_8194# rowon_n[6] a_2874_8154# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2019 a_4274_4178# rowon_n[2] a_3878_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2020 VDD rowon_n[11] a_9902_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2021 vcm a_1962_2170# a_4974_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2022 a_19030_5142# a_2346_5184# a_18938_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2023 a_10298_10202# col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2024 vcm a_1962_1166# a_18026_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2025 a_30074_18194# a_2346_18236# a_29982_18194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2026 a_16018_8154# a_2346_8196# a_15926_8154# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2027 a_19942_7150# row_n[5] a_20434_7512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2028 a_25054_6146# a_2346_6188# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2029 a_30986_18194# VDD a_31478_18556# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2030 vcm a_1962_14218# a_31078_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2031 a_30474_7512# col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2032 a_1962_5182# sample_n VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2033 VDD rowon_n[2] a_3878_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2034 vcm a_1962_15222# a_17022_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2035 VSS row_n[7] a_34394_9198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2036 VDD rowon_n[5] a_15926_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2037 a_8290_6186# rowon_n[4] a_7894_6146# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2038 vcm a_1962_15222# a_6982_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2039 vcm a_1962_9198# a_28066_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2040 a_1962_11206# sample_n VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2041 a_23350_2170# col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2042 VDD rowon_n[0] a_13918_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2043 a_21038_15182# a_2346_15224# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2044 VSS row_n[0] a_33390_2170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2045 a_25358_8194# rowon_n[6] a_24962_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2046 a_7986_7150# a_2346_7192# a_7894_7150# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2047 a_14314_4178# col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2048 a_25054_14178# a_2346_14220# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2049 a_13310_8194# col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2050 a_29070_8154# a_2346_8196# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2051 vcm a_1962_2170# a_27062_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2052 a_24962_5142# row_n[3] a_25454_5504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2053 a_16018_13174# a_2346_13216# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2054 a_34490_9520# col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2055 a_35494_5504# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2056 a_5978_13174# a_2346_13216# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2057 a_28370_12210# col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2058 VSS row_n[8] a_32386_10202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2059 a_2874_8154# row_n[6] a_3366_8516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2060 vcm a_1962_8194# a_17022_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2061 a_32994_11166# a_1962_11206# a_33086_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2062 a_31990_7150# a_1962_7190# a_32082_7150# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2063 a_27366_18234# col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2064 VSS row_n[14] a_31382_16226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2065 a_12002_1126# a_2346_1168# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2066 a_27462_14540# col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2067 VDD rowon_n[10] a_30986_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2068 a_27062_10162# a_2346_10204# a_26970_10162# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2069 a_6282_3174# col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2070 a_13918_4138# row_n[2] a_14410_4500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2071 a_5278_7190# col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2072 a_26058_16186# a_2346_16228# a_25966_16186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2073 a_27974_10162# row_n[8] a_28466_10524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2074 a_18330_6186# col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2075 VDD VDD a_29982_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2076 vcm a_1962_7190# a_8990_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2077 a_26970_16186# row_n[14] a_27462_16548# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2078 a_30378_15222# col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2079 a_7894_6146# row_n[4] a_8386_6508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2080 a_13918_14178# a_1962_14218# a_14010_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2081 a_3878_14178# a_1962_14218# a_3970_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2082 a_23046_6146# a_2346_6188# a_22954_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2083 a_5886_1126# VDD a_6378_1488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2084 vcm a_1962_15222# a_25054_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2085 a_8990_17190# a_2346_17232# a_8898_17190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2086 a_29982_13174# row_n[11] a_30474_13536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2087 a_12914_1126# a_1962_1166# a_13006_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2088 vcm a_1962_10202# a_16018_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2089 VSS row_n[2] a_24354_4178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2090 a_9390_17552# col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2091 a_5886_14178# row_n[12] a_6378_14540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2092 a_15926_14178# row_n[12] a_16418_14540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2093 a_27366_12210# rowon_n[10] a_26970_12170# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2094 vcm a_1962_10202# a_5978_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2095 a_10394_8516# col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2096 a_10998_8154# a_2346_8196# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2097 a_33390_8194# rowon_n[6] a_32994_8154# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2098 a_27366_7190# col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2099 a_34394_4178# rowon_n[2] a_33998_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2100 vcm a_1962_2170# a_35094_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2101 a_19030_15182# a_2346_15224# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2102 a_27062_8154# a_2346_8196# a_26970_8154# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2103 a_28066_4138# a_2346_4180# a_27974_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2104 a_19030_3134# a_2346_3176# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2105 VDD rowon_n[8] a_26970_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2106 a_22954_9158# a_1962_9198# a_23046_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2107 VSS row_n[5] a_12306_7190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2108 VSS row_n[1] a_13310_3174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2109 a_33086_9158# a_2346_9200# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2110 VDD rowon_n[2] a_33998_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2111 a_24450_4500# col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2112 VSS row_n[15] a_25358_17230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2113 a_2966_7150# a_2346_7192# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2114 a_15414_6508# col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2115 a_16018_6146# a_2346_6188# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2116 a_21950_2130# a_1962_2170# a_22042_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2117 VSS row_n[14] a_29374_16226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2118 a_33390_14218# rowon_n[12] a_32994_14178# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2119 a_26362_13214# col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2120 VSS row_n[9] a_30378_11206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2121 a_13406_1488# col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2122 a_12002_17190# a_2346_17232# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2123 a_34090_17190# a_2346_17232# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2124 VSS row_n[10] a_16322_12210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2125 a_21038_12170# a_2346_12212# a_20946_12170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2126 a_11910_8154# a_1962_8194# a_12002_8154# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2127 a_32386_1166# col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2128 a_31382_5182# col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2129 a_19334_5182# rowon_n[3] a_18938_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2130 a_1962_17230# sample_n VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2131 a_9294_15222# rowon_n[13] a_8898_15182# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2132 a_35002_13174# a_1962_13214# a_35094_13174# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2133 VSS row_n[10] a_6282_12210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2134 VSS row_n[0] a_5278_2170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2135 VDD VDD a_27974_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2136 a_25454_15544# col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2137 a_21950_12170# row_n[10] a_22442_12532# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2138 a_25054_11166# a_2346_11208# a_24962_11166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2139 VSS row_n[3] a_17326_5182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2140 VSS en_bit_n[1] a_18330_1166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2141 a_5978_10162# a_2346_10204# a_5886_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2142 a_16018_10162# a_2346_10204# a_15926_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2143 VDD rowon_n[12] a_14922_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2144 a_25966_11166# row_n[9] a_26458_11528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2145 a_32994_8154# row_n[6] a_33486_8516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2146 a_7382_5504# col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2147 a_7986_5142# a_2346_5184# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2148 a_14010_3134# a_2346_3176# a_13918_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2149 VDD rowon_n[12] a_4882_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2150 VDD rowon_n[11] a_8898_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2151 a_6378_10524# col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2152 a_16418_10524# col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2153 vcm a_1962_1166# a_10998_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2154 a_30986_3134# row_n[1] a_31478_3496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2155 VDD rowon_n[1] a_18938_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2156 a_14314_17230# col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2157 a_3878_7150# a_1962_7190# a_3970_7150# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2158 vcm a_1962_5182# a_9994_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2159 a_4274_17230# col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2160 a_16930_6146# a_1962_6186# a_17022_6146# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2161 a_17422_3496# col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2162 a_18330_16226# col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2163 vcm a_1962_16226# a_23046_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2164 VSS row_n[7] a_28370_9198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2165 a_35398_7190# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2166 a_9902_18194# a_1962_18234# a_9994_18194# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2167 a_17022_18194# a_2346_18236# a_16930_18194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2168 a_8290_16226# col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2169 a_6982_18194# a_2346_18236# a_6890_18194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2170 a_23350_3174# rowon_n[1] a_22954_3134# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2171 a_17422_18556# col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2172 a_13918_15182# row_n[13] a_14410_15544# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2173 a_25358_13214# rowon_n[11] a_24962_13174# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2174 vcm a_1962_11206# a_14010_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2175 a_7382_18556# col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2176 a_3878_15182# row_n[13] a_4370_15544# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2177 vcm a_1962_11206# a_3970_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2178 a_13310_9198# rowon_n[7] a_12914_9158# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2179 vcm a_1962_9198# a_21038_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2180 a_31078_9158# a_2346_9200# a_30986_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2181 a_8898_5142# a_1962_5182# a_8990_5142# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2182 a_9390_2492# col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2183 vcm a_1962_3174# a_15014_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2184 a_28466_9520# col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2185 a_26970_12170# a_1962_12210# a_27062_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2186 a_22042_8154# a_2346_8196# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2187 VDD VSS a_22954_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2188 a_29982_2130# a_1962_2170# a_30074_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2189 a_12306_2170# rowon_n[0] a_11910_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2190 a_23046_4138# a_2346_4180# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2191 VSS row_n[10] a_24354_12210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2192 VDD sample a_2346_11208# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2193 VDD rowon_n[9] a_24962_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2194 a_28370_1166# VSS a_27974_1126# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2195 VDD rowon_n[7] a_12914_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2196 VDD rowon_n[3] a_13918_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2197 a_6282_4178# rowon_n[2] a_5886_4138# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2198 VSS VDD a_23350_18234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2199 VDD rowon_n[12] a_22954_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2200 a_24354_14218# col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2201 a_19030_12170# a_2346_12212# a_18938_12170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2202 a_8290_10202# rowon_n[8] a_7894_10162# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2203 a_32082_18194# a_2346_18236# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2204 a_24450_10524# col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2205 a_5978_5142# a_2346_5184# a_5886_5142# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2206 a_7286_16226# rowon_n[14] a_6890_16186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2207 a_17326_16226# rowon_n[14] a_16930_16186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2208 a_18026_8154# a_2346_8196# a_17934_8154# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2209 a_11302_6186# col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2210 a_27062_6146# a_2346_6188# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2211 a_23446_16548# col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2212 a_32994_14178# a_1962_14218# a_33086_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2213 a_32482_7512# col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2214 VDD rowon_n[2] a_5886_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2215 a_18938_15182# a_1962_15222# a_19030_15182# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2216 a_8898_15182# a_1962_15222# a_8990_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2217 a_30474_2492# col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2218 a_19942_2130# row_n[0] a_20434_2492# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2219 a_3270_12210# col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2220 a_13310_12210# col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2221 a_25358_2170# col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2222 VDD rowon_n[0] a_15926_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2223 a_12306_18234# col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2224 a_35002_14178# row_n[12] a_35494_14540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2225 vcm a_1962_10202# a_35094_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2226 a_27366_8194# rowon_n[6] a_26970_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2227 a_9994_7150# a_2346_7192# a_9902_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2228 a_3270_5182# col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2229 VSS row_n[0] a_35398_2170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2230 a_4274_1166# en_C0_n VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2231 a_15318_8194# col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2232 vcm a_1962_2170# a_29070_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2233 a_16322_4178# col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2234 vcm a_1962_16226# a_34090_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2235 a_12402_14540# col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2236 a_21038_10162# a_2346_10204# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2237 vcm a_1962_5182# a_6982_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2238 a_12914_10162# row_n[8] a_13406_10524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2239 a_4882_8154# row_n[6] a_5374_8516# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2240 a_2874_10162# row_n[8] a_3366_10524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2241 vcm a_1962_8194# a_19030_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2242 a_20034_8154# a_2346_8196# a_19942_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2243 a_21038_4138# a_2346_4180# a_20946_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2244 a_11910_16186# row_n[14] a_12402_16548# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2245 a_33998_7150# a_1962_7190# a_34090_7150# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2246 a_2874_3134# row_n[1] a_3366_3496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2247 VDD rowon_n[10] a_18938_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2248 a_14010_1126# a_2346_1168# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2249 a_8290_3174# col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2250 a_15926_4138# row_n[2] a_16418_4500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2251 a_21342_17230# rowon_n[15] a_20946_17190# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2252 a_28066_16186# a_2346_16228# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2253 vcm a_1962_15222# a_9994_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2254 a_9902_3134# a_1962_3174# a_9994_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2255 VSS row_n[11] a_22346_13214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2256 a_31382_6186# rowon_n[4] a_30986_6146# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2257 VSS row_n[10] a_35398_12210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2258 a_12306_12210# rowon_n[10] a_11910_12170# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2259 a_25054_6146# a_2346_6188# a_24962_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2260 a_7894_1126# VDD a_8386_1488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2261 VDD rowon_n[13] a_20946_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2262 a_6282_11206# rowon_n[9] a_5886_11166# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2263 a_16322_11206# rowon_n[9] a_15926_11166# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2264 a_26970_8154# row_n[6] a_27462_8516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2265 VDD rowon_n[12] a_33998_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2266 VSS row_n[3] a_10298_5182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2267 VSS VDD a_11302_1166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2268 a_22442_11528# col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2269 a_35494_10524# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2270 a_14922_1126# a_1962_1166# a_15014_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2271 a_20338_18234# col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2272 a_33390_17230# col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2273 VDD rowon_n[8] a_11910_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2274 a_12402_8516# col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2275 a_13006_8154# a_2346_8196# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2276 a_29374_7190# col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2277 VSS row_n[15] a_10298_17230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2278 a_6890_16186# a_1962_16226# a_6982_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2279 a_16930_16186# a_1962_16226# a_17022_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2280 a_29070_8154# a_2346_8196# a_28978_8154# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2281 VSS row_n[14] a_14314_16226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2282 a_11302_13214# col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2283 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.64e+07u l=1.6e+07u
X2284 a_10394_3496# col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2285 vcm a_1962_17230# a_28066_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2286 VSS row_n[14] a_4274_16226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2287 a_32082_15182# a_2346_15224# a_31990_15182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2288 VSS row_n[7] a_21342_9198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2289 a_19942_16186# row_n[14] a_20434_16548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2290 a_19030_10162# a_2346_10204# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2291 VSS row_n[1] a_15318_3174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2292 a_32994_15182# row_n[13] a_33486_15544# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2293 a_14010_14178# a_2346_14220# a_13918_14178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2294 vcm a_1962_11206# a_33086_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2295 a_24962_9158# a_1962_9198# a_25054_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2296 a_35094_9158# a_2346_9200# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2297 VSS row_n[5] a_14314_7190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2298 vcm a_1962_7190# a_32082_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2299 VDD VDD a_12914_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2300 a_10394_15544# col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2301 a_3970_14178# a_2346_14220# a_3878_14178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2302 a_4370_7512# col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2303 VDD rowon_n[4] a_18938_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2304 a_30986_6146# row_n[4] a_31478_6508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2305 VDD VDD a_2874_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2306 vcm a_1962_12210# a_8990_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2307 vcm a_1962_12210# a_19030_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2308 a_4974_7150# a_2346_7192# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2309 a_17422_6508# col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2310 a_12002_1126# a_2346_1168# a_11910_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2311 a_5978_3134# a_2346_3176# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2312 a_10906_11166# row_n[9] a_11398_11528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2313 a_18026_6146# a_2346_6188# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2314 a_23958_2130# a_1962_2170# a_24050_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2315 VSS sample a_2346_9200# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2316 VDD sample_n a_1962_5182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2317 ctop sw analog_in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.9e+06u l=220000u
X2318 a_23046_12170# a_2346_12212# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2319 a_21438_9520# col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2320 a_13918_8154# a_1962_8194# a_14010_8154# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2321 a_15414_1488# col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2322 VSS row_n[0] a_7286_2170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2323 a_33390_5182# col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2324 a_32386_17230# rowon_n[15] a_31990_17190# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2325 a_35002_8154# row_n[6] a_35494_8516# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2326 a_9390_5504# col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2327 a_21342_1166# VSS a_20946_1126# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2328 a_9994_5142# a_2346_5184# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2329 a_29374_15222# col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2330 VSS row_n[12] a_20338_14218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2331 VSS row_n[11] a_33390_13214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2332 a_20946_17190# a_1962_17230# a_21038_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2333 a_5886_7150# a_1962_7190# a_5978_7150# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2334 vcm a_1962_1166# a_13006_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2335 a_32994_3134# row_n[1] a_33486_3496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2336 a_6890_3134# a_1962_3174# a_6982_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2337 a_10298_13214# rowon_n[11] a_9902_13174# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2338 a_26458_7512# col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2339 a_18938_6146# a_1962_6186# a_19030_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2340 a_24962_16186# a_1962_16226# a_25054_16186# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2341 a_8990_18194# a_2346_18236# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2342 a_28466_17552# col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2343 VDD rowon_n[13] a_31990_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2344 a_28066_13174# a_2346_13216# a_27974_13174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2345 a_10998_8154# a_2346_8196# a_10906_8154# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2346 a_20034_6146# a_2346_6188# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2347 a_11910_12170# a_1962_12210# a_12002_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2348 a_28978_13174# row_n[11] a_29470_13536# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2349 VDD sample_n a_1962_12210# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2350 a_33486_11528# col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2351 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.64e+07u l=1.6e+07u
X2352 VDD rowon_n[9] a_9902_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2353 VDD rowon_n[5] a_10906_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2354 a_3270_6186# rowon_n[4] a_2874_6146# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2355 a_31382_18234# col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2356 vcm a_1962_9198# a_23046_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2357 a_19030_3134# a_2346_3176# a_18938_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2358 a_33086_9158# a_2346_9200# a_32994_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2359 vcm a_1962_18234# a_26058_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2360 a_30074_16186# a_2346_16228# a_29982_16186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2361 a_20338_8194# rowon_n[6] a_19942_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2362 a_2966_7150# a_2346_7192# a_2874_7150# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2363 a_24050_8154# a_2346_8196# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2364 a_16018_6146# a_2346_6188# a_15926_6146# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2365 vcm a_1962_2170# a_22042_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2366 a_14314_2170# rowon_n[0] a_13918_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2367 a_25054_4138# a_2346_4180# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2368 a_19942_5142# row_n[3] a_20434_5504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2369 a_30986_16186# row_n[14] a_31478_16548# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2370 a_2346_14220# sample VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2371 a_1962_3174# sample_n VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2372 a_30474_5504# col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2373 vcm a_1962_8194# a_12002_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2374 a_16930_17190# row_n[15] a_17422_17552# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2375 vcm a_1962_13214# a_17022_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2376 VDD rowon_n[3] a_15926_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2377 a_8290_4178# rowon_n[2] a_7894_4138# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2378 a_6890_17190# row_n[15] a_7382_17552# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2379 vcm a_1962_13214# a_6982_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2380 a_21038_13174# a_2346_13216# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2381 a_25358_6186# rowon_n[4] a_24962_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2382 a_7986_5142# a_2346_5184# a_7894_5142# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2383 a_13310_6186# col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2384 a_29070_6146# a_2346_6188# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2385 a_31382_12210# rowon_n[10] a_30986_12170# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2386 vcm a_1962_7190# a_3970_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2387 a_34490_7512# col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2388 a_2874_6146# row_n[4] a_3366_6508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2389 a_28370_10202# col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2390 vcm a_1962_6186# a_17022_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2391 VDD rowon_n[2] a_7894_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2392 a_30378_18234# VDD a_29982_18194# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2393 a_19942_12170# a_1962_12210# a_20034_12170# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2394 a_32482_2492# col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2395 a_31990_5142# a_1962_5182# a_32082_5142# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2396 a_27366_16226# col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2397 VSS row_n[12] a_31382_14218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2398 a_18938_10162# a_1962_10202# a_19030_10162# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2399 a_31990_17190# a_1962_17230# a_32082_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2400 a_27462_12532# col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2401 a_8898_10162# a_1962_10202# a_8990_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2402 VDD rowon_n[8] a_30986_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2403 VSS row_n[6] a_19334_8194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2404 a_6282_1166# col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2405 a_29374_8194# rowon_n[6] a_28978_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2406 a_5278_5182# col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2407 a_26058_14178# a_2346_14220# a_25966_14178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2408 a_18330_4178# col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2409 a_26458_18556# col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2410 VDD rowon_n[14] a_29982_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2411 vcm a_1962_5182# a_8990_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2412 a_30378_13214# col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2413 a_22346_7190# col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2414 vcm a_1962_2170# a_30074_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2415 VSS row_n[15] a_9294_17230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2416 a_24050_17190# a_2346_17232# a_23958_17190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2417 a_22042_8154# a_2346_8196# a_21950_8154# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2418 a_4882_3134# row_n[1] a_5374_3496# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2419 a_23046_4138# a_2346_4180# a_22954_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2420 vcm a_1962_13214# a_25054_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2421 a_24962_17190# row_n[15] a_25454_17552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2422 a_17934_4138# row_n[2] a_18426_4500# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2423 a_8990_15182# a_2346_15224# a_8898_15182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2424 a_29982_11166# row_n[9] a_30474_11528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2425 a_9390_15544# col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2426 a_5886_12170# row_n[10] a_6378_12532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2427 a_15926_12170# row_n[10] a_16418_12532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2428 a_28066_11166# a_2346_11208# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2429 a_27366_10202# rowon_n[8] a_26970_10162# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2430 a_10394_6508# col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2431 a_10998_6146# a_2346_6188# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2432 a_33390_6186# rowon_n[4] a_32994_6146# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2433 a_27366_5182# col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2434 a_19030_13174# a_2346_13216# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2435 a_27062_6146# a_2346_6188# a_26970_6146# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2436 a_28978_8154# row_n[6] a_29470_8516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2437 a_19030_1126# a_2346_1168# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2438 vcm a_1962_17230# a_13006_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2439 VSS row_n[3] a_12306_5182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2440 VSS VDD a_13310_1166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2441 vcm a_1962_17230# a_2966_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2442 a_26970_3134# row_n[1] a_27462_3496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2443 a_28370_18234# VDD a_27974_18194# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2444 VSS row_n[13] a_25358_15222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2445 a_22346_12210# col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2446 a_2966_5142# a_2346_5184# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2447 a_14410_8516# col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2448 a_16018_4138# a_2346_4180# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2449 VSS row_n[12] a_29374_14218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2450 a_26362_11206# col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2451 a_2346_8196# sample VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2452 a_15014_8154# a_2346_8196# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2453 VSS sample_n a_1962_17230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2454 VDD rowon_n[15] a_23958_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2455 a_12002_15182# a_2346_15224# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2456 a_34090_15182# a_2346_15224# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2457 a_21438_14540# col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2458 a_30986_12170# a_1962_12210# a_31078_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2459 VSS row_n[8] a_16322_10202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2460 a_21038_10162# a_2346_10204# a_20946_10162# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2461 a_18330_7190# rowon_n[5] a_17934_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2462 a_11910_6146# a_1962_6186# a_12002_6146# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2463 a_31382_3174# col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2464 a_19334_3174# rowon_n[1] a_18938_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2465 a_12402_3496# col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2466 a_1962_15222# sample_n VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2467 a_9294_13214# rowon_n[11] a_8898_13174# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2468 a_6890_11166# a_1962_11206# a_6982_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2469 a_16930_11166# a_1962_11206# a_17022_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2470 VSS row_n[8] a_6282_10202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2471 VSS row_n[7] a_23350_9198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2472 a_30378_7190# col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2473 VDD rowon_n[14] a_27974_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2474 a_25454_13536# col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2475 a_21950_10162# row_n[8] a_22442_10524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2476 VSS row_n[1] a_17326_3174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2477 vcm a_1962_7190# a_34090_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2478 a_32994_6146# row_n[4] a_33486_6508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2479 VDD rowon_n[10] a_14922_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2480 a_14010_1126# a_2346_1168# a_13918_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2481 a_7986_3134# a_2346_3176# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2482 VDD rowon_n[10] a_4882_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2483 a_6982_7150# a_2346_7192# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2484 a_25966_2130# a_1962_2170# a_26058_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2485 VDD rowon_n[9] a_8898_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2486 VDD en_bit_n[2] a_18938_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2487 a_30986_1126# VDD a_31478_1488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2488 VSS VDD a_17326_18234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2489 a_22042_18194# a_2346_18236# a_21950_18194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2490 a_14314_15222# col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2491 a_3878_5142# a_1962_5182# a_3970_5142# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2492 a_4370_2492# col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2493 vcm a_1962_3174# a_9994_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2494 VSS VDD a_7286_18234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2495 a_13006_17190# a_2346_17232# a_12914_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2496 a_35094_17190# a_2346_17232# a_35002_17190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2497 a_4274_15222# col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2498 a_23446_9520# col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2499 a_15926_8154# a_1962_8194# a_16018_8154# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2500 a_17422_1488# col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2501 a_16930_4138# a_1962_4178# a_17022_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2502 a_22954_18194# VDD a_23446_18556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2503 a_2966_17190# a_2346_17232# a_2874_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2504 a_18330_14218# col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2505 vcm a_1962_14218# a_23046_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2506 VSS row_n[0] a_9294_2170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2507 VSS sample a_2346_4180# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2508 a_35398_5182# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2509 a_9902_16186# a_1962_16226# a_9994_16186# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2510 a_17022_16186# a_2346_16228# a_16930_16186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2511 a_8290_14218# col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2512 a_13406_17552# col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2513 a_6982_16186# a_2346_16228# a_6890_16186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2514 a_23350_1166# VSS a_22954_1126# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2515 a_3366_17552# col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2516 a_17422_16548# col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2517 a_13918_13174# row_n[11] a_14410_13536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2518 a_25358_11206# rowon_n[9] a_24962_11166# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2519 a_7382_16548# col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2520 a_3878_13174# row_n[11] a_4370_13536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2521 a_35002_3134# row_n[1] a_35494_3496# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2522 a_7894_7150# a_1962_7190# a_7986_7150# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2523 vcm a_1962_1166# a_15014_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2524 a_8898_3134# a_1962_3174# a_8990_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2525 a_28466_7512# col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2526 a_13006_8154# a_2346_8196# a_12914_8154# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2527 a_22042_6146# a_2346_6188# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2528 ctop sw_n analog_in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.102e+12p ps=8.76e+06u w=1.9e+06u l=220000u
X2529 VSS row_n[8] a_24354_10202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2530 a_26458_2492# col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2531 vcm a_1962_18234# a_10998_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2532 a_24962_11166# a_1962_11206# a_25054_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2533 VDD rowon_n[5] a_12914_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2534 VSS row_n[14] a_23350_16226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2535 a_19430_14540# col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2536 VDD rowon_n[10] a_22954_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2537 a_19030_10162# a_2346_10204# a_18938_10162# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2538 vcm a_1962_9198# a_25054_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2539 a_35094_9158# a_2346_9200# a_35002_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2540 a_20338_2170# col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2541 VDD rowon_n[0] a_10906_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2542 a_27974_18194# a_1962_18234# a_28066_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2543 a_32082_16186# a_2346_16228# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2544 a_22346_8194# rowon_n[6] a_21950_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2545 a_4974_7150# a_2346_7192# a_4882_7150# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2546 VSS row_n[0] a_30378_2170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2547 a_5978_3134# a_2346_3176# a_5886_3134# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2548 VDD VDD a_21950_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2549 VDD rowon_n[15] a_35002_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2550 a_7286_14218# rowon_n[12] a_6890_14178# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2551 a_17326_14218# rowon_n[12] a_16930_14178# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2552 a_10298_8194# col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2553 a_18026_6146# a_2346_6188# a_17934_6146# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2554 vcm a_1962_2170# a_24050_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2555 a_16322_2170# rowon_n[0] a_15926_2130# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2556 a_27062_4138# a_2346_4180# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2557 a_11302_4178# col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2558 analog_in sw_n ctop VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.9e+06u l=220000u
X2559 a_32482_5504# col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2560 a_8898_13174# a_1962_13214# a_8990_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2561 a_18938_13174# a_1962_13214# a_19030_13174# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2562 vcm a_1962_8194# a_14010_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2563 a_34090_12170# a_2346_12212# a_33998_12170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2564 a_3270_10202# col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2565 a_13310_10202# col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2566 a_12002_12170# a_2346_12212# a_11910_12170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2567 a_12306_16226# col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2568 a_35002_12170# row_n[10] a_35494_12532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2569 a_27366_6186# rowon_n[4] a_26970_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2570 a_9994_5142# a_2346_5184# a_9902_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2571 a_3270_3174# col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2572 a_10906_4138# row_n[2] a_11398_4500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2573 a_10998_18194# a_2346_18236# a_10906_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2574 a_33086_18194# a_2346_18236# a_32994_18194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2575 a_5278_9198# rowon_n[7] a_4882_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2576 a_15318_6186# col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2577 a_33998_18194# VDD a_34490_18556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2578 vcm a_1962_14218# a_34090_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2579 a_12402_12532# col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2580 a_19334_12210# rowon_n[10] a_18938_12170# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2581 vcm a_1962_3174# a_6982_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2582 vcm a_1962_7190# a_5978_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2583 a_4882_6146# row_n[4] a_5374_6508# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2584 a_11398_18556# col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2585 vcm a_1962_6186# a_19030_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2586 a_20034_6146# a_2346_6188# a_19942_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2587 a_34490_2492# col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2588 a_2874_1126# VDD a_3366_1488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2589 a_33998_5142# a_1962_5182# a_34090_5142# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2590 VDD rowon_n[8] a_18938_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2591 a_21950_8154# row_n[6] a_22442_8516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2592 VDD rowon_n[7] a_4882_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2593 a_8290_1166# col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2594 a_9902_17190# row_n[15] a_10394_17552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2595 a_21342_15222# rowon_n[13] a_20946_15182# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2596 a_28066_14178# a_2346_14220# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2597 vcm a_1962_13214# a_9994_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2598 a_9902_1126# a_1962_1166# a_9994_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2599 VSS row_n[9] a_22346_11206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2600 a_31382_4178# rowon_n[2] a_30986_4138# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2601 VSS row_n[8] a_35398_10202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2602 a_24354_7190# col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2603 a_12306_10202# rowon_n[8] a_11910_10162# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2604 a_24050_8154# a_2346_8196# a_23958_8154# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2605 a_25054_4138# a_2346_4180# a_24962_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2606 VDD rowon_n[11] a_20946_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2607 a_26970_6146# row_n[4] a_27462_6508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2608 VDD rowon_n[10] a_33998_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2609 VSS row_n[1] a_10298_3174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2610 a_19942_9158# a_1962_9198# a_20034_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2611 a_30074_9158# a_2346_9200# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2612 a_20338_16226# col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2613 VDD rowon_n[2] a_30986_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2614 a_33390_15222# col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2615 a_12402_6508# col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2616 a_16930_14178# a_1962_14218# a_17022_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2617 a_13006_6146# a_2346_6188# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2618 a_29374_5182# col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2619 a_3270_18234# VDD a_2874_18194# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2620 a_13310_18234# VDD a_12914_18194# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2621 VSS row_n[13] a_10298_15222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2622 a_6890_14178# a_1962_14218# a_6982_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2623 a_7286_8194# col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2624 a_29070_6146# a_2346_6188# a_28978_6146# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2625 VSS row_n[12] a_14314_14218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2626 a_11302_11206# col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2627 a_10394_1488# col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2628 a_32482_17552# col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2629 vcm a_1962_15222# a_28066_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2630 VSS row_n[12] a_4274_14218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2631 a_32082_13174# a_2346_13216# a_31990_13174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2632 a_4882_17190# a_1962_17230# a_4974_17190# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2633 a_14922_17190# a_1962_17230# a_15014_17190# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2634 VSS row_n[3] a_14314_5182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2635 VSS VDD a_15318_1166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2636 a_32994_13174# row_n[11] a_33486_13536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2637 a_28978_3134# row_n[1] a_29470_3496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2638 vcm a_1962_5182# a_32082_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2639 VDD rowon_n[14] a_12914_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2640 a_10394_13536# col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2641 vcm a_1962_10202# a_19030_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2642 VDD rowon_n[6] a_17934_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2643 a_29982_8154# row_n[6] a_30474_8516# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2644 a_4370_5504# col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2645 VDD rowon_n[14] a_2874_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2646 a_8898_14178# row_n[12] a_9390_14540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2647 a_18938_14178# row_n[12] a_19430_14540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2648 vcm a_1962_10202# a_8990_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2649 a_4974_5142# a_2346_5184# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2650 a_5978_1126# a_2346_1168# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2651 a_17022_8154# a_2346_8196# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2652 a_18026_4138# a_2346_4180# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2653 VDD sample_n a_1962_3174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2654 vcm a_1962_18234# a_30074_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2655 a_21438_7512# col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2656 a_13918_6146# a_1962_6186# a_14010_6146# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2657 analog_in sw ctop VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.9e+06u l=220000u
X2658 a_14410_3496# col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2659 a_33390_3174# col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2660 VSS row_n[7] a_25358_9198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2661 a_35398_9198# rowon_n[7] a_35002_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2662 a_12002_10162# a_2346_10204# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2663 a_34090_10162# a_2346_10204# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2664 VSS row_n[15] a_28370_17230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2665 a_32386_15222# rowon_n[13] a_31990_15182# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2666 a_1962_10202# sample_n VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2667 a_35002_6146# row_n[4] a_35494_6508# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2668 a_8990_7150# a_2346_7192# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2669 a_9994_3134# a_2346_3176# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2670 a_29374_13214# col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2671 VSS row_n[9] a_33390_11206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2672 a_27974_2130# a_1962_2170# a_28066_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2673 a_24050_18194# a_2346_18236# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2674 a_20946_15182# a_1962_15222# a_21038_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2675 a_5886_5142# a_1962_5182# a_5978_5142# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2676 a_6890_1126# a_1962_1166# a_6982_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2677 a_32994_1126# VDD a_33486_1488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2678 a_15014_17190# a_2346_17232# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2679 a_10298_11206# rowon_n[9] a_9902_11166# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2680 a_25454_9520# col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2681 a_17934_8154# a_1962_8194# a_18026_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2682 a_18938_4138# a_1962_4178# a_19030_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2683 a_26458_5504# col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2684 a_4974_17190# a_2346_17232# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2685 a_24962_14178# a_1962_14218# a_25054_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2686 VDD rowon_n[7] a_35002_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2687 a_8990_16186# a_2346_16228# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2688 a_28466_15544# col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2689 VDD rowon_n[11] a_31990_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2690 a_28066_11166# a_2346_11208# a_27974_11166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2691 a_10998_6146# a_2346_6188# a_10906_6146# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2692 a_20034_4138# a_2346_4180# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2693 a_28978_11166# row_n[9] a_29470_11528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2694 a_9902_11166# a_1962_11206# a_9994_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2695 VDD rowon_n[3] a_10906_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2696 a_3270_4178# rowon_n[2] a_2874_4138# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2697 a_31382_16226# col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2698 VSS row_n[5] a_6282_7190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2699 a_19030_1126# a_2346_1168# a_18938_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2700 vcm a_1962_17230# a_22042_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2701 a_7286_17230# col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2702 a_17326_17230# col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2703 vcm a_1962_16226# a_26058_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2704 a_30074_14178# a_2346_14220# a_29982_14178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2705 a_20338_6186# rowon_n[4] a_19942_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2706 a_2966_5142# a_2346_5184# a_2874_5142# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2707 a_12914_18194# a_1962_18234# a_13006_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2708 a_30474_18556# col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2709 a_15014_8154# a_2346_8196# a_14922_8154# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2710 a_24050_6146# a_2346_6188# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2711 a_16018_4138# a_2346_4180# a_15926_4138# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2712 a_2874_18194# a_1962_18234# a_2966_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2713 a_9994_18194# a_2346_18236# a_9902_18194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2714 a_2346_12212# sample VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2715 a_1962_1166# sample_n VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2716 a_28466_2492# col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2717 vcm a_1962_6186# a_12002_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2718 VDD rowon_n[2] a_2874_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2719 a_16930_15182# row_n[13] a_17422_15544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2720 vcm a_1962_11206# a_17022_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2721 a_6890_15182# row_n[13] a_7382_15544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2722 vcm a_1962_11206# a_6982_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2723 VDD rowon_n[0] a_12914_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2724 VSS row_n[0] a_32386_2170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2725 a_24354_8194# rowon_n[6] a_23958_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2726 a_6982_7150# a_2346_7192# a_6890_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2727 a_7986_3134# a_2346_3176# a_7894_3134# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2728 a_25358_4178# rowon_n[2] a_24962_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2729 VSS row_n[10] a_27366_12210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2730 vcm a_1962_2170# a_26058_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2731 a_29070_4138# a_2346_4180# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2732 a_13310_4178# col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2733 a_32082_11166# a_2346_11208# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2734 a_31382_10202# rowon_n[8] a_30986_10162# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2735 vcm a_1962_5182# a_3970_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2736 a_34490_5504# col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2737 vcm a_1962_8194# a_16018_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2738 vcm a_1962_4178# a_17022_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2739 VSS VDD a_26362_18234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2740 a_30378_16226# rowon_n[14] a_29982_16186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2741 VDD rowon_n[12] a_25966_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2742 a_14010_12170# a_2346_12212# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2743 a_30986_7150# a_1962_7190# a_31078_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2744 a_31990_3134# a_1962_3174# a_32082_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2745 a_27366_14218# col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2746 a_3970_12170# a_2346_12212# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2747 VDD rowon_n[2] a_24962_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2748 a_35094_18194# a_2346_18236# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2749 a_31990_15182# a_1962_15222# a_32082_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2750 a_27462_10524# col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2751 VSS row_n[4] a_19334_6186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2752 a_12914_4138# row_n[2] a_13406_4500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2753 a_2966_18194# a_2346_18236# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2754 a_13006_18194# a_2346_18236# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2755 a_29374_6186# rowon_n[4] a_28978_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2756 a_5278_3174# col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2757 a_25358_17230# col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2758 a_26458_16548# col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2759 a_7286_9198# rowon_n[7] a_6890_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2760 vcm a_1962_7190# a_7986_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2761 vcm a_1962_3174# a_8990_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2762 a_30378_11206# col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2763 ctop sw analog_in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.9e+06u l=220000u
X2764 a_22346_5182# col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2765 VSS row_n[13] a_9294_15222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2766 a_24050_15182# a_2346_15224# a_23958_15182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2767 a_6282_12210# col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2768 a_16322_12210# col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2769 vcm a_1962_12210# a_21038_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2770 a_22042_6146# a_2346_6188# a_21950_6146# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2771 a_4882_1126# VDD a_5374_1488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2772 vcm a_1962_11206# a_25054_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2773 a_23958_8154# row_n[6] a_24450_8516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2774 a_24962_15182# row_n[13] a_25454_15544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2775 a_8990_13174# a_2346_13216# a_8898_13174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2776 VDD rowon_n[7] a_6890_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2777 VDD rowon_n[15] a_7894_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2778 a_5374_14540# col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2779 a_15414_14540# col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2780 VSS sample_n a_1962_8194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2781 a_21950_3134# row_n[1] a_22442_3496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2782 a_9390_13536# col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2783 a_5886_10162# row_n[8] a_6378_10524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2784 a_15926_10162# row_n[8] a_16418_10524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2785 a_26362_7190# col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2786 a_27366_3174# col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2787 a_33390_4178# rowon_n[2] a_32994_4138# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2788 a_10998_4138# a_2346_4180# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2789 a_17326_9198# col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2790 a_27062_4138# a_2346_4180# a_26970_4138# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2791 a_28978_6146# row_n[4] a_29470_6508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2792 a_24354_17230# rowon_n[15] a_23958_17190# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2793 vcm a_1962_15222# a_13006_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2794 VSS row_n[1] a_12306_3174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2795 vcm a_1962_15222# a_2966_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2796 a_32082_9158# a_2346_9200# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2797 a_26970_1126# VDD a_27462_1488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2798 a_28370_16226# rowon_n[14] a_27974_16186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2799 VSS row_n[11] a_25358_13214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2800 a_22346_10202# col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2801 a_2966_3134# a_2346_3176# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2802 VDD rowon_n[2] a_32994_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2803 a_1962_7190# sample_n VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2804 a_14410_6508# col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2805 a_20946_2130# a_1962_2170# a_21038_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2806 a_15318_12210# rowon_n[10] a_14922_12170# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2807 a_16930_9158# row_n[7] a_17422_9520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2808 a_9294_8194# col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2809 a_2346_6188# sample VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2810 a_15014_6146# a_2346_6188# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2811 a_31078_2130# a_2346_2172# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2812 a_5278_12210# rowon_n[10] a_4882_12170# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2813 VSS sample_n a_1962_15222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2814 VDD rowon_n[13] a_23958_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2815 a_12002_13174# a_2346_13216# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2816 a_34090_13174# a_2346_13216# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2817 a_21438_12532# col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2818 a_10906_8154# a_1962_8194# a_10998_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2819 a_18330_5182# rowon_n[3] a_17934_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2820 a_12402_1488# col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2821 a_19334_1166# en_bit_n[2] a_18938_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2822 a_31382_1166# col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2823 a_11910_4138# a_1962_4178# a_12002_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2824 a_1962_13214# sample_n VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2825 a_9294_11206# rowon_n[9] a_8898_11166# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2826 VSS row_n[0] a_4274_2170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2827 a_30378_5182# col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2828 a_25454_11528# col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2829 VSS VDD a_17326_1166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2830 a_23350_18234# col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2831 vcm a_1962_5182# a_34090_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2832 VDD rowon_n[8] a_14922_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2833 a_7986_1126# a_2346_1168# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2834 VDD rowon_n[8] a_4882_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2835 a_6982_5142# a_2346_5184# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2836 VSS row_n[15] a_3270_17230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2837 VSS row_n[15] a_13310_17230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2838 a_29982_3134# row_n[1] a_30474_3496# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2839 VDD rowon_n[1] a_17934_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2840 VSS row_n[14] a_17326_16226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2841 a_22042_16186# a_2346_16228# a_21950_16186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2842 a_14314_13214# col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2843 a_2874_7150# a_1962_7190# a_2966_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2844 vcm a_1962_1166# a_9994_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2845 a_3878_3134# a_1962_3174# a_3970_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2846 VSS row_n[14] a_7286_16226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2847 a_13006_15182# a_2346_15224# a_12914_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2848 a_35094_15182# a_2346_15224# a_35002_15182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2849 a_4274_13214# col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2850 vcm a_1962_12210# a_32082_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2851 a_23446_7512# col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2852 a_15926_6146# a_1962_6186# a_16018_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2853 a_22954_16186# row_n[14] a_23446_16548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2854 a_2966_15182# a_2346_15224# a_2874_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2855 VSS row_n[7] a_27366_9198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2856 VSS sample a_2346_2172# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2857 a_35398_3174# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2858 a_9902_14178# a_1962_14218# a_9994_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2859 a_17022_14178# a_2346_14220# a_16930_14178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2860 a_21438_2492# col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2861 VDD VDD a_15926_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2862 a_13406_15544# col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2863 a_6982_14178# a_2346_14220# a_6890_14178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2864 VDD VDD a_5886_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2865 a_3366_15544# col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2866 VSS row_n[0] a_26362_2170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2867 a_13918_11166# row_n[9] a_14410_11528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2868 a_3878_11166# row_n[9] a_4370_11528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2869 vcm a_1962_9198# a_20034_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2870 a_35002_1126# VDD a_35494_1488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2871 a_26058_12170# a_2346_12212# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2872 a_30074_9158# a_2346_9200# a_29982_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2873 VSS row_n[6] a_16322_8194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2874 a_7894_5142# a_1962_5182# a_7986_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2875 a_8898_1126# a_1962_1166# a_8990_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2876 a_27462_9520# col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2877 a_28466_5504# col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2878 a_23350_12210# rowon_n[10] a_22954_12170# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2879 a_20946_10162# a_1962_10202# a_21038_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2880 a_6378_8516# col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2881 a_13006_6146# a_2346_6188# a_12914_6146# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2882 a_11302_2170# rowon_n[0] a_10906_2130# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2883 a_22042_4138# a_2346_4180# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2884 a_22346_18234# VDD a_21950_18194# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2885 vcm a_1962_16226# a_10998_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2886 a_35398_17230# rowon_n[15] a_35002_17190# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2887 VDD rowon_n[3] a_12914_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2888 VSS row_n[12] a_23350_14218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2889 a_8990_11166# a_2346_11208# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2890 a_23958_17190# a_1962_17230# a_24050_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2891 a_19430_12532# col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2892 VDD rowon_n[8] a_22954_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2893 VSS row_n[5] a_8290_7190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2894 a_27974_16186# a_1962_16226# a_28066_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2895 a_32082_14178# a_2346_14220# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2896 a_22346_6186# rowon_n[4] a_21950_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2897 a_4974_5142# a_2346_5184# a_4882_5142# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2898 a_5978_1126# a_2346_1168# a_5886_1126# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2899 VDD rowon_n[14] a_21950_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2900 VDD rowon_n[13] a_35002_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2901 a_10298_6186# col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2902 a_18026_4138# a_2346_4180# a_17934_4138# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2903 a_35398_12210# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2904 a_17022_8154# a_2346_8196# a_16930_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2905 VSS row_n[10] a_12306_12210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2906 vcm a_1962_6186# a_14010_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2907 a_34394_18234# col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2908 VSS VDD a_11302_18234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2909 a_34490_14540# col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2910 a_34090_10162# a_2346_10204# a_33998_10162# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2911 a_12002_10162# a_2346_10204# a_11910_10162# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2912 vcm a_1962_18234# a_29070_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2913 VDD rowon_n[12] a_10906_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2914 a_12306_14218# col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2915 a_35002_10162# row_n[8] a_35494_10524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2916 VSS row_n[0] a_34394_2170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2917 a_3270_1166# col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2918 a_9994_3134# a_2346_3176# a_9902_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2919 a_27366_4178# rowon_n[2] a_26970_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2920 a_10998_16186# a_2346_16228# a_10906_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2921 a_33086_16186# a_2346_16228# a_32994_16186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2922 a_19334_10202# rowon_n[8] a_18938_10162# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2923 a_26362_8194# rowon_n[6] a_25966_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2924 a_8990_7150# a_2346_7192# a_8898_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2925 vcm a_1962_2170# a_28066_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2926 a_15318_4178# col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2927 a_33998_16186# row_n[14] a_34490_16548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2928 a_12402_10524# col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2929 vcm a_1962_1166# a_6982_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2930 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X2931 a_10298_17230# col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2932 vcm a_1962_5182# a_5978_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2933 a_11398_16548# col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2934 vcm a_1962_8194# a_18026_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2935 vcm a_1962_4178# a_19030_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2936 a_20034_4138# a_2346_4180# a_19942_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2937 a_26058_9158# a_2346_9200# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2938 a_15318_7190# rowon_n[5] a_14922_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2939 a_32994_7150# a_1962_7190# a_33086_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2940 a_33998_3134# a_1962_3174# a_34090_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2941 a_21950_6146# row_n[4] a_22442_6508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2942 VDD rowon_n[2] a_26970_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2943 VDD rowon_n[5] a_4882_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2944 a_14922_4138# row_n[2] a_15414_4500# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2945 a_9902_15182# row_n[13] a_10394_15544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2946 a_21342_13214# rowon_n[11] a_20946_13174# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2947 vcm a_1962_11206# a_9994_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2948 a_34394_12210# rowon_n[10] a_33998_12170# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2949 a_31990_10162# a_1962_10202# a_32082_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2950 a_9294_9198# rowon_n[7] a_8898_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2951 a_1962_18234# sample_n VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2952 a_22954_12170# a_1962_12210# a_23046_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2953 a_24354_5182# col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2954 a_24050_6146# a_2346_6188# a_23958_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2955 a_21950_18194# a_1962_18234# a_22042_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2956 VDD rowon_n[9] a_20946_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2957 VDD rowon_n[8] a_33998_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2958 a_25966_8154# row_n[6] a_26458_8516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2959 VDD rowon_n[7] a_8898_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2960 VSS VDD a_10298_1166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2961 VSS row_n[15] a_32386_17230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2962 a_23958_3134# row_n[1] a_24450_3496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2963 a_20338_14218# col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2964 a_33390_13214# col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2965 a_12002_8154# a_2346_8196# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2966 a_28370_7190# col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2967 a_29374_3174# col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2968 a_13006_4138# a_2346_4180# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2969 a_27062_17190# a_2346_17232# a_26970_17190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2970 a_3270_16226# rowon_n[14] a_2874_16186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2971 a_13310_16226# rowon_n[14] a_12914_16186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2972 VSS row_n[11] a_10298_13214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2973 a_7286_6186# col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2974 a_29070_4138# a_2346_4180# a_28978_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2975 a_19334_9198# col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2976 a_27974_17190# row_n[15] a_28466_17552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2977 a_32482_15544# col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2978 vcm a_1962_13214# a_28066_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2979 a_32082_11166# a_2346_11208# a_31990_11166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2980 a_4882_15182# a_1962_15222# a_4974_15182# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2981 a_14922_15182# a_1962_15222# a_15014_15182# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2982 VSS row_n[7] a_20338_9198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2983 a_30378_9198# rowon_n[7] a_29982_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2984 VSS row_n[1] a_14314_3174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2985 a_32994_11166# row_n[9] a_33486_11528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2986 a_28978_1126# VDD a_29470_1488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2987 vcm a_1962_3174# a_32082_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2988 a_10394_11528# col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2989 a_34090_9158# a_2346_9200# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2990 vcm a_1962_7190# a_31078_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2991 VDD rowon_n[4] a_17934_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2992 a_29982_6146# row_n[4] a_30474_6508# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2993 a_8898_12170# row_n[10] a_9390_12532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2994 a_18938_12170# row_n[10] a_19430_12532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2995 a_3970_7150# a_2346_7192# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2996 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X2997 a_4974_3134# a_2346_3176# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2998 a_17022_6146# a_2346_6188# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2999 a_22954_2130# a_1962_2170# a_23046_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3000 a_18938_9158# row_n[7] a_19430_9520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3001 VDD sample_n a_1962_1166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3002 a_33086_2130# a_2346_2172# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3003 vcm a_1962_16226# a_30074_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3004 a_20434_9520# col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3005 a_12914_8154# a_1962_8194# a_13006_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3006 a_14410_1488# col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3007 a_13918_4138# a_1962_4178# a_14010_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3008 a_21438_5504# col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3009 VSS sample a_2346_14220# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3010 VDD rowon_n[7] a_29982_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3011 a_33390_1166# col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3012 vcm a_1962_17230# a_16018_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3013 vcm a_1962_17230# a_5978_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3014 VSS row_n[13] a_28370_15222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3015 a_32386_13214# rowon_n[11] a_31990_13174# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3016 a_20034_17190# a_2346_17232# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3017 a_8990_5142# a_2346_5184# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3018 a_9994_1126# a_2346_1168# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3019 a_29374_11206# col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3020 a_24050_16186# a_2346_16228# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3021 a_20946_13174# a_1962_13214# a_21038_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3022 a_4882_7150# a_1962_7190# a_4974_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3023 a_5886_3134# a_1962_3174# a_5978_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3024 VDD rowon_n[15] a_26970_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3025 a_15014_15182# a_2346_15224# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3026 a_33998_12170# a_1962_12210# a_34090_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3027 a_25454_7512# col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3028 a_17934_6146# a_1962_6186# a_18026_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3029 a_4974_15182# a_2346_15224# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3030 VDD rowon_n[5] a_35002_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3031 a_8990_14178# a_2346_14220# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3032 a_28466_13536# col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3033 VDD rowon_n[9] a_31990_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3034 VSS row_n[7] a_29374_9198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3035 a_10998_4138# a_2346_4180# a_10906_4138# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3036 a_23446_2492# col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3037 VSS VDD a_30378_18234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3038 VSS row_n[0] a_28370_2170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3039 a_31382_14218# col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3040 a_32386_8194# col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3041 VSS row_n[3] a_6282_5182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3042 a_25054_18194# a_2346_18236# a_24962_18194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3043 vcm a_1962_15222# a_22042_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3044 a_32082_9158# a_2346_9200# a_31990_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3045 VSS row_n[6] a_18330_8194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3046 a_16018_17190# a_2346_17232# a_15926_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3047 a_7286_15222# col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3048 a_17326_15222# col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3049 a_29470_9520# col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3050 a_25966_18194# VDD a_26458_18556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3051 a_5978_17190# a_2346_17232# a_5886_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3052 vcm a_1962_14218# a_26058_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3053 a_8386_8516# col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3054 a_2966_3134# a_2346_3176# a_2874_3134# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3055 a_20338_4178# rowon_n[2] a_19942_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3056 a_12914_16186# a_1962_16226# a_13006_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3057 a_30474_16548# col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3058 a_15014_6146# a_2346_6188# a_14922_6146# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3059 vcm a_1962_2170# a_21038_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3060 a_13310_2170# rowon_n[0] a_12914_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3061 a_24050_4138# a_2346_4180# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3062 a_2874_16186# a_1962_16226# a_2966_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3063 a_9994_16186# a_2346_16228# a_9902_16186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3064 a_2346_10204# sample VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3065 a_26970_7150# a_1962_7190# a_27062_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3066 a_31078_2130# a_2346_2172# a_30986_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3067 a_6378_17552# col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3068 a_16418_17552# col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3069 vcm a_1962_8194# a_10998_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3070 a_6378_3496# col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3071 vcm a_1962_4178# a_12002_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3072 a_16930_13174# row_n[11] a_17422_13536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3073 a_6890_13174# row_n[11] a_7382_13536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3074 VDD rowon_n[2] a_19942_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3075 vcm a_1962_12210# a_15014_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3076 vcm a_1962_12210# a_4974_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3077 a_24354_6186# rowon_n[4] a_23958_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3078 a_6982_5142# a_2346_5184# a_6890_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3079 a_7986_1126# a_2346_1168# a_7894_1126# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3080 VSS row_n[8] a_27366_10202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3081 vcm a_1962_18234# a_3970_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3082 vcm a_1962_18234# a_14010_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3083 a_27974_11166# a_1962_11206# a_28066_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3084 vcm a_1962_7190# a_2966_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3085 vcm a_1962_3174# a_3970_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3086 vcm a_1962_6186# a_16018_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3087 VSS row_n[14] a_26362_16226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3088 a_30378_14218# rowon_n[12] a_29982_14178# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3089 VDD rowon_n[10] a_25966_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3090 a_31990_1126# a_1962_1166# a_32082_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3091 a_30986_5142# a_1962_5182# a_31078_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3092 a_31078_17190# a_2346_17232# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3093 a_35094_16186# a_2346_16228# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3094 a_31990_13174# a_1962_13214# a_32082_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3095 a_5278_1166# col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3096 VSS row_n[2] a_19334_4178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3097 VDD VDD a_24962_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3098 a_2966_16186# a_2346_16228# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3099 a_13006_16186# a_2346_16228# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3100 a_28370_8194# rowon_n[6] a_27974_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3101 a_29374_4178# rowon_n[2] a_28978_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3102 a_25358_15222# col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3103 VDD rowon_n[6] a_14922_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3104 vcm a_1962_5182# a_7986_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3105 vcm a_1962_1166# a_8990_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3106 a_21342_7190# col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3107 a_22346_3174# col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3108 a_8290_17230# rowon_n[15] a_7894_17190# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3109 VSS row_n[5] a_31382_7190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3110 ctop sw_n ctop VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.9e+06u l=220000u
X3111 a_24450_17552# col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3112 a_20946_14178# row_n[12] a_21438_14540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3113 VSS row_n[11] a_9294_13214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3114 a_24050_13174# a_2346_13216# a_23958_13174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3115 a_6282_10202# col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3116 a_16322_10202# col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3117 vcm a_1962_10202# a_21038_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3118 a_12306_9198# col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3119 a_35002_7150# a_1962_7190# a_35094_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3120 a_22042_4138# a_2346_4180# a_21950_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3121 a_4974_12170# a_2346_12212# a_4882_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3122 a_15014_12170# a_2346_12212# a_14922_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3123 a_28066_9158# a_2346_9200# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3124 a_17326_7190# rowon_n[5] a_16930_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3125 a_23958_6146# row_n[4] a_24450_6508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3126 VDD rowon_n[2] a_28978_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3127 a_19430_4500# col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3128 a_24962_13174# row_n[11] a_25454_13536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3129 a_8990_11166# a_2346_11208# a_8898_11166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3130 VDD rowon_n[5] a_6890_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3131 VDD rowon_n[13] a_7894_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3132 a_5374_12532# col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3133 a_15414_12532# col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3134 VSS sample_n a_1962_6186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3135 a_21950_1126# VDD a_22442_1488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3136 VDD rowon_n[0] a_4882_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3137 a_9390_11528# col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3138 a_27366_1166# col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3139 a_26362_5182# col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3140 a_11910_9158# row_n[7] a_12402_9520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3141 a_4274_8194# col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3142 vcm a_1962_17230# a_35094_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3143 a_27974_8154# row_n[6] a_28466_8516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3144 a_12914_17190# row_n[15] a_13406_17552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3145 a_24354_15222# rowon_n[13] a_23958_15182# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3146 vcm a_1962_13214# a_13006_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3147 VSS row_n[10] a_21342_12210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3148 VSS VDD a_12306_1166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3149 a_2874_17190# row_n[15] a_3366_17552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3150 vcm a_1962_13214# a_2966_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3151 a_25966_3134# row_n[1] a_26458_3496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3152 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.64e+07u l=1.6e+07u
X3153 a_28370_14218# rowon_n[12] a_27974_14178# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3154 VSS row_n[9] a_25358_11206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3155 a_1962_5182# sample_n VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3156 a_2966_1126# a_2346_1168# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3157 a_15014_4138# a_2346_4180# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3158 a_29070_17190# a_2346_17232# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3159 VDD rowon_n[12] a_19942_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3160 a_30074_12170# a_2346_12212# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3161 a_15318_10202# rowon_n[8] a_14922_10162# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3162 a_14010_8154# a_2346_8196# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3163 a_16930_7150# row_n[5] a_17422_7512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3164 a_9294_6186# col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3165 a_5278_10202# rowon_n[8] a_4882_10162# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3166 VSS sample_n a_1962_13214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3167 VDD rowon_n[11] a_23958_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3168 a_21438_10524# col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3169 a_10906_6146# a_1962_6186# a_10998_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3170 a_18330_3174# rowon_n[1] a_17934_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3171 VSS row_n[7] a_22346_9198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3172 a_30378_3174# col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3173 a_32386_9198# rowon_n[7] a_31990_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3174 a_23350_16226# col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3175 vcm a_1962_7190# a_33086_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3176 vcm a_1962_3174# a_34090_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3177 a_14922_10162# a_1962_10202# a_15014_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3178 a_26058_9158# a_2346_9200# a_25966_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3179 VSS row_n[0] a_21342_2170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3180 a_6982_3134# a_2346_3176# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3181 a_4882_10162# a_1962_10202# a_4974_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3182 a_6282_18234# VDD a_5886_18194# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3183 a_16322_18234# VDD a_15926_18194# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3184 VSS row_n[13] a_3270_15222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3185 VSS row_n[13] a_13310_15222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3186 a_35094_2130# a_2346_2172# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3187 a_3878_1126# a_1962_1166# a_3970_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3188 VDD en_bit_n[1] a_17934_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3189 a_29982_1126# VDD a_30474_1488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3190 a_24962_2130# a_1962_2170# a_25054_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3191 a_22442_18556# col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3192 VSS row_n[12] a_17326_14218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3193 a_22042_14178# a_2346_14220# a_21950_14178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3194 a_14314_11206# col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3195 VSS row_n[6] a_11302_8194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3196 a_2874_5142# a_1962_5182# a_2966_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3197 a_35494_17552# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3198 VSS row_n[12] a_7286_14218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3199 a_31990_14178# row_n[12] a_32482_14540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3200 a_13006_13174# a_2346_13216# a_12914_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3201 a_35094_13174# a_2346_13216# a_35002_13174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3202 a_4274_11206# col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3203 vcm a_1962_10202# a_32082_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3204 a_22442_9520# col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3205 a_14922_8154# a_1962_8194# a_15014_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3206 a_35398_1166# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3207 a_15926_4138# a_1962_4178# a_16018_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3208 a_23446_5504# col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3209 a_17934_17190# a_1962_17230# a_18026_17190# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3210 a_2966_13174# a_2346_13216# a_2874_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3211 VDD rowon_n[7] a_31990_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3212 a_7894_17190# a_1962_17230# a_7986_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3213 VDD rowon_n[15] a_11910_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3214 VDD rowon_n[14] a_15926_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3215 a_13406_13536# col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3216 VDD rowon_n[14] a_5886_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3217 a_3366_13536# col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3218 VSS row_n[5] a_3270_7190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3219 vcm a_1962_18234# a_33086_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3220 VSS row_n[4] a_16322_6186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3221 a_7894_3134# a_1962_3174# a_7986_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3222 VSS row_n[10] a_19334_12210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3223 a_27462_7512# col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3224 a_24050_11166# a_2346_11208# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3225 a_23350_10202# rowon_n[8] a_22954_10162# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3226 a_6378_6508# col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3227 a_13006_4138# a_2346_4180# a_12914_4138# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3228 a_15014_10162# a_2346_10204# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3229 a_12002_8154# a_2346_8196# a_11910_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3230 a_25454_2492# col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3231 a_10906_18194# VDD a_11398_18556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3232 a_22346_16226# rowon_n[14] a_21950_16186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3233 a_35398_15222# rowon_n[13] a_35002_15182# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3234 vcm a_1962_14218# a_10998_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3235 a_4974_10162# a_2346_10204# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3236 VDD rowon_n[0] a_35002_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3237 VDD rowon_n[12] a_17934_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3238 a_34394_8194# col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3239 a_27062_18194# a_2346_18236# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3240 a_23958_15182# a_1962_15222# a_24050_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3241 a_19430_10524# col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3242 VSS row_n[3] a_8290_5182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3243 a_18026_17190# a_2346_17232# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3244 a_34090_9158# a_2346_9200# a_33998_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3245 a_7986_17190# a_2346_17232# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3246 a_27974_14178# a_1962_14218# a_28066_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3247 a_21342_8194# rowon_n[6] a_20946_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3248 a_4974_3134# a_2346_3176# a_4882_3134# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3249 a_22346_4178# rowon_n[2] a_21950_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3250 VDD rowon_n[11] a_35002_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3251 a_3970_7150# a_2346_7192# a_3878_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3252 vcm a_1962_2170# a_23046_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3253 a_10298_4178# col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3254 a_35398_10202# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3255 a_17022_6146# a_2346_6188# a_16930_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3256 a_33086_2130# a_2346_2172# a_32994_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3257 a_28978_7150# a_1962_7190# a_29070_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3258 a_8386_3496# col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3259 VSS row_n[8] a_12306_10202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3260 vcm a_1962_8194# a_13006_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3261 vcm a_1962_4178# a_14010_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3262 a_34394_16226# col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3263 a_2874_11166# a_1962_11206# a_2966_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3264 a_12914_11166# a_1962_11206# a_13006_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3265 VSS row_n[14] a_11302_16226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3266 a_34490_12532# col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3267 a_21038_9158# a_2346_9200# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3268 a_10298_7190# rowon_n[5] a_9902_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3269 VDD rowon_n[2] a_21950_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3270 vcm a_1962_16226# a_29070_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3271 a_33086_14178# a_2346_14220# a_32994_14178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3272 VDD rowon_n[10] a_10906_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3273 a_26362_6186# rowon_n[4] a_25966_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3274 a_9994_1126# a_2346_1168# a_9902_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3275 a_9902_4138# row_n[2] a_10394_4500# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3276 a_33486_18556# col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3277 a_10998_14178# a_2346_14220# a_10906_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3278 a_8990_5142# a_2346_5184# a_8898_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3279 a_5886_18194# a_1962_18234# a_5978_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3280 VDD VDD a_9902_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3281 a_15926_18194# a_1962_18234# a_16018_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3282 a_4274_9198# rowon_n[7] a_3878_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3283 a_10298_15222# col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3284 vcm a_1962_7190# a_4974_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3285 vcm a_1962_3174# a_5978_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3286 vcm a_1962_6186# a_18026_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3287 a_15318_5182# rowon_n[3] a_14922_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3288 a_32994_5142# a_1962_5182# a_33086_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3289 a_20946_8154# row_n[6] a_21438_8516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3290 VDD rowon_n[7] a_3878_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3291 a_31478_8516# col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3292 VDD rowon_n[3] a_4882_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3293 a_9902_13174# row_n[11] a_10394_13536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3294 a_21342_11206# rowon_n[9] a_20946_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3295 VDD rowon_n[6] a_16930_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3296 a_35094_11166# a_2346_11208# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3297 a_34394_10202# rowon_n[8] a_33998_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3298 a_2966_11166# a_2346_11208# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3299 a_13006_11166# a_2346_11208# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3300 a_1962_16226# sample_n VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3301 a_23350_7190# col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3302 a_24354_3174# col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3303 VDD rowon_n[1] a_14922_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3304 VDD rowon_n[12] a_28978_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3305 a_17022_12170# a_2346_12212# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3306 VSS row_n[5] a_33390_7190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3307 a_24050_4138# a_2346_4180# a_23958_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3308 a_6982_12170# a_2346_12212# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3309 a_14314_9198# col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3310 vcm a_1962_7190# a_27062_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3311 a_21950_16186# a_1962_16226# a_22042_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3312 a_25966_6146# row_n[4] a_26458_6508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3313 a_5978_18194# a_2346_18236# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3314 a_16018_18194# a_2346_18236# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3315 VDD rowon_n[5] a_8898_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3316 a_28370_17230# col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3317 VSS row_n[13] a_32386_15222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3318 a_23958_1126# VDD a_24450_1488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3319 a_33390_11206# col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3320 VDD rowon_n[0] a_6890_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3321 a_13310_14218# rowon_n[12] a_12914_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3322 a_12002_6146# a_2346_6188# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3323 a_29374_1166# col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3324 a_28370_5182# col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3325 VDD rowon_n[15] a_30986_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3326 a_27062_15182# a_2346_15224# a_26970_15182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3327 a_3270_14218# rowon_n[12] a_2874_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3328 a_9294_12210# col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3329 a_19334_12210# col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3330 vcm a_1962_12210# a_24050_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3331 VSS row_n[9] a_10298_11206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3332 a_13918_9158# row_n[7] a_14410_9520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3333 a_6282_8194# col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3334 a_7286_4178# col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3335 vcm a_1962_11206# a_28066_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3336 a_27974_15182# row_n[13] a_28466_15544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3337 a_32482_13536# col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3338 a_4882_13174# a_1962_13214# a_4974_13174# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3339 a_14922_13174# a_1962_13214# a_15014_13174# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3340 VSS VDD a_14314_1166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3341 a_8386_14540# col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3342 a_18426_14540# col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3343 vcm a_1962_1166# a_32082_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3344 a_27974_3134# row_n[1] a_28466_3496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3345 vcm a_1962_5182# a_31078_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3346 a_8898_10162# row_n[8] a_9390_10524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3347 a_18938_10162# row_n[8] a_19430_10524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3348 a_3970_5142# a_2346_5184# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3349 a_4974_1126# a_2346_1168# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3350 a_6890_4138# row_n[2] a_7382_4500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3351 a_17022_4138# a_2346_4180# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3352 a_18938_7150# row_n[5] a_19430_7512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3353 a_29982_18194# VDD a_30474_18556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3354 vcm a_1962_14218# a_30074_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3355 a_20434_7512# col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3356 a_12914_6146# a_1962_6186# a_13006_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3357 VSS sample a_2346_12212# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3358 VDD rowon_n[5] a_29982_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3359 a_16930_2130# row_n[0] a_17422_2492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3360 a_27366_17230# rowon_n[15] a_26970_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3361 vcm a_1962_15222# a_16018_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3362 VSS row_n[7] a_24354_9198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3363 vcm a_1962_15222# a_5978_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3364 a_34394_9198# rowon_n[7] a_33998_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3365 VSS row_n[11] a_28370_13214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3366 a_32386_11206# rowon_n[9] a_31990_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3367 a_28066_9158# a_2346_9200# a_27974_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3368 vcm a_1962_7190# a_35094_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3369 a_20034_15182# a_2346_15224# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3370 VSS row_n[0] a_23350_2170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3371 a_8990_3134# a_2346_3176# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3372 a_24050_14178# a_2346_14220# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3373 VSS row_n[6] a_13310_8194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3374 a_19030_8154# a_2346_8196# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3375 a_4882_5142# a_1962_5182# a_4974_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3376 a_5886_1126# a_1962_1166# a_5978_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3377 VDD rowon_n[13] a_26970_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3378 a_15014_13174# a_2346_13216# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3379 a_24450_9520# col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3380 a_17934_4138# a_1962_4178# a_18026_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3381 a_25454_5504# col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3382 a_4974_13174# a_2346_13216# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3383 VDD rowon_n[7] a_33998_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3384 a_3366_8516# col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3385 VDD rowon_n[3] a_35002_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3386 a_28466_11528# col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3387 a_21950_7150# a_1962_7190# a_22042_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3388 a_26362_18234# col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3389 VSS row_n[14] a_30378_16226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3390 VSS row_n[15] a_6282_17230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3391 VSS row_n[15] a_16322_17230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3392 a_21038_17190# a_2346_17232# a_20946_17190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3393 VSS row_n[5] a_5278_7190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3394 a_32386_6186# col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3395 VSS row_n[1] a_6282_3174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3396 a_35002_18194# a_1962_18234# a_35094_18194# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X3397 a_25054_16186# a_2346_16228# a_24962_16186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3398 a_17326_13214# col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3399 vcm a_1962_13214# a_22042_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3400 VSS row_n[4] a_18330_6186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3401 a_21950_17190# row_n[15] a_22442_17552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3402 a_16018_15182# a_2346_15224# a_15926_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3403 a_7286_13214# col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3404 a_29470_7512# col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3405 a_25966_16186# row_n[14] a_26458_16548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3406 a_5978_15182# a_2346_15224# a_5886_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3407 a_8386_6508# col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3408 a_2966_1126# a_2346_1168# a_2874_1126# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3409 a_12914_14178# a_1962_14218# a_13006_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3410 a_14010_8154# a_2346_8196# a_13918_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3411 a_15014_4138# a_2346_4180# a_14922_4138# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3412 a_16418_15544# col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3413 a_2874_14178# a_1962_14218# a_2966_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3414 a_9994_14178# a_2346_14220# a_9902_14178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3415 a_27462_2492# col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3416 a_26970_5142# a_1962_5182# a_27062_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3417 VDD VDD a_8898_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3418 a_6378_15544# col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3419 vcm a_1962_6186# a_10998_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3420 a_6378_1488# col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3421 a_16930_11166# row_n[9] a_17422_11528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3422 a_6890_11166# row_n[9] a_7382_11528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3423 vcm a_1962_10202# a_15014_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3424 a_4882_14178# row_n[12] a_5374_14540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3425 a_14922_14178# row_n[12] a_15414_14540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3426 a_26362_12210# rowon_n[10] a_25966_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3427 vcm a_1962_10202# a_4974_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3428 a_23958_10162# a_1962_10202# a_24050_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3429 a_23350_8194# rowon_n[6] a_22954_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3430 a_6982_3134# a_2346_3176# a_6890_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3431 a_24354_4178# rowon_n[2] a_23958_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3432 VDD rowon_n[6] a_9902_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3433 vcm a_1962_2170# a_25054_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3434 a_25358_18234# VDD a_24962_18194# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3435 vcm a_1962_16226# a_3970_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3436 vcm a_1962_16226# a_14010_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3437 vcm a_1962_5182# a_2966_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3438 a_35094_2130# a_2346_2172# a_35002_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3439 vcm a_1962_1166# a_3970_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3440 vcm a_1962_8194# a_15014_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3441 vcm a_1962_4178# a_16018_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3442 VSS row_n[12] a_26362_14218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3443 a_26970_17190# a_1962_17230# a_27062_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3444 VDD rowon_n[8] a_25966_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3445 a_29982_7150# a_1962_7190# a_30074_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3446 a_30986_3134# a_1962_3174# a_31078_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3447 a_31078_15182# a_2346_15224# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3448 a_23046_9158# a_2346_9200# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3449 a_12306_7190# rowon_n[5] a_11910_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3450 VDD rowon_n[2] a_23958_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3451 VSS row_n[15] a_24354_17230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3452 a_35094_14178# a_2346_14220# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3453 VDD rowon_n[14] a_24962_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3454 a_2966_14178# a_2346_14220# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3455 a_13006_14178# a_2346_14220# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3456 a_28370_6186# rowon_n[4] a_27974_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3457 a_25358_13214# col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3458 a_6282_9198# rowon_n[7] a_5886_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3459 VDD rowon_n[4] a_14922_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3460 vcm a_1962_3174# a_7986_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3461 a_19030_17190# a_2346_17232# a_18938_17190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3462 VSS row_n[10] a_15318_12210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3463 a_20034_12170# a_2346_12212# a_19942_12170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3464 a_22346_1166# col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3465 a_21342_5182# col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3466 a_8290_15222# rowon_n[13] a_7894_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3467 VSS row_n[10] a_5278_12210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3468 a_5278_2170# rowon_n[0] a_4882_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3469 VSS row_n[3] a_31382_5182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3470 a_24450_15544# col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3471 a_20946_12170# row_n[10] a_21438_12532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3472 VSS row_n[9] a_9294_11206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3473 a_24050_11166# a_2346_11208# a_23958_11166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3474 ctop sw_n ctop VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.9e+06u l=220000u
X3475 a_35002_5142# a_1962_5182# a_35094_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3476 a_4974_10162# a_2346_10204# a_4882_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3477 a_15014_10162# a_2346_10204# a_14922_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3478 a_22954_8154# row_n[6] a_23446_8516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3479 a_17326_5182# rowon_n[3] a_16930_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3480 VDD rowon_n[12] a_13918_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3481 a_24962_11166# row_n[9] a_25454_11528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3482 a_33486_8516# col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3483 VDD rowon_n[12] a_3878_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3484 VDD rowon_n[7] a_5886_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3485 VDD rowon_n[3] a_6890_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3486 VDD rowon_n[11] a_7894_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3487 a_5374_10524# col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3488 a_15414_10524# col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3489 a_20946_3134# row_n[1] a_21438_3496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3490 VSS sample_n a_1962_4178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3491 a_13310_17230# col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3492 a_31478_3496# col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3493 a_3270_17230# col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3494 a_26362_3174# col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3495 VDD rowon_n[1] a_16930_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3496 a_11910_7150# row_n[5] a_12402_7512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3497 a_25358_7190# col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3498 VSS row_n[5] a_35398_7190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3499 a_4274_6186# col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3500 vcm a_1962_15222# a_35094_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3501 a_16322_9198# col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3502 vcm a_1962_7190# a_29070_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3503 a_27974_6146# row_n[4] a_28466_6508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3504 a_12914_15182# row_n[13] a_13406_15544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3505 a_24354_13214# rowon_n[11] a_23958_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3506 vcm a_1962_11206# a_13006_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3507 VSS row_n[8] a_21342_10202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3508 a_2874_15182# row_n[13] a_3366_15544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3509 vcm a_1962_11206# a_2966_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3510 a_21950_11166# a_1962_11206# a_22042_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3511 a_25966_1126# VDD a_26458_1488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3512 a_2346_14220# sample VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3513 a_21038_9158# a_2346_9200# a_20946_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3514 VDD rowon_n[0] a_8898_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3515 a_1962_3174# sample_n VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3516 VDD rowon_n[15] a_18938_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3517 a_29070_15182# a_2346_15224# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3518 VDD rowon_n[10] a_19942_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3519 a_25966_12170# a_1962_12210# a_26058_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3520 a_15926_9158# row_n[7] a_16418_9520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3521 a_14010_6146# a_2346_6188# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3522 a_16930_5142# row_n[3] a_17422_5504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3523 a_30074_2130# a_2346_2172# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3524 a_19942_2130# a_1962_2170# a_20034_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3525 a_9294_4178# col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3526 a_8290_8194# col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3527 VSS sample_n a_1962_11206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3528 VDD rowon_n[9] a_23958_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3529 a_9902_8154# a_1962_8194# a_9994_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3530 a_18330_1166# en_bit_n[1] a_17934_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3531 a_30378_1166# col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3532 a_10906_4138# a_1962_4178# a_10998_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3533 VSS VDD a_22346_18234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3534 VSS row_n[15] a_35398_17230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3535 a_23350_14218# col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3536 vcm a_1962_5182# a_33086_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3537 a_12306_17230# rowon_n[15] a_11910_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3538 a_6982_1126# a_2346_1168# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3539 a_8898_4138# row_n[2] a_9390_4500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3540 a_6282_16226# rowon_n[14] a_5886_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3541 a_16322_16226# rowon_n[14] a_15926_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3542 VSS row_n[11] a_3270_13214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3543 VSS row_n[11] a_13310_13214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3544 a_31078_12170# a_2346_12212# a_30986_12170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3545 a_22442_16548# col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3546 VSS row_n[4] a_11302_6186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3547 a_2874_3134# a_1962_3174# a_2966_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3548 a_35494_15544# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3549 a_31990_12170# row_n[10] a_32482_12532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3550 a_13006_11166# a_2346_11208# a_12914_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3551 a_35094_11166# a_2346_11208# a_35002_11166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3552 a_22442_7512# col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3553 a_14922_6146# a_1962_6186# a_15014_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3554 a_7894_15182# a_1962_15222# a_7986_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3555 a_17934_15182# a_1962_15222# a_18026_15182# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3556 a_2966_11166# a_2346_11208# a_2874_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3557 VDD rowon_n[5] a_31990_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3558 a_18938_2130# row_n[0] a_19430_2492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3559 VDD rowon_n[13] a_11910_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3560 a_20434_2492# col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3561 a_13406_11528# col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3562 VDD rowon_n[0] a_29982_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3563 a_3366_11528# col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3564 a_11302_18234# col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3565 a_35398_2170# rowon_n[0] a_35002_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3566 VSS row_n[0] a_25358_2170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3567 VSS row_n[3] a_3270_5182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3568 vcm a_1962_16226# a_33086_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3569 a_20034_10162# a_2346_10204# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3570 VSS row_n[6] a_15318_8194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3571 a_7894_1126# a_1962_1166# a_7986_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3572 VSS row_n[2] a_16322_4178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3573 VSS row_n[8] a_19334_10202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3574 a_27462_5504# col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3575 vcm a_1962_17230# a_19030_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3576 a_5374_8516# col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3577 a_5978_8154# a_2346_8196# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3578 vcm a_1962_17230# a_8990_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3579 a_12002_6146# a_2346_6188# a_11910_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3580 a_10906_16186# row_n[14] a_11398_16548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3581 a_22346_14218# rowon_n[12] a_21950_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3582 a_35398_13214# rowon_n[11] a_35002_13174# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3583 a_23958_7150# a_1962_7190# a_24050_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3584 a_3366_3496# col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3585 a_23046_17190# a_2346_17232# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3586 VDD rowon_n[10] a_17934_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3587 a_34394_6186# col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3588 a_16418_4500# col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3589 a_27062_16186# a_2346_16228# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3590 a_23958_13174# a_1962_13214# a_24050_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3591 VSS row_n[5] a_7286_7190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3592 VSS row_n[1] a_8290_3174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3593 a_18026_15182# a_2346_15224# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3594 a_7986_15182# a_2346_15224# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3595 a_21342_6186# rowon_n[4] a_20946_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3596 a_4974_1126# a_2346_1168# a_4882_1126# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3597 VSS row_n[10] a_34394_12210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3598 VDD rowon_n[9] a_35002_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3599 a_3970_5142# a_2346_5184# a_3878_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3600 a_11302_12210# rowon_n[10] a_10906_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3601 a_17022_4138# a_2346_4180# a_16930_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3602 VSS VDD a_33390_18234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3603 a_8386_1488# col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3604 a_29470_2492# col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3605 a_28978_5142# a_1962_5182# a_29070_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3606 a_29070_12170# a_2346_12212# a_28978_12170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3607 a_6890_8154# a_1962_8194# a_6982_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3608 vcm a_1962_6186# a_13006_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3609 a_10298_18234# VDD a_9902_18194# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3610 VDD rowon_n[12] a_32994_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3611 a_34394_14218# col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3612 a_28066_18194# a_2346_18236# a_27974_18194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3613 VSS row_n[12] a_11302_14218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3614 a_34490_10524# col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3615 a_10298_5182# rowon_n[3] a_9902_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3616 a_28978_18194# VDD a_29470_18556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3617 VDD sample_n a_1962_17230# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3618 a_11910_17190# a_1962_17230# a_12002_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3619 vcm a_1962_14218# a_29070_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3620 VDD rowon_n[8] a_10906_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3621 a_26362_4178# rowon_n[2] a_25966_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3622 a_15926_16186# a_1962_16226# a_16018_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3623 a_33486_16548# col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3624 VDD rowon_n[6] a_11910_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3625 a_8990_3134# a_2346_3176# a_8898_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3626 a_5886_16186# a_1962_16226# a_5978_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3627 VDD rowon_n[14] a_9902_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3628 a_19030_8154# a_2346_8196# a_18938_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3629 a_10298_13214# col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3630 vcm a_1962_5182# a_4974_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3631 vcm a_1962_1166# a_5978_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3632 VDD rowon_n[1] a_9902_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3633 vcm a_1962_4178# a_18026_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3634 a_25054_9158# a_2346_9200# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3635 a_14314_7190# rowon_n[5] a_13918_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3636 vcm a_1962_7190# a_22042_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3637 a_32994_3134# a_1962_3174# a_33086_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3638 a_15318_3174# rowon_n[1] a_14922_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3639 vcm a_1962_12210# a_18026_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3640 a_20946_6146# row_n[4] a_21438_6508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3641 VDD rowon_n[2] a_25966_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3642 vcm a_1962_12210# a_7986_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3643 a_1962_8194# sample_n VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3644 VDD rowon_n[5] a_3878_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3645 a_31478_6508# col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3646 a_9902_11166# row_n[9] a_10394_11528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3647 a_31078_10162# a_2346_10204# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3648 VDD rowon_n[4] a_16930_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3649 VDD sample a_2346_4180# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3650 vcm a_1962_18234# a_6982_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3651 vcm a_1962_18234# a_17022_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3652 a_8290_9198# rowon_n[7] a_7894_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3653 a_22042_12170# a_2346_12212# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3654 a_2346_9200# sample VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3655 a_1962_14218# sample_n VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3656 VDD VSS a_14922_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3657 a_24354_1166# col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3658 a_23350_5182# col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3659 a_21038_18194# a_2346_18236# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3660 VDD rowon_n[10] a_28978_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3661 a_7286_2170# rowon_n[0] a_6890_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3662 VSS row_n[3] a_33390_5182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3663 vcm a_1962_5182# a_27062_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3664 a_31382_17230# rowon_n[15] a_30986_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3665 a_21950_14178# a_1962_14218# a_22042_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3666 a_24962_8154# row_n[6] a_25454_8516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3667 a_5978_16186# a_2346_16228# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3668 a_16018_16186# a_2346_16228# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3669 VDD rowon_n[7] a_7894_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3670 a_35494_8516# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3671 VDD rowon_n[3] a_8898_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3672 a_28370_15222# col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3673 VSS row_n[11] a_32386_13214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3674 a_19942_17190# a_1962_17230# a_20034_17190# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X3675 a_33486_3496# col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3676 a_22954_3134# row_n[1] a_23446_3496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3677 a_28370_3174# col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3678 a_12002_4138# a_2346_4180# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3679 a_27462_17552# col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3680 VDD rowon_n[13] a_30986_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3681 a_23958_14178# row_n[12] a_24450_14540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3682 a_27062_13174# a_2346_13216# a_26970_13174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3683 a_9294_10202# col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3684 a_19334_10202# col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3685 vcm a_1962_10202# a_24050_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3686 a_13918_7150# row_n[5] a_14410_7512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3687 a_6282_6186# col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3688 a_7986_12170# a_2346_12212# a_7894_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3689 a_10906_12170# a_1962_12210# a_10998_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3690 a_18026_12170# a_2346_12212# a_17934_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3691 a_18330_9198# col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3692 a_27974_13174# row_n[11] a_28466_13536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3693 a_32482_11528# col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3694 a_11910_2130# row_n[0] a_12402_2492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3695 a_30378_18234# col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3696 a_8386_12532# col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3697 a_18426_12532# col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3698 a_17326_2170# col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3699 a_23046_9158# a_2346_9200# a_22954_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3700 vcm a_1962_7190# a_30074_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3701 a_27974_1126# VDD a_28466_1488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3702 vcm a_1962_3174# a_31078_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3703 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X3704 a_3970_3134# a_2346_3176# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3705 vcm a_1962_18234# a_25054_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3706 a_17934_9158# row_n[7] a_18426_9520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3707 a_18938_5142# row_n[3] a_19430_5504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3708 a_32082_2130# a_2346_2172# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3709 a_29982_16186# row_n[14] a_30474_16548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3710 a_12914_4138# a_1962_4178# a_13006_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3711 a_20434_5504# col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3712 VSS sample a_2346_10204# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3713 a_29070_10162# a_2346_10204# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3714 VDD rowon_n[3] a_29982_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3715 a_15926_17190# row_n[15] a_16418_17552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3716 a_27366_15222# rowon_n[13] a_26970_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3717 vcm a_1962_13214# a_16018_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3718 a_5886_17190# row_n[15] a_6378_17552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3719 vcm a_1962_13214# a_5978_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3720 VSS row_n[9] a_28370_11206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3721 vcm a_1962_5182# a_35094_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3722 a_19030_18194# a_2346_18236# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3723 a_20034_13174# a_2346_13216# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3724 a_8990_1126# a_2346_1168# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3725 a_10998_12170# a_2346_12212# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3726 a_33086_12170# a_2346_12212# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3727 VSS row_n[4] a_13310_6186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3728 a_19030_6146# a_2346_6188# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3729 a_4882_3134# a_1962_3174# a_4974_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3730 VDD rowon_n[11] a_26970_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3731 a_24450_7512# col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3732 VDD rowon_n[5] a_33998_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3733 a_3366_6508# col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3734 a_22346_17230# col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3735 a_16018_9158# a_2346_9200# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3736 a_22442_2492# col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3737 a_21950_5142# a_1962_5182# a_22042_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3738 a_26362_16226# col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3739 VSS row_n[12] a_30378_14218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3740 a_17934_10162# a_1962_10202# a_18026_10162# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3741 VDD rowon_n[0] a_31990_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3742 a_30986_17190# a_1962_17230# a_31078_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3743 a_7894_10162# a_1962_10202# a_7986_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3744 VSS row_n[0] a_27366_2170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3745 a_9294_18234# VDD a_8898_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3746 VSS row_n[13] a_6282_15222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3747 VSS row_n[13] a_16322_15222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3748 a_21038_15182# a_2346_15224# a_20946_15182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3749 a_19334_8194# rowon_n[6] a_18938_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3750 a_31382_8194# col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3751 VSS row_n[3] a_5278_5182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3752 VSS VDD a_6282_1166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3753 a_32386_4178# col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3754 a_35002_16186# a_1962_16226# a_35094_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3755 a_25054_14178# a_2346_14220# a_24962_14178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3756 a_17326_11206# col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3757 vcm a_1962_11206# a_22042_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3758 VSS row_n[2] a_18330_4178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3759 a_25454_18556# col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3760 a_21950_15182# row_n[13] a_22442_15544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3761 a_16018_13174# a_2346_13216# a_15926_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3762 a_7286_11206# col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3763 VSS row_n[6] a_17326_8194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3764 a_29470_5504# col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3765 a_5978_13174# a_2346_13216# a_5886_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3766 a_7382_8516# col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3767 VDD rowon_n[15] a_4882_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3768 VDD rowon_n[15] a_14922_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3769 a_7986_8154# a_2346_8196# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3770 a_14010_6146# a_2346_6188# a_13918_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3771 vcm a_1962_2170# a_20034_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3772 a_16418_13536# col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3773 a_25966_7150# a_1962_7190# a_26058_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3774 a_30074_2130# a_2346_2172# a_29982_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3775 a_26970_3134# a_1962_3174# a_27062_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3776 VDD rowon_n[14] a_8898_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3777 a_6378_13536# col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3778 vcm a_1962_8194# a_9994_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3779 a_5374_3496# col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3780 a_31990_4138# row_n[2] a_32482_4500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3781 vcm a_1962_4178# a_10998_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3782 a_16930_9158# a_1962_9198# a_17022_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3783 a_18426_4500# col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3784 VSS row_n[5] a_9294_7190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3785 a_4882_12170# row_n[10] a_5374_12532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3786 a_14922_12170# row_n[10] a_15414_12532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3787 a_27062_11166# a_2346_11208# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3788 a_26362_10202# rowon_n[8] a_25966_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3789 a_23350_6186# rowon_n[4] a_22954_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3790 a_6982_1126# a_2346_1168# a_6890_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3791 a_18026_10162# a_2346_10204# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3792 VDD rowon_n[4] a_9902_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3793 a_3878_18194# VDD a_4370_18556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3794 a_13918_18194# VDD a_14410_18556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3795 a_25358_16226# rowon_n[14] a_24962_16186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3796 vcm a_1962_14218# a_3970_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3797 vcm a_1962_14218# a_14010_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3798 a_7986_10162# a_2346_10204# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3799 vcm a_1962_3174# a_2966_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3800 a_8898_8154# a_1962_8194# a_8990_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3801 vcm a_1962_6186# a_15014_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3802 a_26970_15182# a_1962_15222# a_27062_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3803 a_31078_13174# a_2346_13216# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3804 a_30986_1126# a_1962_1166# a_31078_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3805 a_29982_5142# a_1962_5182# a_30074_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3806 a_12306_5182# rowon_n[3] a_11910_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3807 VSS row_n[13] a_24354_15222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3808 a_21342_12210# col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3809 a_28370_4178# rowon_n[2] a_27974_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3810 a_25358_11206# col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3811 VDD rowon_n[6] a_13918_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3812 vcm a_1962_1166# a_7986_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3813 VDD rowon_n[15] a_22954_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3814 a_19030_15182# a_2346_15224# a_18938_15182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3815 a_20434_14540# col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3816 a_29982_12170# a_1962_12210# a_30074_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3817 VSS row_n[8] a_15318_10202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3818 a_20034_10162# a_2346_10204# a_19942_10162# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3819 a_21342_3174# col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3820 VDD rowon_n[1] a_11910_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3821 a_8290_13214# rowon_n[11] a_7894_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3822 a_5886_11166# a_1962_11206# a_5978_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3823 a_15926_11166# a_1962_11206# a_16018_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3824 VSS row_n[8] a_5278_10202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3825 a_20338_7190# col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3826 VSS row_n[5] a_30378_7190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3827 VSS row_n[1] a_31382_3174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3828 a_24450_13536# col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3829 a_20946_10162# row_n[8] a_21438_10524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3830 a_5978_8154# a_2346_8196# a_5886_8154# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3831 a_35002_3134# a_1962_3174# a_35094_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3832 a_11302_9198# col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3833 a_27062_9158# a_2346_9200# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3834 a_16322_7190# rowon_n[5] a_15926_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3835 vcm a_1962_7190# a_24050_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3836 a_22954_6146# row_n[4] a_23446_6508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3837 a_17326_3174# rowon_n[1] a_16930_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3838 VDD rowon_n[10] a_13918_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3839 a_33486_6508# col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3840 VDD rowon_n[2] a_27974_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3841 VDD rowon_n[10] a_3878_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3842 VDD rowon_n[5] a_5886_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3843 a_8898_18194# a_1962_18234# a_8990_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3844 a_18938_18194# a_1962_18234# a_19030_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3845 VDD rowon_n[9] a_7894_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3846 a_20946_1126# VDD a_21438_1488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3847 a_26058_2130# a_2346_2172# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3848 a_13310_15222# col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3849 a_31478_1488# col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3850 VDD rowon_n[0] a_3878_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3851 a_12002_17190# a_2346_17232# a_11910_17190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3852 a_34090_17190# a_2346_17232# a_33998_17190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3853 a_3270_15222# col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3854 VDD VSS a_16930_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3855 a_26362_1166# col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3856 a_10906_9158# row_n[7] a_11398_9520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3857 a_11910_5142# row_n[3] a_12402_5504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3858 a_4274_4178# col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3859 VSS row_n[3] a_35398_5182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3860 a_25358_5182# col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3861 a_35002_17190# row_n[15] a_35494_17552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3862 vcm a_1962_13214# a_35094_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3863 a_3270_8194# col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3864 a_9294_2170# rowon_n[0] a_8898_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3865 a_2346_4180# sample VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3866 a_12402_17552# col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3867 a_19334_17230# rowon_n[15] a_18938_17190# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3868 vcm a_1962_5182# a_29070_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3869 a_20338_12210# rowon_n[10] a_19942_12170# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3870 vcm a_1962_8194# a_6982_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3871 a_12914_13174# row_n[11] a_13406_13536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3872 a_24354_11206# rowon_n[9] a_23958_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3873 a_2874_13174# row_n[11] a_3366_13536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3874 a_24962_3134# row_n[1] a_25454_3496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3875 a_2346_12212# sample VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3876 a_5978_11166# a_2346_11208# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3877 a_16018_11166# a_2346_11208# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3878 a_1962_1166# sample_n VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3879 a_35494_3496# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3880 a_29070_13174# a_2346_13216# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3881 a_3878_4138# row_n[2] a_4370_4500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3882 VDD rowon_n[13] a_18938_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3883 VDD rowon_n[8] a_19942_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3884 a_15926_7150# row_n[5] a_16418_7512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3885 a_14010_4138# a_2346_4180# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3886 a_9994_12170# a_2346_12212# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3887 a_8290_6186# col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3888 vcm a_1962_18234# a_9994_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3889 a_9902_6146# a_1962_6186# a_9994_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3890 a_13918_2130# row_n[0] a_14410_2492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3891 VSS row_n[14] a_22346_16226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3892 VSS row_n[13] a_35398_15222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3893 a_32386_12210# col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3894 a_31382_9198# rowon_n[7] a_30986_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3895 a_19334_2170# col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3896 vcm a_1962_3174# a_33086_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3897 a_12306_15222# rowon_n[13] a_11910_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3898 a_25054_9158# a_2346_9200# a_24962_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3899 a_30378_2170# rowon_n[0] a_29982_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3900 VSS row_n[0] a_20338_2170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3901 VDD VDD a_20946_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3902 VDD rowon_n[15] a_33998_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3903 a_6282_14218# rowon_n[12] a_5886_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3904 a_16322_14218# rowon_n[12] a_15926_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3905 a_31478_14540# col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3906 vcm a_1962_12210# a_27062_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3907 VSS row_n[9] a_3270_11206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3908 VSS row_n[9] a_13310_11206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3909 a_31078_10162# a_2346_10204# a_30986_10162# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3910 VSS row_n[6] a_10298_8194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3911 a_34090_2130# a_2346_2172# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3912 a_2874_1126# a_1962_1166# a_2966_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3913 VSS row_n[2] a_11302_4178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3914 a_35494_13536# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3915 a_31990_10162# row_n[8] a_32482_10524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3916 a_14922_4138# a_1962_4178# a_15014_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3917 a_22442_5504# col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3918 a_7894_13174# a_1962_13214# a_7986_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3919 a_17934_13174# a_1962_13214# a_18026_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3920 VDD rowon_n[7] a_30986_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3921 VDD rowon_n[3] a_31990_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3922 VDD rowon_n[11] a_11910_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3923 a_11302_16226# col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3924 a_11398_4500# col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3925 a_32082_18194# a_2346_18236# a_31990_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3926 VSS row_n[1] a_3270_3174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3927 a_32994_18194# VDD a_33486_18556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3928 vcm a_1962_14218# a_33086_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3929 a_18330_12210# rowon_n[10] a_17934_12170# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3930 VSS row_n[4] a_15318_6186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3931 a_10394_18556# col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3932 vcm a_1962_15222# a_19030_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3933 a_5374_6508# col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3934 a_5978_6146# a_2346_6188# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3935 a_12002_4138# a_2346_4180# a_11910_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3936 vcm a_1962_15222# a_8990_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3937 a_35398_11206# rowon_n[9] a_35002_11166# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3938 a_18026_9158# a_2346_9200# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3939 VDD rowon_n[0] a_33998_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3940 a_3366_1488# col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3941 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X3942 a_24450_2492# col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3943 a_23958_5142# a_1962_5182# a_24050_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3944 a_23046_15182# a_2346_15224# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3945 VDD rowon_n[8] a_17934_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3946 VDD sample_n a_1962_8194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3947 VSS row_n[0] a_29374_2170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3948 a_34394_4178# col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3949 a_27062_14178# a_2346_14220# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3950 a_33390_8194# col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3951 VSS row_n[3] a_7286_5182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3952 VSS VDD a_8290_1166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3953 a_18026_13174# a_2346_13216# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3954 a_7986_13174# a_2346_13216# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3955 a_3970_3134# a_2346_3176# a_3878_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3956 a_21342_4178# rowon_n[2] a_20946_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3957 a_35002_11166# a_1962_11206# a_35094_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3958 VSS row_n[8] a_34394_10202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3959 a_9390_8516# col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3960 a_11302_10202# rowon_n[8] a_10906_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3961 a_9994_8154# a_2346_8196# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3962 a_32082_2130# a_2346_2172# a_31990_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3963 a_29374_18234# col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3964 VSS row_n[14] a_33390_16226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3965 a_27974_7150# a_1962_7190# a_28066_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3966 a_28978_3134# a_1962_3174# a_29070_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3967 a_10298_16226# rowon_n[14] a_9902_16186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3968 a_29470_14540# col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3969 VDD rowon_n[10] a_32994_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3970 a_29070_10162# a_2346_10204# a_28978_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3971 a_6890_6146# a_1962_6186# a_6982_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3972 a_7382_3496# col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3973 a_33998_4138# row_n[2] a_34490_4500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3974 vcm a_1962_4178# a_13006_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3975 a_18938_9158# a_1962_9198# a_19030_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3976 a_28066_16186# a_2346_16228# a_27974_16186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3977 a_20034_9158# a_2346_9200# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3978 a_10298_3174# rowon_n[1] a_9902_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3979 VDD VDD a_31990_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3980 VDD rowon_n[2] a_20946_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3981 a_28978_16186# row_n[14] a_29470_16548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3982 VDD sample_n a_1962_15222# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3983 a_11910_15182# a_1962_15222# a_12002_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3984 a_8990_1126# a_2346_1168# a_8898_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3985 a_15926_14178# a_1962_14218# a_16018_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3986 VDD rowon_n[4] a_11910_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3987 a_5886_14178# a_1962_14218# a_5978_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3988 a_3270_9198# rowon_n[7] a_2874_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3989 a_19030_6146# a_2346_6188# a_18938_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3990 a_10298_11206# col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3991 vcm a_1962_3174# a_4974_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3992 VDD VSS a_9902_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3993 a_16018_9158# a_2346_9200# a_15926_9158# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3994 a_14314_5182# rowon_n[3] a_13918_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3995 a_15318_1166# VSS a_14922_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3996 a_32994_1126# a_1962_1166# a_33086_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3997 vcm a_1962_5182# a_22042_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3998 a_2346_17232# sample VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3999 vcm a_1962_10202# a_18026_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4000 a_19942_8154# row_n[6] a_20434_8516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4001 a_7894_14178# row_n[12] a_8386_14540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4002 a_17934_14178# row_n[12] a_18426_14540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4003 a_29374_12210# rowon_n[10] a_28978_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4004 vcm a_1962_10202# a_7986_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4005 a_26970_10162# a_1962_10202# a_27062_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4006 VDD rowon_n[7] a_2874_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4007 a_30474_8516# col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4008 a_1962_6186# sample_n VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4009 VDD rowon_n[3] a_3878_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4010 VDD rowon_n[6] a_15926_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4011 VDD sample a_2346_2172# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4012 vcm a_1962_16226# a_6982_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4013 vcm a_1962_16226# a_17022_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4014 a_23350_3174# col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4015 VDD rowon_n[1] a_13918_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4016 a_21038_16186# a_2346_16228# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4017 VDD rowon_n[8] a_28978_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4018 a_25358_9198# rowon_n[7] a_24962_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4019 a_7986_8154# a_2346_8196# a_7894_8154# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4020 VSS row_n[5] a_32386_7190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4021 VSS row_n[1] a_33390_3174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4022 a_13310_9198# col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4023 vcm a_1962_3174# a_27062_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4024 VSS row_n[15] a_27366_17230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4025 a_31382_15222# rowon_n[13] a_30986_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4026 a_29070_9158# a_2346_9200# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4027 vcm a_1962_7190# a_26058_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4028 a_24962_6146# row_n[4] a_25454_6508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4029 a_5978_14178# a_2346_14220# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4030 a_16018_14178# a_2346_14220# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4031 VDD rowon_n[5] a_7894_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4032 a_35494_6508# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4033 a_28370_13214# col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4034 VSS row_n[9] a_32386_11206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4035 vcm a_1962_9198# a_17022_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4036 a_12306_2170# col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4037 a_19942_15182# a_1962_15222# a_20034_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4038 a_22954_1126# VDD a_23446_1488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4039 a_33486_1488# col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4040 a_28066_2130# a_2346_2172# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4041 a_14010_17190# a_2346_17232# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4042 VSS row_n[10] a_18330_12210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4043 a_23046_12170# a_2346_12212# a_22954_12170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4044 a_31990_8154# a_1962_8194# a_32082_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4045 VDD rowon_n[0] a_5886_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4046 a_3970_17190# a_2346_17232# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4047 VSS row_n[10] a_8290_12210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4048 VDD rowon_n[7] a_24962_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4049 a_28370_1166# col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4050 a_27462_15544# col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4051 VDD rowon_n[11] a_30986_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4052 a_23958_12170# row_n[10] a_24450_12532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4053 a_27062_11166# a_2346_11208# a_26970_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4054 a_12914_9158# row_n[7] a_13406_9520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4055 a_5278_8194# col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4056 a_13918_5142# row_n[3] a_14410_5504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4057 a_6282_4178# col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4058 a_7986_10162# a_2346_10204# a_7894_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4059 a_18026_10162# a_2346_10204# a_17934_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4060 VDD rowon_n[12] a_16930_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4061 a_27974_11166# row_n[9] a_28466_11528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4062 VDD rowon_n[12] a_6890_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4063 vcm a_1962_8194# a_8990_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4064 a_30378_16226# col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4065 a_8386_10524# col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4066 a_18426_10524# col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4067 vcm a_1962_1166# a_31078_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4068 vcm a_1962_17230# a_21038_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4069 vcm a_1962_5182# a_30074_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4070 a_6282_17230# col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4071 a_16322_17230# col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4072 a_3970_1126# a_2346_1168# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4073 vcm a_1962_16226# a_25054_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4074 a_5886_4138# row_n[2] a_6378_4500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4075 a_17934_7150# row_n[5] a_18426_7512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4076 ctop sw_n analog_in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.9e+06u l=220000u
X4077 a_8990_18194# a_2346_18236# a_8898_18194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4078 vcm a_1962_12210# a_12002_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4079 a_15926_2130# row_n[0] a_16418_2492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4080 a_15926_15182# row_n[13] a_16418_15544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4081 a_27366_13214# rowon_n[11] a_26970_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4082 vcm a_1962_11206# a_16018_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4083 a_9390_18556# col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4084 a_5886_15182# row_n[13] a_6378_15544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4085 vcm a_1962_11206# a_5978_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4086 a_10998_9158# a_2346_9200# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4087 a_33390_9198# rowon_n[7] a_32994_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4088 a_27366_8194# col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4089 a_27062_9158# a_2346_9200# a_26970_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4090 vcm a_1962_3174# a_35094_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4091 a_19030_16186# a_2346_16228# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4092 VSS row_n[0] a_22346_2170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4093 a_28978_12170# a_1962_12210# a_29070_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4094 a_32386_2170# rowon_n[0] a_31990_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4095 a_4882_1126# a_1962_1166# a_4974_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4096 a_19030_4138# a_2346_4180# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4097 VSS row_n[2] a_13310_4178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4098 VDD rowon_n[9] a_26970_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4099 VSS row_n[6] a_12306_8194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4100 a_26058_2130# a_2346_2172# a_25966_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4101 a_24450_5504# col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4102 VDD rowon_n[7] a_32994_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4103 VDD rowon_n[3] a_33998_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4104 VSS VDD a_25358_18234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4105 a_22346_15222# col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4106 a_2966_8154# a_2346_8196# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4107 a_26362_14218# col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4108 a_20946_7150# a_1962_7190# a_21038_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4109 a_21950_3134# a_1962_3174# a_22042_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4110 a_15318_17230# rowon_n[15] a_14922_17190# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4111 a_31078_7150# a_2346_7192# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4112 a_34090_18194# a_2346_18236# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4113 a_5278_17230# rowon_n[15] a_4882_17190# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4114 a_30986_15182# a_1962_15222# a_31078_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4115 a_11910_9158# a_1962_9198# a_12002_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4116 a_1962_18234# sample_n VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4117 a_12002_18194# a_2346_18236# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4118 a_21438_17552# col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4119 a_9294_16226# rowon_n[14] a_8898_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4120 VSS row_n[11] a_6282_13214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4121 VSS row_n[11] a_16322_13214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4122 a_21038_13174# a_2346_13216# a_20946_13174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4123 a_19334_6186# rowon_n[4] a_18938_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4124 a_31382_6186# col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4125 VSS row_n[1] a_5278_3174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4126 a_13406_4500# col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4127 a_25454_16548# col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4128 a_35002_14178# a_1962_14218# a_35094_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4129 a_21950_13174# row_n[11] a_22442_13536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4130 VSS row_n[5] a_4274_7190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4131 a_16018_11166# a_2346_11208# a_15926_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4132 VSS row_n[4] a_17326_6186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4133 a_5978_11166# a_2346_11208# a_5886_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4134 a_7382_6508# col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4135 VDD rowon_n[13] a_4882_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4136 VDD rowon_n[13] a_14922_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4137 a_7986_6146# a_2346_6188# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4138 a_14010_4138# a_2346_4180# a_13918_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4139 a_5278_12210# col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4140 a_15318_12210# col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4141 vcm a_1962_12210# a_20034_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4142 a_16418_11528# col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4143 a_26970_1126# a_1962_1166# a_27062_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4144 a_25966_5142# a_1962_5182# a_26058_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4145 a_6378_11528# col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4146 a_3878_8154# a_1962_8194# a_3970_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4147 vcm a_1962_6186# a_9994_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4148 a_5374_1488# col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4149 a_14314_18234# col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4150 a_4274_18234# col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4151 vcm a_1962_17230# a_32082_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4152 a_35398_8194# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4153 a_4370_14540# col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4154 a_14410_14540# col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4155 VSS sample a_2346_7192# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4156 VSS row_n[3] a_9294_5182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4157 a_14922_10162# row_n[8] a_15414_10524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4158 a_23046_10162# a_2346_10204# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4159 a_4882_10162# row_n[8] a_5374_10524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4160 a_23350_4178# rowon_n[2] a_22954_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4161 VSS row_n[5] a_26362_7190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4162 a_3878_16186# row_n[14] a_4370_16548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4163 a_13918_16186# row_n[14] a_14410_16548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4164 a_25358_14218# rowon_n[12] a_24962_14178# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X4165 a_34090_2130# a_2346_2172# a_33998_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4166 vcm a_1962_1166# a_2966_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4167 a_8898_6146# a_1962_6186# a_8990_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4168 a_9390_3496# col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4169 vcm a_1962_4178# a_15014_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4170 a_26058_17190# a_2346_17232# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4171 a_23350_17230# rowon_n[15] a_22954_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4172 a_26970_13174# a_1962_13214# a_27062_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4173 a_29982_3134# a_1962_3174# a_30074_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4174 a_22042_9158# a_2346_9200# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4175 a_11302_7190# rowon_n[5] a_10906_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4176 a_12306_3174# rowon_n[1] a_11910_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4177 VSS row_n[11] a_24354_13214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4178 a_21342_10202# col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4179 VDD rowon_n[2] a_22954_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4180 VDD sample a_2346_14220# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4181 a_14314_12210# rowon_n[10] a_13918_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4182 VDD rowon_n[4] a_13918_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4183 a_21038_2130# a_2346_2172# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4184 a_4274_12210# rowon_n[10] a_3878_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4185 a_11910_10162# a_1962_10202# a_12002_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4186 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.64e+07u l=1.6e+07u
X4187 a_19430_17552# col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4188 VDD rowon_n[13] a_22954_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4189 a_19030_13174# a_2346_13216# a_18938_13174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4190 a_20434_12532# col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4191 VDD sample_n a_1962_10202# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4192 VDD VSS a_11910_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4193 a_21342_1166# col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4194 a_8290_11206# rowon_n[9] a_7894_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4195 VSS VDD a_31382_1166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4196 VSS row_n[3] a_30378_5182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4197 a_20338_5182# col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4198 a_24450_11528# col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4199 a_5978_6146# a_2346_6188# a_5886_6146# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4200 a_35002_1126# a_1962_1166# a_35094_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4201 a_4274_2170# rowon_n[0] a_3878_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4202 a_18026_9158# a_2346_9200# a_17934_9158# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4203 a_16322_5182# rowon_n[3] a_15926_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4204 a_17326_1166# VSS a_16930_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4205 vcm a_1962_5182# a_24050_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4206 a_35398_17230# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4207 VDD rowon_n[8] a_13918_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4208 a_32482_8516# col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4209 VDD rowon_n[8] a_3878_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4210 VDD rowon_n[3] a_5886_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4211 VSS row_n[15] a_12306_17230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4212 a_8898_16186# a_1962_16226# a_8990_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4213 a_18938_16186# a_1962_16226# a_19030_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4214 a_19942_3134# row_n[1] a_20434_3496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4215 a_13310_13214# col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4216 a_30474_3496# col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4217 a_12002_15182# a_2346_15224# a_11910_15182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4218 a_34090_15182# a_2346_15224# a_33998_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4219 a_3270_13214# col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4220 vcm a_1962_12210# a_31078_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4221 a_25358_3174# col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4222 a_10906_7150# row_n[5] a_11398_7512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4223 VSS row_n[1] a_35398_3174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4224 VDD rowon_n[1] a_15926_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4225 a_35002_15182# row_n[13] a_35494_15544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4226 vcm a_1962_11206# a_35094_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4227 a_27366_9198# rowon_n[7] a_26970_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4228 a_9994_8154# a_2346_8196# a_9902_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4229 VSS row_n[5] a_34394_7190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4230 a_3270_6186# col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4231 a_2346_2172# sample VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4232 a_12402_15544# col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4233 a_19334_15222# rowon_n[13] a_18938_15182# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X4234 a_20338_10202# rowon_n[8] a_19942_10162# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X4235 a_15318_9198# col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4236 vcm a_1962_7190# a_28066_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4237 vcm a_1962_3174# a_29070_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4238 a_21038_11166# a_2346_11208# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4239 vcm a_1962_6186# a_6982_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4240 a_12914_11166# row_n[9] a_13406_11528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4241 vcm a_1962_9198# a_19030_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4242 a_2874_11166# row_n[9] a_3366_11528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4243 a_24962_1126# VDD a_25454_1488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4244 a_14314_2170# col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4245 a_25054_12170# a_2346_12212# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4246 a_20034_9158# a_2346_9200# a_19942_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4247 a_33998_8154# a_1962_8194# a_34090_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4248 a_35494_1488# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4249 VDD rowon_n[0] a_7894_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4250 VDD rowon_n[11] a_18938_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4251 a_19942_10162# a_1962_10202# a_20034_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4252 a_14922_9158# row_n[7] a_15414_9520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4253 VDD rowon_n[7] a_26970_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4254 a_15926_5142# row_n[3] a_16418_5504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4255 a_8290_4178# col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4256 a_21342_18234# VDD a_20946_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4257 vcm a_1962_16226# a_9994_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4258 a_9902_4138# a_1962_4178# a_9994_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4259 a_34394_17230# rowon_n[15] a_33998_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4260 VSS row_n[12] a_22346_14218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4261 VSS row_n[11] a_35398_13214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4262 a_32386_10202# col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4263 a_22954_17190# a_1962_17230# a_23046_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4264 vcm a_1962_1166# a_33086_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4265 a_12306_13214# rowon_n[11] a_11910_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4266 a_7894_4138# row_n[2] a_8386_4500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4267 VDD rowon_n[14] a_20946_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4268 VDD rowon_n[13] a_33998_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4269 a_26970_14178# row_n[12] a_27462_14540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4270 a_31478_12532# col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4271 vcm a_1962_10202# a_27062_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4272 a_13918_12170# a_1962_12210# a_14010_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4273 VSS row_n[4] a_10298_6186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4274 a_3878_12170# a_1962_12210# a_3970_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4275 a_35494_11528# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4276 VDD rowon_n[5] a_30986_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4277 a_17934_2130# row_n[0] a_18426_2492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4278 a_33390_18234# col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4279 VDD rowon_n[9] a_11910_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4280 a_29374_8194# col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4281 VSS VDD a_10298_18234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4282 a_13006_9158# a_2346_9200# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4283 a_29070_9158# a_2346_9200# a_28978_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4284 vcm a_1962_18234# a_28066_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4285 a_32082_16186# a_2346_16228# a_31990_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4286 a_11302_14218# col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4287 VSS row_n[0] a_24354_2170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4288 a_18330_10202# rowon_n[8] a_17934_10162# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X4289 a_34394_2170# rowon_n[0] a_33998_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4290 VSS VDD a_3270_1166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4291 a_32994_16186# row_n[14] a_33486_16548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4292 a_19030_11166# a_2346_11208# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4293 VSS row_n[6] a_14314_8194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4294 a_28066_2130# a_2346_2172# a_27974_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4295 VSS row_n[2] a_15318_4178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4296 vcm a_1962_8194# a_32082_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4297 a_18938_17190# row_n[15] a_19430_17552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4298 a_10394_16548# col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4299 vcm a_1962_13214# a_19030_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4300 a_4370_8516# col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4301 a_5978_4138# a_2346_4180# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4302 a_8898_17190# row_n[15] a_9390_17552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4303 vcm a_1962_13214# a_8990_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4304 a_4974_8154# a_2346_8196# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4305 a_23958_3134# a_1962_3174# a_24050_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4306 a_22954_7150# a_1962_7190# a_23046_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4307 a_23046_13174# a_2346_13216# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4308 a_33086_7150# a_2346_7192# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4309 VDD sample_n a_1962_6186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4310 a_13918_9158# a_1962_9198# a_14010_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4311 a_33390_6186# col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4312 VSS row_n[1] a_7286_3174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4313 a_15414_4500# col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4314 a_33390_12210# rowon_n[10] a_32994_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4315 a_30986_10162# a_1962_10202# a_31078_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4316 a_3970_1126# a_2346_1168# a_3878_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4317 a_32386_18234# VDD a_31990_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4318 a_9390_6508# col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4319 a_9994_6146# a_2346_6188# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4320 a_28978_1126# a_1962_1166# a_29070_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4321 a_29374_16226# col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4322 VSS row_n[12] a_33390_14218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4323 a_27974_5142# a_1962_5182# a_28066_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4324 a_20946_18194# a_1962_18234# a_21038_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4325 a_33998_17190# a_1962_17230# a_34090_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4326 a_10298_14218# rowon_n[12] a_9902_14178# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X4327 a_29470_12532# col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4328 VDD rowon_n[8] a_32994_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4329 a_5886_8154# a_1962_8194# a_5978_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4330 a_7382_1488# col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4331 a_6890_4138# a_1962_4178# a_6982_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4332 a_26458_8516# col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4333 a_28066_14178# a_2346_14220# a_27974_14178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4334 a_10998_9158# a_2346_9200# a_10906_9158# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4335 a_10298_1166# VSS a_9902_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4336 a_28466_18556# col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4337 VDD rowon_n[14] a_31990_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4338 VDD sample_n a_1962_13214# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4339 a_11910_13174# a_1962_13214# a_12002_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4340 VDD rowon_n[6] a_10906_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4341 VSS row_n[5] a_28370_7190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4342 a_19030_4138# a_2346_4180# a_18938_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4343 vcm a_1962_1166# a_4974_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4344 a_20338_9198# rowon_n[7] a_19942_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4345 a_2966_8154# a_2346_8196# a_2874_8154# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4346 a_13310_7190# rowon_n[5] a_12914_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4347 vcm a_1962_3174# a_22042_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4348 a_14314_3174# rowon_n[1] a_13918_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4349 a_2346_15224# sample VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4350 a_24050_9158# a_2346_9200# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4351 vcm a_1962_7190# a_21038_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4352 a_31078_7150# a_2346_7192# a_30986_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4353 a_19942_6146# row_n[4] a_20434_6508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4354 a_7894_12170# row_n[10] a_8386_12532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4355 a_17934_12170# row_n[10] a_18426_12532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4356 a_29374_10202# rowon_n[8] a_28978_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4357 VDD rowon_n[5] a_2874_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4358 a_30474_6508# col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4359 a_1962_4178# sample_n VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4360 vcm a_1962_9198# a_12002_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4361 VDD rowon_n[4] a_15926_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4362 a_16930_18194# VDD a_17422_18556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4363 vcm a_1962_14218# a_6982_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4364 vcm a_1962_14218# a_17022_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4365 a_23046_2130# a_2346_2172# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4366 a_6890_18194# VDD a_7382_18556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4367 VDD rowon_n[7] a_19942_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4368 VDD VSS a_13918_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4369 a_23350_1166# col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4370 vcm a_1962_17230# a_15014_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4371 a_21038_14178# a_2346_14220# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4372 a_7986_6146# a_2346_6188# a_7894_6146# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4373 VSS VDD a_33390_1166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4374 a_6282_2170# rowon_n[0] a_5886_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4375 VSS row_n[3] a_32386_5182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4376 vcm a_1962_17230# a_4974_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4377 vcm a_1962_1166# a_27062_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4378 VSS row_n[13] a_27366_15222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4379 a_31382_13214# rowon_n[11] a_30986_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4380 a_24354_12210# col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4381 vcm a_1962_5182# a_26058_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4382 vcm a_1962_8194# a_3970_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4383 a_34490_8516# col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4384 VDD rowon_n[3] a_7894_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4385 a_28370_11206# col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4386 a_19942_13174# a_1962_13214# a_20034_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4387 VDD rowon_n[15] a_25966_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4388 a_14010_15182# a_2346_15224# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4389 a_23446_14540# col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4390 a_32994_12170# a_1962_12210# a_33086_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4391 VSS row_n[8] a_18330_10202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4392 a_23046_10162# a_2346_10204# a_22954_10162# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4393 a_31990_6146# a_1962_6186# a_32082_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4394 a_32482_3496# col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4395 a_3970_15182# a_2346_15224# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4396 a_8898_11166# a_1962_11206# a_8990_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4397 a_18938_11166# a_1962_11206# a_19030_11166# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X4398 VSS row_n[8] a_8290_10202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4399 VDD rowon_n[5] a_24962_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4400 a_31990_18194# a_1962_18234# a_32082_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4401 a_27462_13536# col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4402 VDD rowon_n[9] a_30986_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4403 a_23958_10162# row_n[8] a_24450_10524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4404 VSS row_n[7] a_19334_9198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4405 a_12914_7150# row_n[5] a_13406_7512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4406 a_5278_6186# col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4407 a_29374_9198# rowon_n[7] a_28978_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4408 VDD rowon_n[10] a_16930_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4409 a_10906_2130# row_n[0] a_11398_2492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4410 VDD rowon_n[10] a_6890_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4411 vcm a_1962_6186# a_8990_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4412 a_30378_14218# col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4413 a_22346_8194# col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4414 a_24050_18194# a_2346_18236# a_23958_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4415 a_16322_15222# col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4416 vcm a_1962_15222# a_21038_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4417 a_22042_9158# a_2346_9200# a_21950_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4418 a_16322_2170# col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4419 vcm a_1962_3174# a_30074_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4420 VSS VDD a_9294_18234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4421 a_15014_17190# a_2346_17232# a_14922_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4422 a_6282_15222# col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4423 a_19430_9520# col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4424 a_24962_18194# VDD a_25454_18556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4425 a_4974_17190# a_2346_17232# a_4882_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4426 vcm a_1962_14218# a_25054_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4427 VDD rowon_n[7] a_28978_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4428 a_17934_5142# row_n[3] a_18426_5504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4429 a_15414_17552# col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4430 a_8990_16186# a_2346_16228# a_8898_16186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4431 vcm a_1962_10202# a_12002_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4432 a_21038_2130# a_2346_2172# a_20946_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4433 a_5374_17552# col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4434 a_11910_14178# row_n[12] a_12402_14540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4435 a_15926_13174# row_n[11] a_16418_13536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4436 a_27366_11206# rowon_n[9] a_26970_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4437 a_9390_16548# col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4438 a_5886_13174# row_n[11] a_6378_13536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4439 a_27366_6186# col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4440 vcm a_1962_1166# a_35094_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4441 a_19030_14178# a_2346_14220# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4442 vcm a_1962_18234# a_2966_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4443 vcm a_1962_18234# a_13006_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4444 VSS row_n[15] a_21342_17230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4445 VSS row_n[4] a_12306_6186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4446 VDD rowon_n[5] a_32994_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4447 VSS row_n[14] a_25358_16226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4448 a_22346_13214# col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4449 a_2966_6146# a_2346_6188# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4450 a_15014_9158# a_2346_9200# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4451 a_21950_1126# a_1962_1166# a_22042_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4452 a_20946_5142# a_1962_5182# a_21038_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4453 a_30074_17190# a_2346_17232# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4454 a_15318_15222# rowon_n[13] a_14922_15182# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4455 VDD rowon_n[0] a_30986_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4456 a_31078_5142# a_2346_5184# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4457 a_34090_16186# a_2346_16228# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4458 a_5278_15222# rowon_n[13] a_4882_15182# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4459 a_30986_13174# a_1962_13214# a_31078_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4460 VSS sample_n a_1962_18234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4461 VDD VDD a_23958_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4462 a_1962_16226# sample_n VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4463 a_12002_16186# a_2346_16228# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4464 a_21438_15544# col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4465 a_9294_14218# rowon_n[12] a_8898_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4466 VSS row_n[9] a_6282_11206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4467 VSS row_n[9] a_16322_11206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4468 a_21038_11166# a_2346_11208# a_20946_11166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4469 a_18330_8194# rowon_n[6] a_17934_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4470 a_30378_8194# col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4471 VSS VDD a_5278_1166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4472 a_31382_4178# col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4473 a_19334_4178# rowon_n[2] a_18938_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4474 a_21950_11166# row_n[9] a_22442_11528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4475 VSS row_n[3] a_4274_5182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4476 VSS row_n[2] a_17326_4178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4477 vcm a_1962_8194# a_34090_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4478 VDD rowon_n[11] a_4882_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4479 VDD rowon_n[11] a_14922_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4480 a_6982_8154# a_2346_8196# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4481 VSS row_n[5] a_21342_7190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4482 a_7986_4138# a_2346_4180# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4483 a_19942_14178# row_n[12] a_20434_14540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4484 a_5278_10202# col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4485 a_15318_10202# col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4486 vcm a_1962_10202# a_20034_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4487 a_24962_7150# a_1962_7190# a_25054_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4488 a_25966_3134# a_1962_3174# a_26058_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4489 a_3970_12170# a_2346_12212# a_3878_12170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4490 a_14010_12170# a_2346_12212# a_13918_12170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4491 a_35094_7150# a_2346_7192# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4492 a_3878_6146# a_1962_6186# a_3970_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4493 a_4370_3496# col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4494 VDD rowon_n[2] a_18938_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4495 vcm a_1962_4178# a_9994_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4496 a_14314_16226# col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4497 a_15926_9158# a_1962_9198# a_16018_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4498 a_30986_4138# row_n[2] a_31478_4500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4499 a_13006_18194# a_2346_18236# a_12914_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4500 a_35094_18194# a_2346_18236# a_35002_18194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4501 a_4274_16226# col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4502 vcm a_1962_15222# a_32082_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4503 a_35398_6186# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4504 VSS row_n[1] a_9294_3174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4505 a_17422_4500# col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4506 a_2966_18194# a_2346_18236# a_2874_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4507 a_4370_12532# col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4508 a_14410_12532# col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4509 VSS sample a_2346_5184# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4510 a_13406_18556# col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4511 a_3366_18556# col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4512 VSS row_n[3] a_26362_5182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4513 a_26058_15182# a_2346_15224# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4514 a_7894_8154# a_1962_8194# a_7986_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4515 a_9390_1488# col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4516 a_8898_4138# a_1962_4178# a_8990_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4517 a_28466_8516# col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4518 VSS row_n[15] a_19334_17230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4519 a_23350_15222# rowon_n[13] a_22954_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4520 VSS row_n[10] a_20338_12210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4521 a_29982_1126# a_1962_1166# a_30074_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4522 a_13006_9158# a_2346_9200# a_12914_9158# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4523 a_11302_5182# rowon_n[3] a_10906_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4524 a_12306_1166# VSS a_11910_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4525 VSS row_n[9] a_24354_11206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4526 a_26458_3496# col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4527 VDD sample a_2346_12212# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4528 a_14314_10202# rowon_n[8] a_13918_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4529 VDD rowon_n[6] a_12914_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4530 a_4274_10202# rowon_n[8] a_3878_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4531 a_19430_15544# col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4532 VDD rowon_n[11] a_22954_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4533 a_19030_11166# a_2346_11208# a_18938_11166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4534 a_20434_10524# col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4535 a_20338_3174# col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4536 VSS row_n[1] a_30378_3174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4537 VDD rowon_n[1] a_10906_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4538 a_22346_9198# rowon_n[7] a_21950_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4539 a_4974_8154# a_2346_8196# a_4882_8154# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4540 a_5978_4138# a_2346_4180# a_5886_4138# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4541 VDD VDD a_35002_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4542 a_10298_9198# col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4543 vcm a_1962_7190# a_23046_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4544 vcm a_1962_3174# a_24050_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4545 a_16322_3174# rowon_n[1] a_15926_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4546 a_35398_15222# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4547 a_33086_7150# a_2346_7192# a_32994_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4548 a_32482_6508# col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4549 vcm a_1962_9198# a_14010_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4550 VSS row_n[13] a_12306_15222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4551 a_8898_14178# a_1962_14218# a_8990_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4552 a_18938_14178# a_1962_14218# a_19030_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4553 a_19942_1126# en_bit_n[0] a_20434_1488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4554 a_25054_2130# a_2346_2172# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4555 a_13310_11206# col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4556 a_30474_1488# col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4557 a_34490_17552# col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4558 a_30986_14178# row_n[12] a_31478_14540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4559 a_12002_13174# a_2346_13216# a_11910_13174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4560 a_34090_13174# a_2346_13216# a_33998_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4561 a_3270_11206# col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4562 vcm a_1962_10202# a_31078_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4563 VDD VSS a_15926_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4564 a_25358_1166# col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4565 VDD rowon_n[0] a_2874_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4566 a_9902_9158# row_n[7] a_10394_9520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4567 VDD rowon_n[7] a_21950_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4568 a_10906_5142# row_n[3] a_11398_5504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4569 VSS VDD a_35398_1166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4570 VDD rowon_n[15] a_10906_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4571 a_35002_13174# row_n[11] a_35494_13536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4572 a_9994_6146# a_2346_6188# a_9902_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4573 a_8290_2170# rowon_n[0] a_7894_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4574 a_3270_4178# col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4575 VSS row_n[3] a_34394_5182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4576 a_12402_13536# col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4577 a_19334_13214# rowon_n[11] a_18938_13174# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X4578 vcm a_1962_1166# a_29070_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4579 vcm a_1962_5182# a_28066_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4580 vcm a_1962_8194# a_5978_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4581 vcm a_1962_4178# a_6982_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4582 a_33998_6146# a_1962_6186# a_34090_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4583 a_34490_3496# col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4584 a_2874_4138# row_n[2] a_3366_4500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4585 VDD rowon_n[9] a_18938_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4586 a_14922_7150# row_n[5] a_15414_7512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4587 VDD rowon_n[5] a_26970_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4588 a_14010_10162# a_2346_10204# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4589 a_9902_18194# VDD a_10394_18556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4590 a_21342_16226# rowon_n[14] a_20946_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4591 a_34394_15222# rowon_n[13] a_33998_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4592 vcm a_1962_14218# a_9994_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4593 VSS row_n[10] a_31382_12210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4594 a_3970_10162# a_2346_10204# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4595 VDD rowon_n[0] a_24962_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4596 a_12914_2130# row_n[0] a_13406_2492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4597 VSS row_n[9] a_35398_11206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4598 a_24354_8194# col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4599 a_22954_15182# a_1962_15222# a_23046_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4600 a_18330_2170# col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4601 a_17022_17190# a_2346_17232# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4602 VDD rowon_n[12] a_29982_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4603 a_26058_12170# a_2346_12212# a_25966_12170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4604 a_12306_11206# rowon_n[9] a_11910_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4605 a_24050_9158# a_2346_9200# a_23958_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4606 a_6982_17190# a_2346_17232# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4607 VDD rowon_n[11] a_33998_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4608 a_26970_12170# row_n[10] a_27462_12532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4609 a_31478_10524# col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4610 a_23046_2130# a_2346_2172# a_22954_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4611 VSS row_n[2] a_10298_4178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4612 VDD rowon_n[3] a_30986_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4613 a_33390_16226# col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4614 a_29374_6186# col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4615 VSS row_n[14] a_10298_16226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4616 a_9294_17230# col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4617 a_19334_17230# col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4618 vcm a_1962_17230# a_24050_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4619 a_7286_9198# col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4620 vcm a_1962_16226# a_28066_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4621 a_32082_14178# a_2346_14220# a_31990_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4622 a_10394_4500# col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4623 a_14922_18194# a_1962_18234# a_15014_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4624 a_32482_18556# col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4625 a_4882_18194# a_1962_18234# a_4974_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4626 VSS row_n[4] a_14314_6186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4627 vcm a_1962_6186# a_32082_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4628 a_18938_15182# row_n[13] a_19430_15544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4629 vcm a_1962_11206# a_19030_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4630 a_4370_6508# col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4631 a_8898_15182# row_n[13] a_9390_15544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4632 vcm a_1962_11206# a_8990_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4633 a_6890_9158# row_n[7] a_7382_9520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4634 a_4974_6146# a_2346_6188# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4635 a_23958_1126# a_1962_1166# a_24050_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4636 a_17022_9158# a_2346_9200# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4637 a_33086_5142# a_2346_5184# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4638 a_22954_5142# a_1962_5182# a_23046_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4639 VDD rowon_n[0] a_32994_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4640 VDD sample_n a_1962_4178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4641 a_21438_8516# col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4642 VSS sample a_2346_17232# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4643 VSS row_n[10] a_29374_12210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4644 VSS VDD a_7286_1166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4645 a_16018_2130# a_2346_2172# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4646 a_33390_4178# col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4647 a_34090_11166# a_2346_11208# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4648 a_33390_10202# rowon_n[8] a_32994_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4649 a_1962_11206# sample_n VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4650 a_12002_11166# a_2346_11208# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4651 VSS VDD a_28370_18234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4652 a_32386_16226# rowon_n[14] a_31990_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4653 VDD rowon_n[12] a_27974_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4654 a_8990_8154# a_2346_8196# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4655 VSS row_n[5] a_23350_7190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4656 a_9994_4138# a_2346_4180# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4657 a_29374_14218# col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4658 a_27974_3134# a_1962_3174# a_28066_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4659 a_20946_16186# a_1962_16226# a_21038_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4660 a_33998_15182# a_1962_15222# a_34090_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4661 a_29470_10524# col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4662 a_5886_6146# a_1962_6186# a_5978_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4663 a_32994_4138# row_n[2] a_33486_4500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4664 a_4974_18194# a_2346_18236# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4665 a_15014_18194# a_2346_18236# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4666 a_17934_9158# a_1962_9198# a_18026_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4667 a_26458_6508# col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4668 a_28466_16548# col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4669 a_16930_2130# a_1962_2170# a_17022_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4670 VDD rowon_n[4] a_10906_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4671 a_8290_12210# col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4672 a_18330_12210# col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4673 vcm a_1962_12210# a_23046_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4674 VSS row_n[3] a_28370_5182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4675 VSS row_n[6] a_6282_8194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4676 a_17326_18234# col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4677 vcm a_1962_18234# a_22042_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4678 a_7286_18234# col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4679 a_2966_6146# a_2346_6188# a_2874_6146# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4680 a_7382_14540# col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4681 a_17422_14540# col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4682 a_13310_5182# rowon_n[3] a_12914_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4683 a_14314_1166# VSS a_13918_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4684 vcm a_1962_1166# a_22042_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4685 a_2346_13216# sample VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4686 a_26058_10162# a_2346_10204# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4687 a_15014_9158# a_2346_9200# a_14922_9158# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4688 a_28466_3496# col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4689 a_31078_5142# a_2346_5184# a_30986_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4690 vcm a_1962_5182# a_21038_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4691 a_7894_10162# row_n[8] a_8386_10524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4692 a_17934_10162# row_n[8] a_18426_10524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4693 VDD rowon_n[3] a_2874_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4694 a_16930_16186# row_n[14] a_17422_16548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4695 a_6890_16186# row_n[14] a_7382_16548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4696 VDD rowon_n[5] a_19942_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4697 VDD rowon_n[1] a_12914_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4698 a_26362_17230# rowon_n[15] a_25966_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4699 vcm a_1962_15222# a_15014_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4700 VSS row_n[1] a_32386_3174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4701 a_7986_4138# a_2346_4180# a_7894_4138# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4702 vcm a_1962_15222# a_4974_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4703 a_24354_9198# rowon_n[7] a_23958_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4704 a_6982_8154# a_2346_8196# a_6890_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4705 VSS row_n[11] a_27366_13214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4706 a_31382_11206# rowon_n[9] a_30986_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4707 a_24354_10202# col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4708 vcm a_1962_7190# a_25054_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4709 vcm a_1962_3174# a_26058_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4710 a_35094_7150# a_2346_7192# a_35002_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4711 vcm a_1962_6186# a_3970_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4712 a_34490_6508# col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4713 a_17326_12210# rowon_n[10] a_16930_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4714 vcm a_1962_9198# a_16018_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4715 a_7286_12210# rowon_n[10] a_6890_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4716 a_27062_2130# a_2346_2172# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4717 a_11302_2170# col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4718 VDD rowon_n[13] a_25966_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4719 a_14010_13174# a_2346_13216# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4720 a_23446_12532# col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4721 a_30986_8154# a_1962_8194# a_31078_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4722 a_32482_1488# col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4723 a_31990_4138# a_1962_4178# a_32082_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4724 a_3970_13174# a_2346_13216# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4725 VDD rowon_n[7] a_23958_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4726 VDD rowon_n[3] a_24962_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4727 a_31990_16186# a_1962_16226# a_32082_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4728 a_27462_11528# col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4729 a_12914_5142# row_n[3] a_13406_5504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4730 a_5278_4178# col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4731 a_25358_18234# col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4732 VDD rowon_n[8] a_16930_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4733 VDD rowon_n[8] a_6890_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4734 vcm a_1962_8194# a_7986_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4735 vcm a_1962_4178# a_8990_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4736 VSS row_n[15] a_5278_17230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4737 VSS row_n[15] a_15318_17230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4738 a_20034_17190# a_2346_17232# a_19942_17190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4739 a_22346_6186# col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4740 a_24050_16186# a_2346_16228# a_23958_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4741 a_16322_13214# col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4742 vcm a_1962_13214# a_21038_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4743 a_5278_7190# rowon_n[5] a_4882_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4744 vcm a_1962_1166# a_30074_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4745 a_20946_17190# row_n[15] a_21438_17552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4746 VSS row_n[14] a_9294_16226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4747 a_15014_15182# a_2346_15224# a_14922_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4748 a_6282_13214# col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4749 vcm a_1962_12210# a_34090_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4750 a_19430_7512# col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4751 a_24962_16186# row_n[14] a_25454_16548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4752 a_4974_15182# a_2346_15224# a_4882_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4753 VDD rowon_n[5] a_28978_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4754 a_4882_4138# row_n[2] a_5374_4500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4755 a_15414_15544# col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4756 a_8990_14178# a_2346_14220# a_8898_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4757 a_11910_12170# row_n[10] a_12402_12532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4758 VDD VDD a_7894_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4759 a_5374_15544# col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4760 VSS sample_n a_1962_9198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4761 VDD rowon_n[0] a_26970_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4762 a_15926_11166# row_n[9] a_16418_11528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4763 a_14922_2130# row_n[0] a_15414_2492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4764 a_5886_11166# row_n[9] a_6378_11528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4765 a_26362_8194# col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4766 a_27366_4178# col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4767 a_28066_12170# a_2346_12212# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4768 a_22954_10162# a_1962_10202# a_23046_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4769 a_31382_2170# rowon_n[0] a_30986_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4770 VSS row_n[2] a_12306_4178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4771 a_24354_18234# VDD a_23958_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4772 vcm a_1962_16226# a_2966_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4773 vcm a_1962_16226# a_13006_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4774 VSS row_n[13] a_21342_15222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4775 a_25054_2130# a_2346_2172# a_24962_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4776 a_26970_4138# row_n[2] a_27462_4500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4777 VDD rowon_n[3] a_32994_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4778 VSS row_n[12] a_25358_14218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4779 a_22346_11206# col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4780 a_1962_8194# sample_n VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4781 a_2966_4138# a_2346_4180# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4782 a_25966_17190# a_1962_17230# a_26058_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4783 a_30074_15182# a_2346_15224# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4784 a_19942_7150# a_1962_7190# a_20034_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4785 a_20946_3134# a_1962_3174# a_21038_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4786 VDD rowon_n[15] a_19942_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4787 a_15318_13214# rowon_n[11] a_14922_13174# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4788 a_9294_9198# col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4789 a_30074_7150# a_2346_7192# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4790 a_31078_3134# a_2346_3176# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4791 a_34090_14178# a_2346_14220# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4792 a_5278_13214# rowon_n[11] a_4882_13174# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4793 a_10906_9158# a_1962_9198# a_10998_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4794 VSS sample_n a_1962_16226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4795 VDD rowon_n[14] a_23958_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4796 a_1962_14218# sample_n VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4797 a_12002_14178# a_2346_14220# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4798 a_21438_13536# col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4799 a_18330_6186# rowon_n[4] a_17934_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4800 a_30378_6186# col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4801 VSS row_n[1] a_4274_3174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4802 a_12402_4500# col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4803 a_16930_12170# a_1962_12210# a_17022_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4804 a_6890_12170# a_1962_12210# a_6982_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4805 VSS row_n[10] a_14314_12210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4806 vcm a_1962_6186# a_34090_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4807 VSS row_n[10] a_4274_12210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4808 VDD rowon_n[9] a_4882_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4809 VDD rowon_n[9] a_14922_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4810 a_6982_6146# a_2346_6188# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4811 VSS row_n[3] a_21342_5182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4812 VSS VDD a_13310_18234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4813 a_19942_12170# row_n[10] a_20434_12532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4814 a_8898_9158# row_n[7] a_9390_9520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4815 a_25966_1126# a_1962_1166# a_26058_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4816 a_24962_5142# a_1962_5182# a_25054_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4817 VSS VDD a_3270_18234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4818 a_31078_17190# a_2346_17232# a_30986_17190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4819 a_3970_10162# a_2346_10204# a_3878_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4820 a_14010_10162# a_2346_10204# a_13918_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4821 a_2874_8154# a_1962_8194# a_2966_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4822 a_4370_1488# en_C0_n VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4823 a_3878_4138# a_1962_4178# a_3970_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4824 a_35094_5142# a_2346_5184# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4825 VDD rowon_n[12] a_12914_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4826 a_14314_14218# col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4827 a_23446_8516# col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4828 a_31990_17190# row_n[15] a_32482_17552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4829 a_13006_16186# a_2346_16228# a_12914_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4830 a_35094_16186# a_2346_16228# a_35002_16186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4831 VDD rowon_n[12] a_2874_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4832 a_4274_14218# col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4833 vcm a_1962_13214# a_32082_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4834 VSS VDD a_9294_1166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4835 a_35398_4178# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4836 a_2966_16186# a_2346_16228# a_2874_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4837 a_4370_10524# col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4838 a_14410_10524# col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4839 a_18026_2130# a_2346_2172# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4840 VSS sample a_2346_3176# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4841 a_21438_3496# col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4842 a_13406_16548# col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4843 a_3366_16548# col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4844 VSS row_n[5] a_25358_7190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4845 VSS row_n[1] a_26362_3174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4846 a_35398_7190# rowon_n[5] a_35002_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4847 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X4848 a_26058_13174# a_2346_13216# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4849 VSS row_n[7] a_16322_9198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4850 a_7894_6146# a_1962_6186# a_7986_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4851 a_28466_6508# col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4852 a_35002_4138# row_n[2] a_35494_4500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4853 VSS row_n[13] a_19334_15222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4854 a_23350_13214# rowon_n[11] a_22954_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4855 VSS row_n[8] a_20338_10202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4856 a_20946_11166# a_1962_11206# a_21038_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4857 a_11302_3174# rowon_n[1] a_10906_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4858 a_33998_10162# a_1962_10202# a_34090_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4859 a_26458_1488# col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4860 a_35398_18234# VDD a_35002_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4861 a_18938_2130# a_1962_2170# a_19030_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4862 VDD rowon_n[15] a_17934_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4863 a_24962_12170# a_1962_12210# a_25054_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4864 VDD rowon_n[4] a_12914_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4865 a_20034_2130# a_2346_2172# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4866 a_16418_9520# col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4867 VSS row_n[6] a_8290_8194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4868 a_23958_18194# a_1962_18234# a_24050_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4869 a_19430_13536# col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4870 VDD rowon_n[9] a_22954_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4871 VDD VSS a_10906_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4872 a_20338_1166# en_bit_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4873 VSS VDD a_30378_1166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4874 VSS row_n[15] a_34394_17230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4875 a_4974_6146# a_2346_6188# a_4882_6146# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4876 a_3270_2170# rowon_n[0] a_2874_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4877 VDD rowon_n[14] a_35002_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4878 a_17022_9158# a_2346_9200# a_16930_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4879 a_16322_1166# VSS a_15926_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4880 vcm a_1962_1166# a_24050_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4881 vcm a_1962_5182# a_23046_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4882 a_11302_17230# rowon_n[15] a_10906_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4883 a_35398_13214# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4884 a_33086_5142# a_2346_5184# a_32994_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4885 a_29070_17190# a_2346_17232# a_28978_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4886 VSS row_n[11] a_12306_13214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4887 a_30074_12170# a_2346_12212# a_29982_12170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4888 a_16018_2130# a_2346_2172# a_15926_2130# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4889 a_34490_15544# col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4890 a_30986_12170# row_n[10] a_31478_12532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4891 a_12002_11166# a_2346_11208# a_11910_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4892 a_34090_11166# a_2346_11208# a_33998_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4893 a_9902_7150# row_n[5] a_10394_7512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4894 VDD rowon_n[5] a_21950_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4895 VSS row_n[1] a_34394_3174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4896 VDD rowon_n[13] a_10906_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4897 a_35002_11166# row_n[9] a_35494_11528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4898 a_26362_9198# rowon_n[7] a_25966_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4899 a_8990_8154# a_2346_8196# a_8898_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4900 a_9994_4138# a_2346_4180# a_9902_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4901 a_12402_11528# col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4902 a_19334_11206# rowon_n[9] a_18938_11166# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X4903 VDD rowon_n[0] a_19942_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4904 vcm a_1962_3174# a_28066_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4905 vcm a_1962_6186# a_5978_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4906 a_10298_18234# col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4907 vcm a_1962_9198# a_18026_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4908 a_25358_2170# rowon_n[0] a_24962_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4909 a_13310_2170# col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4910 a_32994_8154# a_1962_8194# a_33086_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4911 a_29070_2130# a_2346_2172# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4912 a_33998_4138# a_1962_4178# a_34090_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4913 a_15318_8194# rowon_n[6] a_14922_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4914 vcm a_1962_17230# a_18026_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4915 VDD rowon_n[7] a_25966_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4916 a_14922_5142# row_n[3] a_15414_5504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4917 vcm a_1962_2170# a_17022_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4918 VDD rowon_n[3] a_26970_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4919 vcm a_1962_17230# a_7986_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4920 VDD rowon_n[6] a_4882_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4921 a_9902_16186# row_n[14] a_10394_16548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4922 a_21342_14218# rowon_n[12] a_20946_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4923 a_34394_13214# rowon_n[11] a_33998_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4924 a_27366_12210# col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4925 VSS row_n[8] a_31382_10202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4926 VDD sample a_2346_9200# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4927 a_22042_17190# a_2346_17232# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4928 a_31990_11166# a_1962_11206# a_32082_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4929 a_24354_6186# col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4930 a_22954_13174# a_1962_13214# a_23046_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4931 VDD rowon_n[15] a_28978_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4932 a_17022_15182# a_2346_15224# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4933 a_26458_14540# col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4934 VDD rowon_n[10] a_29982_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4935 a_26058_10162# a_2346_10204# a_25966_10162# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4936 a_7286_7190# rowon_n[5] a_6890_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4937 a_6982_15182# a_2346_15224# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4938 VDD rowon_n[9] a_33998_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4939 a_26970_10162# row_n[8] a_27462_10524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4940 VSS VDD a_32386_18234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4941 VDD rowon_n[0] a_28978_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4942 a_19430_2492# col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4943 a_33390_14218# col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4944 a_29374_4178# col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4945 a_27062_18194# a_2346_18236# a_26970_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4946 vcm a_1962_15222# a_24050_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4947 VSS row_n[12] a_10298_14218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4948 a_12002_9158# a_2346_9200# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4949 a_28370_8194# col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4950 a_18026_17190# a_2346_17232# a_17934_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4951 a_9294_15222# col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4952 a_19334_15222# col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4953 a_27974_18194# VDD a_28466_18556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4954 a_7986_17190# a_2346_17232# a_7894_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4955 a_10906_17190# a_1962_17230# a_10998_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4956 vcm a_1962_14218# a_28066_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4957 a_14922_16186# a_1962_16226# a_15014_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4958 a_32482_16548# col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4959 a_33390_2170# rowon_n[0] a_32994_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4960 a_10998_2130# a_2346_2172# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4961 a_4882_16186# a_1962_16226# a_4974_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4962 a_27062_2130# a_2346_2172# a_26970_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4963 VSS row_n[2] a_14314_4178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4964 a_8386_17552# col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4965 a_18426_17552# col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4966 vcm a_1962_8194# a_31078_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4967 a_17326_7190# col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4968 vcm a_1962_4178# a_32082_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4969 a_18938_13174# row_n[11] a_19430_13536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4970 a_28978_4138# row_n[2] a_29470_4500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4971 a_8898_13174# row_n[11] a_9390_13536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4972 a_3970_8154# a_2346_8196# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4973 a_6890_7150# row_n[5] a_7382_7512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4974 a_4974_4138# a_2346_4180# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4975 a_33086_3134# a_2346_3176# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4976 a_22954_3134# a_1962_3174# a_23046_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4977 a_32082_7150# a_2346_7192# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4978 a_12914_9158# a_1962_9198# a_13006_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4979 a_21438_6508# col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4980 VSS sample a_2346_15224# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4981 a_30074_10162# a_2346_10204# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4982 VSS row_n[8] a_29374_10202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4983 a_14410_4500# col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4984 vcm a_1962_18234# a_5978_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4985 vcm a_1962_18234# a_16018_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4986 a_2346_4180# sample VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4987 a_11910_2130# a_1962_2170# a_12002_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4988 VSS row_n[14] a_28370_16226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4989 a_32386_14218# rowon_n[12] a_31990_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4990 a_20034_18194# a_2346_18236# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4991 VDD rowon_n[10] a_27974_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4992 a_8990_6146# a_2346_6188# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4993 VSS row_n[3] a_23350_5182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4994 a_10998_17190# a_2346_17232# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4995 a_33086_17190# a_2346_17232# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4996 a_27974_1126# a_1962_1166# a_28066_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4997 a_20946_14178# a_1962_14218# a_21038_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4998 a_33998_13174# a_1962_13214# a_34090_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4999 a_4882_8154# a_1962_8194# a_4974_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5000 a_5886_4138# a_1962_4178# a_5978_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5001 VDD VDD a_26970_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5002 a_4974_16186# a_2346_16228# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5003 a_15014_16186# a_2346_16228# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5004 a_25454_8516# col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5005 VDD rowon_n[6] a_35002_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5006 a_23446_3496# col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5007 a_22954_14178# row_n[12] a_23446_14540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5008 a_8290_10202# col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5009 a_18330_10202# col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5010 vcm a_1962_10202# a_23046_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5011 a_32386_9198# col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5012 VSS row_n[5] a_27366_7190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5013 VSS row_n[1] a_28370_3174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5014 a_6982_12170# a_2346_12212# a_6890_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5015 a_9902_12170# a_1962_12210# a_9994_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5016 a_17022_12170# a_2346_12212# a_16930_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5017 VSS row_n[4] a_6282_6186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5018 a_17326_16226# col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5019 vcm a_1962_16226# a_22042_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5020 VSS row_n[7] a_18330_9198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5021 a_16018_18194# a_2346_18236# a_15926_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5022 a_7286_16226# col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5023 a_2966_4138# a_2346_4180# a_2874_4138# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5024 a_5978_18194# a_2346_18236# a_5886_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5025 a_7382_12532# col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5026 a_17422_12532# col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5027 a_13310_3174# rowon_n[1] a_12914_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5028 a_2346_11208# sample VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5029 vcm a_1962_7190# a_20034_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5030 a_28466_1488# col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5031 a_31078_3134# a_2346_3176# a_30986_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5032 vcm a_1962_3174# a_21038_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5033 a_16418_18556# col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5034 a_26970_8154# a_1962_8194# a_27062_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5035 a_30074_7150# a_2346_7192# a_29982_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5036 a_6378_18556# col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5037 vcm a_1962_9198# a_10998_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5038 a_31990_9158# row_n[7] a_32482_9520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5039 a_22042_2130# a_2346_2172# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5040 a_18426_9520# col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5041 VDD VSS a_12914_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5042 VDD rowon_n[3] a_19942_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5043 a_14922_17190# row_n[15] a_15414_17552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5044 a_26362_15222# rowon_n[13] a_25966_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5045 vcm a_1962_13214# a_15014_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5046 VSS row_n[10] a_23350_12210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5047 VSS VDD a_32386_1166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5048 a_4882_17190# row_n[15] a_5374_17552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5049 vcm a_1962_13214# a_4974_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5050 a_6982_6146# a_2346_6188# a_6890_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5051 vcm a_1962_1166# a_26058_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5052 VSS row_n[9] a_27366_11206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5053 vcm a_1962_5182# a_25054_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5054 vcm a_1962_8194# a_2966_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5055 vcm a_1962_4178# a_3970_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5056 a_35094_5142# a_2346_5184# a_35002_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5057 VDD rowon_n[12] a_21950_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5058 a_32082_12170# a_2346_12212# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5059 a_17326_10202# rowon_n[8] a_16930_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5060 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X5061 a_7286_10202# rowon_n[8] a_6890_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5062 a_18026_2130# a_2346_2172# a_17934_2130# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5063 a_31078_18194# a_2346_18236# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5064 VDD rowon_n[11] a_25966_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5065 a_23446_10524# col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5066 a_30986_6146# a_1962_6186# a_31078_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5067 VDD rowon_n[5] a_23958_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5068 a_21342_17230# col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5069 a_31990_14178# a_1962_14218# a_32082_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5070 a_25358_16226# col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5071 a_28370_9198# rowon_n[7] a_27974_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5072 VDD rowon_n[0] a_21950_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5073 a_29982_17190# a_1962_17230# a_30074_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5074 vcm a_1962_6186# a_7986_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5075 a_9902_2130# row_n[0] a_10394_2492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5076 a_8290_18234# VDD a_7894_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5077 VSS row_n[13] a_5278_15222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5078 VSS row_n[13] a_15318_15222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5079 a_20034_15182# a_2346_15224# a_19942_15182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5080 a_12306_12210# col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5081 a_21342_8194# col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5082 a_27366_2170# rowon_n[0] a_26970_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5083 a_22346_4178# col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5084 a_24450_18556# col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5085 a_24050_14178# a_2346_14220# a_23958_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5086 a_16322_11206# col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5087 vcm a_1962_11206# a_21038_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5088 VSS row_n[6] a_31382_8194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5089 a_5278_5182# rowon_n[3] a_4882_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5090 a_15318_2170# col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5091 a_20946_15182# row_n[13] a_21438_15544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5092 VSS row_n[12] a_9294_14218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5093 a_33998_14178# row_n[12] a_34490_14540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5094 a_15014_13174# a_2346_13216# a_14922_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5095 a_6282_11206# col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5096 vcm a_1962_10202# a_34090_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5097 a_17326_8194# rowon_n[6] a_16930_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5098 a_35002_8154# a_1962_8194# a_35094_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5099 a_19430_5504# col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5100 a_4974_13174# a_2346_13216# a_4882_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5101 VDD rowon_n[7] a_27974_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5102 vcm a_1962_2170# a_19030_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5103 VDD rowon_n[3] a_28978_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5104 VDD rowon_n[15] a_3878_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5105 VDD rowon_n[15] a_13918_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5106 a_11398_14540# col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5107 VDD rowon_n[6] a_6890_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5108 a_15414_13536# col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5109 a_11910_10162# row_n[8] a_12402_10524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5110 a_20034_2130# a_2346_2172# a_19942_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5111 VDD rowon_n[14] a_7894_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5112 a_5374_13536# col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5113 a_26058_7150# a_2346_7192# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5114 a_21950_4138# row_n[2] a_22442_4500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5115 VDD rowon_n[1] a_4882_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5116 a_26362_6186# col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5117 vcm a_1962_18234# a_35094_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5118 a_4274_9198# col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5119 a_9294_7190# rowon_n[5] a_8898_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5120 a_20338_17230# rowon_n[15] a_19942_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5121 a_17022_10162# a_2346_10204# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5122 a_2874_18194# VDD a_3366_18556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5123 a_12914_18194# VDD a_13406_18556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5124 a_24354_16226# rowon_n[14] a_23958_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5125 vcm a_1962_14218# a_2966_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5126 vcm a_1962_14218# a_13006_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5127 VSS row_n[11] a_21342_13214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5128 a_6982_10162# a_2346_10204# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5129 a_2346_17232# sample VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5130 a_1962_6186# sample_n VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5131 a_29070_18194# a_2346_18236# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5132 a_25966_15182# a_1962_15222# a_26058_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5133 a_30074_13174# a_2346_13216# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5134 a_3878_9158# row_n[7] a_4370_9520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5135 a_14010_9158# a_2346_9200# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5136 a_20946_1126# a_1962_1166# a_21038_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5137 a_19942_5142# a_1962_5182# a_20034_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5138 VDD rowon_n[13] a_19942_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5139 a_5278_11206# rowon_n[9] a_4882_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5140 a_15318_11206# rowon_n[9] a_14922_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5141 a_16930_8154# row_n[6] a_17422_8516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5142 a_31078_1126# a_2346_1168# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5143 a_30074_5142# a_2346_5184# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5144 a_9994_17190# a_2346_17232# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5145 a_20338_12210# col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5146 VSS sample_n a_1962_14218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5147 a_21438_11528# col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5148 VSS en_C0_n a_4274_1166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5149 a_30378_4178# col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5150 a_18330_4178# rowon_n[2] a_17934_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5151 a_13006_2130# a_2346_2172# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5152 a_32386_17230# col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5153 a_29070_2130# a_2346_2172# a_28978_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5154 VSS row_n[8] a_14314_10202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5155 vcm a_1962_8194# a_33086_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5156 a_19334_7190# col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5157 vcm a_1962_4178# a_34090_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5158 a_4882_11166# a_1962_11206# a_4974_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5159 a_14922_11166# a_1962_11206# a_15014_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5160 VSS row_n[8] a_4274_10202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5161 VSS row_n[5] a_20338_7190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5162 VSS row_n[1] a_21342_3174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5163 a_6982_4138# a_2346_4180# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5164 VSS row_n[14] a_13310_16226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5165 a_19942_10162# row_n[8] a_20434_10524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5166 a_8898_7150# row_n[5] a_9390_7512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5167 a_30378_7190# rowon_n[5] a_29982_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5168 a_24962_3134# a_1962_3174# a_25054_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5169 vcm a_1962_17230# a_27062_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5170 VSS row_n[14] a_3270_16226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5171 a_31078_15182# a_2346_15224# a_30986_15182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5172 VSS row_n[7] a_11302_9198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5173 a_34090_7150# a_2346_7192# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5174 a_2874_6146# a_1962_6186# a_2966_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5175 a_35094_3134# a_2346_3176# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5176 VDD rowon_n[10] a_12914_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5177 a_23446_6508# col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5178 a_6890_2130# row_n[0] a_7382_2492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5179 a_29982_4138# row_n[2] a_30474_4500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5180 VDD rowon_n[2] a_17934_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5181 a_35494_18556# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5182 a_31990_15182# row_n[13] a_32482_15544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5183 a_13006_14178# a_2346_14220# a_12914_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5184 a_35094_14178# a_2346_14220# a_35002_14178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5185 VDD rowon_n[10] a_2874_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5186 vcm a_1962_11206# a_32082_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5187 a_14922_9158# a_1962_9198# a_15014_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5188 VSS sample a_2346_1168# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5189 a_7894_18194# a_1962_18234# a_7986_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5190 VDD VDD a_11910_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5191 a_17934_18194# a_1962_18234# a_18026_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5192 a_2966_14178# a_2346_14220# a_2874_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5193 a_21438_1488# col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5194 a_13918_2130# a_1962_2170# a_14010_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5195 VSS VDD a_26362_1166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5196 VSS row_n[3] a_25358_5182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5197 a_11398_9520# col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5198 VSS row_n[6] a_3270_8194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5199 a_35398_5182# rowon_n[3] a_35002_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5200 a_18330_17230# rowon_n[15] a_17934_17190# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X5201 a_7894_4138# a_1962_4178# a_7986_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5202 a_27462_8516# col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5203 VSS row_n[11] a_19334_13214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5204 a_23350_11206# rowon_n[9] a_22954_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5205 a_12002_9158# a_2346_9200# a_11910_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5206 a_11302_1166# VSS a_10906_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5207 a_4974_11166# a_2346_11208# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5208 a_15014_11166# a_2346_11208# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5209 a_25454_3496# col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5210 a_35398_16226# rowon_n[14] a_35002_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5211 VDD rowon_n[1] a_35002_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5212 VDD rowon_n[13] a_17934_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5213 a_10998_2130# a_2346_2172# a_10906_2130# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5214 a_8990_12170# a_2346_12212# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5215 a_34394_9198# col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5216 a_16418_7512# col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5217 VSS row_n[5] a_29374_7190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5218 VSS row_n[4] a_8290_6186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5219 a_23958_16186# a_1962_16226# a_24050_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5220 a_19430_11528# col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5221 a_7986_18194# a_2346_18236# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5222 a_18026_18194# a_2346_18236# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5223 VSS row_n[13] a_34394_15222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5224 a_31382_12210# col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5225 a_21342_9198# rowon_n[7] a_20946_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5226 a_3970_8154# a_2346_8196# a_3878_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5227 a_4974_4138# a_2346_4180# a_4882_4138# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5228 vcm a_1962_3174# a_23046_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5229 a_11302_15222# rowon_n[13] a_10906_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5230 a_35398_11206# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5231 a_28978_8154# a_1962_8194# a_29070_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5232 a_32082_7150# a_2346_7192# a_31990_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5233 a_33086_3134# a_2346_3176# a_32994_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5234 vcm a_1962_9198# a_13006_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5235 a_20338_2170# rowon_n[0] a_19942_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5236 VDD rowon_n[15] a_32994_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5237 a_29070_15182# a_2346_15224# a_28978_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5238 a_30474_14540# col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5239 vcm a_1962_12210# a_26058_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5240 VSS row_n[9] a_12306_11206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5241 a_30074_10162# a_2346_10204# a_29982_10162# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5242 a_33998_9158# row_n[7] a_34490_9520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5243 a_24050_2130# a_2346_2172# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5244 a_34490_13536# col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5245 a_30986_10162# row_n[8] a_31478_10524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5246 a_10298_8194# rowon_n[6] a_9902_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5247 VDD rowon_n[3] a_21950_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5248 VDD rowon_n[7] a_20946_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5249 a_9902_5142# row_n[3] a_10394_5504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5250 vcm a_1962_2170# a_12002_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5251 VDD rowon_n[11] a_10906_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5252 a_8990_6146# a_2346_6188# a_8898_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5253 vcm a_1962_1166# a_28066_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5254 vcm a_1962_8194# a_4974_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5255 vcm a_1962_4178# a_5978_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5256 a_10298_16226# col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5257 a_32994_6146# a_1962_6186# a_33086_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5258 a_15318_6186# rowon_n[4] a_14922_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5259 a_29374_17230# rowon_n[15] a_28978_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5260 vcm a_1962_15222# a_18026_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5261 VDD rowon_n[5] a_25966_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5262 vcm a_1962_15222# a_7986_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5263 a_30378_12210# rowon_n[10] a_29982_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5264 VDD rowon_n[4] a_4882_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5265 a_34394_11206# rowon_n[9] a_33998_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5266 a_27366_10202# col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5267 VDD sample a_2346_7192# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5268 VDD rowon_n[0] a_23958_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5269 a_22042_15182# a_2346_15224# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5270 VSS row_n[0] a_19334_2170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5271 a_24354_4178# col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5272 a_23350_8194# col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5273 VSS row_n[6] a_33390_8194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5274 a_29374_2170# rowon_n[0] a_28978_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5275 VDD rowon_n[13] a_28978_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5276 a_17022_13174# a_2346_13216# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5277 a_26458_12532# col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5278 VDD rowon_n[8] a_29982_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5279 a_7286_5182# rowon_n[3] a_6890_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5280 a_6982_13174# a_2346_13216# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5281 vcm a_1962_8194# a_27062_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5282 VDD rowon_n[6] a_8898_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5283 a_22042_2130# a_2346_2172# a_21950_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5284 a_28370_18234# col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5285 VSS row_n[14] a_32386_16226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5286 a_12306_7190# col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5287 a_28066_7150# a_2346_7192# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5288 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X5289 VDD rowon_n[1] a_6890_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5290 a_23958_4138# row_n[2] a_24450_4500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5291 VSS row_n[15] a_8290_17230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5292 VSS row_n[15] a_18330_17230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5293 a_23046_17190# a_2346_17232# a_22954_17190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5294 a_27062_16186# a_2346_16228# a_26970_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5295 vcm a_1962_13214# a_24050_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5296 a_28370_6186# col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5297 VDD VDD a_30986_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5298 a_23958_17190# row_n[15] a_24450_17552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5299 a_18026_15182# a_2346_15224# a_17934_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5300 a_9294_13214# col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5301 a_19334_13214# col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5302 a_6282_9198# col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5303 a_27974_16186# row_n[14] a_28466_16548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5304 a_7986_15182# a_2346_15224# a_7894_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5305 a_10906_15182# a_1962_15222# a_10998_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5306 a_14922_14178# a_1962_14218# a_15014_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5307 a_4882_14178# a_1962_14218# a_4974_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5308 a_8386_15544# col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5309 a_18426_15544# col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5310 vcm a_1962_6186# a_31078_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5311 a_17326_5182# col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5312 a_18938_11166# row_n[9] a_19430_11528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5313 a_8898_11166# row_n[9] a_9390_11528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5314 a_5886_9158# row_n[7] a_6378_9520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5315 a_3970_6146# a_2346_6188# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5316 a_6890_5142# row_n[3] a_7382_5504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5317 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.64e+07u l=1.6e+07u
X5318 a_18938_8154# row_n[6] a_19430_8516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5319 a_22954_1126# a_1962_1166# a_23046_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5320 a_33086_1126# a_2346_1168# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5321 a_32082_5142# a_2346_5184# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5322 vcm a_1962_17230# a_12002_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5323 a_28370_12210# rowon_n[10] a_27974_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5324 a_25966_10162# a_1962_10202# a_26058_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5325 a_20434_8516# col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5326 VSS sample a_2346_13216# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5327 VDD rowon_n[6] a_29982_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5328 a_15014_2130# a_2346_2172# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5329 a_16930_3134# row_n[1] a_17422_3496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5330 a_27366_18234# VDD a_26970_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5331 vcm a_1962_16226# a_5978_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5332 vcm a_1962_16226# a_16018_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5333 a_2346_2172# sample VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5334 vcm a_1962_8194# a_35094_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5335 VSS row_n[12] a_28370_14218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5336 a_28978_17190# a_1962_17230# a_29070_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5337 a_20034_16186# a_2346_16228# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5338 VDD rowon_n[8] a_27974_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5339 VSS row_n[5] a_22346_7190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5340 VSS row_n[1] a_23350_3174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5341 a_8990_4138# a_2346_4180# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5342 a_10998_15182# a_2346_15224# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5343 a_33086_15182# a_2346_15224# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5344 a_32386_7190# rowon_n[5] a_31990_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5345 VSS row_n[7] a_13310_9198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5346 a_19030_9158# a_2346_9200# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5347 a_26058_7150# a_2346_7192# a_25966_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5348 a_4882_6146# a_1962_6186# a_4974_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5349 VDD rowon_n[14] a_26970_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5350 a_4974_14178# a_2346_14220# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5351 a_15014_14178# a_2346_14220# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5352 a_25454_6508# col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5353 a_8898_2130# row_n[0] a_9390_2492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5354 VDD rowon_n[4] a_35002_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5355 a_23446_1488# col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5356 VSS row_n[10] a_17326_12210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5357 a_22042_12170# a_2346_12212# a_21950_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5358 a_21950_8154# a_1962_8194# a_22042_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5359 a_15926_2130# a_1962_2170# a_16018_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5360 VSS row_n[10] a_7286_12210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5361 VSS VDD a_16322_18234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5362 a_21038_18194# a_2346_18236# a_20946_18194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5363 a_22954_12170# row_n[10] a_23446_12532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5364 VSS VDD a_28370_1166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5365 VSS row_n[3] a_27366_5182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5366 VSS VDD a_6282_18234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5367 a_6982_10162# a_2346_10204# a_6890_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5368 a_17022_10162# a_2346_10204# a_16930_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5369 a_13406_9520# col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5370 VSS row_n[6] a_5278_8194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5371 VSS row_n[2] a_6282_4178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5372 a_21950_18194# VDD a_22442_18556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5373 VDD rowon_n[12] a_15926_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5374 a_17326_14218# col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5375 vcm a_1962_14218# a_22042_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5376 a_16018_16186# a_2346_16228# a_15926_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5377 VDD rowon_n[12] a_5886_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5378 a_7286_14218# col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5379 a_29470_8516# col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5380 a_5978_16186# a_2346_16228# a_5886_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5381 a_7382_10524# col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5382 a_17422_10524# col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5383 a_13310_1166# VSS a_12914_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5384 vcm a_1962_1166# a_21038_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5385 a_15318_17230# col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5386 vcm a_1962_17230# a_20034_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5387 a_14010_9158# a_2346_9200# a_13918_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5388 a_31078_1126# a_2346_1168# a_30986_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5389 vcm a_1962_5182# a_20034_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5390 a_5278_17230# col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5391 a_16418_16548# col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5392 a_26970_6146# a_1962_6186# a_27062_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5393 a_27462_3496# col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5394 a_30074_5142# a_2346_5184# a_29982_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5395 a_6378_16548# col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5396 a_31990_7150# row_n[5] a_32482_7512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5397 a_6378_4500# col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5398 a_13006_2130# a_2346_2172# a_12914_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5399 vcm a_1962_12210# a_10998_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5400 a_18426_7512# col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5401 a_14922_15182# row_n[13] a_15414_15544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5402 a_26362_13214# rowon_n[11] a_25966_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5403 vcm a_1962_11206# a_15014_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5404 VSS row_n[8] a_23350_10202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5405 a_16418_2492# col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5406 a_4882_15182# row_n[13] a_5374_15544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5407 vcm a_1962_11206# a_4974_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5408 a_23958_11166# a_1962_11206# a_24050_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5409 a_23350_9198# rowon_n[7] a_22954_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5410 a_6982_4138# a_2346_4180# a_6890_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5411 a_35094_3134# a_2346_3176# a_35002_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5412 vcm a_1962_3174# a_25054_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5413 a_34090_7150# a_2346_7192# a_33998_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5414 vcm a_1962_6186# a_2966_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5415 VDD rowon_n[10] a_21950_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5416 a_27974_12170# a_1962_12210# a_28066_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5417 vcm a_1962_9198# a_15014_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5418 a_22346_2170# rowon_n[0] a_21950_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5419 a_10298_2170# col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5420 a_26970_18194# a_1962_18234# a_27062_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5421 a_31078_16186# a_2346_16228# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5422 VDD rowon_n[9] a_25966_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5423 a_12306_8194# rowon_n[6] a_11910_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5424 a_29982_8154# a_1962_8194# a_30074_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5425 a_30986_4138# a_1962_4178# a_31078_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5426 VDD rowon_n[7] a_22954_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5427 vcm a_1962_2170# a_14010_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5428 VDD rowon_n[3] a_23958_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5429 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.64e+07u l=1.6e+07u
X5430 VSS VDD a_24354_18234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5431 a_21342_15222# col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5432 a_25358_14218# col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5433 a_14314_17230# rowon_n[15] a_13918_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5434 a_21038_7150# a_2346_7192# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5435 a_19030_18194# a_2346_18236# a_18938_18194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5436 a_4274_17230# rowon_n[15] a_3878_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5437 a_29982_15182# a_1962_15222# a_30074_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5438 vcm a_1962_4178# a_7986_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5439 a_20434_17552# col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5440 a_8290_16226# rowon_n[14] a_7894_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5441 VSS row_n[11] a_5278_13214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5442 VSS row_n[11] a_15318_13214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5443 a_20034_13174# a_2346_13216# a_19942_13174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5444 a_33086_12170# a_2346_12212# a_32994_12170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5445 a_12306_10202# col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5446 a_21342_6186# col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5447 a_24450_16548# col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5448 a_20946_13174# row_n[11] a_21438_13536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5449 a_10998_12170# a_2346_12212# a_10906_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5450 a_4274_7190# rowon_n[5] a_3878_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5451 VSS row_n[4] a_31382_6186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5452 a_5278_3174# rowon_n[1] a_4882_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5453 a_33998_12170# row_n[10] a_34490_12532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5454 a_15014_11166# a_2346_11208# a_14922_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5455 a_17326_6186# rowon_n[4] a_16930_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5456 a_35002_6146# a_1962_6186# a_35094_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5457 a_4974_11166# a_2346_11208# a_4882_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5458 VDD rowon_n[5] a_27974_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5459 VDD rowon_n[13] a_3878_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5460 VDD rowon_n[13] a_13918_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5461 a_11398_12532# col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5462 VDD rowon_n[4] a_6890_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5463 a_15414_11528# col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5464 a_5374_11528# col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5465 VDD rowon_n[0] a_25966_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5466 a_26058_5142# a_2346_5184# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5467 a_13310_18234# col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5468 VDD VSS a_4882_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5469 a_3270_18234# col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5470 vcm a_1962_17230# a_31078_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5471 a_25358_8194# col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5472 a_26362_4178# col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5473 vcm a_1962_16226# a_35094_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5474 a_11910_8154# row_n[6] a_12402_8516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5475 VSS row_n[6] a_35398_8194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5476 a_2346_7192# sample VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5477 a_9294_5182# rowon_n[3] a_8898_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5478 a_22042_10162# a_2346_10204# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5479 a_20338_15222# rowon_n[13] a_19942_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5480 vcm a_1962_8194# a_29070_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5481 a_2874_16186# row_n[14] a_3366_16548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5482 a_12914_16186# row_n[14] a_13406_16548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5483 a_24354_14218# rowon_n[12] a_23958_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5484 VSS row_n[9] a_21342_11206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5485 a_24050_2130# a_2346_2172# a_23958_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5486 a_25054_17190# a_2346_17232# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5487 a_2346_15224# sample VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5488 a_14314_7190# col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5489 VDD rowon_n[1] a_8898_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5490 a_25966_4138# row_n[2] a_26458_4500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5491 a_1962_4178# sample_n VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5492 a_29070_16186# a_2346_16228# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5493 a_25966_13174# a_1962_13214# a_26058_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5494 a_3878_7150# row_n[5] a_4370_7512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5495 a_19942_3134# a_1962_3174# a_20034_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5496 VDD VDD a_18938_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5497 VDD rowon_n[11] a_19942_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5498 a_8290_9198# col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5499 a_16930_6146# row_n[4] a_17422_6508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5500 a_30074_3134# a_2346_3176# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5501 a_9994_15182# a_2346_15224# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5502 a_20338_10202# col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5503 a_9902_9158# a_1962_9198# a_9994_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5504 a_13310_12210# rowon_n[10] a_12914_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5505 VSS VDD a_35398_18234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5506 a_32386_15222# col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5507 a_3270_12210# rowon_n[10] a_2874_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5508 a_10906_10162# a_1962_10202# a_10998_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5509 a_7286_2170# col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5510 vcm a_1962_6186# a_33086_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5511 a_19334_5182# col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5512 a_12306_18234# VDD a_11910_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5513 VSS VDD a_21342_1166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5514 VSS row_n[3] a_20338_5182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5515 VSS row_n[12] a_13310_14218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5516 a_7894_9158# row_n[7] a_8386_9520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5517 a_8898_5142# row_n[3] a_9390_5504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5518 a_24962_1126# a_1962_1166# a_25054_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5519 a_30378_5182# rowon_n[3] a_29982_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5520 a_31478_17552# col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5521 vcm a_1962_15222# a_27062_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5522 VSS row_n[12] a_3270_14218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5523 a_31078_13174# a_2346_13216# a_30986_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5524 a_35094_1126# a_2346_1168# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5525 a_2874_4138# a_1962_4178# a_2966_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5526 a_34090_5142# a_2346_5184# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5527 a_3878_17190# a_1962_17230# a_3970_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5528 a_13918_17190# a_1962_17230# a_14010_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5529 VDD rowon_n[8] a_12914_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5530 a_22442_8516# col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5531 a_35494_16548# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5532 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.64e+07u l=1.6e+07u
X5533 a_31990_13174# row_n[11] a_32482_13536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5534 VDD rowon_n[8] a_2874_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5535 VDD rowon_n[6] a_31990_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5536 a_18938_3134# row_n[1] a_19430_3496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5537 a_7894_16186# a_1962_16226# a_7986_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5538 VDD rowon_n[14] a_11910_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5539 a_17934_16186# a_1962_16226# a_18026_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5540 a_17022_2130# a_2346_2172# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5541 a_20434_3496# col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5542 vcm a_1962_12210# a_30074_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5543 VDD rowon_n[1] a_29982_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5544 VSS row_n[1] a_25358_3174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5545 a_11398_7512# col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5546 VSS row_n[5] a_24354_7190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5547 a_34394_7190# rowon_n[5] a_33998_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5548 VSS row_n[4] a_3270_6186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5549 a_35398_3174# rowon_n[1] a_35002_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5550 a_18330_15222# rowon_n[13] a_17934_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5551 a_20034_11166# a_2346_11208# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5552 VSS row_n[7] a_15318_9198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5553 a_28066_7150# a_2346_7192# a_27974_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5554 a_27462_6508# col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5555 VSS row_n[9] a_19334_11206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5556 a_10998_10162# a_2346_10204# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5557 a_33086_10162# a_2346_10204# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5558 vcm a_1962_18234# a_19030_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5559 a_5978_9158# a_2346_9200# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5560 vcm a_1962_18234# a_8990_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5561 a_24050_12170# a_2346_12212# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5562 a_23958_8154# a_1962_8194# a_24050_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5563 a_25454_1488# col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5564 a_35398_14218# rowon_n[12] a_35002_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5565 VDD VSS a_35002_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5566 analog_in sw_n ctop VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.9e+06u l=220000u
X5567 a_17934_2130# a_1962_2170# a_18026_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5568 a_23046_18194# a_2346_18236# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5569 VDD rowon_n[11] a_17934_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5570 VSS row_n[3] a_29374_5182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5571 a_15414_9520# col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5572 a_16418_5504# col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5573 VSS row_n[2] a_8290_4178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5574 a_33390_17230# rowon_n[15] a_32994_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5575 a_23958_14178# a_1962_14218# a_24050_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5576 VSS row_n[6] a_7286_8194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5577 a_7986_16186# a_2346_16228# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5578 a_18026_16186# a_2346_16228# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5579 VSS row_n[11] a_34394_13214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5580 a_31382_10202# col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5581 a_3970_6146# a_2346_6188# a_3878_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5582 vcm a_1962_1166# a_23046_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5583 a_11302_13214# rowon_n[11] a_10906_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5584 a_28978_6146# a_1962_6186# a_29070_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5585 a_33086_1126# a_2346_1168# a_32994_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5586 a_29470_3496# col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5587 a_32082_5142# a_2346_5184# a_31990_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5588 a_6890_9158# a_1962_9198# a_6982_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5589 a_29470_17552# col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5590 VDD rowon_n[13] a_32994_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5591 a_25966_14178# row_n[12] a_26458_14540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5592 a_29070_13174# a_2346_13216# a_28978_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5593 a_30474_12532# col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5594 vcm a_1962_10202# a_26058_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5595 a_33998_7150# row_n[5] a_34490_7512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5596 a_8386_4500# col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5597 a_9994_12170# a_2346_12212# a_9902_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5598 a_12914_12170# a_1962_12210# a_13006_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5599 a_15014_2130# a_2346_2172# a_14922_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5600 a_2874_12170# a_1962_12210# a_2966_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5601 a_34490_11528# col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5602 a_10298_6186# rowon_n[4] a_9902_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5603 a_31990_2130# row_n[0] a_32482_2492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5604 a_11910_18194# a_1962_18234# a_12002_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5605 VDD rowon_n[9] a_10906_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5606 VDD rowon_n[5] a_20946_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5607 VDD sample_n a_1962_18234# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5608 a_18426_2492# col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5609 a_8990_4138# a_2346_4180# a_8898_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5610 a_19030_9158# a_2346_9200# a_18938_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5611 vcm a_1962_6186# a_4974_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5612 a_10298_14218# col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5613 a_24354_2170# rowon_n[0] a_23958_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5614 a_32994_4138# a_1962_4178# a_33086_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5615 a_14314_8194# rowon_n[6] a_13918_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5616 vcm a_1962_8194# a_22042_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5617 a_15318_4178# rowon_n[2] a_14922_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5618 a_17934_17190# row_n[15] a_18426_17552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5619 a_29374_15222# rowon_n[13] a_28978_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5620 vcm a_1962_13214# a_18026_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5621 VSS row_n[10] a_26362_12210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5622 vcm a_1962_2170# a_16018_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5623 VDD rowon_n[3] a_25966_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5624 a_7894_17190# row_n[15] a_8386_17552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5625 vcm a_1962_13214# a_7986_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5626 a_31078_11166# a_2346_11208# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5627 a_30378_10202# rowon_n[8] a_29982_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5628 a_1962_9198# sample_n VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5629 VDD rowon_n[6] a_3878_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5630 VDD sample a_2346_5184# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5631 a_22042_13174# a_2346_13216# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5632 a_23046_7150# a_2346_7192# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5633 VDD rowon_n[12] a_24962_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5634 a_13006_12170# a_2346_12212# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5635 a_35094_12170# a_2346_12212# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5636 a_2966_12170# a_2346_12212# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5637 a_23350_6186# col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5638 VSS row_n[4] a_33390_6186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5639 VDD rowon_n[2] a_14922_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5640 VDD rowon_n[11] a_28978_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5641 a_26458_10524# col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5642 a_29982_10162# a_1962_10202# a_30074_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5643 a_6282_7190# rowon_n[5] a_5886_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5644 a_7286_3174# rowon_n[1] a_6890_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5645 vcm a_1962_6186# a_27062_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5646 a_31382_18234# VDD a_30986_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5647 a_24354_17230# col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5648 VDD rowon_n[4] a_8898_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5649 a_28370_16226# col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5650 VSS row_n[12] a_32386_14218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5651 a_12306_5182# col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5652 VDD rowon_n[0] a_27974_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5653 a_28066_5142# a_2346_5184# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5654 a_19942_18194# a_1962_18234# a_20034_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5655 a_32994_17190# a_1962_17230# a_33086_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5656 VDD VSS a_6890_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5657 VSS row_n[13] a_8290_15222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5658 VSS row_n[13] a_18330_15222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5659 a_23046_15182# a_2346_15224# a_22954_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5660 a_27062_14178# a_2346_14220# a_26970_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5661 a_19334_11206# col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5662 vcm a_1962_11206# a_24050_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5663 a_13918_8154# row_n[6] a_14410_8516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5664 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X5665 a_28370_4178# col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5666 a_27462_18556# col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5667 VDD rowon_n[14] a_30986_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5668 a_23958_15182# row_n[13] a_24450_15544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5669 a_18026_13174# a_2346_13216# a_17934_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5670 a_9294_11206# col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5671 VSS sample_n a_1962_2170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5672 a_7986_13174# a_2346_13216# a_7894_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5673 a_10906_13174# a_1962_13214# a_10998_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5674 VDD rowon_n[15] a_6890_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5675 VDD rowon_n[15] a_16930_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5676 a_11910_3134# row_n[1] a_12402_3496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5677 a_18426_13536# col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5678 a_8386_13536# col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5679 vcm a_1962_8194# a_30074_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5680 a_16322_7190# col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5681 a_17326_3174# col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5682 vcm a_1962_4178# a_31078_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5683 ctop sw ctop VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.9e+06u l=220000u
X5684 a_27974_4138# row_n[2] a_28466_4500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5685 a_5886_7150# row_n[5] a_6378_7512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5686 a_3970_4138# a_2346_4180# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5687 a_18938_6146# row_n[4] a_19430_6508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5688 a_2346_10204# sample VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5689 a_21038_7150# a_2346_7192# a_20946_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5690 a_32082_3134# a_2346_3176# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5691 vcm a_1962_15222# a_12002_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5692 a_29070_11166# a_2346_11208# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5693 a_28370_10202# rowon_n[8] a_27974_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5694 a_20434_6508# col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5695 a_3878_2130# row_n[0] a_4370_2492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5696 VSS sample a_2346_11208# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5697 VDD rowon_n[4] a_29982_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5698 a_16930_1126# VDD a_17422_1488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5699 a_15926_18194# VDD a_16418_18556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5700 a_27366_16226# rowon_n[14] a_26970_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5701 vcm a_1962_14218# a_5978_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5702 vcm a_1962_14218# a_16018_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5703 a_9994_10162# a_2346_10204# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5704 a_9294_2170# col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5705 a_5886_18194# VDD a_6378_18556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5706 vcm a_1962_6186# a_35094_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5707 a_10906_2130# a_1962_2170# a_10998_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5708 a_28978_15182# a_1962_15222# a_29070_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5709 a_20034_14178# a_2346_14220# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5710 VSS VDD a_23350_1166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5711 VSS row_n[3] a_22346_5182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5712 a_10998_13174# a_2346_13216# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5713 a_33086_13174# a_2346_13216# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5714 a_32386_5182# rowon_n[3] a_31990_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5715 a_23350_12210# col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5716 a_4882_4138# a_1962_4178# a_4974_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5717 a_26058_5142# a_2346_5184# a_25966_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5718 a_24450_8516# col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5719 a_22346_18234# col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5720 VDD rowon_n[6] a_33998_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5721 a_22442_14540# col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5722 VSS row_n[8] a_17326_10202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5723 a_22042_10162# a_2346_10204# a_21950_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5724 a_21950_6146# a_1962_6186# a_22042_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5725 VDD rowon_n[1] a_31990_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5726 a_22442_3496# col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5727 a_7894_11166# a_1962_11206# a_7986_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5728 a_17934_11166# a_1962_11206# a_18026_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5729 VSS row_n[8] a_7286_10202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5730 a_30986_18194# a_1962_18234# a_31078_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5731 VSS row_n[14] a_16322_16226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5732 a_21038_16186# a_2346_16228# a_20946_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5733 a_22954_10162# row_n[8] a_23446_10524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5734 VSS row_n[1] a_27366_3174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5735 VSS row_n[14] a_6282_16226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5736 a_19334_9198# rowon_n[7] a_18938_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5737 a_31382_9198# col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5738 a_13406_7512# col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5739 VSS row_n[4] a_5278_6186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5740 a_21950_16186# row_n[14] a_22442_16548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5741 VDD rowon_n[10] a_15926_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5742 VSS row_n[7] a_17326_9198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5743 a_16018_14178# a_2346_14220# a_15926_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5744 VDD rowon_n[10] a_5886_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5745 a_29470_6508# col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5746 a_11398_2492# col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5747 VDD VDD a_14922_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5748 a_5978_14178# a_2346_14220# a_5886_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5749 VDD VDD a_4882_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5750 a_15318_15222# col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5751 vcm a_1962_15222# a_20034_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5752 a_7986_9158# a_2346_9200# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5753 VSS row_n[0] a_16322_2170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5754 a_30074_3134# a_2346_3176# a_29982_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5755 vcm a_1962_3174# a_20034_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5756 a_14010_17190# a_2346_17232# a_13918_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5757 a_5278_15222# col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5758 a_25966_8154# a_1962_8194# a_26058_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5759 a_27462_1488# col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5760 a_26970_4138# a_1962_4178# a_27062_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5761 a_3970_17190# a_2346_17232# a_3878_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5762 vcm a_1962_9198# a_9994_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5763 VDD rowon_n[7] a_18938_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5764 a_30986_9158# row_n[7] a_31478_9520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5765 a_31990_5142# row_n[3] a_32482_5504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5766 a_14410_17552# col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5767 a_10906_14178# row_n[12] a_11398_14540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5768 vcm a_1962_10202# a_10998_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5769 a_17422_9520# col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5770 VSS row_n[6] a_9294_8194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5771 a_18426_5504# col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5772 a_4370_17552# col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5773 a_22346_12210# rowon_n[10] a_21950_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5774 a_14922_13174# row_n[11] a_15414_13536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5775 a_26362_11206# rowon_n[9] a_25966_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5776 a_4882_13174# row_n[11] a_5374_13536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5777 a_18026_11166# a_2346_11208# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5778 vcm a_1962_1166# a_25054_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5779 a_35094_1126# a_2346_1168# a_35002_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5780 a_7986_11166# a_2346_11208# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5781 vcm a_1962_4178# a_2966_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5782 a_34090_5142# a_2346_5184# a_33998_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5783 VDD rowon_n[8] a_21950_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5784 a_8898_9158# a_1962_9198# a_8990_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5785 a_17022_2130# a_2346_2172# a_16930_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5786 VSS row_n[15] a_20338_17230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5787 a_26970_16186# a_1962_16226# a_27062_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5788 a_31078_14178# a_2346_14220# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5789 a_12306_6186# rowon_n[4] a_11910_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5790 a_29982_6146# a_1962_6186# a_30074_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5791 VDD rowon_n[5] a_22954_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5792 a_33998_2130# row_n[0] a_34490_2492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5793 VSS row_n[14] a_24354_16226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5794 a_21342_13214# col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5795 a_34394_12210# col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5796 VDD sample a_2346_17232# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5797 a_14314_15222# rowon_n[13] a_13918_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5798 VSS row_n[10] a_11302_12210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5799 VDD rowon_n[0] a_20946_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5800 a_21038_5142# a_2346_5184# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5801 a_19030_16186# a_2346_16228# a_18938_16186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5802 a_4274_15222# rowon_n[13] a_3878_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5803 a_29982_13174# a_1962_13214# a_30074_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5804 VDD VDD a_22954_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5805 a_20434_15544# col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5806 a_8290_14218# rowon_n[12] a_7894_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5807 a_33486_14540# col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5808 vcm a_1962_12210# a_29070_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5809 VSS row_n[9] a_5278_11206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5810 VSS row_n[9] a_15318_11206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5811 a_20034_11166# a_2346_11208# a_19942_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5812 a_33086_10162# a_2346_10204# a_32994_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5813 a_20338_8194# col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5814 a_26362_2170# rowon_n[0] a_25966_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5815 a_21342_4178# col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5816 a_20946_11166# row_n[9] a_21438_11528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5817 a_10998_10162# a_2346_10204# a_10906_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5818 a_5978_9158# a_2346_9200# a_5886_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5819 VSS row_n[6] a_30378_8194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5820 a_4274_5182# rowon_n[3] a_3878_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5821 a_5278_1166# VSS a_4882_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5822 VSS row_n[2] a_31382_4178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5823 VDD rowon_n[12] a_9902_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5824 a_33998_10162# row_n[8] a_34490_10524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5825 a_35002_4138# a_1962_4178# a_35094_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5826 a_17326_4178# rowon_n[2] a_16930_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5827 a_16322_8194# rowon_n[6] a_15926_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5828 vcm a_1962_8194# a_24050_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5829 vcm a_1962_2170# a_18026_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5830 VDD rowon_n[3] a_27974_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5831 VDD rowon_n[11] a_3878_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5832 VDD rowon_n[11] a_13918_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5833 a_11398_10524# col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5834 VDD rowon_n[6] a_5886_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5835 a_25054_7150# a_2346_7192# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5836 a_26058_3134# a_2346_3176# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5837 a_13310_16226# col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5838 VDD rowon_n[1] a_3878_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5839 a_31478_4500# col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5840 a_20946_4138# row_n[2] a_21438_4500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5841 a_12002_18194# a_2346_18236# a_11910_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5842 a_34090_18194# a_2346_18236# a_33998_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5843 a_3270_16226# col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5844 vcm a_1962_15222# a_31078_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5845 a_25358_6186# col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5846 a_35002_18194# VDD a_35494_18556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5847 vcm a_1962_14218# a_35094_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5848 a_3270_9198# col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5849 a_11910_6146# row_n[4] a_12402_6508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5850 VSS row_n[4] a_35398_6186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5851 a_2346_5184# sample VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5852 a_9294_3174# rowon_n[1] a_8898_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5853 VDD rowon_n[2] a_16930_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5854 a_8290_7190# rowon_n[5] a_7894_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5855 a_12402_18556# col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5856 a_19334_18234# VDD a_18938_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5857 a_20338_13214# rowon_n[11] a_19942_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5858 vcm a_1962_6186# a_29070_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5859 a_1962_12210# sample_n VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5860 vcm a_1962_9198# a_6982_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5861 a_25054_15182# a_2346_15224# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5862 a_2346_13216# sample VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5863 a_21950_12170# a_1962_12210# a_22042_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5864 a_14314_5182# col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5865 VDD VSS a_8898_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5866 a_29070_14178# a_2346_14220# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5867 a_2874_9158# row_n[7] a_3366_9520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5868 a_3878_5142# row_n[3] a_4370_5504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5869 a_19942_1126# a_1962_1166# a_20034_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5870 VDD rowon_n[14] a_18938_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5871 VDD rowon_n[9] a_19942_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5872 a_15926_8154# row_n[6] a_16418_8516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5873 a_30074_1126# a_2346_1168# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5874 a_9994_13174# a_2346_13216# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5875 VSS row_n[15] a_31382_17230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5876 a_13918_3134# row_n[1] a_14410_3496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5877 a_13310_10202# rowon_n[8] a_12914_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5878 a_12002_2130# a_2346_2172# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5879 VSS row_n[14] a_35398_16226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5880 a_32386_13214# col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5881 a_3270_10202# rowon_n[8] a_2874_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5882 a_18330_7190# col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5883 a_19334_3174# col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5884 vcm a_1962_4178# a_33086_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5885 a_26058_17190# a_2346_17232# a_25966_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5886 a_12306_16226# rowon_n[14] a_11910_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5887 VSS row_n[1] a_20338_3174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5888 a_7894_7150# row_n[5] a_8386_7512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5889 a_30378_3174# rowon_n[1] a_29982_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5890 VDD VDD a_33998_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5891 a_26970_17190# row_n[15] a_27462_17552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5892 a_31478_15544# col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5893 vcm a_1962_13214# a_27062_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5894 a_31078_11166# a_2346_11208# a_30986_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5895 a_34090_3134# a_2346_3176# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5896 a_3878_15182# a_1962_15222# a_3970_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5897 a_13918_15182# a_1962_15222# a_14010_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5898 VSS row_n[7] a_10298_9198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5899 a_23046_7150# a_2346_7192# a_22954_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5900 a_22442_6508# col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5901 a_5886_2130# row_n[0] a_6378_2492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5902 a_17934_14178# a_1962_14218# a_18026_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5903 a_31990_11166# row_n[9] a_32482_11528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5904 VDD rowon_n[4] a_31990_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5905 a_18938_1126# en_bit_n[2] a_19430_1488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5906 a_7894_14178# a_1962_14218# a_7986_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5907 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.64e+07u l=1.6e+07u
X5908 a_20434_1488# en_bit_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5909 a_29982_14178# row_n[12] a_30474_14540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5910 vcm a_1962_10202# a_30074_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5911 VDD VSS a_29982_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5912 a_12914_2130# a_1962_2170# a_13006_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5913 VSS VDD a_25358_1166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5914 VSS row_n[3] a_24354_5182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5915 a_10394_9520# col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5916 a_11398_5504# col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5917 a_35398_1166# VSS a_35002_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5918 VSS row_n[2] a_3270_4178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5919 a_34394_5182# rowon_n[3] a_33998_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5920 a_18330_13214# rowon_n[11] a_17934_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5921 a_28978_10162# a_1962_10202# a_29070_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5922 a_28066_5142# a_2346_5184# a_27974_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5923 vcm a_1962_16226# a_8990_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5924 vcm a_1962_16226# a_19030_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5925 a_23958_6146# a_1962_6186# a_24050_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5926 a_24450_3496# col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5927 VDD sample_n a_1962_9198# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5928 VDD rowon_n[1] a_33998_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5929 a_23046_16186# a_2346_16228# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5930 VDD rowon_n[9] a_17934_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5931 VSS row_n[1] a_29374_3174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5932 a_3366_4500# col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5933 a_33390_9198# col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5934 a_15414_7512# col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5935 VSS row_n[15] a_29374_17230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5936 a_33390_15222# rowon_n[13] a_32994_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5937 VSS row_n[10] a_30378_12210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5938 a_16018_7150# a_2346_7192# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5939 VSS row_n[4] a_7286_6186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5940 a_7986_14178# a_2346_14220# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5941 a_18026_14178# a_2346_14220# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5942 VSS row_n[9] a_34394_11206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5943 a_32386_2170# col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5944 a_13406_2492# col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5945 a_3970_4138# a_2346_4180# a_3878_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5946 a_9994_9158# a_2346_9200# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5947 a_25054_12170# a_2346_12212# a_24962_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5948 a_11302_11206# rowon_n[9] a_10906_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5949 a_27974_8154# a_1962_8194# a_28066_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5950 a_29470_1488# col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5951 VSS row_n[0] a_18330_2170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5952 a_32082_3134# a_2346_3176# a_31990_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5953 a_28978_4138# a_1962_4178# a_29070_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5954 a_29470_15544# col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5955 VDD rowon_n[11] a_32994_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5956 a_25966_12170# row_n[10] a_26458_12532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5957 a_29070_11166# a_2346_11208# a_28978_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5958 a_30474_10524# col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5959 a_32994_9158# row_n[7] a_33486_9520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5960 a_33998_5142# row_n[3] a_34490_5504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5961 a_9994_10162# a_2346_10204# a_9902_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5962 a_10298_4178# rowon_n[2] a_9902_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5963 a_11910_16186# a_1962_16226# a_12002_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5964 VDD rowon_n[12] a_8898_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5965 vcm a_1962_2170# a_10998_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5966 VDD rowon_n[3] a_20946_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5967 VDD sample_n a_1962_16226# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5968 a_16930_7150# a_1962_7190# a_17022_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5969 vcm a_1962_17230# a_23046_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5970 a_8290_17230# col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5971 a_18330_17230# col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5972 vcm a_1962_4178# a_4974_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5973 VDD rowon_n[2] a_9902_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5974 vcm a_1962_12210# a_14010_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5975 vcm a_1962_12210# a_3970_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5976 a_14314_6186# rowon_n[4] a_13918_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5977 vcm a_1962_6186# a_22042_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5978 a_2346_18236# sample VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5979 a_17934_15182# row_n[13] a_18426_15544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5980 a_29374_13214# rowon_n[11] a_28978_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5981 vcm a_1962_11206# a_18026_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5982 VSS row_n[8] a_26362_10202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5983 a_7894_15182# row_n[13] a_8386_15544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5984 vcm a_1962_11206# a_7986_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5985 a_26970_11166# a_1962_11206# a_27062_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5986 VDD rowon_n[4] a_3878_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5987 VDD rowon_n[0] a_22954_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5988 VDD sample a_2346_3176# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5989 a_23046_5142# a_2346_5184# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5990 VDD rowon_n[10] a_24962_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5991 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.64e+07u l=1.6e+07u
X5992 a_28370_2170# rowon_n[0] a_27974_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5993 VSS row_n[2] a_33390_4178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5994 a_23350_4178# col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5995 VDD rowon_n[9] a_28978_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5996 a_7986_9158# a_2346_9200# a_7894_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5997 VSS row_n[6] a_32386_8194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5998 a_6282_5182# rowon_n[3] a_5886_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5999 a_7286_1166# VSS a_6890_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6000 vcm a_1962_8194# a_26058_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6001 vcm a_1962_4178# a_27062_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6002 VSS VDD a_27366_18234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6003 a_31382_16226# rowon_n[14] a_30986_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6004 a_24354_15222# col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6005 VDD rowon_n[6] a_7894_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6006 a_17326_17230# rowon_n[15] a_16930_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6007 a_28370_14218# col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6008 a_11302_7190# col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6009 a_28066_3134# a_2346_3176# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6010 a_12306_3174# col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6011 a_7286_17230# rowon_n[15] a_6890_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6012 a_19942_16186# a_1962_16226# a_20034_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6013 a_32994_15182# a_1962_15222# a_33086_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6014 a_31990_9158# a_1962_9198# a_32082_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6015 a_27062_7150# a_2346_7192# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6016 a_22954_4138# row_n[2] a_23446_4500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6017 a_3970_18194# a_2346_18236# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6018 a_14010_18194# a_2346_18236# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6019 a_23446_17552# col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6020 VSS row_n[11] a_8290_13214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6021 VSS row_n[11] a_18330_13214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6022 a_23046_13174# a_2346_13216# a_22954_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6023 VDD rowon_n[1] a_5886_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6024 a_33486_4500# col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6025 a_13918_6146# row_n[4] a_14410_6508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6026 a_27462_16548# col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6027 a_23958_13174# row_n[11] a_24450_13536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6028 a_18026_11166# a_2346_11208# a_17934_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6029 a_5278_9198# col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6030 a_7986_11166# a_2346_11208# a_7894_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6031 VDD rowon_n[13] a_6890_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6032 VDD rowon_n[13] a_16930_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6033 vcm a_1962_9198# a_8990_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6034 a_11910_1126# VDD a_12402_1488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6035 a_18426_11528# col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6036 a_4274_2170# col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6037 a_8386_11528# col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6038 vcm a_1962_6186# a_30074_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6039 a_16322_5182# col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6040 a_17326_1166# col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6041 a_16322_18234# col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6042 vcm a_1962_18234# a_21038_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6043 a_6282_18234# col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6044 vcm a_1962_17230# a_34090_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6045 a_5886_5142# row_n[3] a_6378_5504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6046 a_4882_9158# row_n[7] a_5374_9520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6047 a_17934_8154# row_n[6] a_18426_8516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6048 a_25054_10162# a_2346_10204# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6049 a_32082_1126# a_2346_1168# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6050 a_21038_5142# a_2346_5184# a_20946_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6051 a_11910_17190# row_n[15] a_12402_17552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6052 vcm a_1962_13214# a_12002_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6053 a_14010_2130# a_2346_2172# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6054 a_15926_3134# row_n[1] a_16418_3496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6055 a_5886_16186# row_n[14] a_6378_16548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6056 a_15926_16186# row_n[14] a_16418_16548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6057 a_27366_14218# rowon_n[12] a_26970_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6058 a_27366_9198# col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6059 vcm a_1962_4178# a_35094_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6060 a_28066_17190# a_2346_17232# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6061 a_28978_13174# a_1962_13214# a_29070_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6062 VSS row_n[1] a_22346_3174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6063 a_31382_7190# rowon_n[5] a_30986_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6064 a_32386_3174# rowon_n[1] a_31990_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6065 a_23350_10202# col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6066 VSS row_n[7] a_12306_9198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6067 a_26058_3134# a_2346_3176# a_25966_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6068 a_25054_7150# a_2346_7192# a_24962_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6069 a_24450_6508# col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6070 a_7894_2130# row_n[0] a_8386_2492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6071 a_22346_16226# col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6072 a_16322_12210# rowon_n[10] a_15926_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6073 a_26970_9158# row_n[7] a_27462_9520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6074 VDD rowon_n[4] a_33998_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6075 a_6282_12210# rowon_n[10] a_5886_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6076 a_13918_10162# a_1962_10202# a_14010_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6077 a_2966_9158# a_2346_9200# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6078 VSS row_n[0] a_11302_2170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6079 a_22442_12532# col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6080 a_3878_10162# a_1962_10202# a_3970_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6081 a_20946_8154# a_1962_8194# a_21038_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6082 a_22442_1488# col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6083 VDD VSS a_31990_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6084 a_21950_4138# a_1962_4178# a_22042_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6085 a_5278_18234# VDD a_4882_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6086 a_15318_18234# VDD a_14922_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6087 a_31078_8154# a_2346_8196# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6088 a_14922_2130# a_1962_2170# a_15014_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6089 a_21438_18556# col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6090 a_30986_16186# a_1962_16226# a_31078_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6091 VSS row_n[12] a_16322_14218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6092 a_21038_14178# a_2346_14220# a_20946_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6093 VSS VDD a_27366_1166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6094 VSS row_n[12] a_6282_14218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6095 a_12402_9520# col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6096 VSS row_n[6] a_4274_8194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6097 a_13406_5504# col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6098 VSS row_n[2] a_5278_4178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6099 a_16930_17190# a_1962_17230# a_17022_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6100 VDD rowon_n[8] a_15926_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6101 a_6890_17190# a_1962_17230# a_6982_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6102 VDD rowon_n[8] a_5886_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6103 VSS row_n[15] a_4274_17230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6104 VSS row_n[15] a_14314_17230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6105 VDD rowon_n[14] a_14922_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6106 VDD rowon_n[14] a_4882_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6107 a_15318_13214# col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6108 vcm a_1962_13214# a_20034_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6109 vcm a_1962_1166# a_20034_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6110 a_30074_1126# a_2346_1168# a_29982_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6111 a_19942_17190# row_n[15] a_20434_17552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6112 a_14010_15182# a_2346_15224# a_13918_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6113 a_5278_13214# col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6114 vcm a_1962_12210# a_33086_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6115 a_25966_6146# a_1962_6186# a_26058_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
C0 m2_1732_946# vcm 0.42fF
C1 a_1962_10202# a_23046_10162# 0.27fF
C2 a_2346_9200# rowoff_n[7] 4.09fF
C3 a_12306_5182# vcm 0.22fF
C4 a_1962_8194# row_n[6] 25.57fF
C5 a_32082_15182# vcm 0.62fF
C6 a_6890_15182# rowoff_n[13] 0.24fF
C7 m2_1732_18014# m3_1864_17142# 0.15fF
C8 m2_12776_18014# m3_13912_18146# 0.13fF
C9 a_12914_7150# rowoff_n[5] 0.24fF
C10 a_2346_7192# a_18026_7150# 0.19fF
C11 a_1962_7190# a_16322_7190# 0.14fF
C12 a_14010_15182# m2_14208_15430# 0.16fF
C13 a_27062_8154# a_27062_7150# 1.00fF
C14 a_25358_9198# vcm 0.22fF
C15 a_28066_17190# a_29070_17190# 0.97fF
C16 a_16018_3134# m2_16216_3382# 0.16fF
C17 a_22954_5142# rowoff_n[3] 0.24fF
C18 a_6982_3134# ctop 3.57fF
C19 a_1962_9198# col_n[15] 0.13fF
C20 a_34090_9158# row_n[7] 0.17fF
C21 a_35002_11166# m2_34864_10986# 0.16fF
C22 a_15014_14178# col[12] 0.29fF
C23 a_14922_11166# VDD 0.23fF
C24 a_1962_9198# a_29374_9198# 0.14fF
C25 a_16930_9158# a_17022_9158# 0.26fF
C26 a_2346_9200# a_31078_9158# 0.19fF
C27 a_1962_3174# col[6] 0.11fF
C28 a_32994_3134# rowoff_n[1] 0.24fF
C29 ctop col[13] 1.98fF
C30 col[3] col[4] 0.20fF
C31 a_1962_16226# col[8] 0.11fF
C32 a_2346_1168# a_7894_1126# 0.35fF
C33 a_33086_10162# col[30] 0.29fF
C34 a_20034_7150# ctop 3.58fF
C35 a_2346_2172# col[26] 0.15fF
C36 a_6982_17190# rowon_n[15] 0.14fF
C37 a_2346_15224# col[28] 0.15fF
C38 a_27974_15182# VDD 0.23fF
C39 a_22042_7150# rowon_n[5] 0.14fF
C40 a_10998_3134# a_12002_3134# 0.97fF
C41 a_2346_3176# a_20946_3134# 0.35fF
C42 a_2346_1168# m2_25828_946# 0.19fF
C43 a_33086_11166# ctop 3.57fF
C44 a_1962_18234# col[18] 0.11fF
C45 a_10998_16186# m2_11196_16434# 0.16fF
C46 a_15014_16186# col_n[12] 0.28fF
C47 a_29982_13174# a_30074_13174# 0.26fF
C48 a_13006_13174# a_13006_12170# 1.00fF
C49 a_14010_10162# vcm 0.62fF
C50 a_21038_11166# rowoff_n[9] 0.10fF
C51 a_16018_3134# col[13] 0.29fF
C52 a_1962_17230# a_7986_17190# 0.27fF
C53 m2_15788_18014# m2_16216_18442# 0.16fF
C54 a_13006_4138# m2_13204_4386# 0.16fF
C55 a_1962_5182# col_n[6] 0.13fF
C56 m2_1732_2954# m3_1864_4090# 0.15fF
C57 a_17022_3134# VDD 0.52fF
C58 m3_10900_18146# ctop 0.23fF
C59 a_2346_5184# a_33998_5142# 0.35fF
C60 a_35494_13536# VDD 0.11fF
C61 a_33086_12170# col_n[30] 0.28fF
C62 a_31078_9158# rowoff_n[7] 0.10fF
C63 a_7286_4178# vcm 0.22fF
C64 a_2346_14220# a_2874_14178# 0.35fF
C65 a_27062_14178# vcm 0.62fF
C66 a_1962_2170# a_28066_2130# 0.27fF
C67 a_30074_7150# VDD 0.52fF
C68 a_24050_7150# a_25054_7150# 0.97fF
C69 a_2966_14178# m2_1732_13998# 0.96fF
C70 a_2346_11208# col[19] 0.15fF
C71 a_19030_10162# row_n[8] 0.17fF
C72 a_20338_8194# vcm 0.22fF
C73 col[18] rowoff_n[13] 0.11fF
C74 a_1962_16226# a_14314_16226# 0.14fF
C75 a_26058_17190# a_26058_16186# 1.00fF
C76 a_2346_16228# a_16018_16186# 0.19fF
C77 VDD rowoff_n[4] 1.17fF
C78 vcm rowoff_n[8] 0.20fF
C79 sample_n rowoff_n[5] 0.38fF
C80 a_16018_5142# col_n[13] 0.28fF
C81 m2_22816_946# vcm 0.42fF
C82 a_9902_10162# VDD 0.23fF
C83 a_7986_17190# m2_8184_17438# 0.16fF
C84 a_1962_7190# col[26] 0.11fF
C85 a_8898_12170# rowoff_n[10] 0.24fF
C86 a_33390_12210# vcm 0.22fF
C87 a_9994_5142# m2_10192_5390# 0.16fF
C88 a_6982_8154# rowon_n[6] 0.14fF
C89 a_1962_14218# col_n[0] 0.13fF
C90 a_15014_6146# ctop 3.58fF
C91 m3_34996_10114# VDD 0.26fF
C92 a_22954_14178# VDD 0.23fF
C93 a_31078_15182# col[28] 0.29fF
C94 a_2346_10204# a_5886_10162# 0.35fF
C95 a_5886_2130# rowoff_n[0] 0.24fF
C96 col[2] rowoff_n[14] 0.11fF
C97 a_22954_16186# rowoff_n[14] 0.24fF
C98 m2_17796_18014# ctop 0.18fF
C99 a_8990_3134# a_8990_2130# 1.00fF
C100 a_25966_3134# a_26058_3134# 0.26fF
C101 a_28066_10162# ctop 3.58fF
C102 a_2346_7192# col[10] 0.15fF
C103 a_2346_12212# a_18938_12170# 0.35fF
C104 a_9994_12170# a_10998_12170# 0.97fF
C105 a_26058_11166# rowon_n[9] 0.14fF
C106 a_1962_9198# col_n[26] 0.13fF
C107 a_8990_9158# vcm 0.62fF
C108 a_12002_2130# VDD 0.55fF
C109 a_14010_8154# col[11] 0.29fF
C110 a_1962_3174# col[17] 0.11fF
C111 VDD col_n[2] 4.94fF
C112 sample vcm 13.47fF
C113 a_1962_9198# a_13006_9158# 0.27fF
C114 a_1962_16226# col[19] 0.11fF
C115 ctop col[24] 1.98fF
C116 a_3970_11166# row_n[9] 0.17fF
C117 a_2346_14220# a_31990_14178# 0.35fF
C118 a_31078_17190# col_n[28] 0.28fF
C119 a_22042_13174# vcm 0.62fF
C120 a_32082_4138# col[29] 0.29fF
C121 a_6982_6146# m2_7180_6394# 0.16fF
C122 a_25054_6146# VDD 0.52fF
C123 a_1962_6186# a_6282_6186# 0.14fF
C124 a_22042_7150# a_22042_6146# 1.00fF
C125 a_2346_6188# a_7986_6146# 0.19fF
C126 a_3970_8154# rowoff_n[6] 0.10fF
C127 a_1962_11206# a_26058_11166# 0.27fF
C128 a_15318_7190# vcm 0.22fF
C129 a_23046_16186# a_24050_16186# 0.97fF
C130 a_35094_17190# vcm 0.12fF
C131 a_9994_17190# rowoff_n[15] 0.10fF
C132 a_1962_18234# col[29] 0.11fF
C133 a_14010_6146# rowoff_n[4] 0.10fF
C134 a_2346_3176# a_1962_3174# 2.62fF
C135 a_2346_3176# col[1] 0.15fF
C136 a_4882_9158# VDD 0.23fF
C137 a_2346_16228# col[3] 0.15fF
C138 a_1962_8194# a_19334_8194# 0.14fF
C139 a_2346_8196# a_21038_8154# 0.19fF
C140 a_11910_8154# a_12002_8154# 0.26fF
C141 a_23046_14178# row_n[12] 0.17fF
C142 a_14010_10162# col_n[11] 0.28fF
C143 m2_1732_1950# m2_1732_946# 0.99fF
C144 a_1962_5182# col_n[17] 0.13fF
C145 a_24050_4138# rowoff_n[2] 0.10fF
C146 a_28370_11206# vcm 0.22fF
C147 a_2966_11166# rowoff_n[9] 0.10fF
C148 a_9994_5142# ctop 3.58fF
C149 m2_16792_946# vcm 0.42fF
C150 a_17934_13174# VDD 0.23fF
C151 a_32082_6146# col_n[29] 0.28fF
C152 a_1962_12210# col[10] 0.11fF
C153 a_1962_10202# a_32386_10202# 0.14fF
C154 a_2346_10204# a_34090_10162# 0.19fF
C155 a_34090_2130# rowoff_n[0] 0.10fF
C156 m2_33860_946# vcm 0.23fF
C157 a_10998_12170# rowon_n[10] 0.14fF
C158 a_3970_7150# m2_4168_7398# 0.16fF
C159 a_5978_2130# a_6982_2130# 0.97fF
C160 a_2346_2172# a_10906_2130# 0.35fF
C161 a_2346_11208# col[30] 0.15fF
C162 m2_27836_18014# m3_26964_18146# 0.13fF
C163 a_23046_9158# ctop 3.58fF
C164 a_30986_17190# VDD 0.24fF
C165 a_26058_2130# rowon_n[0] 0.14fF
C166 col[29] rowoff_n[13] 0.11fF
C167 a_24962_12170# a_25054_12170# 0.26fF
C168 a_7986_12170# a_7986_11166# 1.00fF
C169 a_3970_8154# vcm 0.62fF
C170 a_1962_10202# m2_34864_9982# 0.17fF
C171 a_2346_4180# a_23958_4138# 0.35fF
C172 a_2346_12212# ctop 1.59fF
C173 a_3970_2130# row_n[0] 0.17fF
C174 a_12002_13174# col[9] 0.29fF
C175 a_1962_1166# col_n[8] 0.13fF
C176 a_22954_10162# rowoff_n[8] 0.24fF
C177 a_30074_15182# rowon_n[13] 0.14fF
C178 a_1962_14218# col_n[10] 0.13fF
C179 a_17022_12170# vcm 0.62fF
C180 a_24962_13174# rowoff_n[11] 0.24fF
C181 a_1962_1166# a_18026_1126# 0.26fF
C182 a_20034_5142# VDD 0.52fF
C183 m2_24824_946# VDD 0.62fF
C184 a_19030_6146# a_20034_6146# 0.97fF
C185 a_1962_6186# a_1962_5182# 0.16fF
C186 a_1962_8194# col[1] 0.11fF
C187 col[13] rowoff_n[14] 0.11fF
C188 a_30074_9158# col[27] 0.29fF
C189 a_32994_8154# rowoff_n[6] 0.24fF
C190 VDD rowoff_n[10] 1.17fF
C191 a_7986_15182# row_n[13] 0.17fF
C192 a_10298_6186# vcm 0.22fF
C193 a_2346_15224# a_5978_15182# 0.19fF
C194 a_1962_15222# a_4274_15222# 0.14fF
C195 a_21038_16186# a_21038_15182# 1.00fF
C196 a_30074_16186# vcm 0.62fF
C197 a_2346_7192# col[21] 0.15fF
C198 a_23046_5142# row_n[3] 0.17fF
C199 a_1962_3174# a_31078_3134# 0.27fF
C200 a_33086_9158# VDD 0.52fF
C201 a_23350_10202# vcm 0.22fF
C202 a_1962_17230# a_17326_17230# 0.14fF
C203 a_2346_17232# a_19030_17190# 0.19fF
C204 a_10906_17190# a_10998_17190# 0.26fF
C205 a_12002_15182# col_n[9] 0.28fF
C206 m2_1732_1950# m3_1864_1078# 0.15fF
C207 m2_2736_1950# m3_2868_2082# 2.75fF
C208 a_4974_4138# ctop 3.58fF
C209 a_1962_3174# col[28] 0.11fF
C210 col_n[4] col_n[5] 0.10fF
C211 vcm col_n[9] 2.80fF
C212 m3_1864_8106# ctop 0.23fF
C213 VDD col_n[13] 4.94fF
C214 a_13006_2130# col[10] 0.29fF
C215 a_1962_16226# col[30] 0.11fF
C216 col[14] col[15] 0.20fF
C217 a_12914_12170# VDD 0.23fF
C218 a_32082_10162# a_33086_10162# 0.97fF
C219 a_30074_11166# col_n[27] 0.28fF
C220 a_1962_10202# col_n[1] 0.13fF
C221 a_10998_3134# rowon_n[1] 0.14fF
C222 a_12002_14178# rowoff_n[12] 0.10fF
C223 a_20946_2130# a_21038_2130# 0.26fF
C224 a_3970_2130# a_3970_1126# 1.00fF
C225 a_18026_8154# ctop 3.58fF
C226 a_1962_17230# ctop 1.30fF
C227 a_25966_16186# VDD 0.23fF
C228 m2_34864_10986# vcm 0.51fF
C229 a_2346_11208# a_8898_11166# 0.35fF
C230 a_4974_11166# a_5978_11166# 0.97fF
C231 a_2346_3176# col[12] 0.15fF
C232 a_15014_16186# rowon_n[14] 0.14fF
C233 a_2346_16228# col[14] 0.15fF
C234 a_32082_10162# m2_32280_10410# 0.16fF
C235 a_31078_12170# ctop 3.58fF
C236 a_2346_8196# a_2966_8154# 0.21fF
C237 a_30074_6146# rowon_n[4] 0.14fF
C238 a_1962_5182# col_n[28] 0.13fF
C239 a_13006_4138# col_n[10] 0.28fF
C240 a_2346_13216# a_21950_13174# 0.35fF
C241 a_12002_11166# vcm 0.62fF
C242 a_1962_12210# col[21] 0.11fF
C243 a_15014_4138# VDD 0.52fF
C244 a_2966_12170# m2_3164_12418# 0.16fF
C245 m3_26964_1078# VDD 0.14fF
C246 a_33998_6146# a_34090_6146# 0.26fF
C247 a_17022_6146# a_17022_5142# 1.00fF
C248 a_7986_6146# row_n[4] 0.17fF
C249 a_1962_10202# a_16018_10162# 0.27fF
C250 a_5278_5182# vcm 0.22fF
C251 a_28066_14178# col[25] 0.29fF
C252 a_2346_15224# a_35002_15182# 0.35fF
C253 a_18026_15182# a_19030_15182# 0.97fF
C254 a_25054_15182# vcm 0.62fF
C255 m2_3740_18014# m3_3872_18146# 2.78fF
C256 a_28066_8154# VDD 0.52fF
C257 a_5886_7150# rowoff_n[5] 0.24fF
C258 a_1962_7190# a_9294_7190# 0.14fF
C259 a_6890_7150# a_6982_7150# 0.26fF
C260 a_2346_7192# a_10998_7150# 0.19fF
C261 a_1962_12210# a_29070_12170# 0.27fF
C262 m2_1732_1950# sample 0.19fF
C263 a_18330_9198# vcm 0.22fF
C264 m2_1732_12994# sample_n 0.15fF
C265 a_2966_3134# m2_2736_1950# 0.99fF
C266 a_2346_12212# col[5] 0.15fF
C267 a_15926_5142# rowoff_n[3] 0.24fF
C268 a_27062_9158# row_n[7] 0.17fF
C269 a_29070_11166# m2_29268_11414# 0.16fF
C270 a_7894_11166# VDD 0.23fF
C271 a_1962_1166# col_n[19] 0.13fF
C272 a_30074_10162# a_30074_9158# 1.00fF
C273 a_2346_9200# a_24050_9158# 0.19fF
C274 a_1962_9198# a_22346_9198# 0.14fF
C275 a_10998_7150# col[8] 0.29fF
C276 a_1962_14218# col_n[21] 0.13fF
C277 a_25966_3134# rowoff_n[1] 0.24fF
C278 m2_34864_5966# m2_35292_6394# 0.16fF
C279 a_31382_13214# vcm 0.22fF
C280 col[24] rowoff_n[14] 0.11fF
C281 m2_15788_18014# col_n[13] 0.25fF
C282 a_1962_8194# col[12] 0.11fF
C283 a_28066_16186# col_n[25] 0.28fF
C284 a_13006_7150# ctop 3.58fF
C285 a_2346_13216# row_n[11] 0.35fF
C286 a_34090_14178# m2_34864_13998# 0.96fF
C287 a_29070_3134# col[26] 0.29fF
C288 a_20946_15182# VDD 0.23fF
C289 a_19942_11166# a_20034_11166# 0.26fF
C290 a_3878_18194# m2_3740_18014# 0.16fF
C291 a_15014_7150# rowon_n[5] 0.14fF
C292 a_2346_3176# a_13918_3134# 0.35fF
C293 a_26058_11166# ctop 3.58fF
C294 a_28066_2130# m2_27836_946# 0.99fF
C295 a_1962_9198# rowon_n[7] 1.18fF
C296 a_14010_11166# rowoff_n[9] 0.10fF
C297 a_6982_10162# vcm 0.62fF
C298 a_10998_9158# col_n[8] 0.28fF
C299 vcm col_n[20] 2.80fF
C300 VDD col_n[24] 4.99fF
C301 col[8] rowoff_n[15] 0.11fF
C302 m2_8760_18014# m2_9188_18442# 0.16fF
C303 m2_5748_946# col_n[3] 0.37fF
C304 a_9994_3134# VDD 0.52fF
C305 a_14010_5142# a_15014_5142# 0.97fF
C306 a_26058_12170# m2_26256_12418# 0.16fF
C307 a_2346_5184# a_26970_5142# 0.35fF
C308 a_1962_10202# col_n[12] 0.13fF
C309 a_34090_10162# rowon_n[8] 0.14fF
C310 a_24050_9158# rowoff_n[7] 0.10fF
C311 a_29070_5142# col_n[26] 0.28fF
C312 a_16018_15182# a_16018_14178# 1.00fF
C313 a_32994_15182# a_33086_15182# 0.26fF
C314 a_2966_7150# col_n[0] 0.28fF
C315 a_20034_14178# vcm 0.62fF
C316 a_28066_15182# rowoff_n[13] 0.10fF
C317 a_1962_4178# col[3] 0.11fF
C318 a_1962_2170# a_21038_2130# 0.27fF
C319 a_1962_17230# col[5] 0.11fF
C320 a_23046_7150# VDD 0.52fF
C321 a_34090_7150# rowoff_n[5] 0.10fF
C322 a_12002_10162# row_n[8] 0.17fF
C323 a_2346_3176# col[23] 0.15fF
C324 a_13310_8194# vcm 0.22fF
C325 a_5886_16186# a_5978_16186# 0.26fF
C326 a_1962_16226# a_7286_16226# 0.14fF
C327 a_2346_16228# col[25] 0.15fF
C328 a_2346_16228# a_8990_16186# 0.19fF
C329 a_33086_18194# vcm 0.12fF
C330 a_1962_4178# a_34090_4138# 0.27fF
C331 a_2346_10204# VDD 32.63fF
C332 a_1962_17230# m2_1732_17010# 0.15fF
C333 a_27062_9158# a_28066_9158# 0.97fF
C334 a_2874_13174# a_2966_13174# 0.26fF
C335 a_2346_13216# a_3878_13174# 0.35fF
C336 a_2346_4180# row_n[2] 0.35fF
C337 a_8990_12170# col[6] 0.29fF
C338 a_26362_12210# vcm 0.22fF
C339 a_1962_1166# a_27366_1166# 0.14fF
C340 a_7986_6146# ctop 3.58fF
C341 a_31078_13174# row_n[11] 0.17fF
C342 m3_22948_18146# VDD 0.38fF
C343 a_23046_13174# m2_23244_13422# 0.16fF
C344 a_1962_6186# col_n[3] 0.13fF
C345 a_15926_14178# VDD 0.23fF
C346 a_27062_8154# col[24] 0.29fF
C347 a_15926_16186# rowoff_n[14] 0.24fF
C348 m2_3740_18014# ctop 0.18fF
C349 a_29070_2130# m3_28972_1078# 0.15fF
C350 a_24962_1126# m2_24824_946# 0.16fF
C351 a_21038_10162# ctop 3.58fF
C352 a_28978_18194# VDD 0.33fF
C353 m2_32856_18014# vcm 0.28fF
C354 a_2346_12212# a_11910_12170# 0.35fF
C355 a_2346_12212# col[16] 0.15fF
C356 a_19030_11166# rowon_n[9] 0.14fF
C357 a_34394_10202# vcm 0.22fF
C358 a_4974_2130# VDD 0.55fF
C359 m3_29976_1078# ctop 0.23fF
C360 a_1962_1166# col_n[30] 0.14fF
C361 a_28978_5142# a_29070_5142# 0.26fF
C362 a_12002_5142# a_12002_4138# 1.00fF
C363 a_8990_14178# col_n[6] 0.28fF
C364 a_34090_14178# ctop 3.42fF
C365 a_1962_9198# a_5978_9158# 0.27fF
C366 a_13006_14178# a_14010_14178# 0.97fF
C367 a_2346_14220# a_24962_14178# 0.35fF
C368 a_1962_8194# col[23] 0.11fF
C369 a_2346_18236# a_33998_18194# 0.35fF
C370 a_15014_13174# vcm 0.62fF
C371 a_27062_10162# col_n[24] 0.28fF
C372 a_18026_6146# VDD 0.52fF
C373 a_20034_14178# m2_20232_14426# 0.16fF
C374 a_1962_15222# VDD 2.73fF
C375 a_1962_11206# a_19030_11166# 0.27fF
C376 a_8290_7190# vcm 0.22fF
C377 a_2966_16186# a_2966_15182# 1.00fF
C378 m2_34864_8978# row_n[7] 0.15fF
C379 a_2874_17190# rowoff_n[15] 0.24fF
C380 a_28066_17190# vcm 0.60fF
C381 m2_23820_18014# VDD 1.04fF
C382 a_6982_6146# rowoff_n[4] 0.10fF
C383 a_31078_10162# VDD 0.52fF
C384 a_1962_8194# a_12306_8194# 0.14fF
C385 a_2346_8196# a_14010_8154# 0.19fF
C386 a_25054_9158# a_25054_8154# 1.00fF
C387 a_16018_14178# row_n[12] 0.17fF
C388 vcm col_n[31] 2.78fF
C389 sample row_n[15] 1.03fF
C390 VDD row_n[14] 2.93fF
C391 a_1962_13214# a_32082_13174# 0.27fF
C392 col[25] col[26] 0.21fF
C393 col[19] rowoff_n[15] 0.11fF
C394 a_2346_8196# col[7] 0.15fF
C395 a_9994_3134# col_n[7] 0.28fF
C396 a_17022_4138# rowoff_n[2] 0.10fF
C397 a_30074_12170# rowoff_n[10] 0.10fF
C398 a_21342_11206# vcm 0.22fF
C399 a_31078_4138# row_n[2] 0.17fF
C400 a_1962_10202# col_n[23] 0.13fF
C401 a_6982_17190# col[4] 0.29fF
C402 a_10906_13174# VDD 0.23fF
C403 a_2346_18236# m2_33860_18014# 0.19fF
C404 m2_9764_946# vcm 0.42fF
C405 a_1962_10202# a_25358_10202# 0.14fF
C406 a_14922_10162# a_15014_10162# 0.26fF
C407 a_2346_10204# a_27062_10162# 0.19fF
C408 a_27062_2130# rowoff_n[0] 0.10fF
C409 a_1962_4178# col[14] 0.11fF
C410 a_1962_17230# col[16] 0.11fF
C411 a_35398_15222# vcm 0.23fF
C412 a_25054_13174# col[22] 0.29fF
C413 a_3970_12170# rowon_n[10] 0.14fF
C414 m2_17796_18014# m3_18932_18146# 0.13fF
C415 a_16018_9158# ctop 3.58fF
C416 a_17022_15182# m2_17220_15430# 0.16fF
C417 a_23958_17190# VDD 0.24fF
C418 a_19030_2130# rowon_n[0] 0.14fF
C419 m2_1732_13998# vcm 0.45fF
C420 a_19030_3134# m2_19228_3382# 0.16fF
C421 a_33998_2130# VDD 0.21fF
C422 a_2346_4180# a_16930_4138# 0.35fF
C423 a_8990_4138# a_9994_4138# 0.97fF
C424 a_29070_13174# ctop 3.58fF
C425 a_27974_14178# a_28066_14178# 0.26fF
C426 a_10998_14178# a_10998_13174# 1.00fF
C427 a_15926_10162# rowoff_n[8] 0.24fF
C428 a_2346_17232# col[0] 0.15fF
C429 a_23046_15182# rowon_n[13] 0.14fF
C430 a_7986_6146# col[5] 0.29fF
C431 a_9994_12170# vcm 0.62fF
C432 a_17934_13174# rowoff_n[11] 0.24fF
C433 a_1962_6186# col_n[14] 0.13fF
C434 a_13006_5142# VDD 0.52fF
C435 a_2346_6188# a_29982_6146# 0.35fF
C436 a_25054_15182# col_n[22] 0.28fF
C437 a_25966_8154# rowoff_n[6] 0.24fF
C438 m2_15788_946# a_1962_1166# 0.18fF
C439 a_26058_2130# col[23] 0.29fF
C440 a_3270_6186# vcm 0.22fF
C441 a_1962_13214# col[7] 0.11fF
C442 a_23046_16186# vcm 0.62fF
C443 a_31990_17190# rowoff_n[15] 0.24fF
C444 m2_30848_18014# col[28] 0.28fF
C445 a_16018_5142# row_n[3] 0.17fF
C446 a_1962_3174# a_24050_3134# 0.27fF
C447 a_1962_1166# m2_32856_946# 0.18fF
C448 a_2966_10162# ctop 3.42fF
C449 a_26058_9158# VDD 0.52fF
C450 a_14010_16186# m2_14208_16434# 0.16fF
C451 a_22042_8154# a_23046_8154# 0.97fF
C452 a_2346_12212# col[27] 0.15fF
C453 a_33086_1126# vcm 0.12fF
C454 a_16322_10202# vcm 0.22fF
C455 a_2346_17232# a_12002_17190# 0.19fF
C456 a_1962_17230# a_10298_17230# 0.14fF
C457 a_16018_4138# m2_16216_4386# 0.16fF
C458 m3_25960_18146# ctop 0.23fF
C459 a_7986_8154# col_n[5] 0.28fF
C460 a_35002_12170# m2_34864_11990# 0.16fF
C461 a_5886_12170# VDD 0.23fF
C462 a_3970_3134# rowon_n[1] 0.14fF
C463 a_29374_14218# vcm 0.22fF
C464 a_4974_14178# rowoff_n[12] 0.10fF
C465 a_26058_4138# col_n[23] 0.28fF
C466 a_1962_2170# a_30378_2170# 0.14fF
C467 a_2346_2172# a_32082_2130# 0.19fF
C468 a_1962_2170# col_n[5] 0.13fF
C469 a_34090_3134# a_34090_2130# 1.00fF
C470 a_1962_15222# col_n[7] 0.13fF
C471 a_10998_8154# ctop 3.58fF
C472 a_18938_16186# VDD 0.23fF
C473 a_28978_1126# VDD 0.44fF
C474 a_7986_16186# rowon_n[14] 0.14fF
C475 a_2874_18194# m2_2736_18014# 0.16fF
C476 a_6982_4138# a_6982_3134# 1.00fF
C477 a_23958_4138# a_24050_4138# 0.26fF
C478 a_24050_12170# ctop 3.58fF
C479 col_n[3] row_n[12] 0.23fF
C480 col_n[9] row_n[15] 0.23fF
C481 col_n[0] row_n[10] 0.23fF
C482 VDD rowon_n[8] 2.61fF
C483 col_n[7] row_n[14] 0.23fF
C484 col_n[5] row_n[13] 0.23fF
C485 col_n[1] row_n[11] 0.23fF
C486 vcm rowon_n[10] 0.50fF
C487 a_2346_8196# col[18] 0.15fF
C488 col[30] rowoff_n[15] 0.11fF
C489 a_10998_17190# m2_11196_17438# 0.16fF
C490 a_21038_17190# m2_20808_18014# 1.00fF
C491 a_23046_6146# rowon_n[4] 0.14fF
C492 a_7986_13174# a_8990_13174# 0.97fF
C493 a_2346_13216# a_14922_13174# 0.35fF
C494 a_4974_11166# vcm 0.62fF
C495 a_13006_5142# m2_13204_5390# 0.16fF
C496 a_7986_4138# VDD 0.52fF
C497 m2_2736_1950# row_n[0] 0.15fF
C498 a_5978_11166# col[3] 0.29fF
C499 m3_1864_2082# VDD 0.25fF
C500 a_1962_10202# a_8990_10162# 0.27fF
C501 a_1962_4178# col[25] 0.11fF
C502 a_1962_17230# col[27] 0.11fF
C503 a_2346_15224# a_27974_15182# 0.35fF
C504 a_18026_15182# vcm 0.62fF
C505 a_24050_7150# col[21] 0.29fF
C506 a_1962_11206# sample 0.14fF
C507 a_21038_8154# VDD 0.52fF
C508 a_2346_7192# a_3970_7150# 0.19fF
C509 a_20034_8154# a_20034_7150# 1.00fF
C510 a_2966_15182# m2_1732_15002# 0.96fF
C511 sample_n rowoff_n[12] 0.38fF
C512 a_1962_12210# a_22042_12170# 0.27fF
C513 m2_13780_946# m3_13912_1078# 2.79fF
C514 a_11302_9198# vcm 0.22fF
C515 a_21038_17190# a_22042_17190# 0.97fF
C516 a_8898_5142# rowoff_n[3] 0.24fF
C517 a_20034_9158# row_n[7] 0.17fF
C518 a_2346_4180# col[9] 0.15fF
C519 a_34090_12170# VDD 0.54fF
C520 m2_24824_946# m3_25960_1078# 0.13fF
C521 a_1962_9198# a_15318_9198# 0.14fF
C522 a_2346_17232# col[11] 0.15fF
C523 a_2346_9200# a_17022_9158# 0.19fF
C524 a_9902_9158# a_9994_9158# 0.26fF
C525 a_5978_13174# col_n[3] 0.28fF
C526 m2_1732_3958# rowoff_n[2] 0.12fF
C527 a_18938_3134# rowoff_n[1] 0.24fF
C528 a_1962_6186# col_n[25] 0.13fF
C529 a_33998_14178# rowoff_n[12] 0.24fF
C530 a_24354_13214# vcm 0.22fF
C531 a_31078_2130# a_32082_2130# 0.97fF
C532 a_9994_6146# m2_10192_6394# 0.16fF
C533 a_5978_7150# ctop 3.58fF
C534 a_24050_9158# col_n[21] 0.28fF
C535 a_13918_15182# VDD 0.23fF
C536 a_1962_13214# col[18] 0.11fF
C537 a_1962_11206# a_28370_11206# 0.14fF
C538 a_33086_12170# a_33086_11166# 1.00fF
C539 a_2346_11208# a_30074_11166# 0.19fF
C540 a_5978_17190# m3_5880_18146# 0.15fF
C541 rowon_n[5] rowoff_n[5] 20.27fF
C542 a_7986_7150# rowon_n[5] 0.14fF
C543 a_2346_3176# a_6890_3134# 0.35fF
C544 a_3970_3134# a_4974_3134# 0.97fF
C545 a_19030_11166# ctop 3.58fF
C546 a_22954_13174# a_23046_13174# 0.26fF
C547 a_5978_13174# a_5978_12170# 1.00fF
C548 a_6982_11166# rowoff_n[9] 0.10fF
C549 m2_1732_18014# m2_2160_18442# 0.16fF
C550 a_2874_3134# VDD 0.24fF
C551 a_6982_2130# col_n[4] 0.28fF
C552 a_2346_5184# a_19942_5142# 0.35fF
C553 a_32082_15182# ctop 3.58fF
C554 a_2346_13216# col[2] 0.15fF
C555 a_27062_10162# rowon_n[8] 0.14fF
C556 a_17022_9158# rowoff_n[7] 0.10fF
C557 a_3970_16186# col[1] 0.29fF
C558 m2_28840_946# col_n[26] 0.42fF
C559 a_1962_2170# col_n[16] 0.13fF
C560 a_1962_15222# col_n[18] 0.13fF
C561 a_21038_15182# rowoff_n[13] 0.10fF
C562 a_13006_14178# vcm 0.62fF
C563 a_6982_7150# m2_7180_7398# 0.16fF
C564 a_1962_2170# a_14010_2130# 0.27fF
C565 m2_32856_18014# m3_31984_18146# 0.13fF
C566 a_16018_7150# VDD 0.52fF
C567 a_27062_7150# rowoff_n[5] 0.10fF
C568 a_2346_7192# a_32994_7150# 0.35fF
C569 a_17022_7150# a_18026_7150# 0.97fF
C570 a_22042_12170# col[19] 0.29fF
C571 a_4974_10162# row_n[8] 0.17fF
C572 a_1962_9198# col[9] 0.11fF
C573 a_2346_14220# rowon_n[12] 0.26fF
C574 a_6282_8194# vcm 0.22fF
C575 a_19030_17190# a_19030_16186# 1.00fF
C576 a_26058_18194# vcm 0.12fF
C577 col_n[12] row_n[11] 0.23fF
C578 col_n[20] row_n[15] 0.23fF
C579 col_n[10] row_n[10] 0.23fF
C580 col_n[2] row_n[6] 0.23fF
C581 vcm row_n[5] 0.49fF
C582 sample row_n[4] 1.03fF
C583 col_n[26] col_n[27] 0.10fF
C584 col_n[16] row_n[13] 0.23fF
C585 VDD row_n[3] 2.93fF
C586 col_n[14] row_n[12] 0.23fF
C587 col_n[18] row_n[14] 0.23fF
C588 col_n[4] row_n[7] 0.23fF
C589 col_n[6] row_n[8] 0.23fF
C590 col_n[8] row_n[9] 0.23fF
C591 a_2346_8196# col[29] 0.15fF
C592 a_1962_4178# a_27062_4138# 0.27fF
C593 a_29070_11166# VDD 0.52fF
C594 m3_25960_1078# m3_26964_1078# 0.22fF
C595 a_2346_2172# vcm 0.40fF
C596 a_19334_12210# vcm 0.22fF
C597 a_1962_1166# a_20338_1166# 0.19fF
C598 a_24050_13174# row_n[11] 0.17fF
C599 a_4974_5142# col[2] 0.29fF
C600 a_8898_14178# VDD 0.23fF
C601 m2_34864_10986# rowon_n[9] 0.13fF
C602 a_30074_11166# a_31078_11166# 0.97fF
C603 a_22042_14178# col_n[19] 0.28fF
C604 a_1962_11206# col_n[9] 0.13fF
C605 a_32386_16226# vcm 0.22fF
C606 a_8898_16186# rowoff_n[14] 0.24fF
C607 a_3970_8154# m2_4168_8402# 0.16fF
C608 a_18938_3134# a_19030_3134# 0.26fF
C609 a_1962_3174# a_33390_3174# 0.14fF
C610 a_14010_10162# ctop 3.58fF
C611 a_2966_8154# VDD 0.56fF
C612 a_1962_5182# col[0] 0.11fF
C613 a_21950_18194# VDD 0.33fF
C614 m2_18800_18014# vcm 0.28fF
C615 a_2346_12212# a_4882_12170# 0.35fF
C616 a_12002_11166# rowon_n[9] 0.14fF
C617 a_2346_4180# col[20] 0.15fF
C618 a_31990_3134# VDD 0.23fF
C619 a_2346_17232# col[22] 0.15fF
C620 a_1962_11206# m2_34864_10986# 0.17fF
C621 a_27062_14178# ctop 3.58fF
C622 a_4974_7150# col_n[2] 0.28fF
C623 a_2346_14220# a_17934_14178# 0.35fF
C624 a_2346_18236# a_26970_18194# 0.35fF
C625 a_7986_13174# vcm 0.62fF
C626 m2_1732_4962# VDD 1.02fF
C627 a_10998_6146# VDD 0.52fF
C628 a_2346_5184# rowon_n[3] 0.26fF
C629 a_1962_13214# col[29] 0.11fF
C630 a_15014_7150# a_15014_6146# 1.00fF
C631 a_31990_7150# a_32082_7150# 0.26fF
C632 a_23046_3134# col_n[20] 0.28fF
C633 ctop rowoff_n[8] 0.60fF
C634 a_31078_14178# rowon_n[12] 0.14fF
C635 a_1962_11206# a_12002_11166# 0.27fF
C636 m2_22816_946# ctop 0.18fF
C637 a_20034_17190# col[17] 0.29fF
C638 a_1962_7190# vcm 6.95fF
C639 a_2346_16228# a_30986_16186# 0.35fF
C640 a_16018_16186# a_17022_16186# 0.97fF
C641 m2_1732_12994# row_n[11] 0.13fF
C642 a_21038_17190# vcm 0.60fF
C643 m2_9764_18014# VDD 0.93fF
C644 a_1962_18234# m2_24824_18014# 0.18fF
C645 a_24050_10162# VDD 0.52fF
C646 a_1962_8194# a_5278_8194# 0.14fF
C647 a_2346_8196# a_6982_8154# 0.19fF
C648 a_4882_8154# a_4974_8154# 0.26fF
C649 a_8990_14178# row_n[12] 0.17fF
C650 a_31078_2130# vcm 0.62fF
C651 a_1962_13214# a_25054_13174# 0.27fF
C652 a_9994_4138# rowoff_n[2] 0.10fF
C653 a_24050_4138# row_n[2] 0.17fF
C654 a_14314_11206# vcm 0.22fF
C655 a_23046_12170# rowoff_n[10] 0.10fF
C656 a_2346_13216# col[13] 0.15fF
C657 a_2346_18236# m2_19804_18014# 0.19fF
C658 a_1962_10202# a_18330_10202# 0.14fF
C659 a_28066_11166# a_28066_10162# 1.00fF
C660 a_2346_10204# a_20034_10162# 0.19fF
C661 a_1962_2170# col_n[27] 0.13fF
C662 a_20034_2130# rowoff_n[0] 0.10fF
C663 a_1962_15222# col_n[29] 0.13fF
C664 m2_1732_8978# m2_2160_9406# 0.16fF
C665 a_2966_15182# rowoff_n[13] 0.10fF
C666 a_27366_15222# vcm 0.22fF
C667 m2_8760_18014# m3_8892_18146# 2.78fF
C668 a_28066_17190# row_n[15] 0.17fF
C669 a_1962_9198# col[20] 0.11fF
C670 a_8990_9158# ctop 3.58fF
C671 a_21038_6146# col[18] 0.29fF
C672 a_16930_17190# VDD 0.24fF
C673 a_12002_2130# rowon_n[0] 0.14fF
C674 a_1962_12210# a_31382_12210# 0.14fF
C675 a_2346_12212# a_33086_12170# 0.19fF
C676 a_17934_12170# a_18026_12170# 0.26fF
C677 col_n[13] row_n[6] 0.23fF
C678 col_n[19] row_n[9] 0.23fF
C679 col_n[9] row_n[4] 0.23fF
C680 VDD en_bit_n[1] 0.15fF
C681 col_n[3] row_n[1] 0.23fF
C682 col_n[17] row_n[8] 0.23fF
C683 col_n[15] row_n[7] 0.23fF
C684 col_n[1] row_n[0] 0.22fF
C685 sample ctop 0.11fF
C686 col_n[21] row_n[10] 0.23fF
C687 col_n[31] row_n[15] 0.23fF
C688 col_n[5] row_n[2] 0.23fF
C689 col_n[23] row_n[11] 0.23fF
C690 col_n[25] row_n[12] 0.23fF
C691 col_n[11] row_n[5] 0.23fF
C692 col_n[27] row_n[13] 0.23fF
C693 col_n[7] row_n[3] 0.23fF
C694 col_n[29] row_n[14] 0.23fF
C695 a_26970_2130# VDD 0.23fF
C696 a_2346_4180# a_9902_4138# 0.35fF
C697 a_32082_11166# m2_32280_11414# 0.16fF
C698 a_22042_13174# ctop 3.58fF
C699 m3_34996_7102# m3_34996_6098# 0.22fF
C700 a_19942_18194# m2_19804_18014# 0.16fF
C701 a_8898_10162# rowoff_n[8] 0.24fF
C702 a_16018_15182# rowon_n[13] 0.14fF
C703 a_10906_13174# rowoff_n[11] 0.24fF
C704 a_1962_1166# a_3970_1126# 0.27fF
C705 a_2346_9200# col[4] 0.15fF
C706 a_5978_5142# VDD 0.52fF
C707 a_31078_5142# rowon_n[3] 0.14fF
C708 a_2966_13174# m2_3164_13422# 0.16fF
C709 a_12002_6146# a_13006_6146# 0.97fF
C710 a_2346_6188# a_22954_6146# 0.35fF
C711 a_1962_18234# col_n[3] 0.13fF
C712 a_18938_8154# rowoff_n[6] 0.24fF
C713 a_1962_11206# col_n[20] 0.13fF
C714 a_21038_8154# col_n[18] 0.28fF
C715 a_14010_16186# a_14010_15182# 1.00fF
C716 a_30986_16186# a_31078_16186# 0.26fF
C717 a_1962_1166# m2_8760_946# 0.18fF
C718 m2_34864_12994# m2_34864_11990# 0.99fF
C719 a_24962_17190# rowoff_n[15] 0.24fF
C720 a_16018_16186# vcm 0.62fF
C721 a_8990_5142# row_n[3] 0.17fF
C722 a_1962_5182# col[11] 0.11fF
C723 a_1962_3174# a_17022_3134# 0.27fF
C724 a_28978_6146# rowoff_n[4] 0.24fF
C725 a_19030_9158# VDD 0.52fF
C726 m2_16792_946# ctop 0.22fF
C727 a_26058_1126# vcm 0.12fF
C728 a_2966_15182# col[0] 0.29fF
C729 a_2346_4180# col[31] 0.15fF
C730 a_9294_10202# vcm 0.22fF
C731 a_2346_17232# a_4974_17190# 0.19fF
C732 a_1962_17230# a_3270_17230# 0.14fF
C733 m2_33860_946# ctop 0.68fF
C734 a_29070_12170# m2_29268_12418# 0.16fF
C735 a_1962_5182# a_30074_5142# 0.27fF
C736 a_32082_13174# VDD 0.52fF
C737 a_25054_10162# a_26058_10162# 0.97fF
C738 a_3970_1126# col_n[1] 0.31fF
C739 a_28066_8154# row_n[6] 0.17fF
C740 a_22346_14218# vcm 0.22fF
C741 a_13918_2130# a_14010_2130# 0.26fF
C742 a_1962_2170# a_23350_2170# 0.14fF
C743 a_2346_2172# a_25054_2130# 0.19fF
C744 col[2] rowoff_n[5] 0.11fF
C745 col[1] rowoff_n[4] 0.11fF
C746 col[4] rowoff_n[7] 0.11fF
C747 col[6] rowoff_n[9] 0.11fF
C748 col[5] rowoff_n[8] 0.11fF
C749 a_3970_8154# ctop 3.57fF
C750 m2_34864_17010# m3_34996_18146# 0.15fF
C751 col[0] rowoff_n[3] 0.11fF
C752 col[3] rowoff_n[6] 0.11fF
C753 a_34090_15182# m2_34864_15002# 0.96fF
C754 a_11910_16186# VDD 0.23fF
C755 a_1962_7190# col_n[11] 0.13fF
C756 a_19030_11166# col[16] 0.29fF
C757 m2_9764_18014# col_n[7] 0.25fF
C758 a_2346_2172# m2_1732_1950# 0.12fF
C759 a_2966_17190# vcm 0.60fF
C760 a_21950_1126# VDD 0.44fF
C761 a_1962_1166# col[2] 0.11fF
C762 a_1962_14218# col[4] 0.11fF
C763 a_17022_12170# ctop 3.58fF
C764 a_16018_6146# rowon_n[4] 0.14fF
C765 a_2346_13216# a_7894_13174# 0.35fF
C766 a_2346_13216# col[24] 0.15fF
C767 a_35002_5142# VDD 0.29fF
C768 a_26970_6146# a_27062_6146# 0.26fF
C769 a_9994_6146# a_9994_5142# 1.00fF
C770 a_26058_13174# m2_26256_13422# 0.16fF
C771 m3_1864_16138# VDD 0.25fF
C772 a_30074_16186# ctop 3.57fF
C773 a_2346_15224# a_20946_15182# 0.35fF
C774 a_10998_15182# a_12002_15182# 0.97fF
C775 a_1962_9198# col[31] 0.11fF
C776 a_10998_15182# vcm 0.62fF
C777 a_19030_13174# col_n[16] 0.28fF
C778 a_32082_2130# m3_31984_1078# 0.15fF
C779 a_14010_8154# VDD 0.52fF
C780 a_1962_3174# col_n[2] 0.13fF
C781 col_n[26] row_n[7] 0.23fF
C782 col_n[16] row_n[2] 0.23fF
C783 col_n[14] row_n[1] 0.23fF
C784 col_n[30] row_n[9] 0.23fF
C785 col_n[18] row_n[3] 0.23fF
C786 col_n[9] ctop 2.02fF
C787 col_n[20] row_n[4] 0.23fF
C788 a_1962_16226# col_n[4] 0.13fF
C789 vcm col[3] 5.84fF
C790 VDD col[7] 4.17fF
C791 col_n[28] row_n[8] 0.23fF
C792 col_n[1] col[2] 6.01fF
C793 col_n[22] row_n[5] 0.23fF
C794 col_n[12] row_n[0] 0.23fF
C795 col_n[24] row_n[6] 0.23fF
C796 a_1962_12210# a_15014_12170# 0.27fF
C797 a_4274_9198# vcm 0.22fF
C798 a_2346_17232# a_33998_17190# 0.35fF
C799 m2_8760_946# m3_9896_1078# 0.13fF
C800 a_13006_9158# row_n[7] 0.17fF
C801 a_27062_12170# VDD 0.52fF
C802 m3_21944_18146# m3_22948_18146# 0.22fF
C803 a_2346_9200# a_9994_9158# 0.19fF
C804 a_23046_10162# a_23046_9158# 1.00fF
C805 a_1962_9198# a_8290_9198# 0.14fF
C806 a_34090_4138# vcm 0.62fF
C807 a_1962_14218# a_28066_14178# 0.27fF
C808 a_11910_3134# rowoff_n[1] 0.24fF
C809 a_2346_9200# col[15] 0.15fF
C810 m2_1732_17010# sample 0.19fF
C811 m2_34864_10986# ctop 0.17fF
C812 a_26970_14178# rowoff_n[12] 0.24fF
C813 a_17326_13214# vcm 0.22fF
C814 m2_34864_13998# m3_34996_15134# 0.15fF
C815 a_1962_18234# col_n[14] 0.13fF
C816 a_2966_6146# a_3970_6146# 0.97fF
C817 a_23046_14178# m2_23244_14426# 0.16fF
C818 a_1962_11206# col_n[31] 0.13fF
C819 a_6890_15182# VDD 0.23fF
C820 a_1962_11206# a_21342_11206# 0.14fF
C821 a_12914_11166# a_13006_11166# 0.26fF
C822 a_2346_11208# a_23046_11166# 0.19fF
C823 m2_12776_946# a_13006_2130# 0.99fF
C824 a_20034_2130# col_n[17] 0.26fF
C825 a_1962_5182# col[22] 0.11fF
C826 a_32082_12170# row_n[10] 0.17fF
C827 a_30378_17230# vcm 0.22fF
C828 a_17022_16186# col[14] 0.29fF
C829 a_12002_11166# ctop 3.58fF
C830 a_2346_13216# a_2346_12212# 0.22fF
C831 a_1962_13214# a_35398_13214# 0.14fF
C832 a_29982_4138# VDD 0.23fF
C833 a_2346_5184# a_12914_5142# 0.35fF
C834 a_6982_5142# a_7986_5142# 0.97fF
C835 a_25054_15182# ctop 3.58fF
C836 a_20034_10162# rowon_n[8] 0.14fF
C837 a_9994_9158# rowoff_n[7] 0.10fF
C838 a_2346_5184# col[6] 0.15fF
C839 a_8990_15182# a_8990_14178# 1.00fF
C840 a_25966_15182# a_26058_15182# 0.26fF
C841 col[8] rowoff_n[0] 0.11fF
C842 col[10] rowoff_n[2] 0.11fF
C843 col[9] rowoff_n[1] 0.11fF
C844 col[16] rowoff_n[8] 0.11fF
C845 col[15] rowoff_n[7] 0.11fF
C846 col[17] rowoff_n[9] 0.11fF
C847 col[12] rowoff_n[4] 0.11fF
C848 col[11] rowoff_n[3] 0.11fF
C849 col[13] rowoff_n[5] 0.11fF
C850 col[14] rowoff_n[6] 0.11fF
C851 a_5978_14178# vcm 0.62fF
C852 a_14010_15182# rowoff_n[13] 0.10fF
C853 a_1962_2170# a_6982_2130# 0.27fF
C854 m2_22816_18014# m3_23952_18146# 0.13fF
C855 a_8990_7150# VDD 0.52fF
C856 a_1962_7190# col_n[22] 0.13fF
C857 a_20034_7150# rowoff_n[5] 0.10fF
C858 a_2346_7192# a_25966_7150# 0.35fF
C859 a_20034_15182# m2_20232_15430# 0.16fF
C860 a_18026_5142# col[15] 0.29fF
C861 a_1962_1166# col[13] 0.11fF
C862 a_1962_14218# col[15] 0.11fF
C863 a_22042_3134# m2_22240_3382# 0.16fF
C864 a_30074_5142# rowoff_n[3] 0.10fF
C865 a_19030_18194# vcm 0.12fF
C866 a_3878_1126# VDD 0.39fF
C867 a_1962_4178# a_20034_4138# 0.27fF
C868 a_22042_11166# VDD 0.52fF
C869 m3_11904_1078# m3_12908_1078# 0.22fF
C870 a_20034_9158# a_21038_9158# 0.97fF
C871 a_29070_3134# vcm 0.62fF
C872 col[1] rowoff_n[10] 0.11fF
C873 a_12306_12210# vcm 0.22fF
C874 a_1962_1166# a_13310_1166# 0.14fF
C875 m2_34864_10986# m3_34996_12122# 0.15fF
C876 a_17022_13174# row_n[11] 0.17fF
C877 a_1962_6186# a_33086_6146# 0.27fF
C878 m2_1732_15002# rowon_n[13] 0.11fF
C879 a_32082_3134# row_n[1] 0.17fF
C880 a_2346_15224# a_1962_15222# 2.62fF
C881 m2_22816_946# m3_22948_1078# 2.79fF
C882 a_25358_16226# vcm 0.22fF
C883 a_18026_7150# col_n[15] 0.28fF
C884 a_1962_3174# a_26362_3174# 0.14fF
C885 a_32082_4138# a_32082_3134# 1.00fF
C886 a_2346_3176# a_28066_3134# 0.19fF
C887 a_1962_3174# col_n[13] 0.13fF
C888 a_6982_10162# ctop 3.58fF
C889 col_n[25] row_n[1] 0.23fF
C890 col_n[31] row_n[4] 0.23fF
C891 col_n[27] row_n[2] 0.23fF
C892 VDD col[18] 4.17fF
C893 col_n[20] ctop 2.02fF
C894 col_n[23] row_n[0] 0.23fF
C895 vcm col[14] 5.84fF
C896 col_n[7] col[7] 0.72fF
C897 rowon_n[10] rowon_n[9] 0.15fF
C898 a_1962_16226# col_n[15] 0.13fF
C899 col_n[29] row_n[3] 0.23fF
C900 a_17022_16186# m2_17220_16434# 0.16fF
C901 a_14922_18194# VDD 0.34fF
C902 m2_4744_18014# vcm 0.28fF
C903 a_33086_13174# a_34090_13174# 0.97fF
C904 a_4974_11166# rowon_n[9] 0.14fF
C905 a_28978_11166# rowoff_n[9] 0.24fF
C906 a_1962_10202# col[6] 0.11fF
C907 a_19030_4138# m2_19228_4386# 0.16fF
C908 a_24962_3134# VDD 0.23fF
C909 m3_34996_15134# ctop 0.23fF
C910 a_33086_17190# col[30] 0.29fF
C911 a_4974_5142# a_4974_4138# 1.00fF
C912 a_21950_5142# a_22042_5142# 0.26fF
C913 a_20034_14178# ctop 3.58fF
C914 m2_27836_946# m2_28840_946# 0.96fF
C915 a_2346_9200# col[26] 0.15fF
C916 a_2346_14220# a_10906_14178# 0.35fF
C917 a_5978_14178# a_6982_14178# 0.97fF
C918 a_2346_18236# a_19942_18194# 0.35fF
C919 a_1962_18234# col_n[25] 0.13fF
C920 a_1962_2170# a_34394_2170# 0.14fF
C921 m2_1732_15002# m3_1864_15134# 2.76fF
C922 a_3970_6146# VDD 0.52fF
C923 a_3878_11166# a_3970_11166# 0.26fF
C924 a_1962_11206# a_4974_11166# 0.27fF
C925 a_24050_14178# rowon_n[12] 0.14fF
C926 a_2346_16228# a_23958_16186# 0.35fF
C927 a_16018_10162# col[13] 0.29fF
C928 a_14010_17190# vcm 0.60fF
C929 a_1962_18234# m2_10768_18014# 0.18fF
C930 a_1962_12210# col_n[6] 0.13fF
C931 a_17022_10162# VDD 0.52fF
C932 a_18026_9158# a_18026_8154# 1.00fF
C933 a_14010_17190# m2_14208_17438# 0.16fF
C934 a_24050_2130# vcm 0.62fF
C935 a_1962_13214# a_18026_13174# 0.27fF
C936 m2_24824_18014# col[22] 0.28fF
C937 a_34090_6146# col[31] 0.29fF
C938 a_17022_4138# row_n[2] 0.17fF
C939 a_7286_11206# vcm 0.22fF
C940 a_2874_4138# rowoff_n[2] 0.24fF
C941 a_16018_12170# rowoff_n[10] 0.10fF
C942 a_16018_5142# m2_16216_5390# 0.16fF
C943 m2_34864_7974# m3_34996_9110# 0.15fF
C944 a_35002_13174# m2_34864_12994# 0.16fF
C945 m3_13912_1078# VDD 0.14fF
C946 a_2346_18236# m2_5748_18014# 0.19fF
C947 a_30074_14178# VDD 0.52fF
C948 a_2346_5184# col[17] 0.15fF
C949 a_1962_10202# a_11302_10202# 0.14fF
C950 a_7894_10162# a_7986_10162# 0.26fF
C951 a_2346_10204# a_13006_10162# 0.19fF
C952 a_13006_2130# rowoff_n[0] 0.10fF
C953 col[26] rowoff_n[7] 0.11fF
C954 col[20] rowoff_n[1] 0.11fF
C955 col[22] rowoff_n[3] 0.11fF
C956 col[28] rowoff_n[9] 0.11fF
C957 col[27] rowoff_n[8] 0.11fF
C958 col[21] rowoff_n[2] 0.11fF
C959 col[24] rowoff_n[5] 0.11fF
C960 col[23] rowoff_n[4] 0.11fF
C961 col[19] rowoff_n[0] 0.11fF
C962 col[25] rowoff_n[6] 0.11fF
C963 a_1962_15222# a_31078_15182# 0.27fF
C964 a_30074_16186# rowoff_n[14] 0.10fF
C965 m2_32856_18014# ctop 0.18fF
C966 a_20338_15222# vcm 0.22fF
C967 a_29070_3134# a_30074_3134# 0.97fF
C968 a_21038_17190# row_n[15] 0.17fF
C969 a_16018_12170# col_n[13] 0.28fF
C970 a_4974_2130# rowon_n[0] 0.14fF
C971 a_9902_17190# VDD 0.24fF
C972 a_1962_1166# col[24] 0.11fF
C973 a_1962_12210# a_24354_12210# 0.14fF
C974 a_31078_13174# a_31078_12170# 1.00fF
C975 a_2346_12212# a_26058_12170# 0.19fF
C976 a_1962_14218# col[26] 0.11fF
C977 a_19942_2130# VDD 0.23fF
C978 a_34090_8154# col_n[31] 0.28fF
C979 a_15014_13174# ctop 3.58fF
C980 m3_34996_14130# m3_34996_13126# 0.22fF
C981 m2_29844_946# m3_30980_1078# 0.13fF
C982 col[12] rowoff_n[10] 0.11fF
C983 a_3970_14178# a_3970_13174# 1.00fF
C984 a_20946_14178# a_21038_14178# 0.26fF
C985 a_8990_15182# rowon_n[13] 0.14fF
C986 a_13006_6146# m2_13204_6394# 0.16fF
C987 m2_1732_11990# m3_1864_12122# 2.76fF
C988 a_32994_6146# VDD 0.23fF
C989 a_24050_5142# rowon_n[3] 0.14fF
C990 a_2346_6188# a_15926_6146# 0.35fF
C991 a_28066_17190# ctop 3.39fF
C992 a_2346_1168# col[8] 0.14fF
C993 a_11910_8154# rowoff_n[6] 0.24fF
C994 a_2346_14220# col[10] 0.15fF
C995 a_8990_17190# m3_8892_18146# 0.15fF
C996 a_1962_3174# col_n[24] 0.13fF
C997 col_n[12] col[13] 5.98fF
C998 rowon_n[7] row_n[7] 19.75fF
C999 col_n[31] ctop 1.93fF
C1000 vcm col[25] 5.84fF
C1001 VDD col[29] 4.18fF
C1002 a_8990_16186# vcm 0.62fF
C1003 a_17934_17190# rowoff_n[15] 0.24fF
C1004 a_1962_16226# col_n[26] 0.13fF
C1005 m2_34864_17010# VDD 1.05fF
C1006 a_21950_6146# rowoff_n[4] 0.24fF
C1007 a_1962_3174# a_9994_3134# 0.27fF
C1008 a_12002_9158# VDD 0.52fF
C1009 a_2966_16186# m2_1732_16006# 0.96fF
C1010 a_15014_8154# a_16018_8154# 0.97fF
C1011 a_2346_8196# a_28978_8154# 0.35fF
C1012 a_14010_15182# col[11] 0.29fF
C1013 a_1962_10202# col[17] 0.11fF
C1014 a_19030_1126# vcm 0.59fF
C1015 a_31990_4138# rowoff_n[2] 0.24fF
C1016 m2_9764_946# ctop 0.18fF
C1017 m2_34864_4962# m3_34996_6098# 0.15fF
C1018 a_32082_11166# col[29] 0.29fF
C1019 a_1962_5182# a_23046_5142# 0.27fF
C1020 a_25054_13174# VDD 0.52fF
C1021 a_32082_5142# vcm 0.62fF
C1022 a_21038_8154# row_n[6] 0.17fF
C1023 m2_1732_13998# ctop 0.17fF
C1024 a_15318_14218# vcm 0.22fF
C1025 a_9994_7150# m2_10192_7398# 0.16fF
C1026 a_1962_2170# a_16322_2170# 0.14fF
C1027 a_27062_3134# a_27062_2130# 1.00fF
C1028 a_2346_2172# a_18026_2130# 0.19fF
C1029 a_2346_10204# col[1] 0.15fF
C1030 a_4882_16186# VDD 0.23fF
C1031 a_28066_12170# a_29070_12170# 0.97fF
C1032 a_14010_17190# col_n[11] 0.28fF
C1033 a_1962_12210# col_n[17] 0.13fF
C1034 a_15014_4138# col[12] 0.29fF
C1035 a_28370_18234# vcm 0.22fF
C1036 a_14922_1126# VDD 0.44fF
C1037 a_1962_4178# a_29374_4178# 0.14fF
C1038 a_2346_4180# a_31078_4138# 0.19fF
C1039 a_16930_4138# a_17022_4138# 0.26fF
C1040 a_9994_12170# ctop 3.58fF
C1041 a_8990_6146# rowon_n[4] 0.14fF
C1042 a_1962_6186# col[8] 0.11fF
C1043 a_32082_13174# col_n[29] 0.28fF
C1044 a_30074_10162# rowoff_n[8] 0.10fF
C1045 a_32082_13174# rowoff_n[11] 0.10fF
C1046 rowon_n[13] rowoff_n[13] 20.27fF
C1047 m2_1732_8978# m3_1864_9110# 2.76fF
C1048 a_2346_5184# col[28] 0.15fF
C1049 a_27974_5142# VDD 0.23fF
C1050 m3_9896_18146# VDD 0.25fF
C1051 col[30] rowoff_n[0] 0.11fF
C1052 col[31] rowoff_n[1] 0.11fF
C1053 a_23046_16186# ctop 3.57fF
C1054 a_2346_15224# a_13918_15182# 0.35fF
C1055 a_3970_15182# vcm 0.62fF
C1056 a_6982_8154# m2_7180_8402# 0.16fF
C1057 a_2966_17190# row_n[15] 0.16fF
C1058 a_6982_8154# VDD 0.52fF
C1059 a_28066_9158# rowon_n[7] 0.14fF
C1060 a_15014_6146# col_n[12] 0.28fF
C1061 a_29982_8154# a_30074_8154# 0.26fF
C1062 a_13006_8154# a_13006_7150# 1.00fF
C1063 a_1962_18234# a_31382_18234# 0.14fF
C1064 a_1962_12210# a_7986_12170# 0.27fF
C1065 m2_11772_946# col[9] 0.39fF
C1066 a_2346_17232# a_26970_17190# 0.35fF
C1067 a_14010_17190# a_15014_17190# 0.97fF
C1068 a_1962_8194# col_n[8] 0.13fF
C1069 m2_33860_18014# m2_34864_18014# 0.96fF
C1070 a_35494_3496# VDD 0.11fF
C1071 a_33086_2130# col_n[30] 0.29fF
C1072 m3_16924_1078# ctop 0.24fF
C1073 a_5978_9158# row_n[7] 0.17fF
C1074 col[23] rowoff_n[10] 0.11fF
C1075 a_20034_12170# VDD 0.52fF
C1076 m3_7888_18146# m3_8892_18146# 0.22fF
C1077 a_2346_9200# a_2874_9158# 0.35fF
C1078 a_30074_16186# col[27] 0.29fF
C1079 a_1962_15222# col[1] 0.11fF
C1080 a_27062_4138# vcm 0.62fF
C1081 m2_1732_3958# row_n[2] 0.13fF
C1082 a_1962_14218# a_21038_14178# 0.27fF
C1083 a_4882_3134# rowoff_n[1] 0.24fF
C1084 a_10298_13214# vcm 0.22fF
C1085 a_19942_14178# rowoff_n[12] 0.24fF
C1086 a_24050_2130# a_25054_2130# 0.97fF
C1087 a_2346_1168# col[19] 0.14fF
C1088 a_2346_14220# col[21] 0.15fF
C1089 a_33086_16186# VDD 0.52fF
C1090 a_1962_11206# a_14314_11206# 0.14fF
C1091 a_2346_11208# a_16018_11166# 0.19fF
C1092 a_26058_12170# a_26058_11166# 1.00fF
C1093 col_n[18] col[18] 0.72fF
C1094 rowon_n[10] ctop 1.40fF
C1095 a_1962_16226# a_34090_16186# 0.27fF
C1096 a_25054_12170# row_n[10] 0.17fF
C1097 a_23350_17230# vcm 0.22fF
C1098 col[7] rowoff_n[11] 0.11fF
C1099 a_3878_6146# rowoff_n[4] 0.24fF
C1100 a_3970_9158# m2_4168_9406# 0.16fF
C1101 a_4974_11166# ctop 3.58fF
C1102 a_1962_10202# col[28] 0.11fF
C1103 a_13006_9158# col[10] 0.29fF
C1104 a_33390_2170# vcm 0.22fF
C1105 a_1962_13214# a_27366_13214# 0.14fF
C1106 a_15926_13174# a_16018_13174# 0.26fF
C1107 a_2346_13216# a_29070_13174# 0.19fF
C1108 a_1962_4178# col_n[0] 0.13fF
C1109 a_1962_17230# col_n[1] 0.13fF
C1110 m2_1732_5966# m3_1864_6098# 2.76fF
C1111 a_31078_5142# col[28] 0.29fF
C1112 a_22954_4138# VDD 0.23fF
C1113 a_2346_5184# a_5886_5142# 0.35fF
C1114 a_1962_12210# m2_34864_11990# 0.17fF
C1115 a_18026_15182# ctop 3.58fF
C1116 m2_2736_946# vcm 0.41fF
C1117 a_13006_10162# rowon_n[8] 0.14fF
C1118 a_2874_9158# rowoff_n[7] 0.24fF
C1119 a_2966_8154# row_n[6] 0.16fF
C1120 a_6982_15182# rowoff_n[13] 0.10fF
C1121 a_2346_10204# col[12] 0.15fF
C1122 m2_13780_18014# m3_13912_18146# 2.78fF
C1123 a_13006_7150# rowoff_n[5] 0.10fF
C1124 a_9994_7150# a_10998_7150# 0.97fF
C1125 a_2346_7192# a_18938_7150# 0.35fF
C1126 a_1962_12210# col_n[28] 0.13fF
C1127 a_13006_11166# col_n[10] 0.28fF
C1128 a_12002_17190# a_12002_16186# 1.00fF
C1129 a_28978_17190# a_29070_17190# 0.26fF
C1130 m2_1732_16006# m2_1732_15002# 0.99fF
C1131 a_23046_5142# rowoff_n[3] 0.10fF
C1132 a_12002_18194# vcm 0.12fF
C1133 a_1962_4178# a_13006_4138# 0.27fF
C1134 a_1962_6186# col[19] 0.11fF
C1135 a_32082_13174# rowon_n[11] 0.14fF
C1136 a_15014_11166# VDD 0.52fF
C1137 a_2346_9200# a_31990_9158# 0.35fF
C1138 a_31078_7150# col_n[28] 0.28fF
C1139 a_22042_3134# vcm 0.62fF
C1140 a_33086_3134# rowoff_n[1] 0.10fF
C1141 a_5278_12210# vcm 0.22fF
C1142 a_1962_1166# a_6282_1166# 0.14fF
C1143 a_9994_13174# row_n[11] 0.17fF
C1144 a_1962_6186# a_26058_6146# 0.27fF
C1145 a_28066_15182# VDD 0.52fF
C1146 m2_34864_6970# vcm 0.51fF
C1147 a_23046_11166# a_24050_11166# 0.97fF
C1148 a_25054_3134# row_n[1] 0.17fF
C1149 a_35094_7150# vcm 0.12fF
C1150 a_18330_16226# vcm 0.22fF
C1151 a_2346_6188# col[3] 0.15fF
C1152 a_2346_3176# a_21038_3134# 0.19fF
C1153 a_1962_3174# a_19334_3174# 0.14fF
C1154 a_11910_3134# a_12002_3134# 0.26fF
C1155 a_2346_1168# m2_26832_946# 0.19fF
C1156 a_33086_2130# m2_32856_946# 0.99fF
C1157 a_7894_18194# VDD 0.33fF
C1158 a_1962_8194# col_n[19] 0.13fF
C1159 a_28370_1166# vcm 0.23fF
C1160 a_10998_14178# col[8] 0.29fF
C1161 a_21950_11166# rowoff_n[9] 0.24fF
C1162 a_29070_16186# row_n[14] 0.17fF
C1163 m2_1732_2954# m3_1864_3086# 2.76fF
C1164 a_17934_3134# VDD 0.23fF
C1165 m3_12908_18146# ctop 0.23fF
C1166 a_1962_2170# col[10] 0.11fF
C1167 a_2346_5184# a_34090_5142# 0.19fF
C1168 a_32082_12170# m2_32280_12418# 0.16fF
C1169 a_1962_5182# a_32386_5182# 0.14fF
C1170 a_1962_15222# col[12] 0.11fF
C1171 a_13006_14178# ctop 3.58fF
C1172 a_29070_10162# col[26] 0.29fF
C1173 a_31990_9158# rowoff_n[7] 0.24fF
C1174 a_1962_14218# a_2966_14178# 0.27fF
C1175 a_2346_1168# col[30] 0.14fF
C1176 a_2346_18236# a_12914_18194# 0.35fF
C1177 a_2346_18236# col[4] 0.14fF
C1178 a_30986_7150# VDD 0.23fF
C1179 a_7986_7150# a_7986_6146# 1.00fF
C1180 a_2966_14178# m2_3164_14426# 0.16fF
C1181 a_24962_7150# a_25054_7150# 0.26fF
C1182 row_n[5] ctop 1.65fF
C1183 col_n[23] col[24] 5.98fF
C1184 a_17022_14178# rowon_n[12] 0.14fF
C1185 col[18] rowoff_n[11] 0.11fF
C1186 a_8990_16186# a_9994_16186# 0.97fF
C1187 a_2346_16228# a_16930_16186# 0.35fF
C1188 m2_1732_8978# sample_n 0.15fF
C1189 a_4974_2130# m2_5172_2378# 0.16fF
C1190 a_32082_4138# rowon_n[2] 0.14fF
C1191 a_2346_2172# ctop 1.36fF
C1192 a_6982_17190# vcm 0.60fF
C1193 a_10998_16186# col_n[8] 0.28fF
C1194 a_2966_3134# m3_1864_3086# 0.14fF
C1195 a_12002_3134# col[9] 0.29fF
C1196 a_9994_10162# VDD 0.52fF
C1197 a_1962_4178# col_n[10] 0.13fF
C1198 a_17022_2130# vcm 0.62fF
C1199 a_1962_13214# a_10998_13174# 0.27fF
C1200 a_1962_17230# col_n[12] 0.13fF
C1201 m2_34864_3958# m2_35292_4386# 0.16fF
C1202 a_9994_4138# row_n[2] 0.17fF
C1203 a_29070_12170# col_n[26] 0.28fF
C1204 a_8990_12170# rowoff_n[10] 0.10fF
C1205 a_19030_1126# a_20034_1126# 0.97fF
C1206 a_2966_14178# col_n[0] 0.28fF
C1207 a_1962_11206# col[3] 0.11fF
C1208 m3_34996_9110# VDD 0.26fF
C1209 a_29070_13174# m2_29268_13422# 0.16fF
C1210 a_23046_14178# VDD 0.52fF
C1211 a_21038_11166# a_21038_10162# 1.00fF
C1212 a_2346_10204# a_5978_10162# 0.19fF
C1213 a_1962_10202# a_4274_10202# 0.14fF
C1214 a_5978_2130# rowoff_n[0] 0.10fF
C1215 col[2] rowoff_n[12] 0.11fF
C1216 a_30074_6146# vcm 0.62fF
C1217 a_1962_15222# a_24050_15182# 0.27fF
C1218 a_2346_10204# col[23] 0.15fF
C1219 a_13310_15222# vcm 0.22fF
C1220 m2_18800_18014# ctop 0.18fF
C1221 a_23046_16186# rowoff_n[14] 0.10fF
C1222 a_29982_1126# m2_29844_946# 0.16fF
C1223 a_14010_17190# row_n[15] 0.17fF
C1224 a_34090_16186# m2_34864_16006# 0.96fF
C1225 a_2346_17232# VDD 32.69fF
C1226 a_1962_12210# a_17326_12210# 0.14fF
C1227 a_2346_12212# a_19030_12170# 0.19fF
C1228 a_10906_12170# a_10998_12170# 0.26fF
C1229 a_29070_7150# row_n[5] 0.17fF
C1230 a_12002_5142# col_n[9] 0.28fF
C1231 a_2346_3176# m2_1732_2954# 0.12fF
C1232 a_1962_6186# col[30] 0.11fF
C1233 a_12914_2130# VDD 0.23fF
C1234 a_32082_5142# a_33086_5142# 0.97fF
C1235 a_7986_13174# ctop 3.58fF
C1236 m2_3740_18014# col_n[1] 0.25fF
C1237 a_1962_13214# col_n[3] 0.13fF
C1238 a_1962_14218# a_30378_14218# 0.14fF
C1239 a_34090_15182# a_34090_14178# 1.00fF
C1240 a_2346_14220# a_32082_14178# 0.19fF
C1241 a_27062_15182# col[24] 0.29fF
C1242 a_1962_7190# ctop 1.49fF
C1243 a_25966_6146# VDD 0.23fF
C1244 a_17022_5142# rowon_n[3] 0.14fF
C1245 a_2346_6188# a_8898_6146# 0.35fF
C1246 a_4974_6146# a_5978_6146# 0.97fF
C1247 a_26058_14178# m2_26256_14426# 0.16fF
C1248 a_21038_17190# ctop 3.39fF
C1249 a_4882_8154# rowoff_n[6] 0.24fF
C1250 m2_21812_946# col[19] 0.39fF
C1251 a_23958_16186# a_24050_16186# 0.26fF
C1252 a_6982_16186# a_6982_15182# 1.00fF
C1253 a_2346_6188# col[14] 0.15fF
C1254 a_31078_2130# ctop 3.39fF
C1255 a_10906_17190# rowoff_n[15] 0.24fF
C1256 a_34394_17230# vcm 0.22fF
C1257 a_14922_6146# rowoff_n[4] 0.24fF
C1258 a_2346_3176# a_2966_3134# 0.21fF
C1259 a_4974_9158# VDD 0.52fF
C1260 a_1962_8194# col_n[30] 0.13fF
C1261 a_2346_8196# a_21950_8154# 0.35fF
C1262 a_12002_1126# vcm 0.12fF
C1263 a_9994_8154# col[7] 0.29fF
C1264 a_24962_4138# rowoff_n[2] 0.24fF
C1265 a_3878_11166# rowoff_n[9] 0.24fF
C1266 a_1962_2170# col[21] 0.11fF
C1267 a_1962_15222# col[23] 0.11fF
C1268 a_27062_17190# col_n[24] 0.28fF
C1269 a_1962_5182# a_16018_5142# 0.27fF
C1270 a_18026_13174# VDD 0.52fF
C1271 a_28066_4138# col[25] 0.29fF
C1272 a_2346_10204# a_35002_10162# 0.35fF
C1273 a_18026_10162# a_19030_10162# 0.97fF
C1274 a_35002_2130# rowoff_n[0] 0.24fF
C1275 a_25054_5142# vcm 0.62fF
C1276 a_14010_8154# row_n[6] 0.17fF
C1277 a_8290_14218# vcm 0.22fF
C1278 a_2346_18236# col[15] 0.14fF
C1279 a_6890_2130# a_6982_2130# 0.26fF
C1280 a_1962_2170# a_9294_2170# 0.14fF
C1281 a_2346_2172# a_10998_2130# 0.19fF
C1282 m2_27836_18014# m3_28972_18146# 0.13fF
C1283 sw ctop 0.23fF
C1284 col_n[29] col[29] 0.78fF
C1285 a_23046_15182# m2_23244_15430# 0.16fF
C1286 a_1962_7190# a_29070_7150# 0.27fF
C1287 a_31078_17190# VDD 0.55fF
C1288 col[29] rowoff_n[11] 0.11fF
C1289 a_2346_2172# col[5] 0.15fF
C1290 a_2346_15224# col[7] 0.15fF
C1291 a_25054_3134# m2_25252_3382# 0.16fF
C1292 a_9994_10162# col_n[7] 0.28fF
C1293 a_21342_18234# vcm 0.22fF
C1294 a_7894_1126# VDD 0.44fF
C1295 a_2346_4180# a_24050_4138# 0.19fF
C1296 a_1962_4178# a_22346_4178# 0.14fF
C1297 a_30074_5142# a_30074_4138# 1.00fF
C1298 m2_1732_5966# rowon_n[4] 0.11fF
C1299 a_1962_4178# col_n[21] 0.13fF
C1300 a_1962_17230# col_n[23] 0.13fF
C1301 a_6982_17190# m2_6752_18014# 1.00fF
C1302 a_33086_11166# row_n[9] 0.17fF
C1303 a_31382_3174# vcm 0.22fF
C1304 a_31078_14178# a_32082_14178# 0.97fF
C1305 a_23046_10162# rowoff_n[8] 0.10fF
C1306 a_28066_6146# col_n[25] 0.28fF
C1307 a_25054_13174# rowoff_n[11] 0.10fF
C1308 a_1962_11206# col[14] 0.11fF
C1309 a_20946_5142# VDD 0.23fF
C1310 a_19942_6146# a_20034_6146# 0.26fF
C1311 m2_25828_946# VDD 0.62fF
C1312 col[13] rowoff_n[12] 0.11fF
C1313 a_16018_16186# ctop 3.57fF
C1314 a_33086_8154# rowoff_n[6] 0.10fF
C1315 a_3970_15182# a_4974_15182# 0.97fF
C1316 a_2346_15224# a_6890_15182# 0.35fF
C1317 m2_14784_946# m2_15212_1374# 0.16fF
C1318 a_21038_9158# rowon_n[7] 0.14fF
C1319 a_33998_9158# VDD 0.23fF
C1320 a_20034_16186# m2_20232_16434# 0.16fF
C1321 a_1962_18234# a_24354_18234# 0.14fF
C1322 a_2346_17232# a_19942_17190# 0.35fF
C1323 a_3970_1126# en_C0_n 0.26fF
C1324 a_22042_4138# m2_22240_4386# 0.16fF
C1325 m2_26832_18014# m2_27836_18014# 0.96fF
C1326 a_7986_13174# col[5] 0.29fF
C1327 m3_1864_7102# ctop 0.23fF
C1328 a_1962_13214# col_n[14] 0.13fF
C1329 a_13006_12170# VDD 0.52fF
C1330 m2_31852_946# m2_32280_1374# 0.16fF
C1331 a_32994_10162# a_33086_10162# 0.26fF
C1332 a_16018_10162# a_16018_9158# 1.00fF
C1333 a_20034_4138# vcm 0.62fF
C1334 a_1962_14218# a_14010_14178# 0.27fF
C1335 a_26058_9158# col[23] 0.29fF
C1336 a_1962_7190# col[5] 0.11fF
C1337 a_12914_14178# rowoff_n[12] 0.24fF
C1338 a_3270_13214# vcm 0.22fF
C1339 a_2966_17190# ctop 3.24fF
C1340 a_26058_16186# VDD 0.52fF
C1341 a_2346_6188# col[25] 0.15fF
C1342 m2_1732_9982# vcm 0.45fF
C1343 a_2346_11208# a_8990_11166# 0.19fF
C1344 a_1962_11206# a_7286_11206# 0.14fF
C1345 a_5886_11166# a_5978_11166# 0.26fF
C1346 a_33086_8154# vcm 0.62fF
C1347 a_1962_16226# a_27062_16186# 0.27fF
C1348 a_5978_2130# m2_5748_946# 0.99fF
C1349 a_18026_12170# row_n[10] 0.17fF
C1350 a_16322_17230# vcm 0.22fF
C1351 a_27062_4138# a_28066_4138# 0.97fF
C1352 a_33086_2130# row_n[0] 0.17fF
C1353 a_7986_15182# col_n[5] 0.28fF
C1354 a_17022_17190# m2_17220_17438# 0.16fF
C1355 a_26058_17190# m2_25828_18014# 1.00fF
C1356 a_2346_8196# a_3878_8154# 0.35fF
C1357 a_2874_8154# a_2966_8154# 0.26fF
C1358 a_2966_12170# m3_1864_12122# 0.14fF
C1359 a_8990_2130# col[6] 0.29fF
C1360 a_2346_13216# a_22042_13174# 0.19fF
C1361 a_26362_2170# vcm 0.22fF
C1362 a_1962_13214# a_20338_13214# 0.14fF
C1363 a_29070_14178# a_29070_13174# 1.00fF
C1364 a_19030_5142# m2_19228_5390# 0.16fF
C1365 a_15926_4138# VDD 0.23fF
C1366 a_26058_11166# col_n[23] 0.28fF
C1367 m3_28972_1078# VDD 0.14fF
C1368 a_1962_9198# col_n[5] 0.13fF
C1369 a_10998_15182# ctop 3.58fF
C1370 a_5978_10162# rowon_n[8] 0.14fF
C1371 a_2346_18236# col[26] 0.14fF
C1372 a_1962_15222# a_33390_15222# 0.14fF
C1373 a_18938_15182# a_19030_15182# 0.26fF
C1374 ctop col[3] 1.98fF
C1375 m2_4744_18014# m3_3872_18146# 0.13fF
C1376 a_28978_8154# VDD 0.23fF
C1377 a_5978_7150# rowoff_n[5] 0.10fF
C1378 a_2346_7192# a_11910_7150# 0.35fF
C1379 a_2346_2172# col[16] 0.15fF
C1380 a_2346_15224# col[18] 0.15fF
C1381 a_16018_5142# rowoff_n[3] 0.10fF
C1382 a_8990_4138# col_n[6] 0.28fF
C1383 a_4974_18194# vcm 0.12fF
C1384 a_34090_4138# ctop 3.42fF
C1385 a_1962_4178# a_5978_4138# 0.27fF
C1386 a_25054_13174# rowon_n[11] 0.14fF
C1387 a_7986_11166# VDD 0.52fF
C1388 a_2346_9200# a_24962_9158# 0.35fF
C1389 a_13006_9158# a_14010_9158# 0.97fF
C1390 a_1962_18234# col[8] 0.11fF
C1391 a_1962_11206# col[25] 0.11fF
C1392 a_15014_3134# vcm 0.62fF
C1393 a_26058_3134# rowoff_n[1] 0.10fF
C1394 a_16018_6146# m2_16216_6394# 0.16fF
C1395 col[24] rowoff_n[12] 0.11fF
C1396 a_1962_5182# VDD 2.73fF
C1397 a_24050_14178# col[21] 0.29fF
C1398 a_1962_6186# a_19030_6146# 0.27fF
C1399 a_35002_14178# m2_34864_13998# 0.16fF
C1400 a_21038_15182# VDD 0.52fF
C1401 m2_18800_18014# col[16] 0.28fF
C1402 a_2966_11166# a_2966_10162# 1.00fF
C1403 a_12002_17190# m3_11904_18146# 0.15fF
C1404 a_18026_3134# row_n[1] 0.17fF
C1405 a_28066_7150# vcm 0.62fF
C1406 a_1962_1166# m2_1732_946# 0.15fF
C1407 a_11302_16226# vcm 0.22fF
C1408 a_1962_3174# a_12306_3174# 0.14fF
C1409 a_2346_3176# a_14010_3134# 0.19fF
C1410 a_25054_4138# a_25054_3134# 1.00fF
C1411 a_2966_9158# rowon_n[7] 0.13fF
C1412 a_1962_8194# a_32082_8154# 0.27fF
C1413 a_2346_11208# col[9] 0.15fF
C1414 a_21342_1166# vcm 0.23fF
C1415 a_26058_13174# a_27062_13174# 0.97fF
C1416 a_14922_11166# rowoff_n[9] 0.24fF
C1417 col[8] rowoff_n[13] 0.11fF
C1418 a_22042_16186# row_n[14] 0.17fF
C1419 a_6982_7150# col[4] 0.29fF
C1420 a_1962_13214# col_n[25] 0.13fF
C1421 a_10906_3134# VDD 0.23fF
C1422 a_1962_5182# a_25358_5182# 0.14fF
C1423 a_14922_5142# a_15014_5142# 0.26fF
C1424 a_2346_5184# a_27062_5142# 0.19fF
C1425 a_5978_14178# ctop 3.58fF
C1426 m2_8760_946# col[6] 0.39fF
C1427 a_24050_16186# col_n[21] 0.28fF
C1428 a_24962_9158# rowoff_n[7] 0.24fF
C1429 a_1962_7190# col[16] 0.11fF
C1430 a_35398_5182# vcm 0.23fF
C1431 a_25054_3134# col[22] 0.29fF
C1432 a_2346_18236# a_5886_18194# 0.35fF
C1433 a_28978_15182# rowoff_n[13] 0.24fF
C1434 a_13006_7150# m2_13204_7398# 0.16fF
C1435 a_23958_7150# VDD 0.23fF
C1436 a_35002_7150# rowoff_n[5] 0.24fF
C1437 a_9994_14178# rowon_n[12] 0.14fF
C1438 a_2346_16228# a_9902_16186# 0.35fF
C1439 a_25054_4138# rowon_n[2] 0.14fF
C1440 a_29070_3134# ctop 3.57fF
C1441 a_2874_10162# VDD 0.24fF
C1442 a_6982_9158# col_n[4] 0.28fF
C1443 a_2966_17190# m2_1732_17010# 0.96fF
C1444 a_10998_9158# a_10998_8154# 1.00fF
C1445 a_27974_9158# a_28066_9158# 0.26fF
C1446 a_2346_7192# col[0] 0.15fF
C1447 a_9994_2130# vcm 0.62fF
C1448 a_1962_13214# a_3970_13174# 0.27fF
C1449 a_1962_9198# col_n[16] 0.13fF
C1450 a_2346_1168# a_29982_1126# 0.35fF
C1451 a_25054_5142# col_n[22] 0.28fF
C1452 m3_24956_18146# VDD 0.24fF
C1453 a_29070_17190# rowon_n[15] 0.14fF
C1454 a_16018_14178# VDD 0.52fF
C1455 a_1962_3174# col[7] 0.11fF
C1456 ctop col[14] 1.98fF
C1457 a_1962_16226# col[9] 0.11fF
C1458 a_23046_6146# vcm 0.62fF
C1459 a_1962_15222# a_17022_15182# 0.27fF
C1460 a_16018_16186# rowoff_n[14] 0.10fF
C1461 a_6282_15222# vcm 0.22fF
C1462 m2_4744_18014# ctop 0.18fF
C1463 a_22042_3134# a_23046_3134# 0.97fF
C1464 a_9994_8154# m2_10192_8402# 0.16fF
C1465 a_2346_2172# col[27] 0.15fF
C1466 a_6982_17190# row_n[15] 0.17fF
C1467 a_2346_15224# col[29] 0.15fF
C1468 a_2346_12212# a_12002_12170# 0.19fF
C1469 a_24050_13174# a_24050_12170# 1.00fF
C1470 a_1962_12210# a_10298_12210# 0.14fF
C1471 m2_33860_18014# vcm 0.28fF
C1472 a_22042_7150# row_n[5] 0.17fF
C1473 a_2346_9200# vcm 0.40fF
C1474 a_1962_17230# a_30074_17190# 0.27fF
C1475 m2_4744_946# m3_4876_1078# 2.79fF
C1476 a_5886_2130# VDD 0.23fF
C1477 m3_31984_1078# ctop 0.23fF
C1478 a_1962_18234# col[19] 0.11fF
C1479 a_4974_12170# col[2] 0.29fF
C1480 a_5886_18194# m2_5748_18014# 0.16fF
C1481 a_29374_4178# vcm 0.22fF
C1482 a_2346_14220# a_25054_14178# 0.19fF
C1483 a_13918_14178# a_14010_14178# 0.26fF
C1484 a_1962_14218# a_23350_14218# 0.14fF
C1485 a_1962_1166# m2_22816_946# 0.18fF
C1486 a_1962_5182# col_n[7] 0.13fF
C1487 a_23046_8154# col[20] 0.29fF
C1488 a_18938_6146# VDD 0.23fF
C1489 a_9994_5142# rowon_n[3] 0.14fF
C1490 a_14010_17190# ctop 3.39fF
C1491 a_2966_15182# VDD 0.56fF
C1492 a_1962_12210# col[0] 0.11fF
C1493 a_24050_2130# ctop 3.39fF
C1494 m2_24824_18014# VDD 0.91fF
C1495 a_7894_6146# rowoff_n[4] 0.24fF
C1496 a_6982_9158# m2_7180_9406# 0.16fF
C1497 a_2346_11208# col[20] 0.15fF
C1498 a_31990_10162# VDD 0.23fF
C1499 a_7986_8154# a_8990_8154# 0.97fF
C1500 a_2346_8196# a_14922_8154# 0.35fF
C1501 a_4974_1126# vcm 0.12fF
C1502 col[19] rowoff_n[13] 0.11fF
C1503 a_4974_14178# col_n[2] 0.28fF
C1504 a_17934_4138# rowoff_n[2] 0.24fF
C1505 a_30986_12170# rowoff_n[10] 0.24fF
C1506 sample_n rowoff_n[4] 0.38fF
C1507 vcm rowoff_n[7] 0.20fF
C1508 VDD rowoff_n[3] 1.17fF
C1509 a_29070_8154# rowon_n[6] 0.14fF
C1510 a_1962_5182# a_8990_5142# 0.27fF
C1511 a_1962_7190# col[27] 0.11fF
C1512 a_2346_18236# m2_34864_18014# 0.17fF
C1513 a_10998_13174# VDD 0.52fF
C1514 m2_10768_946# vcm 0.42fF
C1515 a_2346_10204# a_27974_10162# 0.35fF
C1516 a_23046_10162# col_n[20] 0.28fF
C1517 a_27974_2130# rowoff_n[0] 0.24fF
C1518 a_18026_5142# vcm 0.62fF
C1519 a_1962_1166# sample 0.14fF
C1520 a_6982_8154# row_n[6] 0.17fF
C1521 a_1962_14218# vcm 6.95fF
C1522 a_20034_3134# a_20034_2130# 1.00fF
C1523 a_2346_2172# a_3970_2130# 0.19fF
C1524 m2_18800_18014# m3_18932_18146# 2.78fF
C1525 a_1962_7190# a_22042_7150# 0.27fF
C1526 a_24050_17190# VDD 0.55fF
C1527 col[3] rowoff_n[14] 0.11fF
C1528 a_21038_12170# a_22042_12170# 0.97fF
C1529 a_31078_9158# vcm 0.62fF
C1530 a_14314_18234# vcm 0.22fF
C1531 a_34090_2130# VDD 0.59fF
C1532 a_2346_7192# col[11] 0.15fF
C1533 a_3970_10162# m2_4168_10410# 0.16fF
C1534 a_2346_4180# a_17022_4138# 0.19fF
C1535 a_9902_4138# a_9994_4138# 0.26fF
C1536 a_1962_4178# a_15318_4178# 0.14fF
C1537 a_5978_3134# col_n[3] 0.28fF
C1538 a_24962_18194# m2_24824_18014# 0.16fF
C1539 a_26058_11166# row_n[9] 0.17fF
C1540 a_24354_3174# vcm 0.22fF
C1541 a_1962_9198# col_n[27] 0.13fF
C1542 a_16018_10162# rowoff_n[8] 0.10fF
C1543 a_18026_13174# rowoff_n[11] 0.10fF
C1544 a_13918_5142# VDD 0.23fF
C1545 a_1962_3174# col[18] 0.11fF
C1546 a_2346_6188# a_30074_6146# 0.19fF
C1547 a_33086_7150# a_33086_6146# 1.00fF
C1548 a_1962_13214# m2_34864_12994# 0.17fF
C1549 a_1962_6186# a_28370_6186# 0.14fF
C1550 col_n[0] vcm 2.80fF
C1551 VDD col_n[3] 4.94fF
C1552 col[9] col[10] 0.20fF
C1553 ctop col[25] 1.98fF
C1554 a_1962_16226# col[20] 0.11fF
C1555 a_8990_16186# ctop 3.57fF
C1556 a_26058_8154# rowoff_n[6] 0.10fF
C1557 a_21038_13174# col[18] 0.29fF
C1558 m2_16792_946# a_1962_1166# 0.18fF
C1559 a_32082_17190# rowoff_n[15] 0.10fF
C1560 a_19030_1126# ctop 1.70fF
C1561 a_1962_1166# m2_33860_946# 0.10fF
C1562 a_2346_1168# m2_34864_946# 0.17fF
C1563 a_26970_9158# VDD 0.23fF
C1564 a_14010_9158# rowon_n[7] 0.14fF
C1565 a_5978_8154# a_5978_7150# 1.00fF
C1566 a_22954_8154# a_23046_8154# 0.26fF
C1567 a_1962_18234# a_17326_18234# 0.14fF
C1568 a_2346_17232# a_12914_17190# 0.35fF
C1569 a_6982_17190# a_7986_17190# 0.97fF
C1570 m2_19804_18014# m2_20808_18014# 0.96fF
C1571 a_1962_18234# col[30] 0.11fF
C1572 a_32082_5142# ctop 3.58fF
C1573 a_2346_3176# col[2] 0.15fF
C1574 m3_27968_18146# ctop 0.23fF
C1575 a_2346_16228# col[4] 0.15fF
C1576 a_34090_6146# m3_34996_6098# 0.13fF
C1577 a_3970_6146# col[1] 0.29fF
C1578 a_5978_12170# VDD 0.52fF
C1579 m2_24824_946# m2_25252_1374# 0.16fF
C1580 a_1962_5182# col_n[18] 0.13fF
C1581 a_1962_14218# a_6982_14178# 0.27fF
C1582 a_13006_4138# vcm 0.62fF
C1583 m2_1732_6970# m2_2160_7398# 0.16fF
C1584 a_21038_15182# col_n[18] 0.28fF
C1585 a_5886_14178# rowoff_n[12] 0.24fF
C1586 a_33086_12170# rowon_n[10] 0.14fF
C1587 a_17022_2130# a_18026_2130# 0.97fF
C1588 a_2346_2172# a_32994_2130# 0.35fF
C1589 a_22042_2130# col[19] 0.29fF
C1590 a_1962_12210# col[11] 0.11fF
C1591 a_19030_16186# VDD 0.52fF
C1592 a_19030_12170# a_19030_11166# 1.00fF
C1593 a_26058_8154# vcm 0.62fF
C1594 a_1962_16226# a_20034_16186# 0.27fF
C1595 a_10998_12170# row_n[10] 0.17fF
C1596 a_7986_2130# m2_8184_2378# 0.16fF
C1597 a_2346_11208# col[31] 0.15fF
C1598 a_9294_17230# vcm 0.22fF
C1599 a_26058_2130# row_n[0] 0.17fF
C1600 col[30] rowoff_n[13] 0.11fF
C1601 a_19334_2170# vcm 0.22fF
C1602 a_1962_13214# a_13310_13214# 0.14fF
C1603 a_2346_13216# a_15014_13174# 0.19fF
C1604 a_8898_13174# a_8990_13174# 0.26fF
C1605 a_3970_8154# col_n[1] 0.28fF
C1606 a_8898_4138# VDD 0.23fF
C1607 m3_34996_2082# VDD 0.27fF
C1608 a_32082_13174# m2_32280_13422# 0.16fF
C1609 a_30074_6146# a_31078_6146# 0.97fF
C1610 a_3970_15182# ctop 3.57fF
C1611 a_22042_4138# col_n[19] 0.28fF
C1612 a_1962_1166# col_n[9] 0.13fF
C1613 a_1962_14218# col_n[11] 0.13fF
C1614 a_30074_15182# row_n[13] 0.17fF
C1615 a_32082_16186# a_32082_15182# 1.00fF
C1616 a_2346_15224# a_28066_15182# 0.19fF
C1617 a_32386_6186# vcm 0.22fF
C1618 a_1962_15222# a_26362_15222# 0.14fF
C1619 m2_34864_10986# m2_34864_9982# 0.99fF
C1620 col[14] rowoff_n[14] 0.11fF
C1621 a_1962_8194# col[2] 0.11fF
C1622 a_21950_8154# VDD 0.23fF
C1623 a_2346_7192# a_4882_7150# 0.35fF
C1624 a_2966_15182# m2_3164_15430# 0.16fF
C1625 sample_n rowoff_n[10] 0.38fF
C1626 m2_14784_946# m3_13912_1078# 0.13fF
C1627 a_4974_17190# a_4974_16186# 1.00fF
C1628 a_21950_17190# a_22042_17190# 0.26fF
C1629 a_2346_7192# col[22] 0.15fF
C1630 a_8990_5142# rowoff_n[3] 0.10fF
C1631 a_27062_4138# ctop 3.58fF
C1632 a_18026_13174# rowon_n[11] 0.14fF
C1633 a_35002_12170# VDD 0.29fF
C1634 m2_25828_946# m3_25960_1078# 2.79fF
C1635 a_2346_9200# a_17934_9158# 0.35fF
C1636 a_7986_3134# vcm 0.62fF
C1637 a_1962_14218# a_34394_14218# 0.14fF
C1638 a_19030_3134# rowoff_n[1] 0.10fF
C1639 a_33086_3134# rowon_n[1] 0.14fF
C1640 a_34090_14178# rowoff_n[12] 0.10fF
C1641 a_1962_3174# col[29] 0.11fF
C1642 VDD col_n[14] 4.94fF
C1643 vcm col_n[10] 2.80fF
C1644 a_31990_2130# a_32082_2130# 0.26fF
C1645 a_1962_16226# col[31] 0.11fF
C1646 analog_in col[31] 0.10fF
C1647 a_29070_14178# m2_29268_14426# 0.16fF
C1648 a_1962_6186# a_12002_6146# 0.27fF
C1649 a_14010_15182# VDD 0.52fF
C1650 a_20034_7150# col[17] 0.29fF
C1651 a_16018_11166# a_17022_11166# 0.97fF
C1652 a_2346_11208# a_30986_11166# 0.35fF
C1653 a_1962_10202# col_n[2] 0.13fF
C1654 a_10998_3134# row_n[1] 0.17fF
C1655 a_21038_7150# vcm 0.62fF
C1656 a_4274_16226# vcm 0.22fF
C1657 a_2346_3176# a_6982_3134# 0.19fF
C1658 a_1962_3174# a_5278_3174# 0.14fF
C1659 a_4882_3134# a_4974_3134# 0.26fF
C1660 a_34090_17190# m2_34864_17010# 0.96fF
C1661 a_1962_8194# a_25054_8154# 0.27fF
C1662 a_14314_1166# vcm 0.23fF
C1663 a_7894_11166# rowoff_n[9] 0.24fF
C1664 a_2346_3176# col[13] 0.15fF
C1665 a_34090_11166# vcm 0.62fF
C1666 a_2346_16228# col[15] 0.15fF
C1667 a_15014_16186# row_n[14] 0.17fF
C1668 a_2346_4180# m2_1732_3958# 0.12fF
C1669 a_2346_5184# a_20034_5142# 0.19fF
C1670 a_28066_6146# a_28066_5142# 1.00fF
C1671 a_1962_5182# a_18330_5182# 0.14fF
C1672 a_30074_6146# row_n[4] 0.17fF
C1673 a_1962_5182# col_n[29] 0.13fF
C1674 a_17934_9158# rowoff_n[7] 0.24fF
C1675 a_27366_5182# vcm 0.22fF
C1676 a_29070_15182# a_30074_15182# 0.97fF
C1677 a_20034_9158# col_n[17] 0.28fF
C1678 a_21950_15182# rowoff_n[13] 0.24fF
C1679 a_1962_12210# col[22] 0.11fF
C1680 m2_31852_946# col[29] 0.39fF
C1681 m2_32856_18014# m3_33992_18146# 0.13fF
C1682 a_16930_7150# VDD 0.23fF
C1683 a_27974_7150# rowoff_n[5] 0.24fF
C1684 a_17934_7150# a_18026_7150# 0.26fF
C1685 a_1962_7190# a_31382_7190# 0.14fF
C1686 a_26058_15182# m2_26256_15430# 0.16fF
C1687 a_2346_7192# a_33086_7150# 0.19fF
C1688 a_28066_3134# m2_28264_3382# 0.16fF
C1689 a_18026_4138# rowon_n[2] 0.14fF
C1690 a_22042_3134# ctop 3.57fF
C1691 a_29982_11166# VDD 0.23fF
C1692 m3_26964_1078# m3_27968_1078# 0.22fF
C1693 m2_1732_12994# sample 0.19fF
C1694 m2_34864_6970# ctop 0.17fF
C1695 a_2346_12212# col[6] 0.15fF
C1696 a_2346_1168# a_22954_1126# 0.35fF
C1697 a_1962_1166# col_n[20] 0.13fF
C1698 a_22042_17190# rowon_n[15] 0.14fF
C1699 a_8990_14178# VDD 0.52fF
C1700 a_1962_14218# col_n[22] 0.13fF
C1701 a_14010_11166# a_14010_10162# 1.00fF
C1702 a_30986_11166# a_31078_11166# 0.26fF
C1703 m2_14784_946# a_14922_1126# 0.16fF
C1704 a_16018_6146# vcm 0.62fF
C1705 a_1962_15222# a_9994_15182# 0.27fF
C1706 a_18026_12170# col[15] 0.29fF
C1707 a_1962_8194# col[13] 0.11fF
C1708 a_8990_16186# rowoff_n[14] 0.10fF
C1709 col[25] rowoff_n[14] 0.11fF
C1710 a_3878_8154# VDD 0.23fF
C1711 a_23046_16186# m2_23244_16434# 0.16fF
C1712 a_2966_5142# col[0] 0.29fF
C1713 m2_19804_18014# vcm 0.28fF
C1714 a_2346_12212# a_4974_12170# 0.19fF
C1715 a_1962_12210# a_3270_12210# 0.14fF
C1716 a_15014_7150# row_n[5] 0.17fF
C1717 a_1962_17230# a_23046_17190# 0.27fF
C1718 a_29070_10162# vcm 0.62fF
C1719 a_25054_4138# m2_25252_4386# 0.16fF
C1720 m2_30848_18014# m2_31276_18442# 0.16fF
C1721 a_32082_3134# VDD 0.52fF
C1722 m3_3872_1078# ctop 0.35fF
C1723 a_1962_9198# row_n[7] 25.57fF
C1724 a_25054_5142# a_26058_5142# 0.97fF
C1725 a_34090_15182# m3_34996_15134# 0.13fF
C1726 a_27062_15182# a_27062_14178# 1.00fF
C1727 a_1962_14218# a_16322_14218# 0.14fF
C1728 a_2346_14220# a_18026_14178# 0.19fF
C1729 a_22346_4178# vcm 0.22fF
C1730 vcm col_n[21] 2.80fF
C1731 col_n[10] col_n[11] 0.10fF
C1732 VDD col_n[25] 4.95fF
C1733 col[9] rowoff_n[15] 0.11fF
C1734 col[20] col[21] 0.20fF
C1735 a_18026_14178# col_n[15] 0.28fF
C1736 a_11910_6146# VDD 0.23fF
C1737 a_1962_10202# col_n[13] 0.13fF
C1738 a_34090_10162# row_n[8] 0.17fF
C1739 a_6982_17190# ctop 3.39fF
C1740 a_19030_1126# col[16] 0.38fF
C1741 a_2966_7150# vcm 0.61fF
C1742 a_1962_16226# a_29374_16226# 0.14fF
C1743 a_2346_16228# a_31078_16186# 0.19fF
C1744 a_16930_16186# a_17022_16186# 0.26fF
C1745 a_1962_4178# col[4] 0.11fF
C1746 a_17022_2130# ctop 3.39fF
C1747 a_1962_17230# col[6] 0.11fF
C1748 m2_10768_18014# VDD 1.27fF
C1749 a_1962_18234# m2_25828_18014# 0.18fF
C1750 a_24962_10162# VDD 0.23fF
C1751 a_2346_8196# a_7894_8154# 0.35fF
C1752 a_20034_17190# m2_20232_17438# 0.16fF
C1753 a_2346_3176# col[24] 0.15fF
C1754 a_2346_16228# col[26] 0.15fF
C1755 a_10906_4138# rowoff_n[2] 0.24fF
C1756 a_23958_12170# rowoff_n[10] 0.24fF
C1757 a_22042_5142# m2_22240_5390# 0.16fF
C1758 a_22042_8154# rowon_n[6] 0.14fF
C1759 a_30074_6146# ctop 3.58fF
C1760 a_3970_13174# VDD 0.52fF
C1761 a_2346_18236# m2_20808_18014# 0.19fF
C1762 a_2346_10204# a_20946_10162# 0.35fF
C1763 a_10998_10162# a_12002_10162# 0.97fF
C1764 a_20946_2130# rowoff_n[0] 0.24fF
C1765 a_10998_5142# vcm 0.62fF
C1766 a_19030_3134# col_n[16] 0.28fF
C1767 a_3878_15182# rowoff_n[13] 0.24fF
C1768 m2_9764_18014# m3_8892_18146# 0.13fF
C1769 a_16018_17190# col[13] 0.29fF
C1770 a_1962_6186# col_n[4] 0.13fF
C1771 a_1962_7190# a_15014_7150# 0.27fF
C1772 a_17022_17190# VDD 0.55fF
C1773 a_2346_12212# a_33998_12170# 0.35fF
C1774 a_24050_9158# vcm 0.62fF
C1775 a_34090_13174# col[31] 0.29fF
C1776 a_7286_18234# vcm 0.22fF
C1777 a_27062_2130# VDD 0.55fF
C1778 a_1962_4178# a_8290_4178# 0.14fF
C1779 a_23046_5142# a_23046_4138# 1.00fF
C1780 a_2346_4180# a_9994_4138# 0.19fF
C1781 m3_1864_6098# m3_1864_5094# 0.22fF
C1782 a_1962_9198# a_28066_9158# 0.27fF
C1783 a_2346_12212# col[17] 0.15fF
C1784 a_19030_11166# row_n[9] 0.17fF
C1785 a_17326_3174# vcm 0.22fF
C1786 a_24050_14178# a_25054_14178# 0.97fF
C1787 a_8990_10162# rowoff_n[8] 0.10fF
C1788 a_10998_13174# rowoff_n[11] 0.10fF
C1789 a_19030_6146# m2_19228_6394# 0.16fF
C1790 a_6890_5142# VDD 0.23fF
C1791 a_1962_6186# a_21342_6186# 0.14fF
C1792 a_2346_6188# a_23046_6146# 0.19fF
C1793 a_12914_6146# a_13006_6146# 0.26fF
C1794 a_19030_8154# rowoff_n[6] 0.10fF
C1795 a_15014_17190# m3_14916_18146# 0.15fF
C1796 a_1962_8194# col[24] 0.11fF
C1797 a_30378_7190# vcm 0.22fF
C1798 a_17022_6146# col[14] 0.29fF
C1799 a_1962_1166# m2_9764_946# 0.18fF
C1800 a_25054_17190# rowoff_n[15] 0.10fF
C1801 a_29070_6146# rowoff_n[4] 0.10fF
C1802 a_19942_9158# VDD 0.23fF
C1803 a_6982_9158# rowon_n[7] 0.14fF
C1804 a_2346_8196# a_2346_7192# 0.22fF
C1805 a_1962_8194# a_35398_8194# 0.14fF
C1806 a_34090_15182# col_n[31] 0.28fF
C1807 a_1962_18234# a_10298_18234# 0.14fF
C1808 m2_7756_946# m2_8184_1374# 0.16fF
C1809 a_2346_17232# a_5886_17190# 0.35fF
C1810 m2_12776_18014# m2_13780_18014# 0.96fF
C1811 a_25054_5142# ctop 3.58fF
C1812 a_32994_13174# VDD 0.23fF
C1813 a_8990_10162# a_8990_9158# 1.00fF
C1814 a_25966_10162# a_26058_10162# 0.26fF
C1815 col_n[0] row_n[15] 0.23fF
C1816 vcm rowon_n[15] 0.50fF
C1817 VDD rowon_n[13] 2.61fF
C1818 col[20] rowoff_n[15] 0.11fF
C1819 a_2346_8196# col[8] 0.15fF
C1820 a_5978_4138# vcm 0.62fF
C1821 a_26058_12170# rowon_n[10] 0.14fF
C1822 a_1962_10202# col_n[24] 0.13fF
C1823 a_2346_2172# a_25966_2130# 0.35fF
C1824 a_16018_7150# m2_16216_7398# 0.16fF
C1825 m2_34864_17010# m3_34996_17142# 2.76fF
C1826 a_17022_8154# col_n[14] 0.28fF
C1827 a_35002_15182# m2_34864_15002# 0.16fF
C1828 a_12002_16186# VDD 0.52fF
C1829 a_1962_4178# col[15] 0.11fF
C1830 a_1962_17230# col[17] 0.11fF
C1831 a_1962_16226# a_13006_16186# 0.27fF
C1832 a_19030_8154# vcm 0.62fF
C1833 a_3970_12170# row_n[10] 0.17fF
C1834 a_2346_2172# m2_2736_1950# 0.20fF
C1835 m2_12776_18014# col[10] 0.28fF
C1836 a_20034_4138# a_21038_4138# 0.97fF
C1837 a_19030_2130# row_n[0] 0.17fF
C1838 a_1962_13214# a_6282_13214# 0.14fF
C1839 a_12306_2170# vcm 0.22fF
C1840 a_22042_14178# a_22042_13174# 1.00fF
C1841 a_2346_13216# a_7986_13174# 0.19fF
C1842 a_32082_12170# vcm 0.62fF
C1843 m3_1864_15134# VDD 0.25fF
C1844 a_2346_10204# a_1962_10202# 2.62fF
C1845 a_2346_17232# col[1] 0.15fF
C1846 a_23046_15182# row_n[13] 0.17fF
C1847 a_25358_6186# vcm 0.22fF
C1848 a_1962_15222# a_19334_15222# 0.14fF
C1849 a_11910_15182# a_12002_15182# 0.26fF
C1850 a_2346_15224# a_21038_15182# 0.19fF
C1851 a_1962_6186# col_n[15] 0.13fF
C1852 m2_34864_12994# VDD 1.01fF
C1853 a_13006_8154# m2_13204_8402# 0.16fF
C1854 a_15014_11166# col[12] 0.29fF
C1855 a_14922_8154# VDD 0.23fF
C1856 a_33086_8154# a_34090_8154# 0.97fF
C1857 m2_28840_18014# col_n[26] 0.25fF
C1858 a_1962_13214# col[8] 0.11fF
C1859 a_2346_17232# a_34090_17190# 0.19fF
C1860 a_1962_17230# a_32386_17230# 0.14fF
C1861 a_33086_7150# col[30] 0.29fF
C1862 m2_9764_946# m3_9896_1078# 2.79fF
C1863 a_20034_4138# ctop 3.58fF
C1864 a_10998_13174# rowon_n[11] 0.14fF
C1865 a_2346_12212# col[28] 0.15fF
C1866 a_27974_12170# VDD 0.23fF
C1867 m3_22948_18146# m3_23952_18146# 0.22fF
C1868 a_5978_9158# a_6982_9158# 0.97fF
C1869 a_2346_9200# a_10906_9158# 0.35fF
C1870 a_26058_3134# rowon_n[1] 0.14fF
C1871 a_12002_3134# rowoff_n[1] 0.10fF
C1872 a_27062_14178# rowoff_n[12] 0.10fF
C1873 m2_1732_9982# ctop 0.17fF
C1874 a_33086_8154# ctop 3.57fF
C1875 m2_34864_13998# m3_34996_14130# 2.76fF
C1876 a_1962_6186# a_4974_6146# 0.27fF
C1877 a_3878_6146# a_3970_6146# 0.26fF
C1878 a_6982_15182# VDD 0.52fF
C1879 a_2346_11208# a_23958_11166# 0.35fF
C1880 a_15014_13174# col_n[12] 0.28fF
C1881 a_3970_3134# row_n[1] 0.17fF
C1882 a_14010_7150# vcm 0.62fF
C1883 m2_22816_946# m2_23820_946# 0.96fF
C1884 a_1962_2170# col_n[6] 0.13fF
C1885 a_1962_15222# col_n[8] 0.13fF
C1886 a_30074_16186# rowon_n[14] 0.14fF
C1887 a_18026_4138# a_18026_3134# 1.00fF
C1888 a_9994_9158# m2_10192_9406# 0.16fF
C1889 a_35494_10524# VDD 0.11fF
C1890 a_33086_9158# col_n[30] 0.28fF
C1891 a_1962_8194# a_18026_8154# 0.27fF
C1892 a_7286_1166# vcm 0.23fF
C1893 a_19030_13174# a_20034_13174# 0.97fF
C1894 a_1962_13214# a_1962_12210# 0.16fF
C1895 a_27062_11166# vcm 0.62fF
C1896 a_7986_16186# row_n[14] 0.17fF
C1897 a_2346_18236# vcm 0.24fF
C1898 a_30074_4138# VDD 0.52fF
C1899 col_n[4] row_n[12] 0.23fF
C1900 col_n[10] row_n[15] 0.23fF
C1901 vcm row_n[10] 0.49fF
C1902 VDD row_n[8] 2.93fF
C1903 a_1962_5182# a_11302_5182# 0.14fF
C1904 col_n[2] row_n[11] 0.23fF
C1905 col_n[6] row_n[13] 0.23fF
C1906 col_n[21] col_n[22] 0.10fF
C1907 col_n[8] row_n[14] 0.23fF
C1908 a_7894_5142# a_7986_5142# 0.26fF
C1909 a_2346_5184# a_13006_5142# 0.19fF
C1910 sample row_n[9] 1.03fF
C1911 col[31] rowoff_n[15] 0.11fF
C1912 a_2346_8196# col[19] 0.15fF
C1913 a_23046_6146# row_n[4] 0.17fF
C1914 a_1962_10202# a_31078_10162# 0.27fF
C1915 a_10906_9158# rowoff_n[7] 0.24fF
C1916 a_20338_5182# vcm 0.22fF
C1917 a_14922_15182# rowoff_n[13] 0.24fF
C1918 a_16018_2130# col_n[13] 0.28fF
C1919 m2_23820_18014# m3_23952_18146# 2.79fF
C1920 a_9902_7150# VDD 0.23fF
C1921 a_20946_7150# rowoff_n[5] 0.24fF
C1922 a_31078_8154# a_31078_7150# 1.00fF
C1923 a_2346_7192# a_26058_7150# 0.19fF
C1924 a_1962_7190# a_24354_7190# 0.14fF
C1925 a_1962_4178# col[26] 0.11fF
C1926 a_1962_17230# col[28] 0.11fF
C1927 a_13006_16186# col[10] 0.29fF
C1928 a_33390_9198# vcm 0.22fF
C1929 a_32082_17190# a_33086_17190# 0.97fF
C1930 a_10998_4138# rowon_n[2] 0.14fF
C1931 a_30986_5142# rowoff_n[3] 0.24fF
C1932 a_1962_11206# col_n[0] 0.13fF
C1933 a_15014_3134# ctop 3.57fF
C1934 a_6982_10162# m2_7180_10410# 0.16fF
C1935 a_22954_11166# VDD 0.23fF
C1936 a_31078_12170# col[28] 0.29fF
C1937 m3_12908_1078# m3_13912_1078# 0.22fF
C1938 a_20946_9158# a_21038_9158# 0.26fF
C1939 a_3970_9158# a_3970_8154# 1.00fF
C1940 a_2346_1168# a_15926_1126# 0.35fF
C1941 m2_34864_10986# m3_34996_11118# 2.76fF
C1942 a_28066_7150# ctop 3.58fF
C1943 a_2346_4180# col[10] 0.15fF
C1944 a_15014_17190# rowon_n[15] 0.14fF
C1945 a_2346_17232# col[12] 0.15fF
C1946 a_1962_6186# col_n[26] 0.13fF
C1947 a_2346_15224# a_2966_15182# 0.21fF
C1948 a_8990_6146# vcm 0.62fF
C1949 a_30074_7150# rowon_n[5] 0.14fF
C1950 a_2346_3176# a_28978_3134# 0.35fF
C1951 a_14010_5142# col[11] 0.29fF
C1952 a_15014_3134# a_16018_3134# 0.97fF
C1953 a_1962_13214# col[19] 0.11fF
C1954 a_33998_13174# a_34090_13174# 0.26fF
C1955 a_17022_13174# a_17022_12170# 1.00fF
C1956 m2_5748_18014# vcm 0.28fF
C1957 a_7986_7150# row_n[5] 0.17fF
C1958 a_31078_14178# col_n[28] 0.28fF
C1959 a_22042_10162# vcm 0.62fF
C1960 a_29070_11166# rowoff_n[9] 0.10fF
C1961 a_1962_17230# a_16018_17190# 0.27fF
C1962 m2_23820_18014# m2_24248_18442# 0.16fF
C1963 a_25054_3134# VDD 0.52fF
C1964 m3_34996_14130# ctop 0.23fF
C1965 a_3970_11166# m2_4168_11414# 0.16fF
C1966 a_15318_4178# vcm 0.22fF
C1967 a_1962_14218# a_9294_14218# 0.14fF
C1968 a_2346_14220# a_10998_14178# 0.19fF
C1969 a_6890_14178# a_6982_14178# 0.26fF
C1970 a_35094_14178# vcm 0.12fF
C1971 m2_1732_15002# m3_1864_14130# 0.15fF
C1972 a_4882_6146# VDD 0.23fF
C1973 a_2346_13216# col[3] 0.15fF
C1974 a_28066_7150# a_29070_7150# 0.97fF
C1975 a_1962_14218# m2_34864_13998# 0.17fF
C1976 a_27062_10162# row_n[8] 0.17fF
C1977 a_14010_7150# col_n[11] 0.28fF
C1978 m2_15788_946# col_n[13] 0.37fF
C1979 a_1962_2170# col_n[17] 0.13fF
C1980 a_28370_8194# vcm 0.22fF
C1981 a_1962_16226# a_22346_16226# 0.14fF
C1982 a_1962_15222# col_n[19] 0.13fF
C1983 a_2346_16228# a_24050_16186# 0.19fF
C1984 a_30074_17190# a_30074_16186# 1.00fF
C1985 a_10998_2130# m2_11196_2378# 0.16fF
C1986 m2_1732_13998# m2_1732_12994# 0.99fF
C1987 a_9994_2130# ctop 3.39fF
C1988 a_1962_18234# m2_11772_18014# 0.18fF
C1989 a_32082_3134# col_n[29] 0.28fF
C1990 a_17934_10162# VDD 0.23fF
C1991 a_1962_9198# col[10] 0.11fF
C1992 a_2346_14220# row_n[12] 0.35fF
C1993 a_29070_17190# col[26] 0.29fF
C1994 a_16930_12170# rowoff_n[10] 0.24fF
C1995 col_n[1] row_n[5] 0.23fF
C1996 col_n[0] row_n[4] 0.23fF
C1997 col_n[3] row_n[6] 0.23fF
C1998 col_n[13] row_n[11] 0.23fF
C1999 col_n[7] row_n[8] 0.23fF
C2000 VDD rowon_n[2] 2.61fF
C2001 col_n[19] row_n[14] 0.23fF
C2002 col_n[5] row_n[7] 0.23fF
C2003 col_n[21] row_n[15] 0.23fF
C2004 col_n[9] row_n[9] 0.23fF
C2005 vcm rowon_n[4] 0.50fF
C2006 col_n[15] row_n[12] 0.23fF
C2007 col_n[17] row_n[13] 0.23fF
C2008 col_n[11] row_n[10] 0.23fF
C2009 a_2346_8196# col[30] 0.15fF
C2010 a_15014_8154# rowon_n[6] 0.14fF
C2011 m2_34864_7974# m3_34996_8106# 2.76fF
C2012 a_23046_6146# ctop 3.58fF
C2013 m3_15920_1078# VDD 0.14fF
C2014 a_2346_18236# m2_6752_18014# 0.19fF
C2015 a_30986_14178# VDD 0.23fF
C2016 m2_34864_2954# vcm 0.50fF
C2017 a_2346_10204# a_13918_10162# 0.35fF
C2018 a_1962_10202# rowon_n[8] 1.18fF
C2019 a_13918_2130# rowoff_n[0] 0.24fF
C2020 a_3970_5142# vcm 0.62fF
C2021 m2_33860_18014# ctop 0.18fF
C2022 a_30986_16186# rowoff_n[14] 0.24fF
C2023 a_13006_3134# a_13006_2130# 1.00fF
C2024 a_29982_3134# a_30074_3134# 0.26fF
C2025 a_2346_9200# ctop 1.59fF
C2026 a_1962_7190# a_7986_7150# 0.27fF
C2027 m2_34864_10986# row_n[9] 0.15fF
C2028 a_12002_10162# col[9] 0.29fF
C2029 a_9994_17190# VDD 0.55fF
C2030 a_14010_12170# a_15014_12170# 0.97fF
C2031 a_2346_12212# a_26970_12170# 0.35fF
C2032 m2_20808_946# m3_19936_1078# 0.12fF
C2033 a_1962_11206# col_n[10] 0.13fF
C2034 a_34090_11166# rowon_n[9] 0.14fF
C2035 a_17022_9158# vcm 0.62fF
C2036 a_20034_2130# VDD 0.54fF
C2037 a_2346_4180# a_2874_4138# 0.35fF
C2038 a_1962_5182# col[1] 0.11fF
C2039 a_30074_6146# col[27] 0.29fF
C2040 m2_30848_946# m3_30980_1078# 2.79fF
C2041 m3_1864_13126# m3_1864_12122# 0.22fF
C2042 a_1962_9198# a_21038_9158# 0.27fF
C2043 a_10298_3174# vcm 0.22fF
C2044 a_12002_11166# row_n[9] 0.17fF
C2045 a_30074_13174# vcm 0.62fF
C2046 a_3970_13174# rowoff_n[11] 0.10fF
C2047 a_2346_4180# col[21] 0.15fF
C2048 a_2346_17232# col[23] 0.15fF
C2049 m2_1732_11990# m3_1864_11118# 0.15fF
C2050 a_33086_6146# VDD 0.52fF
C2051 a_1962_6186# a_14314_6186# 0.14fF
C2052 a_2346_6188# a_16018_6146# 0.19fF
C2053 a_32082_14178# m2_32280_14426# 0.16fF
C2054 a_26058_7150# a_26058_6146# 1.00fF
C2055 a_12002_8154# rowoff_n[6] 0.10fF
C2056 a_1962_11206# a_34090_11166# 0.27fF
C2057 m2_20808_946# a_21038_2130# 0.99fF
C2058 a_23350_7190# vcm 0.22fF
C2059 a_27062_16186# a_28066_16186# 0.97fF
C2060 a_12002_12170# col_n[9] 0.28fF
C2061 m2_1732_4962# sample_n 0.15fF
C2062 a_18026_17190# rowoff_n[15] 0.10fF
C2063 m2_1732_16006# VDD 1.02fF
C2064 a_1962_13214# col[30] 0.11fF
C2065 a_2346_5184# row_n[3] 0.35fF
C2066 a_22042_6146# rowoff_n[4] 0.10fF
C2067 a_3970_2130# m3_3872_1078# 0.12fF
C2068 a_12914_9158# VDD 0.23fF
C2069 ctop rowoff_n[7] 0.60fF
C2070 rowon_n[1] rowoff_n[1] 20.27fF
C2071 a_15926_8154# a_16018_8154# 0.26fF
C2072 a_1962_8194# a_27366_8194# 0.14fF
C2073 a_2346_8196# a_29070_8154# 0.19fF
C2074 a_2966_16186# m2_3164_16434# 0.16fF
C2075 a_31078_14178# row_n[12] 0.17fF
C2076 a_1962_18234# a_3270_18234# 0.14fF
C2077 a_30074_8154# col_n[27] 0.28fF
C2078 a_1962_7190# col_n[1] 0.13fF
C2079 a_32082_4138# rowoff_n[2] 0.10fF
C2080 m2_10768_946# ctop 0.18fF
C2081 m2_5748_18014# m2_6752_18014# 0.96fF
C2082 m2_34864_4962# m3_34996_5094# 2.76fF
C2083 a_18026_5142# ctop 3.58fF
C2084 a_1962_14218# ctop 1.49fF
C2085 a_25966_13174# VDD 0.23fF
C2086 a_2346_13216# col[14] 0.15fF
C2087 a_19030_12170# rowon_n[10] 0.14fF
C2088 a_9994_2130# a_10998_2130# 0.97fF
C2089 a_2346_2172# a_18938_2130# 0.35fF
C2090 a_31078_9158# ctop 3.58fF
C2091 a_29070_15182# m2_29268_15430# 0.16fF
C2092 a_1962_2170# col_n[28] 0.13fF
C2093 a_4974_16186# VDD 0.52fF
C2094 a_34090_2130# rowon_n[0] 0.14fF
C2095 a_1962_15222# col_n[30] 0.13fF
C2096 a_28978_12170# a_29070_12170# 0.26fF
C2097 a_12002_12170# a_12002_11166# 1.00fF
C2098 a_12002_8154# vcm 0.62fF
C2099 a_1962_16226# a_5978_16186# 0.27fF
C2100 a_9994_15182# col[7] 0.29fF
C2101 a_31078_3134# m2_31276_3382# 0.16fF
C2102 a_1962_9198# col[21] 0.11fF
C2103 a_2346_4180# a_31990_4138# 0.35fF
C2104 a_12002_2130# row_n[0] 0.17fF
C2105 a_12002_17190# m2_11772_18014# 1.00fF
C2106 a_28066_11166# col[25] 0.29fF
C2107 a_5278_2170# vcm 0.22fF
C2108 col_n[8] row_n[3] 0.23fF
C2109 col_n[2] row_n[0] 0.23fF
C2110 rowon_n[15] row_n[15] 19.75fF
C2111 col_n[4] row_n[1] 0.23fF
C2112 col_n[10] row_n[4] 0.23fF
C2113 col_n[14] row_n[6] 0.23fF
C2114 col_n[26] row_n[12] 0.23fF
C2115 col_n[28] row_n[13] 0.23fF
C2116 col_n[12] row_n[5] 0.23fF
C2117 col_n[0] ctop 1.81fF
C2118 col_n[30] row_n[14] 0.23fF
C2119 col_n[16] row_n[7] 0.23fF
C2120 col_n[6] row_n[2] 0.23fF
C2121 col_n[24] row_n[11] 0.23fF
C2122 col_n[18] row_n[8] 0.23fF
C2123 VDD en_bit_n[2] 0.15fF
C2124 col_n[22] row_n[10] 0.23fF
C2125 col_n[20] row_n[9] 0.23fF
C2126 a_30986_10162# rowoff_n[8] 0.24fF
C2127 a_32994_13174# rowoff_n[11] 0.24fF
C2128 a_25054_12170# vcm 0.62fF
C2129 a_2346_5184# m2_1732_4962# 0.12fF
C2130 m2_1732_8978# m3_1864_8106# 0.15fF
C2131 a_28066_5142# VDD 0.52fF
C2132 m3_11904_18146# VDD 0.30fF
C2133 a_23046_6146# a_24050_6146# 0.97fF
C2134 a_16018_15182# row_n[13] 0.17fF
C2135 a_18330_6186# vcm 0.22fF
C2136 a_1962_15222# a_12306_15222# 0.14fF
C2137 a_2346_15224# a_14010_15182# 0.19fF
C2138 a_25054_16186# a_25054_15182# 1.00fF
C2139 a_2346_9200# col[5] 0.15fF
C2140 a_31078_5142# row_n[3] 0.17fF
C2141 a_9994_17190# col_n[7] 0.28fF
C2142 a_7894_8154# VDD 0.23fF
C2143 a_1962_18234# col_n[4] 0.13fF
C2144 a_26058_16186# m2_26256_16434# 0.16fF
C2145 a_1962_11206# col_n[21] 0.13fF
C2146 a_10998_4138# col[8] 0.29fF
C2147 a_31382_10202# vcm 0.22fF
C2148 m2_25828_946# col[23] 0.39fF
C2149 a_1962_17230# a_25358_17230# 0.14fF
C2150 a_14922_17190# a_15014_17190# 0.26fF
C2151 a_2346_17232# a_27062_17190# 0.19fF
C2152 a_28066_4138# m2_28264_4386# 0.16fF
C2153 a_28066_13174# col_n[25] 0.28fF
C2154 a_1962_5182# col[12] 0.11fF
C2155 a_13006_4138# ctop 3.58fF
C2156 m3_18932_1078# ctop 0.31fF
C2157 a_3970_13174# rowon_n[11] 0.14fF
C2158 a_20946_12170# VDD 0.23fF
C2159 m3_8892_18146# m3_9896_18146# 0.22fF
C2160 a_1962_9198# a_2966_9158# 0.27fF
C2161 a_19030_3134# rowon_n[1] 0.14fF
C2162 a_4974_3134# rowoff_n[1] 0.10fF
C2163 a_20034_14178# rowoff_n[12] 0.10fF
C2164 a_24962_2130# a_25054_2130# 0.26fF
C2165 a_26058_8154# ctop 3.58fF
C2166 a_33998_16186# VDD 0.23fF
C2167 a_2346_11208# a_16930_11166# 0.35fF
C2168 a_8990_11166# a_9994_11166# 0.97fF
C2169 a_6982_7150# vcm 0.62fF
C2170 a_10998_6146# col_n[8] 0.28fF
C2171 a_10998_2130# m2_10768_946# 0.99fF
C2172 col[7] rowoff_n[9] 0.11fF
C2173 col[4] rowoff_n[6] 0.11fF
C2174 col[3] rowoff_n[5] 0.11fF
C2175 col[2] rowoff_n[4] 0.11fF
C2176 col[1] rowoff_n[3] 0.11fF
C2177 col[0] rowoff_n[2] 0.11fF
C2178 col[6] rowoff_n[8] 0.11fF
C2179 col[5] rowoff_n[7] 0.11fF
C2180 a_23046_16186# rowon_n[14] 0.14fF
C2181 a_1962_7190# col_n[12] 0.13fF
C2182 a_23046_17190# m2_23244_17438# 0.16fF
C2183 a_1962_8194# a_10998_8154# 0.27fF
C2184 a_31078_17190# m2_30848_18014# 1.00fF
C2185 a_2346_13216# a_29982_13174# 0.35fF
C2186 a_29070_2130# col_n[26] 0.29fF
C2187 a_2966_4138# col_n[0] 0.28fF
C2188 a_20034_11166# vcm 0.62fF
C2189 a_1962_1166# col[3] 0.11fF
C2190 a_26058_16186# col[23] 0.29fF
C2191 a_25054_5142# m2_25252_5390# 0.16fF
C2192 a_1962_14218# col[5] 0.11fF
C2193 m2_1732_5966# m3_1864_5094# 0.15fF
C2194 a_23046_4138# VDD 0.52fF
C2195 a_2346_5184# a_5978_5142# 0.19fF
C2196 a_1962_5182# a_4274_5182# 0.14fF
C2197 a_21038_6146# a_21038_5142# 1.00fF
C2198 a_16018_6146# row_n[4] 0.17fF
C2199 a_1962_10202# a_24050_10162# 0.27fF
C2200 a_2346_13216# col[25] 0.15fF
C2201 a_13310_5182# vcm 0.22fF
C2202 a_22042_15182# a_23046_15182# 0.97fF
C2203 a_33086_15182# vcm 0.62fF
C2204 a_7894_15182# rowoff_n[13] 0.24fF
C2205 m2_14784_18014# m3_13912_18146# 0.13fF
C2206 a_2346_7192# VDD 32.63fF
C2207 a_13918_7150# rowoff_n[5] 0.24fF
C2208 a_1962_7190# a_17326_7190# 0.14fF
C2209 a_10906_7150# a_10998_7150# 0.26fF
C2210 a_2346_7192# a_19030_7150# 0.19fF
C2211 a_8990_9158# col[6] 0.29fF
C2212 a_26362_9198# vcm 0.22fF
C2213 a_23958_5142# rowoff_n[3] 0.24fF
C2214 a_3970_4138# rowon_n[2] 0.14fF
C2215 a_7986_3134# ctop 3.57fF
C2216 a_1962_3174# col_n[3] 0.13fF
C2217 a_15926_11166# VDD 0.23fF
C2218 m3_1864_2082# m3_2868_2082# 0.22fF
C2219 m3_34996_3086# m3_34996_2082# 0.22fF
C2220 col_n[23] row_n[5] 0.23fF
C2221 col_n[25] row_n[6] 0.23fF
C2222 col_n[17] row_n[2] 0.23fF
C2223 col_n[10] ctop 2.02fF
C2224 col_n[31] row_n[9] 0.23fF
C2225 col_n[21] row_n[4] 0.23fF
C2226 col_n[29] row_n[8] 0.23fF
C2227 col_n[2] col[2] 0.72fF
C2228 col_n[19] row_n[3] 0.23fF
C2229 col_n[27] row_n[7] 0.23fF
C2230 VDD col[8] 4.17fF
C2231 vcm col[4] 5.84fF
C2232 col_n[13] row_n[0] 0.23fF
C2233 col_n[15] row_n[1] 0.23fF
C2234 a_1962_9198# a_30378_9198# 0.14fF
C2235 a_2346_9200# a_32082_9158# 0.19fF
C2236 a_1962_16226# col_n[5] 0.13fF
C2237 a_34090_10162# a_34090_9158# 1.00fF
C2238 a_27062_5142# col[24] 0.29fF
C2239 a_33998_3134# rowoff_n[1] 0.24fF
C2240 a_18026_1126# en_bit_n[1] 0.25fF
C2241 a_22042_6146# m2_22240_6394# 0.16fF
C2242 a_2346_1168# a_8898_1126# 0.35fF
C2243 a_21038_7150# ctop 3.58fF
C2244 a_7986_17190# rowon_n[15] 0.14fF
C2245 a_28978_15182# VDD 0.23fF
C2246 a_6982_11166# a_6982_10162# 1.00fF
C2247 a_23958_11166# a_24050_11166# 0.26fF
C2248 m2_1732_5966# vcm 0.45fF
C2249 a_18026_17190# m3_17928_18146# 0.15fF
C2250 a_2346_9200# col[16] 0.15fF
C2251 a_34394_7190# vcm 0.22fF
C2252 a_23046_7150# rowon_n[5] 0.14fF
C2253 a_7894_1126# m2_7756_946# 0.16fF
C2254 a_1962_18234# col_n[15] 0.13fF
C2255 a_2346_3176# a_21950_3134# 0.35fF
C2256 a_8990_11166# col_n[6] 0.28fF
C2257 a_2346_1168# m2_27836_946# 0.19fF
C2258 a_34090_11166# ctop 3.42fF
C2259 a_1962_5182# col[23] 0.11fF
C2260 a_1962_17230# a_8990_17190# 0.27fF
C2261 a_22042_11166# rowoff_n[9] 0.10fF
C2262 a_15014_10162# vcm 0.62fF
C2263 a_27062_7150# col_n[24] 0.28fF
C2264 m2_16792_18014# m2_17220_18442# 0.16fF
C2265 m2_1732_2954# m3_1864_2082# 0.15fF
C2266 a_18026_3134# VDD 0.52fF
C2267 m3_14916_18146# ctop 0.23fF
C2268 a_18026_5142# a_19030_5142# 0.97fF
C2269 a_2346_5184# a_35002_5142# 0.35fF
C2270 a_1962_12210# VDD 2.73fF
C2271 a_32082_9158# rowoff_n[7] 0.10fF
C2272 a_20034_15182# a_20034_14178# 1.00fF
C2273 a_2346_14220# a_3970_14178# 0.19fF
C2274 a_8290_4178# vcm 0.22fF
C2275 m2_34864_12994# rowon_n[11] 0.13fF
C2276 a_28066_14178# vcm 0.62fF
C2277 a_1962_2170# a_29070_2130# 0.27fF
C2278 a_19030_7150# m2_19228_7398# 0.16fF
C2279 a_31078_7150# VDD 0.52fF
C2280 a_20034_10162# row_n[8] 0.17fF
C2281 m2_1732_13998# rowoff_n[12] 0.12fF
C2282 a_2346_5184# col[7] 0.15fF
C2283 col[12] rowoff_n[3] 0.11fF
C2284 col[11] rowoff_n[2] 0.11fF
C2285 col[14] rowoff_n[5] 0.11fF
C2286 col[13] rowoff_n[4] 0.11fF
C2287 col[15] rowoff_n[6] 0.11fF
C2288 col[9] rowoff_n[0] 0.11fF
C2289 col[10] rowoff_n[1] 0.11fF
C2290 a_21342_8194# vcm 0.22fF
C2291 col[17] rowoff_n[8] 0.11fF
C2292 col[18] rowoff_n[9] 0.11fF
C2293 col[16] rowoff_n[7] 0.11fF
C2294 a_2346_16228# a_17022_16186# 0.19fF
C2295 a_9902_16186# a_9994_16186# 0.26fF
C2296 a_1962_16226# a_15318_16226# 0.14fF
C2297 a_1962_7190# col_n[23] 0.13fF
C2298 a_6982_14178# col[4] 0.29fF
C2299 a_10906_10162# VDD 0.23fF
C2300 a_31078_9158# a_32082_9158# 0.97fF
C2301 a_1962_1166# col[14] 0.11fF
C2302 a_1962_14218# col[16] 0.11fF
C2303 a_35398_12210# vcm 0.23fF
C2304 a_9902_12170# rowoff_n[10] 0.24fF
C2305 a_25054_10162# col[22] 0.29fF
C2306 a_19942_1126# a_20034_1126# 0.26fF
C2307 a_7986_8154# rowon_n[6] 0.14fF
C2308 a_16018_6146# ctop 3.58fF
C2309 m3_34996_8106# VDD 0.26fF
C2310 a_23958_14178# VDD 0.23fF
C2311 a_2346_10204# a_6890_10162# 0.35fF
C2312 a_3970_10162# a_4974_10162# 0.97fF
C2313 a_6890_2130# rowoff_n[0] 0.24fF
C2314 col[2] rowoff_n[10] 0.11fF
C2315 a_23958_16186# rowoff_n[14] 0.24fF
C2316 m2_19804_18014# ctop 0.18fF
C2317 a_16018_8154# m2_16216_8402# 0.16fF
C2318 a_29070_10162# ctop 3.58fF
C2319 m2_1732_15002# row_n[13] 0.13fF
C2320 a_35002_16186# m2_34864_16006# 0.16fF
C2321 a_2874_17190# VDD 0.24fF
C2322 a_6982_16186# col_n[4] 0.28fF
C2323 a_2346_12212# a_19942_12170# 0.35fF
C2324 a_2346_14220# col[0] 0.15fF
C2325 a_7986_3134# col[5] 0.29fF
C2326 a_27062_11166# rowon_n[9] 0.14fF
C2327 a_9994_9158# vcm 0.62fF
C2328 a_1962_3174# col_n[14] 0.13fF
C2329 a_13006_2130# VDD 0.55fF
C2330 col_n[7] col[8] 5.98fF
C2331 vcm col[15] 5.84fF
C2332 a_1962_16226# col_n[16] 0.13fF
C2333 col_n[17] en_bit_n[0] 0.17fF
C2334 col_n[26] row_n[1] 0.23fF
C2335 col_n[24] row_n[0] 0.23fF
C2336 col_n[21] ctop 2.02fF
C2337 col_n[28] row_n[2] 0.23fF
C2338 VDD col[19] 4.17fF
C2339 col_n[30] row_n[3] 0.23fF
C2340 a_16018_5142# a_16018_4138# 1.00fF
C2341 a_32994_5142# a_33086_5142# 0.26fF
C2342 a_25054_12170# col_n[22] 0.28fF
C2343 a_10906_18194# m2_10768_18014# 0.16fF
C2344 a_1962_9198# a_14010_9158# 0.27fF
C2345 a_3270_3174# vcm 0.22fF
C2346 a_4974_11166# row_n[9] 0.17fF
C2347 a_17022_14178# a_18026_14178# 0.97fF
C2348 a_2346_14220# a_32994_14178# 0.35fF
C2349 a_1962_10202# col[7] 0.11fF
C2350 m2_6752_18014# col[4] 0.28fF
C2351 a_2346_15224# rowon_n[13] 0.26fF
C2352 a_23046_13174# vcm 0.62fF
C2353 a_2966_7150# ctop 3.42fF
C2354 a_26058_6146# VDD 0.52fF
C2355 a_2346_6188# a_8990_6146# 0.19fF
C2356 a_1962_6186# a_7286_6186# 0.14fF
C2357 a_5886_6146# a_5978_6146# 0.26fF
C2358 a_2346_9200# col[27] 0.15fF
C2359 a_4974_8154# rowoff_n[6] 0.10fF
C2360 a_1962_11206# a_27062_11166# 0.27fF
C2361 a_16322_7190# vcm 0.22fF
C2362 a_1962_18234# col_n[26] 0.13fF
C2363 a_2346_16228# vcm 0.40fF
C2364 a_10998_17190# rowoff_n[15] 0.10fF
C2365 a_15014_6146# rowoff_n[4] 0.10fF
C2366 a_13006_9158# m2_13204_9406# 0.16fF
C2367 a_7986_5142# col_n[5] 0.28fF
C2368 a_2346_3176# a_3878_3134# 0.35fF
C2369 a_2874_3134# a_2966_3134# 0.26fF
C2370 a_5886_9158# VDD 0.23fF
C2371 a_29070_9158# a_29070_8154# 1.00fF
C2372 a_2346_8196# a_22042_8154# 0.19fF
C2373 a_1962_8194# a_20338_8194# 0.14fF
C2374 a_24050_14178# row_n[12] 0.17fF
C2375 m2_2736_1950# m2_2736_946# 0.99fF
C2376 a_25054_4138# rowoff_n[2] 0.10fF
C2377 a_29374_11206# vcm 0.22fF
C2378 a_1962_12210# col_n[7] 0.13fF
C2379 a_10998_5142# ctop 3.58fF
C2380 m2_22816_18014# col_n[20] 0.25fF
C2381 a_23046_15182# col[20] 0.29fF
C2382 a_18938_13174# VDD 0.23fF
C2383 a_1962_10202# a_33390_10202# 0.14fF
C2384 a_18938_10162# a_19030_10162# 0.26fF
C2385 a_12002_12170# rowon_n[10] 0.14fF
C2386 a_2346_2172# a_11910_2130# 0.35fF
C2387 m2_28840_18014# m3_28972_18146# 2.78fF
C2388 a_24050_9158# ctop 3.58fF
C2389 a_2346_5184# col[18] 0.15fF
C2390 a_27062_2130# rowon_n[0] 0.14fF
C2391 a_31990_17190# VDD 0.24fF
C2392 col[29] rowoff_n[9] 0.11fF
C2393 col[22] rowoff_n[2] 0.11fF
C2394 col[21] rowoff_n[1] 0.11fF
C2395 col[26] rowoff_n[6] 0.11fF
C2396 col[25] rowoff_n[5] 0.11fF
C2397 col[24] rowoff_n[4] 0.11fF
C2398 col[23] rowoff_n[3] 0.11fF
C2399 col[20] rowoff_n[0] 0.11fF
C2400 col[27] rowoff_n[7] 0.11fF
C2401 col[28] rowoff_n[8] 0.11fF
C2402 a_4974_8154# vcm 0.62fF
C2403 a_5978_8154# col[3] 0.29fF
C2404 a_9994_10162# m2_10192_10410# 0.16fF
C2405 a_2346_4180# a_24962_4138# 0.35fF
C2406 a_13006_4138# a_14010_4138# 0.97fF
C2407 a_4974_2130# row_n[0] 0.17fF
C2408 a_1962_1166# col[25] 0.11fF
C2409 a_29982_18194# m2_29844_18014# 0.16fF
C2410 a_2346_6188# rowon_n[4] 0.26fF
C2411 a_1962_14218# col[27] 0.11fF
C2412 a_31990_14178# a_32082_14178# 0.26fF
C2413 a_15014_14178# a_15014_13174# 1.00fF
C2414 a_23958_10162# rowoff_n[8] 0.24fF
C2415 a_23046_17190# col_n[20] 0.28fF
C2416 a_31078_15182# rowon_n[13] 0.14fF
C2417 a_25966_13174# rowoff_n[11] 0.24fF
C2418 a_18026_12170# vcm 0.62fF
C2419 a_24050_4138# col[21] 0.29fF
C2420 a_1962_1166# a_19030_1126# 0.26fF
C2421 a_1962_8194# sample 0.14fF
C2422 a_21038_5142# VDD 0.52fF
C2423 a_2966_18194# vcm 0.12fF
C2424 m2_26832_946# VDD 0.62fF
C2425 a_2966_6146# a_2966_5142# 1.00fF
C2426 col[13] rowoff_n[10] 0.11fF
C2427 a_33998_8154# rowoff_n[6] 0.24fF
C2428 a_8990_15182# row_n[13] 0.17fF
C2429 a_11302_6186# vcm 0.22fF
C2430 a_1962_15222# a_5278_15222# 0.14fF
C2431 a_4882_15182# a_4974_15182# 0.26fF
C2432 a_2346_15224# a_6982_15182# 0.19fF
C2433 a_31078_16186# vcm 0.62fF
C2434 a_1962_3174# a_32082_3134# 0.27fF
C2435 a_24050_5142# row_n[3] 0.17fF
C2436 a_2346_1168# col[9] 0.14fF
C2437 a_34090_9158# VDD 0.54fF
C2438 a_2346_14220# col[11] 0.15fF
C2439 a_26058_8154# a_27062_8154# 0.97fF
C2440 a_5978_10162# col_n[3] 0.28fF
C2441 a_1962_3174# col_n[25] 0.13fF
C2442 a_24354_10202# vcm 0.22fF
C2443 a_1962_17230# a_18330_17230# 0.14fF
C2444 a_2346_17232# a_20034_17190# 0.19fF
C2445 a_1962_16226# col_n[27] 0.13fF
C2446 col_n[13] col[13] 0.72fF
C2447 rowon_n[15] ctop 1.19fF
C2448 VDD col[30] 4.17fF
C2449 vcm col[26] 5.84fF
C2450 rowon_n[7] rowon_n[6] 0.15fF
C2451 a_5978_4138# ctop 3.58fF
C2452 m3_1864_6098# ctop 0.23fF
C2453 a_6982_11166# m2_7180_11414# 0.16fF
C2454 a_24050_6146# col_n[21] 0.28fF
C2455 a_13918_12170# VDD 0.23fF
C2456 a_1962_10202# col[18] 0.11fF
C2457 a_12002_3134# rowon_n[1] 0.14fF
C2458 a_13006_14178# rowoff_n[12] 0.10fF
C2459 a_19030_8154# ctop 3.58fF
C2460 a_26970_16186# VDD 0.23fF
C2461 a_2346_11208# a_9902_11166# 0.35fF
C2462 a_14010_2130# m2_14208_2378# 0.16fF
C2463 a_2346_18236# a_3878_18194# 0.35fF
C2464 a_16018_16186# rowon_n[14] 0.14fF
C2465 a_10998_4138# a_10998_3134# 1.00fF
C2466 a_27974_4138# a_28066_4138# 0.26fF
C2467 a_32082_12170# ctop 3.58fF
C2468 a_2346_10204# col[2] 0.15fF
C2469 a_1962_8194# a_3970_8154# 0.27fF
C2470 a_3970_13174# col[1] 0.29fF
C2471 a_31078_6146# rowon_n[4] 0.14fF
C2472 a_12002_13174# a_13006_13174# 0.97fF
C2473 a_2346_13216# a_22954_13174# 0.35fF
C2474 a_1962_12210# col_n[18] 0.13fF
C2475 a_13006_11166# vcm 0.62fF
C2476 a_16018_4138# VDD 0.52fF
C2477 a_3970_12170# m2_4168_12418# 0.16fF
C2478 m3_30980_1078# VDD 0.14fF
C2479 a_22042_9158# col[19] 0.29fF
C2480 a_1962_6186# col[9] 0.11fF
C2481 a_8990_6146# row_n[4] 0.17fF
C2482 a_1962_10202# a_17022_10162# 0.27fF
C2483 a_6282_5182# vcm 0.22fF
C2484 a_26058_15182# vcm 0.62fF
C2485 a_2346_5184# col[29] 0.15fF
C2486 m2_4744_18014# m3_5880_18146# 0.13fF
C2487 col[31] rowoff_n[0] 0.11fF
C2488 a_29070_8154# VDD 0.52fF
C2489 a_6890_7150# rowoff_n[5] 0.24fF
C2490 a_2346_7192# a_12002_7150# 0.19fF
C2491 a_1962_7190# a_10298_7190# 0.14fF
C2492 a_1962_15222# m2_34864_15002# 0.17fF
C2493 a_24050_8154# a_24050_7150# 1.00fF
C2494 a_1962_12210# a_30074_12170# 0.27fF
C2495 a_19334_9198# vcm 0.22fF
C2496 a_25054_17190# a_26058_17190# 0.97fF
C2497 a_3970_15182# col_n[1] 0.28fF
C2498 a_16930_5142# rowoff_n[3] 0.24fF
C2499 a_4974_2130# col[2] 0.29fF
C2500 a_28066_9158# row_n[7] 0.17fF
C2501 a_8898_11166# VDD 0.23fF
C2502 a_2346_9200# a_25054_9158# 0.19fF
C2503 a_13918_9158# a_14010_9158# 0.26fF
C2504 a_1962_9198# a_23350_9198# 0.14fF
C2505 a_22042_11166# col_n[19] 0.28fF
C2506 a_26970_3134# rowoff_n[1] 0.24fF
C2507 a_1962_8194# col_n[9] 0.13fF
C2508 m2_1732_4962# m2_2160_5390# 0.16fF
C2509 a_32386_13214# vcm 0.22fF
C2510 col[24] rowoff_n[10] 0.11fF
C2511 a_14010_7150# ctop 3.58fF
C2512 a_2966_5142# VDD 0.56fF
C2513 a_1962_2170# col[0] 0.11fF
C2514 a_1962_15222# col[2] 0.11fF
C2515 a_21950_15182# VDD 0.23fF
C2516 a_16018_7150# rowon_n[5] 0.14fF
C2517 a_1962_1166# m2_2736_946# 0.18fF
C2518 a_2346_1168# col[20] 0.14fF
C2519 a_2346_14220# col[22] 0.15fF
C2520 a_2346_3176# a_14922_3134# 0.35fF
C2521 a_7986_3134# a_8990_3134# 0.97fF
C2522 a_27062_11166# ctop 3.58fF
C2523 a_6982_2130# m3_6884_1078# 0.15fF
C2524 a_2346_18236# ctop 0.22fF
C2525 a_4974_4138# col_n[2] 0.28fF
C2526 row_n[10] ctop 1.65fF
C2527 col_n[18] col[19] 5.98fF
C2528 rowon_n[4] row_n[4] 19.75fF
C2529 a_26970_13174# a_27062_13174# 0.26fF
C2530 a_9994_13174# a_9994_12170# 1.00fF
C2531 a_7986_10162# vcm 0.62fF
C2532 a_15014_11166# rowoff_n[9] 0.10fF
C2533 col[8] rowoff_n[11] 0.11fF
C2534 m2_9764_18014# m2_10192_18442# 0.16fF
C2535 a_10998_3134# VDD 0.52fF
C2536 a_1962_10202# col[29] 0.11fF
C2537 a_2346_5184# a_27974_5142# 0.35fF
C2538 a_25054_9158# rowoff_n[7] 0.10fF
C2539 a_20034_14178# col[17] 0.29fF
C2540 a_1962_4178# vcm 6.95fF
C2541 a_1962_17230# col_n[2] 0.13fF
C2542 m2_34864_8978# m2_34864_7974# 0.99fF
C2543 m2_1732_17010# rowon_n[15] 0.11fF
C2544 a_29070_15182# rowoff_n[13] 0.10fF
C2545 a_21038_14178# vcm 0.62fF
C2546 a_1962_2170# a_22042_2130# 0.27fF
C2547 a_24050_7150# VDD 0.52fF
C2548 a_21038_7150# a_22042_7150# 0.97fF
C2549 a_32082_15182# m2_32280_15430# 0.16fF
C2550 a_13006_10162# row_n[8] 0.17fF
C2551 a_23046_17190# a_23046_16186# 1.00fF
C2552 a_14314_8194# vcm 0.22fF
C2553 a_1962_16226# a_8290_16226# 0.14fF
C2554 a_2346_16228# a_9994_16186# 0.19fF
C2555 a_34090_3134# m2_34288_3382# 0.16fF
C2556 a_34090_18194# vcm 0.12fF
C2557 a_2346_10204# col[13] 0.15fF
C2558 a_2966_17190# m2_3164_17438# 0.16fF
C2559 a_1962_12210# col_n[29] 0.13fF
C2560 a_2966_13174# a_3970_13174# 0.97fF
C2561 a_27366_12210# vcm 0.22fF
C2562 a_2346_12212# rowoff_n[10] 4.09fF
C2563 a_1962_1166# a_28370_1166# 0.14fF
C2564 a_20034_16186# col_n[17] 0.28fF
C2565 a_1962_6186# col[20] 0.11fF
C2566 a_8990_6146# ctop 3.58fF
C2567 a_32082_13174# row_n[11] 0.17fF
C2568 m3_26964_18146# VDD 0.38fF
C2569 a_21038_3134# col[18] 0.29fF
C2570 a_16930_14178# VDD 0.23fF
C2571 m2_20232_1374# a_20034_1126# 0.16fF
C2572 m2_5748_18014# ctop 0.18fF
C2573 a_16930_16186# rowoff_n[14] 0.24fF
C2574 a_22954_3134# a_23046_3134# 0.26fF
C2575 a_5978_3134# a_5978_2130# 1.00fF
C2576 a_22042_10162# ctop 3.58fF
C2577 a_29070_16186# m2_29268_16434# 0.16fF
C2578 a_29982_18194# VDD 0.33fF
C2579 m2_34864_18014# vcm 0.34fF
C2580 a_2346_12212# a_12914_12170# 0.35fF
C2581 a_6982_12170# a_7986_12170# 0.97fF
C2582 a_20034_11166# rowon_n[9] 0.14fF
C2583 a_2346_6188# col[4] 0.15fF
C2584 a_31078_4138# m2_31276_4386# 0.16fF
C2585 m2_5748_946# m3_4876_1078# 0.13fF
C2586 a_5978_2130# VDD 0.55fF
C2587 m3_33992_1078# ctop 0.37fF
C2588 a_1962_9198# a_6982_9158# 0.27fF
C2589 a_1962_8194# col_n[20] 0.13fF
C2590 a_21038_5142# col_n[18] 0.28fF
C2591 a_2346_14220# a_25966_14178# 0.35fF
C2592 a_2346_18236# a_35002_18194# 0.35fF
C2593 a_16018_13174# vcm 0.62fF
C2594 a_2346_6188# m2_1732_5966# 0.12fF
C2595 a_1962_2170# col[11] 0.11fF
C2596 a_1962_15222# col[13] 0.11fF
C2597 a_19030_6146# VDD 0.52fF
C2598 a_19030_7150# a_19030_6146# 1.00fF
C2599 a_3878_15182# VDD 0.23fF
C2600 a_1962_11206# a_20034_11166# 0.27fF
C2601 a_2966_12170# col[0] 0.29fF
C2602 a_9294_7190# vcm 0.22fF
C2603 a_20034_16186# a_21038_16186# 0.97fF
C2604 a_3970_17190# rowoff_n[15] 0.10fF
C2605 a_29070_17190# vcm 0.60fF
C2606 m2_25828_18014# VDD 0.93fF
C2607 a_2346_18236# col[5] 0.14fF
C2608 a_7986_6146# rowoff_n[4] 0.10fF
C2609 a_32082_10162# VDD 0.52fF
C2610 col_n[24] col[24] 0.72fF
C2611 rowon_n[4] ctop 1.40fF
C2612 a_8898_8154# a_8990_8154# 0.26fF
C2613 a_1962_8194# a_13310_8194# 0.14fF
C2614 a_2346_8196# a_15014_8154# 0.19fF
C2615 a_26058_17190# m2_26256_17438# 0.16fF
C2616 a_17022_14178# row_n[12] 0.17fF
C2617 a_1962_13214# a_33086_13174# 0.27fF
C2618 col[19] rowoff_n[11] 0.11fF
C2619 m2_1732_8978# sample 0.19fF
C2620 a_18026_4138# rowoff_n[2] 0.10fF
C2621 m2_34864_2954# ctop 0.17fF
C2622 a_32082_4138# row_n[2] 0.17fF
C2623 a_31078_12170# rowoff_n[10] 0.10fF
C2624 a_22346_11206# vcm 0.22fF
C2625 a_28066_5142# m2_28264_5390# 0.16fF
C2626 a_3970_5142# ctop 3.57fF
C2627 a_11910_13174# VDD 0.23fF
C2628 a_1962_4178# col_n[11] 0.13fF
C2629 a_1962_10202# a_26362_10202# 0.14fF
C2630 a_2346_10204# a_28066_10162# 0.19fF
C2631 a_32082_11166# a_32082_10162# 1.00fF
C2632 a_1962_17230# col_n[13] 0.13fF
C2633 a_28066_2130# rowoff_n[0] 0.10fF
C2634 a_19030_8154# col[16] 0.29fF
C2635 a_2966_14178# vcm 0.61fF
C2636 a_4974_12170# rowon_n[10] 0.14fF
C2637 a_2346_2172# a_4882_2130# 0.35fF
C2638 a_1962_11206# col[4] 0.11fF
C2639 m2_19804_18014# m3_18932_18146# 0.13fF
C2640 a_17022_9158# ctop 3.58fF
C2641 a_20034_2130# rowon_n[0] 0.14fF
C2642 a_24962_17190# VDD 0.24fF
C2643 col[3] rowoff_n[12] 0.11fF
C2644 a_21950_12170# a_22042_12170# 0.26fF
C2645 a_4974_12170# a_4974_11166# 1.00fF
C2646 a_2346_10204# col[24] 0.15fF
C2647 a_35002_2130# VDD 0.30fF
C2648 a_2346_4180# a_17934_4138# 0.35fF
C2649 a_30074_13174# ctop 3.58fF
C2650 a_1962_9198# a_34394_9198# 0.14fF
C2651 a_16930_10162# rowoff_n[8] 0.24fF
C2652 a_24050_15182# rowon_n[13] 0.14fF
C2653 a_1962_6186# col[31] 0.11fF
C2654 a_10998_12170# vcm 0.62fF
C2655 a_18938_13174# rowoff_n[11] 0.24fF
C2656 a_19030_10162# col_n[16] 0.28fF
C2657 a_25054_6146# m2_25252_6394# 0.16fF
C2658 a_14010_5142# VDD 0.52fF
C2659 a_2346_6188# a_30986_6146# 0.35fF
C2660 a_16018_6146# a_17022_6146# 0.97fF
C2661 a_26970_8154# rowoff_n[6] 0.24fF
C2662 a_1962_13214# col_n[4] 0.13fF
C2663 a_21038_17190# m3_20940_18146# 0.15fF
C2664 a_4274_6186# vcm 0.22fF
C2665 a_18026_16186# a_18026_15182# 1.00fF
C2666 a_32994_17190# rowoff_n[15] 0.24fF
C2667 a_24050_16186# vcm 0.62fF
C2668 a_1962_3174# a_25054_3134# 0.27fF
C2669 a_17022_5142# row_n[3] 0.17fF
C2670 a_27062_9158# VDD 0.52fF
C2671 a_35094_1126# vcm 0.12fF
C2672 a_2346_6188# col[15] 0.15fF
C2673 m2_34864_3958# rowon_n[2] 0.13fF
C2674 a_17326_10202# vcm 0.22fF
C2675 a_2346_17232# a_13006_17190# 0.19fF
C2676 a_1962_17230# a_11302_17230# 0.14fF
C2677 a_7894_17190# a_7986_17190# 0.26fF
C2678 m3_29976_18146# ctop 0.23fF
C2679 a_1962_8194# col_n[31] 0.13fF
C2680 a_6890_12170# VDD 0.23fF
C2681 a_29070_10162# a_30074_10162# 0.97fF
C2682 a_4974_3134# rowon_n[1] 0.14fF
C2683 a_1962_2170# col[22] 0.11fF
C2684 a_1962_15222# col[24] 0.11fF
C2685 a_5978_14178# rowoff_n[12] 0.10fF
C2686 a_30378_14218# vcm 0.22fF
C2687 a_17022_13174# col[14] 0.29fF
C2688 a_1962_2170# a_31382_2170# 0.14fF
C2689 a_2346_2172# a_33086_2130# 0.19fF
C2690 a_17934_2130# a_18026_2130# 0.26fF
C2691 a_22042_7150# m2_22240_7398# 0.16fF
C2692 a_12002_8154# ctop 3.58fF
C2693 a_19942_16186# VDD 0.23fF
C2694 a_2346_18236# col[16] 0.14fF
C2695 col_n[29] col[30] 5.92fF
C2696 sw_n ctop 0.25fF
C2697 a_29982_1126# VDD 0.44fF
C2698 a_8990_16186# rowon_n[14] 0.14fF
C2699 a_25054_12170# ctop 3.58fF
C2700 col[30] rowoff_n[11] 0.11fF
C2701 a_24050_6146# rowon_n[4] 0.14fF
C2702 a_2346_2172# col[6] 0.15fF
C2703 a_2346_13216# a_15926_13174# 0.35fF
C2704 a_2346_15224# col[8] 0.15fF
C2705 a_5978_11166# vcm 0.62fF
C2706 m2_1732_5966# row_n[4] 0.13fF
C2707 a_1962_4178# col_n[22] 0.13fF
C2708 a_8990_4138# VDD 0.52fF
C2709 m3_2868_1078# VDD 0.17fF
C2710 a_30986_6146# a_31078_6146# 0.26fF
C2711 a_1962_17230# col_n[24] 0.13fF
C2712 a_14010_6146# a_14010_5142# 1.00fF
C2713 a_17022_15182# col_n[14] 0.28fF
C2714 a_1962_10202# a_9994_10162# 0.27fF
C2715 a_18026_2130# col[15] 0.29fF
C2716 a_15014_15182# a_16018_15182# 0.97fF
C2717 a_2346_15224# a_28978_15182# 0.35fF
C2718 a_1962_11206# col[15] 0.11fF
C2719 a_19030_15182# vcm 0.62fF
C2720 a_19030_8154# m2_19228_8402# 0.16fF
C2721 a_22042_8154# VDD 0.52fF
C2722 col[14] rowoff_n[12] 0.11fF
C2723 a_1962_7190# a_3270_7190# 0.14fF
C2724 a_2346_7192# a_4974_7150# 0.19fF
C2725 a_1962_12210# a_23046_12170# 0.27fF
C2726 m2_14784_946# m3_15920_1078# 0.13fF
C2727 a_12306_9198# vcm 0.22fF
C2728 a_9902_5142# rowoff_n[3] 0.24fF
C2729 a_21038_9158# row_n[7] 0.17fF
C2730 m2_26832_946# m3_25960_1078# 0.13fF
C2731 a_1962_9198# a_16322_9198# 0.14fF
C2732 a_2346_9200# a_18026_9158# 0.19fF
C2733 a_27062_10162# a_27062_9158# 1.00fF
C2734 a_19942_3134# rowoff_n[1] 0.24fF
C2735 a_35002_14178# rowoff_n[12] 0.24fF
C2736 a_25358_13214# vcm 0.22fF
C2737 a_18026_4138# col_n[15] 0.28fF
C2738 a_6982_7150# ctop 3.58fF
C2739 a_1962_13214# col_n[15] 0.13fF
C2740 a_14922_15182# VDD 0.23fF
C2741 a_1962_11206# a_29374_11206# 0.14fF
C2742 a_2346_11208# a_31078_11166# 0.19fF
C2743 a_16930_11166# a_17022_11166# 0.26fF
C2744 a_8990_7150# rowon_n[5] 0.14fF
C2745 a_1962_7190# col[6] 0.11fF
C2746 a_33086_14178# col[30] 0.29fF
C2747 a_2346_3176# a_7894_3134# 0.35fF
C2748 a_16018_9158# m2_16216_9406# 0.16fF
C2749 a_24050_2130# m2_23820_946# 0.99fF
C2750 a_20034_11166# ctop 3.58fF
C2751 a_35002_17190# m2_34864_17010# 0.16fF
C2752 a_2346_6188# col[26] 0.15fF
C2753 a_7986_11166# rowoff_n[9] 0.10fF
C2754 m2_2736_18014# m2_3164_18442# 0.16fF
C2755 a_3970_3134# VDD 0.52fF
C2756 a_10998_5142# a_12002_5142# 0.97fF
C2757 a_2346_5184# a_20946_5142# 0.35fF
C2758 a_33086_15182# ctop 3.57fF
C2759 a_28066_10162# rowon_n[8] 0.14fF
C2760 a_18026_9158# rowoff_n[7] 0.10fF
C2761 a_13006_15182# a_13006_14178# 1.00fF
C2762 a_29982_15182# a_30074_15182# 0.26fF
C2763 a_14010_14178# vcm 0.62fF
C2764 a_22042_15182# rowoff_n[13] 0.10fF
C2765 a_16018_7150# col[13] 0.29fF
C2766 m2_34864_8978# VDD 1.01fF
C2767 a_1962_2170# a_15014_2130# 0.27fF
C2768 a_1962_9198# col_n[6] 0.13fF
C2769 m2_33860_18014# m3_33992_18146# 2.78fF
C2770 a_17022_7150# VDD 0.52fF
C2771 a_28066_7150# rowoff_n[5] 0.10fF
C2772 a_2346_7192# a_33998_7150# 0.35fF
C2773 a_5978_10162# row_n[8] 0.17fF
C2774 a_35494_17552# VDD 0.11fF
C2775 a_33086_16186# col_n[30] 0.28fF
C2776 a_2346_18236# col[27] 0.14fF
C2777 a_34090_3134# col[31] 0.29fF
C2778 ctop col[4] 1.98fF
C2779 a_7286_8194# vcm 0.22fF
C2780 a_2346_16228# a_2874_16186# 0.35fF
C2781 a_27062_18194# vcm 0.12fF
C2782 a_1962_4178# a_28066_4138# 0.27fF
C2783 a_13006_10162# m2_13204_10410# 0.16fF
C2784 a_30074_11166# VDD 0.52fF
C2785 m3_27968_1078# m3_28972_1078# 0.22fF
C2786 a_2346_2172# col[17] 0.15fF
C2787 a_24050_9158# a_25054_9158# 0.97fF
C2788 a_2346_15224# col[19] 0.15fF
C2789 m2_2736_1950# col_n[0] 0.28fF
C2790 m2_1732_5966# ctop 0.17fF
C2791 a_20338_12210# vcm 0.22fF
C2792 a_1962_1166# a_21342_1166# 0.14fF
C2793 a_25054_13174# row_n[11] 0.17fF
C2794 m2_34864_946# VDD 1.11fF
C2795 a_16018_9158# col_n[13] 0.28fF
C2796 a_1962_18234# col[9] 0.11fF
C2797 a_9902_14178# VDD 0.23fF
C2798 a_1962_11206# col[26] 0.11fF
C2799 a_9902_16186# rowoff_n[14] 0.24fF
C2800 a_33390_16226# vcm 0.22fF
C2801 col[25] rowoff_n[12] 0.11fF
C2802 m2_16792_18014# col_n[14] 0.25fF
C2803 a_34090_5142# col_n[31] 0.28fF
C2804 a_2346_3176# a_2346_2172# 0.22fF
C2805 a_1962_3174# a_35398_3174# 0.14fF
C2806 a_15014_10162# ctop 3.58fF
C2807 a_22954_18194# VDD 0.34fF
C2808 m2_20808_18014# vcm 0.28fF
C2809 a_2346_12212# a_5886_12170# 0.35fF
C2810 a_13006_11166# rowon_n[9] 0.14fF
C2811 a_32994_3134# VDD 0.23fF
C2812 a_2966_9158# row_n[7] 0.16fF
C2813 m3_5880_1078# ctop 0.23fF
C2814 a_8990_5142# a_8990_4138# 1.00fF
C2815 a_25966_5142# a_26058_5142# 0.26fF
C2816 a_9994_11166# m2_10192_11414# 0.16fF
C2817 a_28066_14178# ctop 3.58fF
C2818 a_2346_11208# col[10] 0.15fF
C2819 a_9994_14178# a_10998_14178# 0.97fF
C2820 a_2346_14220# a_18938_14178# 0.35fF
C2821 col[9] rowoff_n[13] 0.11fF
C2822 a_2346_18236# a_27974_18194# 0.35fF
C2823 a_1962_13214# col_n[26] 0.13fF
C2824 a_8990_13174# vcm 0.62fF
C2825 m2_6752_946# col_n[4] 0.37fF
C2826 a_12002_6146# VDD 0.52fF
C2827 a_14010_12170# col[11] 0.29fF
C2828 a_1962_7190# col[17] 0.11fF
C2829 a_32082_14178# rowon_n[12] 0.14fF
C2830 a_1962_11206# a_13006_11166# 0.27fF
C2831 a_2346_16228# a_31990_16186# 0.35fF
C2832 a_17022_2130# m2_17220_2378# 0.16fF
C2833 a_22042_17190# vcm 0.60fF
C2834 m2_11772_18014# VDD 1.06fF
C2835 a_32082_8154# col[29] 0.29fF
C2836 a_1962_18234# m2_26832_18014# 0.18fF
C2837 a_25054_10162# VDD 0.52fF
C2838 a_1962_8194# a_6282_8194# 0.14fF
C2839 a_2346_8196# a_7986_8154# 0.19fF
C2840 a_22042_9158# a_22042_8154# 1.00fF
C2841 a_9994_14178# row_n[12] 0.17fF
C2842 a_1962_13214# a_26058_13174# 0.27fF
C2843 a_32082_2130# vcm 0.62fF
C2844 a_24050_12170# rowoff_n[10] 0.10fF
C2845 a_25054_4138# row_n[2] 0.17fF
C2846 a_10998_4138# rowoff_n[2] 0.10fF
C2847 a_15318_11206# vcm 0.22fF
C2848 a_2346_5184# a_1962_5182# 2.62fF
C2849 a_6982_12170# m2_7180_12418# 0.16fF
C2850 a_2346_7192# col[1] 0.15fF
C2851 a_2346_18236# m2_21812_18014# 0.19fF
C2852 a_4882_13174# VDD 0.23fF
C2853 a_11910_10162# a_12002_10162# 0.26fF
C2854 a_1962_10202# a_19334_10202# 0.14fF
C2855 a_2346_10204# a_21038_10162# 0.19fF
C2856 a_21038_2130# rowoff_n[0] 0.10fF
C2857 a_14010_14178# col_n[11] 0.28fF
C2858 a_1962_9198# col_n[17] 0.13fF
C2859 a_28370_15222# vcm 0.22fF
C2860 a_33086_3134# a_34090_3134# 0.97fF
C2861 a_20034_1126# m3_20940_1078# 0.14fF
C2862 m2_9764_18014# m3_10900_18146# 0.13fF
C2863 a_9994_9158# ctop 3.58fF
C2864 a_29070_17190# row_n[15] 0.17fF
C2865 a_1962_3174# col[8] 0.11fF
C2866 a_32082_10162# col_n[29] 0.28fF
C2867 a_13006_2130# rowon_n[0] 0.14fF
C2868 a_17934_17190# VDD 0.24fF
C2869 ctop col[15] 1.99fF
C2870 col[4] col[5] 0.20fF
C2871 a_1962_16226# col[10] 0.11fF
C2872 a_2346_12212# a_34090_12170# 0.19fF
C2873 a_1962_12210# a_32386_12210# 0.14fF
C2874 a_27974_2130# VDD 0.23fF
C2875 a_2346_2172# col[28] 0.15fF
C2876 a_2346_4180# a_10906_4138# 0.35fF
C2877 a_2346_15224# col[30] 0.15fF
C2878 a_5978_4138# a_6982_4138# 0.97fF
C2879 a_23046_13174# ctop 3.58fF
C2880 m3_34996_6098# m3_34996_5094# 0.22fF
C2881 a_7986_14178# a_7986_13174# 1.00fF
C2882 a_24962_14178# a_25054_14178# 0.26fF
C2883 a_9902_10162# rowoff_n[8] 0.24fF
C2884 a_17022_15182# rowon_n[13] 0.14fF
C2885 a_3970_12170# vcm 0.62fF
C2886 a_11910_13174# rowoff_n[11] 0.24fF
C2887 a_3878_1126# a_3970_1126# 0.26fF
C2888 a_1962_18234# col[20] 0.11fF
C2889 a_6982_5142# VDD 0.52fF
C2890 a_32082_5142# rowon_n[3] 0.14fF
C2891 a_15014_3134# col_n[12] 0.28fF
C2892 a_2346_6188# a_23958_6146# 0.35fF
C2893 a_3970_13174# m2_4168_13422# 0.16fF
C2894 a_2346_16228# ctop 1.57fF
C2895 a_19942_8154# rowoff_n[6] 0.24fF
C2896 a_12002_17190# col[9] 0.29fF
C2897 a_1962_5182# col_n[8] 0.13fF
C2898 m2_1732_11990# m2_1732_10986# 0.99fF
C2899 a_1962_1166# m2_10768_946# 0.18fF
C2900 a_25966_17190# rowoff_n[15] 0.24fF
C2901 a_17022_16186# vcm 0.62fF
C2902 a_9994_5142# row_n[3] 0.17fF
C2903 a_29982_6146# rowoff_n[4] 0.24fF
C2904 a_1962_3174# a_18026_3134# 0.27fF
C2905 a_9994_2130# m3_9896_1078# 0.15fF
C2906 a_20034_9158# VDD 0.52fF
C2907 a_1962_16226# m2_34864_16006# 0.17fF
C2908 a_1962_8194# a_1962_7190# 0.16fF
C2909 a_19030_8154# a_20034_8154# 0.97fF
C2910 a_1962_12210# col[1] 0.11fF
C2911 a_30074_13174# col[27] 0.29fF
C2912 a_27062_1126# vcm 0.12fF
C2913 m2_1732_7974# rowon_n[6] 0.11fF
C2914 a_10298_10202# vcm 0.22fF
C2915 a_2346_17232# a_5978_17190# 0.19fF
C2916 a_1962_17230# a_4274_17230# 0.14fF
C2917 a_2346_11208# col[21] 0.15fF
C2918 a_1962_5182# a_31078_5142# 0.27fF
C2919 a_33086_13174# VDD 0.52fF
C2920 col[20] rowoff_n[13] 0.11fF
C2921 VDD rowoff_n[2] 1.17fF
C2922 vcm rowoff_n[6] 0.20fF
C2923 sample_n rowoff_n[3] 0.38fF
C2924 a_29070_8154# row_n[6] 0.17fF
C2925 a_23350_14218# vcm 0.22fF
C2926 a_1962_2170# a_24354_2170# 0.14fF
C2927 a_31078_3134# a_31078_2130# 1.00fF
C2928 a_2346_2172# a_26058_2130# 0.19fF
C2929 a_4974_8154# ctop 3.58fF
C2930 m2_34864_17010# m3_34996_16138# 0.15fF
C2931 a_1962_7190# col[28] 0.11fF
C2932 a_13006_6146# col[10] 0.29fF
C2933 a_12914_16186# VDD 0.23fF
C2934 a_32082_12170# a_33086_12170# 0.97fF
C2935 a_1962_1166# col_n[0] 0.13fF
C2936 a_30074_15182# col_n[27] 0.28fF
C2937 a_1962_14218# col_n[1] 0.13fF
C2938 a_2874_2130# m2_2736_1950# 0.16fF
C2939 a_31078_2130# col[28] 0.29fF
C2940 a_22954_1126# VDD 0.44fF
C2941 a_3970_4138# a_3970_3134# 1.00fF
C2942 a_20946_4138# a_21038_4138# 0.26fF
C2943 a_18026_12170# ctop 3.58fF
C2944 col[4] rowoff_n[14] 0.11fF
C2945 a_17022_17190# m2_16792_18014# 1.00fF
C2946 a_17022_6146# rowon_n[4] 0.14fF
C2947 a_4974_13174# a_5978_13174# 0.97fF
C2948 a_2346_13216# a_8898_13174# 0.35fF
C2949 a_2346_7192# col[12] 0.15fF
C2950 m3_1864_14130# VDD 0.25fF
C2951 a_31078_16186# ctop 3.57fF
C2952 a_2346_10204# a_2966_10162# 0.21fF
C2953 a_1962_9198# col_n[28] 0.13fF
C2954 a_13006_8154# col_n[10] 0.28fF
C2955 a_2346_15224# a_21950_15182# 0.35fF
C2956 a_12002_15182# vcm 0.62fF
C2957 m2_1732_11990# VDD 1.02fF
C2958 a_1962_3174# col[19] 0.11fF
C2959 VDD col_n[4] 4.98fF
C2960 ctop col[26] 1.98fF
C2961 a_15014_8154# VDD 0.52fF
C2962 a_1962_16226# col[21] 0.11fF
C2963 a_33998_8154# a_34090_8154# 0.26fF
C2964 a_17022_8154# a_17022_7150# 1.00fF
C2965 a_32082_16186# m2_32280_16434# 0.16fF
C2966 a_31078_4138# col_n[28] 0.28fF
C2967 a_1962_12210# a_16018_12170# 0.27fF
C2968 a_5278_9198# vcm 0.22fF
C2969 a_2346_17232# a_35002_17190# 0.35fF
C2970 a_18026_17190# a_19030_17190# 0.97fF
C2971 m2_31852_18014# col[29] 0.28fF
C2972 a_34090_4138# m2_34288_4386# 0.16fF
C2973 a_2346_5184# rowoff_n[3] 4.09fF
C2974 m2_10768_946# m3_9896_1078# 0.13fF
C2975 a_14010_9158# row_n[7] 0.17fF
C2976 a_28066_12170# VDD 0.52fF
C2977 m3_23952_18146# m3_24956_18146# 0.22fF
C2978 a_6890_9158# a_6982_9158# 0.26fF
C2979 a_2346_9200# a_10998_9158# 0.19fF
C2980 a_1962_9198# a_9294_9198# 0.14fF
C2981 a_35094_4138# vcm 0.12fF
C2982 a_1962_14218# a_29070_14178# 0.27fF
C2983 a_12914_3134# rowoff_n[1] 0.24fF
C2984 a_1962_18234# col[31] 0.11fF
C2985 a_18330_13214# vcm 0.22fF
C2986 a_27974_14178# rowoff_n[12] 0.24fF
C2987 a_2346_3176# col[3] 0.15fF
C2988 a_28066_2130# a_29070_2130# 0.97fF
C2989 a_2346_16228# col[5] 0.15fF
C2990 m2_34864_13998# m3_34996_13126# 0.15fF
C2991 a_2966_8154# m3_1864_8106# 0.14fF
C2992 a_7894_15182# VDD 0.23fF
C2993 a_1962_5182# col_n[19] 0.13fF
C2994 a_1962_11206# a_22346_11206# 0.14fF
C2995 a_30074_12170# a_30074_11166# 1.00fF
C2996 a_2346_11208# a_24050_11166# 0.19fF
C2997 a_10998_11166# col[8] 0.29fF
C2998 a_33086_12170# row_n[10] 0.17fF
C2999 a_31382_17230# vcm 0.22fF
C3000 a_1962_12210# col[12] 0.11fF
C3001 a_13006_11166# ctop 3.58fF
C3002 a_29070_17190# m2_29268_17438# 0.16fF
C3003 a_29070_7150# col[26] 0.29fF
C3004 a_19942_13174# a_20034_13174# 0.26fF
C3005 a_31078_5142# m2_31276_5390# 0.16fF
C3006 a_30986_4138# VDD 0.23fF
C3007 a_2346_5184# a_13918_5142# 0.35fF
C3008 col[31] rowoff_n[13] 0.11fF
C3009 a_26058_15182# ctop 3.58fF
C3010 a_21038_10162# rowon_n[8] 0.14fF
C3011 a_10998_9158# rowoff_n[7] 0.10fF
C3012 a_15014_15182# rowoff_n[13] 0.10fF
C3013 a_6982_14178# vcm 0.62fF
C3014 a_10998_13174# col_n[8] 0.28fF
C3015 a_2346_7192# m2_1732_6970# 0.12fF
C3016 a_1962_2170# a_7986_2130# 0.27fF
C3017 m2_24824_18014# m3_23952_18146# 0.13fF
C3018 m2_1732_17010# m3_1864_18146# 0.15fF
C3019 a_9994_7150# VDD 0.52fF
C3020 a_21038_7150# rowoff_n[5] 0.10fF
C3021 a_2346_7192# a_26970_7150# 0.35fF
C3022 a_14010_7150# a_15014_7150# 0.97fF
C3023 a_1962_1166# col_n[10] 0.13fF
C3024 a_1962_14218# col_n[12] 0.13fF
C3025 a_16018_17190# a_16018_16186# 1.00fF
C3026 a_32994_17190# a_33086_17190# 0.26fF
C3027 a_29070_9158# col_n[26] 0.28fF
C3028 a_31078_5142# rowoff_n[3] 0.10fF
C3029 a_2966_11166# col_n[0] 0.28fF
C3030 a_20034_18194# vcm 0.12fF
C3031 col[15] rowoff_n[14] 0.11fF
C3032 a_1962_8194# col[3] 0.11fF
C3033 a_1962_4178# a_21038_4138# 0.27fF
C3034 a_23046_11166# VDD 0.52fF
C3035 m3_13912_1078# m3_14916_1078# 0.22fF
C3036 a_30074_3134# vcm 0.62fF
C3037 a_2346_7192# col[23] 0.15fF
C3038 a_13310_12210# vcm 0.22fF
C3039 a_1962_1166# a_14314_1166# 0.14fF
C3040 a_28066_6146# m2_28264_6394# 0.16fF
C3041 m2_34864_10986# m3_34996_10114# 0.15fF
C3042 a_18026_13174# row_n[11] 0.17fF
C3043 a_1962_6186# a_34090_6146# 0.27fF
C3044 a_2346_14220# VDD 32.63fF
C3045 a_27062_11166# a_28066_11166# 0.97fF
C3046 a_33086_3134# row_n[1] 0.17fF
C3047 a_24050_17190# m3_23952_18146# 0.15fF
C3048 a_12002_2130# col_n[9] 0.28fF
C3049 a_2874_15182# a_2966_15182# 0.26fF
C3050 a_2346_15224# a_3878_15182# 0.35fF
C3051 a_1962_3174# col[30] 0.11fF
C3052 col_n[5] col_n[6] 0.10fF
C3053 vcm col_n[11] 2.80fF
C3054 VDD col_n[15] 4.67fF
C3055 col[15] col[16] 0.20fF
C3056 a_8990_16186# col[6] 0.29fF
C3057 a_26362_16226# vcm 0.22fF
C3058 a_2346_16228# rowoff_n[14] 4.09fF
C3059 m2_11772_946# m2_12776_946# 0.96fF
C3060 a_15926_3134# a_16018_3134# 0.26fF
C3061 a_2346_3176# a_29070_3134# 0.19fF
C3062 a_1962_3174# a_27366_3174# 0.14fF
C3063 a_7986_10162# ctop 3.58fF
C3064 a_1962_10202# col_n[3] 0.13fF
C3065 a_15926_18194# VDD 0.33fF
C3066 m2_6752_18014# vcm 0.28fF
C3067 a_27062_12170# col[24] 0.29fF
C3068 a_5978_11166# rowon_n[9] 0.14fF
C3069 a_29982_11166# rowoff_n[9] 0.24fF
C3070 a_1962_4178# ctop 1.49fF
C3071 a_25966_3134# VDD 0.23fF
C3072 m3_34996_13126# ctop 0.23fF
C3073 a_21038_14178# ctop 3.58fF
C3074 m2_28840_946# m2_29844_946# 0.96fF
C3075 a_2346_14220# a_11910_14178# 0.35fF
C3076 a_2346_3176# col[14] 0.15fF
C3077 a_2346_16228# col[16] 0.15fF
C3078 a_2346_18236# a_20946_18194# 0.35fF
C3079 a_34394_14218# vcm 0.22fF
C3080 a_25054_7150# m2_25252_7398# 0.16fF
C3081 a_4974_6146# VDD 0.52fF
C3082 a_1962_5182# col_n[30] 0.13fF
C3083 a_12002_7150# a_12002_6146# 1.00fF
C3084 a_28978_7150# a_29070_7150# 0.26fF
C3085 a_1962_11206# a_5978_11166# 0.27fF
C3086 a_25054_14178# rowon_n[12] 0.14fF
C3087 a_9994_5142# col[7] 0.29fF
C3088 m2_29844_946# col_n[27] 0.43fF
C3089 a_13006_16186# a_14010_16186# 0.97fF
C3090 a_2346_16228# a_24962_16186# 0.35fF
C3091 a_1962_12210# col[23] 0.11fF
C3092 a_15014_17190# vcm 0.60fF
C3093 a_27062_14178# col_n[24] 0.28fF
C3094 a_1962_18234# m2_12776_18014# 0.18fF
C3095 a_18026_10162# VDD 0.52fF
C3096 a_25054_2130# vcm 0.62fF
C3097 a_1962_13214# a_19030_13174# 0.27fF
C3098 a_18026_4138# row_n[2] 0.17fF
C3099 a_3970_4138# rowoff_n[2] 0.10fF
C3100 a_8290_11206# vcm 0.22fF
C3101 a_17022_12170# rowoff_n[10] 0.10fF
C3102 m2_34864_7974# m3_34996_7102# 0.15fF
C3103 a_31078_14178# VDD 0.52fF
C3104 a_2346_18236# m2_7756_18014# 0.19fF
C3105 m2_1732_1950# vcm 0.45fF
C3106 a_25054_11166# a_25054_10162# 1.00fF
C3107 a_1962_10202# a_12306_10202# 0.14fF
C3108 a_2346_10204# a_14010_10162# 0.19fF
C3109 a_2966_10162# rowon_n[8] 0.13fF
C3110 a_14010_2130# rowoff_n[0] 0.10fF
C3111 a_1962_15222# a_32082_15182# 0.27fF
C3112 a_2346_12212# col[7] 0.15fF
C3113 a_9994_7150# col_n[7] 0.28fF
C3114 a_31078_16186# rowoff_n[14] 0.10fF
C3115 a_21342_15222# vcm 0.22fF
C3116 a_22042_8154# m2_22240_8402# 0.16fF
C3117 a_1962_1166# col_n[21] 0.13fF
C3118 a_22042_17190# row_n[15] 0.17fF
C3119 a_2966_7150# rowoff_n[5] 0.10fF
C3120 a_1962_14218# col_n[23] 0.13fF
C3121 a_5978_2130# rowon_n[0] 0.14fF
C3122 a_10906_17190# VDD 0.24fF
C3123 a_14922_12170# a_15014_12170# 0.26fF
C3124 a_2346_12212# a_27062_12170# 0.19fF
C3125 a_1962_12210# a_25358_12210# 0.14fF
C3126 m2_20808_946# m3_21944_1078# 0.13fF
C3127 a_28066_3134# col_n[25] 0.28fF
C3128 col[26] rowoff_n[14] 0.11fF
C3129 a_1962_8194# col[14] 0.11fF
C3130 m2_34864_17010# m2_35292_17438# 0.16fF
C3131 a_20946_2130# VDD 0.23fF
C3132 a_25054_17190# col[22] 0.29fF
C3133 a_1962_4178# a_2966_4138# 0.27fF
C3134 a_16018_13174# ctop 3.58fF
C3135 m3_34996_13126# m3_34996_12122# 0.22fF
C3136 m2_31852_946# m3_30980_1078# 0.13fF
C3137 a_15926_18194# m2_15788_18014# 0.16fF
C3138 a_2346_10204# rowoff_n[8] 4.09fF
C3139 a_9994_15182# rowon_n[13] 0.14fF
C3140 a_4882_13174# rowoff_n[11] 0.24fF
C3141 a_33998_6146# VDD 0.23fF
C3142 a_25054_5142# rowon_n[3] 0.14fF
C3143 a_2346_6188# a_16930_6146# 0.35fF
C3144 a_8990_6146# a_9994_6146# 0.97fF
C3145 a_29070_17190# ctop 3.39fF
C3146 a_12914_8154# rowoff_n[6] 0.24fF
C3147 a_2966_17190# m3_1864_17142# 0.14fF
C3148 VDD col_n[26] 4.96fF
C3149 vcm col_n[22] 2.80fF
C3150 col[10] rowoff_n[15] 0.11fF
C3151 a_27974_16186# a_28066_16186# 0.26fF
C3152 a_10998_16186# a_10998_15182# 1.00fF
C3153 a_34090_2130# m2_34864_1950# 0.96fF
C3154 a_7986_10162# col[5] 0.29fF
C3155 a_18938_17190# rowoff_n[15] 0.24fF
C3156 a_9994_16186# vcm 0.62fF
C3157 a_22954_6146# rowoff_n[4] 0.24fF
C3158 a_1962_3174# a_10998_3134# 0.27fF
C3159 a_19030_9158# m2_19228_9406# 0.16fF
C3160 a_1962_10202# col_n[14] 0.13fF
C3161 a_13006_9158# VDD 0.52fF
C3162 a_2346_8196# a_29982_8154# 0.35fF
C3163 a_20034_1126# vcm 0.59fF
C3164 m2_34864_1950# m2_35292_2378# 0.16fF
C3165 a_26058_6146# col[23] 0.29fF
C3166 a_1962_4178# col[5] 0.11fF
C3167 a_3270_10202# vcm 0.22fF
C3168 a_32994_4138# rowoff_n[2] 0.24fF
C3169 a_1962_17230# col[7] 0.11fF
C3170 m2_34864_4962# m3_34996_4090# 0.15fF
C3171 a_1962_5182# a_24050_5142# 0.27fF
C3172 a_2966_14178# ctop 3.42fF
C3173 a_26058_13174# VDD 0.52fF
C3174 a_2346_3176# col[25] 0.15fF
C3175 a_22042_10162# a_23046_10162# 0.97fF
C3176 a_2346_16228# col[27] 0.15fF
C3177 a_33086_5142# vcm 0.62fF
C3178 a_22042_8154# row_n[6] 0.17fF
C3179 a_16322_14218# vcm 0.22fF
C3180 a_10906_2130# a_10998_2130# 0.26fF
C3181 a_2346_2172# a_19030_2130# 0.19fF
C3182 a_1962_2170# a_17326_2170# 0.14fF
C3183 a_7986_12170# col_n[5] 0.28fF
C3184 a_5886_16186# VDD 0.23fF
C3185 a_29374_18234# vcm 0.22fF
C3186 a_15926_1126# VDD 0.44fF
C3187 a_26058_8154# col_n[23] 0.28fF
C3188 a_16018_10162# m2_16216_10410# 0.16fF
C3189 a_2346_4180# a_32082_4138# 0.19fF
C3190 a_34090_5142# a_34090_4138# 1.00fF
C3191 a_1962_6186# col_n[5] 0.13fF
C3192 a_1962_4178# a_30378_4178# 0.14fF
C3193 a_10998_12170# ctop 3.58fF
C3194 a_35002_18194# m2_34864_18014# 0.16fF
C3195 a_9994_6146# rowon_n[4] 0.14fF
C3196 a_31078_10162# rowoff_n[8] 0.10fF
C3197 a_33086_13174# rowoff_n[11] 0.10fF
C3198 a_28978_5142# VDD 0.23fF
C3199 m3_13912_18146# VDD 0.25fF
C3200 a_6982_6146# a_6982_5142# 1.00fF
C3201 a_23958_6146# a_24050_6146# 0.26fF
C3202 a_24050_16186# ctop 3.57fF
C3203 a_2346_12212# col[18] 0.15fF
C3204 a_2346_15224# a_14922_15182# 0.35fF
C3205 a_7986_15182# a_8990_15182# 0.97fF
C3206 a_4974_15182# vcm 0.62fF
C3207 a_29070_9158# rowon_n[7] 0.14fF
C3208 a_7986_8154# VDD 0.52fF
C3209 a_5978_15182# col[3] 0.29fF
C3210 a_1962_8194# col[25] 0.11fF
C3211 a_1962_12210# a_8990_12170# 0.27fF
C3212 a_1962_18234# a_32386_18234# 0.14fF
C3213 a_2346_17232# a_27974_17190# 0.35fF
C3214 m2_34864_1950# m3_34996_2082# 2.76fF
C3215 m2_1732_946# m3_1864_2082# 0.15fF
C3216 a_24050_11166# col[21] 0.29fF
C3217 a_1962_2170# VDD 2.76fF
C3218 m3_20940_1078# ctop 0.23fF
C3219 a_6982_9158# row_n[7] 0.17fF
C3220 a_1962_15222# sample 0.14fF
C3221 a_13006_11166# m2_13204_11414# 0.16fF
C3222 a_21038_12170# VDD 0.52fF
C3223 m3_9896_18146# m3_10900_18146# 0.22fF
C3224 a_2346_9200# a_3970_9158# 0.19fF
C3225 a_20034_10162# a_20034_9158# 1.00fF
C3226 a_28066_4138# vcm 0.62fF
C3227 a_1962_14218# a_22042_14178# 0.27fF
C3228 a_5886_3134# rowoff_n[1] 0.24fF
C3229 a_11302_13214# vcm 0.22fF
C3230 a_20946_14178# rowoff_n[12] 0.24fF
C3231 VDD row_n[13] 2.93fF
C3232 vcm row_n[15] 0.49fF
C3233 sample row_n[14] 1.03fF
C3234 a_2346_8196# col[9] 0.15fF
C3235 col[21] rowoff_n[15] 0.11fF
C3236 a_34090_16186# VDD 0.54fF
C3237 col[26] col[27] 0.20fF
C3238 a_2346_11208# a_17022_11166# 0.19fF
C3239 a_1962_11206# a_15318_11206# 0.14fF
C3240 a_9902_11166# a_9994_11166# 0.26fF
C3241 a_5978_17190# col_n[3] 0.28fF
C3242 a_6982_4138# col[4] 0.29fF
C3243 a_20034_2130# m2_20232_2378# 0.16fF
C3244 a_26058_12170# row_n[10] 0.17fF
C3245 a_1962_10202# col_n[25] 0.13fF
C3246 a_24354_17230# vcm 0.22fF
C3247 a_31078_4138# a_32082_4138# 0.97fF
C3248 a_5978_11166# ctop 3.58fF
C3249 a_24050_13174# col_n[21] 0.28fF
C3250 a_1962_4178# col[16] 0.11fF
C3251 a_1962_17230# col[18] 0.11fF
C3252 a_35398_2170# vcm 0.23fF
C3253 a_1962_13214# a_28370_13214# 0.14fF
C3254 a_33086_14178# a_33086_13174# 1.00fF
C3255 a_2346_13216# a_30074_13174# 0.19fF
C3256 m2_10768_18014# col_n[8] 0.25fF
C3257 a_23958_4138# VDD 0.23fF
C3258 a_3970_5142# a_4974_5142# 0.97fF
C3259 a_2346_5184# a_6890_5142# 0.35fF
C3260 a_9994_12170# m2_10192_12418# 0.16fF
C3261 a_19030_15182# ctop 3.58fF
C3262 a_14010_10162# rowon_n[8] 0.14fF
C3263 a_3970_9158# rowoff_n[7] 0.10fF
C3264 a_5978_15182# a_5978_14178# 1.00fF
C3265 a_22954_15182# a_23046_15182# 0.26fF
C3266 a_7986_15182# rowoff_n[13] 0.10fF
C3267 m2_14784_18014# m3_15920_18146# 0.13fF
C3268 a_2874_7150# VDD 0.24fF
C3269 a_6982_6146# col_n[4] 0.28fF
C3270 a_14010_7150# rowoff_n[5] 0.10fF
C3271 a_2346_7192# a_19942_7150# 0.35fF
C3272 a_2346_4180# col[0] 0.15fF
C3273 a_2346_17232# col[2] 0.15fF
C3274 a_1962_6186# col_n[16] 0.13fF
C3275 a_24050_5142# rowoff_n[3] 0.10fF
C3276 a_13006_18194# vcm 0.12fF
C3277 a_25054_2130# col_n[22] 0.28fF
C3278 a_1962_4178# a_14010_4138# 0.27fF
C3279 a_33086_13174# rowon_n[11] 0.14fF
C3280 a_16018_11166# VDD 0.52fF
C3281 m3_1864_2082# m3_1864_1078# 0.22fF
C3282 a_17022_9158# a_18026_9158# 0.97fF
C3283 a_2346_9200# a_32994_9158# 0.35fF
C3284 a_22042_16186# col[19] 0.29fF
C3285 a_1962_13214# col[9] 0.11fF
C3286 a_23046_3134# vcm 0.62fF
C3287 a_34090_3134# rowoff_n[1] 0.10fF
C3288 rowon_n[8] rowoff_n[8] 20.27fF
C3289 a_6282_12210# vcm 0.22fF
C3290 a_1962_1166# a_7286_1166# 0.14fF
C3291 a_10998_13174# row_n[11] 0.17fF
C3292 a_2346_12212# col[29] 0.15fF
C3293 a_1962_6186# a_27062_6146# 0.27fF
C3294 a_6982_13174# m2_7180_13422# 0.16fF
C3295 a_29070_15182# VDD 0.52fF
C3296 m2_11772_946# a_2346_1168# 0.19fF
C3297 a_26058_3134# row_n[1] 0.17fF
C3298 a_2346_6188# vcm 0.40fF
C3299 a_19334_16226# vcm 0.22fF
C3300 a_29070_4138# a_29070_3134# 1.00fF
C3301 a_2346_3176# a_22042_3134# 0.19fF
C3302 a_1962_3174# a_20338_3174# 0.14fF
C3303 a_13006_2130# m3_12908_1078# 0.15fF
C3304 a_2346_1168# m2_28840_946# 0.19fF
C3305 a_4974_9158# col[2] 0.29fF
C3306 a_8898_18194# VDD 0.33fF
C3307 a_30074_13174# a_31078_13174# 0.97fF
C3308 a_29374_1166# vcm 0.23fF
C3309 a_22954_11166# rowoff_n[9] 0.24fF
C3310 a_1962_2170# col_n[7] 0.13fF
C3311 a_1962_15222# col_n[9] 0.13fF
C3312 a_30074_16186# row_n[14] 0.17fF
C3313 a_23046_5142# col[20] 0.29fF
C3314 a_18938_3134# VDD 0.23fF
C3315 m3_16924_18146# ctop 0.23fF
C3316 a_1962_5182# a_33390_5182# 0.14fF
C3317 a_18938_5142# a_19030_5142# 0.26fF
C3318 a_14010_14178# ctop 3.58fF
C3319 a_2966_12170# VDD 0.56fF
C3320 a_1962_9198# col[0] 0.11fF
C3321 a_32994_9158# rowoff_n[7] 0.24fF
C3322 a_2346_14220# a_4882_14178# 0.35fF
C3323 a_2346_18236# a_13918_18194# 0.35fF
C3324 vcm rowon_n[9] 0.50fF
C3325 col_n[11] row_n[15] 0.23fF
C3326 col_n[0] row_n[9] 0.23fF
C3327 col_n[3] row_n[11] 0.23fF
C3328 col_n[5] row_n[12] 0.23fF
C3329 VDD rowon_n[7] 2.61fF
C3330 col_n[7] row_n[13] 0.23fF
C3331 col_n[1] row_n[10] 0.23fF
C3332 col_n[9] row_n[14] 0.23fF
C3333 a_2346_8196# col[20] 0.15fF
C3334 a_31990_7150# VDD 0.23fF
C3335 a_3970_14178# m2_4168_14426# 0.16fF
C3336 a_18026_14178# rowon_n[12] 0.14fF
C3337 a_4974_11166# col_n[2] 0.28fF
C3338 a_2346_16228# a_17934_16186# 0.35fF
C3339 a_33086_4138# rowon_n[2] 0.14fF
C3340 a_7986_17190# vcm 0.60fF
C3341 a_1962_4178# col[27] 0.11fF
C3342 a_10998_10162# VDD 0.52fF
C3343 a_1962_17230# col[29] 0.11fF
C3344 a_31990_9158# a_32082_9158# 0.26fF
C3345 a_1962_17230# m2_34864_17010# 0.17fF
C3346 a_15014_9158# a_15014_8154# 1.00fF
C3347 a_23046_7150# col_n[20] 0.28fF
C3348 a_18026_2130# vcm 0.62fF
C3349 a_1962_13214# a_12002_13174# 0.27fF
C3350 m2_1732_2954# m2_2160_3382# 0.16fF
C3351 a_10998_4138# row_n[2] 0.17fF
C3352 a_9994_12170# rowoff_n[10] 0.10fF
C3353 a_1962_11206# vcm 6.95fF
C3354 m3_34996_7102# VDD 0.26fF
C3355 a_24050_14178# VDD 0.52fF
C3356 a_2346_10204# a_6982_10162# 0.19fF
C3357 a_1962_10202# a_5278_10202# 0.14fF
C3358 a_4882_10162# a_4974_10162# 0.26fF
C3359 a_6982_2130# rowoff_n[0] 0.10fF
C3360 a_31078_6146# vcm 0.62fF
C3361 a_1962_15222# a_25054_15182# 0.27fF
C3362 m2_20808_18014# ctop 0.18fF
C3363 a_14314_15222# vcm 0.22fF
C3364 a_24050_16186# rowoff_n[14] 0.10fF
C3365 a_26058_3134# a_27062_3134# 0.97fF
C3366 a_2346_4180# col[11] 0.15fF
C3367 a_2346_17232# col[13] 0.15fF
C3368 a_15014_17190# row_n[15] 0.17fF
C3369 a_34090_11166# m3_34996_11118# 0.13fF
C3370 a_28066_13174# a_28066_12170# 1.00fF
C3371 a_1962_12210# a_18330_12210# 0.14fF
C3372 a_2346_12212# a_20034_12170# 0.19fF
C3373 a_30074_7150# row_n[5] 0.17fF
C3374 a_1962_6186# col_n[27] 0.13fF
C3375 a_13918_2130# VDD 0.23fF
C3376 a_1962_13214# col[20] 0.11fF
C3377 a_8990_13174# ctop 3.58fF
C3378 a_21038_10162# col[18] 0.29fF
C3379 a_1962_14218# a_31382_14218# 0.14fF
C3380 a_17934_14178# a_18026_14178# 0.26fF
C3381 a_2346_14220# a_33086_14178# 0.19fF
C3382 m2_34864_6970# m2_34864_5966# 0.99fF
C3383 a_26970_6146# VDD 0.23fF
C3384 a_18026_5142# rowon_n[3] 0.14fF
C3385 a_2346_6188# a_9902_6146# 0.35fF
C3386 a_22042_17190# ctop 3.39fF
C3387 a_5886_8154# rowoff_n[6] 0.24fF
C3388 a_32082_2130# ctop 3.39fF
C3389 a_11910_17190# rowoff_n[15] 0.24fF
C3390 a_2346_13216# col[4] 0.15fF
C3391 a_15926_6146# rowoff_n[4] 0.24fF
C3392 a_1962_3174# a_3970_3134# 0.27fF
C3393 a_3970_3134# col[1] 0.29fF
C3394 a_5978_9158# VDD 0.52fF
C3395 rowon_n[10] rowoff_n[10] 20.27fF
C3396 a_12002_8154# a_13006_8154# 0.97fF
C3397 a_32082_17190# m2_32280_17438# 0.16fF
C3398 a_2346_8196# a_22954_8154# 0.35fF
C3399 a_1962_2170# col_n[18] 0.13fF
C3400 a_13006_1126# vcm 0.12fF
C3401 a_1962_15222# col_n[20] 0.13fF
C3402 a_21038_12170# col_n[18] 0.28fF
C3403 a_25966_4138# rowoff_n[2] 0.24fF
C3404 a_34090_5142# m2_34288_5390# 0.16fF
C3405 a_1962_5182# a_17022_5142# 0.27fF
C3406 a_1962_9198# col[11] 0.11fF
C3407 a_19030_13174# VDD 0.52fF
C3408 m2_25828_18014# col[23] 0.28fF
C3409 a_26058_5142# vcm 0.62fF
C3410 VDD row_n[2] 2.93fF
C3411 vcm row_n[4] 0.49fF
C3412 col_n[18] row_n[13] 0.23fF
C3413 sample row_n[3] 1.03fF
C3414 col_n[12] row_n[10] 0.23fF
C3415 col_n[4] row_n[6] 0.23fF
C3416 col_n[14] row_n[11] 0.23fF
C3417 col_n[22] row_n[15] 0.23fF
C3418 col_n[10] row_n[9] 0.23fF
C3419 col_n[27] col_n[28] 0.10fF
C3420 col_n[6] row_n[7] 0.23fF
C3421 col_n[20] row_n[14] 0.23fF
C3422 col_n[8] row_n[8] 0.23fF
C3423 col_n[2] row_n[5] 0.23fF
C3424 col_n[16] row_n[12] 0.23fF
C3425 a_2346_8196# col[31] 0.15fF
C3426 a_15014_8154# row_n[6] 0.17fF
C3427 a_9294_14218# vcm 0.22fF
C3428 a_24050_3134# a_24050_2130# 1.00fF
C3429 a_2346_2172# a_12002_2130# 0.19fF
C3430 a_1962_2170# a_10298_2170# 0.14fF
C3431 m2_29844_18014# m3_28972_18146# 0.13fF
C3432 a_1962_7190# a_30074_7150# 0.27fF
C3433 a_1962_10202# row_n[8] 25.57fF
C3434 a_32082_17190# VDD 0.55fF
C3435 a_25054_12170# a_26058_12170# 0.97fF
C3436 m2_34864_13998# vcm 0.51fF
C3437 a_3970_5142# col_n[1] 0.28fF
C3438 a_22346_18234# vcm 0.22fF
C3439 a_8898_1126# VDD 0.44fF
C3440 a_1962_4178# a_23350_4178# 0.14fF
C3441 a_13918_4138# a_14010_4138# 0.26fF
C3442 a_2346_4180# a_25054_4138# 0.19fF
C3443 a_3970_12170# ctop 3.57fF
C3444 a_1962_11206# col_n[11] 0.13fF
C3445 a_34090_11166# row_n[9] 0.17fF
C3446 a_32386_3174# vcm 0.22fF
C3447 a_24050_10162# rowoff_n[8] 0.10fF
C3448 a_19030_15182# col[16] 0.29fF
C3449 a_26058_13174# rowoff_n[11] 0.10fF
C3450 a_31078_6146# m2_31276_6394# 0.16fF
C3451 a_21950_5142# VDD 0.23fF
C3452 a_1962_5182# col[2] 0.11fF
C3453 m2_27836_946# VDD 0.62fF
C3454 a_17022_16186# ctop 3.57fF
C3455 a_34090_8154# rowoff_n[6] 0.10fF
C3456 a_27062_17190# m3_26964_18146# 0.15fF
C3457 a_2346_15224# a_7894_15182# 0.35fF
C3458 a_2346_4180# col[22] 0.15fF
C3459 a_2346_17232# col[24] 0.15fF
C3460 m2_15788_946# m2_16216_1374# 0.16fF
C3461 a_2346_8196# m2_1732_7974# 0.12fF
C3462 a_22042_9158# rowon_n[7] 0.14fF
C3463 a_35002_9158# VDD 0.29fF
C3464 a_9994_8154# a_9994_7150# 1.00fF
C3465 a_26970_8154# a_27062_8154# 0.26fF
C3466 a_1962_18234# a_25358_18234# 0.14fF
C3467 m2_1732_4962# sample 0.19fF
C3468 a_2346_17232# a_20946_17190# 0.35fF
C3469 a_10998_17190# a_12002_17190# 0.97fF
C3470 m2_1732_16006# sample_n 0.15fF
C3471 m2_27836_18014# m2_28840_18014# 0.96fF
C3472 a_1962_13214# col[31] 0.11fF
C3473 a_19030_17190# col_n[16] 0.28fF
C3474 m3_1864_5094# ctop 0.23fF
C3475 ctop rowoff_n[6] 0.60fF
C3476 a_14010_12170# VDD 0.52fF
C3477 m2_32856_946# m2_33284_1374# 0.16fF
C3478 a_20034_4138# col[17] 0.29fF
C3479 a_1962_7190# col_n[2] 0.13fF
C3480 a_21038_4138# vcm 0.62fF
C3481 a_1962_14218# a_15014_14178# 0.27fF
C3482 a_13918_14178# rowoff_n[12] 0.24fF
C3483 a_4274_13214# vcm 0.22fF
C3484 a_21038_2130# a_22042_2130# 0.97fF
C3485 a_28066_7150# m2_28264_7398# 0.16fF
C3486 a_27062_16186# VDD 0.52fF
C3487 a_1962_11206# a_8290_11206# 0.14fF
C3488 a_2346_11208# a_9994_11166# 0.19fF
C3489 a_23046_12170# a_23046_11166# 1.00fF
C3490 a_34090_8154# vcm 0.62fF
C3491 a_1962_16226# a_28066_16186# 0.27fF
C3492 a_2346_13216# col[15] 0.15fF
C3493 a_19030_12170# row_n[10] 0.17fF
C3494 a_17326_17230# vcm 0.22fF
C3495 a_1962_2170# col_n[29] 0.13fF
C3496 a_34090_2130# row_n[0] 0.17fF
C3497 a_2966_8154# a_3970_8154# 0.97fF
C3498 a_1962_15222# col_n[31] 0.13fF
C3499 a_2346_13216# a_23046_13174# 0.19fF
C3500 a_1962_13214# a_21342_13214# 0.14fF
C3501 a_27366_2170# vcm 0.22fF
C3502 a_12914_13174# a_13006_13174# 0.26fF
C3503 a_20034_6146# col_n[17] 0.28fF
C3504 a_1962_9198# col[22] 0.11fF
C3505 a_16930_4138# VDD 0.23fF
C3506 m3_32988_1078# VDD 0.14fF
C3507 a_12002_15182# ctop 3.58fF
C3508 a_6982_10162# rowon_n[8] 0.14fF
C3509 col_n[7] row_n[2] 0.23fF
C3510 col_n[3] row_n[0] 0.23fF
C3511 col_n[19] row_n[8] 0.23fF
C3512 VDD en_bit_n[0] 0.15fF
C3513 vcm ctop 33.18fF
C3514 col_n[25] row_n[11] 0.23fF
C3515 col_n[13] row_n[5] 0.23fF
C3516 col_n[17] row_n[7] 0.23fF
C3517 rowon_n[15] rowon_n[14] 0.15fF
C3518 col_n[11] row_n[4] 0.23fF
C3519 col_n[31] row_n[14] 0.23fF
C3520 col_n[23] row_n[10] 0.23fF
C3521 col_n[9] row_n[3] 0.23fF
C3522 col_n[21] row_n[9] 0.23fF
C3523 col_n[29] row_n[13] 0.23fF
C3524 col_n[27] row_n[12] 0.23fF
C3525 col_n[15] row_n[6] 0.23fF
C3526 col_n[5] row_n[1] 0.23fF
C3527 a_2346_15224# a_2346_14220# 0.22fF
C3528 a_1962_15222# a_35398_15222# 0.14fF
C3529 a_25054_8154# m2_25252_8402# 0.16fF
C3530 m2_5748_18014# m3_5880_18146# 2.78fF
C3531 a_29982_8154# VDD 0.23fF
C3532 a_6982_7150# rowoff_n[5] 0.10fF
C3533 a_6982_7150# a_7986_7150# 0.97fF
C3534 a_2346_7192# a_12914_7150# 0.35fF
C3535 a_2346_9200# col[6] 0.15fF
C3536 a_25966_17190# a_26058_17190# 0.26fF
C3537 a_8990_17190# a_8990_16186# 1.00fF
C3538 a_17022_5142# rowoff_n[3] 0.10fF
C3539 a_5978_18194# vcm 0.12fF
C3540 a_1962_18234# col_n[5] 0.13fF
C3541 a_1962_4178# a_6982_4138# 0.27fF
C3542 a_26058_13174# rowon_n[11] 0.14fF
C3543 a_1962_11206# col_n[22] 0.13fF
C3544 a_8990_11166# VDD 0.52fF
C3545 m2_23820_946# col_n[21] 0.37fF
C3546 a_2346_9200# a_25966_9158# 0.35fF
C3547 a_16018_3134# vcm 0.62fF
C3548 m2_12776_946# col[10] 0.39fF
C3549 a_27062_3134# rowoff_n[1] 0.10fF
C3550 a_18026_9158# col[15] 0.29fF
C3551 a_1962_5182# col[13] 0.11fF
C3552 a_19030_2130# a_19030_1126# 1.00fF
C3553 a_3970_13174# row_n[11] 0.17fF
C3554 a_3878_5142# VDD 0.23fF
C3555 a_1962_6186# a_20034_6146# 0.27fF
C3556 a_22042_15182# VDD 0.52fF
C3557 a_20034_11166# a_21038_11166# 0.97fF
C3558 a_19030_3134# row_n[1] 0.17fF
C3559 a_29070_7150# vcm 0.62fF
C3560 a_2346_1168# m2_4744_946# 0.19fF
C3561 a_12306_16226# vcm 0.22fF
C3562 a_22042_9158# m2_22240_9406# 0.16fF
C3563 a_2346_3176# a_15014_3134# 0.19fF
C3564 a_1962_3174# a_13310_3174# 0.14fF
C3565 a_8898_3134# a_8990_3134# 0.26fF
C3566 a_29070_2130# m2_28840_946# 0.99fF
C3567 a_1962_8194# a_33086_8154# 0.27fF
C3568 a_22346_1166# vcm 0.23fF
C3569 m2_4744_946# m2_5748_946# 0.96fF
C3570 a_2346_17232# a_1962_17230# 2.62fF
C3571 a_15926_11166# rowoff_n[9] 0.24fF
C3572 col[0] rowoff_n[1] 0.11fF
C3573 col[1] rowoff_n[2] 0.11fF
C3574 col[6] rowoff_n[7] 0.11fF
C3575 col[8] rowoff_n[9] 0.11fF
C3576 col[7] rowoff_n[8] 0.11fF
C3577 col[5] rowoff_n[6] 0.11fF
C3578 col[2] rowoff_n[3] 0.11fF
C3579 col[3] rowoff_n[4] 0.11fF
C3580 col[4] rowoff_n[5] 0.11fF
C3581 a_23046_16186# row_n[14] 0.17fF
C3582 a_11910_3134# VDD 0.23fF
C3583 a_18026_11166# col_n[15] 0.28fF
C3584 a_1962_5182# a_26362_5182# 0.14fF
C3585 a_32082_6146# a_32082_5142# 1.00fF
C3586 a_2346_5184# a_28066_5142# 0.19fF
C3587 a_1962_7190# col_n[13] 0.13fF
C3588 a_6982_14178# ctop 3.58fF
C3589 a_25966_9158# rowoff_n[7] 0.24fF
C3590 a_33086_15182# a_34090_15182# 0.97fF
C3591 a_2966_4138# vcm 0.61fF
C3592 a_1962_1166# col[4] 0.11fF
C3593 a_2346_18236# a_6890_18194# 0.35fF
C3594 a_1962_14218# col[6] 0.11fF
C3595 a_29982_15182# rowoff_n[13] 0.24fF
C3596 a_24962_7150# VDD 0.23fF
C3597 a_4974_7150# a_4974_6146# 1.00fF
C3598 a_21950_7150# a_22042_7150# 0.26fF
C3599 a_10998_14178# rowon_n[12] 0.14fF
C3600 a_2346_13216# col[26] 0.15fF
C3601 a_5978_16186# a_6982_16186# 0.97fF
C3602 a_2346_16228# a_10906_16186# 0.35fF
C3603 a_26058_4138# rowon_n[2] 0.14fF
C3604 a_30074_3134# ctop 3.57fF
C3605 a_19030_10162# m2_19228_10410# 0.16fF
C3606 a_1962_4178# a_34394_4178# 0.14fF
C3607 a_3970_10162# VDD 0.52fF
C3608 a_10998_2130# vcm 0.62fF
C3609 a_3878_13174# a_3970_13174# 0.26fF
C3610 a_1962_13214# a_4974_13174# 0.27fF
C3611 a_3970_4138# row_n[2] 0.17fF
C3612 a_2874_12170# rowoff_n[10] 0.24fF
C3613 a_2346_1168# a_30986_1126# 0.35fF
C3614 a_16018_14178# col[13] 0.29fF
C3615 a_1962_3174# col_n[4] 0.13fF
C3616 m3_28972_18146# VDD 0.24fF
C3617 col_n[14] row_n[0] 0.23fF
C3618 col_n[24] row_n[5] 0.23fF
C3619 col_n[20] row_n[3] 0.23fF
C3620 col_n[28] row_n[7] 0.23fF
C3621 rowon_n[12] row_n[12] 19.75fF
C3622 col_n[30] row_n[8] 0.23fF
C3623 VDD col[9] 4.19fF
C3624 col_n[26] row_n[6] 0.23fF
C3625 vcm col[5] 5.84fF
C3626 col_n[22] row_n[4] 0.23fF
C3627 col_n[2] col[3] 5.98fF
C3628 col_n[16] row_n[1] 0.23fF
C3629 col_n[18] row_n[2] 0.23fF
C3630 col_n[11] ctop 2.02fF
C3631 a_1962_16226# col_n[6] 0.13fF
C3632 a_30074_17190# rowon_n[15] 0.14fF
C3633 a_17022_14178# VDD 0.52fF
C3634 a_18026_11166# a_18026_10162# 1.00fF
C3635 a_24050_6146# vcm 0.62fF
C3636 a_1962_15222# a_18026_15182# 0.27fF
C3637 a_34090_10162# col[31] 0.29fF
C3638 a_17022_16186# rowoff_n[14] 0.10fF
C3639 a_7286_15222# vcm 0.22fF
C3640 m2_6752_18014# ctop 0.18fF
C3641 a_7986_17190# row_n[15] 0.17fF
C3642 a_25966_1126# m2_25828_946# 0.16fF
C3643 a_2346_9200# col[17] 0.15fF
C3644 a_2346_12212# a_13006_12170# 0.19fF
C3645 m2_1732_17010# vcm 0.44fF
C3646 a_7894_12170# a_7986_12170# 0.26fF
C3647 a_1962_12210# a_11302_12210# 0.14fF
C3648 a_23046_7150# row_n[5] 0.17fF
C3649 a_1962_17230# a_31078_17190# 0.27fF
C3650 a_1962_18234# col_n[16] 0.13fF
C3651 m2_5748_946# m3_6884_1078# 0.13fF
C3652 a_6890_2130# VDD 0.23fF
C3653 a_29070_5142# a_30074_5142# 0.97fF
C3654 a_16018_11166# m2_16216_11414# 0.16fF
C3655 a_16018_16186# col_n[13] 0.28fF
C3656 a_1962_5182# col[24] 0.11fF
C3657 a_30378_4178# vcm 0.22fF
C3658 a_2346_14220# a_26058_14178# 0.19fF
C3659 a_31078_15182# a_31078_14178# 1.00fF
C3660 a_1962_14218# a_24354_14218# 0.14fF
C3661 a_17022_3134# col[14] 0.29fF
C3662 m2_34864_4962# VDD 1.01fF
C3663 a_19942_6146# VDD 0.23fF
C3664 a_10998_5142# rowon_n[3] 0.14fF
C3665 a_34090_12170# col_n[31] 0.28fF
C3666 a_15014_17190# ctop 3.39fF
C3667 a_3970_16186# a_3970_15182# 1.00fF
C3668 a_20946_16186# a_21038_16186# 0.26fF
C3669 m2_34864_12994# row_n[11] 0.15fF
C3670 a_23046_2130# m2_23244_2378# 0.16fF
C3671 a_25054_2130# ctop 3.39fF
C3672 a_4882_17190# rowoff_n[15] 0.24fF
C3673 m2_26832_18014# VDD 1.32fF
C3674 a_8898_6146# rowoff_n[4] 0.24fF
C3675 a_32994_10162# VDD 0.23fF
C3676 a_2346_8196# a_15926_8154# 0.35fF
C3677 a_2346_5184# col[8] 0.15fF
C3678 a_5978_1126# vcm 0.12fF
C3679 col[18] rowoff_n[8] 0.11fF
C3680 col[17] rowoff_n[7] 0.11fF
C3681 col[19] rowoff_n[9] 0.11fF
C3682 col[12] rowoff_n[2] 0.11fF
C3683 col[11] rowoff_n[1] 0.11fF
C3684 col[10] rowoff_n[0] 0.11fF
C3685 col[15] rowoff_n[5] 0.11fF
C3686 col[16] rowoff_n[6] 0.11fF
C3687 col[13] rowoff_n[3] 0.11fF
C3688 col[14] rowoff_n[4] 0.11fF
C3689 a_31990_12170# rowoff_n[10] 0.24fF
C3690 a_18938_4138# rowoff_n[2] 0.24fF
C3691 a_30074_8154# rowon_n[6] 0.14fF
C3692 a_1962_7190# col_n[24] 0.13fF
C3693 a_17022_5142# col_n[14] 0.28fF
C3694 a_1962_5182# a_9994_5142# 0.27fF
C3695 a_13006_12170# m2_13204_12418# 0.16fF
C3696 a_12002_13174# VDD 0.52fF
C3697 a_2346_10204# a_28978_10162# 0.35fF
C3698 a_15014_10162# a_16018_10162# 0.97fF
C3699 a_28978_2130# rowoff_n[0] 0.24fF
C3700 a_1962_1166# col[15] 0.11fF
C3701 a_1962_14218# col[17] 0.11fF
C3702 a_19030_5142# vcm 0.62fF
C3703 a_7986_8154# row_n[6] 0.17fF
C3704 a_2346_2172# a_4974_2130# 0.19fF
C3705 a_1962_2170# a_3270_2170# 0.14fF
C3706 vcm rowoff_n[14] 0.20fF
C3707 m2_19804_18014# m3_20940_18146# 0.13fF
C3708 a_32082_15182# col[29] 0.29fF
C3709 a_1962_7190# a_23046_7150# 0.27fF
C3710 a_25054_17190# VDD 0.55fF
C3711 col[3] rowoff_n[10] 0.11fF
C3712 a_32082_9158# vcm 0.62fF
C3713 a_15318_18234# vcm 0.22fF
C3714 a_1962_4178# a_16322_4178# 0.14fF
C3715 a_27062_5142# a_27062_4138# 1.00fF
C3716 a_2346_4180# a_18026_4138# 0.19fF
C3717 a_2346_14220# col[1] 0.15fF
C3718 a_2346_18236# a_2874_18194# 0.35fF
C3719 a_28066_14178# a_29070_14178# 0.97fF
C3720 a_25358_3174# vcm 0.22fF
C3721 a_27062_11166# row_n[9] 0.17fF
C3722 a_17022_10162# rowoff_n[8] 0.10fF
C3723 a_19030_13174# rowoff_n[11] 0.10fF
C3724 a_1962_3174# col_n[15] 0.13fF
C3725 VDD col[20] 4.17fF
C3726 col_n[29] row_n[2] 0.23fF
C3727 col_n[8] col[8] 0.72fF
C3728 vcm col[16] 5.84fF
C3729 col_n[25] row_n[0] 0.23fF
C3730 col_n[27] row_n[1] 0.23fF
C3731 col_n[31] row_n[3] 0.23fF
C3732 col_n[22] ctop 2.02fF
C3733 a_1962_16226# col_n[17] 0.13fF
C3734 a_15014_8154# col[12] 0.29fF
C3735 a_14922_5142# VDD 0.23fF
C3736 a_16930_6146# a_17022_6146# 0.26fF
C3737 a_9994_13174# m2_10192_13422# 0.16fF
C3738 a_1962_6186# a_29374_6186# 0.14fF
C3739 a_2346_6188# a_31078_6146# 0.19fF
C3740 m2_4744_18014# col_n[2] 0.25fF
C3741 a_9994_16186# ctop 3.57fF
C3742 a_27062_8154# rowoff_n[6] 0.10fF
C3743 m2_20808_946# a_2346_1168# 0.19fF
C3744 a_1962_10202# col[8] 0.11fF
C3745 a_32082_17190# col_n[29] 0.28fF
C3746 a_2346_15224# row_n[13] 0.35fF
C3747 a_33086_4138# col[30] 0.29fF
C3748 a_20034_1126# ctop 0.65fF
C3749 a_33086_17190# rowoff_n[15] 0.10fF
C3750 a_16018_2130# m3_15920_1078# 0.15fF
C3751 a_2346_9200# col[28] 0.15fF
C3752 a_15014_9158# rowon_n[7] 0.14fF
C3753 a_27974_9158# VDD 0.23fF
C3754 a_33390_1166# vcm 0.22fF
C3755 a_1962_18234# a_18330_18234# 0.14fF
C3756 a_1962_18234# col_n[27] 0.13fF
C3757 a_1962_11206# rowon_n[9] 1.18fF
C3758 a_2346_17232# a_13918_17190# 0.35fF
C3759 m2_20808_18014# m2_21812_18014# 0.96fF
C3760 a_33086_5142# ctop 3.57fF
C3761 m3_31984_18146# ctop 0.23fF
C3762 a_6982_12170# VDD 0.52fF
C3763 m2_25828_946# m2_26256_1374# 0.16fF
C3764 a_15014_10162# col_n[12] 0.28fF
C3765 a_29982_10162# a_30074_10162# 0.26fF
C3766 a_13006_10162# a_13006_9158# 1.00fF
C3767 a_14010_4138# vcm 0.62fF
C3768 a_1962_14218# a_7986_14178# 0.27fF
C3769 a_6890_14178# rowoff_n[12] 0.24fF
C3770 a_1962_12210# col_n[8] 0.13fF
C3771 a_34090_12170# rowon_n[10] 0.14fF
C3772 a_2346_2172# a_33998_2130# 0.35fF
C3773 a_35494_7512# VDD 0.11fF
C3774 a_33086_6146# col_n[30] 0.28fF
C3775 a_6982_14178# m2_7180_14426# 0.16fF
C3776 a_20034_16186# VDD 0.52fF
C3777 a_2346_11208# a_2874_11166# 0.35fF
C3778 a_27062_8154# vcm 0.62fF
C3779 a_1962_16226# a_21038_16186# 0.27fF
C3780 a_12002_12170# row_n[10] 0.17fF
C3781 a_10298_17230# vcm 0.22fF
C3782 a_24050_4138# a_25054_4138# 0.97fF
C3783 a_2346_5184# col[19] 0.15fF
C3784 a_27062_2130# row_n[0] 0.17fF
C3785 a_22042_17190# m2_21812_18014# 1.00fF
C3786 col[27] rowoff_n[6] 0.11fF
C3787 col[21] rowoff_n[0] 0.11fF
C3788 col[28] rowoff_n[7] 0.11fF
C3789 col[30] rowoff_n[9] 0.11fF
C3790 col[22] rowoff_n[1] 0.11fF
C3791 col[29] rowoff_n[8] 0.11fF
C3792 col[23] rowoff_n[2] 0.11fF
C3793 col[24] rowoff_n[3] 0.11fF
C3794 col[25] rowoff_n[4] 0.11fF
C3795 col[26] rowoff_n[5] 0.11fF
C3796 a_20338_2170# vcm 0.22fF
C3797 a_2346_13216# a_16018_13174# 0.19fF
C3798 a_26058_14178# a_26058_13174# 1.00fF
C3799 a_1962_13214# a_14314_13214# 0.14fF
C3800 a_9902_4138# VDD 0.23fF
C3801 m3_4876_1078# VDD 0.14fF
C3802 a_1962_1166# col[26] 0.11fF
C3803 a_4974_15182# ctop 3.58fF
C3804 a_2346_6188# row_n[4] 0.35fF
C3805 a_1962_14218# col[28] 0.11fF
C3806 a_13006_13174# col[10] 0.29fF
C3807 a_31078_15182# row_n[13] 0.17fF
C3808 a_15926_15182# a_16018_15182# 0.26fF
C3809 a_2346_15224# a_29070_15182# 0.19fF
C3810 a_33390_6186# vcm 0.22fF
C3811 a_1962_15222# a_27366_15222# 0.14fF
C3812 m2_1732_9982# m2_1732_8978# 0.99fF
C3813 a_1962_8194# col_n[0] 0.13fF
C3814 col[14] rowoff_n[10] 0.11fF
C3815 a_22954_8154# VDD 0.23fF
C3816 a_31078_9158# col[28] 0.29fF
C3817 a_2346_7192# a_5886_7150# 0.35fF
C3818 a_3970_15182# m2_4168_15430# 0.16fF
C3819 a_1962_2170# rowon_n[0] 1.18fF
C3820 m2_15788_946# m3_15920_1078# 2.79fF
C3821 a_5978_3134# m2_6176_3382# 0.16fF
C3822 a_9994_5142# rowoff_n[3] 0.10fF
C3823 a_28066_4138# ctop 3.58fF
C3824 a_2346_1168# col[10] 0.14fF
C3825 a_2346_14220# col[12] 0.15fF
C3826 a_19030_13174# rowon_n[11] 0.14fF
C3827 m2_26832_946# m3_27968_1078# 0.13fF
C3828 a_2346_9200# a_18938_9158# 0.35fF
C3829 a_9994_9158# a_10998_9158# 0.97fF
C3830 a_1962_3174# col_n[26] 0.13fF
C3831 a_8990_3134# vcm 0.62fF
C3832 a_34090_3134# rowon_n[1] 0.14fF
C3833 a_20034_3134# rowoff_n[1] 0.10fF
C3834 row_n[15] ctop 1.37fF
C3835 VDD col[31] 4.08fF
C3836 vcm col[27] 5.84fF
C3837 a_1962_16226# col_n[28] 0.13fF
C3838 col_n[13] col[14] 5.98fF
C3839 a_13006_15182# col_n[10] 0.28fF
C3840 a_14010_2130# col[11] 0.29fF
C3841 a_1962_6186# a_13006_6146# 0.27fF
C3842 a_1962_10202# col[19] 0.11fF
C3843 a_15014_15182# VDD 0.52fF
C3844 a_2346_11208# a_31990_11166# 0.35fF
C3845 a_12002_3134# row_n[1] 0.17fF
C3846 a_31078_11166# col_n[28] 0.28fF
C3847 a_22042_7150# vcm 0.62fF
C3848 a_5278_16226# vcm 0.22fF
C3849 a_1962_3174# a_6282_3174# 0.14fF
C3850 a_22042_4138# a_22042_3134# 1.00fF
C3851 a_2346_3176# a_7986_3134# 0.19fF
C3852 a_1962_8194# a_26058_8154# 0.27fF
C3853 a_15318_1166# vcm 0.23fF
C3854 a_23046_13174# a_24050_13174# 0.97fF
C3855 a_35094_11166# vcm 0.12fF
C3856 a_8898_11166# rowoff_n[9] 0.24fF
C3857 a_16018_16186# row_n[14] 0.17fF
C3858 a_4882_3134# VDD 0.23fF
C3859 a_2346_10204# col[3] 0.15fF
C3860 a_2346_5184# a_21038_5142# 0.19fF
C3861 a_1962_5182# a_19334_5182# 0.14fF
C3862 a_11910_5142# a_12002_5142# 0.26fF
C3863 a_31078_6146# row_n[4] 0.17fF
C3864 a_14010_4138# col_n[11] 0.28fF
C3865 a_18938_9158# rowoff_n[7] 0.24fF
C3866 a_1962_12210# col_n[19] 0.13fF
C3867 a_28370_5182# vcm 0.22fF
C3868 a_22954_15182# rowoff_n[13] 0.24fF
C3869 m2_1732_7974# VDD 1.02fF
C3870 m2_34864_18014# m3_33992_18146# 0.13fF
C3871 a_17934_7150# VDD 0.23fF
C3872 a_1962_6186# col[10] 0.11fF
C3873 a_28978_7150# rowoff_n[5] 0.24fF
C3874 a_1962_7190# a_32386_7190# 0.14fF
C3875 a_2346_7192# a_34090_7150# 0.19fF
C3876 a_3970_14178# rowon_n[12] 0.14fF
C3877 a_29070_14178# col[26] 0.29fF
C3878 a_1962_16226# a_2966_16186# 0.27fF
C3879 a_2346_5184# col[30] 0.15fF
C3880 a_19030_4138# rowon_n[2] 0.14fF
C3881 a_23046_3134# ctop 3.57fF
C3882 a_30986_11166# VDD 0.23fF
C3883 m3_28972_1078# m3_29976_1078# 0.22fF
C3884 a_7986_9158# a_7986_8154# 1.00fF
C3885 a_24962_9158# a_25054_9158# 0.26fF
C3886 a_3970_2130# vcm 0.62fF
C3887 a_2346_1168# a_23958_1126# 0.35fF
C3888 a_34090_6146# m2_34288_6394# 0.16fF
C3889 a_2346_6188# ctop 1.59fF
C3890 m3_1046_19620# VDD 0.13fF
C3891 a_23046_17190# rowon_n[15] 0.14fF
C3892 a_9994_14178# VDD 0.52fF
C3893 a_12002_7150# col[9] 0.29fF
C3894 m2_34864_15002# rowon_n[13] 0.13fF
C3895 a_30074_17190# m3_29976_18146# 0.15fF
C3896 a_1962_8194# col_n[10] 0.13fF
C3897 a_17022_6146# vcm 0.62fF
C3898 a_1962_15222# a_10998_15182# 0.27fF
C3899 col[25] rowoff_n[10] 0.11fF
C3900 a_9994_16186# rowoff_n[14] 0.10fF
C3901 a_29070_16186# col_n[26] 0.28fF
C3902 m2_20808_946# m2_21812_946# 0.96fF
C3903 a_19030_3134# a_20034_3134# 0.97fF
C3904 a_1962_3174# a_1962_2170# 0.16fF
C3905 a_30074_3134# col[27] 0.29fF
C3906 a_1962_2170# col[1] 0.11fF
C3907 m2_19804_18014# col[17] 0.28fF
C3908 a_1962_15222# col[3] 0.11fF
C3909 m2_21812_18014# vcm 0.28fF
C3910 a_21038_13174# a_21038_12170# 1.00fF
C3911 a_1962_12210# a_4274_12210# 0.14fF
C3912 a_2346_12212# a_5978_12170# 0.19fF
C3913 a_16018_7150# row_n[5] 0.17fF
C3914 a_30074_10162# vcm 0.62fF
C3915 a_1962_17230# a_24050_17190# 0.27fF
C3916 a_2346_1168# col[21] 0.14fF
C3917 a_2346_14220# col[23] 0.15fF
C3918 m2_31852_18014# m2_32280_18442# 0.16fF
C3919 a_33086_3134# VDD 0.52fF
C3920 m3_7888_1078# ctop 0.23fF
C3921 rowon_n[9] ctop 1.40fF
C3922 rowon_n[4] rowon_n[3] 0.15fF
C3923 col_n[19] col[19] 0.72fF
C3924 a_10906_14178# a_10998_14178# 0.26fF
C3925 a_2346_14220# a_19030_14178# 0.19fF
C3926 a_1962_14218# a_17326_14218# 0.14fF
C3927 a_23350_4178# vcm 0.22fF
C3928 a_12002_9158# col_n[9] 0.28fF
C3929 col[9] rowoff_n[11] 0.11fF
C3930 a_1962_10202# col[30] 0.11fF
C3931 a_31078_7150# m2_31276_7398# 0.16fF
C3932 a_12914_6146# VDD 0.23fF
C3933 a_3970_5142# rowon_n[3] 0.14fF
C3934 a_32082_7150# a_33086_7150# 0.97fF
C3935 m2_9764_946# col[7] 0.39fF
C3936 a_7986_17190# ctop 3.39fF
C3937 a_30074_5142# col_n[27] 0.28fF
C3938 a_1962_4178# col_n[1] 0.13fF
C3939 a_1962_17230# col_n[3] 0.13fF
C3940 m2_1732_17010# row_n[15] 0.13fF
C3941 a_2346_16228# a_32082_16186# 0.19fF
C3942 a_1962_16226# a_30378_16226# 0.14fF
C3943 a_34090_17190# a_34090_16186# 1.00fF
C3944 a_18026_2130# ctop 3.46fF
C3945 m2_12776_18014# VDD 0.91fF
C3946 a_1962_18234# m2_27836_18014# 0.18fF
C3947 a_2346_9200# m2_1732_8978# 0.12fF
C3948 a_1962_11206# ctop 1.49fF
C3949 a_25966_10162# VDD 0.23fF
C3950 a_2346_8196# a_8898_8154# 0.35fF
C3951 a_4974_8154# a_5978_8154# 0.97fF
C3952 a_11910_4138# rowoff_n[2] 0.24fF
C3953 a_24962_12170# rowoff_n[10] 0.24fF
C3954 a_2346_10204# col[14] 0.15fF
C3955 a_23046_8154# rowon_n[6] 0.14fF
C3956 a_31078_6146# ctop 3.58fF
C3957 a_2346_5184# a_2966_5142# 0.21fF
C3958 a_2346_18236# m2_22816_18014# 0.19fF
C3959 a_4974_13174# VDD 0.52fF
C3960 a_1962_12210# col_n[30] 0.13fF
C3961 a_2346_10204# a_21950_10162# 0.35fF
C3962 a_21950_2130# rowoff_n[0] 0.24fF
C3963 a_12002_5142# vcm 0.62fF
C3964 a_9994_12170# col[7] 0.29fF
C3965 a_1962_6186# col[21] 0.11fF
C3966 a_17022_3134# a_17022_2130# 1.00fF
C3967 a_33998_3134# a_34090_3134# 0.26fF
C3968 a_28066_8154# m2_28264_8402# 0.16fF
C3969 m2_10768_18014# m3_10900_18146# 2.78fF
C3970 a_1962_7190# a_16018_7150# 0.27fF
C3971 a_18026_17190# VDD 0.55fF
C3972 a_18026_12170# a_19030_12170# 0.97fF
C3973 a_28066_8154# col[25] 0.29fF
C3974 a_2346_12212# a_35002_12170# 0.35fF
C3975 a_25054_9158# vcm 0.62fF
C3976 a_8290_18234# vcm 0.22fF
C3977 a_28066_2130# VDD 0.55fF
C3978 a_6890_4138# a_6982_4138# 0.26fF
C3979 a_1962_4178# a_9294_4178# 0.14fF
C3980 a_2346_4180# a_10998_4138# 0.19fF
C3981 m2_1732_8978# rowoff_n[7] 0.12fF
C3982 m3_1864_5094# m3_1864_4090# 0.22fF
C3983 a_1962_9198# a_29070_9158# 0.27fF
C3984 a_20946_18194# m2_20808_18014# 0.16fF
C3985 a_20034_11166# row_n[9] 0.17fF
C3986 a_18330_3174# vcm 0.22fF
C3987 a_9994_10162# rowoff_n[8] 0.10fF
C3988 a_2346_6188# col[5] 0.15fF
C3989 a_12002_13174# rowoff_n[11] 0.10fF
C3990 a_9994_14178# col_n[7] 0.28fF
C3991 a_7894_5142# VDD 0.23fF
C3992 a_2346_6188# a_24050_6146# 0.19fF
C3993 a_30074_7150# a_30074_6146# 1.00fF
C3994 a_1962_6186# a_22346_6186# 0.14fF
C3995 a_1962_8194# col_n[21] 0.13fF
C3996 a_20034_8154# rowoff_n[6] 0.10fF
C3997 a_31078_16186# a_32082_16186# 0.97fF
C3998 a_31382_7190# vcm 0.22fF
C3999 a_28066_10162# col_n[25] 0.28fF
C4000 a_1962_2170# col[12] 0.11fF
C4001 a_26058_17190# rowoff_n[15] 0.10fF
C4002 a_1962_15222# col[14] 0.11fF
C4003 a_30074_6146# rowoff_n[4] 0.10fF
C4004 a_25054_9158# m2_25252_9406# 0.16fF
C4005 a_20946_9158# VDD 0.23fF
C4006 a_7986_9158# rowon_n[7] 0.14fF
C4007 a_19942_8154# a_20034_8154# 0.26fF
C4008 a_1962_18234# a_11302_18234# 0.14fF
C4009 m2_8760_946# m2_9188_1374# 0.16fF
C4010 a_2346_17232# a_6890_17190# 0.35fF
C4011 a_3970_17190# a_4974_17190# 0.97fF
C4012 m2_13780_18014# m2_14784_18014# 0.96fF
C4013 a_2346_18236# col[6] 0.14fF
C4014 a_26058_5142# ctop 3.58fF
C4015 m3_3872_18146# ctop 0.23fF
C4016 col_n[24] col[25] 5.98fF
C4017 row_n[4] ctop 1.65fF
C4018 rowon_n[1] row_n[1] 19.75fF
C4019 a_33998_13174# VDD 0.23fF
C4020 col[20] rowoff_n[11] 0.11fF
C4021 a_6982_4138# vcm 0.62fF
C4022 a_10998_3134# col_n[8] 0.28fF
C4023 m2_34864_13998# ctop 0.17fF
C4024 a_27062_12170# rowon_n[10] 0.14fF
C4025 a_2346_2172# a_26970_2130# 0.35fF
C4026 a_14010_2130# a_15014_2130# 0.97fF
C4027 a_7986_17190# col[5] 0.29fF
C4028 a_1962_4178# col_n[12] 0.13fF
C4029 a_1962_17230# col_n[14] 0.13fF
C4030 a_13006_16186# VDD 0.52fF
C4031 a_16018_12170# a_16018_11166# 1.00fF
C4032 a_32994_12170# a_33086_12170# 0.26fF
C4033 a_1962_16226# a_14010_16186# 0.27fF
C4034 a_20034_8154# vcm 0.62fF
C4035 m2_34864_15002# m2_35292_15430# 0.16fF
C4036 a_4974_12170# row_n[10] 0.17fF
C4037 a_26058_13174# col[23] 0.29fF
C4038 a_1962_11206# col[5] 0.11fF
C4039 a_3270_17230# vcm 0.22fF
C4040 a_2346_16228# rowon_n[14] 0.26fF
C4041 a_22042_10162# m2_22240_10410# 0.16fF
C4042 a_20034_2130# row_n[0] 0.17fF
C4043 col[4] rowoff_n[12] 0.11fF
C4044 a_2346_13216# a_8990_13174# 0.19fF
C4045 a_5886_13174# a_5978_13174# 0.26fF
C4046 a_2346_10204# col[25] 0.15fF
C4047 a_13310_2170# vcm 0.22fF
C4048 a_1962_13214# a_7286_13214# 0.14fF
C4049 a_33086_12170# vcm 0.62fF
C4050 a_2346_4180# VDD 32.63fF
C4051 m3_1864_13126# VDD 0.25fF
C4052 a_27062_6146# a_28066_6146# 0.97fF
C4053 a_2346_10204# a_3878_10162# 0.35fF
C4054 a_2874_10162# a_2966_10162# 0.26fF
C4055 a_3878_2130# rowoff_n[0] 0.24fF
C4056 a_24050_15182# row_n[13] 0.17fF
C4057 a_26362_6186# vcm 0.22fF
C4058 a_8990_6146# col[6] 0.29fF
C4059 a_2346_15224# a_22042_15182# 0.19fF
C4060 a_29070_16186# a_29070_15182# 1.00fF
C4061 a_1962_15222# a_20338_15222# 0.14fF
C4062 a_15926_8154# VDD 0.23fF
C4063 a_26058_15182# col_n[23] 0.28fF
C4064 a_1962_13214# col_n[5] 0.13fF
C4065 a_27062_2130# col[24] 0.29fF
C4066 a_1962_17230# a_33390_17230# 0.14fF
C4067 a_18938_17190# a_19030_17190# 0.26fF
C4068 a_2874_5142# rowoff_n[3] 0.24fF
C4069 a_21038_4138# ctop 3.58fF
C4070 m2_10768_946# m3_11904_1078# 0.13fF
C4071 a_19030_11166# m2_19228_11414# 0.16fF
C4072 a_12002_13174# rowon_n[11] 0.14fF
C4073 a_28978_12170# VDD 0.23fF
C4074 m3_24956_18146# m3_25960_18146# 0.22fF
C4075 a_2346_9200# a_11910_9158# 0.35fF
C4076 a_2346_6188# col[16] 0.15fF
C4077 m2_34864_3958# row_n[2] 0.15fF
C4078 a_34394_4178# vcm 0.22fF
C4079 a_13006_3134# rowoff_n[1] 0.10fF
C4080 a_27062_3134# rowon_n[1] 0.14fF
C4081 a_28066_14178# rowoff_n[12] 0.10fF
C4082 a_28978_2130# a_29070_2130# 0.26fF
C4083 a_8990_8154# col_n[6] 0.28fF
C4084 a_34090_8154# ctop 3.42fF
C4085 a_1962_6186# a_5978_6146# 0.27fF
C4086 a_7986_15182# VDD 0.52fF
C4087 a_2346_11208# a_24962_11166# 0.35fF
C4088 a_13006_11166# a_14010_11166# 0.97fF
C4089 m2_13780_946# a_14010_2130# 0.99fF
C4090 a_4974_3134# row_n[1] 0.17fF
C4091 a_1962_2170# col[23] 0.11fF
C4092 a_2346_7192# rowon_n[5] 0.26fF
C4093 a_1962_15222# col[25] 0.11fF
C4094 a_15014_7150# vcm 0.62fF
C4095 a_26058_2130# m2_26256_2378# 0.16fF
C4096 a_27062_4138# col_n[24] 0.28fF
C4097 a_31078_16186# rowon_n[14] 0.14fF
C4098 a_1962_9198# VDD 2.73fF
C4099 a_1962_8194# a_19030_8154# 0.27fF
C4100 a_8290_1166# vcm 0.23fF
C4101 a_2966_13174# a_2966_12170# 1.00fF
C4102 a_2346_18236# col[17] 0.14fF
C4103 a_28066_11166# vcm 0.62fF
C4104 col_n[30] col[30] 0.86fF
C4105 a_8990_16186# row_n[14] 0.17fF
C4106 a_31078_4138# VDD 0.52fF
C4107 a_1962_5182# a_12306_5182# 0.14fF
C4108 a_16018_12170# m2_16216_12418# 0.16fF
C4109 a_25054_6146# a_25054_5142# 1.00fF
C4110 a_2346_5184# a_14010_5142# 0.19fF
C4111 col[31] rowoff_n[11] 0.11fF
C4112 a_24050_6146# row_n[4] 0.17fF
C4113 a_1962_10202# a_32082_10162# 0.27fF
C4114 a_2346_2172# col[7] 0.15fF
C4115 a_11910_9158# rowoff_n[7] 0.24fF
C4116 a_2346_15224# col[9] 0.15fF
C4117 a_26058_15182# a_27062_15182# 0.97fF
C4118 a_21342_5182# vcm 0.22fF
C4119 a_15926_15182# rowoff_n[13] 0.24fF
C4120 a_1962_4178# col_n[23] 0.13fF
C4121 a_6982_11166# col[4] 0.29fF
C4122 a_1962_17230# col_n[25] 0.13fF
C4123 m2_24824_18014# m3_25960_18146# 0.13fF
C4124 a_10906_7150# VDD 0.23fF
C4125 a_21950_7150# rowoff_n[5] 0.24fF
C4126 a_1962_7190# a_25358_7190# 0.14fF
C4127 a_2346_7192# a_27062_7150# 0.19fF
C4128 a_14922_7150# a_15014_7150# 0.26fF
C4129 a_1962_11206# col[16] 0.11fF
C4130 a_35398_9198# vcm 0.23fF
C4131 a_25054_7150# col[22] 0.29fF
C4132 a_31990_5142# rowoff_n[3] 0.24fF
C4133 a_12002_4138# rowon_n[2] 0.14fF
C4134 a_16018_3134# ctop 3.57fF
C4135 col[15] rowoff_n[12] 0.11fF
C4136 a_23958_11166# VDD 0.23fF
C4137 m3_14916_1078# m3_15920_1078# 0.22fF
C4138 a_2346_1168# a_16930_1126# 0.35fF
C4139 a_29070_7150# ctop 3.58fF
C4140 a_13006_13174# m2_13204_13422# 0.16fF
C4141 a_16018_17190# rowon_n[15] 0.14fF
C4142 a_2874_14178# VDD 0.24fF
C4143 a_6982_13174# col_n[4] 0.28fF
C4144 a_10998_11166# a_10998_10162# 1.00fF
C4145 a_27974_11166# a_28066_11166# 0.26fF
C4146 a_2346_11208# col[0] 0.15fF
C4147 a_1962_15222# a_3970_15182# 0.27fF
C4148 a_9994_6146# vcm 0.62fF
C4149 a_31078_7150# rowon_n[5] 0.14fF
C4150 a_2874_16186# rowoff_n[14] 0.24fF
C4151 a_1962_13214# col_n[16] 0.13fF
C4152 a_2346_3176# a_29982_3134# 0.35fF
C4153 a_25054_9158# col_n[22] 0.28fF
C4154 m2_7756_18014# vcm 0.28fF
C4155 a_1962_7190# col[7] 0.11fF
C4156 a_8990_7150# row_n[5] 0.17fF
C4157 a_30074_11166# rowoff_n[9] 0.10fF
C4158 a_23046_10162# vcm 0.62fF
C4159 a_1962_17230# a_17022_17190# 0.27fF
C4160 m2_24824_18014# m2_25252_18442# 0.16fF
C4161 a_2966_4138# ctop 3.41fF
C4162 a_26058_3134# VDD 0.52fF
C4163 m3_34996_12122# ctop 0.23fF
C4164 a_22042_5142# a_23046_5142# 0.97fF
C4165 a_2346_6188# col[27] 0.15fF
C4166 a_16322_4178# vcm 0.22fF
C4167 a_1962_14218# a_10298_14218# 0.14fF
C4168 a_2346_14220# a_12002_14178# 0.19fF
C4169 a_24050_15182# a_24050_14178# 1.00fF
C4170 a_2346_13216# vcm 0.40fF
C4171 a_7986_2130# col_n[5] 0.28fF
C4172 a_5886_6146# VDD 0.23fF
C4173 a_9994_14178# m2_10192_14426# 0.16fF
C4174 a_28066_10162# row_n[8] 0.17fF
C4175 a_4974_16186# col[2] 0.29fF
C4176 a_13918_16186# a_14010_16186# 0.26fF
C4177 a_1962_16226# a_23350_16226# 0.14fF
C4178 a_29374_8194# vcm 0.22fF
C4179 a_2346_16228# a_25054_16186# 0.19fF
C4180 m2_32856_946# col[30] 0.38fF
C4181 a_10998_2130# ctop 3.39fF
C4182 a_1962_9198# col_n[7] 0.13fF
C4183 a_1962_18234# m2_13780_18014# 0.18fF
C4184 a_23046_12170# col[20] 0.29fF
C4185 a_18938_10162# VDD 0.23fF
C4186 a_2346_18236# col[28] 0.14fF
C4187 a_1962_16226# col[0] 0.11fF
C4188 ctop col[5] 1.98fF
C4189 a_4882_4138# rowoff_n[2] 0.24fF
C4190 a_17934_12170# rowoff_n[10] 0.24fF
C4191 a_16018_8154# rowon_n[6] 0.14fF
C4192 a_24050_6146# ctop 3.58fF
C4193 m3_19936_1078# VDD 0.10fF
C4194 a_2346_2172# col[18] 0.15fF
C4195 a_2346_15224# col[20] 0.15fF
C4196 a_2346_18236# m2_8760_18014# 0.19fF
C4197 a_31990_14178# VDD 0.23fF
C4198 m2_2736_1950# vcm 0.44fF
C4199 a_7986_10162# a_8990_10162# 0.97fF
C4200 a_2346_10204# a_14922_10162# 0.35fF
C4201 a_14922_2130# rowoff_n[0] 0.24fF
C4202 a_4974_5142# vcm 0.62fF
C4203 m2_1732_17010# ctop 0.17fF
C4204 a_31990_16186# rowoff_n[14] 0.24fF
C4205 a_5978_5142# col[3] 0.29fF
C4206 a_3878_7150# rowoff_n[5] 0.24fF
C4207 a_1962_18234# col[10] 0.11fF
C4208 a_1962_7190# a_8990_7150# 0.27fF
C4209 a_6982_15182# m2_7180_15430# 0.16fF
C4210 a_1962_11206# col[27] 0.11fF
C4211 a_10998_17190# VDD 0.55fF
C4212 a_2346_12212# a_27974_12170# 0.35fF
C4213 a_23046_14178# col_n[20] 0.28fF
C4214 m2_21812_946# m3_21944_1078# 2.79fF
C4215 a_18026_9158# vcm 0.62fF
C4216 col[26] rowoff_n[12] 0.11fF
C4217 a_8990_3134# m2_9188_3382# 0.16fF
C4218 a_1962_5182# sample 0.14fF
C4219 a_2346_3176# m2_34864_2954# 0.17fF
C4220 a_21038_2130# VDD 0.55fF
C4221 a_20034_5142# a_20034_4138# 1.00fF
C4222 a_2346_4180# a_3970_4138# 0.19fF
C4223 m3_1864_12122# m3_1864_11118# 0.22fF
C4224 m2_31852_946# m3_32988_1078# 0.13fF
C4225 a_1962_9198# a_22042_9158# 0.27fF
C4226 a_21038_14178# a_22042_14178# 0.97fF
C4227 a_13006_11166# row_n[9] 0.17fF
C4228 a_11302_3174# vcm 0.22fF
C4229 a_2874_10162# rowoff_n[8] 0.24fF
C4230 a_31078_13174# vcm 0.62fF
C4231 a_4974_13174# rowoff_n[11] 0.10fF
C4232 a_34090_6146# VDD 0.54fF
C4233 a_2346_11208# col[11] 0.15fF
C4234 a_9902_6146# a_9994_6146# 0.26fF
C4235 a_2346_6188# a_17022_6146# 0.19fF
C4236 a_1962_6186# a_15318_6186# 0.14fF
C4237 a_13006_8154# rowoff_n[6] 0.10fF
C4238 a_5978_7150# col_n[3] 0.28fF
C4239 col[10] rowoff_n[13] 0.11fF
C4240 a_24354_7190# vcm 0.22fF
C4241 a_1962_13214# col_n[27] 0.13fF
C4242 a_35002_2130# m2_34864_1950# 0.16fF
C4243 a_19030_17190# rowoff_n[15] 0.10fF
C4244 a_23046_6146# rowoff_n[4] 0.10fF
C4245 a_24050_3134# col_n[21] 0.28fF
C4246 a_13918_9158# VDD 0.23fF
C4247 a_2346_8196# a_30074_8154# 0.19fF
C4248 a_1962_7190# col[18] 0.11fF
C4249 a_3970_16186# m2_4168_16434# 0.16fF
C4250 a_33086_9158# a_33086_8154# 1.00fF
C4251 a_1962_8194# a_28370_8194# 0.14fF
C4252 a_32082_14178# row_n[12] 0.17fF
C4253 a_21038_17190# col[18] 0.29fF
C4254 a_1962_18234# a_4274_18234# 0.14fF
C4255 a_33086_4138# rowoff_n[2] 0.10fF
C4256 m2_6752_18014# m2_7756_18014# 0.96fF
C4257 a_5978_4138# m2_6176_4386# 0.16fF
C4258 a_19030_5142# ctop 3.58fF
C4259 a_26970_13174# VDD 0.23fF
C4260 a_5978_10162# a_5978_9158# 1.00fF
C4261 a_22954_10162# a_23046_10162# 0.26fF
C4262 ctop rowoff_n[14] 0.60fF
C4263 a_20034_12170# rowon_n[10] 0.14fF
C4264 a_2346_2172# a_19942_2130# 0.35fF
C4265 a_32082_9158# ctop 3.58fF
C4266 a_2346_7192# col[2] 0.15fF
C4267 a_3970_10162# col[1] 0.29fF
C4268 a_5978_16186# VDD 0.52fF
C4269 a_1962_9198# col_n[18] 0.13fF
C4270 a_13006_8154# vcm 0.62fF
C4271 a_1962_16226# a_6982_16186# 0.27fF
C4272 a_2346_4180# a_32994_4138# 0.35fF
C4273 a_17022_4138# a_18026_4138# 0.97fF
C4274 a_22042_6146# col[19] 0.29fF
C4275 m2_34864_5966# rowon_n[4] 0.13fF
C4276 a_1962_3174# col[9] 0.11fF
C4277 a_13006_2130# row_n[0] 0.17fF
C4278 a_1962_16226# col[11] 0.11fF
C4279 ctop col[16] 2.03fF
C4280 a_6282_2170# vcm 0.22fF
C4281 a_19030_14178# a_19030_13174# 1.00fF
C4282 a_31990_10162# rowoff_n[8] 0.24fF
C4283 m2_34864_4962# m2_34864_3958# 0.99fF
C4284 a_26058_12170# vcm 0.62fF
C4285 a_33998_13174# rowoff_n[11] 0.24fF
C4286 a_2346_2172# col[29] 0.15fF
C4287 a_2346_15224# col[31] 0.15fF
C4288 a_29070_5142# VDD 0.52fF
C4289 m3_15920_18146# VDD 0.29fF
C4290 a_33086_17190# m3_32988_18146# 0.15fF
C4291 a_17022_15182# row_n[13] 0.17fF
C4292 a_1962_15222# a_13310_15222# 0.14fF
C4293 a_8898_15182# a_8990_15182# 0.26fF
C4294 a_19334_6186# vcm 0.22fF
C4295 a_2346_15224# a_15014_15182# 0.19fF
C4296 a_3970_12170# col_n[1] 0.28fF
C4297 a_1962_18234# col[21] 0.11fF
C4298 a_32082_5142# row_n[3] 0.17fF
C4299 a_8898_8154# VDD 0.23fF
C4300 a_30074_8154# a_31078_8154# 0.97fF
C4301 a_22042_8154# col_n[19] 0.28fF
C4302 a_1962_5182# col_n[9] 0.13fF
C4303 a_32386_10202# vcm 0.22fF
C4304 a_1962_17230# a_26362_17230# 0.14fF
C4305 a_2346_17232# a_28066_17190# 0.19fF
C4306 a_14010_4138# ctop 3.58fF
C4307 m3_22948_1078# ctop 0.23fF
C4308 a_4974_13174# rowon_n[11] 0.14fF
C4309 a_21950_12170# VDD 0.23fF
C4310 a_1962_12210# col[2] 0.11fF
C4311 m3_10900_18146# m3_11904_18146# 0.22fF
C4312 a_2346_9200# a_4882_9158# 0.35fF
C4313 m2_1732_7974# row_n[6] 0.13fF
C4314 a_5978_3134# rowoff_n[1] 0.10fF
C4315 a_20034_3134# rowon_n[1] 0.14fF
C4316 a_21038_14178# rowoff_n[12] 0.10fF
C4317 a_2346_11208# col[22] 0.15fF
C4318 a_34090_7150# m2_34288_7398# 0.16fF
C4319 a_27062_8154# ctop 3.58fF
C4320 col[21] rowoff_n[13] 0.11fF
C4321 a_35002_16186# VDD 0.29fF
C4322 m2_34864_9982# vcm 0.51fF
C4323 a_2346_11208# a_17934_11166# 0.35fF
C4324 sample_n rowoff_n[2] 0.38fF
C4325 VDD rowoff_n[1] 1.17fF
C4326 vcm rowoff_n[5] 0.20fF
C4327 a_7986_7150# vcm 0.62fF
C4328 a_1962_16226# a_34394_16226# 0.14fF
C4329 a_24050_16186# rowon_n[14] 0.14fF
C4330 a_1962_7190# col[29] 0.11fF
C4331 a_15014_4138# a_15014_3134# 1.00fF
C4332 a_31990_4138# a_32082_4138# 0.26fF
C4333 a_1962_8194# a_12002_8154# 0.27fF
C4334 a_20034_11166# col[17] 0.29fF
C4335 a_16018_13174# a_17022_13174# 0.97fF
C4336 a_1962_1166# vcm 7.69fF
C4337 a_2346_13216# a_30986_13174# 0.35fF
C4338 a_1962_14218# col_n[2] 0.13fF
C4339 m2_1732_1950# m2_2736_1950# 0.96fF
C4340 a_21038_11166# vcm 0.62fF
C4341 m2_13780_18014# col[11] 0.28fF
C4342 a_24050_4138# VDD 0.52fF
C4343 a_1962_5182# a_5278_5182# 0.14fF
C4344 a_2346_5184# a_6982_5142# 0.19fF
C4345 a_4882_5142# a_4974_5142# 0.26fF
C4346 col[5] rowoff_n[14] 0.11fF
C4347 a_17022_6146# row_n[4] 0.17fF
C4348 a_1962_10202# a_25054_10162# 0.27fF
C4349 a_4882_9158# rowoff_n[7] 0.24fF
C4350 a_14314_5182# vcm 0.22fF
C4351 a_2346_7192# col[13] 0.15fF
C4352 a_8898_15182# rowoff_n[13] 0.24fF
C4353 a_34090_15182# vcm 0.62fF
C4354 a_31078_8154# m2_31276_8402# 0.16fF
C4355 m2_15788_18014# m3_15920_18146# 2.79fF
C4356 a_14922_7150# rowoff_n[5] 0.24fF
C4357 a_28066_8154# a_28066_7150# 1.00fF
C4358 a_1962_7190# a_18330_7190# 0.14fF
C4359 a_2346_7192# a_20034_7150# 0.19fF
C4360 a_1962_9198# col_n[29] 0.13fF
C4361 a_29070_17190# a_30074_17190# 0.97fF
C4362 a_27366_9198# vcm 0.22fF
C4363 m2_1732_11990# sample_n 0.15fF
C4364 a_20034_13174# col_n[17] 0.28fF
C4365 a_24962_5142# rowoff_n[3] 0.24fF
C4366 a_4974_4138# rowon_n[2] 0.14fF
C4367 a_1962_3174# col[20] 0.11fF
C4368 a_8990_3134# ctop 3.57fF
C4369 VDD col_n[5] 4.94fF
C4370 vcm col_n[1] 2.79fF
C4371 ctop col[27] 1.98fF
C4372 col[10] col[11] 0.20fF
C4373 a_1962_16226# col[22] 0.11fF
C4374 a_2346_10204# m2_1732_9982# 0.12fF
C4375 a_16930_11166# VDD 0.23fF
C4376 m3_2868_2082# m3_2868_1078# 0.22fF
C4377 a_2346_9200# a_33086_9158# 0.19fF
C4378 a_1962_9198# a_31382_9198# 0.14fF
C4379 a_17934_9158# a_18026_9158# 0.26fF
C4380 m2_29844_18014# col_n[27] 0.25fF
C4381 a_35002_3134# rowoff_n[1] 0.24fF
C4382 a_2346_1168# a_9902_1126# 0.35fF
C4383 a_22042_7150# ctop 3.58fF
C4384 a_8990_17190# rowon_n[15] 0.14fF
C4385 a_29982_15182# VDD 0.23fF
C4386 m2_12776_946# a_2346_1168# 0.19fF
C4387 a_24050_7150# rowon_n[5] 0.14fF
C4388 a_2346_3176# col[4] 0.15fF
C4389 a_2346_16228# col[6] 0.15fF
C4390 a_2346_3176# a_22954_3134# 0.35fF
C4391 a_28066_9158# m2_28264_9406# 0.16fF
C4392 a_12002_3134# a_13006_3134# 0.97fF
C4393 a_2346_1168# m2_29844_946# 0.19fF
C4394 a_34090_2130# m2_33860_946# 0.99fF
C4395 a_1962_5182# col_n[20] 0.13fF
C4396 a_21038_2130# col_n[18] 0.28fF
C4397 a_30986_13174# a_31078_13174# 0.26fF
C4398 a_14010_13174# a_14010_12170# 1.00fF
C4399 a_1962_17230# a_9994_17190# 0.27fF
C4400 a_16018_10162# vcm 0.62fF
C4401 a_23046_11166# rowoff_n[9] 0.10fF
C4402 a_18026_16186# col[15] 0.29fF
C4403 m2_17796_18014# m2_18224_18442# 0.16fF
C4404 m2_34864_1950# m2_34864_946# 0.99fF
C4405 a_1962_12210# col[13] 0.11fF
C4406 a_19030_3134# VDD 0.52fF
C4407 m3_18932_18146# ctop 0.23fF
C4408 a_3878_12170# VDD 0.23fF
C4409 a_2966_9158# col[0] 0.29fF
C4410 a_33086_9158# rowoff_n[7] 0.10fF
C4411 a_9294_4178# vcm 0.22fF
C4412 a_2346_14220# a_4974_14178# 0.19fF
C4413 a_1962_14218# a_3270_14218# 0.14fF
C4414 a_2966_14178# rowoff_n[12] 0.10fF
C4415 a_29070_14178# vcm 0.62fF
C4416 a_1962_2170# a_30074_2130# 0.27fF
C4417 a_32082_7150# VDD 0.52fF
C4418 a_25054_7150# a_26058_7150# 0.97fF
C4419 a_21038_10162# row_n[8] 0.17fF
C4420 a_22346_8194# vcm 0.22fF
C4421 a_1962_16226# a_16322_16226# 0.14fF
C4422 a_2346_16228# a_18026_16186# 0.19fF
C4423 a_27062_17190# a_27062_16186# 1.00fF
C4424 a_3970_2130# ctop 3.27fF
C4425 a_25054_10162# m2_25252_10410# 0.16fF
C4426 a_11910_10162# VDD 0.23fF
C4427 a_1962_1166# col_n[11] 0.13fF
C4428 a_1962_14218# col_n[13] 0.13fF
C4429 a_19030_5142# col[16] 0.29fF
C4430 a_10906_12170# rowoff_n[10] 0.24fF
C4431 a_2966_11166# vcm 0.61fF
C4432 a_1962_8194# col[4] 0.11fF
C4433 a_8990_8154# rowon_n[6] 0.14fF
C4434 col[16] rowoff_n[14] 0.11fF
C4435 a_17022_6146# ctop 3.58fF
C4436 m3_34996_6098# VDD 0.26fF
C4437 a_24962_14178# VDD 0.23fF
C4438 a_2346_10204# a_7894_10162# 0.35fF
C4439 a_7894_2130# rowoff_n[0] 0.24fF
C4440 a_2346_7192# col[24] 0.15fF
C4441 a_24962_16186# rowoff_n[14] 0.24fF
C4442 m2_21812_18014# ctop 0.18fF
C4443 a_9994_3134# a_9994_2130# 1.00fF
C4444 a_26970_3134# a_27062_3134# 0.26fF
C4445 a_30074_10162# ctop 3.58fF
C4446 a_30986_1126# m2_30848_946# 0.16fF
C4447 a_3970_17190# VDD 0.56fF
C4448 a_2346_12212# a_20946_12170# 0.35fF
C4449 a_10998_12170# a_12002_12170# 0.97fF
C4450 m2_11772_946# m3_10900_1078# 0.13fF
C4451 a_1962_3174# col[31] 0.11fF
C4452 a_28066_11166# rowon_n[9] 0.14fF
C4453 vcm col_n[12] 2.80fF
C4454 a_10998_9158# vcm 0.62fF
C4455 VDD col_n[16] 4.70fF
C4456 col[0] rowoff_n[15] 0.11fF
C4457 a_19030_7150# col_n[16] 0.28fF
C4458 a_14010_2130# VDD 0.55fF
C4459 a_22042_11166# m2_22240_11414# 0.16fF
C4460 a_1962_10202# col_n[4] 0.13fF
C4461 a_1962_9198# a_15014_9158# 0.27fF
C4462 a_4274_3174# vcm 0.22fF
C4463 a_5978_11166# row_n[9] 0.17fF
C4464 a_2346_14220# a_33998_14178# 0.35fF
C4465 a_24050_13174# vcm 0.62fF
C4466 a_34090_17190# col[31] 0.29fF
C4467 a_27062_6146# VDD 0.52fF
C4468 a_23046_7150# a_23046_6146# 1.00fF
C4469 a_2346_6188# a_9994_6146# 0.19fF
C4470 a_1962_6186# a_8290_6186# 0.14fF
C4471 a_5978_8154# rowoff_n[6] 0.10fF
C4472 a_1962_11206# a_28066_11166# 0.27fF
C4473 a_2346_3176# col[15] 0.15fF
C4474 a_2346_16228# col[17] 0.15fF
C4475 a_17326_7190# vcm 0.22fF
C4476 a_24050_16186# a_25054_16186# 0.97fF
C4477 a_29070_2130# m2_29268_2378# 0.16fF
C4478 a_12002_17190# rowoff_n[15] 0.10fF
C4479 a_16018_6146# rowoff_n[4] 0.10fF
C4480 a_2966_3134# a_3970_3134# 0.97fF
C4481 a_1962_5182# col_n[31] 0.13fF
C4482 a_6890_9158# VDD 0.23fF
C4483 a_12914_8154# a_13006_8154# 0.26fF
C4484 a_1962_8194# a_21342_8194# 0.14fF
C4485 a_2346_8196# a_23046_8154# 0.19fF
C4486 a_25054_14178# row_n[12] 0.17fF
C4487 m2_16792_946# col_n[14] 0.37fF
C4488 a_1962_12210# col[24] 0.11fF
C4489 a_30378_11206# vcm 0.22fF
C4490 a_26058_4138# rowoff_n[2] 0.10fF
C4491 a_17022_10162# col[14] 0.29fF
C4492 a_12002_5142# ctop 3.58fF
C4493 a_19030_12170# m2_19228_12418# 0.16fF
C4494 a_19942_13174# VDD 0.23fF
C4495 a_2346_10204# a_2346_9200# 0.22fF
C4496 a_1962_10202# a_35398_10202# 0.14fF
C4497 a_13006_12170# rowon_n[10] 0.14fF
C4498 a_2346_2172# a_12914_2130# 0.35fF
C4499 a_6982_2130# a_7986_2130# 0.97fF
C4500 m2_29844_18014# m3_30980_18146# 0.13fF
C4501 a_25054_9158# ctop 3.58fF
C4502 a_2966_10162# row_n[8] 0.16fF
C4503 a_28066_2130# rowon_n[0] 0.14fF
C4504 a_32994_17190# VDD 0.24fF
C4505 m2_1732_12994# vcm 0.45fF
C4506 a_8990_12170# a_8990_11166# 1.00fF
C4507 a_25966_12170# a_26058_12170# 0.26fF
C4508 a_2346_12212# col[8] 0.15fF
C4509 a_5978_8154# vcm 0.62fF
C4510 a_1962_1166# col_n[22] 0.13fF
C4511 a_2346_4180# a_25966_4138# 0.35fF
C4512 a_1962_14218# col_n[24] 0.13fF
C4513 m2_1732_9982# rowon_n[8] 0.11fF
C4514 a_17022_12170# col_n[14] 0.28fF
C4515 a_5978_2130# row_n[0] 0.17fF
C4516 a_7986_17190# m2_7756_18014# 1.00fF
C4517 m2_11772_946# VDD 0.62fF
C4518 a_24962_10162# rowoff_n[8] 0.24fF
C4519 col[27] rowoff_n[14] 0.11fF
C4520 a_1962_8194# col[15] 0.11fF
C4521 a_32082_15182# rowon_n[13] 0.14fF
C4522 a_19030_12170# vcm 0.62fF
C4523 a_26970_13174# rowoff_n[11] 0.24fF
C4524 a_1962_1166# a_20034_1126# 0.26fF
C4525 a_22042_5142# VDD 0.52fF
C4526 m2_28840_946# VDD 0.62fF
C4527 a_16018_13174# m2_16216_13422# 0.16fF
C4528 a_20034_6146# a_21038_6146# 0.97fF
C4529 a_35002_8154# rowoff_n[6] 0.24fF
C4530 a_9994_15182# row_n[13] 0.17fF
C4531 a_12306_6186# vcm 0.22fF
C4532 a_1962_15222# a_6282_15222# 0.14fF
C4533 a_22042_16186# a_22042_15182# 1.00fF
C4534 a_2346_15224# a_7986_15182# 0.19fF
C4535 a_32082_16186# vcm 0.62fF
C4536 a_1962_3174# a_33086_3134# 0.27fF
C4537 a_25054_5142# row_n[3] 0.17fF
C4538 a_22042_2130# m3_21944_1078# 0.15fF
C4539 col_n[11] col_n[12] 0.10fF
C4540 VDD col_n[27] 4.97fF
C4541 vcm col_n[23] 2.80fF
C4542 col[21] col[22] 0.20fF
C4543 col[11] rowoff_n[15] 0.11fF
C4544 a_2346_12212# a_1962_12210# 2.62fF
C4545 a_2346_17232# a_21038_17190# 0.19fF
C4546 a_25358_10202# vcm 0.22fF
C4547 a_1962_17230# a_19334_17230# 0.14fF
C4548 a_11910_17190# a_12002_17190# 0.26fF
C4549 a_18026_1126# col_n[15] 0.31fF
C4550 a_6982_4138# ctop 3.58fF
C4551 a_1962_10202# col_n[15] 0.13fF
C4552 m3_1864_4090# ctop 0.23fF
C4553 a_15014_15182# col[12] 0.29fF
C4554 a_14922_12170# VDD 0.23fF
C4555 a_33086_10162# a_34090_10162# 0.97fF
C4556 a_1962_4178# col[6] 0.11fF
C4557 a_13006_3134# rowon_n[1] 0.14fF
C4558 a_1962_17230# col[8] 0.11fF
C4559 a_14010_14178# rowoff_n[12] 0.10fF
C4560 a_33086_11166# col[30] 0.29fF
C4561 a_21950_2130# a_22042_2130# 0.26fF
C4562 a_20034_8154# ctop 3.58fF
C4563 a_13006_14178# m2_13204_14426# 0.16fF
C4564 a_2346_3176# col[26] 0.15fF
C4565 a_27974_16186# VDD 0.23fF
C4566 a_2346_16228# col[28] 0.15fF
C4567 a_5978_11166# a_6982_11166# 0.97fF
C4568 a_2346_11208# a_10906_11166# 0.35fF
C4569 a_6982_2130# m2_6752_946# 0.99fF
C4570 a_17022_16186# rowon_n[14] 0.14fF
C4571 a_33086_12170# ctop 3.57fF
C4572 a_27062_17190# m2_26832_18014# 1.00fF
C4573 a_1962_8194# a_4974_8154# 0.27fF
C4574 a_3878_8154# a_3970_8154# 0.26fF
C4575 a_32082_6146# rowon_n[4] 0.14fF
C4576 a_15014_17190# col_n[12] 0.28fF
C4577 a_2346_13216# a_23958_13174# 0.35fF
C4578 a_16018_4138# col[13] 0.29fF
C4579 a_14010_11166# vcm 0.62fF
C4580 a_1962_6186# col_n[6] 0.13fF
C4581 a_17022_4138# VDD 0.52fF
C4582 a_18026_6146# a_18026_5142# 1.00fF
C4583 a_9994_6146# row_n[4] 0.17fF
C4584 a_35494_14540# VDD 0.11fF
C4585 a_33086_13174# col_n[30] 0.28fF
C4586 a_1962_10202# a_18026_10162# 0.27fF
C4587 a_1962_15222# a_1962_14218# 0.16fF
C4588 a_19030_15182# a_20034_15182# 0.97fF
C4589 a_7286_5182# vcm 0.22fF
C4590 a_27062_15182# vcm 0.62fF
C4591 m2_6752_18014# m3_5880_18146# 0.13fF
C4592 a_18026_1126# m3_17928_1078# 2.08fF
C4593 a_30074_8154# VDD 0.52fF
C4594 a_7894_7150# rowoff_n[5] 0.24fF
C4595 a_7894_7150# a_7986_7150# 0.26fF
C4596 a_9994_15182# m2_10192_15430# 0.16fF
C4597 a_1962_7190# a_11302_7190# 0.14fF
C4598 a_2346_7192# a_13006_7150# 0.19fF
C4599 a_2346_12212# col[19] 0.15fF
C4600 a_1962_12210# a_31078_12170# 0.27fF
C4601 a_20338_9198# vcm 0.22fF
C4602 a_12002_3134# m2_12200_3382# 0.16fF
C4603 a_17934_5142# rowoff_n[3] 0.24fF
C4604 a_29070_9158# row_n[7] 0.17fF
C4605 a_16018_6146# col_n[13] 0.28fF
C4606 a_2966_4138# m3_1864_4090# 0.14fF
C4607 a_9902_11166# VDD 0.23fF
C4608 a_31078_10162# a_31078_9158# 1.00fF
C4609 a_2346_9200# a_26058_9158# 0.19fF
C4610 a_1962_9198# a_24354_9198# 0.14fF
C4611 a_1962_8194# col[26] 0.11fF
C4612 m2_26832_946# col[24] 0.39fF
C4613 a_27974_3134# rowoff_n[1] 0.24fF
C4614 a_33390_13214# vcm 0.22fF
C4615 a_34090_2130# col_n[31] 0.33fF
C4616 a_1962_15222# col_n[0] 0.13fF
C4617 a_15014_7150# ctop 3.58fF
C4618 a_31078_16186# col[28] 0.29fF
C4619 a_22954_15182# VDD 0.23fF
C4620 a_20946_11166# a_21038_11166# 0.26fF
C4621 a_3970_11166# a_3970_10162# 1.00fF
C4622 a_17022_7150# rowon_n[5] 0.14fF
C4623 a_2346_1168# m2_5748_946# 0.19fF
C4624 a_2346_3176# a_15926_3134# 0.35fF
C4625 a_28066_11166# ctop 3.58fF
C4626 vcm rowon_n[14] 0.50fF
C4627 VDD rowon_n[12] 2.61fF
C4628 col_n[0] row_n[14] 0.23fF
C4629 col_n[1] row_n[15] 0.23fF
C4630 a_2346_8196# col[10] 0.15fF
C4631 col[22] rowoff_n[15] 0.11fF
C4632 a_6982_16186# m2_7180_16434# 0.16fF
C4633 a_16018_11166# rowoff_n[9] 0.10fF
C4634 a_8990_10162# vcm 0.62fF
C4635 a_1962_10202# col_n[26] 0.13fF
C4636 a_2346_17232# a_2966_17190# 0.21fF
C4637 a_8990_4138# m2_9188_4386# 0.16fF
C4638 m2_10768_18014# m2_11196_18442# 0.16fF
C4639 a_2346_4180# m2_34864_3958# 0.17fF
C4640 a_12002_3134# VDD 0.52fF
C4641 a_2346_5184# a_28978_5142# 0.35fF
C4642 a_14010_9158# col[11] 0.29fF
C4643 a_15014_5142# a_16018_5142# 0.97fF
C4644 a_1962_4178# col[17] 0.11fF
C4645 a_1962_17230# col[19] 0.11fF
C4646 a_26058_9158# rowoff_n[7] 0.10fF
C4647 a_17022_15182# a_17022_14178# 1.00fF
C4648 a_33998_15182# a_34090_15182# 0.26fF
C4649 m2_1732_7974# m2_1732_6970# 0.99fF
C4650 a_22042_14178# vcm 0.62fF
C4651 a_30074_15182# rowoff_n[13] 0.10fF
C4652 a_32082_5142# col[29] 0.29fF
C4653 a_1962_2170# a_23046_2130# 0.27fF
C4654 a_25054_7150# VDD 0.52fF
C4655 a_14010_10162# row_n[8] 0.17fF
C4656 a_1962_16226# a_9294_16226# 0.14fF
C4657 a_6890_16186# a_6982_16186# 0.26fF
C4658 a_15318_8194# vcm 0.22fF
C4659 a_2346_16228# a_10998_16186# 0.19fF
C4660 a_35094_18194# vcm 0.12fF
C4661 a_2346_4180# col[1] 0.15fF
C4662 a_4882_10162# VDD 0.23fF
C4663 a_2346_17232# col[3] 0.15fF
C4664 a_3970_17190# m2_4168_17438# 0.16fF
C4665 a_28066_9158# a_29070_9158# 0.97fF
C4666 a_14010_11166# col_n[11] 0.28fF
C4667 a_1962_6186# col_n[17] 0.13fF
C4668 a_28370_12210# vcm 0.22fF
C4669 a_5978_5142# m2_6176_5390# 0.16fF
C4670 a_1962_1166# a_29374_1166# 0.14fF
C4671 a_9994_6146# ctop 3.58fF
C4672 a_33086_13174# row_n[11] 0.17fF
C4673 m3_30980_18146# VDD 0.38fF
C4674 a_17934_14178# VDD 0.23fF
C4675 a_32082_7150# col_n[29] 0.28fF
C4676 a_1962_13214# col[10] 0.11fF
C4677 m2_7756_18014# ctop 0.18fF
C4678 a_17934_16186# rowoff_n[14] 0.24fF
C4679 a_2346_12212# col[30] 0.15fF
C4680 a_23046_10162# ctop 3.58fF
C4681 a_3970_1126# m3_2868_1078# 0.15fF
C4682 a_30986_18194# VDD 0.34fF
C4683 a_2346_12212# a_13918_12170# 0.35fF
C4684 a_21038_11166# rowon_n[9] 0.14fF
C4685 a_3970_9158# vcm 0.62fF
C4686 m2_6752_946# m3_6884_1078# 2.79fF
C4687 a_6982_2130# VDD 0.55fF
C4688 a_29982_5142# a_30074_5142# 0.26fF
C4689 a_13006_5142# a_13006_4138# 1.00fF
C4690 a_2346_13216# ctop 1.59fF
C4691 m3_1864_18146# m3_1864_17142# 0.22fF
C4692 a_6890_18194# m2_6752_18014# 0.16fF
C4693 a_1962_9198# a_7986_9158# 0.27fF
C4694 a_12002_14178# col[9] 0.29fF
C4695 a_2346_14220# a_26970_14178# 0.35fF
C4696 a_14010_14178# a_15014_14178# 0.97fF
C4697 a_1962_2170# col_n[8] 0.13fF
C4698 a_1962_15222# col_n[10] 0.13fF
C4699 a_17022_13174# vcm 0.62fF
C4700 m2_1732_3958# VDD 1.02fF
C4701 a_20034_6146# VDD 0.52fF
C4702 a_2346_6188# a_2874_6146# 0.35fF
C4703 a_30074_10162# col[27] 0.29fF
C4704 a_1962_9198# col[1] 0.11fF
C4705 a_1962_11206# a_21038_11166# 0.27fF
C4706 a_10298_7190# vcm 0.22fF
C4707 col_n[6] row_n[12] 0.23fF
C4708 col_n[22] col_n[23] 0.10fF
C4709 VDD row_n[7] 2.93fF
C4710 vcm row_n[9] 0.49fF
C4711 col_n[4] row_n[11] 0.23fF
C4712 col_n[2] row_n[10] 0.23fF
C4713 col_n[12] row_n[15] 0.23fF
C4714 col_n[8] row_n[13] 0.23fF
C4715 sample row_n[8] 1.03fF
C4716 col_n[10] row_n[14] 0.23fF
C4717 a_30074_17190# vcm 0.60fF
C4718 a_4974_17190# rowoff_n[15] 0.10fF
C4719 a_2346_8196# col[21] 0.15fF
C4720 m2_27836_18014# VDD 1.04fF
C4721 a_8990_6146# rowoff_n[4] 0.10fF
C4722 a_33086_10162# VDD 0.52fF
C4723 a_26058_9158# a_26058_8154# 1.00fF
C4724 a_2346_8196# a_16018_8154# 0.19fF
C4725 a_1962_8194# a_14314_8194# 0.14fF
C4726 a_18026_14178# row_n[12] 0.17fF
C4727 a_1962_13214# a_34090_13174# 0.27fF
C4728 a_19030_4138# rowoff_n[2] 0.10fF
C4729 a_33086_4138# row_n[2] 0.17fF
C4730 m2_2736_1950# ctop 0.36fF
C4731 a_32082_12170# rowoff_n[10] 0.10fF
C4732 a_23350_11206# vcm 0.22fF
C4733 a_12002_16186# col_n[9] 0.28fF
C4734 a_4974_5142# ctop 3.58fF
C4735 a_1962_4178# col[28] 0.11fF
C4736 a_13006_3134# col[10] 0.29fF
C4737 a_1962_17230# col[30] 0.11fF
C4738 a_12914_13174# VDD 0.23fF
C4739 a_2346_10204# a_29070_10162# 0.19fF
C4740 a_1962_10202# a_27366_10202# 0.14fF
C4741 a_15926_10162# a_16018_10162# 0.26fF
C4742 a_29070_2130# rowoff_n[0] 0.10fF
C4743 a_1962_11206# col_n[1] 0.13fF
C4744 a_30074_12170# col_n[27] 0.28fF
C4745 m2_23820_946# vcm 0.42fF
C4746 a_5978_12170# rowon_n[10] 0.14fF
C4747 a_2346_2172# a_5886_2130# 0.35fF
C4748 a_34090_8154# m2_34288_8402# 0.16fF
C4749 a_18026_9158# ctop 3.58fF
C4750 vcm rowoff_n[12] 0.20fF
C4751 m2_20808_18014# m3_20940_18146# 2.78fF
C4752 a_21038_2130# rowon_n[0] 0.14fF
C4753 a_25966_17190# VDD 0.24fF
C4754 a_2346_4180# col[12] 0.15fF
C4755 a_2346_17232# col[14] 0.15fF
C4756 a_2346_4180# a_18938_4138# 0.35fF
C4757 a_9994_4138# a_10998_4138# 0.97fF
C4758 a_31078_13174# ctop 3.58fF
C4759 a_25966_18194# m2_25828_18014# 0.16fF
C4760 a_1962_6186# col_n[28] 0.13fF
C4761 a_2966_13174# m3_1864_13126# 0.14fF
C4762 a_13006_5142# col_n[10] 0.28fF
C4763 a_12002_14178# a_12002_13174# 1.00fF
C4764 a_28978_14178# a_29070_14178# 0.26fF
C4765 a_17934_10162# rowoff_n[8] 0.24fF
C4766 a_25054_15182# rowon_n[13] 0.14fF
C4767 a_12002_12170# vcm 0.62fF
C4768 a_19942_13174# rowoff_n[11] 0.24fF
C4769 m2_4744_946# VDD 0.61fF
C4770 a_1962_13214# col[21] 0.11fF
C4771 a_15014_5142# VDD 0.52fF
C4772 a_2346_6188# a_31990_6146# 0.35fF
C4773 rowon_n[4] rowoff_n[4] 20.27fF
C4774 a_27974_8154# rowoff_n[6] 0.24fF
C4775 m2_21812_946# a_2346_1168# 0.19fF
C4776 m2_7756_18014# col[5] 0.28fF
C4777 a_28066_15182# col[25] 0.29fF
C4778 a_5278_6186# vcm 0.22fF
C4779 a_33998_17190# rowoff_n[15] 0.24fF
C4780 a_25054_16186# vcm 0.62fF
C4781 a_18026_5142# row_n[3] 0.17fF
C4782 a_1962_3174# a_26058_3134# 0.27fF
C4783 a_31078_9158# m2_31276_9406# 0.16fF
C4784 a_28066_9158# VDD 0.52fF
C4785 a_23046_8154# a_24050_8154# 0.97fF
C4786 a_2966_11166# rowon_n[9] 0.13fF
C4787 a_18330_10202# vcm 0.22fF
C4788 a_2346_17232# a_14010_17190# 0.19fF
C4789 a_1962_17230# a_12306_17230# 0.14fF
C4790 a_2346_13216# col[5] 0.15fF
C4791 m3_33992_18146# ctop 0.23fF
C4792 a_2346_11208# m2_1732_10986# 0.12fF
C4793 a_7894_12170# VDD 0.23fF
C4794 a_1962_2170# col_n[19] 0.13fF
C4795 a_1962_15222# col_n[21] 0.13fF
C4796 a_10998_8154# col[8] 0.29fF
C4797 a_5978_3134# rowon_n[1] 0.14fF
C4798 a_31382_14218# vcm 0.22fF
C4799 a_6982_14178# rowoff_n[12] 0.10fF
C4800 a_1962_2170# a_32386_2170# 0.14fF
C4801 a_2346_2172# a_34090_2130# 0.19fF
C4802 a_1962_9198# col[12] 0.11fF
C4803 a_28066_17190# col_n[25] 0.28fF
C4804 a_13006_8154# ctop 3.58fF
C4805 m2_23820_18014# col_n[21] 0.25fF
C4806 a_29070_4138# col[26] 0.29fF
C4807 a_20946_16186# VDD 0.23fF
C4808 a_1962_11206# a_2966_11166# 0.27fF
C4809 vcm rowon_n[3] 0.50fF
C4810 col_n[13] row_n[10] 0.23fF
C4811 col_n[19] row_n[13] 0.23fF
C4812 col_n[7] row_n[7] 0.23fF
C4813 col_n[9] row_n[8] 0.23fF
C4814 col_n[17] row_n[12] 0.23fF
C4815 col_n[3] row_n[5] 0.23fF
C4816 col_n[0] row_n[3] 0.23fF
C4817 col_n[21] row_n[14] 0.23fF
C4818 col_n[15] row_n[11] 0.23fF
C4819 col_n[11] row_n[9] 0.23fF
C4820 col_n[1] row_n[4] 0.23fF
C4821 VDD rowon_n[1] 2.61fF
C4822 col_n[5] row_n[6] 0.23fF
C4823 col_n[23] row_n[15] 0.23fF
C4824 a_1962_2170# m2_34864_1950# 0.17fF
C4825 a_30986_1126# VDD 0.44fF
C4826 a_9994_16186# rowon_n[14] 0.14fF
C4827 a_24962_4138# a_25054_4138# 0.26fF
C4828 a_7986_4138# a_7986_3134# 1.00fF
C4829 a_28066_10162# m2_28264_10410# 0.16fF
C4830 a_26058_12170# ctop 3.58fF
C4831 a_25054_6146# rowon_n[4] 0.14fF
C4832 a_8990_13174# a_9994_13174# 0.97fF
C4833 a_2346_13216# a_16930_13174# 0.35fF
C4834 a_6982_11166# vcm 0.62fF
C4835 a_10998_10162# col_n[8] 0.28fF
C4836 a_9994_4138# VDD 0.52fF
C4837 m3_6884_1078# VDD 0.14fF
C4838 a_1962_10202# a_10998_10162# 0.27fF
C4839 a_1962_11206# col_n[12] 0.13fF
C4840 a_29070_6146# col_n[26] 0.28fF
C4841 a_2346_15224# a_29982_15182# 0.35fF
C4842 a_2966_8154# col_n[0] 0.28fF
C4843 a_20034_15182# vcm 0.62fF
C4844 a_1962_5182# col[3] 0.11fF
C4845 a_23046_8154# VDD 0.52fF
C4846 a_21038_8154# a_21038_7150# 1.00fF
C4847 a_2346_7192# a_5978_7150# 0.19fF
C4848 a_1962_7190# a_4274_7190# 0.14fF
C4849 a_1962_12210# a_24050_12170# 0.27fF
C4850 m2_16792_946# m3_15920_1078# 0.13fF
C4851 a_2346_4180# col[23] 0.15fF
C4852 a_22042_17190# a_23046_17190# 0.97fF
C4853 a_13310_9198# vcm 0.22fF
C4854 a_2346_17232# col[25] 0.15fF
C4855 a_10906_5142# rowoff_n[3] 0.24fF
C4856 a_22042_9158# row_n[7] 0.17fF
C4857 a_25054_11166# m2_25252_11414# 0.16fF
C4858 a_2346_11208# VDD 32.63fF
C4859 m2_27836_946# m3_27968_1078# 2.79fF
C4860 a_1962_9198# a_17326_9198# 0.14fF
C4861 a_2346_9200# a_19030_9158# 0.19fF
C4862 a_10906_9158# a_10998_9158# 0.26fF
C4863 a_20946_3134# rowoff_n[1] 0.24fF
C4864 m2_1732_16006# sample 0.19fF
C4865 a_8990_13174# col[6] 0.29fF
C4866 a_26362_13214# vcm 0.22fF
C4867 m2_34864_9982# ctop 0.17fF
C4868 a_32082_2130# a_33086_2130# 0.97fF
C4869 ctop rowoff_n[5] 0.60fF
C4870 a_7986_7150# ctop 3.58fF
C4871 a_1962_7190# col_n[3] 0.13fF
C4872 a_15926_15182# VDD 0.23fF
C4873 a_34090_12170# a_34090_11166# 1.00fF
C4874 a_2346_11208# a_32082_11166# 0.19fF
C4875 a_1962_11206# a_30378_11206# 0.14fF
C4876 a_27062_9158# col[24] 0.29fF
C4877 a_9994_7150# rowon_n[5] 0.14fF
C4878 a_32082_2130# m2_32280_2378# 0.16fF
C4879 m2_34864_12994# m2_35292_13422# 0.16fF
C4880 a_1962_1166# ctop 0.26fF
C4881 a_4974_3134# a_5978_3134# 0.97fF
C4882 a_2346_3176# a_8898_3134# 0.35fF
C4883 a_21038_11166# ctop 3.58fF
C4884 a_6982_13174# a_6982_12170# 1.00fF
C4885 a_23958_13174# a_24050_13174# 0.26fF
C4886 a_2346_13216# col[16] 0.15fF
C4887 a_8990_11166# rowoff_n[9] 0.10fF
C4888 a_34394_11206# vcm 0.22fF
C4889 m2_3740_18014# m2_4168_18442# 0.16fF
C4890 a_4974_3134# VDD 0.52fF
C4891 a_1962_2170# col_n[30] 0.13fF
C4892 a_22042_12170# m2_22240_12418# 0.16fF
C4893 a_2346_5184# a_21950_5142# 0.35fF
C4894 a_8990_15182# col_n[6] 0.28fF
C4895 a_34090_15182# ctop 3.42fF
C4896 a_29070_10162# rowon_n[8] 0.14fF
C4897 a_9994_2130# col[7] 0.29fF
C4898 a_19030_9158# rowoff_n[7] 0.10fF
C4899 a_1962_9198# col[23] 0.11fF
C4900 a_15014_14178# vcm 0.62fF
C4901 a_23046_15182# rowoff_n[13] 0.10fF
C4902 a_27062_11166# col_n[24] 0.28fF
C4903 a_1962_2170# a_16018_2130# 0.27fF
C4904 a_18026_7150# VDD 0.52fF
C4905 a_29070_7150# rowoff_n[5] 0.10fF
C4906 a_2346_7192# a_35002_7150# 0.35fF
C4907 a_18026_7150# a_19030_7150# 0.97fF
C4908 a_6982_10162# row_n[8] 0.17fF
C4909 col_n[12] row_n[4] 0.23fF
C4910 col_n[4] row_n[0] 0.23fF
C4911 col_n[6] row_n[1] 0.23fF
C4912 VDD analog_in 0.48fF
C4913 col_n[28] row_n[12] 0.23fF
C4914 col_n[8] row_n[2] 0.23fF
C4915 col_n[30] row_n[13] 0.23fF
C4916 col_n[14] row_n[5] 0.23fF
C4917 col_n[22] row_n[9] 0.23fF
C4918 col_n[10] row_n[3] 0.23fF
C4919 col_n[24] row_n[10] 0.23fF
C4920 a_1962_16226# VDD 2.73fF
C4921 col_n[18] row_n[7] 0.23fF
C4922 col_n[1] ctop 2.00fF
C4923 col_n[16] row_n[6] 0.23fF
C4924 col_n[20] row_n[8] 0.23fF
C4925 col_n[26] row_n[11] 0.23fF
C4926 a_8290_8194# vcm 0.22fF
C4927 a_20034_17190# a_20034_16186# 1.00fF
C4928 a_2346_16228# a_3970_16186# 0.19fF
C4929 a_28066_18194# vcm 0.12fF
C4930 a_1962_4178# a_29070_4138# 0.27fF
C4931 a_31078_11166# VDD 0.52fF
C4932 m3_29976_1078# m3_30980_1078# 0.22fF
C4933 m2_20808_946# VDD 0.60fF
C4934 a_2346_9200# col[7] 0.15fF
C4935 a_9994_4138# col_n[7] 0.28fF
C4936 a_21342_12210# vcm 0.22fF
C4937 a_1962_1166# a_22346_1166# 0.14fF
C4938 a_1962_18234# col_n[6] 0.13fF
C4939 a_26058_13174# row_n[11] 0.17fF
C4940 a_1962_11206# col_n[23] 0.13fF
C4941 m3_2868_18146# VDD 0.37fF
C4942 a_19030_13174# m2_19228_13422# 0.16fF
C4943 a_10906_14178# VDD 0.23fF
C4944 a_31078_11166# a_32082_11166# 0.97fF
C4945 m2_15788_946# a_15926_1126# 0.16fF
C4946 a_1962_5182# col[14] 0.11fF
C4947 a_35398_16226# vcm 0.23fF
C4948 a_10906_16186# rowoff_n[14] 0.24fF
C4949 a_25054_14178# col[22] 0.29fF
C4950 a_19942_3134# a_20034_3134# 0.26fF
C4951 a_16018_10162# ctop 3.58fF
C4952 a_25054_2130# m3_24956_1078# 0.15fF
C4953 a_23958_18194# VDD 0.33fF
C4954 a_3970_12170# a_4974_12170# 0.97fF
C4955 a_2346_12212# a_6890_12170# 0.35fF
C4956 m2_22816_18014# vcm 0.28fF
C4957 a_14010_11166# rowon_n[9] 0.14fF
C4958 a_33998_3134# VDD 0.23fF
C4959 m3_9896_1078# ctop 0.23fF
C4960 a_29070_14178# ctop 3.58fF
C4961 a_2346_14220# a_19942_14178# 0.35fF
C4962 col[4] rowoff_n[4] 0.11fF
C4963 col[3] rowoff_n[3] 0.11fF
C4964 col[6] rowoff_n[6] 0.11fF
C4965 col[5] rowoff_n[5] 0.11fF
C4966 col[0] rowoff_n[0] 0.11fF
C4967 col[2] rowoff_n[2] 0.11fF
C4968 col[1] rowoff_n[1] 0.11fF
C4969 col[8] rowoff_n[8] 0.11fF
C4970 col[7] rowoff_n[7] 0.11fF
C4971 col[9] rowoff_n[9] 0.11fF
C4972 a_2346_18236# a_28978_18194# 0.35fF
C4973 a_7986_7150# col[5] 0.29fF
C4974 a_9994_13174# vcm 0.62fF
C4975 m2_1732_13998# m3_1864_15134# 0.15fF
C4976 a_1962_7190# col_n[14] 0.13fF
C4977 a_13006_6146# VDD 0.52fF
C4978 a_16018_14178# m2_16216_14426# 0.16fF
C4979 a_16018_7150# a_16018_6146# 1.00fF
C4980 a_32994_7150# a_33086_7150# 0.26fF
C4981 a_25054_16186# col_n[22] 0.28fF
C4982 a_33086_14178# rowon_n[12] 0.14fF
C4983 a_1962_11206# a_14010_11166# 0.27fF
C4984 a_26058_3134# col[23] 0.29fF
C4985 a_1962_1166# col[5] 0.11fF
C4986 a_17022_16186# a_18026_16186# 0.97fF
C4987 a_3270_7190# vcm 0.22fF
C4988 a_2346_16228# a_32994_16186# 0.35fF
C4989 a_1962_14218# col[7] 0.11fF
C4990 m2_1732_5966# rowoff_n[4] 0.12fF
C4991 a_23046_17190# vcm 0.60fF
C4992 m2_13780_18014# VDD 0.93fF
C4993 a_1962_18234# m2_28840_18014# 0.18fF
C4994 a_2966_11166# ctop 3.42fF
C4995 a_26058_10162# VDD 0.52fF
C4996 a_5886_8154# a_5978_8154# 0.26fF
C4997 a_2346_8196# a_8990_8154# 0.19fF
C4998 a_1962_8194# a_7286_8194# 0.14fF
C4999 a_10998_14178# row_n[12] 0.17fF
C5000 a_2346_13216# col[27] 0.15fF
C5001 a_1962_13214# a_27062_13174# 0.27fF
C5002 a_33086_2130# vcm 0.62fF
C5003 a_25054_12170# rowoff_n[10] 0.10fF
C5004 a_16322_11206# vcm 0.22fF
C5005 a_26058_4138# row_n[2] 0.17fF
C5006 a_12002_4138# rowoff_n[2] 0.10fF
C5007 a_2874_5142# a_2966_5142# 0.26fF
C5008 a_2346_5184# a_3878_5142# 0.35fF
C5009 a_7986_9158# col_n[5] 0.28fF
C5010 a_34090_7150# m3_34996_7102# 0.13fF
C5011 a_2346_18236# m2_23820_18014# 0.19fF
C5012 a_5886_13174# VDD 0.23fF
C5013 a_1962_10202# a_20338_10202# 0.14fF
C5014 a_29070_11166# a_29070_10162# 1.00fF
C5015 a_2346_10204# a_22042_10162# 0.19fF
C5016 a_22042_2130# rowoff_n[0] 0.10fF
C5017 a_29374_15222# vcm 0.22fF
C5018 a_26058_5142# col_n[23] 0.28fF
C5019 a_1962_3174# col_n[5] 0.13fF
C5020 col_n[12] ctop 2.02fF
C5021 col_n[21] row_n[3] 0.23fF
C5022 col_n[25] row_n[5] 0.23fF
C5023 col_n[31] row_n[8] 0.23fF
C5024 col_n[15] row_n[0] 0.22fF
C5025 col_n[27] row_n[6] 0.23fF
C5026 col_n[19] row_n[2] 0.23fF
C5027 vcm col[6] 5.84fF
C5028 col_n[23] row_n[4] 0.23fF
C5029 col_n[3] col[3] 0.72fF
C5030 col_n[17] row_n[1] 0.23fF
C5031 VDD col[10] 4.17fF
C5032 rowon_n[12] rowon_n[11] 0.15fF
C5033 col_n[29] row_n[7] 0.23fF
C5034 a_10998_9158# ctop 3.58fF
C5035 a_1962_16226# col_n[7] 0.13fF
C5036 a_30074_17190# row_n[15] 0.17fF
C5037 m2_11772_18014# m3_10900_18146# 0.13fF
C5038 a_13006_15182# m2_13204_15430# 0.16fF
C5039 a_14010_2130# rowon_n[0] 0.14fF
C5040 a_18938_17190# VDD 0.24fF
C5041 a_1962_12210# a_33390_12210# 0.14fF
C5042 a_18938_12170# a_19030_12170# 0.26fF
C5043 a_15014_3134# m2_15212_3382# 0.16fF
C5044 a_28978_2130# VDD 0.23fF
C5045 a_2346_4180# a_11910_4138# 0.35fF
C5046 a_24050_13174# ctop 3.58fF
C5047 m3_34996_5094# m3_34996_4090# 0.22fF
C5048 a_2346_9200# col[18] 0.15fF
C5049 a_10906_10162# rowoff_n[8] 0.24fF
C5050 a_18026_15182# rowon_n[13] 0.14fF
C5051 a_1962_18234# col_n[17] 0.13fF
C5052 a_4974_12170# vcm 0.62fF
C5053 a_12914_13174# rowoff_n[11] 0.24fF
C5054 m2_1732_10986# m3_1864_12122# 0.15fF
C5055 a_7986_5142# VDD 0.52fF
C5056 a_5978_12170# col[3] 0.29fF
C5057 a_33086_5142# rowon_n[3] 0.14fF
C5058 a_13006_6146# a_14010_6146# 0.97fF
C5059 a_2346_6188# a_24962_6146# 0.35fF
C5060 a_20946_8154# rowoff_n[6] 0.24fF
C5061 a_1962_5182# col[25] 0.11fF
C5062 a_31990_16186# a_32082_16186# 0.26fF
C5063 a_15014_16186# a_15014_15182# 1.00fF
C5064 a_18026_16186# vcm 0.62fF
C5065 a_26970_17190# rowoff_n[15] 0.24fF
C5066 a_24050_8154# col[21] 0.29fF
C5067 m2_34864_16006# VDD 1.00fF
C5068 a_1962_3174# a_19030_3134# 0.27fF
C5069 a_10998_5142# row_n[3] 0.17fF
C5070 a_30986_6146# rowoff_n[4] 0.24fF
C5071 a_1962_12210# sample 0.14fF
C5072 a_21038_9158# VDD 0.52fF
C5073 a_2966_8154# a_2966_7150# 1.00fF
C5074 a_9994_16186# m2_10192_16434# 0.16fF
C5075 a_28066_1126# vcm 0.12fF
C5076 a_2346_17232# a_6982_17190# 0.19fF
C5077 a_1962_17230# a_5278_17230# 0.14fF
C5078 a_4882_17190# a_4974_17190# 0.26fF
C5079 a_11302_10202# vcm 0.22fF
C5080 a_12002_4138# m2_12200_4386# 0.16fF
C5081 m3_5880_18146# ctop 0.23fF
C5082 a_1962_5182# a_32082_5142# 0.27fF
C5083 a_2346_5184# col[9] 0.15fF
C5084 a_34090_13174# VDD 0.54fF
C5085 a_26058_10162# a_27062_10162# 0.97fF
C5086 col[12] rowoff_n[1] 0.11fF
C5087 col[14] rowoff_n[3] 0.11fF
C5088 col[16] rowoff_n[5] 0.11fF
C5089 col[15] rowoff_n[4] 0.11fF
C5090 col[13] rowoff_n[2] 0.11fF
C5091 col[17] rowoff_n[6] 0.11fF
C5092 col[18] rowoff_n[7] 0.11fF
C5093 col[11] rowoff_n[0] 0.11fF
C5094 col[19] rowoff_n[8] 0.11fF
C5095 col[20] rowoff_n[9] 0.11fF
C5096 a_5978_14178# col_n[3] 0.28fF
C5097 a_1962_7190# col_n[25] 0.13fF
C5098 a_30074_8154# row_n[6] 0.17fF
C5099 m2_1732_12994# ctop 0.17fF
C5100 a_24354_14218# vcm 0.22fF
C5101 a_14922_2130# a_15014_2130# 0.26fF
C5102 a_1962_2170# a_25358_2170# 0.14fF
C5103 a_2346_2172# a_27062_2130# 0.19fF
C5104 a_5978_8154# ctop 3.58fF
C5105 a_24050_10162# col_n[21] 0.28fF
C5106 a_1962_1166# col[16] 0.11fF
C5107 a_13918_16186# VDD 0.23fF
C5108 a_1962_14218# col[18] 0.11fF
C5109 a_3970_2130# m2_2736_1950# 0.96fF
C5110 a_23958_1126# VDD 0.44fF
C5111 a_19030_12170# ctop 3.58fF
C5112 col[4] rowoff_n[10] 0.11fF
C5113 a_6982_17190# m2_7180_17438# 0.16fF
C5114 a_18026_6146# rowon_n[4] 0.14fF
C5115 a_2346_13216# a_9902_13174# 0.35fF
C5116 a_1962_1166# a_33390_1166# 0.14fF
C5117 a_2346_5184# m2_34864_4962# 0.17fF
C5118 a_8990_5142# m2_9188_5390# 0.16fF
C5119 m2_1732_7974# m3_1864_9110# 0.15fF
C5120 a_2874_4138# VDD 0.24fF
C5121 a_6982_3134# col_n[4] 0.28fF
C5122 m3_1864_12122# VDD 0.25fF
C5123 a_10998_6146# a_10998_5142# 1.00fF
C5124 a_27974_6146# a_28066_6146# 0.26fF
C5125 a_2346_1168# col[0] 0.15fF
C5126 a_32082_16186# ctop 3.57fF
C5127 a_2346_14220# col[2] 0.15fF
C5128 a_1962_10202# a_3970_10162# 0.27fF
C5129 a_3970_17190# col[1] 0.29fF
C5130 a_2346_15224# a_22954_15182# 0.35fF
C5131 a_12002_15182# a_13006_15182# 0.97fF
C5132 a_1962_3174# col_n[16] 0.13fF
C5133 vcm col[17] 5.84fF
C5134 col_n[30] row_n[2] 0.23fF
C5135 VDD col[21] 4.18fF
C5136 col_n[26] row_n[0] 0.23fF
C5137 col_n[28] row_n[1] 0.23fF
C5138 col_n[23] ctop 2.02fF
C5139 col_n[8] col[9] 5.98fF
C5140 rowon_n[9] row_n[9] 19.75fF
C5141 a_1962_16226# col_n[18] 0.13fF
C5142 a_13006_15182# vcm 0.62fF
C5143 a_16018_8154# VDD 0.52fF
C5144 a_22042_13174# col[19] 0.29fF
C5145 a_1962_10202# col[9] 0.11fF
C5146 a_1962_12210# a_17022_12170# 0.27fF
C5147 a_6282_9198# vcm 0.22fF
C5148 m2_20808_946# col_n[18] 0.37fF
C5149 a_2346_9200# col[29] 0.15fF
C5150 a_15014_9158# row_n[7] 0.17fF
C5151 a_29070_12170# VDD 0.52fF
C5152 m3_25960_18146# m3_26964_18146# 0.22fF
C5153 a_1962_9198# a_10298_9198# 0.14fF
C5154 a_24050_10162# a_24050_9158# 1.00fF
C5155 a_2346_9200# a_12002_9158# 0.19fF
C5156 a_1962_18234# col_n[28] 0.13fF
C5157 a_1962_11206# row_n[9] 25.57fF
C5158 a_2346_3176# vcm 0.40fF
C5159 a_1962_14218# a_30074_14178# 0.27fF
C5160 a_13918_3134# rowoff_n[1] 0.24fF
C5161 a_28978_14178# rowoff_n[12] 0.24fF
C5162 a_19334_13214# vcm 0.22fF
C5163 a_5978_6146# m2_6176_6394# 0.16fF
C5164 a_4974_6146# col[2] 0.29fF
C5165 a_8898_15182# VDD 0.23fF
C5166 a_2346_11208# a_25054_11166# 0.19fF
C5167 a_13918_11166# a_14010_11166# 0.26fF
C5168 a_1962_11206# a_23350_11206# 0.14fF
C5169 a_22042_15182# col_n[19] 0.28fF
C5170 a_1962_12210# col_n[9] 0.13fF
C5171 a_34090_12170# row_n[10] 0.17fF
C5172 a_32386_17230# vcm 0.22fF
C5173 a_23046_2130# col[20] 0.29fF
C5174 a_14010_11166# ctop 3.58fF
C5175 a_2966_9158# VDD 0.56fF
C5176 a_1962_6186# col[0] 0.11fF
C5177 m2_1732_4962# m3_1864_6098# 0.15fF
C5178 a_2346_5184# col[20] 0.15fF
C5179 a_31990_4138# VDD 0.23fF
C5180 a_7986_5142# a_8990_5142# 0.97fF
C5181 a_2346_5184# a_14922_5142# 0.35fF
C5182 col[26] rowoff_n[4] 0.11fF
C5183 col[25] rowoff_n[3] 0.11fF
C5184 col[31] rowoff_n[9] 0.11fF
C5185 col[24] rowoff_n[2] 0.11fF
C5186 col[23] rowoff_n[1] 0.11fF
C5187 col[29] rowoff_n[7] 0.11fF
C5188 col[30] rowoff_n[8] 0.11fF
C5189 col[22] rowoff_n[0] 0.11fF
C5190 col[27] rowoff_n[5] 0.11fF
C5191 col[28] rowoff_n[6] 0.11fF
C5192 a_27062_15182# ctop 3.58fF
C5193 a_22042_10162# rowon_n[8] 0.14fF
C5194 a_34090_16186# m3_34996_16138# 0.13fF
C5195 a_4974_8154# col_n[2] 0.28fF
C5196 a_12002_9158# rowoff_n[7] 0.10fF
C5197 a_26970_15182# a_27062_15182# 0.26fF
C5198 a_9994_15182# a_9994_14178# 1.00fF
C5199 a_7986_14178# vcm 0.62fF
C5200 a_16018_15182# rowoff_n[13] 0.10fF
C5201 a_1962_2170# a_8990_2130# 0.27fF
C5202 a_1962_1166# col[27] 0.11fF
C5203 m2_25828_18014# m3_25960_18146# 2.78fF
C5204 a_10998_7150# VDD 0.52fF
C5205 a_1962_14218# col[29] 0.11fF
C5206 a_22042_7150# rowoff_n[5] 0.10fF
C5207 a_2346_7192# a_27974_7150# 0.35fF
C5208 a_23046_4138# col_n[20] 0.28fF
C5209 a_1962_8194# vcm 6.95fF
C5210 a_32082_5142# rowoff_n[3] 0.10fF
C5211 a_21038_18194# vcm 0.12fF
C5212 col[15] rowoff_n[10] 0.11fF
C5213 a_1962_4178# a_22042_4138# 0.27fF
C5214 a_24050_11166# VDD 0.52fF
C5215 a_1962_2170# row_n[0] 25.57fF
C5216 m3_15920_1078# m3_16924_1078# 0.22fF
C5217 a_21038_9158# a_22042_9158# 0.97fF
C5218 a_31078_3134# vcm 0.62fF
C5219 a_14314_12210# vcm 0.22fF
C5220 a_1962_1166# a_15318_1166# 0.14fF
C5221 a_2346_1168# col[11] 0.14fF
C5222 a_2346_14220# col[13] 0.15fF
C5223 a_19030_13174# row_n[11] 0.17fF
C5224 m2_34864_5966# vcm 0.51fF
C5225 a_1962_3174# col_n[27] 0.13fF
C5226 a_34090_3134# row_n[1] 0.17fF
C5227 vcm col[28] 5.84fF
C5228 a_1962_16226# col_n[29] 0.13fF
C5229 VDD rowoff_n[15] 1.22fF
C5230 rowon_n[14] ctop 1.40fF
C5231 col_n[14] col[14] 0.72fF
C5232 a_2966_15182# a_3970_15182# 0.97fF
C5233 a_27366_16226# vcm 0.22fF
C5234 m2_12776_946# m2_13780_946# 0.96fF
C5235 a_1962_3174# a_28370_3174# 0.14fF
C5236 a_2346_3176# a_30074_3134# 0.19fF
C5237 a_33086_4138# a_33086_3134# 1.00fF
C5238 a_34090_9158# m2_34288_9406# 0.16fF
C5239 a_1962_10202# col[20] 0.11fF
C5240 a_8990_10162# ctop 3.58fF
C5241 a_21038_7150# col[18] 0.29fF
C5242 a_16930_18194# VDD 0.33fF
C5243 m2_8760_18014# vcm 0.28fF
C5244 a_6982_11166# rowon_n[9] 0.14fF
C5245 a_30986_11166# rowoff_n[9] 0.24fF
C5246 m2_1732_1950# m3_1864_3086# 0.15fF
C5247 a_26970_3134# VDD 0.23fF
C5248 m3_34996_11118# ctop 0.23fF
C5249 a_5978_5142# a_5978_4138# 1.00fF
C5250 a_22954_5142# a_23046_5142# 0.26fF
C5251 a_22042_14178# ctop 3.58fF
C5252 m2_29844_946# m2_30848_946# 0.96fF
C5253 a_6982_14178# a_7986_14178# 0.97fF
C5254 a_2346_14220# a_12914_14178# 0.35fF
C5255 a_2346_18236# a_21950_18194# 0.35fF
C5256 a_2346_10204# col[4] 0.15fF
C5257 a_5978_6146# VDD 0.52fF
C5258 a_26058_14178# rowon_n[12] 0.14fF
C5259 a_1962_11206# a_6982_11166# 0.27fF
C5260 a_1962_12210# col_n[20] 0.13fF
C5261 a_21038_9158# col_n[18] 0.28fF
C5262 a_2346_16228# a_25966_16186# 0.35fF
C5263 m2_1732_7974# sample_n 0.15fF
C5264 a_16018_17190# vcm 0.60fF
C5265 a_35494_1488# VDD 0.12fF
C5266 a_31078_10162# m2_31276_10410# 0.16fF
C5267 a_1962_6186# col[11] 0.11fF
C5268 a_1962_18234# m2_14784_18014# 0.18fF
C5269 a_19030_10162# VDD 0.52fF
C5270 a_19030_9158# a_19030_8154# 1.00fF
C5271 a_3970_14178# row_n[12] 0.17fF
C5272 a_26058_2130# vcm 0.62fF
C5273 a_1962_13214# a_20034_13174# 0.27fF
C5274 a_2966_16186# col[0] 0.29fF
C5275 a_2346_5184# col[31] 0.15fF
C5276 a_19030_4138# row_n[2] 0.17fF
C5277 a_4974_4138# rowoff_n[2] 0.10fF
C5278 a_18026_12170# rowoff_n[10] 0.10fF
C5279 a_9294_11206# vcm 0.22fF
C5280 a_2346_12212# m2_1732_11990# 0.12fF
C5281 m3_21944_1078# VDD 0.14fF
C5282 a_32082_14178# VDD 0.52fF
C5283 a_2346_18236# m2_9764_18014# 0.19fF
C5284 a_2346_10204# a_15014_10162# 0.19fF
C5285 a_1962_10202# a_13310_10202# 0.14fF
C5286 a_8898_10162# a_8990_10162# 0.26fF
C5287 a_3970_2130# col_n[1] 0.26fF
C5288 a_15014_2130# rowoff_n[0] 0.10fF
C5289 a_1962_15222# a_33086_15182# 0.27fF
C5290 a_22346_15222# vcm 0.22fF
C5291 a_32082_16186# rowoff_n[14] 0.10fF
C5292 a_30074_3134# a_31078_3134# 0.97fF
C5293 a_3970_9158# ctop 3.57fF
C5294 a_23046_17190# row_n[15] 0.17fF
C5295 m2_1732_18014# m3_2868_18146# 0.13fF
C5296 m2_34864_15002# row_n[13] 0.15fF
C5297 a_11910_17190# VDD 0.24fF
C5298 a_6982_2130# rowon_n[0] 0.14fF
C5299 a_1962_8194# col_n[11] 0.13fF
C5300 a_2346_12212# a_28066_12170# 0.19fF
C5301 a_1962_12210# a_26362_12210# 0.14fF
C5302 a_32082_13174# a_32082_12170# 1.00fF
C5303 a_19030_12170# col[16] 0.29fF
C5304 m2_17796_18014# col_n[15] 0.25fF
C5305 col[26] rowoff_n[10] 0.11fF
C5306 m2_1732_16006# m2_2160_16434# 0.16fF
C5307 a_21950_2130# VDD 0.23fF
C5308 a_1962_2170# col[2] 0.11fF
C5309 a_28066_11166# m2_28264_11414# 0.16fF
C5310 a_2346_4180# a_4882_4138# 0.35fF
C5311 a_1962_15222# col[4] 0.11fF
C5312 a_17022_13174# ctop 3.58fF
C5313 m3_34996_12122# m3_34996_11118# 0.22fF
C5314 m2_32856_946# m3_32988_1078# 2.79fF
C5315 a_21950_14178# a_22042_14178# 0.26fF
C5316 a_4974_14178# a_4974_13174# 1.00fF
C5317 a_2346_1168# col[22] 0.14fF
C5318 a_10998_15182# rowon_n[13] 0.14fF
C5319 a_2346_14220# col[24] 0.15fF
C5320 a_5886_13174# rowoff_n[11] 0.24fF
C5321 a_35002_6146# VDD 0.29fF
C5322 a_26058_5142# rowon_n[3] 0.14fF
C5323 a_2346_6188# a_17934_6146# 0.35fF
C5324 col_n[19] col[20] 5.98fF
C5325 row_n[9] ctop 1.65fF
C5326 a_30074_17190# ctop 3.39fF
C5327 a_13918_8154# rowoff_n[6] 0.24fF
C5328 a_1962_11206# a_34394_11206# 0.14fF
C5329 m2_21812_946# a_22042_2130# 0.99fF
C5330 col[10] rowoff_n[11] 0.11fF
C5331 m2_7756_946# col_n[5] 0.37fF
C5332 a_1962_10202# col[31] 0.11fF
C5333 a_19942_17190# rowoff_n[15] 0.24fF
C5334 a_10998_16186# vcm 0.62fF
C5335 a_19030_14178# col_n[16] 0.28fF
C5336 a_1962_3174# a_12002_3134# 0.27fF
C5337 a_23958_6146# rowoff_n[4] 0.24fF
C5338 a_3970_5142# row_n[3] 0.17fF
C5339 a_14010_9158# VDD 0.52fF
C5340 a_20034_1126# col[17] 0.38fF
C5341 a_16018_8154# a_17022_8154# 0.97fF
C5342 a_2346_8196# a_30986_8154# 0.35fF
C5343 a_1962_4178# col_n[2] 0.13fF
C5344 a_1962_17230# col_n[4] 0.13fF
C5345 a_21038_1126# vcm 0.12fF
C5346 m2_1732_946# m2_2160_1374# 0.16fF
C5347 a_33998_4138# rowoff_n[2] 0.24fF
C5348 a_4274_10202# vcm 0.22fF
C5349 m2_23820_946# ctop 0.18fF
C5350 a_1962_5182# a_25054_5142# 0.27fF
C5351 a_25054_12170# m2_25252_12418# 0.16fF
C5352 a_27062_13174# VDD 0.52fF
C5353 ctop rowoff_n[12] 0.60fF
C5354 a_34090_5142# vcm 0.62fF
C5355 a_2346_10204# col[15] 0.15fF
C5356 a_23046_8154# row_n[6] 0.17fF
C5357 a_17326_14218# vcm 0.22fF
C5358 a_28066_3134# a_28066_2130# 1.00fF
C5359 a_2346_2172# a_20034_2130# 0.19fF
C5360 a_1962_2170# a_18330_2170# 0.14fF
C5361 a_1962_12210# col_n[31] 0.13fF
C5362 a_6890_16186# VDD 0.23fF
C5363 m2_1732_15002# rowoff_n[13] 0.12fF
C5364 a_29070_12170# a_30074_12170# 0.97fF
C5365 a_20034_3134# col_n[17] 0.28fF
C5366 a_1962_6186# col[22] 0.11fF
C5367 a_30378_18234# vcm 0.22fF
C5368 a_16930_1126# VDD 0.44fF
C5369 a_17022_17190# col[14] 0.29fF
C5370 a_2346_4180# a_33086_4138# 0.19fF
C5371 a_1962_4178# a_31382_4178# 0.14fF
C5372 a_17934_4138# a_18026_4138# 0.26fF
C5373 a_12002_12170# ctop 3.58fF
C5374 a_13006_17190# m2_12776_18014# 1.00fF
C5375 a_10998_6146# rowon_n[4] 0.14fF
C5376 a_32082_10162# rowoff_n[8] 0.10fF
C5377 a_34090_13174# rowoff_n[11] 0.10fF
C5378 a_29982_5142# VDD 0.23fF
C5379 m3_17928_18146# VDD 0.25fF
C5380 a_22042_13174# m2_22240_13422# 0.16fF
C5381 a_25054_16186# ctop 3.57fF
C5382 a_2346_6188# col[6] 0.15fF
C5383 a_2346_15224# a_15926_15182# 0.35fF
C5384 a_5978_15182# vcm 0.62fF
C5385 a_28066_2130# m3_27968_1078# 0.15fF
C5386 a_8990_8154# VDD 0.52fF
C5387 a_30074_9158# rowon_n[7] 0.14fF
C5388 a_1962_8194# col_n[22] 0.13fF
C5389 rowon_n[14] rowoff_n[14] 20.27fF
C5390 a_14010_8154# a_14010_7150# 1.00fF
C5391 a_30986_8154# a_31078_8154# 0.26fF
C5392 a_1962_12210# a_9994_12170# 0.27fF
C5393 a_1962_18234# a_33390_18234# 0.14fF
C5394 a_18026_6146# col[15] 0.29fF
C5395 a_1962_2170# col[13] 0.11fF
C5396 a_2346_17232# a_28978_17190# 0.35fF
C5397 a_15014_17190# a_16018_17190# 0.97fF
C5398 a_1962_15222# col[15] 0.11fF
C5399 m2_1732_946# m3_2868_1078# 0.13fF
C5400 a_3878_2130# VDD 0.23fF
C5401 m3_24956_1078# ctop 0.23fF
C5402 a_7986_9158# row_n[7] 0.17fF
C5403 a_22042_12170# VDD 0.52fF
C5404 m3_11904_18146# m3_12908_18146# 0.22fF
C5405 a_2346_9200# a_4974_9158# 0.19fF
C5406 a_1962_9198# a_3270_9198# 0.14fF
C5407 a_29070_4138# vcm 0.62fF
C5408 a_1962_14218# a_23046_14178# 0.27fF
C5409 a_6890_3134# rowoff_n[1] 0.24fF
C5410 a_2346_18236# col[7] 0.14fF
C5411 a_12306_13214# vcm 0.22fF
C5412 a_21950_14178# rowoff_n[12] 0.24fF
C5413 a_25054_2130# a_26058_2130# 0.97fF
C5414 rowon_n[3] ctop 1.40fF
C5415 rowon_n[1] rowon_n[0] 0.15fF
C5416 col_n[25] col[25] 0.78fF
C5417 a_19030_14178# m2_19228_14426# 0.16fF
C5418 col[21] rowoff_n[11] 0.11fF
C5419 a_1962_11206# a_16322_11206# 0.14fF
C5420 m2_1732_8978# vcm 0.45fF
C5421 a_2346_11208# a_18026_11166# 0.19fF
C5422 a_27062_12170# a_27062_11166# 1.00fF
C5423 a_27062_12170# row_n[10] 0.17fF
C5424 a_25358_17230# vcm 0.22fF
C5425 a_18026_8154# col_n[15] 0.28fF
C5426 a_1962_4178# col_n[13] 0.13fF
C5427 a_6982_11166# ctop 3.58fF
C5428 a_1962_17230# col_n[15] 0.13fF
C5429 a_32082_17190# m2_31852_18014# 1.00fF
C5430 a_2966_1126# vcm 0.12fF
C5431 a_2346_13216# a_31078_13174# 0.19fF
C5432 a_1962_13214# a_29374_13214# 0.14fF
C5433 a_16930_13174# a_17022_13174# 0.26fF
C5434 a_1962_11206# col[6] 0.11fF
C5435 a_2346_16228# row_n[14] 0.35fF
C5436 a_24962_4138# VDD 0.23fF
C5437 a_2346_5184# a_7894_5142# 0.35fF
C5438 col[5] rowoff_n[12] 0.11fF
C5439 a_20034_15182# ctop 3.58fF
C5440 a_15014_10162# rowon_n[8] 0.14fF
C5441 a_2346_10204# col[26] 0.15fF
C5442 a_4974_9158# rowoff_n[7] 0.10fF
C5443 a_8990_15182# rowoff_n[13] 0.10fF
C5444 a_1962_12210# rowon_n[10] 1.18fF
C5445 m2_16792_18014# m3_15920_18146# 0.13fF
C5446 a_3970_7150# VDD 0.52fF
C5447 a_15014_7150# rowoff_n[5] 0.10fF
C5448 a_16018_15182# m2_16216_15430# 0.16fF
C5449 a_10998_7150# a_12002_7150# 0.97fF
C5450 a_2346_7192# a_20946_7150# 0.35fF
C5451 a_29982_17190# a_30074_17190# 0.26fF
C5452 a_13006_17190# a_13006_16186# 1.00fF
C5453 a_18026_3134# m2_18224_3382# 0.16fF
C5454 a_25054_5142# rowoff_n[3] 0.10fF
C5455 a_16018_11166# col[13] 0.29fF
C5456 a_14010_18194# vcm 0.12fF
C5457 a_1962_4178# a_15014_4138# 0.27fF
C5458 a_1962_13214# col_n[6] 0.13fF
C5459 a_34090_13174# rowon_n[11] 0.14fF
C5460 a_17022_11166# VDD 0.52fF
C5461 m3_1864_1078# m3_2868_1078# 0.22fF
C5462 a_2346_9200# a_33998_9158# 0.35fF
C5463 a_24050_3134# vcm 0.62fF
C5464 m2_32856_18014# col[30] 0.28fF
C5465 a_34090_7150# col[31] 0.29fF
C5466 a_7286_12210# vcm 0.22fF
C5467 a_1962_1166# a_8290_1166# 0.14fF
C5468 a_12002_13174# row_n[11] 0.17fF
C5469 a_1962_6186# a_28066_6146# 0.27fF
C5470 a_30074_15182# VDD 0.52fF
C5471 a_2346_6188# col[17] 0.15fF
C5472 a_24050_11166# a_25054_11166# 0.97fF
C5473 m2_13780_946# a_2346_1168# 0.19fF
C5474 a_27062_3134# row_n[1] 0.17fF
C5475 a_8898_1126# m2_8760_946# 0.16fF
C5476 a_20338_16226# vcm 0.22fF
C5477 a_2346_3176# a_23046_3134# 0.19fF
C5478 a_12914_3134# a_13006_3134# 0.26fF
C5479 a_1962_3174# a_21342_3174# 0.14fF
C5480 a_2346_1168# m2_30848_946# 0.19fF
C5481 a_13006_16186# m2_13204_16434# 0.16fF
C5482 a_16018_13174# col_n[13] 0.28fF
C5483 a_9902_18194# VDD 0.33fF
C5484 a_1962_2170# col[24] 0.11fF
C5485 a_30378_1166# vcm 0.23fF
C5486 a_2346_7192# row_n[5] 0.35fF
C5487 a_1962_15222# col[26] 0.11fF
C5488 a_23958_11166# rowoff_n[9] 0.24fF
C5489 a_31078_16186# row_n[14] 0.17fF
C5490 a_15014_4138# m2_15212_4386# 0.16fF
C5491 a_19942_3134# VDD 0.23fF
C5492 m3_20940_18146# ctop 0.23fF
C5493 a_34090_9158# col_n[31] 0.28fF
C5494 a_2346_5184# a_2346_4180# 0.22fF
C5495 a_1962_5182# a_35398_5182# 0.14fF
C5496 a_15014_14178# ctop 3.58fF
C5497 a_33998_9158# rowoff_n[7] 0.24fF
C5498 a_2346_18236# col[18] 0.14fF
C5499 a_2346_14220# a_5886_14178# 0.35fF
C5500 a_1962_3174# rowon_n[1] 1.18fF
C5501 col_n[30] col[31] 6.04fF
C5502 a_2346_18236# a_14922_18194# 0.35fF
C5503 m2_34864_17010# rowon_n[15] 0.13fF
C5504 a_3878_14178# rowoff_n[12] 0.24fF
C5505 a_32994_7150# VDD 0.23fF
C5506 a_8990_7150# a_8990_6146# 1.00fF
C5507 a_25966_7150# a_26058_7150# 0.26fF
C5508 a_2346_2172# col[8] 0.15fF
C5509 a_2346_15224# col[10] 0.15fF
C5510 a_19030_14178# rowon_n[12] 0.14fF
C5511 a_2346_16228# a_18938_16186# 0.35fF
C5512 a_9994_16186# a_10998_16186# 0.97fF
C5513 a_1962_4178# col_n[24] 0.13fF
C5514 a_34090_4138# rowon_n[2] 0.14fF
C5515 a_1962_17230# col_n[26] 0.13fF
C5516 a_17022_2130# col_n[14] 0.28fF
C5517 a_8990_17190# vcm 0.60fF
C5518 a_12002_10162# VDD 0.52fF
C5519 a_14010_16186# col[11] 0.29fF
C5520 a_9994_17190# m2_10192_17438# 0.16fF
C5521 a_1962_18234# col[0] 0.11fF
C5522 a_1962_11206# col[17] 0.11fF
C5523 a_1962_13214# a_13006_13174# 0.27fF
C5524 a_19030_2130# vcm 0.62fF
C5525 a_10998_12170# rowoff_n[10] 0.10fF
C5526 a_12002_4138# row_n[2] 0.17fF
C5527 col[16] rowoff_n[12] 0.11fF
C5528 a_12002_5142# m2_12200_5390# 0.16fF
C5529 a_32082_12170# col[29] 0.29fF
C5530 m3_34996_5094# VDD 0.26fF
C5531 a_25054_14178# VDD 0.52fF
C5532 a_1962_10202# a_6282_10202# 0.14fF
C5533 a_22042_11166# a_22042_10162# 1.00fF
C5534 a_2346_10204# a_7986_10162# 0.19fF
C5535 a_7986_2130# rowoff_n[0] 0.10fF
C5536 a_32082_6146# vcm 0.62fF
C5537 a_1962_15222# a_26058_15182# 0.27fF
C5538 m2_22816_18014# ctop 0.18fF
C5539 a_25054_16186# rowoff_n[14] 0.10fF
C5540 a_15318_15222# vcm 0.22fF
C5541 a_16018_17190# row_n[15] 0.17fF
C5542 a_2346_7192# a_1962_7190# 2.62fF
C5543 a_2346_11208# col[1] 0.15fF
C5544 a_4882_17190# VDD 0.24fF
C5545 a_2346_12212# a_21038_12170# 0.19fF
C5546 a_1962_12210# a_19334_12210# 0.14fF
C5547 a_11910_12170# a_12002_12170# 0.26fF
C5548 a_31078_7150# row_n[5] 0.17fF
C5549 m2_11772_946# m3_12908_1078# 0.13fF
C5550 col[0] rowoff_n[13] 0.11fF
C5551 a_1962_13214# col_n[17] 0.13fF
C5552 a_15014_5142# col[12] 0.29fF
C5553 a_14922_2130# VDD 0.23fF
C5554 a_33086_5142# a_34090_5142# 0.97fF
C5555 a_9994_13174# ctop 3.58fF
C5556 m2_23820_946# m3_22948_1078# 0.13fF
C5557 a_11910_18194# m2_11772_18014# 0.16fF
C5558 a_1962_7190# col[8] 0.11fF
C5559 a_32082_14178# col_n[29] 0.28fF
C5560 a_2346_14220# a_34090_14178# 0.19fF
C5561 a_1962_14218# a_32386_14218# 0.14fF
C5562 a_3970_15182# rowon_n[13] 0.14fF
C5563 m2_1732_5966# m2_1732_4962# 0.99fF
C5564 a_8990_6146# m2_9188_6394# 0.16fF
C5565 a_2346_6188# m2_34864_5966# 0.17fF
C5566 a_27974_6146# VDD 0.23fF
C5567 a_2346_6188# col[28] 0.15fF
C5568 a_19030_5142# rowon_n[3] 0.14fF
C5569 a_2346_6188# a_10906_6146# 0.35fF
C5570 a_5978_6146# a_6982_6146# 0.97fF
C5571 a_23046_17190# ctop 3.39fF
C5572 a_6890_8154# rowoff_n[6] 0.24fF
C5573 a_4974_17190# m3_4876_18146# 0.15fF
C5574 a_24962_16186# a_25054_16186# 0.26fF
C5575 a_7986_16186# a_7986_15182# 1.00fF
C5576 a_33086_2130# ctop 3.38fF
C5577 a_12914_17190# rowoff_n[15] 0.24fF
C5578 a_3970_16186# vcm 0.62fF
C5579 a_3878_3134# a_3970_3134# 0.26fF
C5580 a_1962_3174# a_4974_3134# 0.27fF
C5581 a_16930_6146# rowoff_n[4] 0.24fF
C5582 a_6982_9158# VDD 0.52fF
C5583 a_2346_8196# a_23958_8154# 0.35fF
C5584 a_15014_7150# col_n[12] 0.28fF
C5585 m2_30848_946# col_n[28] 0.46fF
C5586 a_14010_1126# vcm 0.12fF
C5587 a_26970_4138# rowoff_n[2] 0.24fF
C5588 a_1962_9198# col_n[8] 0.13fF
C5589 a_35494_4500# VDD 0.11fF
C5590 a_33086_3134# col_n[30] 0.28fF
C5591 a_1962_5182# a_18026_5142# 0.27fF
C5592 a_2346_18236# col[29] 0.14fF
C5593 a_20034_13174# VDD 0.52fF
C5594 a_1962_10202# a_1962_9198# 0.16fF
C5595 a_19030_10162# a_20034_10162# 0.97fF
C5596 ctop col[6] 1.98fF
C5597 a_30074_17190# col[27] 0.29fF
C5598 a_1962_16226# col[1] 0.11fF
C5599 a_27062_5142# vcm 0.62fF
C5600 a_16018_8154# row_n[6] 0.17fF
C5601 a_10298_14218# vcm 0.22fF
C5602 a_5978_7150# m2_6176_7398# 0.16fF
C5603 a_2346_2172# a_13006_2130# 0.19fF
C5604 a_1962_2170# a_11302_2170# 0.14fF
C5605 a_7894_2130# a_7986_2130# 0.26fF
C5606 a_2346_2172# col[19] 0.15fF
C5607 m2_30848_18014# m3_30980_18146# 2.78fF
C5608 a_2346_15224# col[21] 0.15fF
C5609 a_1962_7190# a_31078_7150# 0.27fF
C5610 a_33086_17190# VDD 0.55fF
C5611 a_23350_18234# vcm 0.22fF
C5612 a_9902_1126# VDD 0.44fF
C5613 a_1962_18234# col[11] 0.11fF
C5614 a_1962_4178# a_24354_4178# 0.14fF
C5615 a_31078_5142# a_31078_4138# 1.00fF
C5616 a_2346_4180# a_26058_4138# 0.19fF
C5617 a_4974_12170# ctop 3.58fF
C5618 a_1962_11206# col[28] 0.11fF
C5619 a_13006_10162# col[10] 0.29fF
C5620 a_30986_18194# m2_30848_18014# 0.16fF
C5621 a_3970_6146# rowon_n[4] 0.14fF
C5622 m2_12776_946# VDD 0.62fF
C5623 a_33390_3174# vcm 0.22fF
C5624 a_32082_14178# a_33086_14178# 0.97fF
C5625 a_25054_10162# rowoff_n[8] 0.10fF
C5626 col[27] rowoff_n[12] 0.11fF
C5627 a_1962_5182# col_n[0] 0.13fF
C5628 a_27062_13174# rowoff_n[11] 0.10fF
C5629 a_31078_6146# col[28] 0.29fF
C5630 a_22954_5142# VDD 0.23fF
C5631 m2_29844_946# VDD 0.62fF
C5632 a_20946_6146# a_21038_6146# 0.26fF
C5633 a_3970_6146# a_3970_5142# 1.00fF
C5634 a_18026_16186# ctop 3.57fF
C5635 a_4974_15182# a_5978_15182# 0.97fF
C5636 a_2346_15224# a_8898_15182# 0.35fF
C5637 m2_16792_946# m2_17220_1374# 0.16fF
C5638 a_2346_11208# col[12] 0.15fF
C5639 a_23046_9158# rowon_n[7] 0.14fF
C5640 col[11] rowoff_n[13] 0.11fF
C5641 a_2346_12212# a_2966_12170# 0.21fF
C5642 a_1962_18234# a_26362_18234# 0.14fF
C5643 a_1962_13214# col_n[28] 0.13fF
C5644 a_13006_12170# col_n[10] 0.28fF
C5645 a_2346_17232# a_21950_17190# 0.35fF
C5646 m2_28840_18014# m2_29844_18014# 0.96fF
C5647 m3_1864_3086# ctop 0.23fF
C5648 a_1962_7190# col[19] 0.11fF
C5649 a_15014_12170# VDD 0.52fF
C5650 m2_33860_946# m2_34864_946# 0.59fF
C5651 a_33998_10162# a_34090_10162# 0.26fF
C5652 a_17022_10162# a_17022_9158# 1.00fF
C5653 a_31078_8154# col_n[28] 0.28fF
C5654 a_22042_4138# vcm 0.62fF
C5655 a_1962_14218# a_16018_14178# 0.27fF
C5656 a_5278_13214# vcm 0.22fF
C5657 a_14922_14178# rowoff_n[12] 0.24fF
C5658 a_28066_16186# VDD 0.52fF
C5659 a_2346_11208# a_10998_11166# 0.19fF
C5660 a_6890_11166# a_6982_11166# 0.26fF
C5661 a_1962_11206# a_9294_11206# 0.14fF
C5662 a_1962_16226# a_29070_16186# 0.27fF
C5663 a_35094_8154# vcm 0.12fF
C5664 a_20034_12170# row_n[10] 0.17fF
C5665 a_18330_17230# vcm 0.22fF
C5666 a_2346_7192# col[3] 0.15fF
C5667 a_28066_4138# a_29070_4138# 0.97fF
C5668 a_34090_10162# m2_34288_10410# 0.16fF
C5669 a_2346_13216# a_24050_13174# 0.19fF
C5670 a_1962_13214# a_22346_13214# 0.14fF
C5671 a_30074_14178# a_30074_13174# 1.00fF
C5672 a_28370_2170# vcm 0.22fF
C5673 a_1962_9198# col_n[19] 0.13fF
C5674 a_10998_15182# col[8] 0.29fF
C5675 a_17934_4138# VDD 0.23fF
C5676 m2_34864_5966# row_n[4] 0.15fF
C5677 a_1962_3174# col[10] 0.11fF
C5678 ctop col[17] 2.02fF
C5679 col[5] col[6] 0.20fF
C5680 en_bit_n[1] col[15] 0.16fF
C5681 a_1962_16226# col[12] 0.11fF
C5682 a_13006_15182# ctop 3.58fF
C5683 a_29070_11166# col[26] 0.29fF
C5684 a_7986_10162# rowon_n[8] 0.14fF
C5685 a_19942_15182# a_20034_15182# 0.26fF
C5686 a_2346_2172# col[30] 0.15fF
C5687 m2_6752_18014# m3_7888_18146# 0.13fF
C5688 a_30986_8154# VDD 0.23fF
C5689 a_7986_7150# rowoff_n[5] 0.10fF
C5690 a_2346_7192# a_13918_7150# 0.35fF
C5691 a_1962_18234# col[22] 0.11fF
C5692 a_18026_5142# rowoff_n[3] 0.10fF
C5693 a_2346_3176# ctop 1.58fF
C5694 a_6982_18194# vcm 0.12fF
C5695 a_10998_17190# col_n[8] 0.28fF
C5696 a_1962_4178# a_7986_4138# 0.27fF
C5697 a_31078_11166# m2_31276_11414# 0.16fF
C5698 a_27062_13174# rowon_n[11] 0.14fF
C5699 a_12002_4138# col[9] 0.29fF
C5700 a_9994_11166# VDD 0.52fF
C5701 a_14010_9158# a_15014_9158# 0.97fF
C5702 a_2346_9200# a_26970_9158# 0.35fF
C5703 a_1962_5182# col_n[10] 0.13fF
C5704 a_17022_3134# vcm 0.62fF
C5705 a_22954_1126# m2_22816_946# 0.16fF
C5706 a_28066_3134# rowoff_n[1] 0.10fF
C5707 a_29070_13174# col_n[26] 0.28fF
C5708 a_2346_1168# a_2874_1126# 0.35fF
C5709 a_2966_15182# col_n[0] 0.28fF
C5710 a_4974_13174# row_n[11] 0.17fF
C5711 a_1962_12210# col[3] 0.11fF
C5712 a_2346_13216# m2_1732_12994# 0.12fF
C5713 a_1962_6186# a_21038_6146# 0.27fF
C5714 a_2346_17232# rowon_n[15] 0.26fF
C5715 a_23046_15182# VDD 0.52fF
C5716 a_20034_3134# row_n[1] 0.17fF
C5717 a_30074_7150# vcm 0.62fF
C5718 a_2346_1168# m2_6752_946# 0.19fF
C5719 a_2346_11208# col[23] 0.15fF
C5720 a_13310_16226# vcm 0.22fF
C5721 a_1962_3174# a_14314_3174# 0.14fF
C5722 a_2346_3176# a_16018_3134# 0.19fF
C5723 a_26058_4138# a_26058_3134# 1.00fF
C5724 col[22] rowoff_n[13] 0.11fF
C5725 a_1962_8194# a_34090_8154# 0.27fF
C5726 vcm rowoff_n[4] 0.20fF
C5727 a_23350_1166# vcm 0.23fF
C5728 sample_n rowoff_n[1] 0.38fF
C5729 VDD rowoff_n[0] 1.18fF
C5730 a_27062_13174# a_28066_13174# 0.97fF
C5731 a_12002_6146# col_n[9] 0.28fF
C5732 m2_5748_946# m2_6752_946# 0.96fF
C5733 a_2346_17232# a_3878_17190# 0.35fF
C5734 a_16930_11166# rowoff_n[9] 0.24fF
C5735 a_2874_17190# a_2966_17190# 0.26fF
C5736 a_24050_16186# row_n[14] 0.17fF
C5737 a_1962_7190# col[30] 0.11fF
C5738 a_12914_3134# VDD 0.23fF
C5739 a_1962_5182# a_27366_5182# 0.14fF
C5740 a_15926_5142# a_16018_5142# 0.26fF
C5741 a_2346_5184# a_29070_5142# 0.19fF
C5742 a_28066_12170# m2_28264_12418# 0.16fF
C5743 a_7986_14178# ctop 3.58fF
C5744 a_1962_1166# col_n[1] 0.12fF
C5745 a_30074_2130# col_n[27] 0.28fF
C5746 a_26970_9158# rowoff_n[7] 0.24fF
C5747 m2_11772_18014# col_n[9] 0.25fF
C5748 a_1962_14218# col_n[3] 0.13fF
C5749 a_2346_18236# a_7894_18194# 0.35fF
C5750 a_27062_16186# col[24] 0.29fF
C5751 a_30986_15182# rowoff_n[13] 0.24fF
C5752 col[6] rowoff_n[14] 0.11fF
C5753 a_1962_8194# ctop 1.49fF
C5754 a_25966_7150# VDD 0.23fF
C5755 a_12002_14178# rowon_n[12] 0.14fF
C5756 a_2346_16228# a_11910_16186# 0.35fF
C5757 a_2346_7192# col[14] 0.15fF
C5758 a_27062_4138# rowon_n[2] 0.14fF
C5759 a_31078_3134# ctop 3.57fF
C5760 a_34394_18234# vcm 0.22fF
C5761 a_4974_10162# VDD 0.52fF
C5762 a_1962_9198# col_n[30] 0.13fF
C5763 a_12002_9158# a_12002_8154# 1.00fF
C5764 a_28978_9158# a_29070_9158# 0.26fF
C5765 a_12002_2130# vcm 0.62fF
C5766 a_1962_13214# a_5978_13174# 0.27fF
C5767 a_9994_9158# col[7] 0.29fF
C5768 m2_1732_11990# sample 0.19fF
C5769 a_4974_4138# row_n[2] 0.17fF
C5770 m2_34864_5966# ctop 0.17fF
C5771 a_3970_12170# rowoff_n[10] 0.10fF
C5772 a_1962_3174# col[21] 0.11fF
C5773 VDD col_n[6] 4.94fF
C5774 vcm col_n[2] 2.80fF
C5775 a_2346_8196# rowon_n[6] 0.26fF
C5776 a_2346_1168# a_31990_1126# 0.35fF
C5777 ctop col[28] 1.98fF
C5778 a_1962_16226# col[23] 0.11fF
C5779 m3_32988_18146# VDD 0.24fF
C5780 a_25054_13174# m2_25252_13422# 0.16fF
C5781 a_31078_17190# rowon_n[15] 0.14fF
C5782 a_18026_14178# VDD 0.52fF
C5783 a_28066_5142# col[25] 0.29fF
C5784 a_19030_1126# en_bit_n[2] 0.25fF
C5785 a_25054_6146# vcm 0.62fF
C5786 a_1962_15222# a_19030_15182# 0.27fF
C5787 m2_34864_10986# m2_35292_11414# 0.16fF
C5788 a_8290_15222# vcm 0.22fF
C5789 a_18026_16186# rowoff_n[14] 0.10fF
C5790 m2_8760_18014# ctop 0.18fF
C5791 a_23046_3134# a_24050_3134# 0.97fF
C5792 a_3970_1126# m3_4876_1078# 0.14fF
C5793 a_8990_17190# row_n[15] 0.17fF
C5794 a_31078_2130# m3_30980_1078# 0.15fF
C5795 a_25054_13174# a_25054_12170# 1.00fF
C5796 a_1962_12210# a_12306_12210# 0.14fF
C5797 a_2346_12212# a_14010_12170# 0.19fF
C5798 a_24050_7150# row_n[5] 0.17fF
C5799 a_2346_3176# col[5] 0.15fF
C5800 a_1962_17230# a_32082_17190# 0.27fF
C5801 a_2346_16228# col[7] 0.15fF
C5802 m2_7756_946# m3_6884_1078# 0.13fF
C5803 a_9994_11166# col_n[7] 0.28fF
C5804 a_7894_2130# VDD 0.23fF
C5805 a_1962_5182# col_n[21] 0.13fF
C5806 a_31382_4178# vcm 0.22fF
C5807 a_14922_14178# a_15014_14178# 0.26fF
C5808 a_1962_14218# a_25358_14218# 0.14fF
C5809 a_2346_14220# a_27062_14178# 0.19fF
C5810 a_2346_18236# a_2346_17232# 0.22fF
C5811 a_28066_7150# col_n[25] 0.28fF
C5812 a_1962_12210# col[14] 0.11fF
C5813 a_20946_6146# VDD 0.23fF
C5814 a_12002_5142# rowon_n[3] 0.14fF
C5815 a_1962_6186# a_2966_6146# 0.27fF
C5816 a_22042_14178# m2_22240_14426# 0.16fF
C5817 a_16018_17190# ctop 3.39fF
C5818 a_5886_17190# rowoff_n[15] 0.24fF
C5819 a_26058_2130# ctop 3.39fF
C5820 m2_28840_18014# VDD 0.91fF
C5821 a_9902_6146# rowoff_n[4] 0.24fF
C5822 a_33998_10162# VDD 0.23fF
C5823 a_8990_8154# a_9994_8154# 0.97fF
C5824 a_2346_8196# a_16930_8154# 0.35fF
C5825 a_6982_1126# vcm 0.12fF
C5826 a_32994_12170# rowoff_n[10] 0.24fF
C5827 a_19942_4138# rowoff_n[2] 0.24fF
C5828 a_31078_8154# rowon_n[6] 0.14fF
C5829 a_7986_14178# col[5] 0.29fF
C5830 a_1962_5182# a_10998_5142# 0.27fF
C5831 a_1962_1166# col_n[12] 0.13fF
C5832 a_1962_14218# col_n[14] 0.13fF
C5833 a_13006_13174# VDD 0.52fF
C5834 a_2346_10204# a_29982_10162# 0.35fF
C5835 a_29982_2130# rowoff_n[0] 0.24fF
C5836 a_20034_5142# vcm 0.62fF
C5837 m2_24824_946# vcm 0.42fF
C5838 a_26058_10162# col[23] 0.29fF
C5839 a_8990_8154# row_n[6] 0.17fF
C5840 col[17] rowoff_n[14] 0.11fF
C5841 a_1962_8194# col[5] 0.11fF
C5842 a_3270_14218# vcm 0.22fF
C5843 a_21038_3134# a_21038_2130# 1.00fF
C5844 a_1962_2170# a_4274_2170# 0.14fF
C5845 a_2346_2172# a_5978_2130# 0.19fF
C5846 vcm rowoff_n[10] 0.20fF
C5847 m2_21812_18014# m3_20940_18146# 0.13fF
C5848 a_19030_15182# m2_19228_15430# 0.16fF
C5849 a_1962_7190# a_24050_7150# 0.27fF
C5850 a_26058_17190# VDD 0.55fF
C5851 a_2346_7192# col[25] 0.15fF
C5852 a_22042_12170# a_23046_12170# 0.97fF
C5853 a_33086_9158# vcm 0.62fF
C5854 a_21038_3134# m2_21236_3382# 0.16fF
C5855 a_16322_18234# vcm 0.22fF
C5856 a_2346_1168# VDD 36.81fF
C5857 a_1962_4178# a_17326_4178# 0.14fF
C5858 a_2346_4180# a_19030_4138# 0.19fF
C5859 a_10906_4138# a_10998_4138# 0.26fF
C5860 a_7986_16186# col_n[5] 0.28fF
C5861 a_8990_3134# col[6] 0.29fF
C5862 a_26362_3174# vcm 0.22fF
C5863 a_28066_11166# row_n[9] 0.17fF
C5864 vcm col_n[13] 2.80fF
C5865 col_n[6] col_n[7] 0.10fF
C5866 a_18026_10162# rowoff_n[8] 0.10fF
C5867 VDD col_n[17] 4.67fF
C5868 col[1] rowoff_n[15] 0.11fF
C5869 col[16] col[17] 0.20fF
C5870 a_20034_13174# rowoff_n[11] 0.10fF
C5871 m2_5748_946# VDD 0.62fF
C5872 a_15926_5142# VDD 0.23fF
C5873 a_26058_12170# col_n[23] 0.28fF
C5874 a_1962_6186# a_30378_6186# 0.14fF
C5875 a_2346_6188# a_32082_6146# 0.19fF
C5876 a_1962_10202# col_n[5] 0.13fF
C5877 a_34090_7150# a_34090_6146# 1.00fF
C5878 a_10998_16186# ctop 3.57fF
C5879 a_28066_8154# rowoff_n[6] 0.10fF
C5880 a_34090_17190# rowoff_n[15] 0.10fF
C5881 m2_34864_946# col_n[31] 0.30fF
C5882 a_28978_9158# VDD 0.23fF
C5883 a_16018_9158# rowon_n[7] 0.14fF
C5884 a_23958_8154# a_24050_8154# 0.26fF
C5885 a_16018_16186# m2_16216_16434# 0.16fF
C5886 a_6982_8154# a_6982_7150# 1.00fF
C5887 a_2346_3176# col[16] 0.15fF
C5888 a_1962_18234# a_19334_18234# 0.14fF
C5889 a_2346_16228# col[18] 0.15fF
C5890 m2_34864_7974# rowon_n[6] 0.13fF
C5891 a_2346_17232# a_14922_17190# 0.35fF
C5892 a_7986_17190# a_8990_17190# 0.97fF
C5893 m2_21812_18014# m2_22816_18014# 0.96fF
C5894 a_18026_4138# m2_18224_4386# 0.16fF
C5895 a_8990_5142# col_n[6] 0.28fF
C5896 a_34090_5142# ctop 3.42fF
C5897 m3_1864_17142# ctop 0.23fF
C5898 a_7986_12170# VDD 0.52fF
C5899 m2_26832_946# m2_27260_1374# 0.16fF
C5900 a_1962_12210# col[25] 0.11fF
C5901 a_15014_4138# vcm 0.62fF
C5902 a_1962_14218# a_8990_14178# 0.27fF
C5903 a_7894_14178# rowoff_n[12] 0.24fF
C5904 a_18026_2130# a_19030_2130# 0.97fF
C5905 a_2346_2172# a_35002_2130# 0.35fF
C5906 m2_34864_16006# m3_34996_17142# 0.15fF
C5907 a_1962_6186# VDD 2.73fF
C5908 a_24050_15182# col[21] 0.29fF
C5909 a_21038_16186# VDD 0.52fF
C5910 m2_26832_18014# col[24] 0.28fF
C5911 a_2346_11208# a_3970_11166# 0.19fF
C5912 a_20034_12170# a_20034_11166# 1.00fF
C5913 a_28066_8154# vcm 0.62fF
C5914 a_1962_16226# a_22042_16186# 0.27fF
C5915 a_13006_12170# row_n[10] 0.17fF
C5916 a_11302_17230# vcm 0.22fF
C5917 a_28066_2130# row_n[0] 0.17fF
C5918 a_13006_17190# m2_13204_17438# 0.16fF
C5919 a_2346_12212# col[9] 0.15fF
C5920 a_21342_2170# vcm 0.22fF
C5921 a_1962_13214# a_15318_13214# 0.14fF
C5922 a_2346_13216# a_17022_13174# 0.19fF
C5923 a_9902_13174# a_9994_13174# 0.26fF
C5924 a_1962_1166# col_n[23] 0.13fF
C5925 a_6982_8154# col[4] 0.29fF
C5926 a_15014_5142# m2_15212_5390# 0.16fF
C5927 a_1962_14218# col_n[25] 0.13fF
C5928 m2_1732_9982# row_n[8] 0.13fF
C5929 a_10906_4138# VDD 0.23fF
C5930 m3_8892_1078# VDD 0.14fF
C5931 a_31078_6146# a_32082_6146# 0.97fF
C5932 a_5978_15182# ctop 3.58fF
C5933 a_24050_17190# col_n[21] 0.28fF
C5934 col[28] rowoff_n[14] 0.11fF
C5935 a_1962_8194# col[16] 0.11fF
C5936 a_32082_15182# row_n[13] 0.17fF
C5937 a_2346_15224# a_30074_15182# 0.19fF
C5938 a_1962_15222# a_28370_15222# 0.14fF
C5939 a_35398_6186# vcm 0.23fF
C5940 a_33086_16186# a_33086_15182# 1.00fF
C5941 a_25054_4138# col[22] 0.29fF
C5942 m2_34864_11990# VDD 0.99fF
C5943 a_23958_8154# VDD 0.23fF
C5944 a_3970_7150# a_4974_7150# 0.97fF
C5945 a_2346_7192# a_6890_7150# 0.35fF
C5946 m2_16792_946# m3_17928_1078# 0.11fF
C5947 a_22954_17190# a_23046_17190# 0.26fF
C5948 a_5978_17190# a_5978_16186# 1.00fF
C5949 a_10998_5142# rowoff_n[3] 0.10fF
C5950 a_29070_4138# ctop 3.58fF
C5951 a_20034_13174# rowon_n[11] 0.14fF
C5952 a_2874_11166# VDD 0.24fF
C5953 m2_28840_946# m3_27968_1078# 0.13fF
C5954 a_6982_10162# col_n[4] 0.28fF
C5955 a_2346_9200# a_19942_9158# 0.35fF
C5956 VDD col_n[28] 5.01fF
C5957 vcm col_n[24] 2.80fF
C5958 a_2346_8196# col[0] 0.15fF
C5959 col[12] rowoff_n[15] 0.11fF
C5960 a_9994_3134# vcm 0.62fF
C5961 a_21038_3134# rowoff_n[1] 0.10fF
C5962 m2_1732_8978# ctop 0.17fF
C5963 a_1962_10202# col_n[16] 0.13fF
C5964 a_32994_2130# a_33086_2130# 0.26fF
C5965 a_12002_6146# m2_12200_6394# 0.16fF
C5966 m2_34864_12994# m3_34996_14130# 0.15fF
C5967 a_25054_6146# col_n[22] 0.28fF
C5968 a_1962_6186# a_14010_6146# 0.27fF
C5969 a_16018_15182# VDD 0.52fF
C5970 a_2346_11208# a_32994_11166# 0.35fF
C5971 a_17022_11166# a_18026_11166# 0.97fF
C5972 a_1962_4178# col[7] 0.11fF
C5973 a_13006_3134# row_n[1] 0.17fF
C5974 a_7986_17190# m3_7888_18146# 0.15fF
C5975 a_1962_17230# col[9] 0.11fF
C5976 a_23046_7150# vcm 0.62fF
C5977 a_6282_16226# vcm 0.22fF
C5978 a_1962_3174# a_7286_3174# 0.14fF
C5979 a_2346_3176# a_8990_3134# 0.19fF
C5980 a_5886_3134# a_5978_3134# 0.26fF
C5981 a_2346_3176# col[27] 0.15fF
C5982 a_25054_2130# m2_24824_946# 0.99fF
C5983 a_2346_16228# col[29] 0.15fF
C5984 a_1962_8194# a_27062_8154# 0.27fF
C5985 a_16322_1166# vcm 0.23fF
C5986 a_9902_11166# rowoff_n[9] 0.24fF
C5987 a_2346_10204# vcm 0.40fF
C5988 a_17022_16186# row_n[14] 0.17fF
C5989 a_5886_3134# VDD 0.23fF
C5990 a_1962_5182# a_20338_5182# 0.14fF
C5991 a_29070_6146# a_29070_5142# 1.00fF
C5992 a_2346_5184# a_22042_5142# 0.19fF
C5993 a_32082_6146# row_n[4] 0.17fF
C5994 a_4974_13174# col[2] 0.29fF
C5995 a_19942_9158# rowoff_n[7] 0.24fF
C5996 a_29374_5182# vcm 0.22fF
C5997 a_30074_15182# a_31078_15182# 0.97fF
C5998 a_1962_6186# col_n[7] 0.13fF
C5999 a_23958_15182# rowoff_n[13] 0.24fF
C6000 a_2346_7192# m2_34864_6970# 0.17fF
C6001 a_8990_7150# m2_9188_7398# 0.16fF
C6002 m2_1732_17010# m3_1864_17142# 2.76fF
C6003 a_23046_9158# col[20] 0.29fF
C6004 a_18938_7150# VDD 0.23fF
C6005 a_29982_7150# rowoff_n[5] 0.24fF
C6006 a_18938_7150# a_19030_7150# 0.26fF
C6007 a_1962_7190# a_33390_7190# 0.14fF
C6008 a_2966_16186# VDD 0.56fF
C6009 a_4974_14178# rowon_n[12] 0.14fF
C6010 a_1962_13214# col[0] 0.11fF
C6011 a_2346_16228# a_4882_16186# 0.35fF
C6012 a_20034_4138# rowon_n[2] 0.14fF
C6013 a_24050_3134# ctop 3.57fF
C6014 a_2346_12212# col[20] 0.15fF
C6015 a_31990_11166# VDD 0.23fF
C6016 m3_30980_1078# m3_31984_1078# 0.22fF
C6017 m2_21812_946# VDD 0.62fF
C6018 a_4974_2130# vcm 0.62fF
C6019 a_4974_15182# col_n[2] 0.28fF
C6020 a_5978_2130# col[3] 0.29fF
C6021 a_2346_1168# a_24962_1126# 0.35fF
C6022 m2_34864_9982# m3_34996_11118# 0.15fF
C6023 m2_24824_946# col_n[22] 0.37fF
C6024 m3_4876_18146# VDD 0.24fF
C6025 a_24050_17190# rowon_n[15] 0.14fF
C6026 a_1962_8194# col[27] 0.11fF
C6027 a_10998_14178# VDD 0.52fF
C6028 a_15014_11166# a_15014_10162# 1.00fF
C6029 a_31990_11166# a_32082_11166# 0.26fF
C6030 a_23046_11166# col_n[20] 0.28fF
C6031 m2_1732_2954# rowoff_n[1] 0.12fF
C6032 m2_13780_946# col[11] 0.39fF
C6033 a_18026_6146# vcm 0.62fF
C6034 a_1962_15222# a_12002_15182# 0.27fF
C6035 a_1962_2170# sample 0.14fF
C6036 a_10998_16186# rowoff_n[14] 0.10fF
C6037 a_1962_15222# vcm 6.95fF
C6038 a_5978_8154# m2_6176_8402# 0.16fF
C6039 m2_23820_18014# vcm 0.28fF
C6040 a_1962_12210# a_5278_12210# 0.14fF
C6041 a_2346_12212# a_6982_12170# 0.19fF
C6042 a_4882_12170# a_4974_12170# 0.26fF
C6043 a_17022_7150# row_n[5] 0.17fF
C6044 a_31078_10162# vcm 0.62fF
C6045 a_1962_17230# a_25054_17190# 0.27fF
C6046 m2_32856_18014# m2_33284_18442# 0.16fF
C6047 a_34090_3134# VDD 0.54fF
C6048 col_n[2] row_n[15] 0.23fF
C6049 m3_11904_1078# ctop 0.23fF
C6050 VDD row_n[12] 2.93fF
C6051 vcm row_n[14] 0.49fF
C6052 sample row_n[13] 1.03fF
C6053 a_2346_8196# col[11] 0.15fF
C6054 col[27] col[28] 0.20fF
C6055 col[23] rowoff_n[15] 0.11fF
C6056 a_26058_5142# a_27062_5142# 0.97fF
C6057 a_5978_4138# col_n[3] 0.28fF
C6058 a_1962_14218# a_18330_14218# 0.14fF
C6059 a_24354_4178# vcm 0.22fF
C6060 a_28066_15182# a_28066_14178# 1.00fF
C6061 a_2346_14220# a_20034_14178# 0.19fF
C6062 a_1962_10202# col_n[27] 0.13fF
C6063 a_2966_3134# rowoff_n[1] 0.10fF
C6064 m2_1732_13998# m3_1864_14130# 2.76fF
C6065 a_13918_6146# VDD 0.23fF
C6066 a_4974_5142# rowon_n[3] 0.14fF
C6067 a_1962_4178# col[18] 0.11fF
C6068 a_1962_17230# col[20] 0.11fF
C6069 a_8990_17190# ctop 3.39fF
C6070 a_21038_14178# col[18] 0.29fF
C6071 a_17934_16186# a_18026_16186# 0.26fF
C6072 a_1962_16226# a_31382_16226# 0.14fF
C6073 a_2346_16228# a_33086_16186# 0.19fF
C6074 a_19030_2130# ctop 3.50fF
C6075 m2_14784_18014# VDD 1.28fF
C6076 a_2346_6188# rowoff_n[4] 4.09fF
C6077 a_1962_18234# m2_29844_18014# 0.18fF
C6078 a_26970_10162# VDD 0.23fF
C6079 a_2346_8196# a_9902_8154# 0.35fF
C6080 a_12914_4138# rowoff_n[2] 0.24fF
C6081 a_25966_12170# rowoff_n[10] 0.24fF
C6082 a_24050_8154# rowon_n[6] 0.14fF
C6083 a_32082_6146# ctop 3.58fF
C6084 m2_34864_6970# m3_34996_8106# 0.15fF
C6085 a_2346_4180# col[2] 0.15fF
C6086 a_2346_17232# col[4] 0.15fF
C6087 a_1962_5182# a_3970_5142# 0.27fF
C6088 a_3970_7150# col[1] 0.29fF
C6089 a_5978_13174# VDD 0.52fF
C6090 a_2346_18236# m2_24824_18014# 0.19fF
C6091 a_2346_10204# a_22954_10162# 0.35fF
C6092 a_12002_10162# a_13006_10162# 0.97fF
C6093 a_22954_2130# rowoff_n[0] 0.24fF
C6094 a_1962_6186# col_n[18] 0.13fF
C6095 a_13006_5142# vcm 0.62fF
C6096 a_21038_16186# col_n[18] 0.28fF
C6097 a_22042_3134# col[19] 0.29fF
C6098 m2_11772_18014# m3_12908_18146# 0.13fF
C6099 a_1962_7190# a_17022_7150# 0.27fF
C6100 a_1962_13214# col[11] 0.11fF
C6101 a_19030_17190# VDD 0.55fF
C6102 a_26058_9158# vcm 0.62fF
C6103 a_2346_12212# col[31] 0.15fF
C6104 a_9294_18234# vcm 0.22fF
C6105 a_29070_2130# VDD 0.55fF
C6106 a_2346_4180# a_12002_4138# 0.19fF
C6107 a_34090_11166# m2_34288_11414# 0.16fF
C6108 a_24050_5142# a_24050_4138# 1.00fF
C6109 a_1962_4178# a_10298_4178# 0.14fF
C6110 m3_1864_4090# m3_1864_3086# 0.22fF
C6111 a_1962_9198# a_30074_9158# 0.27fF
C6112 a_21038_11166# row_n[9] 0.17fF
C6113 a_19334_3174# vcm 0.22fF
C6114 a_25054_14178# a_26058_14178# 0.97fF
C6115 a_10998_10162# rowoff_n[8] 0.10fF
C6116 a_3970_9158# col_n[1] 0.28fF
C6117 a_13006_13174# rowoff_n[11] 0.10fF
C6118 m2_1732_10986# m3_1864_11118# 2.76fF
C6119 a_8898_5142# VDD 0.23fF
C6120 a_13918_6146# a_14010_6146# 0.26fF
C6121 a_1962_6186# a_23350_6186# 0.14fF
C6122 a_2346_6188# a_25054_6146# 0.19fF
C6123 a_3970_16186# ctop 3.56fF
C6124 a_21038_8154# rowoff_n[6] 0.10fF
C6125 a_22042_5142# col_n[19] 0.28fF
C6126 a_1962_2170# col_n[9] 0.13fF
C6127 a_1962_15222# col_n[11] 0.13fF
C6128 a_32386_7190# vcm 0.22fF
C6129 m2_1732_3958# sample_n 0.15fF
C6130 a_27062_17190# rowoff_n[15] 0.10fF
C6131 m2_1732_15002# VDD 1.02fF
C6132 a_31078_6146# rowoff_n[4] 0.10fF
C6133 a_1962_1166# m2_23820_946# 0.18fF
C6134 a_21950_9158# VDD 0.23fF
C6135 a_8990_9158# rowon_n[7] 0.14fF
C6136 a_1962_9198# col[2] 0.11fF
C6137 a_1962_18234# a_12306_18234# 0.14fF
C6138 m2_1732_11990# rowon_n[10] 0.11fF
C6139 m2_9764_946# m2_10192_1374# 0.16fF
C6140 a_2346_17232# a_7894_17190# 0.35fF
C6141 col_n[13] row_n[15] 0.23fF
C6142 col_n[1] row_n[9] 0.23fF
C6143 col_n[3] row_n[10] 0.23fF
C6144 col_n[0] row_n[8] 0.23fF
C6145 vcm rowon_n[8] 0.50fF
C6146 col_n[7] row_n[12] 0.23fF
C6147 VDD rowon_n[6] 2.61fF
C6148 col_n[5] row_n[11] 0.23fF
C6149 col_n[11] row_n[14] 0.23fF
C6150 col_n[9] row_n[13] 0.23fF
C6151 a_2346_8196# col[22] 0.15fF
C6152 m2_14784_18014# m2_15788_18014# 0.96fF
C6153 a_27062_5142# ctop 3.58fF
C6154 m2_34864_3958# m3_34996_5094# 0.15fF
C6155 m3_7888_18146# ctop 0.23fF
C6156 a_31078_12170# m2_31276_12418# 0.16fF
C6157 a_35002_13174# VDD 0.29fF
C6158 a_9994_10162# a_9994_9158# 1.00fF
C6159 a_26970_10162# a_27062_10162# 0.26fF
C6160 a_7986_4138# vcm 0.62fF
C6161 a_1962_4178# col[29] 0.11fF
C6162 a_28066_12170# rowon_n[10] 0.14fF
C6163 a_2346_2172# a_27974_2130# 0.35fF
C6164 a_1962_17230# col[31] 0.11fF
C6165 a_2346_14220# m2_1732_13998# 0.12fF
C6166 a_14010_16186# VDD 0.52fF
C6167 a_20034_8154# col[17] 0.29fF
C6168 a_1962_11206# col_n[2] 0.13fF
C6169 a_1962_16226# a_15014_16186# 0.27fF
C6170 a_21038_8154# vcm 0.62fF
C6171 a_5978_12170# row_n[10] 0.17fF
C6172 m2_1732_13998# m2_2160_14426# 0.16fF
C6173 a_3970_2130# m2_4168_2378# 0.16fF
C6174 a_4274_17230# vcm 0.22fF
C6175 a_21038_4138# a_22042_4138# 0.97fF
C6176 a_21038_2130# row_n[0] 0.17fF
C6177 a_18026_17190# m2_17796_18014# 1.00fF
C6178 a_2346_13216# a_9994_13174# 0.19fF
C6179 a_1962_13214# a_8290_13214# 0.14fF
C6180 a_23046_14178# a_23046_13174# 1.00fF
C6181 a_14314_2170# vcm 0.22fF
C6182 a_2346_4180# col[13] 0.15fF
C6183 a_34090_12170# vcm 0.62fF
C6184 a_2346_17232# col[15] 0.15fF
C6185 m2_1732_7974# m3_1864_8106# 2.76fF
C6186 m3_1864_11118# VDD 0.25fF
C6187 a_28066_13174# m2_28264_13422# 0.16fF
C6188 a_1962_6186# col_n[29] 0.13fF
C6189 a_2966_10162# a_3970_10162# 0.97fF
C6190 a_25054_15182# row_n[13] 0.17fF
C6191 a_27366_6186# vcm 0.22fF
C6192 a_2346_15224# a_23046_15182# 0.19fF
C6193 a_12914_15182# a_13006_15182# 0.26fF
C6194 a_1962_15222# a_21342_15222# 0.14fF
C6195 a_20034_10162# col_n[17] 0.28fF
C6196 a_1962_13214# col[22] 0.11fF
C6197 a_16930_8154# VDD 0.23fF
C6198 m2_5748_18014# col_n[3] 0.25fF
C6199 a_2346_17232# a_2346_16228# 0.22fF
C6200 a_1962_17230# a_35398_17230# 0.14fF
C6201 m2_34864_18014# m2_34864_17010# 0.99fF
C6202 a_3970_5142# rowoff_n[3] 0.10fF
C6203 a_22042_4138# ctop 3.58fF
C6204 a_13006_13174# rowon_n[11] 0.14fF
C6205 a_29982_12170# VDD 0.23fF
C6206 m3_26964_18146# m3_27968_18146# 0.22fF
C6207 a_6982_9158# a_7986_9158# 0.97fF
C6208 a_2346_9200# a_12914_9158# 0.35fF
C6209 a_2966_11166# row_n[9] 0.16fF
C6210 a_28066_3134# rowon_n[1] 0.14fF
C6211 a_14010_3134# rowoff_n[1] 0.10fF
C6212 a_2346_13216# col[6] 0.15fF
C6213 a_29070_14178# rowoff_n[12] 0.10fF
C6214 a_1962_6186# a_6982_6146# 0.27fF
C6215 a_25054_14178# m2_25252_14426# 0.16fF
C6216 a_1962_2170# col_n[20] 0.13fF
C6217 a_8990_15182# VDD 0.52fF
C6218 a_2966_8154# rowoff_n[6] 0.10fF
C6219 a_1962_15222# col_n[22] 0.13fF
C6220 a_2346_11208# a_25966_11166# 0.35fF
C6221 a_5978_3134# row_n[1] 0.17fF
C6222 a_16018_7150# vcm 0.62fF
C6223 a_18026_13174# col[15] 0.29fF
C6224 a_1962_9198# col[13] 0.11fF
C6225 a_32082_16186# rowon_n[14] 0.14fF
C6226 a_19030_4138# a_19030_3134# 1.00fF
C6227 a_3878_9158# VDD 0.23fF
C6228 a_1962_8194# a_20034_8154# 0.27fF
C6229 a_2966_6146# col[0] 0.29fF
C6230 a_9294_1166# vcm 0.23fF
C6231 col_n[16] row_n[11] 0.23fF
C6232 col_n[22] row_n[14] 0.23fF
C6233 col_n[18] row_n[12] 0.23fF
C6234 col_n[6] row_n[6] 0.23fF
C6235 col_n[12] row_n[9] 0.23fF
C6236 col_n[14] row_n[10] 0.23fF
C6237 col_n[2] row_n[4] 0.23fF
C6238 col_n[10] row_n[8] 0.23fF
C6239 sample row_n[2] 1.03fF
C6240 col_n[4] row_n[5] 0.23fF
C6241 col_n[20] row_n[13] 0.23fF
C6242 col_n[8] row_n[7] 0.23fF
C6243 vcm row_n[3] 0.49fF
C6244 col_n[24] row_n[15] 0.23fF
C6245 VDD row_n[1] 2.93fF
C6246 col_n[28] col_n[29] 0.10fF
C6247 a_20034_13174# a_21038_13174# 0.97fF
C6248 a_2346_11208# rowoff_n[9] 4.09fF
C6249 a_29070_11166# vcm 0.62fF
C6250 a_9994_16186# row_n[14] 0.17fF
C6251 m2_1732_4962# m3_1864_5094# 2.76fF
C6252 a_32082_4138# VDD 0.52fF
C6253 a_1962_5182# a_13310_5182# 0.14fF
C6254 a_8898_5142# a_8990_5142# 0.26fF
C6255 a_2346_5184# a_15014_5142# 0.19fF
C6256 a_25054_6146# row_n[4] 0.17fF
C6257 a_1962_10202# a_33086_10162# 0.27fF
C6258 a_12914_9158# rowoff_n[7] 0.24fF
C6259 a_22346_5182# vcm 0.22fF
C6260 a_16930_15182# rowoff_n[13] 0.24fF
C6261 m2_26832_18014# m3_25960_18146# 0.13fF
C6262 a_1962_18234# VDD 29.26fF
C6263 a_11910_7150# VDD 0.23fF
C6264 a_18026_15182# col_n[15] 0.28fF
C6265 a_22954_7150# rowoff_n[5] 0.24fF
C6266 a_32082_8154# a_32082_7150# 1.00fF
C6267 a_2346_7192# a_28066_7150# 0.19fF
C6268 a_1962_7190# a_26362_7190# 0.14fF
C6269 a_22042_15182# m2_22240_15430# 0.16fF
C6270 a_1962_11206# col_n[13] 0.13fF
C6271 a_19030_2130# col[16] 0.29fF
C6272 a_2966_8154# vcm 0.61fF
C6273 a_33086_17190# a_34090_17190# 0.97fF
C6274 a_24050_3134# m2_24248_3382# 0.16fF
C6275 a_1962_5182# col[4] 0.11fF
C6276 a_32994_5142# rowoff_n[3] 0.24fF
C6277 a_13006_4138# rowon_n[2] 0.14fF
C6278 a_17022_3134# ctop 3.57fF
C6279 a_24962_11166# VDD 0.23fF
C6280 m3_16924_1078# m3_17928_1078# 0.22fF
C6281 a_4974_9158# a_4974_8154# 1.00fF
C6282 a_21950_9158# a_22042_9158# 0.26fF
C6283 a_2346_4180# col[24] 0.15fF
C6284 a_2346_17232# col[26] 0.15fF
C6285 a_2346_1168# a_17934_1126# 0.39fF
C6286 a_30074_7150# ctop 3.58fF
C6287 a_1962_6186# a_34394_6186# 0.14fF
C6288 a_17022_17190# rowon_n[15] 0.14fF
C6289 a_3970_14178# VDD 0.52fF
C6290 m2_1732_4962# vcm 0.45fF
C6291 VDD rowoff_n[13] 1.17fF
C6292 a_10998_6146# vcm 0.62fF
C6293 a_3878_15182# a_3970_15182# 0.26fF
C6294 a_1962_15222# a_4974_15182# 0.27fF
C6295 a_32082_7150# rowon_n[5] 0.14fF
C6296 a_19030_4138# col_n[16] 0.28fF
C6297 rowon_n[0] rowoff_n[0] 20.27fF
C6298 a_3970_16186# rowoff_n[14] 0.10fF
C6299 ctop rowoff_n[4] 0.60fF
C6300 a_2346_3176# a_30986_3134# 0.35fF
C6301 a_16018_3134# a_17022_3134# 0.97fF
C6302 a_1962_7190# col_n[4] 0.13fF
C6303 a_19030_16186# m2_19228_16434# 0.16fF
C6304 m2_9764_18014# vcm 0.28fF
C6305 a_18026_13174# a_18026_12170# 1.00fF
C6306 a_9994_7150# row_n[5] 0.17fF
C6307 a_24050_10162# vcm 0.62fF
C6308 a_31078_11166# rowoff_n[9] 0.10fF
C6309 a_1962_17230# a_18026_17190# 0.27fF
C6310 m2_25828_18014# m2_26256_18442# 0.16fF
C6311 a_21038_4138# m2_21236_4386# 0.16fF
C6312 a_34090_14178# col[31] 0.29fF
C6313 m2_34864_2954# m3_34996_2082# 0.15fF
C6314 m2_1732_1950# m3_1864_2082# 2.76fF
C6315 a_27062_3134# VDD 0.52fF
C6316 m3_34996_10114# ctop 0.23fF
C6317 a_2346_13216# col[17] 0.15fF
C6318 a_17326_4178# vcm 0.22fF
C6319 a_2346_14220# a_13006_14178# 0.19fF
C6320 a_7894_14178# a_7986_14178# 0.26fF
C6321 a_1962_14218# a_11302_14218# 0.14fF
C6322 a_1962_2170# col_n[31] 0.13fF
C6323 a_6890_6146# VDD 0.23fF
C6324 a_29070_7150# a_30074_7150# 0.97fF
C6325 a_29070_10162# row_n[8] 0.17fF
C6326 a_1962_9198# col[24] 0.11fF
C6327 a_31078_17190# a_31078_16186# 1.00fF
C6328 a_30378_8194# vcm 0.22fF
C6329 a_1962_16226# a_24354_16226# 0.14fF
C6330 a_2346_16228# a_26058_16186# 0.19fF
C6331 a_17022_7150# col[14] 0.29fF
C6332 a_12002_2130# ctop 3.39fF
C6333 a_1962_18234# m2_15788_18014# 0.18fF
C6334 a_19942_10162# VDD 0.23fF
C6335 col_n[15] row_n[5] 0.23fF
C6336 VDD col[0] 10.03fF
C6337 col_n[23] row_n[9] 0.23fF
C6338 col_n[13] row_n[4] 0.23fF
C6339 col_n[27] row_n[11] 0.23fF
C6340 col_n[11] row_n[3] 0.23fF
C6341 col_n[25] row_n[10] 0.23fF
C6342 col_n[19] row_n[7] 0.23fF
C6343 col_n[9] row_n[2] 0.23fF
C6344 col_n[5] row_n[0] 0.23fF
C6345 col_n[2] ctop 2.02fF
C6346 col_n[1] en_C0_n 0.17fF
C6347 col_n[29] row_n[12] 0.23fF
C6348 col_n[21] row_n[8] 0.23fF
C6349 col_n[17] row_n[6] 0.23fF
C6350 col_n[7] row_n[1] 0.23fF
C6351 col_n[31] row_n[13] 0.23fF
C6352 a_16018_17190# m2_16216_17438# 0.16fF
C6353 a_34090_16186# col_n[31] 0.28fF
C6354 a_18938_12170# rowoff_n[10] 0.24fF
C6355 a_5886_4138# rowoff_n[2] 0.24fF
C6356 a_17022_8154# rowon_n[6] 0.14fF
C6357 a_18026_5142# m2_18224_5390# 0.16fF
C6358 a_25054_6146# ctop 3.58fF
C6359 m3_23952_1078# VDD 0.14fF
C6360 a_32994_14178# VDD 0.23fF
C6361 a_2346_18236# m2_10768_18014# 0.19fF
C6362 a_2346_10204# a_15926_10162# 0.35fF
C6363 a_2346_9200# col[8] 0.15fF
C6364 a_15926_2130# rowoff_n[0] 0.24fF
C6365 a_5978_5142# vcm 0.62fF
C6366 a_1962_18234# col_n[7] 0.13fF
C6367 a_32994_16186# rowoff_n[14] 0.24fF
C6368 a_14010_3134# a_14010_2130# 1.00fF
C6369 a_1962_11206# col_n[24] 0.13fF
C6370 a_30986_3134# a_31078_3134# 0.26fF
C6371 a_17022_9158# col_n[14] 0.28fF
C6372 m2_2736_18014# m3_2868_18146# 2.78fF
C6373 a_1962_7190# a_9994_7150# 0.27fF
C6374 a_12002_17190# VDD 0.55fF
C6375 a_2346_12212# a_28978_12170# 0.35fF
C6376 a_15014_12170# a_16018_12170# 0.97fF
C6377 a_1962_5182# col[15] 0.11fF
C6378 a_19030_9158# vcm 0.62fF
C6379 a_22042_2130# VDD 0.55fF
C6380 m2_20808_18014# col[18] 0.28fF
C6381 a_1962_4178# a_3270_4178# 0.14fF
C6382 a_2346_4180# a_4974_4138# 0.19fF
C6383 m3_1864_11118# m3_1864_10114# 0.22fF
C6384 a_1962_9198# a_23046_9158# 0.27fF
C6385 a_16930_18194# m2_16792_18014# 0.16fF
C6386 a_14010_11166# row_n[9] 0.17fF
C6387 a_12306_3174# vcm 0.22fF
C6388 a_3970_10162# rowoff_n[8] 0.10fF
C6389 a_5978_13174# rowoff_n[11] 0.10fF
C6390 a_32082_13174# vcm 0.62fF
C6391 a_15014_6146# m2_15212_6394# 0.16fF
C6392 a_2346_6188# a_18026_6146# 0.19fF
C6393 a_1962_6186# a_16322_6186# 0.14fF
C6394 a_27062_7150# a_27062_6146# 1.00fF
C6395 a_14010_8154# rowoff_n[6] 0.10fF
C6396 a_10998_17190# m3_10900_18146# 0.15fF
C6397 col[7] rowoff_n[6] 0.11fF
C6398 col[10] rowoff_n[9] 0.11fF
C6399 col[9] rowoff_n[8] 0.11fF
C6400 col[8] rowoff_n[7] 0.11fF
C6401 col[4] rowoff_n[3] 0.11fF
C6402 col[2] rowoff_n[1] 0.11fF
C6403 col[3] rowoff_n[2] 0.11fF
C6404 col[1] rowoff_n[0] 0.11fF
C6405 col[5] rowoff_n[4] 0.11fF
C6406 col[6] rowoff_n[5] 0.11fF
C6407 a_25358_7190# vcm 0.22fF
C6408 a_28066_16186# a_29070_16186# 0.97fF
C6409 a_20034_17190# rowoff_n[15] 0.10fF
C6410 a_1962_7190# col_n[15] 0.13fF
C6411 a_24050_6146# rowoff_n[4] 0.10fF
C6412 a_15014_12170# col[12] 0.29fF
C6413 m2_10768_946# col[8] 0.39fF
C6414 a_14922_9158# VDD 0.23fF
C6415 a_2346_8196# a_31078_8154# 0.19fF
C6416 a_16930_8154# a_17022_8154# 0.26fF
C6417 a_1962_8194# a_29374_8194# 0.14fF
C6418 a_33086_14178# row_n[12] 0.17fF
C6419 a_1962_1166# col[6] 0.11fF
C6420 a_1962_18234# a_5278_18234# 0.14fF
C6421 a_1962_14218# col[8] 0.11fF
C6422 a_34090_4138# rowoff_n[2] 0.10fF
C6423 a_33086_8154# col[30] 0.29fF
C6424 m2_7756_18014# m2_8760_18014# 0.96fF
C6425 a_20034_5142# ctop 3.58fF
C6426 m2_24824_946# ctop 0.18fF
C6427 a_27974_13174# VDD 0.23fF
C6428 a_2346_13216# col[28] 0.15fF
C6429 ctop rowoff_n[10] 0.60fF
C6430 a_21038_12170# rowon_n[10] 0.14fF
C6431 a_12002_7150# m2_12200_7398# 0.16fF
C6432 a_2346_2172# a_20946_2130# 0.35fF
C6433 a_10998_2130# a_12002_2130# 0.97fF
C6434 a_33086_9158# ctop 3.57fF
C6435 a_2966_9158# m3_1864_9110# 0.14fF
C6436 a_6982_16186# VDD 0.52fF
C6437 a_15014_14178# col_n[12] 0.28fF
C6438 a_29982_12170# a_30074_12170# 0.26fF
C6439 a_13006_12170# a_13006_11166# 1.00fF
C6440 a_14010_8154# vcm 0.62fF
C6441 a_1962_16226# a_7986_16186# 0.27fF
C6442 a_1962_3174# col_n[6] 0.13fF
C6443 col_n[3] col[4] 5.98fF
C6444 col_n[13] ctop 2.02fF
C6445 col_n[18] row_n[1] 0.23fF
C6446 col_n[22] row_n[3] 0.23fF
C6447 col_n[30] row_n[7] 0.23fF
C6448 a_1962_16226# col_n[8] 0.13fF
C6449 col_n[28] row_n[6] 0.23fF
C6450 col_n[20] row_n[2] 0.23fF
C6451 col_n[24] row_n[4] 0.23fF
C6452 col_n[26] row_n[5] 0.23fF
C6453 vcm col[7] 5.84fF
C6454 VDD col[11] 4.17fF
C6455 col_n[16] row_n[0] 0.22fF
C6456 a_2346_4180# a_33998_4138# 0.35fF
C6457 a_35494_11528# VDD 0.11fF
C6458 a_14010_2130# row_n[0] 0.17fF
C6459 a_33086_10162# col_n[30] 0.28fF
C6460 a_7286_2170# vcm 0.22fF
C6461 a_2346_13216# a_2874_13174# 0.35fF
C6462 a_32994_10162# rowoff_n[8] 0.24fF
C6463 m2_1732_3958# m2_1732_2954# 0.99fF
C6464 a_27062_12170# vcm 0.62fF
C6465 a_35002_13174# rowoff_n[11] 0.24fF
C6466 a_30074_5142# VDD 0.52fF
C6467 m3_19936_18146# VDD 0.29fF
C6468 a_24050_6146# a_25054_6146# 0.97fF
C6469 a_2346_9200# col[19] 0.15fF
C6470 a_18026_15182# row_n[13] 0.17fF
C6471 a_1962_18234# col_n[18] 0.13fF
C6472 a_26058_16186# a_26058_15182# 1.00fF
C6473 a_20338_6186# vcm 0.22fF
C6474 a_2346_15224# a_16018_15182# 0.19fF
C6475 a_1962_15222# a_14314_15222# 0.14fF
C6476 a_33086_5142# row_n[3] 0.17fF
C6477 a_2346_8196# m2_34864_7974# 0.17fF
C6478 a_8990_8154# m2_9188_8402# 0.16fF
C6479 a_16018_3134# col_n[13] 0.28fF
C6480 a_9902_8154# VDD 0.23fF
C6481 a_1962_5182# col[26] 0.11fF
C6482 a_13006_17190# col[10] 0.29fF
C6483 a_33390_10202# vcm 0.22fF
C6484 a_2346_17232# a_29070_17190# 0.19fF
C6485 a_15926_17190# a_16018_17190# 0.26fF
C6486 a_1962_17230# a_27366_17230# 0.14fF
C6487 a_1962_12210# col_n[0] 0.13fF
C6488 m2_2736_946# m3_2868_1078# 2.79fF
C6489 a_15014_4138# ctop 3.58fF
C6490 m3_26964_1078# ctop 0.23fF
C6491 a_5978_13174# rowon_n[11] 0.14fF
C6492 a_31078_13174# col[28] 0.29fF
C6493 a_22954_12170# VDD 0.23fF
C6494 m3_12908_18146# m3_13912_18146# 0.22fF
C6495 a_2346_9200# a_5886_9158# 0.35fF
C6496 a_6982_3134# rowoff_n[1] 0.10fF
C6497 a_21038_3134# rowon_n[1] 0.14fF
C6498 a_22042_14178# rowoff_n[12] 0.10fF
C6499 a_25966_2130# a_26058_2130# 0.26fF
C6500 a_28066_8154# ctop 3.58fF
C6501 a_2346_5184# col[10] 0.15fF
C6502 col[20] rowoff_n[8] 0.11fF
C6503 col[19] rowoff_n[7] 0.11fF
C6504 col[12] rowoff_n[0] 0.11fF
C6505 col[21] rowoff_n[9] 0.11fF
C6506 col[17] rowoff_n[5] 0.11fF
C6507 col[18] rowoff_n[6] 0.11fF
C6508 col[13] rowoff_n[1] 0.11fF
C6509 col[14] rowoff_n[2] 0.11fF
C6510 col[15] rowoff_n[3] 0.11fF
C6511 col[16] rowoff_n[4] 0.11fF
C6512 a_9994_11166# a_10998_11166# 0.97fF
C6513 a_2346_11208# a_18938_11166# 0.35fF
C6514 m2_22816_946# col[20] 0.39fF
C6515 a_1962_7190# col_n[26] 0.13fF
C6516 a_8990_7150# vcm 0.62fF
C6517 a_25054_16186# rowon_n[14] 0.14fF
C6518 a_14010_6146# col[11] 0.29fF
C6519 a_5978_9158# m2_6176_9406# 0.16fF
C6520 a_1962_1166# col[17] 0.11fF
C6521 a_1962_8194# a_13006_8154# 0.27fF
C6522 a_1962_14218# col[19] 0.11fF
C6523 a_2346_13216# a_31990_13174# 0.35fF
C6524 a_31078_15182# col_n[28] 0.28fF
C6525 a_22042_11166# vcm 0.62fF
C6526 a_32082_2130# col[29] 0.29fF
C6527 a_25054_4138# VDD 0.52fF
C6528 a_1962_5182# a_6282_5182# 0.14fF
C6529 a_22042_6146# a_22042_5142# 1.00fF
C6530 a_2346_5184# a_7986_5142# 0.19fF
C6531 col[5] rowoff_n[10] 0.11fF
C6532 a_18026_6146# row_n[4] 0.17fF
C6533 a_1962_10202# a_26058_10162# 0.27fF
C6534 a_5886_9158# rowoff_n[7] 0.24fF
C6535 a_15318_5182# vcm 0.22fF
C6536 a_23046_15182# a_24050_15182# 0.97fF
C6537 a_9902_15182# rowoff_n[13] 0.24fF
C6538 a_35094_15182# vcm 0.12fF
C6539 a_2966_12170# rowon_n[10] 0.13fF
C6540 a_2346_2172# a_1962_2170# 2.62fF
C6541 m2_16792_18014# m3_17928_18146# 0.13fF
C6542 a_2346_1168# col[1] 0.14fF
C6543 a_4882_7150# VDD 0.23fF
C6544 a_2346_14220# col[3] 0.15fF
C6545 a_15926_7150# rowoff_n[5] 0.24fF
C6546 a_1962_7190# a_19334_7190# 0.14fF
C6547 a_11910_7150# a_12002_7150# 0.26fF
C6548 a_2346_7192# a_21038_7150# 0.19fF
C6549 a_14010_8154# col_n[11] 0.28fF
C6550 a_1962_3174# col_n[17] 0.13fF
C6551 col_n[31] row_n[2] 0.23fF
C6552 vcm col[18] 5.84fF
C6553 VDD col[22] 4.17fF
C6554 col_n[9] col[9] 0.72fF
C6555 col_n[24] ctop 2.02fF
C6556 col_n[29] row_n[1] 0.23fF
C6557 rowon_n[9] rowon_n[8] 0.15fF
C6558 col_n[27] row_n[0] 0.23fF
C6559 a_1962_16226# col_n[19] 0.13fF
C6560 a_28370_9198# vcm 0.22fF
C6561 a_5978_4138# rowon_n[2] 0.14fF
C6562 a_25966_5142# rowoff_n[3] 0.24fF
C6563 a_9994_3134# ctop 3.57fF
C6564 a_32082_4138# col_n[29] 0.28fF
C6565 a_17934_11166# VDD 0.23fF
C6566 a_1962_10202# col[10] 0.11fF
C6567 m3_2868_1078# m3_3872_1078# 0.14fF
C6568 a_2346_9200# a_34090_9158# 0.19fF
C6569 a_1962_9198# a_32386_9198# 0.14fF
C6570 a_2346_1168# a_10906_1126# 0.35fF
C6571 a_2346_9200# col[30] 0.15fF
C6572 a_23046_7150# ctop 3.58fF
C6573 a_9994_17190# rowon_n[15] 0.14fF
C6574 a_30986_15182# VDD 0.23fF
C6575 a_1962_18234# col_n[29] 0.13fF
C6576 a_7986_11166# a_7986_10162# 1.00fF
C6577 a_24962_11166# a_25054_11166# 0.26fF
C6578 m2_1732_2954# rowon_n[1] 0.11fF
C6579 m2_14784_946# a_2346_1168# 0.19fF
C6580 a_25054_7150# rowon_n[5] 0.14fF
C6581 a_3970_6146# vcm 0.62fF
C6582 a_2346_3176# a_23958_3134# 0.35fF
C6583 a_2346_1168# m2_31852_946# 0.19fF
C6584 a_2346_10204# ctop 1.59fF
C6585 a_12002_11166# col[9] 0.29fF
C6586 a_1962_12210# col_n[10] 0.13fF
C6587 a_17022_10162# vcm 0.62fF
C6588 a_24050_11166# rowoff_n[9] 0.10fF
C6589 a_1962_17230# a_10998_17190# 0.27fF
C6590 m2_18800_18014# m2_19228_18442# 0.16fF
C6591 a_20034_3134# VDD 0.52fF
C6592 m3_22948_18146# ctop 0.23fF
C6593 a_34090_12170# m2_34288_12418# 0.16fF
C6594 a_1962_5182# a_1962_4178# 0.16fF
C6595 a_19030_5142# a_20034_5142# 0.97fF
C6596 a_1962_6186# col[1] 0.11fF
C6597 a_30074_7150# col[27] 0.29fF
C6598 a_34090_9158# rowoff_n[7] 0.10fF
C6599 a_10298_4178# vcm 0.22fF
C6600 a_21038_15182# a_21038_14178# 1.00fF
C6601 a_1962_14218# a_4274_14218# 0.14fF
C6602 a_2346_14220# a_5978_14178# 0.19fF
C6603 a_2966_3134# rowon_n[1] 0.13fF
C6604 a_30074_14178# vcm 0.62fF
C6605 a_2346_5184# col[21] 0.15fF
C6606 a_1962_2170# a_31078_2130# 0.27fF
C6607 col[28] rowoff_n[5] 0.11fF
C6608 col[27] rowoff_n[4] 0.11fF
C6609 col[29] rowoff_n[6] 0.11fF
C6610 col[30] rowoff_n[7] 0.11fF
C6611 col[26] rowoff_n[3] 0.11fF
C6612 col[31] rowoff_n[8] 0.11fF
C6613 col[24] rowoff_n[1] 0.11fF
C6614 col[25] rowoff_n[2] 0.11fF
C6615 col[23] rowoff_n[0] 0.11fF
C6616 a_33086_7150# VDD 0.52fF
C6617 a_22042_10162# row_n[8] 0.17fF
C6618 a_23350_8194# vcm 0.22fF
C6619 a_10906_16186# a_10998_16186# 0.26fF
C6620 a_2346_16228# a_19030_16186# 0.19fF
C6621 a_1962_16226# a_17326_16226# 0.14fF
C6622 a_12002_13174# col_n[9] 0.28fF
C6623 a_6982_2130# m2_7180_2378# 0.16fF
C6624 a_4974_2130# ctop 3.38fF
C6625 a_1962_1166# col[28] 0.11fF
C6626 a_1962_18234# m2_1732_18014# 0.15fF
C6627 a_1962_14218# col[30] 0.11fF
C6628 a_12914_10162# VDD 0.23fF
C6629 a_32082_9158# a_33086_9158# 0.97fF
C6630 a_1962_8194# col_n[1] 0.13fF
C6631 a_30074_9158# col_n[27] 0.28fF
C6632 a_11910_12170# rowoff_n[10] 0.24fF
C6633 a_9994_8154# rowon_n[6] 0.14fF
C6634 col[16] rowoff_n[10] 0.11fF
C6635 a_18026_6146# ctop 3.58fF
C6636 a_31078_13174# m2_31276_13422# 0.16fF
C6637 m3_34996_4090# VDD 0.26fF
C6638 a_1962_15222# ctop 1.49fF
C6639 a_25966_14178# VDD 0.23fF
C6640 a_2346_10204# a_8898_10162# 0.35fF
C6641 a_4974_10162# a_5978_10162# 0.97fF
C6642 a_8898_2130# rowoff_n[0] 0.24fF
C6643 a_2346_1168# col[12] 0.14fF
C6644 m2_23820_18014# ctop 0.18fF
C6645 a_25966_16186# rowoff_n[14] 0.24fF
C6646 a_2346_14220# col[14] 0.15fF
C6647 a_31078_10162# ctop 3.58fF
C6648 a_2346_15224# m2_1732_15002# 0.12fF
C6649 a_2346_7192# a_2966_7150# 0.21fF
C6650 a_1962_3174# col_n[28] 0.13fF
C6651 a_13006_2130# col_n[10] 0.28fF
C6652 a_4974_17190# VDD 0.55fF
C6653 rowon_n[6] row_n[6] 19.75fF
C6654 col_n[14] col[15] 5.99fF
C6655 sample_n rowoff_n[15] 0.38fF
C6656 vcm col[29] 5.84fF
C6657 row_n[14] ctop 1.65fF
C6658 a_1962_16226# col_n[30] 0.13fF
C6659 a_2346_12212# a_21950_12170# 0.35fF
C6660 m2_34864_17010# vcm 0.50fF
C6661 m2_12776_946# m3_12908_1078# 2.79fF
C6662 a_29070_11166# rowon_n[9] 0.14fF
C6663 a_12002_9158# vcm 0.62fF
C6664 col[0] rowoff_n[11] 0.11fF
C6665 a_9994_16186# col[7] 0.29fF
C6666 a_15014_2130# VDD 0.55fF
C6667 a_1962_10202# col[21] 0.11fF
C6668 a_33998_5142# a_34090_5142# 0.26fF
C6669 a_17022_5142# a_17022_4138# 1.00fF
C6670 m2_23820_946# m3_24956_1078# 0.13fF
C6671 a_1962_9198# a_16018_9158# 0.27fF
C6672 a_6982_11166# row_n[9] 0.17fF
C6673 a_28066_12170# col[25] 0.29fF
C6674 a_5278_3174# vcm 0.22fF
C6675 a_2346_14220# a_35002_14178# 0.35fF
C6676 a_18026_14178# a_19030_14178# 0.97fF
C6677 a_25054_13174# vcm 0.62fF
C6678 a_28066_6146# VDD 0.52fF
C6679 a_28066_14178# m2_28264_14426# 0.16fF
C6680 a_2346_6188# a_10998_6146# 0.19fF
C6681 a_6890_6146# a_6982_6146# 0.26fF
C6682 a_1962_6186# a_9294_6186# 0.14fF
C6683 a_6982_8154# rowoff_n[6] 0.10fF
C6684 a_1962_11206# a_29070_11166# 0.27fF
C6685 a_18330_7190# vcm 0.22fF
C6686 a_2346_10204# col[5] 0.15fF
C6687 a_13006_17190# rowoff_n[15] 0.10fF
C6688 a_33998_2130# ctop 0.10fF
C6689 a_17022_6146# rowoff_n[4] 0.10fF
C6690 a_34090_3134# m3_34996_3086# 0.13fF
C6691 a_7894_9158# VDD 0.23fF
C6692 a_2346_8196# a_24050_8154# 0.19fF
C6693 a_1962_8194# a_22346_8194# 0.14fF
C6694 a_30074_9158# a_30074_8154# 1.00fF
C6695 a_26058_14178# row_n[12] 0.17fF
C6696 a_10998_5142# col[8] 0.29fF
C6697 a_1962_12210# col_n[21] 0.13fF
C6698 m2_1732_7974# sample 0.19fF
C6699 a_27062_4138# rowoff_n[2] 0.10fF
C6700 a_31382_11206# vcm 0.22fF
C6701 m2_33860_946# col[31] 0.26fF
C6702 a_1962_6186# col[12] 0.11fF
C6703 a_28066_14178# col_n[25] 0.28fF
C6704 a_13006_5142# ctop 3.58fF
C6705 a_20946_13174# VDD 0.23fF
C6706 a_19942_10162# a_20034_10162# 0.26fF
C6707 m2_34864_8978# m2_35292_9406# 0.16fF
C6708 a_14010_12170# rowon_n[10] 0.14fF
C6709 a_2346_2172# a_13918_2130# 0.35fF
C6710 a_26058_9158# ctop 3.58fF
C6711 m2_31852_18014# m3_30980_18146# 0.13fF
C6712 a_25054_15182# m2_25252_15430# 0.16fF
C6713 a_29070_2130# rowon_n[0] 0.14fF
C6714 a_33998_17190# VDD 0.24fF
C6715 a_6982_8154# vcm 0.62fF
C6716 a_10998_7150# col_n[8] 0.28fF
C6717 a_27062_3134# m2_27260_3382# 0.16fF
C6718 a_14010_4138# a_15014_4138# 0.97fF
C6719 a_2346_4180# a_26970_4138# 0.35fF
C6720 a_6982_2130# row_n[0] 0.17fF
C6721 a_1962_8194# col_n[12] 0.13fF
C6722 m2_13780_946# VDD 0.62fF
C6723 a_16018_14178# a_16018_13174# 1.00fF
C6724 a_29070_3134# col_n[26] 0.28fF
C6725 a_32994_14178# a_33086_14178# 0.26fF
C6726 a_25966_10162# rowoff_n[8] 0.24fF
C6727 col[27] rowoff_n[10] 0.11fF
C6728 a_33086_15182# rowon_n[13] 0.14fF
C6729 a_2966_5142# col_n[0] 0.28fF
C6730 a_20034_12170# vcm 0.62fF
C6731 a_27974_13174# rowoff_n[11] 0.24fF
C6732 a_1962_2170# col[3] 0.11fF
C6733 a_26058_17190# col[23] 0.29fF
C6734 a_1962_15222# col[5] 0.11fF
C6735 a_23046_5142# VDD 0.52fF
C6736 m2_30848_946# VDD 0.62fF
C6737 a_2346_1168# col[23] 0.14fF
C6738 a_10998_15182# row_n[13] 0.17fF
C6739 a_13310_6186# vcm 0.22fF
C6740 a_2346_14220# col[25] 0.15fF
C6741 a_1962_15222# a_7286_15222# 0.14fF
C6742 a_5886_15182# a_5978_15182# 0.26fF
C6743 a_2346_15224# a_8990_15182# 0.19fF
C6744 a_33086_16186# vcm 0.62fF
C6745 a_26058_5142# row_n[3] 0.17fF
C6746 a_1962_3174# a_34090_3134# 0.27fF
C6747 a_2346_8196# VDD 32.63fF
C6748 rowon_n[8] ctop 1.40fF
C6749 col_n[20] col[20] 0.72fF
C6750 a_22042_16186# m2_22240_16434# 0.16fF
C6751 a_27062_8154# a_28066_8154# 0.97fF
C6752 col[11] rowoff_n[11] 0.11fF
C6753 a_2874_12170# a_2966_12170# 0.26fF
C6754 a_2346_12212# a_3878_12170# 0.35fF
C6755 a_26362_10202# vcm 0.22fF
C6756 a_8990_10162# col[6] 0.29fF
C6757 a_1962_17230# a_20338_17230# 0.14fF
C6758 a_2346_17232# a_22042_17190# 0.19fF
C6759 a_24050_4138# m2_24248_4386# 0.16fF
C6760 a_7986_4138# ctop 3.58fF
C6761 a_1962_4178# col_n[3] 0.13fF
C6762 a_15926_12170# VDD 0.23fF
C6763 m2_34864_946# m2_35292_1374# 0.16fF
C6764 a_1962_17230# col_n[5] 0.13fF
C6765 a_27062_6146# col[24] 0.29fF
C6766 a_14010_3134# rowon_n[1] 0.14fF
C6767 a_15014_14178# rowoff_n[12] 0.10fF
C6768 a_21038_8154# ctop 3.58fF
C6769 a_28978_16186# VDD 0.23fF
C6770 a_2346_11208# a_11910_11166# 0.35fF
C6771 a_2346_10204# col[16] 0.15fF
C6772 a_34394_8194# vcm 0.22fF
C6773 a_18026_16186# rowon_n[14] 0.14fF
C6774 a_28978_4138# a_29070_4138# 0.26fF
C6775 a_12002_4138# a_12002_3134# 1.00fF
C6776 a_8990_12170# col_n[6] 0.28fF
C6777 a_34090_12170# ctop 3.42fF
C6778 a_1962_8194# a_5978_8154# 0.27fF
C6779 a_19030_17190# m2_19228_17438# 0.16fF
C6780 a_33086_6146# rowon_n[4] 0.14fF
C6781 a_13006_13174# a_14010_13174# 0.97fF
C6782 a_2346_13216# a_24962_13174# 0.35fF
C6783 a_1962_6186# col[23] 0.11fF
C6784 a_15014_11166# vcm 0.62fF
C6785 a_27062_8154# col_n[24] 0.28fF
C6786 a_21038_5142# m2_21236_5390# 0.16fF
C6787 a_18026_4138# VDD 0.52fF
C6788 a_10998_6146# row_n[4] 0.17fF
C6789 a_1962_13214# VDD 2.73fF
C6790 a_1962_10202# a_19030_10162# 0.27fF
C6791 a_2966_15182# a_2966_14178# 1.00fF
C6792 a_8290_5182# vcm 0.22fF
C6793 a_2346_15224# rowoff_n[13] 4.09fF
C6794 a_28066_15182# vcm 0.62fF
C6795 m2_7756_18014# m3_7888_18146# 2.79fF
C6796 a_31078_8154# VDD 0.52fF
C6797 a_8898_7150# rowoff_n[5] 0.24fF
C6798 a_25054_8154# a_25054_7150# 1.00fF
C6799 a_1962_7190# a_12306_7190# 0.14fF
C6800 a_2346_7192# a_14010_7150# 0.19fF
C6801 a_1962_12210# a_32082_12170# 0.27fF
C6802 a_2346_6188# col[7] 0.15fF
C6803 a_21342_9198# vcm 0.22fF
C6804 a_26058_17190# a_27062_17190# 0.97fF
C6805 a_18938_5142# rowoff_n[3] 0.24fF
C6806 a_1962_8194# col_n[23] 0.13fF
C6807 a_30074_9158# row_n[7] 0.17fF
C6808 a_6982_15182# col[4] 0.29fF
C6809 a_10906_11166# VDD 0.23fF
C6810 a_1962_9198# a_25358_9198# 0.14fF
C6811 a_2346_9200# a_27062_9158# 0.19fF
C6812 a_14922_9158# a_15014_9158# 0.26fF
C6813 a_1962_2170# col[14] 0.11fF
C6814 a_28978_3134# rowoff_n[1] 0.24fF
C6815 a_1962_15222# col[16] 0.11fF
C6816 a_35398_13214# vcm 0.23fF
C6817 a_25054_11166# col[22] 0.29fF
C6818 a_18026_6146# m2_18224_6394# 0.16fF
C6819 a_16018_7150# ctop 3.58fF
C6820 a_23958_15182# VDD 0.23fF
C6821 a_14010_17190# m3_13912_18146# 0.15fF
C6822 a_18026_7150# rowon_n[5] 0.14fF
C6823 a_2346_18236# col[8] 0.14fF
C6824 a_2346_1168# m2_7756_946# 0.19fF
C6825 a_3970_1126# m2_4744_946# 0.96fF
C6826 row_n[3] ctop 1.65fF
C6827 col_n[25] col[26] 5.88fF
C6828 a_8990_3134# a_9994_3134# 0.97fF
C6829 a_2346_3176# a_16930_3134# 0.35fF
C6830 a_30074_2130# m2_29844_946# 0.99fF
C6831 a_29070_11166# ctop 3.58fF
C6832 col[22] rowoff_n[11] 0.11fF
C6833 a_34090_12170# m3_34996_12122# 0.13fF
C6834 a_6982_17190# col_n[4] 0.28fF
C6835 a_27974_13174# a_28066_13174# 0.26fF
C6836 a_10998_13174# a_10998_12170# 1.00fF
C6837 a_2346_15224# col[0] 0.15fF
C6838 a_7986_4138# col[5] 0.29fF
C6839 a_17022_11166# rowoff_n[9] 0.10fF
C6840 a_9994_10162# vcm 0.62fF
C6841 a_1962_17230# a_3970_17190# 0.27fF
C6842 m2_11772_18014# m2_12200_18442# 0.16fF
C6843 a_1962_4178# col_n[14] 0.13fF
C6844 a_13006_3134# VDD 0.52fF
C6845 a_1962_17230# col_n[16] 0.13fF
C6846 a_2346_5184# a_29982_5142# 0.35fF
C6847 a_25054_13174# col_n[22] 0.28fF
C6848 a_27062_9158# rowoff_n[7] 0.10fF
C6849 a_3270_4178# vcm 0.22fF
C6850 a_1962_11206# col[7] 0.11fF
C6851 m2_14784_18014# col[12] 0.28fF
C6852 a_23046_14178# vcm 0.62fF
C6853 a_31078_15182# rowoff_n[13] 0.10fF
C6854 m2_34864_7974# VDD 1.00fF
C6855 a_1962_2170# a_24050_2130# 0.27fF
C6856 a_15014_7150# m2_15212_7398# 0.16fF
C6857 col[6] rowoff_n[12] 0.11fF
C6858 a_2966_8154# ctop 3.42fF
C6859 a_26058_7150# VDD 0.52fF
C6860 a_22042_7150# a_23046_7150# 0.97fF
C6861 a_15014_10162# row_n[8] 0.17fF
C6862 a_2346_10204# col[27] 0.15fF
C6863 a_1962_16226# a_10298_16226# 0.14fF
C6864 a_16322_8194# vcm 0.22fF
C6865 a_2346_16228# a_12002_16186# 0.19fF
C6866 a_24050_17190# a_24050_16186# 1.00fF
C6867 a_1962_12210# row_n[10] 25.57fF
C6868 a_2346_17232# vcm 0.39fF
C6869 a_7986_6146# col_n[5] 0.28fF
C6870 a_5886_10162# VDD 0.23fF
C6871 m2_1732_4962# ctop 0.17fF
C6872 a_29374_12210# vcm 0.22fF
C6873 a_4882_12170# rowoff_n[10] 0.24fF
C6874 m2_4744_946# col[2] 0.39fF
C6875 a_26058_2130# col_n[23] 0.28fF
C6876 a_1962_1166# a_30378_1166# 0.14fF
C6877 a_10998_6146# ctop 3.58fF
C6878 a_1962_13214# col_n[7] 0.13fF
C6879 a_34090_13174# row_n[11] 0.17fF
C6880 m3_34996_18146# VDD 0.46fF
C6881 m2_30848_18014# col_n[28] 0.25fF
C6882 a_23046_16186# col[20] 0.29fF
C6883 a_18938_14178# VDD 0.23fF
C6884 m2_9764_18014# ctop 0.18fF
C6885 a_18938_16186# rowoff_n[14] 0.24fF
C6886 a_23958_3134# a_24050_3134# 0.26fF
C6887 a_6982_3134# a_6982_2130# 1.00fF
C6888 a_12002_8154# m2_12200_8402# 0.16fF
C6889 a_24050_10162# ctop 3.58fF
C6890 a_26970_1126# m2_26832_946# 0.16fF
C6891 a_2346_6188# col[18] 0.15fF
C6892 a_31990_18194# VDD 0.33fF
C6893 a_2346_12212# a_14922_12170# 0.35fF
C6894 a_7986_12170# a_8990_12170# 0.97fF
C6895 a_22042_11166# rowon_n[9] 0.14fF
C6896 a_4974_9158# vcm 0.62fF
C6897 m2_7756_946# m3_8892_1078# 0.13fF
C6898 a_7986_2130# VDD 0.55fF
C6899 a_5978_9158# col[3] 0.29fF
C6900 a_1962_2170# col[25] 0.11fF
C6901 a_1962_9198# a_8990_9158# 0.27fF
C6902 a_1962_15222# col[27] 0.11fF
C6903 a_2346_14220# a_27974_14178# 0.35fF
C6904 a_18026_13174# vcm 0.62fF
C6905 a_24050_5142# col[21] 0.29fF
C6906 a_1962_9198# sample 0.14fF
C6907 a_21038_6146# VDD 0.52fF
C6908 a_2346_6188# a_3970_6146# 0.19fF
C6909 a_20034_7150# a_20034_6146# 1.00fF
C6910 a_2346_18236# col[19] 0.14fF
C6911 a_1962_11206# a_22042_11166# 0.27fF
C6912 a_1962_3174# row_n[1] 25.57fF
C6913 col_n[31] col[31] 0.91fF
C6914 m2_34864_17010# row_n[15] 0.15fF
C6915 a_11302_7190# vcm 0.22fF
C6916 a_21038_16186# a_22042_16186# 0.97fF
C6917 a_31078_17190# vcm 0.60fF
C6918 a_5978_17190# rowoff_n[15] 0.10fF
C6919 m2_29844_18014# VDD 0.93fF
C6920 a_9994_6146# rowoff_n[4] 0.10fF
C6921 a_2346_9200# m2_34864_8978# 0.17fF
C6922 a_8990_9158# m2_9188_9406# 0.16fF
C6923 a_34090_10162# VDD 0.54fF
C6924 a_2346_2172# col[9] 0.15fF
C6925 a_2346_15224# col[11] 0.15fF
C6926 a_1962_8194# a_15318_8194# 0.14fF
C6927 a_2346_8196# a_17022_8154# 0.19fF
C6928 a_9902_8154# a_9994_8154# 0.26fF
C6929 a_19030_14178# row_n[12] 0.17fF
C6930 a_5978_11166# col_n[3] 0.28fF
C6931 a_1962_4178# col_n[25] 0.13fF
C6932 a_34090_4138# row_n[2] 0.17fF
C6933 a_20034_4138# rowoff_n[2] 0.10fF
C6934 a_24354_11206# vcm 0.22fF
C6935 a_33086_12170# rowoff_n[10] 0.10fF
C6936 a_1962_17230# col_n[27] 0.13fF
C6937 a_5978_5142# ctop 3.58fF
C6938 a_1962_18234# col[1] 0.11fF
C6939 a_24050_7150# col_n[21] 0.28fF
C6940 a_13918_13174# VDD 0.23fF
C6941 a_1962_11206# col[18] 0.11fF
C6942 a_33086_11166# a_33086_10162# 1.00fF
C6943 a_1962_10202# a_28370_10202# 0.14fF
C6944 a_2346_10204# a_30074_10162# 0.19fF
C6945 a_30074_2130# rowoff_n[0] 0.10fF
C6946 m2_25828_946# vcm 0.42fF
C6947 col[17] rowoff_n[12] 0.11fF
C6948 a_6982_12170# rowon_n[10] 0.14fF
C6949 a_3970_2130# a_4974_2130# 0.97fF
C6950 a_2346_2172# a_6890_2130# 0.35fF
C6951 m2_21812_18014# m3_22948_18146# 0.13fF
C6952 a_19030_9158# ctop 3.58fF
C6953 a_26970_17190# VDD 0.24fF
C6954 a_22042_2130# rowon_n[0] 0.14fF
C6955 a_5978_12170# a_5978_11166# 1.00fF
C6956 a_22954_12170# a_23046_12170# 0.26fF
C6957 a_2874_1126# VDD 0.44fF
C6958 a_2346_4180# a_19942_4138# 0.35fF
C6959 a_5978_10162# m2_6176_10410# 0.16fF
C6960 a_32082_13174# ctop 3.58fF
C6961 a_2346_11208# col[2] 0.15fF
C6962 a_3970_17190# m2_3740_18014# 1.00fF
C6963 a_3970_14178# col[1] 0.29fF
C6964 a_18938_10162# rowoff_n[8] 0.24fF
C6965 col[1] rowoff_n[13] 0.11fF
C6966 a_26058_15182# rowon_n[13] 0.14fF
C6967 a_1962_13214# col_n[18] 0.13fF
C6968 a_13006_12170# vcm 0.62fF
C6969 a_20946_13174# rowoff_n[11] 0.24fF
C6970 m2_6752_946# VDD 0.62fF
C6971 a_16018_5142# VDD 0.52fF
C6972 a_17022_6146# a_18026_6146# 0.97fF
C6973 a_2346_6188# a_32994_6146# 0.35fF
C6974 a_22042_10162# col[19] 0.29fF
C6975 a_28978_8154# rowoff_n[6] 0.24fF
C6976 a_1962_7190# col[9] 0.11fF
C6977 a_3970_15182# row_n[13] 0.17fF
C6978 a_6282_6186# vcm 0.22fF
C6979 a_19030_16186# a_19030_15182# 1.00fF
C6980 a_35002_17190# rowoff_n[15] 0.24fF
C6981 a_26058_16186# vcm 0.62fF
C6982 a_2346_6188# col[29] 0.15fF
C6983 a_1962_3174# a_27062_3134# 0.27fF
C6984 a_19030_5142# row_n[3] 0.17fF
C6985 a_29070_9158# VDD 0.52fF
C6986 a_19334_10202# vcm 0.22fF
C6987 a_2346_17232# a_15014_17190# 0.19fF
C6988 a_8898_17190# a_8990_17190# 0.26fF
C6989 a_1962_17230# a_13310_17230# 0.14fF
C6990 a_3970_16186# col_n[1] 0.28fF
C6991 a_4974_3134# col[2] 0.29fF
C6992 m3_1864_16138# ctop 0.23fF
C6993 a_8898_12170# VDD 0.23fF
C6994 a_30074_10162# a_31078_10162# 0.97fF
C6995 a_22042_12170# col_n[19] 0.28fF
C6996 a_6982_3134# rowon_n[1] 0.14fF
C6997 a_1962_9198# col_n[9] 0.13fF
C6998 a_32386_14218# vcm 0.22fF
C6999 a_7986_14178# rowoff_n[12] 0.10fF
C7000 a_1962_2170# a_33390_2170# 0.14fF
C7001 a_18938_2130# a_19030_2130# 0.26fF
C7002 a_14010_8154# ctop 3.58fF
C7003 m2_34864_16006# m3_34996_16138# 2.76fF
C7004 a_2966_6146# VDD 0.56fF
C7005 a_2346_18236# col[30] 0.14fF
C7006 a_1962_3174# col[0] 0.11fF
C7007 col[0] col[1] 0.20fF
C7008 ctop col[7] 1.98fF
C7009 a_1962_16226# col[2] 0.11fF
C7010 a_21950_16186# VDD 0.23fF
C7011 a_2346_11208# a_4882_11166# 0.35fF
C7012 a_9994_2130# m2_10192_2378# 0.16fF
C7013 a_2346_2172# col[20] 0.15fF
C7014 a_31990_1126# VDD 0.44fF
C7015 a_10998_16186# rowon_n[14] 0.14fF
C7016 a_2346_15224# col[22] 0.15fF
C7017 a_27062_12170# ctop 3.58fF
C7018 a_23046_17190# m2_22816_18014# 1.00fF
C7019 a_4974_5142# col_n[2] 0.28fF
C7020 a_26058_6146# rowon_n[4] 0.14fF
C7021 a_2346_13216# a_17934_13174# 0.35fF
C7022 a_7986_11166# vcm 0.62fF
C7023 a_1962_18234# col[12] 0.11fF
C7024 a_10998_4138# VDD 0.52fF
C7025 a_1962_11206# col[29] 0.11fF
C7026 m3_10900_1078# VDD 0.14fF
C7027 a_31990_6146# a_32082_6146# 0.26fF
C7028 a_34090_13174# m2_34288_13422# 0.16fF
C7029 a_15014_6146# a_15014_5142# 1.00fF
C7030 a_3970_6146# row_n[4] 0.17fF
C7031 a_1962_10202# a_12002_10162# 0.27fF
C7032 col[28] rowoff_n[12] 0.11fF
C7033 a_20034_15182# col[17] 0.29fF
C7034 a_1962_5182# vcm 6.95fF
C7035 a_2346_15224# a_30986_15182# 0.35fF
C7036 a_16018_15182# a_17022_15182# 0.97fF
C7037 a_21038_15182# vcm 0.62fF
C7038 m2_1732_10986# VDD 1.02fF
C7039 a_35002_1126# m2_34864_946# 0.16fF
C7040 a_24050_8154# VDD 0.52fF
C7041 a_4882_7150# a_4974_7150# 0.26fF
C7042 a_1962_7190# a_5278_7190# 0.14fF
C7043 a_2346_7192# a_6982_7150# 0.19fF
C7044 a_1962_12210# a_25054_12170# 0.27fF
C7045 a_14314_9198# vcm 0.22fF
C7046 a_11910_5142# rowoff_n[3] 0.24fF
C7047 a_2346_11208# col[13] 0.15fF
C7048 a_23046_9158# row_n[7] 0.17fF
C7049 m2_28840_946# m3_29976_1078# 0.13fF
C7050 a_1962_9198# a_18330_9198# 0.14fF
C7051 a_28066_10162# a_28066_9158# 1.00fF
C7052 a_2346_9200# a_20034_9158# 0.19fF
C7053 col[12] rowoff_n[13] 0.11fF
C7054 a_1962_13214# col_n[29] 0.13fF
C7055 a_21950_3134# rowoff_n[1] 0.24fF
C7056 a_27366_13214# vcm 0.22fF
C7057 a_20034_17190# col_n[17] 0.28fF
C7058 a_1962_7190# col[20] 0.11fF
C7059 m2_34864_12994# m3_34996_13126# 2.76fF
C7060 a_8990_7150# ctop 3.58fF
C7061 a_21038_4138# col[18] 0.29fF
C7062 a_31078_14178# m2_31276_14426# 0.16fF
C7063 a_16930_15182# VDD 0.23fF
C7064 a_17934_11166# a_18026_11166# 0.26fF
C7065 a_1962_11206# a_31382_11206# 0.14fF
C7066 a_2346_11208# a_33086_11166# 0.19fF
C7067 a_10998_7150# rowon_n[5] 0.14fF
C7068 m2_1732_11990# m2_2160_12418# 0.16fF
C7069 a_2346_3176# a_9902_3134# 0.35fF
C7070 a_22042_11166# ctop 3.58fF
C7071 a_2346_16228# m2_1732_16006# 0.12fF
C7072 a_9994_11166# rowoff_n[9] 0.10fF
C7073 a_2346_7192# col[4] 0.15fF
C7074 m2_4744_18014# m2_5172_18442# 0.16fF
C7075 a_5978_3134# VDD 0.52fF
C7076 a_12002_5142# a_13006_5142# 0.97fF
C7077 a_2346_5184# a_22954_5142# 0.35fF
C7078 a_1962_9198# col_n[20] 0.13fF
C7079 a_30074_10162# rowon_n[8] 0.14fF
C7080 a_20034_9158# rowoff_n[7] 0.10fF
C7081 a_21038_6146# col_n[18] 0.28fF
C7082 a_30986_15182# a_31078_15182# 0.26fF
C7083 a_14010_15182# a_14010_14178# 1.00fF
C7084 a_16018_14178# vcm 0.62fF
C7085 a_24050_15182# rowoff_n[13] 0.10fF
C7086 a_1962_2170# a_17022_2130# 0.27fF
C7087 a_1962_3174# col[11] 0.11fF
C7088 a_1962_16226# col[13] 0.11fF
C7089 m2_1732_17010# m3_1864_16138# 0.15fF
C7090 ctop col[18] 1.98fF
C7091 a_19030_7150# VDD 0.52fF
C7092 a_30074_7150# rowoff_n[5] 0.10fF
C7093 a_28066_15182# m2_28264_15430# 0.16fF
C7094 a_7986_10162# row_n[8] 0.17fF
C7095 a_3878_16186# VDD 0.23fF
C7096 a_2966_13174# col[0] 0.29fF
C7097 a_2346_2172# col[31] 0.15fF
C7098 a_9294_8194# vcm 0.22fF
C7099 a_2346_16228# a_4974_16186# 0.19fF
C7100 a_1962_16226# a_3270_16226# 0.14fF
C7101 a_30074_3134# m2_30272_3382# 0.16fF
C7102 m2_34864_16006# m2_34864_15002# 0.99fF
C7103 a_29070_18194# vcm 0.12fF
C7104 a_1962_4178# a_30074_4138# 0.27fF
C7105 a_32082_11166# VDD 0.52fF
C7106 m3_31984_1078# m3_32988_1078# 0.22fF
C7107 a_25054_9158# a_26058_9158# 0.97fF
C7108 a_1962_18234# col[23] 0.11fF
C7109 a_22346_12210# vcm 0.22fF
C7110 a_1962_1166# a_23350_1166# 0.14fF
C7111 m2_34864_9982# m3_34996_10114# 2.76fF
C7112 a_3970_6146# ctop 3.57fF
C7113 a_27062_13174# row_n[11] 0.17fF
C7114 m3_6884_18146# VDD 0.36fF
C7115 a_11910_14178# VDD 0.23fF
C7116 a_1962_5182# col_n[11] 0.13fF
C7117 m2_27836_946# col[25] 0.39fF
C7118 a_19030_9158# col[16] 0.29fF
C7119 a_11910_16186# rowoff_n[14] 0.24fF
C7120 a_2966_15182# vcm 0.61fF
C7121 a_1962_12210# col[4] 0.11fF
C7122 a_2346_17232# row_n[15] 0.35fF
C7123 a_17022_10162# ctop 3.58fF
C7124 a_25054_16186# m2_25252_16434# 0.16fF
C7125 a_24962_18194# VDD 0.33fF
C7126 m2_24824_18014# vcm 0.28fF
C7127 a_2346_12212# a_7894_12170# 0.35fF
C7128 a_15014_11166# rowon_n[9] 0.14fF
C7129 a_2346_11208# col[24] 0.15fF
C7130 a_27062_4138# m2_27260_4386# 0.16fF
C7131 a_35002_3134# VDD 0.29fF
C7132 m3_13912_1078# ctop 0.23fF
C7133 col[23] rowoff_n[13] 0.11fF
C7134 a_26970_5142# a_27062_5142# 0.26fF
C7135 a_9994_5142# a_9994_4138# 1.00fF
C7136 a_1962_13214# rowon_n[11] 1.18fF
C7137 a_30074_14178# ctop 3.58fF
C7138 sample_n rowoff_n[0] 0.38fF
C7139 vcm rowoff_n[3] 0.20fF
C7140 a_2346_14220# a_20946_14178# 0.35fF
C7141 a_10998_14178# a_12002_14178# 0.97fF
C7142 a_3878_3134# rowoff_n[1] 0.24fF
C7143 a_2346_18236# a_29982_18194# 0.35fF
C7144 a_1962_7190# col[31] 0.11fF
C7145 a_10998_13174# vcm 0.62fF
C7146 a_19030_11166# col_n[16] 0.28fF
C7147 m2_1732_13998# m3_1864_13126# 0.15fF
C7148 a_14010_6146# VDD 0.52fF
C7149 a_1962_1166# col_n[2] 0.13fF
C7150 a_1962_14218# col_n[4] 0.13fF
C7151 a_1962_11206# a_15014_11166# 0.27fF
C7152 a_34090_14178# rowon_n[12] 0.14fF
C7153 a_2346_16228# a_33998_16186# 0.35fF
C7154 a_4274_7190# vcm 0.22fF
C7155 a_24050_17190# vcm 0.60fF
C7156 col[7] rowoff_n[14] 0.11fF
C7157 m2_15788_18014# VDD 1.05fF
C7158 a_1962_18234# m2_30848_18014# 0.18fF
C7159 a_2874_6146# rowoff_n[4] 0.24fF
C7160 a_27062_10162# VDD 0.52fF
C7161 a_2346_8196# a_9994_8154# 0.19fF
C7162 a_23046_9158# a_23046_8154# 1.00fF
C7163 a_22042_17190# m2_22240_17438# 0.16fF
C7164 a_1962_8194# a_8290_8194# 0.14fF
C7165 a_12002_14178# row_n[12] 0.17fF
C7166 a_1962_13214# a_28066_13174# 0.27fF
C7167 a_34090_2130# vcm 0.62fF
C7168 a_2346_7192# col[15] 0.15fF
C7169 a_17326_11206# vcm 0.22fF
C7170 a_26058_12170# rowoff_n[10] 0.10fF
C7171 a_27062_4138# row_n[2] 0.17fF
C7172 a_13006_4138# rowoff_n[2] 0.10fF
C7173 a_24050_5142# m2_24248_5390# 0.16fF
C7174 m2_34864_6970# m3_34996_7102# 2.76fF
C7175 a_1962_9198# col_n[31] 0.13fF
C7176 a_2966_5142# a_3970_5142# 0.97fF
C7177 a_2346_18236# m2_25828_18014# 0.19fF
C7178 a_6890_13174# VDD 0.23fF
C7179 a_1962_10202# a_21342_10202# 0.14fF
C7180 a_12914_10162# a_13006_10162# 0.26fF
C7181 a_2346_10204# a_23046_10162# 0.19fF
C7182 a_23046_2130# rowoff_n[0] 0.10fF
C7183 a_1962_3174# col[22] 0.11fF
C7184 vcm col_n[3] 2.80fF
C7185 VDD col_n[7] 4.95fF
C7186 a_2346_8196# row_n[6] 0.35fF
C7187 col[11] col[12] 0.20fF
C7188 a_1962_16226# col[24] 0.11fF
C7189 ctop col[29] 1.98fF
C7190 m2_34864_17010# ctop 0.17fF
C7191 a_30378_15222# vcm 0.22fF
C7192 a_17022_14178# col[14] 0.29fF
C7193 a_31078_17190# row_n[15] 0.17fF
C7194 a_12002_9158# ctop 3.58fF
C7195 m2_12776_18014# m3_12908_18146# 2.78fF
C7196 a_15014_2130# rowon_n[0] 0.14fF
C7197 a_19942_17190# VDD 0.24fF
C7198 a_1962_12210# a_35398_12210# 0.14fF
C7199 a_2346_12212# a_2346_11208# 0.22fF
C7200 a_1962_4178# rowon_n[2] 1.18fF
C7201 a_29982_2130# VDD 0.23fF
C7202 a_2346_4180# a_12914_4138# 0.35fF
C7203 a_6982_4138# a_7986_4138# 0.97fF
C7204 a_25054_13174# ctop 3.58fF
C7205 m3_34996_4090# m3_34996_3086# 0.22fF
C7206 a_21950_18194# m2_21812_18014# 0.16fF
C7207 a_25966_14178# a_26058_14178# 0.26fF
C7208 a_8990_14178# a_8990_13174# 1.00fF
C7209 a_2346_3176# col[6] 0.15fF
C7210 a_11910_10162# rowoff_n[8] 0.24fF
C7211 a_2346_16228# col[8] 0.15fF
C7212 a_19030_15182# rowon_n[13] 0.14fF
C7213 a_5978_12170# vcm 0.62fF
C7214 a_13918_13174# rowoff_n[11] 0.24fF
C7215 a_21038_6146# m2_21236_6394# 0.16fF
C7216 m2_1732_10986# m3_1864_10114# 0.15fF
C7217 a_8990_5142# VDD 0.52fF
C7218 a_1962_5182# col_n[22] 0.13fF
C7219 a_34090_5142# rowon_n[3] 0.14fF
C7220 a_2346_6188# a_25966_6146# 0.35fF
C7221 a_17022_16186# col_n[14] 0.28fF
C7222 a_21950_8154# rowoff_n[6] 0.24fF
C7223 a_18026_3134# col[15] 0.29fF
C7224 a_17022_17190# m3_16924_18146# 0.15fF
C7225 a_1962_12210# col[15] 0.11fF
C7226 a_19030_16186# vcm 0.62fF
C7227 a_27974_17190# rowoff_n[15] 0.24fF
C7228 a_31990_6146# rowoff_n[4] 0.24fF
C7229 a_12002_5142# row_n[3] 0.17fF
C7230 a_1962_3174# a_20034_3134# 0.27fF
C7231 a_1962_1166# m2_24824_946# 0.18fF
C7232 a_22042_9158# VDD 0.52fF
C7233 a_20034_8154# a_21038_8154# 0.97fF
C7234 a_29070_1126# vcm 0.12fF
C7235 a_2346_17232# a_7986_17190# 0.19fF
C7236 a_12306_10202# vcm 0.22fF
C7237 a_1962_17230# a_6282_17230# 0.14fF
C7238 m2_34864_3958# m3_34996_4090# 2.76fF
C7239 m3_9896_18146# ctop 0.23fF
C7240 a_1962_5182# a_33086_5142# 0.27fF
C7241 a_2346_14220# a_1962_14218# 2.62fF
C7242 a_31078_8154# row_n[6] 0.17fF
C7243 a_25358_14218# vcm 0.22fF
C7244 a_18026_5142# col_n[15] 0.28fF
C7245 a_2346_2172# a_28066_2130# 0.19fF
C7246 a_32082_3134# a_32082_2130# 1.00fF
C7247 a_18026_7150# m2_18224_7398# 0.16fF
C7248 a_1962_2170# a_26362_2170# 0.14fF
C7249 a_1962_1166# col_n[13] 0.13fF
C7250 a_6982_8154# ctop 3.58fF
C7251 a_1962_14218# col_n[15] 0.13fF
C7252 a_14922_16186# VDD 0.23fF
C7253 a_33086_12170# a_34090_12170# 0.97fF
C7254 a_1962_8194# col[6] 0.11fF
C7255 col[18] rowoff_n[14] 0.11fF
C7256 a_3970_16186# rowon_n[14] 0.14fF
C7257 a_24962_1126# VDD 0.44fF
C7258 a_21950_4138# a_22042_4138# 0.26fF
C7259 a_33086_15182# col[30] 0.29fF
C7260 a_4974_4138# a_4974_3134# 1.00fF
C7261 a_20034_12170# ctop 3.58fF
C7262 a_2346_7192# col[26] 0.15fF
C7263 a_19030_6146# rowon_n[4] 0.14fF
C7264 a_5978_13174# a_6982_13174# 0.97fF
C7265 a_2346_13216# a_10906_13174# 0.35fF
C7266 m2_1732_7974# m3_1864_7102# 0.15fF
C7267 a_3970_4138# VDD 0.52fF
C7268 m3_1864_10114# VDD 0.25fF
C7269 a_33086_16186# ctop 3.56fF
C7270 a_3878_10162# a_3970_10162# 0.26fF
C7271 a_1962_10202# a_4974_10162# 0.27fF
C7272 VDD col_n[18] 4.94fF
C7273 vcm col_n[14] 2.80fF
C7274 col[2] rowoff_n[15] 0.11fF
C7275 a_2346_15224# a_23958_15182# 0.35fF
C7276 a_16018_8154# col[13] 0.29fF
C7277 a_14010_15182# vcm 0.62fF
C7278 a_15014_8154# m2_15212_8402# 0.16fF
C7279 a_1962_10202# col_n[6] 0.13fF
C7280 a_17022_8154# VDD 0.52fF
C7281 a_18026_8154# a_18026_7150# 1.00fF
C7282 a_35494_18556# VDD 0.12fF
C7283 a_33086_17190# col_n[30] 0.28fF
C7284 m2_8760_18014# col[6] 0.28fF
C7285 a_1962_12210# a_18026_12170# 0.27fF
C7286 a_34090_4138# col[31] 0.29fF
C7287 a_7286_9198# vcm 0.22fF
C7288 a_19030_17190# a_20034_17190# 0.97fF
C7289 a_1962_17230# a_1962_16226# 0.16fF
C7290 a_4882_5142# rowoff_n[3] 0.24fF
C7291 a_16018_9158# row_n[7] 0.17fF
C7292 a_30074_12170# VDD 0.52fF
C7293 a_2346_3176# col[17] 0.15fF
C7294 m3_27968_18146# m3_28972_18146# 0.22fF
C7295 a_7894_9158# a_7986_9158# 0.26fF
C7296 a_2346_9200# a_13006_9158# 0.19fF
C7297 a_1962_9198# a_11302_9198# 0.14fF
C7298 a_2346_16228# col[19] 0.15fF
C7299 m2_34864_7974# row_n[6] 0.15fF
C7300 a_1962_14218# a_31078_14178# 0.27fF
C7301 a_14922_3134# rowoff_n[1] 0.24fF
C7302 a_29982_14178# rowoff_n[12] 0.24fF
C7303 a_20338_13214# vcm 0.22fF
C7304 a_29070_2130# a_30074_2130# 0.97fF
C7305 a_16018_10162# col_n[13] 0.28fF
C7306 a_9902_15182# VDD 0.23fF
C7307 a_3878_8154# rowoff_n[6] 0.24fF
C7308 a_2346_11208# a_26058_11166# 0.19fF
C7309 a_1962_11206# a_24354_11206# 0.14fF
C7310 a_31078_12170# a_31078_11166# 1.00fF
C7311 a_1962_12210# col[26] 0.11fF
C7312 m2_14784_946# a_15014_2130# 0.99fF
C7313 a_3970_7150# rowon_n[5] 0.14fF
C7314 a_33390_17230# vcm 0.22fF
C7315 m2_24824_18014# col_n[22] 0.25fF
C7316 a_34090_6146# col_n[31] 0.28fF
C7317 a_12002_9158# m2_12200_9406# 0.16fF
C7318 a_15014_11166# ctop 3.58fF
C7319 a_3970_13174# a_3970_12170# 1.00fF
C7320 a_20946_13174# a_21038_13174# 0.26fF
C7321 a_2874_11166# rowoff_n[9] 0.24fF
C7322 m2_1732_4962# m3_1864_4090# 0.15fF
C7323 a_32994_4138# VDD 0.23fF
C7324 a_2346_5184# a_15926_5142# 0.35fF
C7325 a_28066_15182# ctop 3.58fF
C7326 a_2346_12212# col[10] 0.15fF
C7327 a_23046_10162# rowon_n[8] 0.14fF
C7328 a_13006_9158# rowoff_n[7] 0.10fF
C7329 a_1962_1166# col_n[24] 0.13fF
C7330 a_17022_15182# rowoff_n[13] 0.10fF
C7331 a_8990_14178# vcm 0.62fF
C7332 a_1962_14218# col_n[26] 0.13fF
C7333 a_1962_2170# a_9994_2130# 0.27fF
C7334 m2_26832_18014# m3_27968_18146# 0.13fF
C7335 a_12002_7150# VDD 0.52fF
C7336 a_23046_7150# rowoff_n[5] 0.10fF
C7337 a_2346_7192# a_28978_7150# 0.35fF
C7338 a_15014_7150# a_16018_7150# 0.97fF
C7339 a_14010_13174# col[11] 0.29fF
C7340 col[29] rowoff_n[14] 0.11fF
C7341 a_1962_8194# col[17] 0.11fF
C7342 a_17022_17190# a_17022_16186# 1.00fF
C7343 a_33998_17190# a_34090_17190# 0.26fF
C7344 a_33086_5142# rowoff_n[3] 0.10fF
C7345 a_22042_18194# vcm 0.12fF
C7346 a_32082_9158# col[29] 0.29fF
C7347 a_8990_10162# m2_9188_10410# 0.16fF
C7348 a_1962_4178# a_23046_4138# 0.27fF
C7349 a_2346_10204# m2_34864_9982# 0.17fF
C7350 a_25054_11166# VDD 0.52fF
C7351 m3_34996_2082# m3_34996_1078# 0.22fF
C7352 a_32082_3134# vcm 0.62fF
C7353 a_15318_12210# vcm 0.22fF
C7354 a_1962_1166# a_16322_1166# 0.14fF
C7355 a_2346_1168# a_18026_1126# 0.19fF
C7356 a_20034_13174# row_n[11] 0.17fF
C7357 col_n[12] col_n[13] 0.10fF
C7358 vcm col_n[25] 2.80fF
C7359 VDD col_n[29] 4.96fF
C7360 col[22] col[23] 0.20fF
C7361 col[13] rowoff_n[15] 0.11fF
C7362 a_2346_8196# col[1] 0.15fF
C7363 a_4882_14178# VDD 0.23fF
C7364 a_28066_11166# a_29070_11166# 0.97fF
C7365 m2_11772_946# a_11910_1126# 0.16fF
C7366 VDD rowoff_n[11] 1.17fF
C7367 a_14010_15182# col_n[11] 0.28fF
C7368 a_1962_10202# col_n[17] 0.13fF
C7369 a_15014_2130# col[12] 0.29fF
C7370 a_28370_16226# vcm 0.22fF
C7371 a_4882_16186# rowoff_n[14] 0.24fF
C7372 m2_13780_946# m2_14784_946# 0.96fF
C7373 a_16930_3134# a_17022_3134# 0.26fF
C7374 a_1962_3174# a_29374_3174# 0.14fF
C7375 a_2346_3176# a_31078_3134# 0.19fF
C7376 a_9994_10162# ctop 3.58fF
C7377 a_1962_4178# col[8] 0.11fF
C7378 a_32082_11166# col_n[29] 0.28fF
C7379 a_17934_18194# VDD 0.33fF
C7380 a_1962_17230# col[10] 0.11fF
C7381 m2_10768_18014# vcm 0.28fF
C7382 a_7986_11166# rowon_n[9] 0.14fF
C7383 a_31990_11166# rowoff_n[9] 0.24fF
C7384 m2_2736_1950# m3_1864_2082# 0.13fF
C7385 a_2346_3176# col[28] 0.15fF
C7386 a_27974_3134# VDD 0.23fF
C7387 m3_34996_9110# ctop 0.23fF
C7388 a_2346_16228# col[30] 0.15fF
C7389 a_5978_11166# m2_6176_11414# 0.16fF
C7390 a_23046_14178# ctop 3.58fF
C7391 m2_30848_946# m2_31852_946# 0.96fF
C7392 a_2346_14220# a_13918_14178# 0.35fF
C7393 a_2346_18236# a_22954_18194# 0.35fF
C7394 a_3970_13174# vcm 0.62fF
C7395 a_6982_6146# VDD 0.52fF
C7396 a_15014_4138# col_n[12] 0.28fF
C7397 a_13006_7150# a_13006_6146# 1.00fF
C7398 a_29982_7150# a_30074_7150# 0.26fF
C7399 a_2346_17232# ctop 1.30fF
C7400 a_27062_14178# rowon_n[12] 0.14fF
C7401 a_1962_11206# a_7986_11166# 0.27fF
C7402 a_2346_16228# a_26970_16186# 0.35fF
C7403 a_14010_16186# a_15014_16186# 0.97fF
C7404 a_1962_6186# col_n[8] 0.13fF
C7405 a_13006_2130# m2_13204_2378# 0.16fF
C7406 a_17022_17190# vcm 0.60fF
C7407 m2_1732_18014# VDD 1.37fF
C7408 a_1962_18234# m2_16792_18014# 0.18fF
C7409 a_20034_10162# VDD 0.52fF
C7410 a_2346_8196# a_2874_8154# 0.35fF
C7411 a_4974_14178# row_n[12] 0.17fF
C7412 a_30074_14178# col[27] 0.29fF
C7413 a_1962_13214# col[1] 0.11fF
C7414 a_27062_2130# vcm 0.62fF
C7415 a_1962_13214# a_21038_13174# 0.27fF
C7416 a_10298_11206# vcm 0.22fF
C7417 a_19030_12170# rowoff_n[10] 0.10fF
C7418 a_20034_4138# row_n[2] 0.17fF
C7419 a_5978_4138# rowoff_n[2] 0.10fF
C7420 a_2346_12212# col[21] 0.15fF
C7421 m3_25960_1078# VDD 0.14fF
C7422 a_33086_14178# VDD 0.52fF
C7423 a_2346_18236# m2_11772_18014# 0.19fF
C7424 a_26058_11166# a_26058_10162# 1.00fF
C7425 a_2346_10204# a_16018_10162# 0.19fF
C7426 a_1962_10202# a_14314_10202# 0.14fF
C7427 a_16018_2130# rowoff_n[0] 0.10fF
C7428 a_1962_15222# a_34090_15182# 0.27fF
C7429 a_33086_16186# rowoff_n[14] 0.10fF
C7430 a_23350_15222# vcm 0.22fF
C7431 m2_11772_946# col_n[9] 0.37fF
C7432 m2_3740_18014# m3_2868_18146# 0.13fF
C7433 a_4974_9158# ctop 3.58fF
C7434 a_24050_17190# row_n[15] 0.17fF
C7435 a_1962_8194# col[28] 0.11fF
C7436 a_13006_7150# col[10] 0.29fF
C7437 a_7986_2130# rowon_n[0] 0.14fF
C7438 a_12914_17190# VDD 0.24fF
C7439 a_15926_12170# a_16018_12170# 0.26fF
C7440 a_1962_12210# a_27366_12210# 0.14fF
C7441 a_2346_12212# a_29070_12170# 0.19fF
C7442 a_1962_2170# col_n[0] 0.13fF
C7443 a_30074_16186# col_n[27] 0.28fF
C7444 a_1962_15222# col_n[1] 0.13fF
C7445 a_31078_3134# col[28] 0.29fF
C7446 a_22954_2130# VDD 0.23fF
C7447 a_2346_4180# a_5886_4138# 0.35fF
C7448 a_18026_13174# ctop 3.58fF
C7449 m2_33860_946# m3_34568_1078# 0.82fF
C7450 m3_34996_11118# m3_34996_10114# 0.22fF
C7451 a_4882_10162# rowoff_n[8] 0.24fF
C7452 a_12002_15182# rowon_n[13] 0.14fF
C7453 a_6890_13174# rowoff_n[11] 0.24fF
C7454 VDD rowon_n[11] 2.61fF
C7455 col_n[1] row_n[14] 0.23fF
C7456 col_n[3] row_n[15] 0.23fF
C7457 vcm rowon_n[13] 0.50fF
C7458 col_n[0] row_n[13] 0.23fF
C7459 a_2346_8196# col[12] 0.15fF
C7460 col[24] rowoff_n[15] 0.11fF
C7461 a_27062_5142# rowon_n[3] 0.14fF
C7462 a_9994_6146# a_10998_6146# 0.97fF
C7463 a_2346_6188# a_18938_6146# 0.35fF
C7464 a_34090_14178# m2_34288_14426# 0.16fF
C7465 a_31078_17190# ctop 3.39fF
C7466 a_14922_8154# rowoff_n[6] 0.24fF
C7467 a_1962_10202# col_n[28] 0.13fF
C7468 a_13006_9158# col_n[10] 0.28fF
C7469 a_12002_16186# a_12002_15182# 1.00fF
C7470 a_28978_16186# a_29070_16186# 0.26fF
C7471 a_20946_17190# rowoff_n[15] 0.24fF
C7472 a_12002_16186# vcm 0.62fF
C7473 a_1962_3174# a_13006_3134# 0.27fF
C7474 a_24962_6146# rowoff_n[4] 0.24fF
C7475 a_4974_5142# row_n[3] 0.17fF
C7476 a_1962_4178# col[19] 0.11fF
C7477 a_5978_2130# m3_5880_1078# 0.15fF
C7478 a_2346_9200# rowon_n[7] 0.26fF
C7479 a_15014_9158# VDD 0.52fF
C7480 a_1962_17230# col[21] 0.11fF
C7481 a_2346_8196# a_31990_8154# 0.35fF
C7482 a_31078_5142# col_n[28] 0.28fF
C7483 a_22042_1126# vcm 0.12fF
C7484 m2_2736_946# m2_3164_1374# 0.16fF
C7485 a_5278_10202# vcm 0.22fF
C7486 a_35002_4138# rowoff_n[2] 0.24fF
C7487 m2_25828_946# ctop 0.18fF
C7488 a_1962_5182# a_26058_5142# 0.27fF
C7489 a_28066_13174# VDD 0.52fF
C7490 a_23046_10162# a_24050_10162# 0.97fF
C7491 a_35094_5142# vcm 0.12fF
C7492 a_24050_8154# row_n[6] 0.17fF
C7493 a_18330_14218# vcm 0.22fF
C7494 a_2346_4180# col[3] 0.15fF
C7495 a_2346_2172# a_21038_2130# 0.19fF
C7496 a_1962_2170# a_19334_2170# 0.14fF
C7497 a_11910_2130# a_12002_2130# 0.26fF
C7498 a_2346_17232# col[5] 0.15fF
C7499 a_31078_15182# m2_31276_15430# 0.16fF
C7500 a_7894_16186# VDD 0.23fF
C7501 a_1962_6186# col_n[19] 0.13fF
C7502 m2_34864_12994# vcm 0.51fF
C7503 a_10998_12170# col[8] 0.29fF
C7504 a_33086_3134# m2_33284_3382# 0.16fF
C7505 a_31382_18234# vcm 0.22fF
C7506 a_17934_1126# VDD 0.39fF
C7507 a_1962_4178# a_32386_4178# 0.14fF
C7508 a_2346_4180# a_34090_4138# 0.19fF
C7509 a_1962_13214# col[12] 0.11fF
C7510 m2_34864_9982# rowon_n[8] 0.13fF
C7511 a_13006_12170# ctop 3.58fF
C7512 rowon_n[7] rowoff_n[7] 20.27fF
C7513 a_2346_17232# m2_1732_17010# 0.12fF
C7514 a_29070_8154# col[26] 0.29fF
C7515 a_12002_6146# rowon_n[4] 0.14fF
C7516 a_1962_13214# a_2966_13174# 0.27fF
C7517 a_33086_10162# rowoff_n[8] 0.10fF
C7518 a_30986_5142# VDD 0.23fF
C7519 m3_21944_18146# VDD 0.25fF
C7520 a_24962_6146# a_25054_6146# 0.26fF
C7521 a_7986_6146# a_7986_5142# 1.00fF
C7522 a_26058_16186# ctop 3.57fF
C7523 m2_19228_1374# a_19030_1126# 0.16fF
C7524 a_2346_15224# a_16930_15182# 0.35fF
C7525 a_8990_15182# a_9994_15182# 0.97fF
C7526 a_6982_15182# vcm 0.62fF
C7527 a_10998_14178# col_n[8] 0.28fF
C7528 a_31078_9158# rowon_n[7] 0.14fF
C7529 a_9994_8154# VDD 0.52fF
C7530 a_28066_16186# m2_28264_16434# 0.16fF
C7531 a_1962_2170# col_n[10] 0.13fF
C7532 a_1962_12210# a_10998_12170# 0.27fF
C7533 a_1962_15222# col_n[12] 0.13fF
C7534 a_1962_18234# a_35398_18234# 0.14fF
C7535 m2_1732_3958# sample 0.19fF
C7536 a_29070_10162# col_n[26] 0.28fF
C7537 a_2346_17232# a_29982_17190# 0.35fF
C7538 m2_1732_15002# sample_n 0.15fF
C7539 a_30074_4138# m2_30272_4386# 0.16fF
C7540 a_2966_12170# col_n[0] 0.28fF
C7541 m3_28972_1078# ctop 0.23fF
C7542 a_8990_9158# row_n[7] 0.17fF
C7543 a_1962_9198# col[3] 0.11fF
C7544 a_23046_12170# VDD 0.52fF
C7545 m3_13912_18146# m3_14916_18146# 0.22fF
C7546 a_1962_9198# a_4274_9198# 0.14fF
C7547 a_2346_9200# a_5978_9158# 0.19fF
C7548 a_21038_10162# a_21038_9158# 1.00fF
C7549 m2_1732_11990# row_n[10] 0.13fF
C7550 a_30074_4138# vcm 0.62fF
C7551 a_1962_14218# a_24050_14178# 0.27fF
C7552 a_7894_3134# rowoff_n[1] 0.24fF
C7553 col_n[8] row_n[12] 0.23fF
C7554 col_n[14] row_n[15] 0.23fF
C7555 vcm row_n[8] 0.49fF
C7556 col_n[6] row_n[11] 0.23fF
C7557 col_n[4] row_n[10] 0.23fF
C7558 col_n[12] row_n[14] 0.23fF
C7559 col_n[23] col_n[24] 0.10fF
C7560 sample row_n[7] 1.03fF
C7561 col_n[10] row_n[13] 0.23fF
C7562 col_n[2] row_n[9] 0.23fF
C7563 VDD row_n[6] 2.93fF
C7564 m2_34864_6970# m2_35292_7398# 0.16fF
C7565 a_2346_8196# col[23] 0.15fF
C7566 a_22954_14178# rowoff_n[12] 0.24fF
C7567 a_13310_13214# vcm 0.22fF
C7568 a_2346_15224# VDD 32.63fF
C7569 a_1962_11206# a_17326_11206# 0.14fF
C7570 a_10906_11166# a_10998_11166# 0.26fF
C7571 a_2346_11208# a_19030_11166# 0.19fF
C7572 a_12002_3134# col_n[9] 0.28fF
C7573 a_1962_4178# col[30] 0.11fF
C7574 a_28066_12170# row_n[10] 0.17fF
C7575 a_8990_17190# col[6] 0.29fF
C7576 a_26362_17230# vcm 0.22fF
C7577 a_32082_4138# a_33086_4138# 0.97fF
C7578 a_7986_11166# ctop 3.58fF
C7579 a_25054_17190# m2_25252_17438# 0.16fF
C7580 a_1962_11206# col_n[3] 0.13fF
C7581 a_34090_14178# a_34090_13174# 1.00fF
C7582 a_1962_13214# a_30378_13214# 0.14fF
C7583 a_2346_13216# a_32082_13174# 0.19fF
C7584 a_27062_13174# col[24] 0.29fF
C7585 a_27062_5142# m2_27260_5390# 0.16fF
C7586 a_1962_5182# ctop 1.49fF
C7587 a_25966_4138# VDD 0.23fF
C7588 a_2346_5184# a_8898_5142# 0.35fF
C7589 a_4974_5142# a_5978_5142# 0.97fF
C7590 a_21038_15182# ctop 3.58fF
C7591 a_16018_10162# rowon_n[8] 0.14fF
C7592 a_5978_9158# rowoff_n[7] 0.10fF
C7593 a_23958_15182# a_24050_15182# 0.26fF
C7594 a_6982_15182# a_6982_14178# 1.00fF
C7595 a_2346_4180# col[14] 0.15fF
C7596 a_2346_17232# col[16] 0.15fF
C7597 a_9994_15182# rowoff_n[13] 0.10fF
C7598 a_34394_15222# vcm 0.22fF
C7599 m2_17796_18014# m3_17928_18146# 2.78fF
C7600 a_4974_7150# VDD 0.52fF
C7601 a_16018_7150# rowoff_n[5] 0.10fF
C7602 a_1962_6186# col_n[30] 0.13fF
C7603 a_2346_7192# a_21950_7150# 0.35fF
C7604 a_9994_6146# col[7] 0.29fF
C7605 a_1962_13214# col[23] 0.11fF
C7606 a_26058_5142# rowoff_n[3] 0.10fF
C7607 a_15014_18194# vcm 0.12fF
C7608 a_1962_4178# a_16018_4138# 0.27fF
C7609 a_27062_15182# col_n[24] 0.28fF
C7610 a_18026_11166# VDD 0.52fF
C7611 m3_3872_1078# m3_4876_1078# 0.22fF
C7612 a_28066_2130# col[25] 0.29fF
C7613 a_18026_9158# a_19030_9158# 0.97fF
C7614 a_2346_9200# a_35002_9158# 0.35fF
C7615 a_25054_3134# vcm 0.62fF
C7616 a_8290_12210# vcm 0.22fF
C7617 m2_21812_946# col_n[19] 0.37fF
C7618 a_24050_6146# m2_24248_6394# 0.16fF
C7619 a_1962_1166# a_9294_1166# 0.14fF
C7620 a_13006_13174# row_n[11] 0.17fF
C7621 a_1962_6186# a_29070_6146# 0.27fF
C7622 a_31078_15182# VDD 0.52fF
C7623 m2_15788_946# a_2346_1168# 0.19fF
C7624 a_28066_3134# row_n[1] 0.17fF
C7625 a_20034_17190# m3_19936_18146# 0.15fF
C7626 a_2346_13216# col[7] 0.15fF
C7627 a_21342_16226# vcm 0.22fF
C7628 a_9994_8154# col_n[7] 0.28fF
C7629 a_1962_3174# a_22346_3174# 0.14fF
C7630 a_2346_3176# a_24050_3134# 0.19fF
C7631 a_30074_4138# a_30074_3134# 1.00fF
C7632 a_1962_2170# col_n[21] 0.13fF
C7633 a_2346_1168# m2_32856_946# 0.18fF
C7634 a_1962_15222# col_n[23] 0.13fF
C7635 a_10906_18194# VDD 0.34fF
C7636 a_31078_13174# a_32082_13174# 0.97fF
C7637 a_31382_1166# vcm 0.23fF
C7638 a_28066_4138# col_n[25] 0.28fF
C7639 a_24962_11166# rowoff_n[9] 0.24fF
C7640 a_1962_9198# col[14] 0.11fF
C7641 a_32082_16186# row_n[14] 0.17fF
C7642 a_20946_3134# VDD 0.23fF
C7643 m3_24956_18146# ctop 0.23fF
C7644 a_19942_5142# a_20034_5142# 0.26fF
C7645 a_16018_14178# ctop 3.58fF
C7646 m2_23820_946# m2_24824_946# 0.96fF
C7647 col_n[17] row_n[11] 0.23fF
C7648 col_n[5] row_n[5] 0.23fF
C7649 col_n[21] row_n[13] 0.23fF
C7650 col_n[25] row_n[15] 0.23fF
C7651 VDD rowon_n[0] 2.64fF
C7652 col_n[23] row_n[14] 0.23fF
C7653 col_n[0] row_n[2] 0.23fF
C7654 col_n[3] row_n[4] 0.23fF
C7655 col_n[13] row_n[9] 0.23fF
C7656 col_n[19] row_n[12] 0.23fF
C7657 vcm rowon_n[2] 0.50fF
C7658 col_n[1] row_n[3] 0.23fF
C7659 col_n[15] row_n[10] 0.23fF
C7660 col_n[11] row_n[8] 0.23fF
C7661 col_n[7] row_n[6] 0.23fF
C7662 col_n[9] row_n[7] 0.23fF
C7663 a_35002_9158# rowoff_n[7] 0.24fF
C7664 a_2346_14220# a_6890_14178# 0.35fF
C7665 a_3970_14178# a_4974_14178# 0.97fF
C7666 a_2346_18236# a_15926_18194# 0.35fF
C7667 a_21038_7150# m2_21236_7398# 0.16fF
C7668 a_33998_7150# VDD 0.23fF
C7669 a_20034_14178# rowon_n[12] 0.14fF
C7670 a_2346_16228# a_19942_16186# 0.35fF
C7671 a_7986_11166# col[5] 0.29fF
C7672 a_9994_17190# vcm 0.60fF
C7673 a_1962_18234# m2_2736_18014# 0.18fF
C7674 a_1962_11206# col_n[14] 0.13fF
C7675 a_13006_10162# VDD 0.52fF
C7676 a_16018_9158# a_16018_8154# 1.00fF
C7677 a_32994_9158# a_33086_9158# 0.26fF
C7678 a_20034_2130# vcm 0.62fF
C7679 a_1962_13214# a_14010_13174# 0.27fF
C7680 a_26058_7150# col[23] 0.29fF
C7681 a_1962_5182# col[5] 0.11fF
C7682 a_3270_11206# vcm 0.22fF
C7683 a_12002_12170# rowoff_n[10] 0.10fF
C7684 a_13006_4138# row_n[2] 0.17fF
C7685 m3_34996_3086# VDD 0.26fF
C7686 a_2966_15182# ctop 3.42fF
C7687 a_26058_14178# VDD 0.52fF
C7688 a_2346_10204# a_8990_10162# 0.19fF
C7689 a_1962_10202# a_7286_10202# 0.14fF
C7690 a_2346_4180# col[25] 0.15fF
C7691 a_5886_10162# a_5978_10162# 0.26fF
C7692 a_2346_17232# col[27] 0.15fF
C7693 a_8990_2130# rowoff_n[0] 0.10fF
C7694 a_33086_6146# vcm 0.62fF
C7695 a_1962_15222# a_27062_15182# 0.27fF
C7696 m2_24824_18014# ctop 0.18fF
C7697 a_26058_16186# rowoff_n[14] 0.10fF
C7698 a_16322_15222# vcm 0.22fF
C7699 a_18026_8154# m2_18224_8402# 0.16fF
C7700 a_27062_3134# a_28066_3134# 0.97fF
C7701 a_31990_1126# m2_31852_946# 0.16fF
C7702 a_17022_17190# row_n[15] 0.17fF
C7703 a_2874_7150# a_2966_7150# 0.26fF
C7704 a_2346_7192# a_3878_7150# 0.35fF
C7705 a_7986_13174# col_n[5] 0.28fF
C7706 a_5886_17190# VDD 0.24fF
C7707 sample_n rowoff_n[13] 0.38fF
C7708 m2_1732_16006# vcm 0.45fF
C7709 a_2346_12212# a_22042_12170# 0.19fF
C7710 a_29070_13174# a_29070_12170# 1.00fF
C7711 a_1962_12210# a_20338_12210# 0.14fF
C7712 a_32082_7150# row_n[5] 0.17fF
C7713 m2_13780_946# m3_12908_1078# 0.13fF
C7714 col[0] rowoff_n[9] 0.11fF
C7715 ctop rowoff_n[3] 0.60fF
C7716 a_15926_2130# VDD 0.23fF
C7717 a_26058_9158# col_n[23] 0.28fF
C7718 a_1962_7190# col_n[5] 0.13fF
C7719 a_10998_13174# ctop 3.58fF
C7720 m3_34996_18146# m3_34996_17142# 0.22fF
C7721 m2_24824_946# m3_24956_1078# 2.79fF
C7722 a_1962_14218# a_33390_14218# 0.14fF
C7723 a_18938_14178# a_19030_14178# 0.26fF
C7724 a_4974_15182# rowon_n[13] 0.14fF
C7725 m2_34864_3958# VDD 1.01fF
C7726 a_28978_6146# VDD 0.23fF
C7727 a_20034_5142# rowon_n[3] 0.14fF
C7728 a_2346_6188# a_11910_6146# 0.35fF
C7729 a_24050_17190# ctop 3.39fF
C7730 a_7894_8154# rowoff_n[6] 0.24fF
C7731 a_2346_13216# col[18] 0.15fF
C7732 a_8990_2130# col_n[6] 0.28fF
C7733 a_34090_2130# ctop 3.35fF
C7734 a_4974_16186# vcm 0.62fF
C7735 a_13918_17190# rowoff_n[15] 0.24fF
C7736 a_17934_6146# rowoff_n[4] 0.24fF
C7737 a_1962_3174# a_5978_3134# 0.27fF
C7738 a_15014_9158# m2_15212_9406# 0.16fF
C7739 a_7986_9158# VDD 0.52fF
C7740 a_5978_16186# col[3] 0.29fF
C7741 a_13006_8154# a_14010_8154# 0.97fF
C7742 a_2346_8196# a_24962_8154# 0.35fF
C7743 a_15014_1126# vcm 0.12fF
C7744 a_1962_9198# col[25] 0.11fF
C7745 a_27974_4138# rowoff_n[2] 0.24fF
C7746 a_24050_12170# col[21] 0.29fF
C7747 a_1962_3174# VDD 2.73fF
C7748 col_n[6] row_n[0] 0.23fF
C7749 col_n[24] row_n[9] 0.23fF
C7750 col_n[8] row_n[1] 0.23fF
C7751 col_n[16] row_n[5] 0.23fF
C7752 a_1962_5182# a_19030_5142# 0.27fF
C7753 col_n[14] row_n[4] 0.23fF
C7754 col_n[10] row_n[2] 0.23fF
C7755 col_n[18] row_n[6] 0.23fF
C7756 a_1962_16226# sample 0.14fF
C7757 col_n[3] ctop 2.02fF
C7758 VDD col[1] 4.25fF
C7759 col_n[30] row_n[12] 0.23fF
C7760 col_n[22] row_n[8] 0.23fF
C7761 col_n[20] row_n[7] 0.23fF
C7762 rowon_n[14] row_n[14] 19.75fF
C7763 col_n[12] row_n[3] 0.23fF
C7764 col_n[28] row_n[11] 0.23fF
C7765 col_n[26] row_n[10] 0.23fF
C7766 m2_2736_18014# col[0] 0.28fF
C7767 a_21038_13174# VDD 0.52fF
C7768 a_2966_10162# a_2966_9158# 1.00fF
C7769 rowon_n[11] rowoff_n[11] 20.27fF
C7770 a_28066_5142# vcm 0.62fF
C7771 a_17022_8154# row_n[6] 0.17fF
C7772 a_11302_14218# vcm 0.22fF
C7773 a_1962_2170# a_12306_2170# 0.14fF
C7774 a_2346_2172# a_14010_2130# 0.19fF
C7775 a_25054_3134# a_25054_2130# 1.00fF
C7776 m2_31852_18014# m3_32988_18146# 0.13fF
C7777 a_1962_7190# a_32082_7150# 0.27fF
C7778 a_34090_17190# VDD 0.58fF
C7779 a_2346_9200# col[9] 0.15fF
C7780 a_26058_12170# a_27062_12170# 0.97fF
C7781 a_1962_18234# col_n[8] 0.13fF
C7782 a_6982_5142# col[4] 0.29fF
C7783 a_1962_11206# col_n[25] 0.13fF
C7784 a_24354_18234# vcm 0.22fF
C7785 a_10906_1126# VDD 0.44fF
C7786 a_1962_4178# a_25358_4178# 0.14fF
C7787 a_12002_10162# m2_12200_10410# 0.16fF
C7788 a_14922_4138# a_15014_4138# 0.26fF
C7789 a_2346_4180# a_27062_4138# 0.19fF
C7790 m2_1732_13998# rowon_n[12] 0.11fF
C7791 a_5978_12170# ctop 3.58fF
C7792 a_8990_17190# m2_8760_18014# 1.00fF
C7793 a_4974_6146# rowon_n[4] 0.14fF
C7794 a_24050_14178# col_n[21] 0.28fF
C7795 a_1962_5182# col[16] 0.11fF
C7796 m2_14784_946# VDD 0.62fF
C7797 a_35398_3174# vcm 0.23fF
C7798 a_26058_10162# rowoff_n[8] 0.10fF
C7799 m2_18800_18014# col_n[16] 0.25fF
C7800 a_28066_13174# rowoff_n[11] 0.10fF
C7801 a_23958_5142# VDD 0.23fF
C7802 m2_31852_946# VDD 0.62fF
C7803 a_19030_16186# ctop 3.57fF
C7804 m2_33860_946# analog_in 0.72fF
C7805 a_2346_15224# a_9902_15182# 0.35fF
C7806 a_24050_9158# rowon_n[7] 0.14fF
C7807 a_2874_8154# VDD 0.24fF
C7808 a_6982_7150# col_n[4] 0.28fF
C7809 a_10998_8154# a_10998_7150# 1.00fF
C7810 a_27974_8154# a_28066_8154# 0.26fF
C7811 a_2346_5184# col[0] 0.15fF
C7812 col[6] rowoff_n[4] 0.11fF
C7813 col[5] rowoff_n[3] 0.11fF
C7814 col[2] rowoff_n[0] 0.11fF
C7815 col[11] rowoff_n[9] 0.11fF
C7816 col[4] rowoff_n[2] 0.11fF
C7817 col[3] rowoff_n[1] 0.11fF
C7818 col[8] rowoff_n[6] 0.11fF
C7819 col[7] rowoff_n[5] 0.11fF
C7820 col[10] rowoff_n[8] 0.11fF
C7821 col[9] rowoff_n[7] 0.11fF
C7822 a_1962_18234# a_27366_18234# 0.14fF
C7823 a_1962_12210# a_3970_12170# 0.27fF
C7824 m2_8760_946# col_n[6] 0.37fF
C7825 a_2346_17232# a_22954_17190# 0.35fF
C7826 a_12002_17190# a_13006_17190# 0.97fF
C7827 a_1962_7190# col_n[16] 0.13fF
C7828 m2_29844_18014# m2_30848_18014# 0.96fF
C7829 a_25054_3134# col_n[22] 0.28fF
C7830 m3_34996_2082# ctop 0.23fF
C7831 a_8990_11166# m2_9188_11414# 0.16fF
C7832 a_2346_11208# m2_34864_10986# 0.17fF
C7833 a_16018_12170# VDD 0.52fF
C7834 a_1962_1166# col[7] 0.11fF
C7835 a_22042_17190# col[19] 0.29fF
C7836 a_1962_14218# col[9] 0.11fF
C7837 a_23046_4138# vcm 0.62fF
C7838 a_1962_14218# a_17022_14178# 0.27fF
C7839 a_6282_13214# vcm 0.22fF
C7840 a_15926_14178# rowoff_n[12] 0.24fF
C7841 a_22042_2130# a_23046_2130# 0.97fF
C7842 a_2346_13216# col[29] 0.15fF
C7843 a_29070_16186# VDD 0.52fF
C7844 a_24050_12170# a_24050_11166# 1.00fF
C7845 a_1962_11206# a_10298_11206# 0.14fF
C7846 a_2346_11208# a_12002_11166# 0.19fF
C7847 a_2346_7192# vcm 0.40fF
C7848 a_1962_16226# a_30074_16186# 0.27fF
C7849 a_16018_2130# m2_16216_2378# 0.16fF
C7850 a_7986_2130# m2_7756_946# 0.99fF
C7851 a_21038_12170# row_n[10] 0.17fF
C7852 a_19334_17230# vcm 0.22fF
C7853 a_4974_10162# col[2] 0.29fF
C7854 a_28066_17190# m2_27836_18014# 1.00fF
C7855 a_2346_13216# a_25054_13174# 0.19fF
C7856 a_13918_13174# a_14010_13174# 0.26fF
C7857 a_29374_2170# vcm 0.22fF
C7858 a_1962_13214# a_23350_13214# 0.14fF
C7859 a_1962_3174# col_n[7] 0.13fF
C7860 col_n[29] row_n[6] 0.23fF
C7861 VDD col[12] 4.17fF
C7862 col_n[4] col[4] 0.72fF
C7863 vcm col[8] 5.84fF
C7864 col_n[25] row_n[4] 0.23fF
C7865 a_1962_16226# col_n[9] 0.13fF
C7866 col_n[27] row_n[5] 0.23fF
C7867 col_n[14] ctop 2.02fF
C7868 col_n[23] row_n[3] 0.23fF
C7869 col_n[31] row_n[7] 0.23fF
C7870 col_n[21] row_n[2] 0.23fF
C7871 col_n[19] row_n[1] 0.23fF
C7872 col_n[17] row_n[0] 0.22fF
C7873 a_23046_6146# col[20] 0.29fF
C7874 a_18938_4138# VDD 0.23fF
C7875 a_5978_12170# m2_6176_12418# 0.16fF
C7876 a_14010_15182# ctop 3.58fF
C7877 a_2966_13174# VDD 0.56fF
C7878 a_8990_10162# rowon_n[8] 0.14fF
C7879 a_1962_10202# col[0] 0.11fF
C7880 a_2874_15182# rowoff_n[13] 0.24fF
C7881 m2_8760_18014# m3_7888_18146# 0.13fF
C7882 a_19030_1126# m3_19936_1078# 0.10fF
C7883 a_2346_9200# col[20] 0.15fF
C7884 a_31990_8154# VDD 0.23fF
C7885 a_8990_7150# rowoff_n[5] 0.10fF
C7886 a_2346_7192# a_14922_7150# 0.35fF
C7887 a_7986_7150# a_8990_7150# 0.97fF
C7888 a_1962_18234# col_n[19] 0.13fF
C7889 a_4974_12170# col_n[2] 0.28fF
C7890 a_9994_17190# a_9994_16186# 1.00fF
C7891 a_26970_17190# a_27062_17190# 0.26fF
C7892 a_19030_5142# rowoff_n[3] 0.10fF
C7893 a_7986_18194# vcm 0.12fF
C7894 a_1962_4178# a_8990_4138# 0.27fF
C7895 a_28066_13174# rowon_n[11] 0.14fF
C7896 a_1962_5182# col[27] 0.11fF
C7897 a_10998_11166# VDD 0.52fF
C7898 a_2346_9200# a_27974_9158# 0.35fF
C7899 a_23046_8154# col_n[20] 0.28fF
C7900 a_18026_3134# vcm 0.62fF
C7901 a_29070_3134# rowoff_n[1] 0.10fF
C7902 a_1962_12210# vcm 6.95fF
C7903 a_2346_1168# a_3970_1126# 0.19fF
C7904 a_20034_2130# a_20034_1126# 1.00fF
C7905 a_5978_13174# row_n[11] 0.17fF
C7906 a_1962_6186# a_22042_6146# 0.27fF
C7907 a_24050_15182# VDD 0.52fF
C7908 a_21038_11166# a_22042_11166# 0.97fF
C7909 a_21038_3134# row_n[1] 0.17fF
C7910 a_31078_7150# vcm 0.62fF
C7911 a_2346_1168# m2_8760_946# 0.19fF
C7912 a_4882_1126# m2_4744_946# 0.16fF
C7913 a_14314_16226# vcm 0.22fF
C7914 a_9902_3134# a_9994_3134# 0.26fF
C7915 a_2346_5184# col[11] 0.15fF
C7916 a_2346_3176# a_17022_3134# 0.19fF
C7917 a_1962_3174# a_15318_3174# 0.14fF
C7918 a_8990_2130# m3_8892_1078# 0.15fF
C7919 col[22] rowoff_n[9] 0.11fF
C7920 col[21] rowoff_n[8] 0.11fF
C7921 col[13] rowoff_n[0] 0.11fF
C7922 col[16] rowoff_n[3] 0.11fF
C7923 col[14] rowoff_n[1] 0.11fF
C7924 col[18] rowoff_n[5] 0.11fF
C7925 col[17] rowoff_n[4] 0.11fF
C7926 col[15] rowoff_n[2] 0.11fF
C7927 col[19] rowoff_n[6] 0.11fF
C7928 col[20] rowoff_n[7] 0.11fF
C7929 a_24354_1166# vcm 0.23fF
C7930 a_1962_7190# col_n[27] 0.13fF
C7931 m2_6752_946# m2_7756_946# 0.96fF
C7932 a_2966_17190# a_3970_17190# 0.97fF
C7933 a_17934_11166# rowoff_n[9] 0.24fF
C7934 a_25054_16186# row_n[14] 0.17fF
C7935 a_13918_3134# VDD 0.23fF
C7936 a_1962_5182# a_28370_5182# 0.14fF
C7937 a_1962_1166# col[18] 0.11fF
C7938 a_2346_5184# a_30074_5142# 0.19fF
C7939 a_33086_6146# a_33086_5142# 1.00fF
C7940 a_8990_14178# ctop 3.58fF
C7941 a_1962_14218# col[20] 0.11fF
C7942 a_21038_11166# col[18] 0.29fF
C7943 a_27974_9158# rowoff_n[7] 0.24fF
C7944 a_2346_18236# a_8898_18194# 0.35fF
C7945 a_31990_15182# rowoff_n[13] 0.24fF
C7946 m2_1732_6970# VDD 1.02fF
C7947 col[6] rowoff_n[10] 0.11fF
C7948 a_26970_7150# VDD 0.23fF
C7949 a_34090_15182# m2_34288_15430# 0.16fF
C7950 a_5978_7150# a_5978_6146# 1.00fF
C7951 a_22954_7150# a_23046_7150# 0.26fF
C7952 a_13006_14178# rowon_n[12] 0.14fF
C7953 a_2346_16228# a_12914_16186# 0.35fF
C7954 a_6982_16186# a_7986_16186# 0.97fF
C7955 a_2966_12170# row_n[10] 0.16fF
C7956 a_28066_4138# rowon_n[2] 0.14fF
C7957 a_32082_3134# ctop 3.57fF
C7958 a_2346_1168# col[2] 0.14fF
C7959 a_2346_14220# col[4] 0.15fF
C7960 a_3970_4138# col[1] 0.29fF
C7961 a_5978_10162# VDD 0.52fF
C7962 a_1962_3174# col_n[18] 0.13fF
C7963 a_13006_2130# vcm 0.62fF
C7964 a_1962_13214# a_6982_13174# 0.27fF
C7965 col_n[28] row_n[0] 0.23fF
C7966 col_n[25] ctop 2.02fF
C7967 VDD col[23] 4.17fF
C7968 vcm col[19] 5.84fF
C7969 col_n[9] col[10] 5.98fF
C7970 col_n[30] row_n[1] 0.23fF
C7971 a_1962_16226# col_n[20] 0.13fF
C7972 a_21038_13174# col_n[18] 0.28fF
C7973 a_4974_12170# rowoff_n[10] 0.10fF
C7974 a_5978_4138# row_n[2] 0.17fF
C7975 a_2346_1168# a_32994_1126# 0.35fF
C7976 m3_34996_17142# VDD 0.27fF
C7977 a_1962_10202# col[11] 0.11fF
C7978 a_32082_17190# rowon_n[15] 0.14fF
C7979 a_19030_14178# VDD 0.52fF
C7980 a_19030_11166# a_19030_10162# 1.00fF
C7981 m2_33860_18014# col[31] 0.28fF
C7982 a_1962_15222# a_20034_15182# 0.27fF
C7983 a_26058_6146# vcm 0.62fF
C7984 m2_1732_9982# m2_2160_10410# 0.16fF
C7985 a_2346_9200# col[31] 0.15fF
C7986 m2_10768_18014# ctop 0.18fF
C7987 a_19030_16186# rowoff_n[14] 0.10fF
C7988 a_9294_15222# vcm 0.22fF
C7989 a_9994_17190# row_n[15] 0.17fF
C7990 a_1962_18234# col_n[30] 0.13fF
C7991 a_31078_16186# m2_31276_16434# 0.16fF
C7992 m2_1732_2954# row_n[1] 0.13fF
C7993 a_8898_12170# a_8990_12170# 0.26fF
C7994 a_2346_12212# a_15014_12170# 0.19fF
C7995 a_1962_12210# a_13310_12210# 0.14fF
C7996 a_25054_7150# row_n[5] 0.17fF
C7997 a_3970_6146# col_n[1] 0.28fF
C7998 a_1962_17230# a_33086_17190# 0.27fF
C7999 a_33086_4138# m2_33284_4386# 0.16fF
C8000 m2_8760_946# m3_8892_1078# 2.79fF
C8001 a_8898_2130# VDD 0.23fF
C8002 a_30074_5142# a_31078_5142# 0.97fF
C8003 a_3970_13174# ctop 3.57fF
C8004 a_7894_18194# m2_7756_18014# 0.16fF
C8005 a_22042_2130# col_n[19] 0.28fF
C8006 a_1962_12210# col_n[11] 0.13fF
C8007 a_32386_4178# vcm 0.22fF
C8008 a_2346_14220# a_28066_14178# 0.19fF
C8009 a_1962_14218# a_26362_14218# 0.14fF
C8010 a_32082_15182# a_32082_14178# 1.00fF
C8011 a_19030_16186# col[16] 0.29fF
C8012 a_21950_6146# VDD 0.23fF
C8013 a_1962_6186# col[2] 0.11fF
C8014 a_13006_5142# rowon_n[3] 0.14fF
C8015 a_2346_6188# a_4882_6146# 0.35fF
C8016 a_17022_17190# ctop 3.39fF
C8017 a_2966_3134# row_n[1] 0.16fF
C8018 a_4974_16186# a_4974_15182# 1.00fF
C8019 a_21950_16186# a_22042_16186# 0.26fF
C8020 a_2346_5184# col[22] 0.15fF
C8021 m2_34864_13998# m2_34864_12994# 0.99fF
C8022 a_6890_17190# rowoff_n[15] 0.24fF
C8023 a_27062_2130# ctop 3.39fF
C8024 col[24] rowoff_n[0] 0.11fF
C8025 col[26] rowoff_n[2] 0.11fF
C8026 col[25] rowoff_n[1] 0.11fF
C8027 col[31] rowoff_n[7] 0.11fF
C8028 m2_30848_18014# VDD 1.33fF
C8029 col[28] rowoff_n[4] 0.11fF
C8030 col[27] rowoff_n[3] 0.11fF
C8031 col[30] rowoff_n[6] 0.11fF
C8032 col[29] rowoff_n[5] 0.11fF
C8033 a_10906_6146# rowoff_n[4] 0.24fF
C8034 a_35002_10162# VDD 0.29fF
C8035 a_28066_17190# m2_28264_17438# 0.16fF
C8036 a_2346_8196# a_17934_8154# 0.35fF
C8037 a_1962_13214# a_34394_13214# 0.14fF
C8038 a_7986_1126# vcm 0.12fF
C8039 a_20946_4138# rowoff_n[2] 0.24fF
C8040 a_33998_12170# rowoff_n[10] 0.24fF
C8041 a_1962_1166# col[29] 0.11fF
C8042 a_32082_8154# rowon_n[6] 0.14fF
C8043 a_30074_5142# m2_30272_5390# 0.16fF
C8044 a_1962_14218# col[31] 0.11fF
C8045 a_1962_5182# a_12002_5142# 0.27fF
C8046 a_14010_13174# VDD 0.52fF
C8047 a_20034_5142# col[17] 0.29fF
C8048 a_16018_10162# a_17022_10162# 0.97fF
C8049 a_2346_10204# a_30986_10162# 0.35fF
C8050 a_30986_2130# rowoff_n[0] 0.24fF
C8051 a_1962_8194# col_n[2] 0.13fF
C8052 a_21038_5142# vcm 0.62fF
C8053 m2_26832_946# vcm 0.42fF
C8054 col[17] rowoff_n[10] 0.11fF
C8055 a_9994_8154# row_n[6] 0.17fF
C8056 a_4274_14218# vcm 0.22fF
C8057 a_4882_2130# a_4974_2130# 0.26fF
C8058 a_1962_2170# a_5278_2170# 0.14fF
C8059 a_2346_2172# a_6982_2130# 0.19fF
C8060 m2_22816_18014# m3_22948_18146# 2.78fF
C8061 a_1962_7190# a_25054_7150# 0.27fF
C8062 a_27062_17190# VDD 0.55fF
C8063 a_34090_9158# vcm 0.62fF
C8064 a_2346_1168# col[13] 0.14fF
C8065 a_2346_14220# col[15] 0.15fF
C8066 a_17326_18234# vcm 0.22fF
C8067 a_2346_4180# a_20034_4138# 0.19fF
C8068 a_1962_4178# a_18330_4178# 0.14fF
C8069 a_28066_5142# a_28066_4138# 1.00fF
C8070 a_1962_3174# col_n[29] 0.13fF
C8071 rowon_n[6] rowon_n[5] 0.15fF
C8072 vcm col[30] 5.84fF
C8073 col_n[31] analog_in 0.13fF
C8074 rowon_n[13] ctop 1.40fF
C8075 col_n[15] col[15] 0.64fF
C8076 a_1962_16226# col_n[31] 0.13fF
C8077 a_26970_18194# m2_26832_18014# 0.16fF
C8078 a_29070_11166# row_n[9] 0.17fF
C8079 a_29070_14178# a_30074_14178# 0.97fF
C8080 a_27366_3174# vcm 0.22fF
C8081 a_19030_10162# rowoff_n[8] 0.10fF
C8082 col[1] rowoff_n[11] 0.11fF
C8083 a_20034_7150# col_n[17] 0.28fF
C8084 a_21038_13174# rowoff_n[11] 0.10fF
C8085 m2_7756_946# VDD 0.62fF
C8086 a_1962_10202# col[22] 0.11fF
C8087 a_27062_6146# m2_27260_6394# 0.16fF
C8088 a_16930_5142# VDD 0.23fF
C8089 a_2346_6188# a_33086_6146# 0.19fF
C8090 a_1962_6186# a_31382_6186# 0.14fF
C8091 a_17934_6146# a_18026_6146# 0.26fF
C8092 a_12002_16186# ctop 3.57fF
C8093 a_29070_8154# rowoff_n[6] 0.10fF
C8094 a_23046_17190# m3_22948_18146# 0.15fF
C8095 m2_22816_946# m3_21944_1078# 0.13fF
C8096 a_17022_9158# rowon_n[7] 0.14fF
C8097 a_29982_9158# VDD 0.23fF
C8098 a_1962_18234# a_20338_18234# 0.14fF
C8099 a_2346_17232# a_15926_17190# 0.35fF
C8100 a_2346_10204# col[6] 0.15fF
C8101 m2_22816_18014# m2_23820_18014# 0.96fF
C8102 m3_1864_15134# ctop 0.23fF
C8103 a_2966_5142# m3_1864_5094# 0.14fF
C8104 a_1962_12210# col_n[22] 0.13fF
C8105 a_8990_12170# VDD 0.52fF
C8106 m2_27836_946# m2_28264_1374# 0.16fF
C8107 m2_31852_946# col_n[29] 0.42fF
C8108 a_14010_10162# a_14010_9158# 1.00fF
C8109 a_30986_10162# a_31078_10162# 0.26fF
C8110 a_16018_4138# vcm 0.62fF
C8111 a_1962_14218# a_9994_14178# 0.27fF
C8112 a_18026_10162# col[15] 0.29fF
C8113 m2_34864_12994# ctop 0.17fF
C8114 a_8898_14178# rowoff_n[12] 0.24fF
C8115 a_1962_6186# col[13] 0.11fF
C8116 a_24050_7150# m2_24248_7398# 0.16fF
C8117 m2_34864_16006# m3_34996_15134# 0.15fF
C8118 a_3878_6146# VDD 0.23fF
C8119 a_2966_3134# col[0] 0.29fF
C8120 a_22042_16186# VDD 0.52fF
C8121 a_2346_11208# a_4974_11166# 0.19fF
C8122 a_1962_11206# a_3270_11206# 0.14fF
C8123 a_29070_8154# vcm 0.62fF
C8124 a_1962_16226# a_23046_16186# 0.27fF
C8125 a_14010_12170# row_n[10] 0.17fF
C8126 a_12306_17230# vcm 0.22fF
C8127 a_25054_4138# a_26058_4138# 0.97fF
C8128 a_29070_2130# row_n[0] 0.17fF
C8129 a_22346_2170# vcm 0.22fF
C8130 a_1962_13214# a_16322_13214# 0.14fF
C8131 a_27062_14178# a_27062_13174# 1.00fF
C8132 a_2346_13216# a_18026_13174# 0.19fF
C8133 a_18026_12170# col_n[15] 0.28fF
C8134 a_11910_4138# VDD 0.23fF
C8135 m3_12908_1078# VDD 0.14fF
C8136 a_1962_8194# col_n[13] 0.13fF
C8137 a_6982_15182# ctop 3.58fF
C8138 col[28] rowoff_n[10] 0.11fF
C8139 a_33086_15182# row_n[13] 0.17fF
C8140 a_1962_15222# a_29374_15222# 0.14fF
C8141 a_16930_15182# a_17022_15182# 0.26fF
C8142 a_2966_5142# vcm 0.61fF
C8143 a_2346_15224# a_31078_15182# 0.19fF
C8144 a_1962_2170# col[4] 0.11fF
C8145 a_1962_15222# col[6] 0.11fF
C8146 a_21038_8154# m2_21236_8402# 0.16fF
C8147 a_24962_8154# VDD 0.23fF
C8148 a_2346_7192# a_7894_7150# 0.35fF
C8149 a_2346_1168# col[24] 0.14fF
C8150 a_2346_14220# col[26] 0.15fF
C8151 a_12002_5142# rowoff_n[3] 0.10fF
C8152 a_30074_4138# ctop 3.58fF
C8153 row_n[8] ctop 1.65fF
C8154 col_n[20] col[21] 5.98fF
C8155 rowon_n[3] row_n[3] 19.75fF
C8156 a_21038_13174# rowon_n[11] 0.14fF
C8157 a_3970_11166# VDD 0.52fF
C8158 m2_29844_946# m3_29976_1078# 2.79fF
C8159 a_10998_9158# a_12002_9158# 0.97fF
C8160 a_2346_9200# a_20946_9158# 0.35fF
C8161 col[12] rowoff_n[11] 0.11fF
C8162 a_10998_3134# vcm 0.62fF
C8163 a_22042_3134# rowoff_n[1] 0.10fF
C8164 a_19030_1126# col_n[16] 0.31fF
C8165 a_2966_13174# rowoff_n[11] 0.10fF
C8166 m2_34864_12994# m3_34996_12122# 0.15fF
C8167 a_16018_15182# col[13] 0.29fF
C8168 a_1962_4178# col_n[4] 0.13fF
C8169 a_1962_6186# a_15014_6146# 0.27fF
C8170 a_1962_17230# col_n[6] 0.13fF
C8171 a_17022_15182# VDD 0.52fF
C8172 a_2346_11208# a_33998_11166# 0.35fF
C8173 a_14010_3134# row_n[1] 0.17fF
C8174 a_24050_7150# vcm 0.62fF
C8175 a_34090_11166# col[31] 0.29fF
C8176 a_7286_16226# vcm 0.22fF
C8177 a_23046_4138# a_23046_3134# 1.00fF
C8178 a_1962_3174# a_8290_3174# 0.14fF
C8179 a_18026_9158# m2_18224_9406# 0.16fF
C8180 a_2346_3176# a_9994_3134# 0.19fF
C8181 a_1962_8194# a_28066_8154# 0.27fF
C8182 a_2346_10204# col[17] 0.15fF
C8183 a_17326_1166# vcm 0.23fF
C8184 a_24050_13174# a_25054_13174# 0.97fF
C8185 a_10906_11166# rowoff_n[9] 0.24fF
C8186 a_18026_16186# row_n[14] 0.17fF
C8187 a_6890_3134# VDD 0.23fF
C8188 a_1962_5182# a_21342_5182# 0.14fF
C8189 a_12914_5142# a_13006_5142# 0.26fF
C8190 a_2346_5184# a_23046_5142# 0.19fF
C8191 a_33086_6146# row_n[4] 0.17fF
C8192 a_16018_17190# col_n[13] 0.28fF
C8193 a_20946_9158# rowoff_n[7] 0.24fF
C8194 a_1962_6186# col[24] 0.11fF
C8195 a_30378_5182# vcm 0.22fF
C8196 a_17022_4138# col[14] 0.29fF
C8197 a_24962_15182# rowoff_n[13] 0.24fF
C8198 m2_1732_4962# rowon_n[3] 0.11fF
C8199 a_19942_7150# VDD 0.23fF
C8200 a_30986_7150# rowoff_n[5] 0.24fF
C8201 a_34090_13174# col_n[31] 0.28fF
C8202 a_2346_7192# a_2346_6188# 0.22fF
C8203 a_1962_7190# a_35398_7190# 0.14fF
C8204 a_5978_14178# rowon_n[12] 0.14fF
C8205 a_2346_16228# a_5886_16186# 0.35fF
C8206 a_21038_4138# rowon_n[2] 0.14fF
C8207 a_25054_3134# ctop 3.57fF
C8208 a_15014_10162# m2_15212_10410# 0.16fF
C8209 a_32994_11166# VDD 0.23fF
C8210 m3_32988_1078# m3_33992_1078# 0.21fF
C8211 a_8990_9158# a_8990_8154# 1.00fF
C8212 a_25966_9158# a_26058_9158# 0.26fF
C8213 a_2346_6188# col[8] 0.15fF
C8214 a_5978_2130# vcm 0.62fF
C8215 a_2346_1168# a_25966_1126# 0.35fF
C8216 a_1962_8194# col_n[24] 0.13fF
C8217 a_17022_6146# col_n[14] 0.28fF
C8218 m2_34864_9982# m3_34996_9110# 0.15fF
C8219 m3_8892_18146# VDD 0.24fF
C8220 a_25054_17190# rowon_n[15] 0.14fF
C8221 a_12002_14178# VDD 0.52fF
C8222 m2_16792_946# a_16930_1126# 0.16fF
C8223 a_1962_2170# col[15] 0.11fF
C8224 a_1962_15222# col[17] 0.11fF
C8225 a_19030_6146# vcm 0.62fF
C8226 a_1962_15222# a_13006_15182# 0.27fF
C8227 a_12002_16186# rowoff_n[14] 0.10fF
C8228 a_20034_3134# a_21038_3134# 0.97fF
C8229 a_32082_16186# col[29] 0.29fF
C8230 m2_25828_18014# vcm 0.28fF
C8231 a_2346_12212# a_7986_12170# 0.19fF
C8232 a_22042_13174# a_22042_12170# 1.00fF
C8233 a_1962_12210# a_6282_12210# 0.14fF
C8234 a_2346_18236# col[9] 0.14fF
C8235 a_18026_7150# row_n[5] 0.17fF
C8236 a_1962_17230# a_26058_17190# 0.27fF
C8237 a_32082_10162# vcm 0.62fF
C8238 col_n[26] col[26] 0.78fF
C8239 rowon_n[2] ctop 1.40fF
C8240 m2_33860_18014# m2_34288_18442# 0.16fF
C8241 m3_15920_1078# ctop 0.23fF
C8242 col[23] rowoff_n[11] 0.11fF
C8243 a_12002_11166# m2_12200_11414# 0.16fF
C8244 a_2966_13174# rowon_n[11] 0.13fF
C8245 a_2346_9200# a_1962_9198# 2.62fF
C8246 a_2346_15224# col[1] 0.15fF
C8247 a_2966_14178# m3_1864_14130# 0.14fF
C8248 a_2346_14220# a_21038_14178# 0.19fF
C8249 a_11910_14178# a_12002_14178# 0.26fF
C8250 a_25358_4178# vcm 0.22fF
C8251 a_1962_14218# a_19334_14218# 0.14fF
C8252 a_1962_4178# col_n[15] 0.13fF
C8253 a_1962_17230# col_n[17] 0.13fF
C8254 a_15014_9158# col[12] 0.29fF
C8255 a_14922_6146# VDD 0.23fF
C8256 a_5978_5142# rowon_n[3] 0.14fF
C8257 a_33086_7150# a_34090_7150# 0.97fF
C8258 a_9994_17190# ctop 3.39fF
C8259 m2_12776_18014# col_n[10] 0.25fF
C8260 a_1962_11206# col[8] 0.11fF
C8261 a_2346_16228# a_34090_16186# 0.19fF
C8262 a_1962_16226# a_32386_16226# 0.14fF
C8263 a_33086_5142# col[30] 0.29fF
C8264 a_19030_2130# m2_19228_2378# 0.16fF
C8265 a_20034_2130# ctop 3.43fF
C8266 m2_16792_18014# VDD 0.91fF
C8267 col[7] rowoff_n[12] 0.11fF
C8268 a_1962_18234# m2_31852_18014# 0.18fF
C8269 a_27974_10162# VDD 0.23fF
C8270 a_2346_10204# col[28] 0.15fF
C8271 a_5978_8154# a_6982_8154# 0.97fF
C8272 a_2346_8196# a_10906_8154# 0.35fF
C8273 a_13918_4138# rowoff_n[2] 0.24fF
C8274 a_26970_12170# rowoff_n[10] 0.24fF
C8275 a_25054_8154# rowon_n[6] 0.14fF
C8276 a_33086_6146# ctop 3.57fF
C8277 m2_34864_6970# m3_34996_6098# 0.15fF
C8278 a_1962_5182# a_4974_5142# 0.27fF
C8279 a_2346_12212# m2_34864_11990# 0.17fF
C8280 a_8990_12170# m2_9188_12418# 0.16fF
C8281 a_3878_5142# a_3970_5142# 0.26fF
C8282 a_6982_13174# VDD 0.52fF
C8283 a_2346_18236# m2_26832_18014# 0.19fF
C8284 a_2346_10204# a_23958_10162# 0.35fF
C8285 a_15014_11166# col_n[12] 0.28fF
C8286 a_23958_2130# rowoff_n[0] 0.24fF
C8287 a_14010_5142# vcm 0.62fF
C8288 m2_1732_16006# ctop 0.17fF
C8289 a_1962_13214# col_n[8] 0.13fF
C8290 a_18026_3134# a_18026_2130# 1.00fF
C8291 m2_13780_18014# m3_12908_18146# 0.13fF
C8292 a_35494_8516# VDD 0.11fF
C8293 a_33086_7150# col_n[30] 0.28fF
C8294 a_1962_7190# a_18026_7150# 0.27fF
C8295 a_20034_17190# VDD 0.55fF
C8296 a_1962_12210# a_1962_11206# 0.16fF
C8297 a_19030_12170# a_20034_12170# 0.97fF
C8298 a_27062_9158# vcm 0.62fF
C8299 a_2966_4138# rowon_n[2] 0.13fF
C8300 a_10298_18234# vcm 0.22fF
C8301 a_30074_2130# VDD 0.55fF
C8302 a_7894_4138# a_7986_4138# 0.26fF
C8303 a_1962_4178# a_11302_4178# 0.14fF
C8304 a_2346_4180# a_13006_4138# 0.19fF
C8305 a_2346_6188# col[19] 0.15fF
C8306 m3_1864_3086# m3_1864_2082# 0.22fF
C8307 a_1962_9198# a_31078_9158# 0.27fF
C8308 a_22042_11166# row_n[9] 0.17fF
C8309 a_20338_3174# vcm 0.22fF
C8310 a_12002_10162# rowoff_n[8] 0.10fF
C8311 a_14010_13174# rowoff_n[11] 0.10fF
C8312 a_9902_5142# VDD 0.23fF
C8313 a_5978_13174# m2_6176_13422# 0.16fF
C8314 a_1962_6186# a_24354_6186# 0.14fF
C8315 a_2346_6188# a_26058_6146# 0.19fF
C8316 a_31078_7150# a_31078_6146# 1.00fF
C8317 a_1962_2170# col[26] 0.11fF
C8318 a_4974_16186# ctop 3.57fF
C8319 a_1962_15222# col[28] 0.11fF
C8320 a_22042_8154# rowoff_n[6] 0.10fF
C8321 a_13006_14178# col[10] 0.29fF
C8322 a_32082_16186# a_33086_16186# 0.97fF
C8323 a_33390_7190# vcm 0.22fF
C8324 a_1962_9198# col_n[0] 0.13fF
C8325 a_28066_17190# rowoff_n[15] 0.10fF
C8326 a_32082_6146# rowoff_n[4] 0.10fF
C8327 a_1962_1166# m2_25828_946# 0.18fF
C8328 a_12002_2130# m3_11904_1078# 0.15fF
C8329 a_9994_9158# rowon_n[7] 0.14fF
C8330 a_22954_9158# VDD 0.23fF
C8331 a_31078_10162# col[28] 0.29fF
C8332 a_2346_18236# col[20] 0.14fF
C8333 a_20946_8154# a_21038_8154# 0.26fF
C8334 a_3970_8154# a_3970_7150# 1.00fF
C8335 sw analog_in 0.69fF
C8336 a_1962_18234# a_13310_18234# 0.14fF
C8337 m2_10768_946# m2_11196_1374# 0.16fF
C8338 a_2346_17232# a_8898_17190# 0.35fF
C8339 a_4974_17190# a_5978_17190# 0.97fF
C8340 m2_15788_18014# m2_16792_18014# 0.96fF
C8341 m2_34864_3958# m3_34996_3086# 0.15fF
C8342 a_28066_5142# ctop 3.58fF
C8343 a_2346_2172# col[10] 0.15fF
C8344 m3_11904_18146# ctop 0.23fF
C8345 a_2346_15224# col[12] 0.15fF
C8346 a_1962_4178# col_n[26] 0.13fF
C8347 a_8990_4138# vcm 0.62fF
C8348 a_2346_14220# a_2966_14178# 0.21fF
C8349 a_1962_17230# col_n[28] 0.13fF
C8350 a_13006_16186# col_n[10] 0.28fF
C8351 a_29070_12170# rowon_n[10] 0.14fF
C8352 a_15014_2130# a_16018_2130# 0.97fF
C8353 a_14010_3134# col[11] 0.29fF
C8354 a_2346_2172# a_28978_2130# 0.35fF
C8355 a_1962_18234# col[2] 0.11fF
C8356 a_1962_11206# col[19] 0.11fF
C8357 a_15014_16186# VDD 0.52fF
C8358 a_33998_12170# a_34090_12170# 0.26fF
C8359 a_17022_12170# a_17022_11166# 1.00fF
C8360 a_31078_12170# col_n[28] 0.28fF
C8361 col[18] rowoff_n[12] 0.11fF
C8362 a_22042_8154# vcm 0.62fF
C8363 a_1962_16226# a_16018_16186# 0.27fF
C8364 a_6982_12170# row_n[10] 0.17fF
C8365 a_5278_17230# vcm 0.22fF
C8366 a_22042_2130# row_n[0] 0.17fF
C8367 a_2346_13216# a_10998_13174# 0.19fF
C8368 a_15318_2170# vcm 0.22fF
C8369 a_6890_13174# a_6982_13174# 0.26fF
C8370 a_1962_13214# a_9294_13214# 0.14fF
C8371 a_35094_12170# vcm 0.12fF
C8372 a_4882_4138# VDD 0.23fF
C8373 a_2346_11208# col[3] 0.15fF
C8374 m3_1864_9110# VDD 0.25fF
C8375 a_28066_6146# a_29070_6146# 0.97fF
C8376 a_14010_5142# col_n[11] 0.28fF
C8377 col[2] rowoff_n[13] 0.11fF
C8378 a_26058_15182# row_n[13] 0.17fF
C8379 a_28370_6186# vcm 0.22fF
C8380 a_1962_13214# col_n[19] 0.13fF
C8381 a_30074_16186# a_30074_15182# 1.00fF
C8382 a_1962_15222# a_22346_15222# 0.14fF
C8383 a_2346_15224# a_24050_15182# 0.19fF
C8384 a_17934_8154# VDD 0.23fF
C8385 a_1962_7190# col[10] 0.11fF
C8386 a_34090_16186# m2_34288_16434# 0.16fF
C8387 a_29070_15182# col[26] 0.29fF
C8388 a_19942_17190# a_20034_17190# 0.26fF
C8389 m2_1732_17010# m2_1732_16006# 0.99fF
C8390 a_2346_6188# col[30] 0.15fF
C8391 a_4974_5142# rowoff_n[3] 0.10fF
C8392 a_23046_4138# ctop 3.58fF
C8393 a_14010_13174# rowon_n[11] 0.14fF
C8394 a_30986_12170# VDD 0.23fF
C8395 m3_28972_18146# m3_29976_18146# 0.22fF
C8396 a_2346_9200# a_13918_9158# 0.35fF
C8397 a_3970_3134# vcm 0.62fF
C8398 a_15014_3134# rowoff_n[1] 0.10fF
C8399 a_29070_3134# rowon_n[1] 0.14fF
C8400 a_30074_14178# rowoff_n[12] 0.10fF
C8401 a_29982_2130# a_30074_2130# 0.26fF
C8402 a_2346_7192# ctop 1.59fF
C8403 a_1962_6186# a_7986_6146# 0.27fF
C8404 a_9994_15182# VDD 0.52fF
C8405 a_12002_8154# col[9] 0.29fF
C8406 m2_1732_10986# rowoff_n[9] 0.12fF
C8407 m2_34864_8978# vcm 0.51fF
C8408 a_14010_11166# a_15014_11166# 0.97fF
C8409 a_2346_11208# a_26970_11166# 0.35fF
C8410 a_2966_17190# m3_2868_18146# 0.15fF
C8411 a_6982_3134# row_n[1] 0.17fF
C8412 a_1962_9198# col_n[10] 0.13fF
C8413 a_17022_7150# vcm 0.62fF
C8414 a_29070_17190# col_n[26] 0.28fF
C8415 a_33086_16186# rowon_n[14] 0.14fF
C8416 a_2346_18236# col[31] 0.14fF
C8417 a_2346_3176# a_2874_3134# 0.35fF
C8418 a_30074_4138# col[27] 0.29fF
C8419 a_1962_3174# col[1] 0.11fF
C8420 ctop col[8] 1.98fF
C8421 a_1962_16226# col[3] 0.11fF
C8422 m2_27836_18014# col[25] 0.28fF
C8423 a_31078_17190# m2_31276_17438# 0.16fF
C8424 a_1962_8194# a_21038_8154# 0.27fF
C8425 a_10298_1166# vcm 0.23fF
C8426 a_30074_11166# vcm 0.62fF
C8427 a_2346_2172# col[21] 0.15fF
C8428 a_10998_16186# row_n[14] 0.17fF
C8429 a_33086_5142# m2_33284_5390# 0.16fF
C8430 a_2346_15224# col[23] 0.15fF
C8431 a_33086_4138# VDD 0.52fF
C8432 a_1962_5182# a_14314_5182# 0.14fF
C8433 a_26058_6146# a_26058_5142# 1.00fF
C8434 a_2346_5184# a_16018_5142# 0.19fF
C8435 a_26058_6146# row_n[4] 0.17fF
C8436 a_1962_10202# a_34090_10162# 0.27fF
C8437 a_13918_9158# rowoff_n[7] 0.24fF
C8438 a_27062_15182# a_28066_15182# 0.97fF
C8439 a_23350_5182# vcm 0.22fF
C8440 m2_34864_946# vcm 0.48fF
C8441 a_12002_10162# col_n[9] 0.28fF
C8442 a_1962_18234# col[13] 0.11fF
C8443 a_17934_15182# rowoff_n[13] 0.24fF
C8444 a_1962_11206# col[30] 0.11fF
C8445 m2_27836_18014# m3_27968_18146# 2.78fF
C8446 a_12914_7150# VDD 0.23fF
C8447 a_23958_7150# rowoff_n[5] 0.24fF
C8448 a_1962_7190# a_27366_7190# 0.14fF
C8449 a_2346_7192# a_29070_7150# 0.19fF
C8450 a_15926_7150# a_16018_7150# 0.26fF
C8451 col[29] rowoff_n[12] 0.11fF
C8452 m2_1732_16006# rowoff_n[14] 0.12fF
C8453 a_1962_5182# col_n[1] 0.13fF
C8454 a_30074_6146# col_n[27] 0.28fF
C8455 m2_1732_10986# sample_n 0.15fF
C8456 a_33998_5142# rowoff_n[3] 0.24fF
C8457 a_14010_4138# rowon_n[2] 0.14fF
C8458 a_18026_3134# ctop 3.57fF
C8459 a_1962_12210# ctop 1.49fF
C8460 a_25966_11166# VDD 0.23fF
C8461 m3_18932_1078# m3_19936_1078# 0.13fF
C8462 m2_34864_4962# m2_35292_5390# 0.16fF
C8463 a_2346_11208# col[14] 0.15fF
C8464 a_30074_6146# m2_30272_6394# 0.16fF
C8465 a_2346_1168# a_18938_1126# 0.39fF
C8466 a_31078_7150# ctop 3.58fF
C8467 a_18026_17190# rowon_n[15] 0.14fF
C8468 a_34090_8154# m3_34996_8106# 0.13fF
C8469 col[13] rowoff_n[13] 0.11fF
C8470 a_4974_14178# VDD 0.52fF
C8471 a_1962_13214# col_n[30] 0.13fF
C8472 a_28978_11166# a_29070_11166# 0.26fF
C8473 a_12002_11166# a_12002_10162# 1.00fF
C8474 a_26058_17190# m3_25960_18146# 0.15fF
C8475 VDD rowoff_n[9] 1.17fF
C8476 a_12002_6146# vcm 0.62fF
C8477 a_33086_7150# rowon_n[5] 0.14fF
C8478 a_1962_15222# a_5978_15182# 0.27fF
C8479 a_9994_13174# col[7] 0.29fF
C8480 a_4974_16186# rowoff_n[14] 0.10fF
C8481 a_1962_7190# col[21] 0.11fF
C8482 a_2346_3176# a_31990_3134# 0.35fF
C8483 a_28066_9158# col[25] 0.29fF
C8484 m2_11772_18014# vcm 0.28fF
C8485 a_10998_7150# row_n[5] 0.17fF
C8486 a_32082_11166# rowoff_n[9] 0.10fF
C8487 a_25054_10162# vcm 0.62fF
C8488 a_1962_17230# a_19030_17190# 0.27fF
C8489 m2_26832_18014# m2_27260_18442# 0.16fF
C8490 a_28066_3134# VDD 0.52fF
C8491 m3_34996_8106# ctop 0.23fF
C8492 a_23046_5142# a_24050_5142# 0.97fF
C8493 a_18330_4178# vcm 0.22fF
C8494 a_25054_15182# a_25054_14178# 1.00fF
C8495 a_1962_14218# a_12306_14218# 0.14fF
C8496 a_2346_14220# a_14010_14178# 0.19fF
C8497 a_2346_7192# col[5] 0.15fF
C8498 a_27062_7150# m2_27260_7398# 0.16fF
C8499 a_9994_15182# col_n[7] 0.28fF
C8500 a_7894_6146# VDD 0.23fF
C8501 a_10998_2130# col[8] 0.29fF
C8502 a_1962_9198# col_n[21] 0.13fF
C8503 a_30074_10162# row_n[8] 0.17fF
C8504 a_31382_8194# vcm 0.22fF
C8505 a_1962_16226# a_25358_16226# 0.14fF
C8506 a_14922_16186# a_15014_16186# 0.26fF
C8507 a_2346_16228# a_27062_16186# 0.19fF
C8508 a_1962_3174# col[12] 0.11fF
C8509 a_28066_11166# col_n[25] 0.28fF
C8510 a_13006_2130# ctop 3.39fF
C8511 VDD sample_n 26.64fF
C8512 ctop col[19] 1.98fF
C8513 m2_2736_18014# VDD 1.27fF
C8514 en_bit_n[2] col[16] 0.16fF
C8515 col[6] col[7] 0.20fF
C8516 a_1962_16226# col[14] 0.11fF
C8517 a_1962_18234# m2_17796_18014# 0.18fF
C8518 a_20946_10162# VDD 0.23fF
C8519 a_1962_8194# a_2966_8154# 0.27fF
C8520 a_6890_4138# rowoff_n[2] 0.24fF
C8521 a_19942_12170# rowoff_n[10] 0.24fF
C8522 a_18026_8154# rowon_n[6] 0.14fF
C8523 a_26058_6146# ctop 3.58fF
C8524 m3_27968_1078# VDD 0.14fF
C8525 a_2346_18236# m2_12776_18014# 0.19fF
C8526 a_33998_14178# VDD 0.23fF
C8527 a_8990_10162# a_9994_10162# 0.97fF
C8528 a_2346_10204# a_16930_10162# 0.35fF
C8529 a_16930_2130# rowoff_n[0] 0.24fF
C8530 a_1962_18234# col[24] 0.11fF
C8531 a_6982_5142# vcm 0.62fF
C8532 a_10998_4138# col_n[8] 0.28fF
C8533 a_33998_16186# rowoff_n[14] 0.24fF
C8534 a_24050_8154# m2_24248_8402# 0.16fF
C8535 m2_25828_946# col_n[23] 0.37fF
C8536 m2_3740_18014# m3_4876_18146# 0.13fF
C8537 a_1962_7190# a_10998_7150# 0.27fF
C8538 a_1962_5182# col_n[12] 0.13fF
C8539 m2_14784_946# col[12] 0.39fF
C8540 a_13006_17190# VDD 0.55fF
C8541 a_2346_12212# a_29982_12170# 0.35fF
C8542 a_20034_9158# vcm 0.62fF
C8543 a_26058_14178# col[23] 0.29fF
C8544 a_1962_12210# col[5] 0.11fF
C8545 a_3270_18234# vcm 0.22fF
C8546 a_23046_2130# VDD 0.55fF
C8547 a_2346_4180# a_5978_4138# 0.19fF
C8548 a_1962_4178# a_4274_4178# 0.14fF
C8549 a_21038_5142# a_21038_4138# 1.00fF
C8550 m3_1864_10114# m3_1864_9110# 0.22fF
C8551 m2_34864_946# m3_34996_1078# 2.79fF
C8552 a_1962_9198# a_24050_9158# 0.27fF
C8553 a_2346_11208# col[25] 0.15fF
C8554 a_13310_3174# vcm 0.22fF
C8555 a_22042_14178# a_23046_14178# 0.97fF
C8556 a_15014_11166# row_n[9] 0.17fF
C8557 a_4974_10162# rowoff_n[8] 0.10fF
C8558 a_33086_13174# vcm 0.62fF
C8559 a_6982_13174# rowoff_n[11] 0.10fF
C8560 col[24] rowoff_n[13] 0.11fF
C8561 a_1962_13214# row_n[11] 25.57fF
C8562 a_2346_5184# VDD 32.63fF
C8563 a_10906_6146# a_10998_6146# 0.26fF
C8564 a_1962_6186# a_17326_6186# 0.14fF
C8565 a_2346_6188# a_19030_6146# 0.19fF
C8566 vcm rowoff_n[2] 0.20fF
C8567 a_15014_8154# rowoff_n[6] 0.10fF
C8568 a_8990_7150# col[6] 0.29fF
C8569 a_26362_7190# vcm 0.22fF
C8570 a_2346_1168# m2_1732_946# 0.12fF
C8571 a_21038_17190# rowoff_n[15] 0.10fF
C8572 a_25054_6146# rowoff_n[4] 0.10fF
C8573 a_21038_9158# m2_21236_9406# 0.16fF
C8574 a_1962_1166# col_n[3] 0.13fF
C8575 a_15926_9158# VDD 0.23fF
C8576 a_26058_16186# col_n[23] 0.28fF
C8577 a_34090_9158# a_34090_8154# 1.00fF
C8578 a_1962_14218# col_n[5] 0.13fF
C8579 a_2346_8196# a_32082_8154# 0.19fF
C8580 a_1962_8194# a_30378_8194# 0.14fF
C8581 a_34090_14178# row_n[12] 0.17fF
C8582 a_27062_3134# col[24] 0.29fF
C8583 a_1962_18234# a_6282_18234# 0.14fF
C8584 col[8] rowoff_n[14] 0.11fF
C8585 m2_8760_18014# m2_9764_18014# 0.96fF
C8586 a_21038_5142# ctop 3.58fF
C8587 m2_26832_946# ctop 0.18fF
C8588 a_28978_13174# VDD 0.23fF
C8589 a_23958_10162# a_24050_10162# 0.26fF
C8590 a_6982_10162# a_6982_9158# 1.00fF
C8591 a_2346_7192# col[16] 0.15fF
C8592 a_34394_5182# vcm 0.22fF
C8593 a_22042_12170# rowon_n[10] 0.14fF
C8594 a_2346_2172# a_21950_2130# 0.35fF
C8595 a_8990_9158# col_n[6] 0.28fF
C8596 a_34090_9158# ctop 3.42fF
C8597 a_7986_16186# VDD 0.52fF
C8598 m2_1732_11990# vcm 0.45fF
C8599 a_1962_3174# col[23] 0.11fF
C8600 VDD col_n[8] 4.98fF
C8601 vcm col_n[4] 2.80fF
C8602 ctop col[30] 1.99fF
C8603 a_15014_8154# vcm 0.62fF
C8604 a_1962_16226# col[25] 0.11fF
C8605 a_1962_16226# a_8990_16186# 0.27fF
C8606 a_27062_5142# col_n[24] 0.28fF
C8607 a_18026_1126# VDD 0.59fF
C8608 a_18026_10162# m2_18224_10410# 0.16fF
C8609 a_2346_4180# a_35002_4138# 0.35fF
C8610 a_18026_4138# a_19030_4138# 0.97fF
C8611 a_1962_10202# VDD 2.73fF
C8612 a_15014_2130# row_n[0] 0.17fF
C8613 a_14010_17190# m2_13780_18014# 1.00fF
C8614 a_8290_2170# vcm 0.22fF
C8615 a_2346_13216# a_3970_13174# 0.19fF
C8616 a_20034_14178# a_20034_13174# 1.00fF
C8617 a_33998_10162# rowoff_n[8] 0.24fF
C8618 a_28066_12170# vcm 0.62fF
C8619 a_1962_4178# row_n[2] 25.57fF
C8620 a_31078_5142# VDD 0.52fF
C8621 m3_23952_18146# VDD 0.29fF
C8622 a_2346_3176# col[7] 0.15fF
C8623 a_34090_17190# m3_34996_17142# 0.13fF
C8624 a_2346_16228# col[9] 0.15fF
C8625 a_19030_15182# row_n[13] 0.17fF
C8626 a_21342_6186# vcm 0.22fF
C8627 a_1962_15222# a_15318_15222# 0.14fF
C8628 a_9902_15182# a_9994_15182# 0.26fF
C8629 a_2346_15224# a_17022_15182# 0.19fF
C8630 a_1962_5182# col_n[23] 0.13fF
C8631 a_6982_12170# col[4] 0.29fF
C8632 a_34090_5142# row_n[3] 0.17fF
C8633 a_10906_8154# VDD 0.23fF
C8634 a_31078_8154# a_32082_8154# 0.97fF
C8635 a_1962_18234# a_1962_17230# 0.16fF
C8636 a_1962_12210# col[16] 0.11fF
C8637 a_35398_10202# vcm 0.23fF
C8638 a_1962_17230# a_28370_17230# 0.14fF
C8639 a_2346_17232# a_30074_17190# 0.19fF
C8640 a_25054_8154# col[22] 0.29fF
C8641 a_16018_4138# ctop 3.58fF
C8642 m2_4744_946# m3_3872_1078# 0.12fF
C8643 m3_30980_1078# ctop 0.23fF
C8644 a_15014_11166# m2_15212_11414# 0.16fF
C8645 a_6982_13174# rowon_n[11] 0.14fF
C8646 a_23958_12170# VDD 0.23fF
C8647 m3_14916_18146# m3_15920_18146# 0.22fF
C8648 a_3970_9158# a_4974_9158# 0.97fF
C8649 a_2346_9200# a_6890_9158# 0.35fF
C8650 a_7986_3134# rowoff_n[1] 0.10fF
C8651 a_2346_1168# m2_22816_946# 0.19fF
C8652 a_22042_3134# rowon_n[1] 0.14fF
C8653 a_23046_14178# rowoff_n[12] 0.10fF
C8654 a_29070_8154# ctop 3.58fF
C8655 a_2874_15182# VDD 0.24fF
C8656 a_6982_14178# col_n[4] 0.28fF
C8657 a_2346_11208# a_19942_11166# 0.35fF
C8658 a_2346_12212# col[0] 0.15fF
C8659 a_9994_7150# vcm 0.62fF
C8660 a_22042_2130# m2_22240_2378# 0.16fF
C8661 a_1962_1166# col_n[14] 0.13fF
C8662 a_2966_17190# rowoff_n[15] 0.10fF
C8663 a_26058_16186# rowon_n[14] 0.14fF
C8664 a_1962_14218# col_n[16] 0.13fF
C8665 a_32994_4138# a_33086_4138# 0.26fF
C8666 a_16018_4138# a_16018_3134# 1.00fF
C8667 a_25054_10162# col_n[22] 0.28fF
C8668 a_1962_8194# a_14010_8154# 0.27fF
C8669 a_33086_17190# m2_32856_18014# 1.00fF
C8670 a_2346_13216# a_32994_13174# 0.35fF
C8671 a_17022_13174# a_18026_13174# 0.97fF
C8672 a_3270_1166# vcm 0.23fF
C8673 a_1962_8194# col[7] 0.11fF
C8674 col[19] rowoff_n[14] 0.11fF
C8675 a_23046_11166# vcm 0.62fF
C8676 a_3970_16186# row_n[14] 0.17fF
C8677 a_2966_5142# ctop 3.42fF
C8678 a_26058_4138# VDD 0.52fF
C8679 a_5886_5142# a_5978_5142# 0.26fF
C8680 a_1962_5182# a_7286_5182# 0.14fF
C8681 a_2346_5184# a_8990_5142# 0.19fF
C8682 a_12002_12170# m2_12200_12418# 0.16fF
C8683 a_2346_7192# col[27] 0.15fF
C8684 a_19030_6146# row_n[4] 0.17fF
C8685 a_1962_10202# a_27062_10162# 0.27fF
C8686 a_6890_9158# rowoff_n[7] 0.24fF
C8687 a_16322_5182# vcm 0.22fF
C8688 a_10906_15182# rowoff_n[13] 0.24fF
C8689 a_2346_14220# vcm 0.40fF
C8690 a_7986_3134# col_n[5] 0.28fF
C8691 a_2346_2172# a_3878_2130# 0.35fF
C8692 m2_18800_18014# m3_17928_18146# 0.13fF
C8693 a_5886_7150# VDD 0.23fF
C8694 a_16930_7150# rowoff_n[5] 0.24fF
C8695 a_1962_7190# a_20338_7190# 0.14fF
C8696 a_29070_8154# a_29070_7150# 1.00fF
C8697 a_2346_7192# a_22042_7150# 0.19fF
C8698 col_n[7] col_n[8] 0.10fF
C8699 VDD col_n[19] 4.95fF
C8700 vcm col_n[15] 2.79fF
C8701 a_4974_17190# col[2] 0.29fF
C8702 col[17] col[18] 0.20fF
C8703 col[3] rowoff_n[15] 0.11fF
C8704 a_29374_9198# vcm 0.22fF
C8705 a_30074_17190# a_31078_17190# 0.97fF
C8706 a_26970_5142# rowoff_n[3] 0.24fF
C8707 a_6982_4138# rowon_n[2] 0.14fF
C8708 a_10998_3134# ctop 3.57fF
C8709 a_1962_10202# col_n[7] 0.13fF
C8710 m2_6752_18014# col_n[4] 0.25fF
C8711 a_23046_13174# col[20] 0.29fF
C8712 a_18938_11166# VDD 0.23fF
C8713 m3_4876_1078# m3_5880_1078# 0.22fF
C8714 a_1962_9198# a_33390_9198# 0.14fF
C8715 a_18938_9158# a_19030_9158# 0.26fF
C8716 a_1962_17230# col[0] 0.11fF
C8717 m2_34864_1950# VDD 1.06fF
C8718 a_2346_1168# a_11910_1126# 0.35fF
C8719 a_24050_7150# ctop 3.58fF
C8720 a_2346_3176# col[18] 0.15fF
C8721 a_8990_13174# m2_9188_13422# 0.16fF
C8722 a_2346_13216# m2_34864_12994# 0.17fF
C8723 a_10998_17190# rowon_n[15] 0.14fF
C8724 a_2346_16228# col[20] 0.15fF
C8725 a_31990_15182# VDD 0.23fF
C8726 m2_16792_946# a_2346_1168# 0.19fF
C8727 a_4974_6146# vcm 0.62fF
C8728 a_26058_7150# rowon_n[5] 0.14fF
C8729 a_9902_1126# m2_9764_946# 0.16fF
C8730 a_5978_6146# col[3] 0.29fF
C8731 a_13006_3134# a_14010_3134# 0.97fF
C8732 a_2346_3176# a_24962_3134# 0.35fF
C8733 a_15014_2130# m3_14916_1078# 0.15fF
C8734 a_2346_1168# m2_33860_946# 0.11fF
C8735 m2_11772_946# m2_10768_946# 0.96fF
C8736 a_1962_12210# col[27] 0.11fF
C8737 a_31990_13174# a_32082_13174# 0.26fF
C8738 a_15014_13174# a_15014_12170# 1.00fF
C8739 a_3970_7150# row_n[5] 0.17fF
C8740 a_23046_15182# col_n[20] 0.28fF
C8741 a_18026_10162# vcm 0.62fF
C8742 a_1962_17230# a_12002_17190# 0.27fF
C8743 a_25054_11166# rowoff_n[9] 0.10fF
C8744 a_24050_2130# col[21] 0.29fF
C8745 a_1962_6186# sample 0.14fF
C8746 m2_19804_18014# m2_20232_18442# 0.16fF
C8747 a_21038_3134# VDD 0.52fF
C8748 m3_26964_18146# ctop 0.23fF
C8749 a_2966_5142# a_2966_4138# 1.00fF
C8750 a_4882_14178# a_4974_14178# 0.26fF
C8751 a_2346_14220# a_6982_14178# 0.19fF
C8752 a_1962_14218# a_5278_14218# 0.14fF
C8753 a_11302_4178# vcm 0.22fF
C8754 a_31078_14178# vcm 0.62fF
C8755 a_1962_2170# a_32082_2130# 0.27fF
C8756 a_34090_7150# VDD 0.54fF
C8757 a_26058_7150# a_27062_7150# 0.97fF
C8758 a_5978_14178# m2_6176_14426# 0.16fF
C8759 a_2346_12212# col[11] 0.15fF
C8760 a_23046_10162# row_n[8] 0.17fF
C8761 a_5978_8154# col_n[3] 0.28fF
C8762 a_1962_1166# col_n[25] 0.13fF
C8763 a_24354_8194# vcm 0.22fF
C8764 a_2346_16228# a_20034_16186# 0.19fF
C8765 a_28066_17190# a_28066_16186# 1.00fF
C8766 a_1962_16226# a_18330_16226# 0.14fF
C8767 a_1962_14218# col_n[27] 0.13fF
C8768 a_5978_2130# ctop 3.39fF
C8769 a_1962_18234# m2_3740_18014# 0.18fF
C8770 a_24050_4138# col_n[21] 0.28fF
C8771 a_13918_10162# VDD 0.23fF
C8772 col[30] rowoff_n[14] 0.11fF
C8773 a_1962_8194# col[18] 0.11fF
C8774 a_12914_12170# rowoff_n[10] 0.24fF
C8775 a_10998_8154# rowon_n[6] 0.14fF
C8776 a_19030_6146# ctop 3.58fF
C8777 m3_2868_2082# VDD 0.19fF
C8778 a_26970_14178# VDD 0.23fF
C8779 a_2346_10204# a_9902_10162# 0.35fF
C8780 a_9902_2130# rowoff_n[0] 0.24fF
C8781 m2_25828_18014# ctop 0.18fF
C8782 a_26970_16186# rowoff_n[14] 0.24fF
C8783 a_27974_3134# a_28066_3134# 0.26fF
C8784 a_10998_3134# a_10998_2130# 1.00fF
C8785 a_32082_10162# ctop 3.58fF
C8786 vcm col_n[26] 2.80fF
C8787 VDD col_n[30] 4.97fF
C8788 col[14] rowoff_n[15] 0.11fF
C8789 a_2346_8196# col[2] 0.15fF
C8790 a_1962_7190# a_3970_7150# 0.27fF
C8791 a_3970_11166# col[1] 0.29fF
C8792 a_5978_17190# VDD 0.55fF
C8793 sample_n rowoff_n[11] 0.38fF
C8794 a_2346_12212# a_22954_12170# 0.35fF
C8795 a_12002_12170# a_13006_12170# 0.97fF
C8796 m2_13780_946# m3_14916_1078# 0.13fF
C8797 a_30074_11166# rowon_n[9] 0.14fF
C8798 a_1962_10202# col_n[18] 0.13fF
C8799 a_13006_9158# vcm 0.62fF
C8800 a_4974_3134# m2_5172_3382# 0.16fF
C8801 a_16018_2130# VDD 0.55fF
C8802 a_22042_7150# col[19] 0.29fF
C8803 a_1962_4178# col[9] 0.11fF
C8804 m2_25828_946# m3_24956_1078# 0.13fF
C8805 m3_1864_17142# m3_1864_16138# 0.22fF
C8806 a_1962_9198# a_17022_9158# 0.27fF
C8807 a_1962_17230# col[11] 0.11fF
C8808 a_12914_18194# m2_12776_18014# 0.16fF
C8809 a_7986_11166# row_n[9] 0.17fF
C8810 a_6282_3174# vcm 0.22fF
C8811 a_26058_13174# vcm 0.62fF
C8812 m2_1732_2954# VDD 1.02fF
C8813 a_2346_3176# col[29] 0.15fF
C8814 a_2346_16228# col[31] 0.15fF
C8815 a_29070_6146# VDD 0.52fF
C8816 m2_21812_946# m2_22816_946# 0.96fF
C8817 a_2346_6188# a_12002_6146# 0.19fF
C8818 a_1962_6186# a_10298_6186# 0.14fF
C8819 a_24050_7150# a_24050_6146# 1.00fF
C8820 a_7986_8154# rowoff_n[6] 0.10fF
C8821 a_1962_11206# a_30074_11166# 0.27fF
C8822 a_25054_16186# a_26058_16186# 0.97fF
C8823 a_19334_7190# vcm 0.22fF
C8824 a_3970_13174# col_n[1] 0.28fF
C8825 a_14010_17190# rowoff_n[15] 0.10fF
C8826 a_18026_6146# rowoff_n[4] 0.10fF
C8827 a_8898_9158# VDD 0.23fF
C8828 a_1962_8194# a_23350_8194# 0.14fF
C8829 a_2346_8196# a_25054_8154# 0.19fF
C8830 a_34090_17190# m2_34288_17438# 0.16fF
C8831 a_13918_8154# a_14010_8154# 0.26fF
C8832 a_27062_14178# row_n[12] 0.17fF
C8833 a_22042_9158# col_n[19] 0.28fF
C8834 a_1962_6186# col_n[9] 0.13fF
C8835 a_32386_11206# vcm 0.22fF
C8836 a_28066_4138# rowoff_n[2] 0.10fF
C8837 m2_1732_18014# sample_n 0.13fF
C8838 m2_1732_18014# m2_2736_18014# 0.96fF
C8839 a_14010_5142# ctop 3.58fF
C8840 a_2966_3134# VDD 0.56fF
C8841 a_21950_13174# VDD 0.23fF
C8842 a_1962_13214# col[2] 0.11fF
C8843 m2_1732_7974# m2_2160_8402# 0.16fF
C8844 a_15014_12170# rowon_n[10] 0.14fF
C8845 a_2346_12212# col[22] 0.15fF
C8846 a_7986_2130# a_8990_2130# 0.97fF
C8847 a_2346_2172# a_14922_2130# 0.35fF
C8848 m2_32856_18014# m3_32988_18146# 2.78fF
C8849 a_27062_9158# ctop 3.58fF
C8850 a_4974_2130# col_n[2] 0.28fF
C8851 a_30074_2130# rowon_n[0] 0.14fF
C8852 a_35002_17190# VDD 0.30fF
C8853 a_26970_12170# a_27062_12170# 0.26fF
C8854 a_9994_12170# a_9994_11166# 1.00fF
C8855 a_1962_14218# rowon_n[12] 1.18fF
C8856 a_7986_8154# vcm 0.62fF
C8857 a_1962_8194# col[29] 0.11fF
C8858 a_2346_4180# a_27974_4138# 0.35fF
C8859 a_7986_2130# row_n[0] 0.17fF
C8860 a_31990_18194# m2_31852_18014# 0.16fF
C8861 a_20034_12170# col[17] 0.29fF
C8862 m2_15788_946# VDD 0.62fF
C8863 a_1962_2170# vcm 6.97fF
C8864 a_26970_10162# rowoff_n[8] 0.24fF
C8865 a_1962_15222# col_n[2] 0.13fF
C8866 a_34090_15182# rowon_n[13] 0.14fF
C8867 a_28978_13174# rowoff_n[11] 0.24fF
C8868 a_21038_12170# vcm 0.62fF
C8869 a_33086_6146# m2_33284_6394# 0.16fF
C8870 m2_21812_18014# col[19] 0.28fF
C8871 a_24050_5142# VDD 0.52fF
C8872 m2_32856_946# VDD 0.64fF
C8873 a_21038_6146# a_22042_6146# 0.97fF
C8874 a_29070_17190# m3_28972_18146# 0.15fF
C8875 a_12002_15182# row_n[13] 0.17fF
C8876 a_14314_6186# vcm 0.22fF
C8877 a_1962_15222# a_8290_15222# 0.14fF
C8878 a_2346_15224# a_9994_15182# 0.19fF
C8879 a_23046_16186# a_23046_15182# 1.00fF
C8880 m2_34864_11990# m2_34864_10986# 0.99fF
C8881 sample row_n[12] 1.03fF
C8882 col_n[18] col_n[19] 0.10fF
C8883 col_n[4] row_n[15] 0.23fF
C8884 col_n[2] row_n[14] 0.23fF
C8885 VDD row_n[11] 2.93fF
C8886 vcm row_n[13] 0.49fF
C8887 col[25] rowoff_n[15] 0.11fF
C8888 col[28] col[29] 0.20fF
C8889 a_2346_8196# col[13] 0.15fF
C8890 a_34090_16186# vcm 0.62fF
C8891 a_27062_5142# row_n[3] 0.17fF
C8892 a_1962_10202# col_n[29] 0.13fF
C8893 a_2966_12170# a_3970_12170# 0.97fF
C8894 a_1962_17230# a_21342_17230# 0.14fF
C8895 a_12914_17190# a_13006_17190# 0.26fF
C8896 a_27366_10202# vcm 0.22fF
C8897 a_2346_17232# a_23046_17190# 0.19fF
C8898 a_20034_14178# col_n[17] 0.28fF
C8899 a_8990_4138# ctop 3.58fF
C8900 a_1962_4178# col[20] 0.11fF
C8901 a_1962_17230# col[22] 0.11fF
C8902 a_2346_9200# row_n[7] 0.35fF
C8903 a_16930_12170# VDD 0.23fF
C8904 a_15014_3134# rowon_n[1] 0.14fF
C8905 a_16018_14178# rowoff_n[12] 0.10fF
C8906 a_22954_2130# a_23046_2130# 0.26fF
C8907 a_30074_7150# m2_30272_7398# 0.16fF
C8908 a_22042_8154# ctop 3.58fF
C8909 a_1962_5182# rowon_n[3] 1.18fF
C8910 a_29982_16186# VDD 0.23fF
C8911 a_2346_11208# a_12914_11166# 0.35fF
C8912 a_6982_11166# a_7986_11166# 0.97fF
C8913 a_2346_4180# col[4] 0.15fF
C8914 a_2346_17232# col[6] 0.15fF
C8915 a_19030_16186# rowon_n[14] 0.14fF
C8916 a_1962_8194# a_6982_8154# 0.27fF
C8917 a_1962_6186# col_n[20] 0.13fF
C8918 a_34090_6146# rowon_n[4] 0.14fF
C8919 a_21038_3134# col_n[18] 0.28fF
C8920 a_2346_13216# a_25966_13174# 0.35fF
C8921 a_16018_11166# vcm 0.62fF
C8922 a_18026_17190# col[15] 0.29fF
C8923 a_1962_13214# col[13] 0.11fF
C8924 m2_34864_9982# row_n[8] 0.15fF
C8925 a_19030_4138# VDD 0.52fF
C8926 a_19030_6146# a_19030_5142# 1.00fF
C8927 a_12002_6146# row_n[4] 0.17fF
C8928 a_3878_13174# VDD 0.23fF
C8929 a_1962_10202# a_20034_10162# 0.27fF
C8930 a_2966_10162# col[0] 0.29fF
C8931 a_20034_15182# a_21038_15182# 0.97fF
C8932 a_9294_5182# vcm 0.22fF
C8933 a_29070_15182# vcm 0.62fF
C8934 a_27062_8154# m2_27260_8402# 0.16fF
C8935 m2_8760_18014# m3_9896_18146# 0.13fF
C8936 a_32082_8154# VDD 0.52fF
C8937 a_9902_7150# rowoff_n[5] 0.24fF
C8938 a_2346_7192# a_15014_7150# 0.19fF
C8939 a_8898_7150# a_8990_7150# 0.26fF
C8940 a_1962_7190# a_13310_7190# 0.14fF
C8941 a_1962_12210# a_33086_12170# 0.27fF
C8942 a_22346_9198# vcm 0.22fF
C8943 a_19942_5142# rowoff_n[3] 0.24fF
C8944 a_3970_3134# ctop 3.56fF
C8945 a_31078_9158# row_n[7] 0.17fF
C8946 a_11910_11166# VDD 0.23fF
C8947 a_1962_2170# col_n[11] 0.13fF
C8948 a_2346_9200# a_28066_9158# 0.19fF
C8949 a_1962_9198# a_26362_9198# 0.14fF
C8950 a_32082_10162# a_32082_9158# 1.00fF
C8951 a_1962_15222# col_n[13] 0.13fF
C8952 a_19030_6146# col[16] 0.29fF
C8953 a_29982_3134# rowoff_n[1] 0.24fF
C8954 m2_1732_15002# sample 0.19fF
C8955 m2_34864_8978# ctop 0.17fF
C8956 a_2966_12170# vcm 0.61fF
C8957 a_2346_1168# a_4882_1126# 0.35fF
C8958 a_1962_9198# col[4] 0.11fF
C8959 a_2346_1168# col_n[31] 0.11fF
C8960 a_17022_7150# ctop 3.58fF
C8961 a_3970_17190# rowon_n[15] 0.14fF
C8962 a_24962_15182# VDD 0.23fF
C8963 a_21950_11166# a_22042_11166# 0.26fF
C8964 a_4974_11166# a_4974_10162# 1.00fF
C8965 col_n[7] row_n[11] 0.23fF
C8966 col_n[11] row_n[13] 0.23fF
C8967 col_n[1] row_n[8] 0.23fF
C8968 col_n[5] row_n[10] 0.23fF
C8969 col_n[9] row_n[12] 0.23fF
C8970 col_n[15] row_n[15] 0.23fF
C8971 VDD rowon_n[5] 2.61fF
C8972 col_n[3] row_n[9] 0.23fF
C8973 vcm rowon_n[7] 0.50fF
C8974 col_n[0] row_n[7] 0.23fF
C8975 col_n[13] row_n[14] 0.23fF
C8976 a_2346_8196# col[24] 0.15fF
C8977 a_19030_7150# rowon_n[5] 0.14fF
C8978 a_2346_1168# m2_9764_946# 0.19fF
C8979 a_24050_9158# m2_24248_9406# 0.16fF
C8980 a_2346_3176# a_17934_3134# 0.35fF
C8981 a_30074_11166# ctop 3.58fF
C8982 a_1962_8194# a_34394_8194# 0.14fF
C8983 a_1962_4178# col[31] 0.11fF
C8984 a_18026_11166# rowoff_n[9] 0.10fF
C8985 a_10998_10162# vcm 0.62fF
C8986 a_3878_17190# a_3970_17190# 0.26fF
C8987 a_1962_17230# a_4974_17190# 0.27fF
C8988 a_19030_8154# col_n[16] 0.28fF
C8989 m2_12776_18014# m2_13204_18442# 0.16fF
C8990 a_14010_3134# VDD 0.52fF
C8991 m2_34864_946# ctop 0.11fF
C8992 a_16018_5142# a_17022_5142# 0.97fF
C8993 a_2346_5184# a_30986_5142# 0.35fF
C8994 a_1962_11206# col_n[4] 0.13fF
C8995 a_28066_9158# rowoff_n[7] 0.10fF
C8996 a_4274_4178# vcm 0.22fF
C8997 a_18026_15182# a_18026_14178# 1.00fF
C8998 a_24050_14178# vcm 0.62fF
C8999 a_32082_15182# rowoff_n[13] 0.10fF
C9000 a_1962_2170# a_25054_2130# 0.27fF
C9001 a_27062_7150# VDD 0.52fF
C9002 a_16018_10162# row_n[8] 0.17fF
C9003 a_2346_4180# col[15] 0.15fF
C9004 a_2346_17232# col[17] 0.15fF
C9005 a_2346_16228# a_13006_16186# 0.19fF
C9006 a_7894_16186# a_7986_16186# 0.26fF
C9007 a_1962_16226# a_11302_16226# 0.14fF
C9008 a_17326_8194# vcm 0.22fF
C9009 a_1962_2170# m2_1732_1950# 0.15fF
C9010 a_1962_6186# col_n[31] 0.13fF
C9011 a_21038_10162# m2_21236_10410# 0.16fF
C9012 a_6890_10162# VDD 0.23fF
C9013 a_29070_9158# a_30074_9158# 0.97fF
C9014 a_1962_13214# col[24] 0.11fF
C9015 a_30378_12210# vcm 0.22fF
C9016 a_5886_12170# rowoff_n[10] 0.24fF
C9017 a_17022_11166# col[14] 0.29fF
C9018 rowon_n[3] rowoff_n[3] 20.27fF
C9019 a_3970_8154# rowon_n[6] 0.14fF
C9020 a_17934_1126# a_18026_1126# 0.27fF
C9021 a_1962_1166# a_31382_1166# 0.14fF
C9022 a_12002_6146# ctop 3.58fF
C9023 m3_34996_16138# VDD 0.26fF
C9024 a_19942_14178# VDD 0.23fF
C9025 a_2346_2172# rowoff_n[0] 4.09fF
C9026 m2_11772_18014# ctop 0.18fF
C9027 a_19942_16186# rowoff_n[14] 0.24fF
C9028 a_25054_10162# ctop 3.58fF
C9029 a_32994_18194# VDD 0.33fF
C9030 a_2346_12212# a_15926_12170# 0.35fF
C9031 a_2346_13216# col[8] 0.15fF
C9032 a_23046_11166# rowon_n[9] 0.14fF
C9033 a_5978_9158# vcm 0.62fF
C9034 m2_9764_946# m3_8892_1078# 0.13fF
C9035 a_8990_2130# VDD 0.55fF
C9036 a_1962_2170# col_n[22] 0.13fF
C9037 a_30986_5142# a_31078_5142# 0.26fF
C9038 a_14010_5142# a_14010_4138# 1.00fF
C9039 a_1962_15222# col_n[24] 0.13fF
C9040 a_18026_11166# m2_18224_11414# 0.16fF
C9041 a_17022_13174# col_n[14] 0.28fF
C9042 a_1962_9198# a_9994_9158# 0.27fF
C9043 a_15014_14178# a_16018_14178# 0.97fF
C9044 a_2346_14220# a_28978_14178# 0.35fF
C9045 a_1962_9198# col[15] 0.11fF
C9046 a_19030_13174# vcm 0.62fF
C9047 a_22042_6146# VDD 0.52fF
C9048 a_2346_6188# a_4974_6146# 0.19fF
C9049 a_1962_6186# a_3270_6186# 0.14fF
C9050 col_n[20] row_n[12] 0.23fF
C9051 col_n[16] row_n[10] 0.23fF
C9052 col_n[2] row_n[3] 0.23fF
C9053 sample row_n[1] 1.03fF
C9054 col_n[22] row_n[13] 0.23fF
C9055 col_n[8] row_n[6] 0.23fF
C9056 vcm row_n[2] 0.49fF
C9057 col_n[24] row_n[14] 0.23fF
C9058 col_n[4] row_n[4] 0.23fF
C9059 col_n[12] row_n[8] 0.23fF
C9060 col_n[26] row_n[15] 0.23fF
C9061 VDD row_n[0] 3.02fF
C9062 col_n[6] row_n[5] 0.23fF
C9063 col_n[18] row_n[11] 0.23fF
C9064 col_n[29] col_n[30] 0.11fF
C9065 col_n[10] row_n[7] 0.23fF
C9066 col_n[14] row_n[9] 0.23fF
C9067 a_1962_11206# a_23046_11166# 0.27fF
C9068 a_12306_7190# vcm 0.22fF
C9069 a_25054_2130# m2_25252_2378# 0.16fF
C9070 a_6982_17190# rowoff_n[15] 0.10fF
C9071 a_32082_17190# vcm 0.60fF
C9072 m2_31852_18014# VDD 1.04fF
C9073 a_10998_6146# rowoff_n[4] 0.10fF
C9074 a_2346_8196# a_18026_8154# 0.19fF
C9075 a_27062_9158# a_27062_8154# 1.00fF
C9076 a_1962_8194# a_16322_8194# 0.14fF
C9077 a_20034_14178# row_n[12] 0.17fF
C9078 a_34090_12170# rowoff_n[10] 0.10fF
C9079 a_21038_4138# rowoff_n[2] 0.10fF
C9080 a_25358_11206# vcm 0.22fF
C9081 a_18026_2130# col_n[15] 0.26fF
C9082 a_1962_18234# sample 0.14fF
C9083 a_6982_5142# ctop 3.58fF
C9084 a_1962_11206# col_n[15] 0.13fF
C9085 a_15014_12170# m2_15212_12418# 0.16fF
C9086 a_15014_16186# col[12] 0.29fF
C9087 a_14922_13174# VDD 0.23fF
C9088 a_2346_10204# a_31078_10162# 0.19fF
C9089 a_16930_10162# a_17022_10162# 0.26fF
C9090 a_1962_10202# a_29374_10202# 0.14fF
C9091 a_31078_2130# rowoff_n[0] 0.10fF
C9092 a_1962_5182# col[6] 0.11fF
C9093 m2_27836_946# vcm 0.42fF
C9094 a_7986_12170# rowon_n[10] 0.14fF
C9095 a_2346_2172# a_7894_2130# 0.35fF
C9096 a_33086_12170# col[30] 0.29fF
C9097 m2_23820_18014# m3_22948_18146# 0.13fF
C9098 a_20034_9158# ctop 3.58fF
C9099 a_2346_4180# col[26] 0.15fF
C9100 a_27974_17190# VDD 0.24fF
C9101 a_23046_2130# rowon_n[0] 0.14fF
C9102 a_2346_17232# col[28] 0.15fF
C9103 a_3970_1126# VDD 0.60fF
C9104 a_10998_4138# a_12002_4138# 0.97fF
C9105 a_2346_4180# a_20946_4138# 0.35fF
C9106 a_33086_13174# ctop 3.57fF
C9107 a_29982_14178# a_30074_14178# 0.26fF
C9108 a_13006_14178# a_13006_13174# 1.00fF
C9109 a_19942_10162# rowoff_n[8] 0.24fF
C9110 col[0] rowoff_n[8] 0.11fF
C9111 col[1] rowoff_n[9] 0.11fF
C9112 ctop rowoff_n[2] 0.60fF
C9113 a_27062_15182# rowon_n[13] 0.14fF
C9114 a_16018_5142# col[13] 0.29fF
C9115 a_21950_13174# rowoff_n[11] 0.24fF
C9116 a_14010_12170# vcm 0.62fF
C9117 m2_8760_946# VDD 0.62fF
C9118 a_1962_7190# col_n[6] 0.13fF
C9119 a_17022_5142# VDD 0.52fF
C9120 a_2346_6188# a_33998_6146# 0.35fF
C9121 a_12002_13174# m2_12200_13422# 0.16fF
C9122 a_29982_8154# rowoff_n[6] 0.24fF
C9123 a_35494_15544# VDD 0.11fF
C9124 a_33086_14178# col_n[30] 0.28fF
C9125 a_4974_15182# row_n[13] 0.17fF
C9126 a_7286_6186# vcm 0.22fF
C9127 a_2346_15224# a_2874_15182# 0.35fF
C9128 m2_22816_946# m3_23952_1078# 0.13fF
C9129 a_27062_16186# vcm 0.62fF
C9130 m2_34864_15002# VDD 1.01fF
C9131 a_20034_5142# row_n[3] 0.17fF
C9132 a_1962_3174# a_28066_3134# 0.27fF
C9133 a_30074_9158# VDD 0.52fF
C9134 a_24050_8154# a_25054_8154# 0.97fF
C9135 a_2346_13216# col[19] 0.15fF
C9136 m2_34864_11990# rowon_n[10] 0.13fF
C9137 a_20338_10202# vcm 0.22fF
C9138 a_1962_17230# a_14314_17230# 0.14fF
C9139 a_2346_17232# a_16018_17190# 0.19fF
C9140 m3_1864_14130# ctop 0.23fF
C9141 a_16018_7150# col_n[13] 0.28fF
C9142 a_9902_12170# VDD 0.23fF
C9143 a_1962_9198# col[26] 0.11fF
C9144 a_7986_3134# rowon_n[1] 0.14fF
C9145 m2_1732_11990# ctop 0.17fF
C9146 a_8990_14178# rowoff_n[12] 0.10fF
C9147 a_33390_14218# vcm 0.22fF
C9148 a_2346_2172# a_2346_1168# 0.21fF
C9149 a_1962_2170# a_35398_2170# 0.14fF
C9150 a_34090_3134# col_n[31] 0.28fF
C9151 col_n[23] row_n[8] 0.23fF
C9152 col_n[17] row_n[5] 0.23fF
C9153 col_n[27] row_n[10] 0.23fF
C9154 col_n[29] row_n[11] 0.23fF
C9155 col_n[4] ctop 2.02fF
C9156 col_n[25] row_n[9] 0.23fF
C9157 col_n[21] row_n[7] 0.23fF
C9158 col_n[9] row_n[1] 0.23fF
C9159 VDD col[2] 4.17fF
C9160 col_n[13] row_n[3] 0.23fF
C9161 col_n[15] row_n[4] 0.23fF
C9162 col_n[31] row_n[12] 0.23fF
C9163 rowon_n[14] rowon_n[13] 0.15fF
C9164 col_n[19] row_n[6] 0.23fF
C9165 col_n[11] row_n[2] 0.23fF
C9166 col_n[7] row_n[0] 0.23fF
C9167 a_1962_16226# col_n[0] 0.13fF
C9168 a_15014_8154# ctop 3.58fF
C9169 a_2346_14220# m2_34864_13998# 0.17fF
C9170 a_8990_14178# m2_9188_14426# 0.16fF
C9171 a_31078_17190# col[28] 0.29fF
C9172 a_22954_16186# VDD 0.23fF
C9173 a_2346_11208# a_5886_11166# 0.35fF
C9174 a_32994_1126# VDD 0.45fF
C9175 a_12002_16186# rowon_n[14] 0.14fF
C9176 a_8990_4138# a_8990_3134# 1.00fF
C9177 a_25966_4138# a_26058_4138# 0.26fF
C9178 a_28066_12170# ctop 3.58fF
C9179 a_2346_9200# col[10] 0.15fF
C9180 a_27062_6146# rowon_n[4] 0.14fF
C9181 a_2346_13216# a_18938_13174# 0.35fF
C9182 a_9994_13174# a_10998_13174# 0.97fF
C9183 a_1962_18234# col_n[9] 0.13fF
C9184 a_2966_4138# rowoff_n[2] 0.10fF
C9185 a_1962_11206# col_n[26] 0.13fF
C9186 a_8990_11166# vcm 0.62fF
C9187 m2_1732_13998# row_n[12] 0.13fF
C9188 a_12002_4138# VDD 0.52fF
C9189 m3_14916_1078# VDD 0.14fF
C9190 a_14010_10162# col[11] 0.29fF
C9191 a_4974_6146# row_n[4] 0.17fF
C9192 a_1962_5182# col[17] 0.11fF
C9193 a_1962_10202# a_13006_10162# 0.27fF
C9194 a_2346_10204# rowon_n[8] 0.26fF
C9195 a_2346_15224# a_31990_15182# 0.35fF
C9196 a_22042_15182# vcm 0.62fF
C9197 a_32082_6146# col[29] 0.29fF
C9198 a_25054_8154# VDD 0.52fF
C9199 a_2346_7192# rowoff_n[5] 4.09fF
C9200 a_1962_7190# a_6282_7190# 0.14fF
C9201 a_2346_7192# a_7986_7150# 0.19fF
C9202 a_22042_8154# a_22042_7150# 1.00fF
C9203 a_5978_15182# m2_6176_15430# 0.16fF
C9204 a_1962_12210# a_26058_12170# 0.27fF
C9205 a_15318_9198# vcm 0.22fF
C9206 a_23046_17190# a_24050_17190# 0.97fF
C9207 a_7986_3134# m2_8184_3382# 0.16fF
C9208 a_12914_5142# rowoff_n[3] 0.24fF
C9209 a_24050_9158# row_n[7] 0.17fF
C9210 a_2346_4180# a_1962_4178# 2.62fF
C9211 a_2346_5184# col[1] 0.15fF
C9212 a_4882_11166# VDD 0.23fF
C9213 m2_30848_946# m3_29976_1078# 0.13fF
C9214 a_1962_9198# a_19334_9198# 0.14fF
C9215 a_11910_9158# a_12002_9158# 0.26fF
C9216 a_2346_9200# a_21038_9158# 0.19fF
C9217 col[8] rowoff_n[5] 0.11fF
C9218 col[7] rowoff_n[4] 0.11fF
C9219 col[10] rowoff_n[7] 0.11fF
C9220 col[3] rowoff_n[0] 0.11fF
C9221 col[6] rowoff_n[3] 0.11fF
C9222 col[12] rowoff_n[9] 0.11fF
C9223 col[4] rowoff_n[1] 0.11fF
C9224 col[9] rowoff_n[6] 0.11fF
C9225 col[5] rowoff_n[2] 0.11fF
C9226 col[11] rowoff_n[8] 0.11fF
C9227 a_14010_12170# col_n[11] 0.28fF
C9228 a_22954_3134# rowoff_n[1] 0.24fF
C9229 a_1962_7190# col_n[17] 0.13fF
C9230 a_3878_13174# rowoff_n[11] 0.24fF
C9231 a_28370_13214# vcm 0.22fF
C9232 a_33086_2130# a_34090_2130# 0.97fF
C9233 a_9994_7150# ctop 3.58fF
C9234 a_1962_1166# col[8] 0.11fF
C9235 a_32082_8154# col_n[29] 0.28fF
C9236 a_17934_15182# VDD 0.23fF
C9237 a_1962_14218# col[10] 0.11fF
C9238 a_1962_11206# a_32386_11206# 0.14fF
C9239 a_2346_11208# a_34090_11166# 0.19fF
C9240 a_12002_7150# rowon_n[5] 0.14fF
C9241 a_2346_13216# col[30] 0.15fF
C9242 a_2346_3176# a_10906_3134# 0.35fF
C9243 a_5978_3134# a_6982_3134# 0.97fF
C9244 a_23046_11166# ctop 3.58fF
C9245 a_26058_2130# m2_25828_946# 0.99fF
C9246 a_24962_13174# a_25054_13174# 0.26fF
C9247 a_7986_13174# a_7986_12170# 1.00fF
C9248 a_10998_11166# rowoff_n[9] 0.10fF
C9249 a_3970_10162# vcm 0.62fF
C9250 m2_5748_18014# m2_6176_18442# 0.16fF
C9251 a_4974_4138# m2_5172_4386# 0.16fF
C9252 a_6982_3134# VDD 0.52fF
C9253 a_2346_5184# a_23958_5142# 0.35fF
C9254 a_2346_14220# ctop 1.59fF
C9255 a_31078_10162# rowon_n[8] 0.14fF
C9256 a_21038_9158# rowoff_n[7] 0.10fF
C9257 a_12002_15182# col[9] 0.29fF
C9258 a_1962_3174# col_n[8] 0.13fF
C9259 col_n[20] row_n[1] 0.23fF
C9260 col_n[18] row_n[0] 0.23fF
C9261 a_1962_16226# col_n[10] 0.13fF
C9262 rowon_n[11] row_n[11] 19.75fF
C9263 vcm col[9] 5.84fF
C9264 col_n[26] row_n[4] 0.23fF
C9265 col_n[24] row_n[3] 0.23fF
C9266 VDD col[13] 4.18fF
C9267 col_n[15] ctop 2.04fF
C9268 col_n[28] row_n[5] 0.23fF
C9269 col_n[30] row_n[6] 0.23fF
C9270 col_n[22] row_n[2] 0.23fF
C9271 col_n[4] col[5] 5.98fF
C9272 a_25054_15182# rowoff_n[13] 0.10fF
C9273 a_17022_14178# vcm 0.62fF
C9274 a_1962_2170# a_18026_2130# 0.27fF
C9275 a_20034_7150# VDD 0.52fF
C9276 a_31078_7150# rowoff_n[5] 0.10fF
C9277 a_19030_7150# a_20034_7150# 0.97fF
C9278 a_1962_7190# a_1962_6186# 0.16fF
C9279 a_30074_11166# col[27] 0.29fF
C9280 a_8990_10162# row_n[8] 0.17fF
C9281 a_1962_10202# col[1] 0.11fF
C9282 a_10298_8194# vcm 0.22fF
C9283 a_21038_17190# a_21038_16186# 1.00fF
C9284 a_2346_16228# a_5978_16186# 0.19fF
C9285 a_1962_16226# a_4274_16226# 0.14fF
C9286 m2_1732_15002# m2_1732_13998# 0.99fF
C9287 a_30074_18194# vcm 0.12fF
C9288 a_2346_9200# col[21] 0.15fF
C9289 a_1962_4178# a_31078_4138# 0.27fF
C9290 m2_34864_1950# rowon_n[0] 0.13fF
C9291 a_33086_11166# VDD 0.52fF
C9292 a_1962_18234# col_n[20] 0.13fF
C9293 a_23350_12210# vcm 0.22fF
C9294 a_12002_17190# col_n[9] 0.28fF
C9295 a_1962_1166# a_24354_1166# 0.14fF
C9296 a_4974_6146# ctop 3.58fF
C9297 a_28066_13174# row_n[11] 0.17fF
C9298 a_1962_5182# col[28] 0.11fF
C9299 a_13006_4138# col[10] 0.29fF
C9300 m3_10900_18146# VDD 0.36fF
C9301 a_12914_14178# VDD 0.23fF
C9302 m2_34864_4962# vcm 0.51fF
C9303 a_32082_11166# a_33086_11166# 0.97fF
C9304 a_32082_17190# m3_31984_18146# 0.15fF
C9305 a_1962_12210# col_n[1] 0.13fF
C9306 a_30074_13174# col_n[27] 0.28fF
C9307 a_12914_16186# rowoff_n[14] 0.24fF
C9308 a_3970_3134# a_3970_2130# 1.00fF
C9309 a_20946_3134# a_21038_3134# 0.26fF
C9310 a_18026_10162# ctop 3.58fF
C9311 a_25966_18194# VDD 0.33fF
C9312 m2_26832_18014# vcm 0.28fF
C9313 a_4974_12170# a_5978_12170# 0.97fF
C9314 a_2346_12212# a_8898_12170# 0.35fF
C9315 a_16018_11166# rowon_n[9] 0.14fF
C9316 a_2346_5184# col[12] 0.15fF
C9317 m2_34864_1950# m3_34996_3086# 0.15fF
C9318 m3_17928_1078# ctop 0.39fF
C9319 col[22] rowoff_n[8] 0.11fF
C9320 col[21] rowoff_n[7] 0.11fF
C9321 col[14] rowoff_n[0] 0.11fF
C9322 col[23] rowoff_n[9] 0.11fF
C9323 col[19] rowoff_n[5] 0.11fF
C9324 col[20] rowoff_n[6] 0.11fF
C9325 col[15] rowoff_n[1] 0.11fF
C9326 col[16] rowoff_n[2] 0.11fF
C9327 col[17] rowoff_n[3] 0.11fF
C9328 col[18] rowoff_n[4] 0.11fF
C9329 a_31078_14178# ctop 3.58fF
C9330 a_2346_9200# a_2966_9158# 0.21fF
C9331 a_1962_7190# col_n[28] 0.13fF
C9332 a_13006_6146# col_n[10] 0.28fF
C9333 a_2346_14220# a_21950_14178# 0.35fF
C9334 a_2346_18236# a_30986_18194# 0.35fF
C9335 a_12002_13174# vcm 0.62fF
C9336 a_33086_7150# m2_33284_7398# 0.16fF
C9337 a_1962_1166# col[19] 0.11fF
C9338 a_15014_6146# VDD 0.52fF
C9339 a_1962_14218# col[21] 0.11fF
C9340 a_33998_7150# a_34090_7150# 0.26fF
C9341 a_17022_7150# a_17022_6146# 1.00fF
C9342 a_31078_2130# col_n[28] 0.29fF
C9343 a_1962_11206# a_16018_11166# 0.27fF
C9344 a_2346_16228# a_35002_16186# 0.35fF
C9345 a_18026_16186# a_19030_16186# 0.97fF
C9346 a_5278_7190# vcm 0.22fF
C9347 a_28066_16186# col[25] 0.29fF
C9348 m2_15788_18014# col[13] 0.28fF
C9349 m2_1732_6970# sample_n 0.15fF
C9350 a_25054_17190# vcm 0.60fF
C9351 m2_17796_18014# VDD 0.93fF
C9352 col[7] rowoff_n[10] 0.11fF
C9353 a_3970_6146# rowoff_n[4] 0.10fF
C9354 a_1962_18234# m2_32856_18014# 0.18fF
C9355 a_28066_10162# VDD 0.52fF
C9356 a_1962_8194# a_9294_8194# 0.14fF
C9357 a_2346_8196# a_10998_8154# 0.19fF
C9358 a_6890_8154# a_6982_8154# 0.26fF
C9359 a_13006_14178# row_n[12] 0.17fF
C9360 a_1962_13214# a_29070_13174# 0.27fF
C9361 a_35094_2130# vcm 0.12fF
C9362 m2_34864_2954# m2_35292_3382# 0.16fF
C9363 a_27062_12170# rowoff_n[10] 0.10fF
C9364 a_14010_4138# rowoff_n[2] 0.10fF
C9365 a_18330_11206# vcm 0.22fF
C9366 a_28066_4138# row_n[2] 0.17fF
C9367 a_2346_1168# col[3] 0.14fF
C9368 a_2346_14220# col[5] 0.15fF
C9369 a_7894_13174# VDD 0.23fF
C9370 a_2346_18236# m2_27836_18014# 0.19fF
C9371 a_30074_11166# a_30074_10162# 1.00fF
C9372 a_1962_10202# a_22346_10202# 0.14fF
C9373 a_1962_3174# col_n[19] 0.13fF
C9374 a_2346_10204# a_24050_10162# 0.19fF
C9375 col_n[10] col[10] 0.72fF
C9376 a_24050_2130# rowoff_n[0] 0.10fF
C9377 vcm col[20] 5.84fF
C9378 a_2966_9158# rowoff_n[7] 0.10fF
C9379 a_1962_16226# col_n[21] 0.13fF
C9380 col_n[31] row_n[1] 0.23fF
C9381 a_10998_9158# col[8] 0.29fF
C9382 VDD col[24] 4.17fF
C9383 col_n[29] row_n[0] 0.23fF
C9384 col_n[26] ctop 2.02fF
C9385 m2_5748_946# col[3] 0.39fF
C9386 a_31382_15222# vcm 0.22fF
C9387 a_30074_8154# m2_30272_8402# 0.16fF
C9388 a_1962_10202# col[12] 0.11fF
C9389 a_13006_9158# ctop 3.58fF
C9390 m2_13780_18014# m3_14916_18146# 0.13fF
C9391 a_32082_17190# row_n[15] 0.17fF
C9392 m2_31852_18014# col_n[29] 0.25fF
C9393 a_29070_5142# col[26] 0.29fF
C9394 a_16018_2130# rowon_n[0] 0.14fF
C9395 a_20946_17190# VDD 0.24fF
C9396 a_20034_1126# en_bit_n[0] 0.25fF
C9397 a_19942_12170# a_20034_12170# 0.26fF
C9398 a_30986_2130# VDD 0.23fF
C9399 a_1962_18234# col_n[31] 0.13fF
C9400 a_2346_4180# a_13918_4138# 0.35fF
C9401 a_26058_13174# ctop 3.58fF
C9402 a_12914_10162# rowoff_n[8] 0.24fF
C9403 a_20034_15182# rowon_n[13] 0.14fF
C9404 a_14922_13174# rowoff_n[11] 0.24fF
C9405 a_6982_12170# vcm 0.62fF
C9406 a_10998_11166# col_n[8] 0.28fF
C9407 a_9994_5142# VDD 0.52fF
C9408 a_14010_6146# a_15014_6146# 0.97fF
C9409 a_2346_6188# a_26970_6146# 0.35fF
C9410 a_22954_8154# rowoff_n[6] 0.24fF
C9411 a_1962_12210# col_n[12] 0.13fF
C9412 a_29070_7150# col_n[26] 0.28fF
C9413 a_32994_16186# a_33086_16186# 0.26fF
C9414 a_16018_16186# a_16018_15182# 1.00fF
C9415 a_2966_9158# col_n[0] 0.28fF
C9416 a_28978_17190# rowoff_n[15] 0.24fF
C9417 a_20034_16186# vcm 0.62fF
C9418 a_1962_6186# col[3] 0.11fF
C9419 a_1962_3174# a_21038_3134# 0.27fF
C9420 a_32994_6146# rowoff_n[4] 0.24fF
C9421 a_13006_5142# row_n[3] 0.17fF
C9422 a_27062_9158# m2_27260_9406# 0.16fF
C9423 a_1962_1166# m2_26832_946# 0.18fF
C9424 a_23046_9158# VDD 0.52fF
C9425 a_30074_1126# vcm 0.12fF
C9426 m2_1732_16006# rowon_n[14] 0.11fF
C9427 a_2346_5184# col[23] 0.15fF
C9428 a_1962_17230# a_7286_17230# 0.14fF
C9429 a_13310_10202# vcm 0.22fF
C9430 a_5886_17190# a_5978_17190# 0.26fF
C9431 a_2346_17232# a_8990_17190# 0.19fF
C9432 col[29] rowoff_n[4] 0.11fF
C9433 col[27] rowoff_n[2] 0.11fF
C9434 col[25] rowoff_n[0] 0.11fF
C9435 col[31] rowoff_n[6] 0.11fF
C9436 col[26] rowoff_n[1] 0.11fF
C9437 col[28] rowoff_n[3] 0.11fF
C9438 col[30] rowoff_n[5] 0.11fF
C9439 m3_13912_18146# ctop 0.23fF
C9440 a_1962_5182# a_34090_5142# 0.27fF
C9441 a_2346_12212# VDD 32.63fF
C9442 a_27062_10162# a_28066_10162# 0.97fF
C9443 a_2874_14178# a_2966_14178# 0.26fF
C9444 a_2346_14220# a_3878_14178# 0.35fF
C9445 a_1962_1166# col[30] 0.11fF
C9446 a_32082_8154# row_n[6] 0.17fF
C9447 a_26362_14218# vcm 0.22fF
C9448 a_8990_14178# col[6] 0.29fF
C9449 a_1962_2170# a_27366_2170# 0.14fF
C9450 a_2346_2172# a_29070_2130# 0.19fF
C9451 a_15926_2130# a_16018_2130# 0.26fF
C9452 a_7986_8154# ctop 3.58fF
C9453 a_15926_16186# VDD 0.23fF
C9454 a_1962_8194# col_n[3] 0.13fF
C9455 a_27062_10162# col[24] 0.29fF
C9456 col[18] rowoff_n[10] 0.11fF
C9457 a_1962_2170# ctop 1.18fF
C9458 a_25966_1126# VDD 0.44fF
C9459 a_4974_16186# rowon_n[14] 0.14fF
C9460 a_24050_10162# m2_24248_10410# 0.16fF
C9461 a_21038_12170# ctop 3.58fF
C9462 a_19030_17190# m2_18800_18014# 1.00fF
C9463 a_20034_6146# rowon_n[4] 0.14fF
C9464 a_2346_13216# a_11910_13174# 0.35fF
C9465 a_2346_1168# col[14] 0.14fF
C9466 a_2346_14220# col[16] 0.15fF
C9467 a_34394_12210# vcm 0.22fF
C9468 m2_1732_7974# rowoff_n[6] 0.12fF
C9469 a_4974_4138# VDD 0.52fF
C9470 a_1962_3174# col_n[30] 0.13fF
C9471 m3_1864_8106# VDD 0.25fF
C9472 a_28978_6146# a_29070_6146# 0.26fF
C9473 a_12002_6146# a_12002_5142# 1.00fF
C9474 vcm col[31] 5.56fF
C9475 col_n[15] col[16] 6.03fF
C9476 row_n[13] ctop 1.65fF
C9477 a_8990_16186# col_n[6] 0.28fF
C9478 a_34090_16186# ctop 3.41fF
C9479 a_1962_10202# a_5978_10162# 0.27fF
C9480 a_9994_3134# col[7] 0.29fF
C9481 col[2] rowoff_n[11] 0.11fF
C9482 a_2346_15224# a_24962_15182# 0.35fF
C9483 a_13006_15182# a_14010_15182# 0.97fF
C9484 a_1962_10202# col[23] 0.11fF
C9485 a_15014_15182# vcm 0.62fF
C9486 a_27062_12170# col_n[24] 0.28fF
C9487 a_18026_8154# VDD 0.52fF
C9488 a_1962_17230# VDD 2.78fF
C9489 a_1962_12210# a_19030_12170# 0.27fF
C9490 a_8290_9198# vcm 0.22fF
C9491 a_2966_17190# a_2966_16186# 1.00fF
C9492 a_1962_3174# m2_1732_2954# 0.15fF
C9493 a_5886_5142# rowoff_n[3] 0.24fF
C9494 a_17022_9158# row_n[7] 0.17fF
C9495 a_21038_11166# m2_21236_11414# 0.16fF
C9496 a_31078_12170# VDD 0.52fF
C9497 m3_29976_18146# m3_30980_18146# 0.22fF
C9498 a_1962_9198# a_12306_9198# 0.14fF
C9499 a_2346_9200# a_14010_9158# 0.19fF
C9500 a_25054_10162# a_25054_9158# 1.00fF
C9501 a_1962_14218# a_32082_14178# 0.27fF
C9502 a_2346_10204# col[7] 0.15fF
C9503 a_15926_3134# rowoff_n[1] 0.24fF
C9504 a_9994_5142# col_n[7] 0.28fF
C9505 a_21342_13214# vcm 0.22fF
C9506 a_30986_14178# rowoff_n[12] 0.24fF
C9507 a_1962_12210# col_n[23] 0.13fF
C9508 a_10906_15182# VDD 0.23fF
C9509 m2_1732_7974# vcm 0.45fF
C9510 a_14922_11166# a_15014_11166# 0.26fF
C9511 a_2346_11208# a_27062_11166# 0.19fF
C9512 a_1962_11206# a_25358_11206# 0.14fF
C9513 a_4974_7150# rowon_n[5] 0.14fF
C9514 a_1962_6186# col[14] 0.11fF
C9515 a_28066_2130# m2_28264_2378# 0.16fF
C9516 a_35398_17230# vcm 0.23fF
C9517 a_25054_15182# col[22] 0.29fF
C9518 a_1962_3174# a_2966_3134# 0.27fF
C9519 a_16018_11166# ctop 3.58fF
C9520 a_3970_11166# rowoff_n[9] 0.10fF
C9521 a_33998_4138# VDD 0.23fF
C9522 a_18026_12170# m2_18224_12418# 0.16fF
C9523 a_8990_5142# a_9994_5142# 0.97fF
C9524 a_2346_5184# a_16930_5142# 0.35fF
C9525 a_29070_15182# ctop 3.58fF
C9526 a_24050_10162# rowon_n[8] 0.14fF
C9527 a_14010_9158# rowoff_n[7] 0.10fF
C9528 a_27974_15182# a_28066_15182# 0.26fF
C9529 a_10998_15182# a_10998_14178# 1.00fF
C9530 a_7986_8154# col[5] 0.29fF
C9531 a_9994_14178# vcm 0.62fF
C9532 a_18026_15182# rowoff_n[13] 0.10fF
C9533 a_1962_2170# a_10998_2130# 0.27fF
C9534 m2_28840_18014# m3_27968_18146# 0.13fF
C9535 a_1962_8194# col_n[14] 0.13fF
C9536 a_13006_7150# VDD 0.52fF
C9537 a_24050_7150# rowoff_n[5] 0.10fF
C9538 a_2346_7192# a_29982_7150# 0.35fF
C9539 a_25054_17190# col_n[22] 0.28fF
C9540 col[29] rowoff_n[10] 0.11fF
C9541 a_26058_4138# col[23] 0.29fF
C9542 a_1962_2170# col[5] 0.11fF
C9543 a_3270_8194# vcm 0.22fF
C9544 a_1962_15222# col[7] 0.11fF
C9545 a_34090_5142# rowoff_n[3] 0.10fF
C9546 a_23046_18194# vcm 0.12fF
C9547 a_1962_4178# a_24050_4138# 0.27fF
C9548 a_2966_12170# ctop 3.42fF
C9549 a_26058_11166# VDD 0.52fF
C9550 m3_19936_1078# m3_20940_1078# 0.22fF
C9551 a_2346_1168# col[25] 0.14fF
C9552 a_22042_9158# a_23046_9158# 0.97fF
C9553 a_2346_14220# col[27] 0.15fF
C9554 a_33086_3134# vcm 0.62fF
C9555 a_16322_12210# vcm 0.22fF
C9556 rowon_n[3] rowon_n[2] 0.15fF
C9557 rowon_n[7] ctop 1.40fF
C9558 col_n[21] col[21] 0.72fF
C9559 a_2346_1168# a_19030_1126# 0.19fF
C9560 a_1962_1166# a_17326_1166# 0.14fF
C9561 a_21038_13174# row_n[11] 0.17fF
C9562 a_15014_13174# m2_15212_13422# 0.16fF
C9563 a_7986_10162# col_n[5] 0.28fF
C9564 col[13] rowoff_n[11] 0.11fF
C9565 a_5886_14178# VDD 0.23fF
C9566 m2_34864_2954# rowon_n[1] 0.13fF
C9567 a_29374_16226# vcm 0.22fF
C9568 a_5886_16186# rowoff_n[14] 0.24fF
C9569 a_26058_6146# col_n[23] 0.28fF
C9570 m2_14784_946# m2_15788_946# 0.96fF
C9571 a_1962_3174# a_30378_3174# 0.14fF
C9572 a_1962_4178# col_n[5] 0.13fF
C9573 a_2346_3176# a_32082_3134# 0.19fF
C9574 a_34090_4138# a_34090_3134# 1.00fF
C9575 a_1962_17230# col_n[7] 0.13fF
C9576 a_10998_10162# ctop 3.58fF
C9577 a_21038_2130# m3_20940_1078# 0.15fF
C9578 a_18938_18194# VDD 0.34fF
C9579 m2_12776_18014# vcm 0.28fF
C9580 a_8990_11166# rowon_n[9] 0.14fF
C9581 a_32994_11166# rowoff_n[9] 0.24fF
C9582 m2_2736_1950# m3_2868_1078# 0.15fF
C9583 a_28978_3134# VDD 0.23fF
C9584 m3_34996_7102# ctop 0.23fF
C9585 a_6982_5142# a_6982_4138# 1.00fF
C9586 a_23958_5142# a_24050_5142# 0.26fF
C9587 a_24050_14178# ctop 3.58fF
C9588 m2_31852_946# m2_32856_946# 0.96fF
C9589 a_2346_10204# col[18] 0.15fF
C9590 a_2346_14220# a_14922_14178# 0.35fF
C9591 a_7986_14178# a_8990_14178# 0.97fF
C9592 a_2346_18236# a_23958_18194# 0.35fF
C9593 a_4974_13174# vcm 0.62fF
C9594 a_7986_6146# VDD 0.52fF
C9595 a_5978_13174# col[3] 0.29fF
C9596 a_12002_14178# m2_12200_14426# 0.16fF
C9597 a_1962_6186# col[25] 0.11fF
C9598 a_28066_14178# rowon_n[12] 0.14fF
C9599 a_1962_11206# a_8990_11166# 0.27fF
C9600 a_2346_16228# a_27974_16186# 0.35fF
C9601 m2_1732_4962# row_n[3] 0.13fF
C9602 a_18026_17190# vcm 0.60fF
C9603 m2_3740_18014# VDD 1.09fF
C9604 a_24050_9158# col[21] 0.29fF
C9605 a_1962_18234# m2_18800_18014# 0.18fF
C9606 a_1962_13214# sample 0.14fF
C9607 a_21038_10162# VDD 0.52fF
C9608 a_20034_9158# a_20034_8154# 1.00fF
C9609 a_2346_8196# a_3970_8154# 0.19fF
C9610 a_5978_14178# row_n[12] 0.17fF
C9611 a_28066_2130# vcm 0.62fF
C9612 a_1962_13214# a_22042_13174# 0.27fF
C9613 a_11302_11206# vcm 0.22fF
C9614 a_20034_12170# rowoff_n[10] 0.10fF
C9615 a_6982_4138# rowoff_n[2] 0.10fF
C9616 a_21038_4138# row_n[2] 0.17fF
C9617 m3_29976_1078# VDD 0.14fF
C9618 a_2346_6188# col[9] 0.15fF
C9619 a_34090_14178# VDD 0.54fF
C9620 a_2346_18236# m2_13780_18014# 0.19fF
C9621 a_1962_10202# a_15318_10202# 0.14fF
C9622 a_9902_10162# a_9994_10162# 0.26fF
C9623 a_2346_10204# a_17022_10162# 0.19fF
C9624 a_17022_2130# rowoff_n[0] 0.10fF
C9625 a_5978_15182# col_n[3] 0.28fF
C9626 a_6982_2130# col[4] 0.29fF
C9627 a_1962_8194# col_n[25] 0.13fF
C9628 a_34090_16186# rowoff_n[14] 0.10fF
C9629 a_24354_15222# vcm 0.22fF
C9630 a_31078_3134# a_32082_3134# 0.97fF
C9631 a_5978_9158# ctop 3.58fF
C9632 m2_4744_18014# m3_4876_18146# 2.78fF
C9633 a_25054_17190# row_n[15] 0.17fF
C9634 a_8990_15182# m2_9188_15430# 0.16fF
C9635 a_2346_15224# m2_34864_15002# 0.17fF
C9636 a_24050_11166# col_n[21] 0.28fF
C9637 a_1962_2170# col[16] 0.11fF
C9638 m2_28840_946# col[26] 0.39fF
C9639 a_13918_17190# VDD 0.24fF
C9640 a_8990_2130# rowon_n[0] 0.14fF
C9641 a_33086_13174# a_33086_12170# 1.00fF
C9642 a_1962_15222# col[18] 0.11fF
C9643 a_2346_12212# a_30074_12170# 0.19fF
C9644 a_1962_12210# a_28370_12210# 0.14fF
C9645 a_10998_3134# m2_11196_3382# 0.16fF
C9646 a_23958_2130# VDD 0.23fF
C9647 a_2346_4180# a_6890_4138# 0.35fF
C9648 a_3970_4138# a_4974_4138# 0.97fF
C9649 a_19030_13174# ctop 3.58fF
C9650 m3_34996_10114# m3_34996_9110# 0.22fF
C9651 a_17934_18194# m2_17796_18014# 0.16fF
C9652 a_2346_18236# col[10] 0.14fF
C9653 a_22954_14178# a_23046_14178# 0.26fF
C9654 a_5978_14178# a_5978_13174# 1.00fF
C9655 a_5886_10162# rowoff_n[8] 0.24fF
C9656 rowon_n[0] row_n[0] 19.75fF
C9657 col_n[26] col[27] 5.90fF
C9658 row_n[2] ctop 1.65fF
C9659 a_13006_15182# rowon_n[13] 0.14fF
C9660 a_7894_13174# rowoff_n[11] 0.24fF
C9661 col[24] rowoff_n[11] 0.11fF
C9662 a_2966_13174# row_n[11] 0.16fF
C9663 a_2874_5142# VDD 0.24fF
C9664 a_6982_4138# col_n[4] 0.28fF
C9665 a_28066_5142# rowon_n[3] 0.14fF
C9666 a_2346_6188# a_19942_6146# 0.35fF
C9667 a_2346_2172# col[0] 0.15fF
C9668 a_32082_17190# ctop 3.39fF
C9669 a_2346_15224# col[2] 0.15fF
C9670 a_15926_8154# rowoff_n[6] 0.24fF
C9671 a_1962_4178# col_n[16] 0.13fF
C9672 a_2346_1168# m2_2736_946# 0.20fF
C9673 a_1962_17230# col_n[18] 0.13fF
C9674 a_13006_16186# vcm 0.62fF
C9675 a_21950_17190# rowoff_n[15] 0.24fF
C9676 a_25966_6146# rowoff_n[4] 0.24fF
C9677 a_5978_5142# row_n[3] 0.17fF
C9678 a_1962_3174# a_14010_3134# 0.27fF
C9679 a_16018_9158# VDD 0.52fF
C9680 a_2346_8196# a_32994_8154# 0.35fF
C9681 a_5978_16186# m2_6176_16434# 0.16fF
C9682 a_17022_8154# a_18026_8154# 0.97fF
C9683 a_22042_14178# col[19] 0.29fF
C9684 a_1962_11206# col[9] 0.11fF
C9685 a_23046_1126# vcm 0.12fF
C9686 a_6282_10202# vcm 0.22fF
C9687 col[8] rowoff_n[12] 0.11fF
C9688 a_7986_4138# m2_8184_4386# 0.16fF
C9689 m2_27836_946# ctop 0.18fF
C9690 a_2346_10204# col[29] 0.15fF
C9691 a_1962_5182# a_27062_5142# 0.27fF
C9692 a_29070_13174# VDD 0.52fF
C9693 a_2346_4180# vcm 0.40fF
C9694 a_25054_8154# row_n[6] 0.17fF
C9695 a_19334_14218# vcm 0.22fF
C9696 a_29070_3134# a_29070_2130# 1.00fF
C9697 a_2346_2172# a_22042_2130# 0.19fF
C9698 a_1962_2170# a_20338_2170# 0.14fF
C9699 a_4974_7150# col[2] 0.29fF
C9700 a_8898_16186# VDD 0.23fF
C9701 a_30074_12170# a_31078_12170# 0.97fF
C9702 a_22042_16186# col_n[19] 0.28fF
C9703 a_1962_13214# col_n[9] 0.13fF
C9704 a_32386_18234# vcm 0.22fF
C9705 a_23046_3134# col[20] 0.29fF
C9706 a_18938_1126# VDD 0.39fF
C9707 a_1962_4178# a_33390_4178# 0.14fF
C9708 a_18938_4138# a_19030_4138# 0.26fF
C9709 a_14010_12170# ctop 3.58fF
C9710 a_2966_10162# VDD 0.56fF
C9711 a_1962_7190# col[0] 0.11fF
C9712 a_13006_6146# rowon_n[4] 0.14fF
C9713 a_2346_13216# a_4882_13174# 0.35fF
C9714 a_34090_10162# rowoff_n[8] 0.10fF
C9715 a_2966_4138# row_n[2] 0.16fF
C9716 a_4974_5142# m2_5172_5390# 0.16fF
C9717 a_2346_6188# col[20] 0.15fF
C9718 a_31990_5142# VDD 0.23fF
C9719 m3_25960_18146# VDD 0.25fF
C9720 a_27062_16186# ctop 3.57fF
C9721 a_4974_9158# col_n[2] 0.28fF
C9722 a_2346_15224# a_17934_15182# 0.35fF
C9723 a_7986_15182# vcm 0.62fF
C9724 a_1962_2170# col[27] 0.11fF
C9725 a_10998_8154# VDD 0.52fF
C9726 a_32082_9158# rowon_n[7] 0.14fF
C9727 a_1962_15222# col[29] 0.11fF
C9728 a_15014_8154# a_15014_7150# 1.00fF
C9729 a_31990_8154# a_32082_8154# 0.26fF
C9730 a_23046_5142# col_n[20] 0.28fF
C9731 a_1962_12210# a_12002_12170# 0.27fF
C9732 a_1962_9198# vcm 6.95fF
C9733 a_16018_17190# a_17022_17190# 0.97fF
C9734 a_2346_17232# a_30986_17190# 0.35fF
C9735 m2_4744_946# m3_5880_1078# 0.13fF
C9736 m3_32988_1078# ctop 0.27fF
C9737 a_9994_9158# row_n[7] 0.17fF
C9738 a_2346_18236# col[21] 0.14fF
C9739 a_24050_12170# VDD 0.52fF
C9740 m3_15920_18146# m3_16924_18146# 0.22fF
C9741 a_4882_9158# a_4974_9158# 0.26fF
C9742 a_2346_9200# a_6982_9158# 0.19fF
C9743 a_1962_9198# a_5278_9198# 0.14fF
C9744 rowon_n[15] rowoff_n[15] 20.27fF
C9745 a_31078_4138# vcm 0.62fF
C9746 a_1962_14218# a_25054_14178# 0.27fF
C9747 a_8898_3134# rowoff_n[1] 0.24fF
C9748 m2_1732_5966# m2_2160_6394# 0.16fF
C9749 a_14314_13214# vcm 0.22fF
C9750 a_23958_14178# rowoff_n[12] 0.24fF
C9751 a_2346_2172# col[11] 0.15fF
C9752 a_26058_2130# a_27062_2130# 0.97fF
C9753 a_2346_15224# col[13] 0.15fF
C9754 a_2346_11208# a_20034_11166# 0.19fF
C9755 a_1962_11206# a_18330_11206# 0.14fF
C9756 a_28066_12170# a_28066_11166# 1.00fF
C9757 a_1962_4178# col_n[27] 0.13fF
C9758 a_1962_17230# col_n[29] 0.13fF
C9759 a_29070_12170# row_n[10] 0.17fF
C9760 a_27366_17230# vcm 0.22fF
C9761 a_3878_17190# rowoff_n[15] 0.24fF
C9762 a_1962_18234# col[3] 0.11fF
C9763 a_1962_11206# col[20] 0.11fF
C9764 a_8990_11166# ctop 3.58fF
C9765 a_21038_8154# col[18] 0.29fF
C9766 a_1962_13214# a_31382_13214# 0.14fF
C9767 a_2346_13216# a_33086_13174# 0.19fF
C9768 a_17934_13174# a_18026_13174# 0.26fF
C9769 col[19] rowoff_n[12] 0.11fF
C9770 a_26970_4138# VDD 0.23fF
C9771 a_2346_5184# a_9902_5142# 0.35fF
C9772 a_22042_15182# ctop 3.58fF
C9773 a_17022_10162# rowon_n[8] 0.14fF
C9774 a_6982_9158# rowoff_n[7] 0.10fF
C9775 m2_34864_9982# m2_34864_8978# 0.99fF
C9776 a_10998_15182# rowoff_n[13] 0.10fF
C9777 a_1962_2170# a_3970_2130# 0.27fF
C9778 a_33086_8154# m2_33284_8402# 0.16fF
C9779 a_2346_11208# col[4] 0.15fF
C9780 a_3970_1126# col[1] 0.38fF
C9781 m2_18800_18014# m3_19936_18146# 0.13fF
C9782 a_5978_7150# VDD 0.52fF
C9783 a_17022_7150# rowoff_n[5] 0.10fF
C9784 a_2346_7192# a_22954_7150# 0.35fF
C9785 a_12002_7150# a_13006_7150# 0.97fF
C9786 col[3] rowoff_n[13] 0.11fF
C9787 a_1962_13214# col_n[20] 0.13fF
C9788 a_21038_10162# col_n[18] 0.28fF
C9789 a_14010_17190# a_14010_16186# 1.00fF
C9790 a_30986_17190# a_31078_17190# 0.26fF
C9791 a_27062_5142# rowoff_n[3] 0.10fF
C9792 a_16018_18194# vcm 0.12fF
C9793 a_1962_4178# a_17022_4138# 0.27fF
C9794 a_1962_7190# col[11] 0.11fF
C9795 a_19030_11166# VDD 0.52fF
C9796 m3_5880_1078# m3_6884_1078# 0.22fF
C9797 m2_9764_18014# col[7] 0.28fF
C9798 a_26058_3134# vcm 0.62fF
C9799 a_2966_17190# col[0] 0.29fF
C9800 a_2346_6188# col[31] 0.15fF
C9801 a_9294_12210# vcm 0.22fF
C9802 m2_1732_946# VDD 1.21fF
C9803 a_1962_1166# a_10298_1166# 0.14fF
C9804 a_14010_13174# row_n[11] 0.17fF
C9805 a_1962_6186# a_30074_6146# 0.27fF
C9806 a_32082_15182# VDD 0.52fF
C9807 m2_1732_6970# rowon_n[5] 0.11fF
C9808 a_25054_11166# a_26058_11166# 0.97fF
C9809 a_3970_3134# col_n[1] 0.28fF
C9810 a_29070_3134# row_n[1] 0.17fF
C9811 a_22346_16226# vcm 0.22fF
C9812 a_2346_3176# a_25054_3134# 0.19fF
C9813 a_30074_9158# m2_30272_9406# 0.16fF
C9814 a_13918_3134# a_14010_3134# 0.26fF
C9815 a_1962_3174# a_23350_3174# 0.14fF
C9816 a_3970_10162# ctop 3.57fF
C9817 a_1962_1166# m2_34864_946# 0.17fF
C9818 a_11910_18194# VDD 0.33fF
C9819 a_1962_9198# col_n[11] 0.13fF
C9820 a_32386_1166# vcm 0.23fF
C9821 a_19030_13174# col[16] 0.29fF
C9822 a_25966_11166# rowoff_n[9] 0.24fF
C9823 m2_25828_18014# col_n[23] 0.25fF
C9824 a_33086_16186# row_n[14] 0.17fF
C9825 a_21950_3134# VDD 0.23fF
C9826 a_1962_3174# col[2] 0.11fF
C9827 m3_28972_18146# ctop 0.23fF
C9828 col[1] col[2] 0.20fF
C9829 ctop col[9] 1.98fF
C9830 a_1962_16226# col[4] 0.11fF
C9831 a_17022_14178# ctop 3.58fF
C9832 m2_24824_946# m2_25828_946# 0.96fF
C9833 a_2346_14220# a_7894_14178# 0.35fF
C9834 a_2346_2172# col[22] 0.15fF
C9835 a_2346_18236# a_16930_18194# 0.35fF
C9836 a_2346_15224# col[24] 0.15fF
C9837 a_35002_7150# VDD 0.29fF
C9838 a_9994_7150# a_9994_6146# 1.00fF
C9839 a_26970_7150# a_27062_7150# 0.26fF
C9840 a_21038_14178# rowon_n[12] 0.14fF
C9841 a_10998_16186# a_12002_16186# 0.97fF
C9842 a_2346_16228# a_20946_16186# 0.35fF
C9843 a_1962_18234# col[14] 0.11fF
C9844 a_1962_11206# col[31] 0.11fF
C9845 a_10998_17190# vcm 0.60fF
C9846 a_19030_15182# col_n[16] 0.28fF
C9847 a_1962_18234# m2_4744_18014# 0.18fF
C9848 a_27062_10162# m2_27260_10410# 0.16fF
C9849 a_14010_10162# VDD 0.52fF
C9850 a_20034_2130# col[17] 0.29fF
C9851 col[30] rowoff_n[12] 0.11fF
C9852 a_1962_5182# col_n[2] 0.13fF
C9853 a_21038_2130# vcm 0.62fF
C9854 a_1962_13214# a_15014_13174# 0.27fF
C9855 m2_1732_10986# sample 0.19fF
C9856 a_13006_12170# rowoff_n[10] 0.10fF
C9857 a_14010_4138# row_n[2] 0.17fF
C9858 m2_34864_4962# ctop 0.17fF
C9859 a_4274_11206# vcm 0.22fF
C9860 m3_1864_1078# VDD 0.23fF
C9861 a_27062_14178# VDD 0.52fF
C9862 a_23046_11166# a_23046_10162# 1.00fF
C9863 a_1962_10202# a_8290_10202# 0.14fF
C9864 a_2346_10204# a_9994_10162# 0.19fF
C9865 a_9994_2130# rowoff_n[0] 0.10fF
C9866 a_34090_6146# vcm 0.62fF
C9867 a_1962_15222# a_28066_15182# 0.27fF
C9868 a_2346_11208# col[15] 0.15fF
C9869 m2_26832_18014# ctop 0.18fF
C9870 a_17326_15222# vcm 0.22fF
C9871 a_27062_16186# rowoff_n[14] 0.10fF
C9872 a_18026_17190# row_n[15] 0.17fF
C9873 col[14] rowoff_n[13] 0.11fF
C9874 a_1962_13214# col_n[31] 0.13fF
C9875 a_2966_7150# a_3970_7150# 0.97fF
C9876 a_2966_10162# m3_1864_10114# 0.14fF
C9877 a_6890_17190# VDD 0.24fF
C9878 sample_n rowoff_n[9] 0.38fF
C9879 VDD rowoff_n[8] 1.17fF
C9880 a_12914_12170# a_13006_12170# 0.26fF
C9881 a_2346_12212# a_23046_12170# 0.19fF
C9882 a_1962_12210# a_21342_12210# 0.14fF
C9883 a_33086_7150# row_n[5] 0.17fF
C9884 a_20034_4138# col_n[17] 0.28fF
C9885 m2_14784_946# m3_14916_1078# 2.79fF
C9886 m2_22816_946# VDD 0.62fF
C9887 a_1962_7190# col[22] 0.11fF
C9888 a_16930_2130# VDD 0.23fF
C9889 a_24050_11166# m2_24248_11414# 0.16fF
C9890 a_12002_13174# ctop 3.58fF
C9891 m2_25828_946# m3_26964_1078# 0.13fF
C9892 m3_34996_17142# m3_34996_16138# 0.22fF
C9893 a_1962_14218# a_35398_14218# 0.14fF
C9894 a_2346_14220# a_2346_13216# 0.22fF
C9895 a_5978_15182# rowon_n[13] 0.14fF
C9896 a_29982_6146# VDD 0.23fF
C9897 a_21038_5142# rowon_n[3] 0.14fF
C9898 a_2346_6188# a_12914_6146# 0.35fF
C9899 a_6982_6146# a_7986_6146# 0.97fF
C9900 a_25054_17190# ctop 3.39fF
C9901 a_8898_8154# rowoff_n[6] 0.24fF
C9902 a_2346_7192# col[6] 0.15fF
C9903 a_8990_16186# a_8990_15182# 1.00fF
C9904 a_25966_16186# a_26058_16186# 0.26fF
C9905 a_31078_2130# m2_31276_2378# 0.16fF
C9906 a_14922_17190# rowoff_n[15] 0.24fF
C9907 a_5978_16186# vcm 0.62fF
C9908 a_1962_3174# a_6982_3134# 0.27fF
C9909 a_18938_6146# rowoff_n[4] 0.24fF
C9910 a_8990_9158# VDD 0.52fF
C9911 a_1962_9198# col_n[22] 0.13fF
C9912 a_2346_8196# a_25966_8154# 0.35fF
C9913 a_16018_1126# vcm 0.12fF
C9914 a_18026_7150# col[15] 0.29fF
C9915 a_1962_3174# col[13] 0.11fF
C9916 a_28978_4138# rowoff_n[2] 0.24fF
C9917 VDD sample 5.62fF
C9918 ctop col[20] 1.98fF
C9919 a_1962_16226# col[15] 0.11fF
C9920 a_1962_4178# m2_1732_3958# 0.15fF
C9921 a_3878_3134# VDD 0.23fF
C9922 a_21038_12170# m2_21236_12418# 0.16fF
C9923 a_1962_5182# a_20034_5142# 0.27fF
C9924 a_22042_13174# VDD 0.52fF
C9925 a_20034_10162# a_21038_10162# 0.97fF
C9926 a_29070_5142# vcm 0.62fF
C9927 a_18026_8154# row_n[6] 0.17fF
C9928 a_12306_14218# vcm 0.22fF
C9929 a_1962_2170# a_13310_2170# 0.14fF
C9930 a_2346_2172# a_15014_2130# 0.19fF
C9931 a_8898_2130# a_8990_2130# 0.26fF
C9932 m2_33860_18014# m3_32988_18146# 0.13fF
C9933 a_1962_7190# a_33086_7150# 0.27fF
C9934 a_2966_14178# rowon_n[12] 0.13fF
C9935 a_1962_18234# col[25] 0.11fF
C9936 a_2346_16228# a_1962_16226# 2.62fF
C9937 m2_12776_946# col_n[10] 0.37fF
C9938 a_25358_18234# vcm 0.22fF
C9939 a_18026_9158# col_n[15] 0.28fF
C9940 a_11910_1126# VDD 0.44fF
C9941 a_1962_4178# a_26362_4178# 0.14fF
C9942 a_2346_4180# a_28066_4138# 0.19fF
C9943 a_32082_5142# a_32082_4138# 1.00fF
C9944 a_1962_5182# col_n[13] 0.13fF
C9945 a_6982_12170# ctop 3.58fF
C9946 a_5978_6146# rowon_n[4] 0.14fF
C9947 m2_16792_946# VDD 0.61fF
C9948 a_2966_2130# vcm 0.12fF
C9949 a_33086_14178# a_34090_14178# 0.97fF
C9950 a_27062_10162# rowoff_n[8] 0.10fF
C9951 a_1962_12210# col[6] 0.11fF
C9952 a_29070_13174# rowoff_n[11] 0.10fF
C9953 a_24962_5142# VDD 0.23fF
C9954 m2_33860_946# VDD 0.51fF
C9955 a_4974_6146# a_4974_5142# 1.00fF
C9956 a_21950_6146# a_22042_6146# 0.26fF
C9957 a_18026_13174# m2_18224_13422# 0.16fF
C9958 a_20034_16186# ctop 3.57fF
C9959 a_2346_11208# col[26] 0.15fF
C9960 a_2346_15224# a_10906_15182# 0.35fF
C9961 a_5978_15182# a_6982_15182# 0.97fF
C9962 col[25] rowoff_n[13] 0.11fF
C9963 a_1962_3174# a_34394_3174# 0.14fF
C9964 a_24050_2130# m3_23952_1078# 0.15fF
C9965 vcm rowoff_n[1] 0.20fF
C9966 a_3970_8154# VDD 0.52fF
C9967 a_25054_9158# rowon_n[7] 0.14fF
C9968 a_1962_12210# a_4974_12170# 0.27fF
C9969 a_1962_18234# a_28370_18234# 0.14fF
C9970 a_3878_12170# a_3970_12170# 0.26fF
C9971 a_2346_17232# a_23958_17190# 0.35fF
C9972 m2_30848_18014# m2_31852_18014# 0.96fF
C9973 a_16018_12170# col[13] 0.29fF
C9974 a_1962_1166# col_n[4] 0.13fF
C9975 m3_4876_1078# ctop 0.23fF
C9976 a_1962_14218# col_n[6] 0.13fF
C9977 a_17022_12170# VDD 0.52fF
C9978 m3_1864_18146# m3_2868_18146# 0.22fF
C9979 a_18026_10162# a_18026_9158# 1.00fF
C9980 a_24050_4138# vcm 0.62fF
C9981 a_1962_14218# a_18026_14178# 0.27fF
C9982 col[9] rowoff_n[14] 0.11fF
C9983 a_34090_8154# col[31] 0.29fF
C9984 a_7286_13214# vcm 0.22fF
C9985 a_16930_14178# rowoff_n[12] 0.24fF
C9986 a_2966_5142# rowon_n[3] 0.13fF
C9987 a_15014_14178# m2_15212_14426# 0.16fF
C9988 a_30074_16186# VDD 0.52fF
C9989 a_2346_7192# col[17] 0.15fF
C9990 a_2346_11208# a_13006_11166# 0.19fF
C9991 a_1962_11206# a_11302_11206# 0.14fF
C9992 a_7894_11166# a_7986_11166# 0.26fF
C9993 a_1962_16226# a_31078_16186# 0.27fF
C9994 a_22042_12170# row_n[10] 0.17fF
C9995 a_20338_17230# vcm 0.22fF
C9996 a_29070_4138# a_30074_4138# 0.97fF
C9997 a_16018_14178# col_n[13] 0.28fF
C9998 a_1962_3174# col[24] 0.11fF
C9999 a_1962_13214# a_24354_13214# 0.14fF
C10000 a_31078_14178# a_31078_13174# 1.00fF
C10001 a_2346_13216# a_26058_13174# 0.19fF
C10002 a_30378_2170# vcm 0.22fF
C10003 VDD col_n[9] 4.94fF
C10004 vcm col_n[5] 2.80fF
C10005 col_n[2] col_n[3] 0.10fF
C10006 ctop col[31] 2.13fF
C10007 col[12] col[13] 0.20fF
C10008 a_1962_16226# col[26] 0.11fF
C10009 a_19942_4138# VDD 0.23fF
C10010 a_34090_10162# col_n[31] 0.28fF
C10011 a_15014_15182# ctop 3.58fF
C10012 a_9994_10162# rowon_n[8] 0.14fF
C10013 a_20946_15182# a_21038_15182# 0.26fF
C10014 a_3970_15182# a_3970_14178# 1.00fF
C10015 a_3970_15182# rowoff_n[13] 0.10fF
C10016 m2_34864_10986# VDD 1.01fF
C10017 m2_9764_18014# m3_9896_18146# 2.78fF
C10018 a_20034_1126# m3_19936_1078# 2.44fF
C10019 a_32994_8154# VDD 0.23fF
C10020 a_9994_7150# rowoff_n[5] 0.10fF
C10021 a_12002_15182# m2_12200_15430# 0.16fF
C10022 a_2346_7192# a_15926_7150# 0.35fF
C10023 a_2346_3176# col[8] 0.15fF
C10024 a_2346_16228# col[10] 0.15fF
C10025 a_1962_5182# col_n[24] 0.13fF
C10026 a_14010_3134# m2_14208_3382# 0.16fF
C10027 a_20034_5142# rowoff_n[3] 0.10fF
C10028 a_8990_18194# vcm 0.12fF
C10029 a_17022_3134# col_n[14] 0.28fF
C10030 a_1962_4178# a_9994_4138# 0.27fF
C10031 a_29070_13174# rowon_n[11] 0.14fF
C10032 a_12002_11166# VDD 0.52fF
C10033 a_15014_9158# a_16018_9158# 0.97fF
C10034 a_2346_9200# a_28978_9158# 0.35fF
C10035 a_14010_17190# col[11] 0.29fF
C10036 a_1962_12210# col[17] 0.11fF
C10037 a_19030_3134# vcm 0.62fF
C10038 a_30074_3134# rowoff_n[1] 0.10fF
C10039 m2_1732_7974# ctop 0.17fF
C10040 a_1962_1166# a_3270_1166# 0.14fF
C10041 a_6982_13174# row_n[11] 0.17fF
C10042 a_32082_13174# col[29] 0.29fF
C10043 a_1962_6186# a_23046_6146# 0.27fF
C10044 a_25054_15182# VDD 0.52fF
C10045 a_22042_3134# row_n[1] 0.17fF
C10046 a_32082_7150# vcm 0.62fF
C10047 a_2346_1168# m2_10768_946# 0.19fF
C10048 a_15318_16226# vcm 0.22fF
C10049 a_2346_3176# a_18026_3134# 0.19fF
C10050 a_27062_4138# a_27062_3134# 1.00fF
C10051 a_1962_3174# a_16322_3174# 0.14fF
C10052 a_31078_2130# m2_30848_946# 0.99fF
C10053 a_2346_16228# m2_34864_16006# 0.17fF
C10054 a_8990_16186# m2_9188_16434# 0.16fF
C10055 a_2346_12212# col[1] 0.15fF
C10056 a_4882_18194# VDD 0.33fF
C10057 a_25358_1166# vcm 0.23fF
C10058 a_28066_13174# a_29070_13174# 0.97fF
C10059 m2_7756_946# m2_8760_946# 0.96fF
C10060 a_18938_11166# rowoff_n[9] 0.24fF
C10061 a_1962_1166# col_n[15] 0.12fF
C10062 a_26058_16186# row_n[14] 0.17fF
C10063 a_1962_14218# col_n[17] 0.13fF
C10064 a_10998_4138# m2_11196_4386# 0.16fF
C10065 a_15014_6146# col[12] 0.29fF
C10066 a_14922_3134# VDD 0.23fF
C10067 a_1962_5182# a_29374_5182# 0.14fF
C10068 a_16930_5142# a_17022_5142# 0.26fF
C10069 a_2346_5184# a_31078_5142# 0.19fF
C10070 a_9994_14178# ctop 3.58fF
C10071 col[20] rowoff_n[14] 0.11fF
C10072 a_1962_8194# col[8] 0.11fF
C10073 a_28978_9158# rowoff_n[7] 0.24fF
C10074 a_32082_15182# col_n[29] 0.28fF
C10075 a_33086_2130# col[30] 0.29fF
C10076 a_2346_18236# a_9902_18194# 0.35fF
C10077 a_32994_15182# rowoff_n[13] 0.24fF
C10078 m2_1732_16006# m3_1864_17142# 0.15fF
C10079 a_2346_7192# col[28] 0.15fF
C10080 a_27974_7150# VDD 0.23fF
C10081 a_14010_14178# rowon_n[12] 0.14fF
C10082 a_2346_16228# a_13918_16186# 0.35fF
C10083 a_1962_2170# m2_2736_1950# 0.18fF
C10084 a_29070_4138# rowon_n[2] 0.14fF
C10085 a_33086_3134# ctop 3.56fF
C10086 a_3970_17190# vcm 0.60fF
C10087 a_34090_4138# m3_34996_4090# 0.13fF
C10088 a_6982_10162# VDD 0.52fF
C10089 VDD col_n[20] 4.99fF
C10090 vcm col_n[16] 2.79fF
C10091 col[4] rowoff_n[15] 0.11fF
C10092 a_15014_8154# col_n[12] 0.28fF
C10093 a_5978_17190# m2_6176_17438# 0.16fF
C10094 a_13006_9158# a_13006_8154# 1.00fF
C10095 a_29982_9158# a_30074_9158# 0.26fF
C10096 a_14010_2130# vcm 0.62fF
C10097 a_1962_13214# a_7986_13174# 0.27fF
C10098 a_6982_4138# row_n[2] 0.17fF
C10099 a_5978_12170# rowoff_n[10] 0.10fF
C10100 a_1962_10202# col_n[8] 0.13fF
C10101 a_7986_5142# m2_8184_5390# 0.16fF
C10102 a_2346_1168# a_35002_1126# 0.35fF
C10103 a_35494_5504# VDD 0.11fF
C10104 a_33086_4138# col_n[30] 0.28fF
C10105 m3_34996_15134# VDD 0.26fF
C10106 a_33086_17190# rowon_n[15] 0.14fF
C10107 a_20034_14178# VDD 0.52fF
C10108 a_2346_10204# a_2874_10162# 0.35fF
C10109 a_2874_2130# rowoff_n[0] 0.24fF
C10110 a_1962_17230# col[1] 0.11fF
C10111 a_1962_15222# a_21038_15182# 0.27fF
C10112 a_27062_6146# vcm 0.62fF
C10113 a_10298_15222# vcm 0.22fF
C10114 a_20034_16186# rowoff_n[14] 0.10fF
C10115 m2_12776_18014# ctop 0.18fF
C10116 a_24050_3134# a_25054_3134# 0.97fF
C10117 m2_2736_946# col[0] 0.39fF
C10118 a_2346_3176# col[19] 0.15fF
C10119 a_27974_1126# m2_27836_946# 0.16fF
C10120 a_10998_17190# row_n[15] 0.17fF
C10121 a_2346_16228# col[21] 0.15fF
C10122 a_1962_12210# a_14314_12210# 0.14fF
C10123 a_26058_13174# a_26058_12170# 1.00fF
C10124 a_2346_12212# a_16018_12170# 0.19fF
C10125 a_26058_7150# row_n[5] 0.17fF
C10126 a_1962_17230# a_34090_17190# 0.27fF
C10127 m2_9764_946# m3_10900_1078# 0.13fF
C10128 a_9902_2130# VDD 0.23fF
C10129 a_4974_13174# ctop 3.58fF
C10130 a_1962_12210# col[28] 0.11fF
C10131 a_13006_11166# col[10] 0.29fF
C10132 a_33390_4178# vcm 0.22fF
C10133 a_1962_14218# a_27366_14218# 0.14fF
C10134 a_2346_14220# a_29070_14178# 0.19fF
C10135 a_15926_14178# a_16018_14178# 0.26fF
C10136 a_1962_6186# col_n[0] 0.13fF
C10137 a_4974_6146# m2_5172_6394# 0.16fF
C10138 m2_1732_12994# m3_1864_14130# 0.15fF
C10139 a_31078_7150# col[28] 0.29fF
C10140 a_22954_6146# VDD 0.23fF
C10141 a_14010_5142# rowon_n[3] 0.14fF
C10142 a_2346_6188# a_5886_6146# 0.35fF
C10143 a_18026_17190# ctop 3.39fF
C10144 m2_1732_12994# m2_1732_11990# 0.99fF
C10145 a_7894_17190# rowoff_n[15] 0.24fF
C10146 a_28066_2130# ctop 3.39fF
C10147 m2_32856_18014# VDD 0.91fF
C10148 a_11910_6146# rowoff_n[4] 0.24fF
C10149 a_2346_12212# col[12] 0.15fF
C10150 a_2346_8196# a_18938_8154# 0.35fF
C10151 a_9994_8154# a_10998_8154# 0.97fF
C10152 a_1962_1166# col_n[26] 0.13fF
C10153 a_8990_1126# vcm 0.12fF
C10154 a_1962_14218# col_n[28] 0.13fF
C10155 a_13006_13174# col_n[10] 0.28fF
C10156 a_35002_12170# rowoff_n[10] 0.24fF
C10157 a_21950_4138# rowoff_n[2] 0.24fF
C10158 a_33086_8154# rowon_n[6] 0.14fF
C10159 m2_11772_946# vcm 0.42fF
C10160 a_1962_5182# a_13006_5142# 0.27fF
C10161 a_1962_8194# col[19] 0.11fF
C10162 col[31] rowoff_n[14] 0.11fF
C10163 a_15014_13174# VDD 0.52fF
C10164 a_2346_10204# a_31990_10162# 0.35fF
C10165 a_31990_2130# rowoff_n[0] 0.24fF
C10166 a_31078_9158# col_n[28] 0.28fF
C10167 a_22042_5142# vcm 0.62fF
C10168 m2_28840_946# vcm 0.42fF
C10169 a_10998_8154# row_n[6] 0.17fF
C10170 a_5278_14218# vcm 0.22fF
C10171 a_2346_2172# a_7986_2130# 0.19fF
C10172 a_22042_3134# a_22042_2130# 1.00fF
C10173 a_1962_2170# a_6282_2170# 0.14fF
C10174 m2_23820_18014# m3_24956_18146# 0.13fF
C10175 a_1962_7190# a_26058_7150# 0.27fF
C10176 a_28066_17190# VDD 0.55fF
C10177 a_23046_12170# a_24050_12170# 0.97fF
C10178 a_35094_9158# vcm 0.12fF
C10179 a_18330_18234# vcm 0.22fF
C10180 vcm col_n[27] 2.80fF
C10181 col_n[13] col_n[14] 0.10fF
C10182 VDD col_n[31] 5.07fF
C10183 a_4882_1126# VDD 0.44fF
C10184 col[15] rowoff_n[15] 0.11fF
C10185 a_2346_8196# col[3] 0.15fF
C10186 col[23] col[24] 0.20fF
C10187 a_11910_4138# a_12002_4138# 0.26fF
C10188 a_1962_4178# a_19334_4178# 0.14fF
C10189 a_2346_4180# a_21038_4138# 0.19fF
C10190 a_14010_2130# col_n[11] 0.28fF
C10191 a_4974_17190# m2_4744_18014# 1.00fF
C10192 a_28370_3174# vcm 0.22fF
C10193 a_30074_11166# row_n[9] 0.17fF
C10194 a_1962_10202# col_n[19] 0.13fF
C10195 a_20034_10162# rowoff_n[8] 0.10fF
C10196 a_10998_16186# col[8] 0.29fF
C10197 a_22042_13174# rowoff_n[11] 0.10fF
C10198 m2_9764_946# VDD 0.62fF
C10199 m2_1732_9982# m3_1864_11118# 0.15fF
C10200 a_17934_5142# VDD 0.23fF
C10201 a_1962_4178# col[10] 0.11fF
C10202 a_2346_6188# a_34090_6146# 0.19fF
C10203 a_1962_6186# a_32386_6186# 0.14fF
C10204 a_1962_17230# col[12] 0.11fF
C10205 a_13006_16186# ctop 3.57fF
C10206 a_30074_8154# rowoff_n[6] 0.10fF
C10207 a_29070_12170# col[26] 0.29fF
C10208 a_1962_15222# a_2966_15182# 0.27fF
C10209 m2_1732_2954# sample_n 0.15fF
C10210 a_2346_3176# col[30] 0.15fF
C10211 m2_1732_13998# VDD 1.02fF
C10212 m2_11772_946# m2_12200_1374# 0.16fF
C10213 a_33086_9158# m2_33284_9406# 0.16fF
C10214 a_30986_9158# VDD 0.23fF
C10215 a_18026_9158# rowon_n[7] 0.14fF
C10216 a_7986_8154# a_7986_7150# 1.00fF
C10217 a_24962_8154# a_25054_8154# 0.26fF
C10218 a_1962_18234# a_21342_18234# 0.14fF
C10219 a_2346_17232# a_16930_17190# 0.35fF
C10220 a_8990_17190# a_9994_17190# 0.97fF
C10221 m2_23820_18014# m2_24824_18014# 0.96fF
C10222 a_2346_4180# ctop 1.59fF
C10223 m3_1864_13126# ctop 0.23fF
C10224 a_12002_5142# col[9] 0.29fF
C10225 a_9994_12170# VDD 0.52fF
C10226 m2_28840_946# m2_29268_1374# 0.16fF
C10227 a_1962_6186# col_n[10] 0.13fF
C10228 a_1962_14218# a_10998_14178# 0.27fF
C10229 a_17022_4138# vcm 0.62fF
C10230 m2_1732_18014# sample 0.16fF
C10231 a_29070_14178# col_n[26] 0.28fF
C10232 a_9902_14178# rowoff_n[12] 0.24fF
C10233 a_19030_2130# a_20034_2130# 0.97fF
C10234 a_1962_2170# a_1962_1166# 0.15fF
C10235 a_2966_16186# col_n[0] 0.28fF
C10236 m2_3740_18014# col[1] 0.28fF
C10237 a_1962_13214# col[3] 0.11fF
C10238 a_23046_16186# VDD 0.52fF
C10239 a_2346_11208# a_5978_11166# 0.19fF
C10240 a_1962_11206# a_4274_11206# 0.14fF
C10241 a_21038_12170# a_21038_11166# 1.00fF
C10242 a_30074_8154# vcm 0.62fF
C10243 a_1962_16226# a_24050_16186# 0.27fF
C10244 a_2346_12212# col[23] 0.15fF
C10245 a_15014_12170# row_n[10] 0.17fF
C10246 a_13310_17230# vcm 0.22fF
C10247 a_30074_10162# m2_30272_10410# 0.16fF
C10248 a_30074_2130# row_n[0] 0.17fF
C10249 a_24050_17190# m2_23820_18014# 1.00fF
C10250 a_1962_14218# row_n[12] 25.57fF
C10251 a_34090_13174# m3_34996_13126# 0.13fF
C10252 a_23350_2170# vcm 0.22fF
C10253 a_10906_13174# a_10998_13174# 0.26fF
C10254 a_2346_13216# a_19030_13174# 0.19fF
C10255 a_1962_13214# a_17326_13214# 0.14fF
C10256 a_12002_7150# col_n[9] 0.28fF
C10257 a_3878_4138# rowoff_n[2] 0.24fF
C10258 a_1962_8194# col[30] 0.11fF
C10259 m2_1732_6970# m3_1864_8106# 0.15fF
C10260 a_12914_4138# VDD 0.23fF
C10261 m3_16924_1078# VDD 0.14fF
C10262 a_32082_6146# a_33086_6146# 0.97fF
C10263 a_7986_15182# ctop 3.58fF
C10264 a_1962_2170# col_n[1] 0.13fF
C10265 a_30074_3134# col_n[27] 0.28fF
C10266 m2_19804_18014# col_n[17] 0.25fF
C10267 a_1962_15222# col_n[3] 0.13fF
C10268 a_34090_15182# row_n[13] 0.17fF
C10269 a_2346_15224# a_32082_15182# 0.19fF
C10270 a_1962_15222# a_30378_15222# 0.14fF
C10271 a_34090_16186# a_34090_15182# 1.00fF
C10272 a_27062_17190# col[24] 0.29fF
C10273 a_1962_9198# ctop 1.49fF
C10274 a_25966_8154# VDD 0.23fF
C10275 a_2874_7150# rowoff_n[5] 0.24fF
C10276 a_2346_7192# a_8898_7150# 0.35fF
C10277 a_4974_7150# a_5978_7150# 0.97fF
C10278 m2_20808_946# m3_20940_1078# 2.79fF
C10279 col_n[1] row_n[13] 0.23fF
C10280 VDD rowon_n[10] 2.61fF
C10281 vcm rowon_n[12] 0.50fF
C10282 col_n[3] row_n[14] 0.23fF
C10283 col_n[0] row_n[12] 0.23fF
C10284 col_n[5] row_n[15] 0.23fF
C10285 a_6982_17190# a_6982_16186# 1.00fF
C10286 a_23958_17190# a_24050_17190# 0.26fF
C10287 col[26] rowoff_n[15] 0.11fF
C10288 a_2346_8196# col[14] 0.15fF
C10289 a_13006_5142# rowoff_n[3] 0.10fF
C10290 a_31078_4138# ctop 3.58fF
C10291 a_27062_11166# m2_27260_11414# 0.16fF
C10292 a_2346_4180# a_2966_4138# 0.21fF
C10293 a_22042_13174# rowon_n[11] 0.14fF
C10294 a_4974_11166# VDD 0.52fF
C10295 m2_30848_946# m3_31984_1078# 0.13fF
C10296 a_1962_10202# col_n[30] 0.13fF
C10297 a_2346_9200# a_21950_9158# 0.35fF
C10298 a_12002_3134# vcm 0.62fF
C10299 m2_9764_946# col_n[7] 0.37fF
C10300 a_9994_10162# col[7] 0.29fF
C10301 a_23046_3134# rowoff_n[1] 0.10fF
C10302 a_1962_4178# col[21] 0.11fF
C10303 a_1962_17230# col[23] 0.11fF
C10304 a_33998_2130# a_34090_2130# 0.25fF
C10305 a_1962_6186# a_16018_6146# 0.27fF
C10306 a_18026_15182# VDD 0.52fF
C10307 a_28066_6146# col[25] 0.29fF
C10308 a_18026_11166# a_19030_11166# 0.97fF
C10309 a_2346_11208# a_35002_11166# 0.35fF
C10310 a_15014_3134# row_n[1] 0.17fF
C10311 a_25054_7150# vcm 0.62fF
C10312 a_34090_2130# m2_34288_2378# 0.16fF
C10313 a_8290_16226# vcm 0.22fF
C10314 a_1962_5182# row_n[3] 25.57fF
C10315 a_1962_3174# a_9294_3174# 0.14fF
C10316 a_2346_3176# a_10998_3134# 0.19fF
C10317 a_6890_3134# a_6982_3134# 0.26fF
C10318 a_1962_8194# a_29070_8154# 0.27fF
C10319 a_18330_1166# vcm 0.22fF
C10320 a_2346_4180# col[5] 0.15fF
C10321 a_11910_11166# rowoff_n[9] 0.24fF
C10322 a_2346_17232# col[7] 0.15fF
C10323 a_19030_16186# row_n[14] 0.17fF
C10324 m2_1732_3958# m3_1864_5094# 0.15fF
C10325 a_9994_12170# col_n[7] 0.28fF
C10326 a_7894_3134# VDD 0.23fF
C10327 a_2346_5184# a_24050_5142# 0.19fF
C10328 a_1962_5182# a_22346_5182# 0.14fF
C10329 a_24050_12170# m2_24248_12418# 0.16fF
C10330 a_30074_6146# a_30074_5142# 1.00fF
C10331 a_1962_6186# col_n[21] 0.13fF
C10332 a_34090_6146# row_n[4] 0.17fF
C10333 a_21950_9158# rowoff_n[7] 0.24fF
C10334 a_31382_5182# vcm 0.22fF
C10335 a_31078_15182# a_32082_15182# 0.97fF
C10336 a_28066_8154# col_n[25] 0.28fF
C10337 a_25966_15182# rowoff_n[13] 0.24fF
C10338 a_1962_13214# col[14] 0.11fF
C10339 a_20946_7150# VDD 0.23fF
C10340 a_31990_7150# rowoff_n[5] 0.24fF
C10341 a_19942_7150# a_20034_7150# 0.26fF
C10342 a_6982_14178# rowon_n[12] 0.14fF
C10343 a_3970_16186# a_4974_16186# 0.97fF
C10344 a_2346_16228# a_6890_16186# 0.35fF
C10345 a_22042_4138# rowon_n[2] 0.14fF
C10346 a_26058_3134# ctop 3.57fF
C10347 a_33998_11166# VDD 0.23fF
C10348 m3_34568_1078# m3_34996_1078# 0.21fF
C10349 a_6982_2130# vcm 0.62fF
C10350 a_1962_5182# m2_1732_4962# 0.15fF
C10351 a_2346_1168# a_26970_1126# 0.35fF
C10352 a_7986_15182# col[5] 0.29fF
C10353 m3_12908_18146# VDD 0.24fF
C10354 a_21038_13174# m2_21236_13422# 0.16fF
C10355 a_1962_2170# col_n[12] 0.13fF
C10356 a_26058_17190# rowon_n[15] 0.14fF
C10357 a_1962_15222# col_n[14] 0.13fF
C10358 a_13006_14178# VDD 0.52fF
C10359 m2_1732_3958# vcm 0.45fF
C10360 a_16018_11166# a_16018_10162# 1.00fF
C10361 a_32994_11166# a_33086_11166# 0.26fF
C10362 a_20034_6146# vcm 0.62fF
C10363 a_1962_15222# a_14010_15182# 0.27fF
C10364 a_26058_11166# col[23] 0.29fF
C10365 a_1962_9198# col[5] 0.11fF
C10366 a_3270_15222# vcm 0.22fF
C10367 a_13006_16186# rowoff_n[14] 0.10fF
C10368 a_27062_2130# m3_26964_1078# 0.15fF
C10369 a_3970_17190# row_n[15] 0.17fF
C10370 VDD row_n[5] 2.93fF
C10371 sample row_n[6] 1.03fF
C10372 col_n[8] row_n[11] 0.23fF
C10373 col_n[6] row_n[10] 0.23fF
C10374 vcm row_n[7] 0.49fF
C10375 col_n[24] col_n[25] 0.10fF
C10376 col_n[16] row_n[15] 0.23fF
C10377 col_n[10] row_n[12] 0.23fF
C10378 col_n[14] row_n[14] 0.23fF
C10379 col_n[2] row_n[8] 0.23fF
C10380 col_n[4] row_n[9] 0.23fF
C10381 col_n[12] row_n[13] 0.23fF
C10382 a_2346_8196# col[25] 0.15fF
C10383 m2_27836_18014# vcm 0.28fF
C10384 a_2346_12212# a_8990_12170# 0.19fF
C10385 a_1962_12210# a_7286_12210# 0.14fF
C10386 a_5886_12170# a_5978_12170# 0.26fF
C10387 a_19030_7150# row_n[5] 0.17fF
C10388 a_33086_10162# vcm 0.62fF
C10389 a_1962_17230# a_27062_17190# 0.27fF
C10390 m2_34864_18014# m2_35292_18442# 0.16fF
C10391 a_2346_2172# VDD 32.67fF
C10392 m3_19936_1078# ctop 0.36fF
C10393 a_27062_5142# a_28066_5142# 0.97fF
C10394 a_2874_9158# a_2966_9158# 0.26fF
C10395 a_2346_9200# a_3878_9158# 0.35fF
C10396 a_7986_17190# col_n[5] 0.28fF
C10397 a_26362_4178# vcm 0.22fF
C10398 a_29070_15182# a_29070_14178# 1.00fF
C10399 a_2346_14220# a_22042_14178# 0.19fF
C10400 a_1962_14218# a_20338_14218# 0.14fF
C10401 a_8990_4138# col[6] 0.29fF
C10402 a_15926_6146# VDD 0.23fF
C10403 a_6982_5142# rowon_n[3] 0.14fF
C10404 a_26058_13174# col_n[23] 0.28fF
C10405 a_18026_14178# m2_18224_14426# 0.16fF
C10406 a_1962_11206# col_n[5] 0.13fF
C10407 a_10998_17190# ctop 3.39fF
C10408 a_18938_16186# a_19030_16186# 0.26fF
C10409 a_1962_16226# a_33390_16226# 0.14fF
C10410 a_21038_2130# ctop 3.39fF
C10411 m2_18800_18014# VDD 1.30fF
C10412 a_1962_18234# m2_33860_18014# 0.18fF
C10413 a_4882_6146# rowoff_n[4] 0.24fF
C10414 a_28978_10162# VDD 0.23fF
C10415 a_2346_8196# a_11910_8154# 0.35fF
C10416 a_2346_4180# col[16] 0.15fF
C10417 a_34394_2170# vcm 0.22fF
C10418 a_2346_17232# col[18] 0.15fF
C10419 a_14922_4138# rowoff_n[2] 0.24fF
C10420 a_27974_12170# rowoff_n[10] 0.24fF
C10421 a_26058_8154# rowon_n[6] 0.14fF
C10422 a_8990_6146# col_n[6] 0.28fF
C10423 a_34090_6146# ctop 3.42fF
C10424 a_1962_5182# a_5978_5142# 0.27fF
C10425 a_2346_18236# m2_28840_18014# 0.19fF
C10426 a_7986_13174# VDD 0.52fF
C10427 m2_4744_946# vcm 0.41fF
C10428 a_13006_10162# a_14010_10162# 0.97fF
C10429 a_2346_10204# a_24962_10162# 0.35fF
C10430 a_24962_2130# rowoff_n[0] 0.24fF
C10431 a_3878_9158# rowoff_n[7] 0.24fF
C10432 a_1962_13214# col[25] 0.11fF
C10433 a_15014_5142# vcm 0.62fF
C10434 a_27062_2130# col_n[24] 0.28fF
C10435 a_3970_8154# row_n[6] 0.17fF
C10436 m2_14784_18014# m3_14916_18146# 2.78fF
C10437 a_24050_16186# col[21] 0.29fF
C10438 a_1962_7190# VDD 2.73fF
C10439 a_15014_15182# m2_15212_15430# 0.16fF
C10440 a_1962_7190# a_19030_7150# 0.27fF
C10441 a_21038_17190# VDD 0.55fF
C10442 a_2966_12170# a_2966_11166# 1.00fF
C10443 a_28066_9158# vcm 0.62fF
C10444 a_17022_3134# m2_17220_3382# 0.16fF
C10445 a_11302_18234# vcm 0.22fF
C10446 a_31078_2130# VDD 0.55fF
C10447 a_1962_4178# a_12306_4178# 0.14fF
C10448 a_2346_4180# a_14010_4138# 0.19fF
C10449 a_25054_5142# a_25054_4138# 1.00fF
C10450 a_22954_18194# m2_22816_18014# 0.16fF
C10451 a_1962_9198# a_32082_9158# 0.27fF
C10452 a_2346_13216# col[9] 0.15fF
C10453 a_23046_11166# row_n[9] 0.17fF
C10454 a_21342_3174# vcm 0.22fF
C10455 a_26058_14178# a_27062_14178# 0.97fF
C10456 a_13006_10162# rowoff_n[8] 0.10fF
C10457 a_15014_13174# rowoff_n[11] 0.10fF
C10458 a_1962_2170# col_n[23] 0.13fF
C10459 a_6982_9158# col[4] 0.29fF
C10460 a_1962_15222# col_n[25] 0.13fF
C10461 a_10906_5142# VDD 0.23fF
C10462 a_1962_6186# a_25358_6186# 0.14fF
C10463 a_2346_6188# a_27062_6146# 0.19fF
C10464 a_14922_6146# a_15014_6146# 0.26fF
C10465 a_5978_16186# ctop 3.57fF
C10466 a_23046_8154# rowoff_n[6] 0.10fF
C10467 a_1962_9198# col[16] 0.11fF
C10468 a_35398_7190# vcm 0.23fF
C10469 a_25054_5142# col[22] 0.29fF
C10470 a_29070_17190# rowoff_n[15] 0.10fF
C10471 a_33086_6146# rowoff_n[4] 0.10fF
C10472 a_1962_1166# m2_27836_946# 0.18fF
C10473 col_n[11] row_n[7] 0.23fF
C10474 col_n[9] row_n[6] 0.23fF
C10475 col_n[17] row_n[10] 0.23fF
C10476 col_n[21] row_n[12] 0.23fF
C10477 col_n[3] row_n[3] 0.23fF
C10478 col_n[7] row_n[5] 0.23fF
C10479 col_n[15] row_n[9] 0.23fF
C10480 col_n[23] row_n[13] 0.23fF
C10481 col_n[13] row_n[8] 0.23fF
C10482 col_n[19] row_n[11] 0.23fF
C10483 col_n[1] row_n[2] 0.23fF
C10484 col_n[27] row_n[15] 0.23fF
C10485 vcm rowon_n[1] 0.50fF
C10486 col_n[0] row_n[1] 0.23fF
C10487 col_n[5] row_n[4] 0.23fF
C10488 col_n[25] row_n[14] 0.23fF
C10489 VDD sw 0.22fF
C10490 a_10998_9158# rowon_n[7] 0.14fF
C10491 a_23958_9158# VDD 0.23fF
C10492 a_12002_16186# m2_12200_16434# 0.16fF
C10493 a_1962_18234# a_14314_18234# 0.14fF
C10494 m2_1732_4962# rowoff_n[3] 0.12fF
C10495 a_2346_17232# a_9902_17190# 0.35fF
C10496 m2_16792_18014# m2_17796_18014# 0.96fF
C10497 a_14010_4138# m2_14208_4386# 0.16fF
C10498 a_29070_5142# ctop 3.58fF
C10499 m3_15920_18146# ctop 0.23fF
C10500 a_2874_12170# VDD 0.24fF
C10501 a_6982_11166# col_n[4] 0.28fF
C10502 a_10998_10162# a_10998_9158# 1.00fF
C10503 a_27974_10162# a_28066_10162# 0.26fF
C10504 a_2346_9200# col[0] 0.15fF
C10505 a_9994_4138# vcm 0.62fF
C10506 a_1962_14218# a_3970_14178# 0.27fF
C10507 a_1962_18234# col_n[0] 0.13fF
C10508 a_2346_14220# rowoff_n[12] 4.09fF
C10509 a_30074_12170# rowon_n[10] 0.14fF
C10510 a_1962_11206# col_n[16] 0.13fF
C10511 a_2346_2172# a_29982_2130# 0.35fF
C10512 a_25054_7150# col_n[22] 0.28fF
C10513 a_16018_16186# VDD 0.52fF
C10514 a_1962_5182# col[7] 0.11fF
C10515 a_1962_16226# a_17022_16186# 0.27fF
C10516 a_23046_8154# vcm 0.62fF
C10517 a_7986_12170# row_n[10] 0.17fF
C10518 a_6282_17230# vcm 0.22fF
C10519 a_22042_4138# a_23046_4138# 0.97fF
C10520 a_2346_4180# col[27] 0.15fF
C10521 a_2966_3134# m3_2868_2082# 0.15fF
C10522 a_2346_17232# col[29] 0.15fF
C10523 a_23046_2130# row_n[0] 0.17fF
C10524 a_8990_17190# m2_9188_17438# 0.16fF
C10525 a_2346_17232# m2_34864_17010# 0.17fF
C10526 a_16322_2170# vcm 0.22fF
C10527 a_1962_13214# a_10298_13214# 0.14fF
C10528 a_24050_14178# a_24050_13174# 1.00fF
C10529 a_2346_13216# a_12002_13174# 0.19fF
C10530 a_2346_11208# vcm 0.40fF
C10531 a_10998_5142# m2_11196_5390# 0.16fF
C10532 a_5886_4138# VDD 0.23fF
C10533 m3_1864_7102# VDD 0.25fF
C10534 a_4974_14178# col[2] 0.29fF
C10535 col[0] rowoff_n[7] 0.11fF
C10536 col[2] rowoff_n[9] 0.11fF
C10537 col[1] rowoff_n[8] 0.11fF
C10538 ctop rowoff_n[1] 0.60fF
C10539 a_27062_15182# row_n[13] 0.17fF
C10540 a_29374_6186# vcm 0.22fF
C10541 a_2346_15224# a_25054_15182# 0.19fF
C10542 a_13918_15182# a_14010_15182# 0.26fF
C10543 a_1962_15222# a_23350_15222# 0.14fF
C10544 a_1962_7190# col_n[7] 0.13fF
C10545 a_23046_10162# col[20] 0.29fF
C10546 a_18938_8154# VDD 0.23fF
C10547 a_2966_17190# VDD 0.60fF
C10548 a_1962_14218# col[0] 0.11fF
C10549 a_2966_3134# m2_1732_2954# 0.96fF
C10550 a_5978_5142# rowoff_n[3] 0.10fF
C10551 a_24050_4138# ctop 3.58fF
C10552 a_2346_13216# col[20] 0.15fF
C10553 a_15014_13174# rowon_n[11] 0.14fF
C10554 a_31990_12170# VDD 0.23fF
C10555 m3_30980_18146# m3_31984_18146# 0.22fF
C10556 a_7986_9158# a_8990_9158# 0.97fF
C10557 a_2346_9200# a_14922_9158# 0.35fF
C10558 m2_34864_11990# row_n[10] 0.15fF
C10559 a_4974_3134# vcm 0.62fF
C10560 a_30074_3134# rowon_n[1] 0.14fF
C10561 a_16018_3134# rowoff_n[1] 0.10fF
C10562 a_4974_16186# col_n[2] 0.28fF
C10563 a_1962_15222# rowon_n[13] 1.18fF
C10564 a_31078_14178# rowoff_n[12] 0.10fF
C10565 a_5978_3134# col[3] 0.29fF
C10566 a_7986_6146# m2_8184_6394# 0.16fF
C10567 a_1962_6186# a_8990_6146# 0.27fF
C10568 m2_32856_946# col_n[30] 0.45fF
C10569 a_1962_9198# col[27] 0.11fF
C10570 a_10998_15182# VDD 0.52fF
C10571 a_2346_11208# a_27974_11166# 0.35fF
C10572 a_23046_12170# col_n[20] 0.28fF
C10573 m2_15788_946# a_16018_2130# 0.99fF
C10574 a_7986_3134# row_n[1] 0.17fF
C10575 a_3970_17190# m3_3872_18146# 0.15fF
C10576 a_18026_7150# vcm 0.62fF
C10577 a_1962_3174# sample 0.14fF
C10578 col_n[30] row_n[11] 0.23fF
C10579 col_n[8] row_n[0] 0.23fF
C10580 col_n[14] row_n[3] 0.23fF
C10581 col_n[22] row_n[7] 0.23fF
C10582 col_n[24] row_n[8] 0.23fF
C10583 col_n[12] row_n[2] 0.23fF
C10584 col_n[20] row_n[6] 0.23fF
C10585 VDD col[3] 4.17fF
C10586 col_n[0] col[0] 0.72fF
C10587 col_n[5] ctop 2.02fF
C10588 col_n[10] row_n[1] 0.23fF
C10589 col_n[16] row_n[4] 0.23fF
C10590 col_n[26] row_n[9] 0.23fF
C10591 col_n[28] row_n[10] 0.23fF
C10592 col_n[18] row_n[5] 0.23fF
C10593 a_1962_16226# vcm 6.95fF
C10594 a_34090_16186# rowon_n[14] 0.14fF
C10595 a_20034_4138# a_20034_3134# 1.00fF
C10596 a_2346_3176# a_3970_3134# 0.19fF
C10597 a_1962_8194# a_22042_8154# 0.27fF
C10598 a_11302_1166# vcm 0.23fF
C10599 a_21038_13174# a_22042_13174# 0.97fF
C10600 a_31078_11166# vcm 0.62fF
C10601 a_4882_11166# rowoff_n[9] 0.24fF
C10602 a_12002_16186# row_n[14] 0.17fF
C10603 a_34090_4138# VDD 0.54fF
C10604 m2_20808_946# vcm 0.41fF
C10605 a_2346_9200# col[11] 0.15fF
C10606 a_1962_5182# a_15318_5182# 0.14fF
C10607 a_2346_5184# a_17022_5142# 0.19fF
C10608 a_9902_5142# a_9994_5142# 0.26fF
C10609 a_5978_5142# col_n[3] 0.28fF
C10610 a_27062_6146# row_n[4] 0.17fF
C10611 a_14922_9158# rowoff_n[7] 0.24fF
C10612 a_1962_18234# col_n[10] 0.13fF
C10613 a_24354_5182# vcm 0.22fF
C10614 a_1962_11206# col_n[27] 0.13fF
C10615 a_18938_15182# rowoff_n[13] 0.24fF
C10616 a_4974_7150# m2_5172_7398# 0.16fF
C10617 m2_28840_18014# m3_29976_18146# 0.13fF
C10618 a_13918_7150# VDD 0.23fF
C10619 a_24962_7150# rowoff_n[5] 0.24fF
C10620 a_1962_5182# col[18] 0.11fF
C10621 a_1962_7190# a_28370_7190# 0.14fF
C10622 a_33086_8154# a_33086_7150# 1.00fF
C10623 a_2346_7192# a_30074_7150# 0.19fF
C10624 a_2346_10204# row_n[8] 0.35fF
C10625 a_21038_15182# col[18] 0.29fF
C10626 a_35002_5142# rowoff_n[3] 0.24fF
C10627 a_15014_4138# rowon_n[2] 0.14fF
C10628 a_19030_3134# ctop 3.58fF
C10629 a_26970_11166# VDD 0.23fF
C10630 m3_20940_1078# m3_21944_1078# 0.22fF
C10631 a_22954_9158# a_23046_9158# 0.26fF
C10632 a_5978_9158# a_5978_8154# 1.00fF
C10633 a_1962_6186# rowon_n[4] 1.18fF
C10634 m2_1732_3958# m2_2160_4386# 0.16fF
C10635 a_2346_1168# a_19942_1126# 0.39fF
C10636 a_32082_7150# ctop 3.58fF
C10637 a_2346_5184# col[2] 0.15fF
C10638 a_19030_17190# rowon_n[15] 0.14fF
C10639 a_3970_8154# col[1] 0.29fF
C10640 col[12] rowoff_n[8] 0.11fF
C10641 col[11] rowoff_n[7] 0.11fF
C10642 col[6] rowoff_n[2] 0.11fF
C10643 col[5] rowoff_n[1] 0.11fF
C10644 col[10] rowoff_n[6] 0.11fF
C10645 col[9] rowoff_n[5] 0.11fF
C10646 col[13] rowoff_n[9] 0.11fF
C10647 col[8] rowoff_n[4] 0.11fF
C10648 col[7] rowoff_n[3] 0.11fF
C10649 col[4] rowoff_n[0] 0.11fF
C10650 a_5978_14178# VDD 0.52fF
C10651 m2_12776_946# a_12914_1126# 0.16fF
C10652 a_1962_7190# col_n[18] 0.13fF
C10653 a_34090_7150# rowon_n[5] 0.14fF
C10654 a_13006_6146# vcm 0.62fF
C10655 a_1962_15222# a_6982_15182# 0.27fF
C10656 a_21038_17190# col_n[18] 0.28fF
C10657 a_5978_16186# rowoff_n[14] 0.10fF
C10658 a_17022_3134# a_18026_3134# 0.97fF
C10659 a_2346_3176# a_32994_3134# 0.35fF
C10660 a_22042_4138# col[19] 0.29fF
C10661 a_1962_1166# col[9] 0.11fF
C10662 a_1962_14218# col[11] 0.11fF
C10663 m2_13780_18014# vcm 0.28fF
C10664 a_19030_13174# a_19030_12170# 1.00fF
C10665 a_12002_7150# row_n[5] 0.17fF
C10666 a_26058_10162# vcm 0.62fF
C10667 a_33086_11166# rowoff_n[9] 0.10fF
C10668 a_1962_17230# a_20034_17190# 0.27fF
C10669 m2_27836_18014# m2_28264_18442# 0.16fF
C10670 a_2346_13216# col[31] 0.15fF
C10671 a_29070_3134# VDD 0.52fF
C10672 m3_34996_6098# ctop 0.23fF
C10673 a_19334_4178# vcm 0.22fF
C10674 a_8898_14178# a_8990_14178# 0.26fF
C10675 a_1962_14218# a_13310_14218# 0.14fF
C10676 a_2346_14220# a_15014_14178# 0.19fF
C10677 a_3970_10162# col_n[1] 0.28fF
C10678 m2_34864_7974# m2_34864_6970# 0.99fF
C10679 a_8898_6146# VDD 0.23fF
C10680 a_30074_7150# a_31078_7150# 0.97fF
C10681 a_3970_17190# ctop 3.38fF
C10682 a_31078_10162# row_n[8] 0.17fF
C10683 a_22042_6146# col_n[19] 0.28fF
C10684 a_1962_3174# col_n[9] 0.13fF
C10685 col_n[27] row_n[4] 0.23fF
C10686 col_n[16] ctop 2.04fF
C10687 col_n[5] col[5] 0.72fF
C10688 col_n[21] row_n[1] 0.23fF
C10689 VDD col[14] 4.17fF
C10690 col_n[29] row_n[5] 0.23fF
C10691 col_n[19] row_n[0] 0.23fF
C10692 col_n[25] row_n[3] 0.23fF
C10693 col_n[23] row_n[2] 0.23fF
C10694 col_n[31] row_n[6] 0.23fF
C10695 vcm col[10] 5.84fF
C10696 rowon_n[11] rowon_n[10] 0.15fF
C10697 a_1962_16226# col_n[11] 0.13fF
C10698 a_32386_8194# vcm 0.22fF
C10699 a_1962_16226# a_26362_16226# 0.14fF
C10700 a_32082_17190# a_32082_16186# 1.00fF
C10701 a_2346_16228# a_28066_16186# 0.19fF
C10702 a_14010_2130# ctop 3.39fF
C10703 m2_4744_18014# VDD 0.91fF
C10704 a_33086_10162# m2_33284_10410# 0.16fF
C10705 a_1962_18234# m2_19804_18014# 0.18fF
C10706 a_1962_10202# col[2] 0.11fF
C10707 a_21950_10162# VDD 0.23fF
C10708 a_2346_8196# a_4882_8154# 0.35fF
C10709 a_20946_12170# rowoff_n[10] 0.24fF
C10710 a_7894_4138# rowoff_n[2] 0.24fF
C10711 a_2346_9200# col[22] 0.15fF
C10712 a_19030_8154# rowon_n[6] 0.14fF
C10713 a_27062_6146# ctop 3.58fF
C10714 m2_34864_1950# row_n[0] 0.15fF
C10715 m3_31984_1078# VDD 0.15fF
C10716 a_1962_18234# col_n[21] 0.13fF
C10717 a_2346_18236# m2_14784_18014# 0.19fF
C10718 a_35002_14178# VDD 0.29fF
C10719 a_2346_10204# a_17934_10162# 0.35fF
C10720 a_17934_2130# rowoff_n[0] 0.24fF
C10721 a_7986_5142# vcm 0.62fF
C10722 a_1962_15222# a_34394_15222# 0.14fF
C10723 a_35002_16186# rowoff_n[14] 0.24fF
C10724 a_1962_5182# col[29] 0.11fF
C10725 a_15014_3134# a_15014_2130# 1.00fF
C10726 a_31990_3134# a_32082_3134# 0.26fF
C10727 m2_5748_18014# m3_4876_18146# 0.13fF
C10728 a_1962_7190# a_12002_7150# 0.27fF
C10729 a_14010_17190# VDD 0.55fF
C10730 a_20034_9158# col[17] 0.29fF
C10731 m2_34864_16006# vcm 0.50fF
C10732 a_2346_12212# a_30986_12170# 0.35fF
C10733 a_16018_12170# a_17022_12170# 0.97fF
C10734 a_1962_12210# col_n[2] 0.13fF
C10735 a_21038_9158# vcm 0.62fF
C10736 a_4274_18234# vcm 0.22fF
C10737 a_24050_2130# VDD 0.55fF
C10738 a_30074_11166# m2_30272_11414# 0.16fF
C10739 a_2346_4180# a_6982_4138# 0.19fF
C10740 a_1962_4178# a_5278_4178# 0.14fF
C10741 a_4882_4138# a_4974_4138# 0.26fF
C10742 m3_1864_9110# m3_1864_8106# 0.22fF
C10743 a_1962_9198# a_25054_9158# 0.27fF
C10744 a_14314_3174# vcm 0.22fF
C10745 a_16018_11166# row_n[9] 0.17fF
C10746 a_5978_10162# rowoff_n[8] 0.10fF
C10747 a_34090_13174# vcm 0.62fF
C10748 a_2346_5184# col[13] 0.15fF
C10749 a_7986_13174# rowoff_n[11] 0.10fF
C10750 col[15] rowoff_n[0] 0.11fF
C10751 col[18] rowoff_n[3] 0.11fF
C10752 col[16] rowoff_n[1] 0.11fF
C10753 col[20] rowoff_n[5] 0.11fF
C10754 col[19] rowoff_n[4] 0.11fF
C10755 col[17] rowoff_n[2] 0.11fF
C10756 col[24] rowoff_n[9] 0.11fF
C10757 col[23] rowoff_n[8] 0.11fF
C10758 col[22] rowoff_n[7] 0.11fF
C10759 col[21] rowoff_n[6] 0.11fF
C10760 a_2346_6188# a_20034_6146# 0.19fF
C10761 a_28066_7150# a_28066_6146# 1.00fF
C10762 a_1962_6186# a_18330_6186# 0.14fF
C10763 a_16018_8154# rowoff_n[6] 0.10fF
C10764 a_1962_7190# col_n[29] 0.13fF
C10765 a_27366_7190# vcm 0.22fF
C10766 a_29070_16186# a_30074_16186# 0.97fF
C10767 a_2874_1126# m2_2736_946# 0.16fF
C10768 a_20034_11166# col_n[17] 0.28fF
C10769 a_1962_1166# col[20] 0.11fF
C10770 a_22042_17190# rowoff_n[15] 0.10fF
C10771 a_1962_14218# col[22] 0.11fF
C10772 a_26058_6146# rowoff_n[4] 0.10fF
C10773 a_3970_9158# rowon_n[7] 0.14fF
C10774 a_16930_9158# VDD 0.23fF
C10775 m2_13780_18014# col_n[11] 0.25fF
C10776 a_17934_8154# a_18026_8154# 0.26fF
C10777 a_2346_8196# a_33086_8154# 0.19fF
C10778 a_1962_8194# a_31382_8194# 0.14fF
C10779 m2_11772_946# ctop 0.18fF
C10780 a_1962_18234# a_7286_18234# 0.14fF
C10781 m2_1732_6970# sample 0.19fF
C10782 m2_4744_946# m2_5172_1374# 0.16fF
C10783 col[8] rowoff_n[10] 0.11fF
C10784 m2_9764_18014# m2_10768_18014# 0.96fF
C10785 a_22042_5142# ctop 3.58fF
C10786 m2_28840_946# ctop 0.18fF
C10787 a_27062_12170# m2_27260_12418# 0.16fF
C10788 a_29982_13174# VDD 0.23fF
C10789 a_2346_1168# col[4] 0.14fF
C10790 a_2346_14220# col[6] 0.15fF
C10791 a_23046_12170# rowon_n[10] 0.14fF
C10792 a_2346_2172# a_22954_2130# 0.35fF
C10793 a_12002_2130# a_13006_2130# 0.97fF
C10794 a_1962_3174# col_n[20] 0.13fF
C10795 col_n[10] col[11] 5.98fF
C10796 col_n[27] ctop 2.02fF
C10797 VDD col[25] 4.18fF
C10798 a_8990_16186# VDD 0.52fF
C10799 vcm col[21] 5.84fF
C10800 col_n[30] row_n[0] 0.23fF
C10801 rowon_n[8] row_n[8] 19.75fF
C10802 a_1962_16226# col_n[22] 0.13fF
C10803 a_14010_12170# a_14010_11166# 1.00fF
C10804 a_30986_12170# a_31078_12170# 0.26fF
C10805 a_16018_8154# vcm 0.62fF
C10806 a_1962_16226# a_9994_16186# 0.27fF
C10807 a_18026_14178# col[15] 0.29fF
C10808 a_34090_3134# m2_34864_2954# 0.96fF
C10809 a_1962_10202# col[13] 0.11fF
C10810 a_19030_1126# VDD 0.58fF
C10811 m2_34864_13998# rowon_n[12] 0.13fF
C10812 a_3878_10162# VDD 0.23fF
C10813 a_16018_2130# row_n[0] 0.17fF
C10814 a_2966_7150# col[0] 0.29fF
C10815 a_9294_2170# vcm 0.22fF
C10816 a_1962_13214# a_3270_13214# 0.14fF
C10817 a_2346_13216# a_4974_13174# 0.19fF
C10818 a_35002_10162# rowoff_n[8] 0.24fF
C10819 a_29070_12170# vcm 0.62fF
C10820 a_32082_5142# VDD 0.52fF
C10821 m3_27968_18146# VDD 0.29fF
C10822 a_25054_6146# a_26058_6146# 0.97fF
C10823 a_24050_13174# m2_24248_13422# 0.16fF
C10824 m2_20808_946# a_20034_1126# 0.96fF
C10825 a_20034_15182# row_n[13] 0.17fF
C10826 a_22346_6186# vcm 0.22fF
C10827 a_2346_15224# a_18026_15182# 0.19fF
C10828 a_1962_15222# a_16322_15222# 0.14fF
C10829 a_27062_16186# a_27062_15182# 1.00fF
C10830 a_30074_2130# m3_29976_1078# 0.15fF
C10831 a_11910_8154# VDD 0.23fF
C10832 a_18026_16186# col_n[15] 0.28fF
C10833 a_1962_12210# col_n[13] 0.13fF
C10834 a_19030_3134# col[16] 0.29fF
C10835 a_2966_9158# vcm 0.61fF
C10836 a_1962_17230# a_29374_17230# 0.14fF
C10837 a_2346_17232# a_31078_17190# 0.19fF
C10838 a_16930_17190# a_17022_17190# 0.26fF
C10839 a_1962_6186# col[4] 0.11fF
C10840 a_17022_4138# ctop 3.58fF
C10841 m2_5748_946# m3_5880_1078# 2.79fF
C10842 m3_34568_1078# ctop 0.38fF
C10843 a_7986_13174# rowon_n[11] 0.14fF
C10844 a_24962_12170# VDD 0.23fF
C10845 m3_16924_18146# m3_17928_18146# 0.22fF
C10846 a_2346_9200# a_7894_9158# 0.35fF
C10847 m2_1732_16006# row_n[14] 0.13fF
C10848 a_2346_5184# col[24] 0.15fF
C10849 a_8990_3134# rowoff_n[1] 0.10fF
C10850 a_23046_3134# rowon_n[1] 0.14fF
C10851 col[30] rowoff_n[4] 0.11fF
C10852 col[29] rowoff_n[3] 0.11fF
C10853 col[28] rowoff_n[2] 0.11fF
C10854 col[27] rowoff_n[1] 0.11fF
C10855 col[31] rowoff_n[5] 0.11fF
C10856 col[26] rowoff_n[0] 0.11fF
C10857 a_24050_14178# rowoff_n[12] 0.10fF
C10858 a_1962_6186# m2_1732_5966# 0.15fF
C10859 a_26970_2130# a_27062_2130# 0.26fF
C10860 a_30074_8154# ctop 3.58fF
C10861 a_21038_14178# m2_21236_14426# 0.16fF
C10862 a_3970_15182# VDD 0.52fF
C10863 a_10998_11166# a_12002_11166# 0.97fF
C10864 a_2346_11208# a_20946_11166# 0.35fF
C10865 a_10998_7150# vcm 0.62fF
C10866 a_19030_5142# col_n[16] 0.28fF
C10867 a_27062_16186# rowon_n[14] 0.14fF
C10868 a_1962_8194# col_n[4] 0.13fF
C10869 a_1962_8194# a_15014_8154# 0.27fF
C10870 a_4274_1166# vcm 0.22fF
C10871 a_2346_13216# a_33998_13174# 0.35fF
C10872 col[19] rowoff_n[10] 0.11fF
C10873 a_24050_11166# vcm 0.62fF
C10874 a_4974_16186# row_n[14] 0.17fF
C10875 a_34090_15182# col[31] 0.29fF
C10876 a_27062_4138# VDD 0.52fF
C10877 a_1962_5182# a_8290_5182# 0.14fF
C10878 a_23046_6146# a_23046_5142# 1.00fF
C10879 a_2346_5184# a_9994_5142# 0.19fF
C10880 a_20034_6146# row_n[4] 0.17fF
C10881 a_1962_10202# a_28066_10162# 0.27fF
C10882 a_7894_9158# rowoff_n[7] 0.24fF
C10883 a_2346_1168# col[15] 0.14fF
C10884 a_2346_14220# col[17] 0.15fF
C10885 a_17326_5182# vcm 0.22fF
C10886 a_24050_15182# a_25054_15182# 0.97fF
C10887 a_11910_15182# rowoff_n[13] 0.24fF
C10888 a_1962_3174# col_n[31] 0.13fF
C10889 col_n[16] col[16] 0.64fF
C10890 vcm rowoff_n[15] 0.20fF
C10891 m2_19804_18014# m3_19936_18146# 2.79fF
C10892 rowon_n[12] ctop 1.40fF
C10893 a_6890_7150# VDD 0.23fF
C10894 a_17934_7150# rowoff_n[5] 0.24fF
C10895 a_12914_7150# a_13006_7150# 0.26fF
C10896 a_18026_15182# m2_18224_15430# 0.16fF
C10897 a_1962_7190# a_21342_7190# 0.14fF
C10898 a_2346_7192# a_23046_7150# 0.19fF
C10899 col[3] rowoff_n[11] 0.11fF
C10900 a_1962_10202# col[24] 0.11fF
C10901 a_30378_9198# vcm 0.22fF
C10902 a_17022_8154# col[14] 0.29fF
C10903 a_20034_3134# m2_20232_3382# 0.16fF
C10904 a_7986_4138# rowon_n[2] 0.14fF
C10905 a_27974_5142# rowoff_n[3] 0.24fF
C10906 a_12002_3134# ctop 3.57fF
C10907 a_19942_11166# VDD 0.23fF
C10908 m3_6884_1078# m3_7888_1078# 0.22fF
C10909 a_1962_9198# a_35398_9198# 0.14fF
C10910 a_2346_9200# a_2346_8196# 0.22fF
C10911 a_34090_17190# col_n[31] 0.28fF
C10912 a_2346_18236# a_1962_18234# 2.62fF
C10913 m2_2736_946# VDD 0.65fF
C10914 a_2346_1168# a_12914_1126# 0.35fF
C10915 a_25054_7150# ctop 3.58fF
C10916 a_12002_17190# rowon_n[15] 0.14fF
C10917 a_32994_15182# VDD 0.23fF
C10918 a_25966_11166# a_26058_11166# 0.26fF
C10919 a_8990_11166# a_8990_10162# 1.00fF
C10920 a_2346_10204# col[8] 0.15fF
C10921 a_27062_7150# rowon_n[5] 0.14fF
C10922 a_5978_6146# vcm 0.62fF
C10923 a_1962_12210# col_n[24] 0.13fF
C10924 a_2346_3176# a_25966_3134# 0.35fF
C10925 a_17022_10162# col_n[14] 0.28fF
C10926 a_15014_16186# m2_15212_16434# 0.16fF
C10927 a_4974_7150# row_n[5] 0.17fF
C10928 a_1962_6186# col[15] 0.11fF
C10929 a_2346_11208# rowon_n[9] 0.26fF
C10930 a_26058_11166# rowoff_n[9] 0.10fF
C10931 a_19030_10162# vcm 0.62fF
C10932 a_1962_17230# a_13006_17190# 0.27fF
C10933 a_17022_4138# m2_17220_4386# 0.16fF
C10934 m2_20808_18014# m2_21236_18442# 0.16fF
C10935 a_22042_3134# VDD 0.52fF
C10936 m3_30980_18146# ctop 0.23fF
C10937 a_20034_5142# a_21038_5142# 0.97fF
C10938 m2_28840_18014# col[26] 0.28fF
C10939 a_12306_4178# vcm 0.22fF
C10940 a_2346_14220# a_7986_14178# 0.19fF
C10941 a_1962_14218# a_6282_14218# 0.14fF
C10942 a_22042_15182# a_22042_14178# 1.00fF
C10943 a_32082_14178# vcm 0.62fF
C10944 m2_34864_6970# VDD 1.01fF
C10945 a_1962_2170# a_33086_2130# 0.27fF
C10946 a_24050_10162# row_n[8] 0.17fF
C10947 a_2346_11208# a_1962_11206# 2.62fF
C10948 a_25358_8194# vcm 0.22fF
C10949 a_11910_16186# a_12002_16186# 0.26fF
C10950 a_2346_16228# a_21038_16186# 0.19fF
C10951 a_1962_16226# a_19334_16226# 0.14fF
C10952 a_6982_2130# ctop 3.39fF
C10953 a_1962_8194# col_n[15] 0.13fF
C10954 a_1962_18234# m2_5748_18014# 0.18fF
C10955 a_15014_13174# col[12] 0.29fF
C10956 a_14922_10162# VDD 0.23fF
C10957 col[30] rowoff_n[10] 0.11fF
C10958 a_12002_17190# m2_12200_17438# 0.16fF
C10959 a_33086_9158# a_34090_9158# 0.97fF
C10960 a_1962_2170# col[6] 0.11fF
C10961 a_1962_15222# col[8] 0.11fF
C10962 m2_1732_3958# ctop 0.17fF
C10963 a_13918_12170# rowoff_n[10] 0.24fF
C10964 a_12002_8154# rowon_n[6] 0.14fF
C10965 a_33086_9158# col[30] 0.29fF
C10966 a_14010_5142# m2_14208_5390# 0.16fF
C10967 a_20034_6146# ctop 3.58fF
C10968 m3_3872_1078# VDD 0.11fF
C10969 a_2346_1168# col[26] 0.14fF
C10970 a_27974_14178# VDD 0.23fF
C10971 a_2346_14220# col[28] 0.15fF
C10972 a_5978_10162# a_6982_10162# 0.97fF
C10973 a_2346_10204# a_10906_10162# 0.35fF
C10974 a_10906_2130# rowoff_n[0] 0.24fF
C10975 a_2346_18236# col[0] 0.15fF
C10976 col_n[21] col[22] 5.98fF
C10977 row_n[7] ctop 1.65fF
C10978 a_27974_16186# rowoff_n[14] 0.24fF
C10979 m2_27836_18014# ctop 0.18fF
C10980 a_33086_10162# ctop 3.57fF
C10981 a_32994_1126# m2_32856_946# 0.16fF
C10982 col[14] rowoff_n[11] 0.11fF
C10983 a_1962_7190# a_4974_7150# 0.27fF
C10984 a_3878_7150# a_3970_7150# 0.26fF
C10985 m2_34864_2954# row_n[1] 0.15fF
C10986 a_6982_17190# VDD 0.55fF
C10987 a_2346_2172# rowon_n[0] 0.26fF
C10988 a_15014_15182# col_n[12] 0.28fF
C10989 a_2346_12212# a_23958_12170# 0.35fF
C10990 m2_15788_946# m3_14916_1078# 0.13fF
C10991 a_31078_11166# rowon_n[9] 0.14fF
C10992 a_16018_2130# col[13] 0.29fF
C10993 a_14010_9158# vcm 0.62fF
C10994 a_1962_4178# col_n[6] 0.13fF
C10995 a_1962_17230# col_n[8] 0.13fF
C10996 a_17022_2130# VDD 0.55fF
C10997 a_18026_5142# a_18026_4138# 1.00fF
C10998 a_35494_12532# VDD 0.11fF
C10999 m2_26832_946# m3_26964_1078# 2.79fF
C11000 m3_1864_16138# m3_1864_15134# 0.22fF
C11001 a_33086_11166# col_n[30] 0.28fF
C11002 a_1962_9198# a_18026_9158# 0.27fF
C11003 a_8990_11166# row_n[9] 0.17fF
C11004 a_7286_3174# vcm 0.22fF
C11005 a_1962_14218# a_1962_13214# 0.16fF
C11006 a_19030_14178# a_20034_14178# 0.97fF
C11007 a_27062_13174# vcm 0.62fF
C11008 a_10998_6146# m2_11196_6394# 0.16fF
C11009 a_30074_6146# VDD 0.52fF
C11010 a_2346_6188# a_13006_6146# 0.19fF
C11011 a_1962_6186# a_11302_6186# 0.14fF
C11012 a_7894_6146# a_7986_6146# 0.26fF
C11013 a_2346_10204# col[19] 0.15fF
C11014 a_8990_8154# rowoff_n[6] 0.10fF
C11015 a_1962_11206# a_31078_11166# 0.27fF
C11016 a_6982_17190# m3_6884_18146# 0.15fF
C11017 a_20338_7190# vcm 0.22fF
C11018 a_15014_17190# rowoff_n[15] 0.10fF
C11019 a_19030_6146# rowoff_n[4] 0.10fF
C11020 a_16018_4138# col_n[13] 0.28fF
C11021 a_9902_9158# VDD 0.23fF
C11022 a_1962_8194# a_24354_8194# 0.14fF
C11023 a_2346_8196# a_26058_8154# 0.19fF
C11024 a_31078_9158# a_31078_8154# 1.00fF
C11025 a_28066_14178# row_n[12] 0.17fF
C11026 a_1962_6186# col[26] 0.11fF
C11027 a_33390_11206# vcm 0.22fF
C11028 a_29070_4138# rowoff_n[2] 0.10fF
C11029 m2_4744_946# ctop 0.20fF
C11030 m2_2736_18014# m2_3740_18014# 0.96fF
C11031 a_2966_4138# m2_1732_3958# 0.96fF
C11032 a_1962_13214# col_n[0] 0.13fF
C11033 a_15014_5142# ctop 3.58fF
C11034 a_22954_13174# VDD 0.23fF
C11035 a_31078_14178# col[28] 0.29fF
C11036 a_3970_10162# a_3970_9158# 1.00fF
C11037 a_20946_10162# a_21038_10162# 0.26fF
C11038 a_16018_12170# rowon_n[10] 0.14fF
C11039 a_7986_7150# m2_8184_7398# 0.16fF
C11040 a_2346_2172# a_15926_2130# 0.35fF
C11041 m2_33860_18014# m3_34996_18146# 0.13fF
C11042 a_28066_9158# ctop 3.58fF
C11043 a_2346_6188# col[10] 0.15fF
C11044 a_31078_2130# rowon_n[0] 0.14fF
C11045 a_8990_8154# vcm 0.62fF
C11046 a_1962_8194# col_n[26] 0.13fF
C11047 a_2346_16228# a_2966_16186# 0.21fF
C11048 m2_26832_946# col_n[24] 0.37fF
C11049 a_14010_7150# col[11] 0.29fF
C11050 a_15014_4138# a_16018_4138# 0.97fF
C11051 a_2346_4180# a_28978_4138# 0.35fF
C11052 m2_15788_946# col[13] 0.39fF
C11053 a_8990_2130# row_n[0] 0.17fF
C11054 a_1962_2170# col[17] 0.11fF
C11055 a_9994_17190# m2_9764_18014# 1.00fF
C11056 a_1962_15222# col[19] 0.11fF
C11057 a_17022_14178# a_17022_13174# 1.00fF
C11058 a_33998_14178# a_34090_14178# 0.26fF
C11059 a_27974_10162# rowoff_n[8] 0.24fF
C11060 a_31078_16186# col_n[28] 0.28fF
C11061 a_29982_13174# rowoff_n[11] 0.24fF
C11062 a_22042_12170# vcm 0.62fF
C11063 a_32082_3134# col[29] 0.29fF
C11064 a_25054_5142# VDD 0.52fF
C11065 a_2346_18236# col[11] 0.14fF
C11066 rowon_n[1] ctop 1.39fF
C11067 col_n[27] col[27] 0.77fF
C11068 a_13006_15182# row_n[13] 0.17fF
C11069 a_15318_6186# vcm 0.22fF
C11070 a_6890_15182# a_6982_15182# 0.26fF
C11071 a_2346_15224# a_10998_15182# 0.19fF
C11072 a_1962_15222# a_9294_15222# 0.14fF
C11073 m2_1732_10986# m2_1732_9982# 0.99fF
C11074 col[25] rowoff_n[11] 0.11fF
C11075 a_35094_16186# vcm 0.12fF
C11076 m2_20808_946# m2_21236_1374# 0.16fF
C11077 a_28066_5142# row_n[3] 0.17fF
C11078 a_4974_8154# m2_5172_8402# 0.16fF
C11079 a_2346_2172# col[1] 0.15fF
C11080 a_4882_8154# VDD 0.23fF
C11081 a_2346_15224# col[3] 0.15fF
C11082 a_28066_8154# a_29070_8154# 0.97fF
C11083 a_14010_9158# col_n[11] 0.28fF
C11084 a_1962_4178# col_n[17] 0.13fF
C11085 a_1962_17230# col_n[19] 0.13fF
C11086 a_28370_10202# vcm 0.22fF
C11087 a_2346_17232# a_24050_17190# 0.19fF
C11088 a_1962_17230# a_22346_17230# 0.14fF
C11089 a_9994_4138# ctop 3.58fF
C11090 m3_6884_1078# ctop 0.23fF
C11091 a_32082_5142# col_n[29] 0.28fF
C11092 a_17934_12170# VDD 0.23fF
C11093 m3_2868_18146# m3_3872_18146# 0.22fF
C11094 a_1962_11206# col[10] 0.11fF
C11095 a_16018_3134# rowon_n[1] 0.14fF
C11096 col[9] rowoff_n[12] 0.11fF
C11097 a_17022_14178# rowoff_n[12] 0.10fF
C11098 a_2346_10204# col[30] 0.15fF
C11099 a_23046_8154# ctop 3.58fF
C11100 m2_34864_15002# m3_34996_16138# 0.15fF
C11101 a_30986_16186# VDD 0.23fF
C11102 a_2346_11208# a_13918_11166# 0.35fF
C11103 a_3970_7150# vcm 0.62fF
C11104 a_8990_2130# m2_8760_946# 0.99fF
C11105 a_20034_16186# rowon_n[14] 0.14fF
C11106 a_29982_4138# a_30074_4138# 0.26fF
C11107 a_13006_4138# a_13006_3134# 1.00fF
C11108 a_2346_11208# ctop 1.59fF
C11109 a_1962_8194# a_7986_8154# 0.27fF
C11110 a_29070_17190# m2_28840_18014# 1.00fF
C11111 a_12002_12170# col[9] 0.29fF
C11112 a_2346_13216# a_26970_13174# 0.35fF
C11113 a_14010_13174# a_15014_13174# 0.97fF
C11114 a_1962_13214# col_n[10] 0.13fF
C11115 a_17022_11166# vcm 0.62fF
C11116 a_20034_4138# VDD 0.52fF
C11117 a_2346_5184# a_2874_5142# 0.35fF
C11118 a_1962_7190# col[1] 0.11fF
C11119 a_30074_8154# col[27] 0.29fF
C11120 a_13006_6146# row_n[4] 0.17fF
C11121 a_1962_10202# a_21038_10162# 0.27fF
C11122 a_10298_5182# vcm 0.22fF
C11123 a_30074_15182# vcm 0.62fF
C11124 a_4882_15182# rowoff_n[13] 0.24fF
C11125 m2_1732_9982# VDD 1.02fF
C11126 a_2346_6188# col[21] 0.15fF
C11127 m2_10768_18014# m3_9896_18146# 0.13fF
C11128 a_33086_8154# VDD 0.52fF
C11129 a_10906_7150# rowoff_n[5] 0.24fF
C11130 a_1962_7190# a_14314_7190# 0.14fF
C11131 a_26058_8154# a_26058_7150# 1.00fF
C11132 a_2346_7192# a_16018_7150# 0.19fF
C11133 a_1962_12210# a_34090_12170# 0.27fF
C11134 a_23350_9198# vcm 0.22fF
C11135 a_27062_17190# a_28066_17190# 0.97fF
C11136 a_12002_14178# col_n[9] 0.28fF
C11137 a_20946_5142# rowoff_n[3] 0.24fF
C11138 a_4974_3134# ctop 3.57fF
C11139 a_1962_2170# col[28] 0.11fF
C11140 a_32082_9158# row_n[7] 0.17fF
C11141 a_1962_15222# col[30] 0.11fF
C11142 a_33086_11166# m2_33284_11414# 0.16fF
C11143 a_12914_11166# VDD 0.23fF
C11144 a_15926_9158# a_16018_9158# 0.26fF
C11145 a_1962_9198# a_27366_9198# 0.14fF
C11146 a_2346_9200# a_29070_9158# 0.19fF
C11147 a_30986_3134# rowoff_n[1] 0.24fF
C11148 a_30074_10162# col_n[27] 0.28fF
C11149 a_1962_9198# col_n[1] 0.13fF
C11150 a_2346_1168# a_5886_1126# 0.35fF
C11151 m2_34864_11990# m3_34996_13126# 0.15fF
C11152 a_18026_7150# ctop 3.58fF
C11153 a_2346_18236# col[22] 0.14fF
C11154 a_4974_17190# rowon_n[15] 0.14fF
C11155 a_1962_16226# ctop 1.49fF
C11156 ctop analog_in 0.71fF
C11157 a_25966_15182# VDD 0.23fF
C11158 a_20034_7150# rowon_n[5] 0.14fF
C11159 a_5886_1126# m2_5748_946# 0.16fF
C11160 a_2346_2172# col[12] 0.15fF
C11161 a_2346_15224# col[14] 0.15fF
C11162 a_9994_3134# a_10998_3134# 0.97fF
C11163 a_2346_3176# a_18938_3134# 0.35fF
C11164 a_31078_11166# ctop 3.58fF
C11165 a_1962_4178# col_n[28] 0.13fF
C11166 m2_20808_946# ctop 0.20fF
C11167 a_13006_3134# col_n[10] 0.28fF
C11168 a_1962_17230# col_n[30] 0.13fF
C11169 a_12002_13174# a_12002_12170# 1.00fF
C11170 a_28978_13174# a_29070_13174# 0.26fF
C11171 a_12002_10162# vcm 0.62fF
C11172 a_19030_11166# rowoff_n[9] 0.10fF
C11173 a_1962_17230# a_5978_17190# 0.27fF
C11174 a_9994_17190# col[7] 0.29fF
C11175 a_1962_18234# col[4] 0.11fF
C11176 m2_13780_18014# m2_14208_18442# 0.16fF
C11177 a_15014_3134# VDD 0.52fF
C11178 a_1962_11206# col[21] 0.11fF
C11179 m3_2868_18146# ctop 0.23fF
C11180 a_30074_12170# m2_30272_12418# 0.16fF
C11181 a_2346_5184# a_31990_5142# 0.35fF
C11182 col[20] rowoff_n[12] 0.11fF
C11183 a_29070_9158# rowoff_n[7] 0.10fF
C11184 a_5278_4178# vcm 0.22fF
C11185 a_28066_13174# col[25] 0.29fF
C11186 a_33086_15182# rowoff_n[13] 0.10fF
C11187 a_25054_14178# vcm 0.62fF
C11188 m2_34864_4962# rowon_n[3] 0.13fF
C11189 a_1962_2170# a_26058_2130# 0.27fF
C11190 m2_1732_16006# m3_1864_16138# 2.76fF
C11191 a_28066_7150# VDD 0.52fF
C11192 a_23046_7150# a_24050_7150# 0.97fF
C11193 a_17022_10162# row_n[8] 0.17fF
C11194 a_18330_8194# vcm 0.22fF
C11195 a_1962_16226# a_12306_16226# 0.14fF
C11196 a_2346_16228# a_14010_16186# 0.19fF
C11197 a_25054_17190# a_25054_16186# 1.00fF
C11198 a_2346_11208# col[5] 0.15fF
C11199 a_7894_10162# VDD 0.23fF
C11200 col[4] rowoff_n[13] 0.11fF
C11201 a_10998_6146# col[8] 0.29fF
C11202 a_1962_13214# col_n[21] 0.13fF
C11203 a_31382_12210# vcm 0.22fF
C11204 a_6890_12170# rowoff_n[10] 0.24fF
C11205 m2_7756_18014# col_n[5] 0.25fF
C11206 a_4974_8154# rowon_n[6] 0.14fF
C11207 a_1962_1166# a_32386_1166# 0.14fF
C11208 a_28066_15182# col_n[25] 0.28fF
C11209 a_1962_7190# col[12] 0.11fF
C11210 a_13006_6146# ctop 3.58fF
C11211 m2_34864_8978# m3_34996_10114# 0.15fF
C11212 a_27062_13174# m2_27260_13422# 0.16fF
C11213 m3_34996_14130# VDD 0.26fF
C11214 a_29070_2130# col[26] 0.29fF
C11215 a_20946_14178# VDD 0.23fF
C11216 a_1962_10202# a_2966_10162# 0.27fF
C11217 m2_1732_946# sample_n 0.13fF
C11218 m2_13780_18014# ctop 0.18fF
C11219 a_20946_16186# rowoff_n[14] 0.24fF
C11220 a_7986_3134# a_7986_2130# 1.00fF
C11221 a_24962_3134# a_25054_3134# 0.26fF
C11222 a_26058_10162# ctop 3.58fF
C11223 a_33086_2130# m3_32988_1078# 0.15fF
C11224 m2_1732_6970# row_n[5] 0.13fF
C11225 a_33998_18194# VDD 0.33fF
C11226 a_8990_12170# a_9994_12170# 0.97fF
C11227 a_2346_12212# a_16930_12170# 0.35fF
C11228 a_24050_11166# rowon_n[9] 0.14fF
C11229 a_6982_9158# vcm 0.62fF
C11230 a_10998_8154# col_n[8] 0.28fF
C11231 a_34090_4138# m2_34864_3958# 0.96fF
C11232 m2_10768_946# m3_10900_1078# 2.79fF
C11233 a_9994_2130# VDD 0.55fF
C11234 a_1962_9198# col_n[12] 0.13fF
C11235 a_8898_18194# m2_8760_18014# 0.16fF
C11236 a_1962_9198# a_10998_9158# 0.27fF
C11237 a_29070_4138# col_n[26] 0.28fF
C11238 a_2346_14220# a_29982_14178# 0.35fF
C11239 a_2966_6146# col_n[0] 0.28fF
C11240 a_20034_13174# vcm 0.62fF
C11241 a_1962_3174# col[3] 0.11fF
C11242 ctop col[10] 1.98fF
C11243 a_1962_16226# col[5] 0.11fF
C11244 m2_1732_12994# m3_1864_13126# 2.76fF
C11245 a_23046_6146# VDD 0.52fF
C11246 a_1962_6186# a_4274_6186# 0.14fF
C11247 a_21038_7150# a_21038_6146# 1.00fF
C11248 a_24050_14178# m2_24248_14426# 0.16fF
C11249 a_2346_6188# a_5978_6146# 0.19fF
C11250 a_1962_11206# a_24050_11166# 0.27fF
C11251 a_2346_2172# col[23] 0.15fF
C11252 a_13310_7190# vcm 0.22fF
C11253 a_2346_15224# col[25] 0.15fF
C11254 a_22042_16186# a_23046_16186# 0.97fF
C11255 a_7986_17190# rowoff_n[15] 0.10fF
C11256 a_33086_17190# vcm 0.60fF
C11257 m2_33860_18014# VDD 0.96fF
C11258 a_12002_6146# rowoff_n[4] 0.10fF
C11259 a_2346_9200# VDD 32.63fF
C11260 a_1962_8194# a_17326_8194# 0.14fF
C11261 a_10906_8154# a_10998_8154# 0.26fF
C11262 a_2346_8196# a_19030_8154# 0.19fF
C11263 a_21038_14178# row_n[12] 0.17fF
C11264 a_1962_18234# col[15] 0.11fF
C11265 a_26362_11206# vcm 0.22fF
C11266 a_8990_11166# col[6] 0.29fF
C11267 a_22042_4138# rowoff_n[2] 0.10fF
C11268 m2_34864_5966# m3_34996_7102# 0.15fF
C11269 a_7986_5142# ctop 3.58fF
C11270 m2_12776_946# vcm 0.42fF
C11271 col[31] rowoff_n[12] 0.11fF
C11272 a_1962_5182# col_n[3] 0.13fF
C11273 a_15926_13174# VDD 0.23fF
C11274 a_34090_11166# a_34090_10162# 1.00fF
C11275 a_1962_10202# a_30378_10202# 0.14fF
C11276 a_2346_10204# a_32082_10162# 0.19fF
C11277 a_32082_2130# rowoff_n[0] 0.10fF
C11278 a_27062_7150# col[24] 0.29fF
C11279 m2_29844_946# vcm 0.42fF
C11280 m2_34864_16006# ctop 0.17fF
C11281 a_8990_12170# rowon_n[10] 0.14fF
C11282 a_4974_2130# a_5978_2130# 0.97fF
C11283 a_2346_2172# a_8898_2130# 0.35fF
C11284 a_1962_7190# m2_1732_6970# 0.15fF
C11285 a_21038_9158# ctop 3.58fF
C11286 m2_24824_18014# m3_24956_18146# 2.78fF
C11287 a_21038_15182# m2_21236_15430# 0.16fF
C11288 a_28978_17190# VDD 0.24fF
C11289 a_24050_2130# rowon_n[0] 0.14fF
C11290 a_6982_12170# a_6982_11166# 1.00fF
C11291 a_23958_12170# a_24050_12170# 0.26fF
C11292 a_2346_11208# col[16] 0.15fF
C11293 a_34394_9198# vcm 0.22fF
C11294 m2_34864_16006# m2_35292_16434# 0.16fF
C11295 a_23046_3134# m2_23244_3382# 0.16fF
C11296 col[15] rowoff_n[13] 0.11fF
C11297 a_2346_4180# a_21950_4138# 0.35fF
C11298 a_8990_13174# col_n[6] 0.28fF
C11299 a_34090_13174# ctop 3.42fF
C11300 sample_n rowoff_n[8] 0.38fF
C11301 VDD rowoff_n[7] 1.17fF
C11302 a_27974_18194# m2_27836_18014# 0.16fF
C11303 a_20946_10162# rowoff_n[8] 0.24fF
C11304 a_28066_15182# rowon_n[13] 0.14fF
C11305 a_1962_7190# col[23] 0.11fF
C11306 a_22954_13174# rowoff_n[11] 0.24fF
C11307 a_15014_12170# vcm 0.62fF
C11308 m2_10768_946# VDD 0.62fF
C11309 a_27062_9158# col_n[24] 0.28fF
C11310 m2_1732_9982# m3_1864_10114# 2.76fF
C11311 a_18026_5142# VDD 0.52fF
C11312 a_2346_6188# a_35002_6146# 0.35fF
C11313 a_18026_6146# a_19030_6146# 0.97fF
C11314 a_1962_14218# VDD 2.73fF
C11315 a_30986_8154# rowoff_n[6] 0.24fF
C11316 a_5978_15182# row_n[13] 0.17fF
C11317 a_8290_6186# vcm 0.22fF
C11318 a_20034_16186# a_20034_15182# 1.00fF
C11319 a_2346_15224# a_3970_15182# 0.19fF
C11320 a_28066_16186# vcm 0.62fF
C11321 a_21038_5142# row_n[3] 0.17fF
C11322 a_1962_3174# a_29070_3134# 0.27fF
C11323 a_31078_9158# VDD 0.52fF
C11324 a_18026_16186# m2_18224_16434# 0.16fF
C11325 a_2346_7192# col[7] 0.15fF
C11326 a_21342_10202# vcm 0.22fF
C11327 a_9994_2130# col_n[7] 0.28fF
C11328 a_9902_17190# a_9994_17190# 0.26fF
C11329 a_2346_17232# a_17022_17190# 0.19fF
C11330 a_1962_17230# a_15318_17230# 0.14fF
C11331 a_20034_4138# m2_20232_4386# 0.16fF
C11332 m2_34864_2954# m3_34996_4090# 0.15fF
C11333 a_1962_9198# col_n[23] 0.13fF
C11334 m3_1864_12122# ctop 0.23fF
C11335 a_6982_16186# col[4] 0.29fF
C11336 a_10906_12170# VDD 0.23fF
C11337 a_31078_10162# a_32082_10162# 0.97fF
C11338 a_23046_2130# m2_22816_946# 0.99fF
C11339 a_1962_3174# col[14] 0.11fF
C11340 a_8990_3134# rowon_n[1] 0.14fF
C11341 sample_n sample 7.84fF
C11342 VDD col_n[0] 5.06fF
C11343 en_bit_n[0] col[17] 0.16fF
C11344 ctop col[21] 1.98fF
C11345 col[7] col[8] 0.20fF
C11346 a_1962_16226# col[16] 0.11fF
C11347 a_35398_14218# vcm 0.23fF
C11348 a_9994_14178# rowoff_n[12] 0.10fF
C11349 a_25054_12170# col[22] 0.29fF
C11350 a_19942_2130# a_20034_2130# 0.26fF
C11351 a_16018_8154# ctop 3.58fF
C11352 a_23958_16186# VDD 0.23fF
C11353 a_2346_11208# a_6890_11166# 0.35fF
C11354 a_3970_11166# a_4974_11166# 0.97fF
C11355 a_35002_1126# VDD 0.50fF
C11356 a_13006_16186# rowon_n[14] 0.14fF
C11357 a_29070_12170# ctop 3.58fF
C11358 a_15014_17190# m2_15212_17438# 0.16fF
C11359 a_1962_18234# col[26] 0.11fF
C11360 a_2966_14178# row_n[12] 0.16fF
C11361 a_28066_6146# rowon_n[4] 0.14fF
C11362 a_2346_13216# a_19942_13174# 0.35fF
C11363 a_2346_16228# col[0] 0.15fF
C11364 a_7986_5142# col[5] 0.29fF
C11365 a_9994_11166# vcm 0.62fF
C11366 a_17022_5142# m2_17220_5390# 0.16fF
C11367 m2_1732_6970# m3_1864_7102# 2.76fF
C11368 a_1962_5182# col_n[14] 0.13fF
C11369 a_13006_4138# VDD 0.52fF
C11370 a_16018_6146# a_16018_5142# 1.00fF
C11371 a_32994_6146# a_33086_6146# 0.26fF
C11372 a_5978_6146# row_n[4] 0.17fF
C11373 a_25054_14178# col_n[22] 0.28fF
C11374 a_1962_10202# a_14010_10162# 0.27fF
C11375 a_3270_5182# vcm 0.22fF
C11376 a_17022_15182# a_18026_15182# 0.97fF
C11377 a_2346_15224# a_32994_15182# 0.35fF
C11378 a_1962_12210# col[7] 0.11fF
C11379 m2_22816_18014# col[20] 0.28fF
C11380 a_23046_15182# vcm 0.62fF
C11381 a_2966_9158# ctop 3.42fF
C11382 m2_1046_19620# m3_1046_19620# 0.25fF
C11383 a_26058_8154# VDD 0.52fF
C11384 a_1962_7190# a_7286_7190# 0.14fF
C11385 a_5886_7150# a_5978_7150# 0.26fF
C11386 a_2346_7192# a_8990_7150# 0.19fF
C11387 a_2346_11208# col[27] 0.15fF
C11388 a_1962_12210# a_27062_12170# 0.27fF
C11389 m2_21812_946# m3_20940_1078# 0.13fF
C11390 a_16322_9198# vcm 0.22fF
C11391 col[26] rowoff_n[13] 0.11fF
C11392 a_13918_5142# rowoff_n[3] 0.24fF
C11393 vcm rowoff_n[0] 0.20fF
C11394 a_25054_9158# row_n[7] 0.17fF
C11395 a_7986_7150# col_n[5] 0.28fF
C11396 a_2346_4180# a_3878_4138# 0.35fF
C11397 a_2874_4138# a_2966_4138# 0.26fF
C11398 a_5886_11166# VDD 0.23fF
C11399 m2_31852_946# m3_31984_1078# 2.79fF
C11400 a_29070_10162# a_29070_9158# 1.00fF
C11401 a_2346_9200# a_22042_9158# 0.19fF
C11402 a_1962_9198# a_20338_9198# 0.14fF
C11403 a_23958_3134# rowoff_n[1] 0.24fF
C11404 a_29374_13214# vcm 0.22fF
C11405 a_26058_3134# col_n[23] 0.28fF
C11406 a_1962_1166# col_n[5] 0.13fF
C11407 a_14010_6146# m2_14208_6394# 0.16fF
C11408 a_10998_7150# ctop 3.58fF
C11409 a_1962_14218# col_n[7] 0.13fF
C11410 a_23046_17190# col[20] 0.29fF
C11411 a_18938_15182# VDD 0.23fF
C11412 a_18938_11166# a_19030_11166# 0.26fF
C11413 a_1962_11206# a_33390_11206# 0.14fF
C11414 a_9994_17190# m3_9896_18146# 0.15fF
C11415 col[10] rowoff_n[14] 0.11fF
C11416 a_13006_7150# rowon_n[5] 0.14fF
C11417 a_2346_3176# a_11910_3134# 0.35fF
C11418 a_2966_5142# row_n[3] 0.16fF
C11419 a_24050_11166# ctop 3.58fF
C11420 a_2346_7192# col[18] 0.15fF
C11421 a_12002_11166# rowoff_n[9] 0.10fF
C11422 a_4974_10162# vcm 0.62fF
C11423 m2_6752_18014# m2_7180_18442# 0.16fF
C11424 m2_1732_3958# m3_1864_4090# 2.76fF
C11425 a_7986_3134# VDD 0.52fF
C11426 a_5978_10162# col[3] 0.29fF
C11427 a_13006_5142# a_14010_5142# 0.97fF
C11428 a_2346_5184# a_24962_5142# 0.35fF
C11429 a_1962_3174# col[25] 0.11fF
C11430 vcm col_n[6] 2.80fF
C11431 VDD col_n[10] 4.94fF
C11432 a_32082_10162# rowon_n[8] 0.14fF
C11433 ctop rowoff_n[15] 0.42fF
C11434 a_1962_16226# col[27] 0.11fF
C11435 a_22042_9158# rowoff_n[7] 0.10fF
C11436 a_15014_15182# a_15014_14178# 1.00fF
C11437 a_31990_15182# a_32082_15182# 0.26fF
C11438 a_26058_15182# rowoff_n[13] 0.10fF
C11439 a_18026_14178# vcm 0.62fF
C11440 m2_1732_8978# rowon_n[7] 0.11fF
C11441 a_24050_6146# col[21] 0.29fF
C11442 a_1962_2170# a_19030_2130# 0.27fF
C11443 a_1962_10202# sample 0.14fF
C11444 a_10998_7150# m2_11196_7398# 0.16fF
C11445 a_21038_7150# VDD 0.52fF
C11446 a_32082_7150# rowoff_n[5] 0.10fF
C11447 a_2966_7150# a_2966_6146# 1.00fF
C11448 a_9994_10162# row_n[8] 0.17fF
C11449 a_11302_8194# vcm 0.22fF
C11450 a_4882_16186# a_4974_16186# 0.26fF
C11451 a_1962_16226# a_5278_16226# 0.14fF
C11452 a_2346_16228# a_6982_16186# 0.19fF
C11453 a_31078_18194# vcm 0.12fF
C11454 a_1962_4178# a_32082_4138# 0.27fF
C11455 a_2346_3176# col[9] 0.15fF
C11456 a_34090_11166# VDD 0.54fF
C11457 a_2346_16228# col[11] 0.15fF
C11458 a_26058_9158# a_27062_9158# 0.97fF
C11459 a_5978_12170# col_n[3] 0.28fF
C11460 a_1962_5182# col_n[25] 0.13fF
C11461 a_24354_12210# vcm 0.22fF
C11462 a_1962_1166# a_25358_1166# 0.14fF
C11463 a_2966_5142# m2_1732_4962# 0.96fF
C11464 a_5978_6146# ctop 3.58fF
C11465 a_29070_13174# row_n[11] 0.17fF
C11466 m3_14916_18146# VDD 0.37fF
C11467 a_24050_8154# col_n[21] 0.28fF
C11468 a_13918_14178# VDD 0.23fF
C11469 a_1962_12210# col[18] 0.11fF
C11470 m2_16792_946# a_18026_1126# 0.96fF
C11471 a_13918_16186# rowoff_n[14] 0.24fF
C11472 a_7986_8154# m2_8184_8402# 0.16fF
C11473 a_19030_10162# ctop 3.58fF
C11474 a_34090_2130# m3_34996_2082# 0.13fF
C11475 a_26970_18194# VDD 0.34fF
C11476 m2_28840_18014# vcm 0.28fF
C11477 a_2346_12212# a_9902_12170# 0.35fF
C11478 a_17022_11166# rowon_n[9] 0.14fF
C11479 a_2874_2130# VDD 0.24fF
C11480 m3_21944_1078# ctop 0.23fF
C11481 a_27974_5142# a_28066_5142# 0.26fF
C11482 a_10998_5142# a_10998_4138# 1.00fF
C11483 a_32082_14178# ctop 3.58fF
C11484 a_2346_12212# col[2] 0.15fF
C11485 a_1962_9198# a_3970_9158# 0.27fF
C11486 a_3970_15182# col[1] 0.29fF
C11487 a_12002_14178# a_13006_14178# 0.97fF
C11488 a_2346_14220# a_22954_14178# 0.35fF
C11489 a_1962_1166# col_n[16] 0.12fF
C11490 a_2346_18236# a_31990_18194# 0.35fF
C11491 a_1962_14218# col_n[18] 0.13fF
C11492 a_13006_13174# vcm 0.62fF
C11493 a_16018_6146# VDD 0.52fF
C11494 a_22042_11166# col[19] 0.29fF
C11495 col[21] rowoff_n[14] 0.11fF
C11496 a_1962_8194# col[9] 0.11fF
C11497 m2_1732_11990# rowoff_n[10] 0.12fF
C11498 a_1962_11206# a_17022_11166# 0.27fF
C11499 a_6282_7190# vcm 0.22fF
C11500 a_26058_17190# vcm 0.60fF
C11501 m2_19804_18014# VDD 1.05fF
C11502 a_2346_7192# col[29] 0.15fF
C11503 a_4974_6146# rowoff_n[4] 0.10fF
C11504 a_1962_18234# m2_34864_18014# 0.17fF
C11505 a_4974_9158# m2_5172_9406# 0.16fF
C11506 a_29070_10162# VDD 0.52fF
C11507 a_2346_8196# a_12002_8154# 0.19fF
C11508 a_24050_9158# a_24050_8154# 1.00fF
C11509 a_1962_8194# a_10298_8194# 0.14fF
C11510 a_14010_14178# row_n[12] 0.17fF
C11511 a_2346_1168# vcm 0.37fF
C11512 a_1962_13214# a_30074_13174# 0.27fF
C11513 m2_1732_1950# m2_2160_2378# 0.16fF
C11514 a_28066_12170# rowoff_n[10] 0.10fF
C11515 a_19334_11206# vcm 0.22fF
C11516 a_15014_4138# rowoff_n[2] 0.10fF
C11517 a_29070_4138# row_n[2] 0.17fF
C11518 a_3970_17190# col_n[1] 0.28fF
C11519 a_4974_4138# col[2] 0.29fF
C11520 VDD col_n[21] 4.94fF
C11521 col_n[8] col_n[9] 0.10fF
C11522 vcm col_n[17] 2.79fF
C11523 col[18] col[19] 0.20fF
C11524 col[5] rowoff_n[15] 0.11fF
C11525 a_2966_6146# m3_1864_6098# 0.14fF
C11526 a_8898_13174# VDD 0.23fF
C11527 a_2346_18236# m2_29844_18014# 0.19fF
C11528 m2_5748_946# vcm 0.42fF
C11529 a_13918_10162# a_14010_10162# 0.26fF
C11530 a_2346_10204# a_25054_10162# 0.19fF
C11531 a_1962_10202# a_23350_10202# 0.14fF
C11532 a_25054_2130# rowoff_n[0] 0.10fF
C11533 a_22042_13174# col_n[19] 0.28fF
C11534 a_1962_10202# col_n[9] 0.13fF
C11535 a_32386_15222# vcm 0.22fF
C11536 m2_15788_18014# m3_14916_18146# 0.13fF
C11537 a_33086_17190# row_n[15] 0.17fF
C11538 a_14010_9158# ctop 3.58fF
C11539 a_2966_7150# VDD 0.56fF
C11540 a_1962_4178# col[0] 0.11fF
C11541 m2_1732_1950# rowoff_n[0] 0.12fF
C11542 a_17022_2130# rowon_n[0] 0.14fF
C11543 a_21950_17190# VDD 0.24fF
C11544 a_1962_17230# col[2] 0.11fF
C11545 m2_1732_17010# rowoff_n[15] 0.12fF
C11546 a_2346_3176# col[20] 0.15fF
C11547 a_31990_2130# VDD 0.23fF
C11548 a_2346_16228# col[22] 0.15fF
C11549 a_2346_4180# a_14922_4138# 0.35fF
C11550 a_7986_4138# a_8990_4138# 0.97fF
C11551 a_27062_13174# ctop 3.58fF
C11552 a_4974_6146# col_n[2] 0.28fF
C11553 a_9994_14178# a_9994_13174# 1.00fF
C11554 a_26970_14178# a_27062_14178# 0.26fF
C11555 a_13918_10162# rowoff_n[8] 0.24fF
C11556 m2_34864_5966# m2_34864_4962# 0.99fF
C11557 a_21038_15182# rowon_n[13] 0.14fF
C11558 a_7986_12170# vcm 0.62fF
C11559 a_15926_13174# rowoff_n[11] 0.24fF
C11560 a_10998_5142# VDD 0.52fF
C11561 a_1962_12210# col[29] 0.11fF
C11562 a_2346_6188# a_27974_6146# 0.35fF
C11563 a_23046_2130# col_n[20] 0.28fF
C11564 a_23958_8154# rowoff_n[6] 0.24fF
C11565 m2_11772_946# a_1962_1166# 0.18fF
C11566 a_20034_16186# col[17] 0.29fF
C11567 a_1962_6186# vcm 6.95fF
C11568 a_29982_17190# rowoff_n[15] 0.24fF
C11569 a_21038_16186# vcm 0.62fF
C11570 a_14010_5142# row_n[3] 0.17fF
C11571 a_33998_6146# rowoff_n[4] 0.24fF
C11572 a_1962_3174# a_22042_3134# 0.27fF
C11573 a_1962_1166# m2_28840_946# 0.18fF
C11574 a_24050_9158# VDD 0.52fF
C11575 a_21038_8154# a_22042_8154# 0.97fF
C11576 a_31078_1126# vcm 0.12fF
C11577 a_14314_10202# vcm 0.22fF
C11578 a_1962_17230# a_8290_17230# 0.14fF
C11579 a_2346_17232# a_9994_17190# 0.19fF
C11580 a_2346_12212# col[13] 0.15fF
C11581 m3_17928_18146# ctop 0.23fF
C11582 a_33086_12170# m2_33284_12418# 0.16fF
C11583 a_1962_1166# col_n[27] 0.13fF
C11584 a_1962_14218# col_n[29] 0.13fF
C11585 a_2966_14178# a_3970_14178# 0.97fF
C11586 a_33086_8154# row_n[6] 0.17fF
C11587 a_2874_14178# rowoff_n[12] 0.24fF
C11588 a_27366_14218# vcm 0.22fF
C11589 a_1962_2170# a_28370_2170# 0.14fF
C11590 a_2346_2172# a_30074_2130# 0.19fF
C11591 a_33086_3134# a_33086_2130# 1.00fF
C11592 a_8990_8154# ctop 3.58fF
C11593 a_1962_8194# col[20] 0.11fF
C11594 a_21038_5142# col[18] 0.29fF
C11595 a_16930_16186# VDD 0.23fF
C11596 m2_34864_11990# vcm 0.50fF
C11597 a_5978_2130# m2_6176_2378# 0.16fF
C11598 a_5978_16186# rowon_n[14] 0.14fF
C11599 a_26970_1126# VDD 0.44fF
C11600 a_5978_4138# a_5978_3134# 1.00fF
C11601 a_22954_4138# a_23046_4138# 0.26fF
C11602 a_22042_12170# ctop 3.58fF
C11603 a_21038_6146# rowon_n[4] 0.14fF
C11604 a_6982_13174# a_7986_13174# 0.97fF
C11605 a_2346_13216# a_12914_13174# 0.35fF
C11606 VDD rowon_n[15] 2.78fF
C11607 vcm col_n[28] 2.80fF
C11608 a_2346_8196# col[4] 0.15fF
C11609 col[16] rowoff_n[15] 0.11fF
C11610 a_5978_4138# VDD 0.52fF
C11611 m3_1864_6098# VDD 0.25fF
C11612 a_30074_13174# m2_30272_13422# 0.16fF
C11613 a_1962_10202# a_6982_10162# 0.27fF
C11614 a_1962_10202# col_n[20] 0.13fF
C11615 a_21038_7150# col_n[18] 0.28fF
C11616 a_2346_15224# a_25966_15182# 0.35fF
C11617 a_16018_15182# vcm 0.62fF
C11618 a_1962_4178# col[11] 0.11fF
C11619 a_1962_17230# col[13] 0.11fF
C11620 a_19030_8154# VDD 0.52fF
C11621 a_19030_8154# a_19030_7150# 1.00fF
C11622 a_3878_17190# VDD 0.24fF
C11623 a_1962_12210# a_20034_12170# 0.27fF
C11624 a_2966_14178# col[0] 0.29fF
C11625 m2_1732_2954# sample 0.19fF
C11626 a_2346_3176# col[31] 0.15fF
C11627 a_9294_9198# vcm 0.22fF
C11628 a_20034_17190# a_21038_17190# 0.97fF
C11629 m2_1732_13998# sample_n 0.15fF
C11630 a_2966_3134# m2_3164_3382# 0.16fF
C11631 a_6890_5142# rowoff_n[3] 0.24fF
C11632 a_18026_9158# row_n[7] 0.17fF
C11633 a_32082_12170# VDD 0.52fF
C11634 m3_31984_18146# m3_32988_18146# 0.22fF
C11635 a_2346_9200# a_15014_9158# 0.19fF
C11636 a_8898_9158# a_8990_9158# 0.26fF
C11637 a_1962_9198# a_13310_9198# 0.14fF
C11638 a_1962_14218# a_33086_14178# 0.27fF
C11639 a_16930_3134# rowoff_n[1] 0.24fF
C11640 a_2966_15182# rowon_n[13] 0.13fF
C11641 a_31990_14178# rowoff_n[12] 0.24fF
C11642 a_22346_13214# vcm 0.22fF
C11643 a_30074_2130# a_31078_2130# 0.97fF
C11644 a_3970_7150# ctop 3.57fF
C11645 a_27062_14178# m2_27260_14426# 0.16fF
C11646 a_11910_15182# VDD 0.23fF
C11647 a_1962_6186# col_n[11] 0.13fF
C11648 a_32082_12170# a_32082_11166# 1.00fF
C11649 a_1962_11206# a_26362_11206# 0.14fF
C11650 a_2346_11208# a_28066_11166# 0.19fF
C11651 a_19030_10162# col[16] 0.29fF
C11652 a_5978_7150# rowon_n[5] 0.14fF
C11653 a_2966_16186# vcm 0.61fF
C11654 a_2346_3176# a_4882_3134# 0.35fF
C11655 a_1962_13214# col[4] 0.11fF
C11656 a_17022_11166# ctop 3.58fF
C11657 a_21950_13174# a_22042_13174# 0.26fF
C11658 a_4974_13174# a_4974_12170# 1.00fF
C11659 a_2346_12212# col[24] 0.15fF
C11660 a_4974_11166# rowoff_n[9] 0.10fF
C11661 a_34090_5142# m2_34864_4962# 0.96fF
C11662 a_35002_4138# VDD 0.29fF
C11663 m2_21812_946# vcm 0.42fF
C11664 a_2346_5184# a_17934_5142# 0.35fF
C11665 a_30074_15182# ctop 3.58fF
C11666 a_1962_10202# a_34394_10202# 0.14fF
C11667 a_25054_10162# rowon_n[8] 0.14fF
C11668 a_15014_9158# rowoff_n[7] 0.10fF
C11669 a_2966_15182# m3_1864_15134# 0.14fF
C11670 a_1962_8194# col[31] 0.11fF
C11671 a_19030_15182# rowoff_n[13] 0.10fF
C11672 a_10998_14178# vcm 0.62fF
C11673 a_19030_12170# col_n[16] 0.28fF
C11674 a_1962_2170# a_12002_2130# 0.27fF
C11675 m2_29844_18014# m3_29976_18146# 2.78fF
C11676 a_14010_7150# VDD 0.52fF
C11677 a_25054_7150# rowoff_n[5] 0.10fF
C11678 a_16018_7150# a_17022_7150# 0.97fF
C11679 a_2346_7192# a_30986_7150# 0.35fF
C11680 a_24050_15182# m2_24248_15430# 0.16fF
C11681 a_1962_2170# col_n[2] 0.13fF
C11682 a_1962_15222# col_n[4] 0.13fF
C11683 a_4274_8194# vcm 0.22fF
C11684 a_18026_17190# a_18026_16186# 1.00fF
C11685 a_26058_3134# m2_26256_3382# 0.16fF
C11686 a_24050_18194# vcm 0.12fF
C11687 a_1962_4178# a_25054_4138# 0.27fF
C11688 a_27062_11166# VDD 0.52fF
C11689 m3_21944_1078# m3_22948_1078# 0.22fF
C11690 a_2346_18236# VDD 33.26fF
C11691 a_2966_6146# rowon_n[4] 0.13fF
C11692 a_34090_3134# vcm 0.62fF
C11693 col_n[19] col_n[20] 0.10fF
C11694 col_n[2] row_n[13] 0.23fF
C11695 col_n[6] row_n[15] 0.23fF
C11696 sample row_n[11] 1.03fF
C11697 VDD row_n[10] 2.93fF
C11698 col_n[4] row_n[14] 0.23fF
C11699 vcm row_n[12] 0.49fF
C11700 a_2346_8196# col[15] 0.15fF
C11701 col[27] rowoff_n[15] 0.11fF
C11702 col[29] col[30] 0.20fF
C11703 a_17326_12210# vcm 0.22fF
C11704 a_1962_1166# a_18330_1166# 0.19fF
C11705 a_2346_1168# a_20034_1126# 0.19fF
C11706 a_22042_13174# row_n[11] 0.17fF
C11707 a_1962_10202# col_n[31] 0.13fF
C11708 a_6890_14178# VDD 0.23fF
C11709 a_29070_11166# a_30074_11166# 0.97fF
C11710 a_20034_1126# col_n[17] 0.31fF
C11711 a_1962_4178# col[22] 0.11fF
C11712 a_1962_17230# col[24] 0.11fF
C11713 a_6890_16186# rowoff_n[14] 0.24fF
C11714 a_30378_16226# vcm 0.22fF
C11715 a_17022_15182# col[14] 0.29fF
C11716 m2_15788_946# m2_16792_946# 0.96fF
C11717 a_17934_3134# a_18026_3134# 0.26fF
C11718 a_2346_3176# a_33086_3134# 0.19fF
C11719 a_1962_8194# m2_1732_7974# 0.15fF
C11720 a_1962_3174# a_31382_3174# 0.14fF
C11721 a_12002_10162# ctop 3.58fF
C11722 a_21038_16186# m2_21236_16434# 0.16fF
C11723 a_19942_18194# VDD 0.33fF
C11724 m2_14784_18014# vcm 0.28fF
C11725 a_9994_11166# rowon_n[9] 0.14fF
C11726 a_33998_11166# rowoff_n[9] 0.24fF
C11727 a_23046_4138# m2_23244_4386# 0.16fF
C11728 a_29982_3134# VDD 0.23fF
C11729 m3_34996_5094# ctop 0.23fF
C11730 a_25054_14178# ctop 3.58fF
C11731 m2_32856_946# m2_33860_946# 0.93fF
C11732 a_2346_4180# col[6] 0.15fF
C11733 a_2346_14220# a_15926_14178# 0.35fF
C11734 a_2346_17232# col[8] 0.15fF
C11735 a_2346_18236# a_24962_18194# 0.35fF
C11736 a_5978_13174# vcm 0.62fF
C11737 a_1962_6186# col_n[22] 0.13fF
C11738 a_8990_6146# VDD 0.52fF
C11739 a_30986_7150# a_31078_7150# 0.26fF
C11740 a_14010_7150# a_14010_6146# 1.00fF
C11741 a_17022_17190# col_n[14] 0.28fF
C11742 a_29070_14178# rowon_n[12] 0.14fF
C11743 a_1962_11206# a_9994_11166# 0.27fF
C11744 a_18026_4138# col[15] 0.29fF
C11745 a_2346_16228# a_28978_16186# 0.35fF
C11746 a_15014_16186# a_16018_16186# 0.97fF
C11747 a_1962_13214# col[15] 0.11fF
C11748 a_19030_17190# vcm 0.60fF
C11749 rowon_n[6] rowoff_n[6] 20.27fF
C11750 m2_5748_18014# VDD 0.93fF
C11751 a_1962_18234# m2_20808_18014# 0.18fF
C11752 a_22042_10162# VDD 0.52fF
C11753 a_2346_8196# a_4974_8154# 0.19fF
C11754 a_1962_8194# a_3270_8194# 0.14fF
C11755 a_18026_17190# m2_18224_17438# 0.16fF
C11756 a_6982_14178# row_n[12] 0.17fF
C11757 a_29070_2130# vcm 0.62fF
C11758 a_1962_13214# a_23046_13174# 0.27fF
C11759 a_21038_12170# rowoff_n[10] 0.10fF
C11760 a_7986_4138# rowoff_n[2] 0.10fF
C11761 a_12306_11206# vcm 0.22fF
C11762 a_22042_4138# row_n[2] 0.17fF
C11763 a_20034_5142# m2_20232_5390# 0.16fF
C11764 a_2346_18236# m2_15788_18014# 0.19fF
C11765 a_1962_10202# a_16322_10202# 0.14fF
C11766 a_27062_11166# a_27062_10162# 1.00fF
C11767 a_2346_10204# a_18026_10162# 0.19fF
C11768 a_18026_2130# rowoff_n[0] 0.10fF
C11769 a_25358_15222# vcm 0.22fF
C11770 a_18026_6146# col_n[15] 0.28fF
C11771 a_1962_2170# col_n[13] 0.13fF
C11772 a_6982_9158# ctop 3.58fF
C11773 a_18026_1126# m3_16924_1078# 0.14fF
C11774 m2_5748_18014# m3_6884_18146# 0.13fF
C11775 a_26058_17190# row_n[15] 0.17fF
C11776 a_1962_15222# col_n[15] 0.13fF
C11777 a_9994_2130# rowon_n[0] 0.14fF
C11778 a_14922_17190# VDD 0.24fF
C11779 m2_1732_15002# vcm 0.45fF
C11780 a_2346_12212# a_31078_12170# 0.19fF
C11781 a_16930_12170# a_17022_12170# 0.26fF
C11782 a_1962_12210# a_29374_12210# 0.14fF
C11783 a_1962_9198# col[6] 0.11fF
C11784 a_24962_2130# VDD 0.23fF
C11785 a_2346_4180# a_7894_4138# 0.35fF
C11786 a_33086_16186# col[30] 0.29fF
C11787 a_20034_13174# ctop 3.58fF
C11788 m3_34996_9110# m3_34996_8106# 0.22fF
C11789 col_n[0] row_n[6] 0.23fF
C11790 col_n[7] row_n[10] 0.23fF
C11791 vcm rowon_n[6] 0.50fF
C11792 col_n[5] row_n[9] 0.23fF
C11793 col_n[11] row_n[12] 0.23fF
C11794 col_n[9] row_n[11] 0.23fF
C11795 col_n[1] row_n[7] 0.23fF
C11796 VDD rowon_n[4] 2.61fF
C11797 col_n[15] row_n[14] 0.23fF
C11798 col_n[17] row_n[15] 0.23fF
C11799 col_n[13] row_n[13] 0.23fF
C11800 col_n[3] row_n[8] 0.23fF
C11801 a_2346_8196# col[26] 0.15fF
C11802 a_6890_10162# rowoff_n[8] 0.24fF
C11803 a_14010_15182# rowon_n[13] 0.14fF
C11804 a_8898_13174# rowoff_n[11] 0.24fF
C11805 m2_34864_2954# VDD 1.00fF
C11806 a_17022_6146# m2_17220_6394# 0.16fF
C11807 a_3970_5142# VDD 0.52fF
C11808 a_29070_5142# rowon_n[3] 0.14fF
C11809 a_10998_6146# a_12002_6146# 0.97fF
C11810 a_2346_6188# a_20946_6146# 0.35fF
C11811 a_33086_17190# ctop 3.38fF
C11812 a_16930_8154# rowoff_n[6] 0.24fF
C11813 a_13006_17190# m3_12908_18146# 0.15fF
C11814 a_29982_16186# a_30074_16186# 0.26fF
C11815 a_13006_16186# a_13006_15182# 1.00fF
C11816 a_1962_1166# m2_4744_946# 0.18fF
C11817 a_22954_17190# rowoff_n[15] 0.24fF
C11818 a_14010_16186# vcm 0.62fF
C11819 a_16018_9158# col[13] 0.29fF
C11820 a_26970_6146# rowoff_n[4] 0.24fF
C11821 a_6982_5142# row_n[3] 0.17fF
C11822 a_1962_3174# a_15014_3134# 0.27fF
C11823 a_1962_11206# col_n[6] 0.13fF
C11824 a_17022_9158# VDD 0.52fF
C11825 a_2346_8196# a_33998_8154# 0.35fF
C11826 m2_12776_946# ctop 0.18fF
C11827 a_24050_1126# vcm 0.12fF
C11828 m2_16792_18014# col[14] 0.28fF
C11829 a_34090_5142# col[31] 0.29fF
C11830 a_7286_10202# vcm 0.22fF
C11831 a_2346_17232# a_2874_17190# 0.35fF
C11832 m2_29844_946# ctop 0.18fF
C11833 a_1962_5182# a_28066_5142# 0.27fF
C11834 a_30074_13174# VDD 0.52fF
C11835 a_2346_4180# col[17] 0.15fF
C11836 a_24050_10162# a_25054_10162# 0.97fF
C11837 a_2346_17232# col[19] 0.15fF
C11838 a_26058_8154# row_n[6] 0.17fF
C11839 a_20338_14218# vcm 0.22fF
C11840 a_2346_2172# a_23046_2130# 0.19fF
C11841 a_14010_7150# m2_14208_7398# 0.16fF
C11842 a_12914_2130# a_13006_2130# 0.26fF
C11843 a_1962_2170# a_21342_2170# 0.14fF
C11844 a_16018_11166# col_n[13] 0.28fF
C11845 a_9902_16186# VDD 0.23fF
C11846 a_1962_13214# col[26] 0.11fF
C11847 m2_6752_946# col[4] 0.39fF
C11848 a_35002_3134# m2_34864_2954# 0.16fF
C11849 a_33390_18234# vcm 0.22fF
C11850 a_19942_1126# VDD 0.39fF
C11851 m2_32856_18014# col_n[30] 0.25fF
C11852 a_34090_7150# col_n[31] 0.28fF
C11853 a_2346_4180# a_2346_3176# 0.22fF
C11854 a_1962_4178# a_35398_4178# 0.14fF
C11855 a_15014_12170# ctop 3.58fF
C11856 a_15014_17190# m2_14784_18014# 1.00fF
C11857 a_14010_6146# rowon_n[4] 0.14fF
C11858 a_2346_13216# a_5886_13174# 0.35fF
C11859 a_2966_12170# rowoff_n[10] 0.10fF
C11860 a_32994_5142# VDD 0.23fF
C11861 a_8990_6146# a_8990_5142# 1.00fF
C11862 a_25966_6146# a_26058_6146# 0.26fF
C11863 m3_29976_18146# VDD 0.25fF
C11864 a_28066_16186# ctop 3.57fF
C11865 a_2346_13216# col[10] 0.15fF
C11866 m2_20808_946# a_20946_1126# 0.16fF
C11867 a_9994_15182# a_10998_15182# 0.97fF
C11868 a_2346_15224# a_18938_15182# 0.35fF
C11869 a_1962_2170# col_n[24] 0.13fF
C11870 a_1962_15222# col_n[26] 0.13fF
C11871 a_8990_15182# vcm 0.62fF
C11872 a_10998_8154# m2_11196_8402# 0.16fF
C11873 a_33086_9158# rowon_n[7] 0.14fF
C11874 a_12002_8154# VDD 0.52fF
C11875 a_14010_14178# col[11] 0.29fF
C11876 a_1962_9198# col[17] 0.11fF
C11877 a_1962_12210# a_13006_12170# 0.27fF
C11878 a_2346_17232# a_31990_17190# 0.35fF
C11879 m2_6752_946# m3_5880_1078# 0.13fF
C11880 VDD sw_n 0.25fF
C11881 col_n[10] row_n[6] 0.23fF
C11882 col_n[26] row_n[14] 0.23fF
C11883 sample row_n[0] 1.03fF
C11884 col_n[4] row_n[3] 0.23fF
C11885 col_n[22] row_n[12] 0.23fF
C11886 col_n[16] row_n[9] 0.23fF
C11887 col_n[6] row_n[4] 0.23fF
C11888 a_10998_9158# row_n[7] 0.17fF
C11889 col_n[24] row_n[13] 0.23fF
C11890 col_n[20] row_n[11] 0.23fF
C11891 col_n[28] row_n[15] 0.23fF
C11892 col_n[12] row_n[7] 0.23fF
C11893 col_n[8] row_n[5] 0.23fF
C11894 col_n[18] row_n[10] 0.23fF
C11895 col_n[2] row_n[2] 0.23fF
C11896 col_n[30] col_n[31] 0.12fF
C11897 vcm row_n[1] 0.49fF
C11898 a_32082_10162# col[29] 0.29fF
C11899 col_n[14] row_n[8] 0.23fF
C11900 a_25054_12170# VDD 0.52fF
C11901 m3_17928_18146# m3_18932_18146# 0.22fF
C11902 a_2346_9200# a_7986_9158# 0.19fF
C11903 a_1962_9198# a_6282_9198# 0.14fF
C11904 a_22042_10162# a_22042_9158# 1.00fF
C11905 a_32082_4138# vcm 0.62fF
C11906 a_1962_14218# a_26058_14178# 0.27fF
C11907 a_9902_3134# rowoff_n[1] 0.24fF
C11908 a_15318_13214# vcm 0.22fF
C11909 a_24962_14178# rowoff_n[12] 0.24fF
C11910 a_2966_6146# m2_1732_5966# 0.96fF
C11911 a_2346_6188# a_1962_6186# 2.62fF
C11912 a_2346_9200# col[1] 0.15fF
C11913 a_34090_9158# m3_34996_9110# 0.13fF
C11914 a_4882_15182# VDD 0.23fF
C11915 a_2346_11208# a_21038_11166# 0.19fF
C11916 a_11910_11166# a_12002_11166# 0.26fF
C11917 a_1962_11206# a_19334_11206# 0.14fF
C11918 a_14010_16186# col_n[11] 0.28fF
C11919 a_1962_18234# vcm 7.34fF
C11920 a_1962_11206# col_n[17] 0.13fF
C11921 a_30074_12170# row_n[10] 0.17fF
C11922 a_15014_3134# col[12] 0.29fF
C11923 a_28370_17230# vcm 0.22fF
C11924 a_33086_4138# a_34090_4138# 0.97fF
C11925 a_7986_9158# m2_8184_9406# 0.16fF
C11926 a_9994_11166# ctop 3.58fF
C11927 a_34090_17190# m2_33860_18014# 1.00fF
C11928 a_1962_5182# col[8] 0.11fF
C11929 a_32082_12170# col_n[29] 0.28fF
C11930 a_2346_13216# a_34090_13174# 0.19fF
C11931 a_1962_13214# a_32386_13214# 0.14fF
C11932 a_2346_4180# col[28] 0.15fF
C11933 a_27974_4138# VDD 0.23fF
C11934 a_2346_5184# a_10906_5142# 0.35fF
C11935 a_2346_17232# col[30] 0.15fF
C11936 a_5978_5142# a_6982_5142# 0.97fF
C11937 a_23046_15182# ctop 3.58fF
C11938 a_18026_10162# rowon_n[8] 0.14fF
C11939 a_7986_9158# rowoff_n[7] 0.10fF
C11940 a_24962_15182# a_25054_15182# 0.26fF
C11941 a_7986_15182# a_7986_14178# 1.00fF
C11942 m2_1732_8978# m2_1732_7974# 0.99fF
C11943 a_12002_15182# rowoff_n[13] 0.10fF
C11944 a_3970_14178# vcm 0.62fF
C11945 a_3878_2130# a_3970_2130# 0.26fF
C11946 a_1962_2170# a_4974_2130# 0.27fF
C11947 m2_20808_18014# m3_19936_18146# 0.13fF
C11948 vcm rowoff_n[13] 0.20fF
C11949 a_6982_7150# VDD 0.52fF
C11950 a_18026_7150# rowoff_n[5] 0.10fF
C11951 a_2346_7192# a_23958_7150# 0.35fF
C11952 a_15014_5142# col_n[12] 0.28fF
C11953 ctop rowoff_n[0] 0.51fF
C11954 col[2] rowoff_n[8] 0.11fF
C11955 col[1] rowoff_n[7] 0.11fF
C11956 col[3] rowoff_n[9] 0.11fF
C11957 col[0] rowoff_n[6] 0.11fF
C11958 a_1962_7190# col_n[8] 0.13fF
C11959 a_28066_5142# rowoff_n[3] 0.10fF
C11960 a_17022_18194# vcm 0.12fF
C11961 a_35494_2492# VDD 0.11fF
C11962 a_1962_4178# a_18026_4138# 0.27fF
C11963 a_4974_10162# m2_5172_10410# 0.16fF
C11964 a_20034_11166# VDD 0.52fF
C11965 m3_7888_1078# m3_8892_1078# 0.22fF
C11966 a_19030_9158# a_20034_9158# 0.97fF
C11967 a_2966_17190# m2_2736_18014# 1.00fF
C11968 a_1962_9198# a_1962_8194# 0.16fF
C11969 a_1962_14218# col[1] 0.11fF
C11970 a_30074_15182# col[27] 0.29fF
C11971 a_27062_3134# vcm 0.62fF
C11972 a_10298_12210# vcm 0.22fF
C11973 a_1962_1166# a_11302_1166# 0.14fF
C11974 a_2346_13216# col[21] 0.15fF
C11975 a_15014_13174# row_n[11] 0.17fF
C11976 a_1962_6186# a_31078_6146# 0.27fF
C11977 a_33086_15182# VDD 0.52fF
C11978 m2_20808_946# a_1962_1166# 0.18fF
C11979 a_30074_3134# row_n[1] 0.17fF
C11980 a_1962_15222# row_n[13] 25.57fF
C11981 a_10906_1126# m2_10768_946# 0.16fF
C11982 a_23350_16226# vcm 0.22fF
C11983 a_31078_4138# a_31078_3134# 1.00fF
C11984 a_2346_3176# a_26058_3134# 0.19fF
C11985 a_1962_3174# a_24354_3174# 0.14fF
C11986 a_4974_10162# ctop 3.58fF
C11987 a_1962_9198# col[28] 0.11fF
C11988 a_13006_8154# col[10] 0.29fF
C11989 a_12914_18194# VDD 0.33fF
C11990 a_35398_1166# vcm 0.23fF
C11991 a_32082_13174# a_33086_13174# 0.97fF
C11992 a_1962_3174# col_n[0] 0.13fF
C11993 a_26970_11166# rowoff_n[9] 0.24fF
C11994 col_n[19] row_n[5] 0.23fF
C11995 col_n[31] row_n[11] 0.23fF
C11996 col_n[29] row_n[10] 0.23fF
C11997 vcm col[0] 5.82fF
C11998 col_n[23] row_n[7] 0.23fF
C11999 col_n[13] row_n[2] 0.23fF
C12000 col_n[11] row_n[1] 0.23fF
C12001 col_n[21] row_n[6] 0.23fF
C12002 col_n[27] row_n[9] 0.23fF
C12003 col_n[6] ctop 2.02fF
C12004 col_n[25] row_n[8] 0.23fF
C12005 col_n[15] row_n[3] 0.23fF
C12006 col_n[17] row_n[4] 0.23fF
C12007 col_n[9] row_n[0] 0.23fF
C12008 col_n[0] col[1] 6.01fF
C12009 VDD col[4] 4.17fF
C12010 a_30074_17190# col_n[27] 0.28fF
C12011 a_1962_16226# col_n[1] 0.13fF
C12012 a_34090_16186# row_n[14] 0.17fF
C12013 a_22954_3134# VDD 0.23fF
C12014 a_31078_4138# col[28] 0.29fF
C12015 m3_32988_18146# ctop 0.23fF
C12016 a_20946_5142# a_21038_5142# 0.26fF
C12017 a_3970_5142# a_3970_4138# 1.00fF
C12018 a_18026_14178# ctop 3.58fF
C12019 m2_25828_946# m2_26832_946# 0.96fF
C12020 a_2346_14220# a_8898_14178# 0.35fF
C12021 a_4974_14178# a_5978_14178# 0.97fF
C12022 a_2346_18236# a_17934_18194# 0.35fF
C12023 m2_1732_5966# VDD 1.02fF
C12024 a_2346_9200# col[12] 0.15fF
C12025 a_1962_18234# col_n[11] 0.13fF
C12026 a_22042_14178# rowon_n[12] 0.14fF
C12027 a_2346_11208# a_2966_11166# 0.21fF
C12028 a_1962_11206# col_n[28] 0.13fF
C12029 a_13006_10162# col_n[10] 0.28fF
C12030 a_2346_16228# a_21950_16186# 0.35fF
C12031 a_2346_2172# m2_34864_1950# 0.17fF
C12032 a_8990_2130# m2_9188_2378# 0.16fF
C12033 a_12002_17190# vcm 0.60fF
C12034 a_1962_18234# m2_6752_18014# 0.18fF
C12035 a_1962_5182# col[19] 0.11fF
C12036 a_15014_10162# VDD 0.52fF
C12037 a_33998_9158# a_34090_9158# 0.26fF
C12038 a_17022_9158# a_17022_8154# 1.00fF
C12039 a_31078_6146# col_n[28] 0.28fF
C12040 a_22042_2130# vcm 0.62fF
C12041 a_1962_13214# a_16018_13174# 0.27fF
C12042 a_15014_4138# row_n[2] 0.17fF
C12043 a_14010_12170# rowoff_n[10] 0.10fF
C12044 a_5278_11206# vcm 0.22fF
C12045 m3_5880_1078# VDD 0.14fF
C12046 a_33086_13174# m2_33284_13422# 0.16fF
C12047 a_2346_18236# m2_1732_18014# 0.12fF
C12048 a_28066_14178# VDD 0.52fF
C12049 a_1962_6186# row_n[4] 25.57fF
C12050 a_6890_10162# a_6982_10162# 0.26fF
C12051 a_2346_10204# a_10998_10162# 0.19fF
C12052 a_1962_10202# a_9294_10202# 0.14fF
C12053 a_10998_2130# rowoff_n[0] 0.10fF
C12054 a_35094_6146# vcm 0.12fF
C12055 a_1962_15222# a_29070_15182# 0.27fF
C12056 m2_28840_18014# ctop 0.18fF
C12057 a_18330_15222# vcm 0.22fF
C12058 a_28066_16186# rowoff_n[14] 0.10fF
C12059 a_2346_5184# col[3] 0.15fF
C12060 a_28066_3134# a_29070_3134# 0.97fF
C12061 a_19030_17190# row_n[15] 0.17fF
C12062 col[7] rowoff_n[2] 0.11fF
C12063 col[11] rowoff_n[6] 0.11fF
C12064 col[12] rowoff_n[7] 0.11fF
C12065 col[5] rowoff_n[0] 0.11fF
C12066 col[6] rowoff_n[1] 0.11fF
C12067 col[13] rowoff_n[8] 0.11fF
C12068 col[8] rowoff_n[3] 0.11fF
C12069 col[14] rowoff_n[9] 0.11fF
C12070 col[9] rowoff_n[4] 0.11fF
C12071 col[10] rowoff_n[5] 0.11fF
C12072 a_7894_17190# VDD 0.24fF
C12073 a_30074_13174# a_30074_12170# 1.00fF
C12074 a_2346_12212# a_24050_12170# 0.19fF
C12075 a_1962_7190# col_n[19] 0.13fF
C12076 a_1962_12210# a_22346_12210# 0.14fF
C12077 a_34090_7150# row_n[5] 0.17fF
C12078 a_10998_13174# col[8] 0.29fF
C12079 m2_15788_946# m3_16924_1078# 0.13fF
C12080 a_17934_2130# VDD 0.23fF
C12081 a_1962_1166# col[10] 0.11fF
C12082 a_1962_14218# col[12] 0.11fF
C12083 a_13006_13174# ctop 3.58fF
C12084 m2_27836_946# m3_26964_1078# 0.13fF
C12085 m3_34996_16138# m3_34996_15134# 0.22fF
C12086 a_13918_18194# m2_13780_18014# 0.16fF
C12087 a_29070_9158# col[26] 0.29fF
C12088 a_19942_14178# a_20034_14178# 0.26fF
C12089 a_6982_15182# rowon_n[13] 0.14fF
C12090 a_30986_6146# VDD 0.23fF
C12091 a_22042_5142# rowon_n[3] 0.14fF
C12092 a_30074_14178# m2_30272_14426# 0.16fF
C12093 a_2346_6188# a_13918_6146# 0.35fF
C12094 a_26058_17190# ctop 3.39fF
C12095 a_9902_8154# rowoff_n[6] 0.24fF
C12096 a_2346_1168# ctop 0.38fF
C12097 a_15926_17190# rowoff_n[15] 0.24fF
C12098 a_6982_16186# vcm 0.62fF
C12099 a_10998_15182# col_n[8] 0.28fF
C12100 a_1962_3174# a_7986_3134# 0.27fF
C12101 a_19942_6146# rowoff_n[4] 0.24fF
C12102 a_12002_2130# col[9] 0.29fF
C12103 a_9994_9158# VDD 0.52fF
C12104 a_14010_8154# a_15014_8154# 0.97fF
C12105 a_2346_8196# a_26970_8154# 0.35fF
C12106 a_1962_3174# col_n[10] 0.13fF
C12107 col_n[20] row_n[0] 0.23fF
C12108 col_n[17] ctop 2.01fF
C12109 col_n[30] row_n[5] 0.23fF
C12110 col_n[15] en_bit_n[1] 0.17fF
C12111 a_17022_1126# vcm 0.12fF
C12112 col_n[26] row_n[3] 0.23fF
C12113 col_n[22] row_n[1] 0.23fF
C12114 col_n[28] row_n[4] 0.23fF
C12115 vcm col[11] 5.84fF
C12116 col_n[24] row_n[2] 0.23fF
C12117 VDD col[15] 4.17fF
C12118 col_n[5] col[6] 5.98fF
C12119 a_1962_16226# col_n[12] 0.13fF
C12120 m2_5748_946# ctop 0.18fF
C12121 a_29070_11166# col_n[26] 0.28fF
C12122 a_29982_4138# rowoff_n[2] 0.24fF
C12123 a_2966_4138# m2_3164_4386# 0.16fF
C12124 a_2966_13174# col_n[0] 0.28fF
C12125 a_1962_10202# col[3] 0.11fF
C12126 a_1962_5182# a_21038_5142# 0.27fF
C12127 a_23046_13174# VDD 0.52fF
C12128 a_30074_5142# vcm 0.62fF
C12129 a_2346_9200# col[23] 0.15fF
C12130 a_19030_8154# row_n[6] 0.17fF
C12131 a_13310_14218# vcm 0.22fF
C12132 a_1962_2170# a_14314_2170# 0.14fF
C12133 a_26058_3134# a_26058_2130# 1.00fF
C12134 a_2346_2172# a_16018_2130# 0.19fF
C12135 m2_34864_18014# m3_34996_18146# 2.78fF
C12136 a_1962_18234# col_n[22] 0.13fF
C12137 a_1962_7190# a_34090_7150# 0.27fF
C12138 a_27062_15182# m2_27260_15430# 0.16fF
C12139 a_2346_16228# VDD 32.63fF
C12140 a_27062_12170# a_28066_12170# 0.97fF
C12141 a_12002_4138# col_n[9] 0.28fF
C12142 rowon_n[12] rowoff_n[12] 20.27fF
C12143 a_2874_16186# a_2966_16186# 0.26fF
C12144 a_2346_16228# a_3878_16186# 0.35fF
C12145 a_29070_3134# m2_29268_3382# 0.16fF
C12146 a_1962_5182# col[30] 0.11fF
C12147 a_26362_18234# vcm 0.22fF
C12148 a_12914_1126# VDD 0.44fF
C12149 a_1962_4178# a_27366_4178# 0.14fF
C12150 a_2346_4180# a_29070_4138# 0.19fF
C12151 a_15926_4138# a_16018_4138# 0.26fF
C12152 a_7986_12170# ctop 3.58fF
C12153 m2_29844_946# col[27] 0.39fF
C12154 a_32994_18194# m2_32856_18014# 0.16fF
C12155 a_6982_6146# rowon_n[4] 0.14fF
C12156 a_1962_12210# col_n[3] 0.13fF
C12157 a_28066_10162# rowoff_n[8] 0.10fF
C12158 a_27062_14178# col[24] 0.29fF
C12159 a_30074_13174# rowoff_n[11] 0.10fF
C12160 a_34090_6146# m2_34864_5966# 0.96fF
C12161 a_1962_6186# ctop 1.49fF
C12162 a_25966_5142# VDD 0.23fF
C12163 m3_1864_18146# VDD 0.30fF
C12164 a_21038_16186# ctop 3.57fF
C12165 a_2346_15224# a_11910_15182# 0.35fF
C12166 a_2346_5184# col[14] 0.15fF
C12167 col[22] rowoff_n[6] 0.11fF
C12168 col[21] rowoff_n[5] 0.11fF
C12169 a_34394_16226# vcm 0.22fF
C12170 col[16] rowoff_n[0] 0.11fF
C12171 col[23] rowoff_n[7] 0.11fF
C12172 col[24] rowoff_n[8] 0.11fF
C12173 col[17] rowoff_n[1] 0.11fF
C12174 col[18] rowoff_n[2] 0.11fF
C12175 col[25] rowoff_n[9] 0.11fF
C12176 col[19] rowoff_n[3] 0.11fF
C12177 col[20] rowoff_n[4] 0.11fF
C12178 a_26058_9158# rowon_n[7] 0.14fF
C12179 a_4974_8154# VDD 0.52fF
C12180 a_1962_7190# col_n[30] 0.13fF
C12181 a_12002_8154# a_12002_7150# 1.00fF
C12182 a_24050_16186# m2_24248_16434# 0.16fF
C12183 a_28978_8154# a_29070_8154# 0.26fF
C12184 a_1962_12210# a_5978_12170# 0.27fF
C12185 a_1962_18234# a_29374_18234# 0.14fF
C12186 a_9994_7150# col[7] 0.29fF
C12187 a_2346_17232# a_24962_17190# 0.35fF
C12188 a_13006_17190# a_14010_17190# 0.97fF
C12189 a_1962_1166# col[21] 0.11fF
C12190 a_1962_14218# col[23] 0.11fF
C12191 a_26058_4138# m2_26256_4386# 0.16fF
C12192 m2_31852_18014# m2_32856_18014# 0.96fF
C12193 m3_8892_1078# ctop 0.23fF
C12194 a_3970_9158# row_n[7] 0.17fF
C12195 a_27062_16186# col_n[24] 0.28fF
C12196 a_18026_12170# VDD 0.52fF
C12197 m3_3872_18146# m3_4876_18146# 0.22fF
C12198 a_28066_3134# col[25] 0.29fF
C12199 a_25054_4138# vcm 0.62fF
C12200 a_1962_14218# a_19030_14178# 0.27fF
C12201 a_2346_3176# rowoff_n[1] 4.09fF
C12202 col[9] rowoff_n[10] 0.11fF
C12203 m2_34864_11990# ctop 0.17fF
C12204 a_17934_14178# rowoff_n[12] 0.24fF
C12205 a_8290_13214# vcm 0.22fF
C12206 a_23046_2130# a_24050_2130# 0.97fF
C12207 m2_34864_15002# m3_34996_15134# 2.76fF
C12208 a_31078_16186# VDD 0.52fF
C12209 a_2346_11208# a_14010_11166# 0.19fF
C12210 a_1962_11206# a_12306_11206# 0.14fF
C12211 a_25054_12170# a_25054_11166# 1.00fF
C12212 a_2346_1168# col[5] 0.14fF
C12213 a_1962_16226# a_32082_16186# 0.27fF
C12214 a_2346_14220# col[7] 0.15fF
C12215 a_23046_12170# row_n[10] 0.17fF
C12216 m2_34864_13998# m2_35292_14426# 0.16fF
C12217 a_21342_17230# vcm 0.22fF
C12218 a_9994_9158# col_n[7] 0.28fF
C12219 a_1962_9198# m2_1732_8978# 0.15fF
C12220 a_1962_3174# col_n[21] 0.13fF
C12221 rowon_n[8] rowon_n[7] 0.15fF
C12222 col_n[11] col[11] 0.72fF
C12223 a_1962_16226# col_n[23] 0.13fF
C12224 col_n[31] row_n[0] 0.22fF
C12225 col_n[28] ctop 2.02fF
C12226 vcm col[22] 5.84fF
C12227 VDD col[26] 4.17fF
C12228 a_21038_17190# m2_21236_17438# 0.16fF
C12229 a_31382_2170# vcm 0.22fF
C12230 a_1962_13214# a_25358_13214# 0.14fF
C12231 a_2346_13216# a_27062_13174# 0.19fF
C12232 a_14922_13174# a_15014_13174# 0.26fF
C12233 a_28066_5142# col_n[25] 0.28fF
C12234 a_1962_10202# col[14] 0.11fF
C12235 a_23046_5142# m2_23244_5390# 0.16fF
C12236 m2_34864_13998# row_n[12] 0.15fF
C12237 a_20946_4138# VDD 0.23fF
C12238 a_1962_5182# a_2966_5142# 0.27fF
C12239 a_16018_15182# ctop 3.58fF
C12240 a_10998_10162# rowon_n[8] 0.14fF
C12241 a_4974_15182# rowoff_n[13] 0.10fF
C12242 m2_10768_18014# m3_11904_18146# 0.13fF
C12243 a_33998_8154# VDD 0.23fF
C12244 a_10998_7150# rowoff_n[5] 0.10fF
C12245 a_2346_7192# a_16930_7150# 0.35fF
C12246 a_8990_7150# a_9994_7150# 0.97fF
C12247 a_27974_17190# a_28066_17190# 0.26fF
C12248 a_10998_17190# a_10998_16186# 1.00fF
C12249 a_21038_5142# rowoff_n[3] 0.10fF
C12250 a_7986_12170# col[5] 0.29fF
C12251 a_9994_18194# vcm 0.12fF
C12252 a_1962_4178# a_10998_4138# 0.27fF
C12253 a_1962_12210# col_n[14] 0.13fF
C12254 a_30074_13174# rowon_n[11] 0.14fF
C12255 a_13006_11166# VDD 0.52fF
C12256 a_2346_9200# a_29982_9158# 0.35fF
C12257 a_20034_3134# vcm 0.62fF
C12258 a_31078_3134# rowoff_n[1] 0.10fF
C12259 a_26058_8154# col[23] 0.29fF
C12260 a_1962_6186# col[5] 0.11fF
C12261 a_3270_12210# vcm 0.22fF
C12262 a_1962_1166# a_4274_1166# 0.19fF
C12263 a_20034_6146# m2_20232_6394# 0.16fF
C12264 m2_34864_11990# m3_34996_12122# 2.76fF
C12265 a_7986_13174# row_n[11] 0.17fF
C12266 a_1962_6186# a_24050_6146# 0.27fF
C12267 a_2966_16186# ctop 3.41fF
C12268 a_26058_15182# VDD 0.52fF
C12269 a_2346_5184# col[25] 0.15fF
C12270 a_22042_11166# a_23046_11166# 0.97fF
C12271 a_23046_3134# row_n[1] 0.17fF
C12272 a_16018_17190# m3_15920_18146# 0.15fF
C12273 col[29] rowoff_n[2] 0.11fF
C12274 col[31] rowoff_n[4] 0.11fF
C12275 col[28] rowoff_n[1] 0.11fF
C12276 col[30] rowoff_n[3] 0.11fF
C12277 col[27] rowoff_n[0] 0.11fF
C12278 a_33086_7150# vcm 0.62fF
C12279 a_16322_16226# vcm 0.22fF
C12280 a_2346_3176# a_19030_3134# 0.19fF
C12281 a_1962_3174# a_17326_3174# 0.14fF
C12282 a_10906_3134# a_10998_3134# 0.26fF
C12283 a_7986_14178# col_n[5] 0.28fF
C12284 m2_21812_946# ctop 0.18fF
C12285 a_5886_18194# VDD 0.33fF
C12286 a_26362_1166# vcm 0.23fF
C12287 m2_8760_946# m2_9764_946# 0.96fF
C12288 a_19942_11166# rowoff_n[9] 0.24fF
C12289 a_27062_16186# row_n[14] 0.17fF
C12290 a_15926_3134# VDD 0.23fF
C12291 a_26058_10162# col_n[23] 0.28fF
C12292 m3_4876_18146# ctop 0.23fF
C12293 a_1962_8194# col_n[5] 0.13fF
C12294 a_1962_5182# a_30378_5182# 0.14fF
C12295 a_34090_6146# a_34090_5142# 1.00fF
C12296 a_2346_5184# a_32082_5142# 0.19fF
C12297 a_10998_14178# ctop 3.58fF
C12298 col[20] rowoff_n[10] 0.11fF
C12299 a_29982_9158# rowoff_n[7] 0.24fF
C12300 a_2346_18236# a_10906_18194# 0.35fF
C12301 a_33998_15182# rowoff_n[13] 0.24fF
C12302 a_17022_7150# m2_17220_7398# 0.16fF
C12303 m2_1732_16006# m3_1864_15134# 0.15fF
C12304 a_28978_7150# VDD 0.23fF
C12305 a_6982_7150# a_6982_6146# 1.00fF
C12306 a_23958_7150# a_24050_7150# 0.26fF
C12307 a_2346_1168# col[16] 0.14fF
C12308 a_2346_14220# col[18] 0.15fF
C12309 a_15014_14178# rowon_n[12] 0.14fF
C12310 a_2346_16228# a_14922_16186# 0.35fF
C12311 a_7986_16186# a_8990_16186# 0.97fF
C12312 a_8990_3134# col_n[6] 0.28fF
C12313 a_30074_4138# rowon_n[2] 0.14fF
C12314 a_34090_3134# ctop 3.42fF
C12315 a_4974_17190# vcm 0.60fF
C12316 rowon_n[5] row_n[5] 19.75fF
C12317 a_1962_16226# rowon_n[14] 1.18fF
C12318 col_n[16] col[17] 6.03fF
C12319 row_n[12] ctop 1.65fF
C12320 a_7986_10162# VDD 0.52fF
C12321 a_5978_17190# col[3] 0.29fF
C12322 col[4] rowoff_n[11] 0.11fF
C12323 a_15014_2130# vcm 0.62fF
C12324 a_1962_13214# a_8990_13174# 0.27fF
C12325 a_1962_10202# col[25] 0.11fF
C12326 a_6982_12170# rowoff_n[10] 0.10fF
C12327 a_7986_4138# row_n[2] 0.17fF
C12328 a_18026_1126# a_19030_1126# 0.97fF
C12329 m2_34864_8978# m3_34996_9110# 2.76fF
C12330 a_1962_4178# VDD 2.73fF
C12331 a_24050_13174# col[21] 0.29fF
C12332 m3_34996_13126# VDD 0.26fF
C12333 a_1962_17230# sample 0.14fF
C12334 a_34090_17190# rowon_n[15] 0.14fF
C12335 m2_10768_18014# col[8] 0.28fF
C12336 a_21038_14178# VDD 0.52fF
C12337 a_20034_11166# a_20034_10162# 1.00fF
C12338 a_2346_10204# a_3970_10162# 0.19fF
C12339 a_3970_2130# rowoff_n[0] 0.10fF
C12340 a_28066_6146# vcm 0.62fF
C12341 a_1962_15222# a_22042_15182# 0.27fF
C12342 m2_14784_18014# ctop 0.18fF
C12343 a_21038_16186# rowoff_n[14] 0.10fF
C12344 a_11302_15222# vcm 0.22fF
C12345 a_14010_8154# m2_14208_8402# 0.16fF
C12346 a_12002_17190# row_n[15] 0.17fF
C12347 a_2346_10204# col[9] 0.15fF
C12348 a_1962_12210# a_15318_12210# 0.14fF
C12349 a_2346_12212# a_17022_12170# 0.19fF
C12350 a_9902_12170# a_9994_12170# 0.26fF
C12351 a_27062_7150# row_n[5] 0.17fF
C12352 a_6982_6146# col[4] 0.29fF
C12353 a_35002_4138# m2_34864_3958# 0.16fF
C12354 a_2966_5142# rowoff_n[3] 0.10fF
C12355 a_1962_12210# col_n[25] 0.13fF
C12356 a_10906_2130# VDD 0.23fF
C12357 a_31078_5142# a_32082_5142# 0.97fF
C12358 a_5978_13174# ctop 3.58fF
C12359 a_24050_15182# col_n[21] 0.28fF
C12360 a_1962_6186# col[16] 0.11fF
C12361 a_35398_4178# vcm 0.23fF
C12362 a_1962_14218# a_28370_14218# 0.14fF
C12363 a_33086_15182# a_33086_14178# 1.00fF
C12364 a_2346_11208# row_n[9] 0.35fF
C12365 a_2346_14220# a_30074_14178# 0.19fF
C12366 a_25054_2130# col[22] 0.29fF
C12367 m2_26832_18014# col_n[24] 0.25fF
C12368 m2_1732_12994# m3_1864_12122# 0.15fF
C12369 a_23958_6146# VDD 0.23fF
C12370 a_15014_5142# rowon_n[3] 0.14fF
C12371 a_2346_6188# a_6890_6146# 0.35fF
C12372 a_3970_6146# a_4974_6146# 0.97fF
C12373 a_19030_17190# ctop 3.39fF
C12374 a_2346_8196# rowoff_n[6] 4.09fF
C12375 a_1962_7190# rowon_n[5] 1.18fF
C12376 a_22954_16186# a_23046_16186# 0.26fF
C12377 a_5978_16186# a_5978_15182# 1.00fF
C12378 a_8898_17190# rowoff_n[15] 0.24fF
C12379 a_29070_2130# ctop 3.39fF
C12380 m2_34864_18014# VDD 1.77fF
C12381 a_12914_6146# rowoff_n[4] 0.24fF
C12382 a_10998_9158# m2_11196_9406# 0.16fF
C12383 a_2874_9158# VDD 0.24fF
C12384 a_6982_8154# col_n[4] 0.28fF
C12385 a_2346_8196# a_19942_8154# 0.35fF
C12386 a_2346_6188# col[0] 0.15fF
C12387 a_9994_1126# vcm 0.12fF
C12388 a_22954_4138# rowoff_n[2] 0.24fF
C12389 a_1962_8194# col_n[16] 0.13fF
C12390 a_34090_8154# rowon_n[6] 0.14fF
C12391 m2_34864_5966# m3_34996_6098# 2.76fF
C12392 m2_13780_946# vcm 0.42fF
C12393 a_25054_4138# col_n[22] 0.28fF
C12394 a_1962_5182# a_14010_5142# 0.27fF
C12395 col[31] rowoff_n[10] 0.11fF
C12396 a_16018_13174# VDD 0.52fF
C12397 a_17022_10162# a_18026_10162# 0.97fF
C12398 a_2346_10204# a_32994_10162# 0.35fF
C12399 a_1962_2170# col[7] 0.11fF
C12400 a_32994_2130# rowoff_n[0] 0.24fF
C12401 a_1962_15222# col[9] 0.11fF
C12402 a_23046_5142# vcm 0.62fF
C12403 m2_30848_946# vcm 0.42fF
C12404 a_12002_8154# row_n[6] 0.17fF
C12405 m2_1732_15002# ctop 0.17fF
C12406 a_6282_14218# vcm 0.22fF
C12407 a_2966_7150# m2_1732_6970# 0.96fF
C12408 a_1962_2170# a_7286_2170# 0.14fF
C12409 a_5886_2130# a_5978_2130# 0.26fF
C12410 a_2346_2172# a_8990_2130# 0.19fF
C12411 m2_25828_18014# m3_24956_18146# 0.13fF
C12412 a_2346_1168# col[27] 0.14fF
C12413 a_2346_14220# col[29] 0.15fF
C12414 a_1962_7190# a_27062_7150# 0.27fF
C12415 a_29070_17190# VDD 0.55fF
C12416 a_2346_18236# col[1] 0.15fF
C12417 a_2346_8196# vcm 0.40fF
C12418 col_n[22] col[22] 0.72fF
C12419 rowon_n[6] ctop 1.40fF
C12420 a_19334_18234# vcm 0.22fF
C12421 a_5886_1126# VDD 0.44fF
C12422 col[15] rowoff_n[11] 0.11fF
C12423 a_7986_10162# m2_8184_10410# 0.16fF
C12424 a_1962_4178# a_20338_4178# 0.14fF
C12425 a_2346_4180# a_22042_4138# 0.19fF
C12426 a_29070_5142# a_29070_4138# 1.00fF
C12427 a_4974_11166# col[2] 0.29fF
C12428 a_2346_2172# row_n[0] 0.35fF
C12429 a_29374_3174# vcm 0.22fF
C12430 a_31078_11166# row_n[9] 0.17fF
C12431 a_30074_14178# a_31078_14178# 0.97fF
C12432 a_21038_10162# rowoff_n[8] 0.10fF
C12433 a_23046_13174# rowoff_n[11] 0.10fF
C12434 a_1962_4178# col_n[7] 0.13fF
C12435 a_1962_17230# col_n[9] 0.13fF
C12436 m2_1732_9982# m3_1864_9110# 0.15fF
C12437 a_23046_7150# col[20] 0.29fF
C12438 a_18938_5142# VDD 0.23fF
C12439 a_18938_6146# a_19030_6146# 0.26fF
C12440 a_1962_6186# a_33390_6186# 0.14fF
C12441 a_14010_16186# ctop 3.57fF
C12442 a_2966_14178# VDD 0.56fF
C12443 a_31078_8154# rowoff_n[6] 0.10fF
C12444 a_1962_11206# col[0] 0.11fF
C12445 a_2346_15224# a_4882_15182# 0.35fF
C12446 a_2966_16186# rowoff_n[14] 0.10fF
C12447 m2_12776_946# m2_13204_1374# 0.16fF
C12448 a_2346_10204# col[20] 0.15fF
C12449 a_31990_9158# VDD 0.23fF
C12450 a_19030_9158# rowon_n[7] 0.14fF
C12451 a_1962_18234# a_22346_18234# 0.14fF
C12452 m2_34864_16006# rowon_n[14] 0.13fF
C12453 a_4974_13174# col_n[2] 0.28fF
C12454 a_2346_17232# a_17934_17190# 0.35fF
C12455 m2_24824_18014# m2_25828_18014# 0.96fF
C12456 m2_34864_2954# m3_34996_3086# 2.76fF
C12457 m3_1864_11118# ctop 0.23fF
C12458 a_4974_11166# m2_5172_11414# 0.16fF
C12459 a_1962_6186# col[27] 0.11fF
C12460 a_10998_12170# VDD 0.52fF
C12461 m2_29844_946# m2_30272_1374# 0.16fF
C12462 a_15014_10162# a_15014_9158# 1.00fF
C12463 a_31990_10162# a_32082_10162# 0.26fF
C12464 a_23046_9158# col_n[20] 0.28fF
C12465 a_18026_4138# vcm 0.62fF
C12466 a_1962_14218# a_12002_14178# 0.27fF
C12467 a_10906_14178# rowoff_n[12] 0.24fF
C12468 a_1962_13214# vcm 6.95fF
C12469 a_24050_16186# VDD 0.52fF
C12470 a_1962_11206# a_5278_11206# 0.14fF
C12471 a_2346_11208# a_6982_11166# 0.19fF
C12472 a_4882_11166# a_4974_11166# 0.26fF
C12473 a_31078_8154# vcm 0.62fF
C12474 a_1962_16226# a_25054_16186# 0.27fF
C12475 a_12002_2130# m2_12200_2378# 0.16fF
C12476 a_16018_12170# row_n[10] 0.17fF
C12477 a_14314_17230# vcm 0.22fF
C12478 a_26058_4138# a_27062_4138# 0.97fF
C12479 a_2346_6188# col[11] 0.15fF
C12480 a_5978_2130# col_n[3] 0.28fF
C12481 a_31078_2130# row_n[0] 0.17fF
C12482 a_24354_2170# vcm 0.22fF
C12483 a_1962_13214# a_18330_13214# 0.14fF
C12484 a_2346_13216# a_20034_13174# 0.19fF
C12485 a_28066_14178# a_28066_13174# 1.00fF
C12486 a_1962_8194# col_n[27] 0.13fF
C12487 m2_34864_3958# m2_34864_2954# 0.99fF
C12488 m2_13780_946# col_n[11] 0.37fF
C12489 m2_1732_6970# m3_1864_6098# 0.15fF
C12490 a_13918_4138# VDD 0.23fF
C12491 a_1962_2170# col[18] 0.11fF
C12492 m3_20940_1078# VDD 0.14fF
C12493 a_1962_15222# col[20] 0.11fF
C12494 a_8990_15182# ctop 3.58fF
C12495 m2_22816_946# m2_23244_1374# 0.16fF
C12496 a_21038_12170# col[18] 0.29fF
C12497 a_3970_10162# rowon_n[8] 0.14fF
C12498 a_2346_15224# a_33086_15182# 0.19fF
C12499 a_1962_15222# a_31382_15222# 0.14fF
C12500 a_17934_15182# a_18026_15182# 0.26fF
C12501 m2_1732_18014# m3_1864_18146# 2.79fF
C12502 a_26970_8154# VDD 0.23fF
C12503 a_3970_7150# rowoff_n[5] 0.10fF
C12504 a_2346_18236# col[12] 0.14fF
C12505 a_2346_7192# a_9902_7150# 0.35fF
C12506 row_n[1] ctop 1.64fF
C12507 col_n[27] col[28] 5.90fF
C12508 m2_21812_946# m3_22948_1078# 0.13fF
C12509 col[26] rowoff_n[11] 0.11fF
C12510 a_1962_3174# m2_34864_2954# 0.17fF
C12511 a_14010_5142# rowoff_n[3] 0.10fF
C12512 a_32082_4138# ctop 3.58fF
C12513 a_2346_2172# col[2] 0.15fF
C12514 a_2346_15224# col[4] 0.15fF
C12515 a_1962_4178# a_3970_4138# 0.27fF
C12516 a_23046_13174# rowon_n[11] 0.14fF
C12517 a_3970_5142# col[1] 0.29fF
C12518 a_5978_11166# VDD 0.52fF
C12519 m2_32856_946# m3_31984_1078# 0.13fF
C12520 a_12002_9158# a_13006_9158# 0.97fF
C12521 a_2346_9200# a_22954_9158# 0.35fF
C12522 a_1962_4178# col_n[18] 0.13fF
C12523 a_13006_3134# vcm 0.62fF
C12524 a_24050_3134# rowoff_n[1] 0.10fF
C12525 a_1962_17230# col_n[20] 0.13fF
C12526 a_2966_10162# rowoff_n[8] 0.10fF
C12527 a_21038_14178# col_n[18] 0.28fF
C12528 a_1962_18234# ctop 0.30fF
C12529 a_1962_11206# col[11] 0.11fF
C12530 a_1962_6186# a_17022_6146# 0.27fF
C12531 a_33086_14178# m2_33284_14426# 0.16fF
C12532 a_19030_15182# VDD 0.52fF
C12533 m2_34864_7974# vcm 0.50fF
C12534 a_16018_3134# row_n[1] 0.17fF
C12535 col[10] rowoff_n[12] 0.11fF
C12536 a_26058_7150# vcm 0.62fF
C12537 a_2346_10204# col[31] 0.15fF
C12538 a_9294_16226# vcm 0.22fF
C12539 a_2346_3176# a_12002_3134# 0.19fF
C12540 a_1962_3174# a_10298_3174# 0.14fF
C12541 a_24050_4138# a_24050_3134# 1.00fF
C12542 a_27062_2130# m2_26832_946# 0.99fF
C12543 a_4974_2130# m3_4876_1078# 0.15fF
C12544 a_1962_8194# a_30074_8154# 0.27fF
C12545 a_19334_1166# vcm 0.22fF
C12546 a_25054_13174# a_26058_13174# 0.97fF
C12547 a_3970_7150# col_n[1] 0.28fF
C12548 a_12914_11166# rowoff_n[9] 0.24fF
C12549 a_20034_16186# row_n[14] 0.17fF
C12550 m2_1732_3958# m3_1864_3086# 0.15fF
C12551 a_8898_3134# VDD 0.23fF
C12552 a_13918_5142# a_14010_5142# 0.26fF
C12553 a_1962_5182# a_23350_5182# 0.14fF
C12554 a_2346_5184# a_25054_5142# 0.19fF
C12555 a_3970_14178# ctop 3.57fF
C12556 a_22042_3134# col_n[19] 0.28fF
C12557 a_22954_9158# rowoff_n[7] 0.24fF
C12558 ctop rowoff_n[13] 0.60fF
C12559 a_1962_13214# col_n[11] 0.13fF
C12560 a_32386_5182# vcm 0.22fF
C12561 a_19030_17190# col[16] 0.29fF
C12562 a_26970_15182# rowoff_n[13] 0.24fF
C12563 a_21950_7150# VDD 0.23fF
C12564 a_1962_7190# col[2] 0.11fF
C12565 a_32994_7150# rowoff_n[5] 0.24fF
C12566 a_30074_15182# m2_30272_15430# 0.16fF
C12567 a_7986_14178# rowon_n[12] 0.14fF
C12568 a_2346_16228# a_7894_16186# 0.35fF
C12569 a_2346_6188# col[22] 0.15fF
C12570 m2_1732_9982# sample_n 0.15fF
C12571 a_32082_3134# m2_32280_3382# 0.16fF
C12572 a_23046_4138# rowon_n[2] 0.14fF
C12573 a_27062_3134# ctop 3.57fF
C12574 a_35002_11166# VDD 0.29fF
C12575 a_26970_9158# a_27062_9158# 0.26fF
C12576 a_9994_9158# a_9994_8154# 1.00fF
C12577 a_7986_2130# vcm 0.62fF
C12578 a_1962_2170# col[29] 0.11fF
C12579 a_2346_1168# a_27974_1126# 0.35fF
C12580 a_2966_5142# m2_3164_5390# 0.16fF
C12581 a_1962_15222# col[31] 0.11fF
C12582 m3_16924_18146# VDD 0.24fF
C12583 a_27062_17190# rowon_n[15] 0.14fF
C12584 a_14010_14178# VDD 0.52fF
C12585 a_20034_6146# col[17] 0.29fF
C12586 m2_18224_1374# a_18026_1126# 0.16fF
C12587 a_1962_9198# col_n[2] 0.13fF
C12588 a_21038_6146# vcm 0.62fF
C12589 a_1962_15222# a_15014_15182# 0.27fF
C12590 a_4274_15222# vcm 0.22fF
C12591 a_14010_16186# rowoff_n[14] 0.10fF
C12592 a_2346_18236# col[23] 0.14fF
C12593 a_21038_3134# a_22042_3134# 0.97fF
C12594 a_4974_17190# row_n[15] 0.17fF
C12595 a_23958_1126# m2_23820_946# 0.16fF
C12596 ctop col[0] 1.56fF
C12597 a_27062_16186# m2_27260_16434# 0.16fF
C12598 m2_29844_18014# vcm 0.28fF
C12599 a_1962_12210# a_8290_12210# 0.14fF
C12600 a_23046_13174# a_23046_12170# 1.00fF
C12601 a_2346_12212# a_9994_12170# 0.19fF
C12602 a_20034_7150# row_n[5] 0.17fF
C12603 a_2346_2172# col[13] 0.15fF
C12604 a_34090_10162# vcm 0.62fF
C12605 a_1962_17230# a_28066_17190# 0.27fF
C12606 a_2346_15224# col[15] 0.15fF
C12607 m2_1732_17010# m2_2160_17438# 0.16fF
C12608 a_29070_4138# m2_29268_4386# 0.16fF
C12609 m2_1732_946# m3_1864_1078# 2.79fF
C12610 m2_2736_946# m3_2868_2082# 0.15fF
C12611 m3_23952_1078# ctop 0.23fF
C12612 a_1962_4178# col_n[29] 0.13fF
C12613 a_2966_9158# a_3970_9158# 0.97fF
C12614 a_1962_17230# col_n[31] 0.13fF
C12615 a_27366_4178# vcm 0.22fF
C12616 a_1962_14218# a_21342_14218# 0.14fF
C12617 a_12914_14178# a_13006_14178# 0.26fF
C12618 a_2346_14220# a_23046_14178# 0.19fF
C12619 a_20034_8154# col_n[17] 0.28fF
C12620 a_1962_18234# col[5] 0.11fF
C12621 a_1962_11206# col[22] 0.11fF
C12622 m2_23820_946# col[21] 0.39fF
C12623 a_34090_7150# m2_34864_6970# 0.96fF
C12624 a_16930_6146# VDD 0.23fF
C12625 a_7986_5142# rowon_n[3] 0.14fF
C12626 a_12002_17190# ctop 3.39fF
C12627 col[21] rowoff_n[12] 0.11fF
C12628 a_2346_16228# a_2346_15224# 0.22fF
C12629 a_1962_16226# a_35398_16226# 0.14fF
C12630 m2_34864_4962# row_n[3] 0.15fF
C12631 a_22042_2130# ctop 3.39fF
C12632 m2_20808_18014# VDD 0.91fF
C12633 a_5886_6146# rowoff_n[4] 0.24fF
C12634 a_29982_10162# VDD 0.23fF
C12635 a_6982_8154# a_7986_8154# 0.97fF
C12636 a_24050_17190# m2_24248_17438# 0.16fF
C12637 a_2346_8196# a_12914_8154# 0.35fF
C12638 a_28978_12170# rowoff_n[10] 0.24fF
C12639 a_15926_4138# rowoff_n[2] 0.24fF
C12640 a_2346_11208# col[6] 0.15fF
C12641 a_26058_5142# m2_26256_5390# 0.16fF
C12642 a_27062_8154# rowon_n[6] 0.14fF
C12643 a_1962_5182# a_6982_5142# 0.27fF
C12644 col[5] rowoff_n[13] 0.11fF
C12645 a_8990_13174# VDD 0.52fF
C12646 a_2346_18236# m2_30848_18014# 0.19fF
C12647 a_1962_13214# col_n[22] 0.13fF
C12648 m2_6752_946# vcm 0.42fF
C12649 a_2346_10204# a_25966_10162# 0.35fF
C12650 a_25966_2130# rowoff_n[0] 0.24fF
C12651 a_16018_5142# vcm 0.62fF
C12652 a_18026_11166# col[15] 0.29fF
C12653 a_4974_8154# row_n[6] 0.17fF
C12654 a_1962_7190# col[13] 0.11fF
C12655 a_2346_12212# rowon_n[10] 0.26fF
C12656 a_19030_3134# a_19030_2130# 1.00fF
C12657 m2_15788_18014# m3_16924_18146# 0.13fF
C12658 a_3878_7150# VDD 0.23fF
C12659 a_1962_7190# a_20034_7150# 0.27fF
C12660 a_2966_4138# col[0] 0.29fF
C12661 a_22042_17190# VDD 0.55fF
C12662 a_20034_12170# a_21038_12170# 0.97fF
C12663 m2_1732_946# sample 0.16fF
C12664 a_29070_9158# vcm 0.62fF
C12665 a_12306_18234# vcm 0.22fF
C12666 a_32082_2130# VDD 0.55fF
C12667 a_1962_10202# m2_1732_9982# 0.15fF
C12668 a_2346_4180# a_15014_4138# 0.19fF
C12669 a_1962_4178# a_13310_4178# 0.14fF
C12670 a_8898_4138# a_8990_4138# 0.26fF
C12671 a_1962_9198# a_33086_9158# 0.27fF
C12672 a_22346_3174# vcm 0.22fF
C12673 a_24050_11166# row_n[9] 0.17fF
C12674 a_14010_10162# rowoff_n[8] 0.10fF
C12675 a_16018_13174# rowoff_n[11] 0.10fF
C12676 a_23046_6146# m2_23244_6394# 0.16fF
C12677 a_11910_5142# VDD 0.23fF
C12678 a_18026_13174# col_n[15] 0.28fF
C12679 a_1962_6186# a_26362_6186# 0.14fF
C12680 a_32082_7150# a_32082_6146# 1.00fF
C12681 a_2346_6188# a_28066_6146# 0.19fF
C12682 a_1962_9198# col_n[13] 0.13fF
C12683 a_6982_16186# ctop 3.57fF
C12684 a_24050_8154# rowoff_n[6] 0.10fF
C12685 m2_12776_946# a_1962_1166# 0.18fF
C12686 a_19030_17190# m3_18932_18146# 0.15fF
C12687 a_2966_6146# vcm 0.61fF
C12688 a_33086_16186# a_34090_16186# 0.97fF
C12689 a_1962_3174# col[4] 0.11fF
C12690 a_1962_16226# col[6] 0.11fF
C12691 ctop col[11] 1.98fF
C12692 col[2] col[3] 0.20fF
C12693 a_30074_17190# rowoff_n[15] 0.10fF
C12694 a_34090_6146# rowoff_n[4] 0.10fF
C12695 a_1962_1166# m2_29844_946# 0.18fF
C12696 a_24962_9158# VDD 0.23fF
C12697 a_12002_9158# rowon_n[7] 0.14fF
C12698 a_4974_8154# a_4974_7150# 1.00fF
C12699 a_21950_8154# a_22042_8154# 0.26fF
C12700 a_2346_2172# col[24] 0.15fF
C12701 a_1962_18234# a_15318_18234# 0.14fF
C12702 a_2346_15224# col[26] 0.15fF
C12703 a_2346_17232# a_10906_17190# 0.35fF
C12704 a_5978_17190# a_6982_17190# 0.97fF
C12705 m2_17796_18014# m2_18800_18014# 0.96fF
C12706 a_30074_5142# ctop 3.58fF
C12707 m3_19936_18146# ctop 0.23fF
C12708 a_1962_5182# a_34394_5182# 0.14fF
C12709 a_3970_12170# VDD 0.52fF
C12710 a_1962_18234# col[16] 0.11fF
C12711 a_10998_4138# vcm 0.62fF
C12712 a_1962_14218# a_4974_14178# 0.27fF
C12713 a_3878_14178# a_3970_14178# 0.26fF
C12714 a_2346_3176# rowon_n[1] 0.26fF
C12715 a_19030_2130# col_n[16] 0.26fF
C12716 a_31078_12170# rowon_n[10] 0.14fF
C12717 a_16018_2130# a_17022_2130# 0.97fF
C12718 a_20034_7150# m2_20232_7398# 0.16fF
C12719 a_2346_2172# a_30986_2130# 0.35fF
C12720 a_16018_16186# col[13] 0.29fF
C12721 a_1962_5182# col_n[4] 0.13fF
C12722 a_17022_16186# VDD 0.52fF
C12723 m2_1732_10986# vcm 0.45fF
C12724 a_18026_12170# a_18026_11166# 1.00fF
C12725 a_24050_8154# vcm 0.62fF
C12726 a_1962_16226# a_18026_16186# 0.27fF
C12727 a_8990_12170# row_n[10] 0.17fF
C12728 a_34090_12170# col[31] 0.29fF
C12729 a_7286_17230# vcm 0.22fF
C12730 a_24050_2130# row_n[0] 0.17fF
C12731 a_20034_17190# m2_19804_18014# 1.00fF
C12732 a_2346_11208# col[17] 0.15fF
C12733 a_17326_2170# vcm 0.22fF
C12734 a_1962_13214# a_11302_13214# 0.14fF
C12735 a_2346_13216# a_13006_13174# 0.19fF
C12736 a_7894_13174# a_7986_13174# 0.26fF
C12737 col[16] rowoff_n[13] 0.11fF
C12738 a_6890_4138# VDD 0.23fF
C12739 m3_1864_5094# VDD 0.25fF
C12740 a_29070_6146# a_30074_6146# 0.97fF
C12741 VDD rowoff_n[6] 1.17fF
C12742 sample_n rowoff_n[7] 0.38fF
C12743 a_28066_15182# row_n[13] 0.17fF
C12744 a_1962_7190# col[24] 0.11fF
C12745 a_30378_6186# vcm 0.22fF
C12746 a_1962_15222# a_24354_15222# 0.14fF
C12747 a_2346_15224# a_26058_15182# 0.19fF
C12748 a_31078_16186# a_31078_15182# 1.00fF
C12749 a_17022_5142# col[14] 0.29fF
C12750 a_17022_8154# m2_17220_8402# 0.16fF
C12751 a_19942_8154# VDD 0.23fF
C12752 a_34090_14178# col_n[31] 0.28fF
C12753 m2_11772_946# m3_11904_1078# 2.79fF
C12754 a_20946_17190# a_21038_17190# 0.26fF
C12755 a_3970_17190# a_3970_16186# 1.00fF
C12756 col[0] rowoff_n[14] 0.11fF
C12757 a_6982_5142# rowoff_n[3] 0.10fF
C12758 a_25054_4138# ctop 3.58fF
C12759 a_16018_13174# rowon_n[11] 0.14fF
C12760 a_32994_12170# VDD 0.23fF
C12761 m3_32988_18146# m3_33992_18146# 0.22fF
C12762 m2_34864_946# m3_34996_2082# 0.15fF
C12763 a_2346_9200# a_15926_9158# 0.35fF
C12764 a_2346_7192# col[8] 0.15fF
C12765 a_5978_3134# vcm 0.62fF
C12766 a_31078_3134# rowon_n[1] 0.14fF
C12767 a_17022_3134# rowoff_n[1] 0.10fF
C12768 a_32082_14178# rowoff_n[12] 0.10fF
C12769 a_1962_9198# col_n[24] 0.13fF
C12770 a_30986_2130# a_31078_2130# 0.26fF
C12771 a_17022_7150# col_n[14] 0.28fF
C12772 a_1962_6186# a_9994_6146# 0.27fF
C12773 a_12002_15182# VDD 0.52fF
C12774 a_15014_11166# a_16018_11166# 0.97fF
C12775 a_2346_11208# a_28978_11166# 0.35fF
C12776 a_8990_3134# row_n[1] 0.17fF
C12777 a_1962_3174# col[15] 0.11fF
C12778 VDD vcm 73.66fF
C12779 a_1962_16226# col[17] 0.11fF
C12780 m2_2736_18014# col_n[0] 0.25fF
C12781 ctop col[22] 1.98fF
C12782 a_19030_7150# vcm 0.62fF
C12783 m2_4744_18014# col[2] 0.28fF
C12784 a_2346_3176# a_4974_3134# 0.19fF
C12785 a_14010_9158# m2_14208_9406# 0.16fF
C12786 a_1962_3174# a_3270_3174# 0.14fF
C12787 a_32082_17190# col[29] 0.29fF
C12788 a_1962_8194# a_23046_8154# 0.27fF
C12789 a_12306_1166# vcm 0.23fF
C12790 a_32082_11166# vcm 0.62fF
C12791 a_5886_11166# rowoff_n[9] 0.24fF
C12792 a_13006_16186# row_n[14] 0.17fF
C12793 a_35002_5142# m2_34864_4962# 0.16fF
C12794 a_27062_6146# a_27062_5142# 1.00fF
C12795 a_2346_5184# a_18026_5142# 0.19fF
C12796 a_1962_5182# a_16322_5182# 0.14fF
C12797 a_1962_18234# col[27] 0.11fF
C12798 a_28066_6146# row_n[4] 0.17fF
C12799 a_15926_9158# rowoff_n[7] 0.24fF
C12800 a_2346_16228# col[1] 0.15fF
C12801 a_25358_5182# vcm 0.22fF
C12802 a_28066_15182# a_29070_15182# 0.97fF
C12803 a_19942_15182# rowoff_n[13] 0.24fF
C12804 a_1962_5182# col_n[15] 0.13fF
C12805 a_15014_10162# col[12] 0.29fF
C12806 m2_30848_18014# m3_29976_18146# 0.13fF
C12807 a_14922_7150# VDD 0.23fF
C12808 a_25966_7150# rowoff_n[5] 0.24fF
C12809 a_2346_7192# a_31078_7150# 0.19fF
C12810 a_1962_7190# a_29374_7190# 0.14fF
C12811 a_16930_7150# a_17022_7150# 0.26fF
C12812 m2_20808_18014# col_n[18] 0.25fF
C12813 a_1962_12210# col[8] 0.11fF
C12814 a_33086_6146# col[30] 0.29fF
C12815 a_16018_4138# rowon_n[2] 0.14fF
C12816 a_20034_3134# ctop 3.57fF
C12817 a_10998_10162# m2_11196_10410# 0.16fF
C12818 a_27974_11166# VDD 0.23fF
C12819 a_2346_11208# col[28] 0.15fF
C12820 a_3970_18194# vcm 0.12fF
C12821 m3_22948_1078# m3_23952_1078# 0.22fF
C12822 col[27] rowoff_n[13] 0.11fF
C12823 a_2346_1168# a_20946_1126# 0.35fF
C12824 a_33086_7150# ctop 3.57fF
C12825 a_20034_17190# rowon_n[15] 0.14fF
C12826 a_6982_14178# VDD 0.52fF
C12827 m2_34864_6970# rowon_n[5] 0.13fF
C12828 a_13006_11166# a_13006_10162# 1.00fF
C12829 a_15014_12170# col_n[12] 0.28fF
C12830 a_29982_11166# a_30074_11166# 0.26fF
C12831 m2_10768_946# col_n[8] 0.37fF
C12832 a_14010_6146# vcm 0.62fF
C12833 a_1962_15222# a_7986_15182# 0.27fF
C12834 a_1962_1166# col_n[6] 0.13fF
C12835 a_6982_16186# rowoff_n[14] 0.10fF
C12836 a_1962_14218# col_n[8] 0.13fF
C12837 a_2966_8154# m2_1732_7974# 0.96fF
C12838 a_2346_3176# a_33998_3134# 0.35fF
C12839 a_35494_9520# VDD 0.11fF
C12840 a_33086_8154# col_n[30] 0.28fF
C12841 col[11] rowoff_n[14] 0.11fF
C12842 m2_15788_18014# vcm 0.28fF
C12843 a_2346_12212# a_2874_12170# 0.35fF
C12844 a_13006_7150# row_n[5] 0.17fF
C12845 a_27062_10162# vcm 0.62fF
C12846 a_34090_11166# rowoff_n[9] 0.10fF
C12847 a_1962_17230# a_21038_17190# 0.27fF
C12848 m2_28840_18014# m2_29268_18442# 0.16fF
C12849 a_30074_3134# VDD 0.52fF
C12850 m3_34996_4090# ctop 0.23fF
C12851 a_7986_11166# m2_8184_11414# 0.16fF
C12852 a_24050_5142# a_25054_5142# 0.97fF
C12853 a_2346_7192# col[19] 0.15fF
C12854 a_20338_4178# vcm 0.22fF
C12855 a_26058_15182# a_26058_14178# 1.00fF
C12856 a_1962_14218# a_14314_14218# 0.14fF
C12857 a_2346_14220# a_16018_14178# 0.19fF
C12858 m2_1732_6970# m2_1732_5966# 0.99fF
C12859 a_9902_6146# VDD 0.23fF
C12860 a_1962_3174# col[26] 0.11fF
C12861 VDD col_n[11] 4.95fF
C12862 a_4974_17190# ctop 3.39fF
C12863 a_32082_10162# row_n[8] 0.17fF
C12864 vcm col_n[7] 2.80fF
C12865 col_n[3] col_n[4] 0.10fF
C12866 col[13] col[14] 0.20fF
C12867 a_1962_16226# col[28] 0.11fF
C12868 a_13006_15182# col[10] 0.29fF
C12869 a_33390_8194# vcm 0.22fF
C12870 a_2346_16228# a_29070_16186# 0.19fF
C12871 a_15926_16186# a_16018_16186# 0.26fF
C12872 a_1962_16226# a_27366_16226# 0.14fF
C12873 m2_1732_8978# row_n[7] 0.13fF
C12874 a_15014_2130# m2_15212_2378# 0.16fF
C12875 a_1962_10202# col_n[0] 0.13fF
C12876 a_15014_2130# ctop 3.39fF
C12877 m2_6752_18014# VDD 1.26fF
C12878 a_1962_18234# m2_21812_18014# 0.18fF
C12879 a_22954_10162# VDD 0.23fF
C12880 a_31078_11166# col[28] 0.29fF
C12881 a_2346_8196# a_5886_8154# 0.35fF
C12882 a_21950_12170# rowoff_n[10] 0.24fF
C12883 a_8898_4138# rowoff_n[2] 0.24fF
C12884 a_20034_8154# rowon_n[6] 0.14fF
C12885 a_28066_6146# ctop 3.58fF
C12886 a_2346_3176# col[10] 0.15fF
C12887 a_4974_12170# m2_5172_12418# 0.16fF
C12888 m3_34996_1078# VDD 0.23fF
C12889 a_2346_16228# col[12] 0.15fF
C12890 a_2346_18236# m2_16792_18014# 0.19fF
C12891 a_2346_10204# a_18938_10162# 0.35fF
C12892 a_9994_10162# a_10998_10162# 0.97fF
C12893 a_18938_2130# rowoff_n[0] 0.24fF
C12894 a_1962_5182# col_n[26] 0.13fF
C12895 a_8990_5142# vcm 0.62fF
C12896 a_13006_17190# col_n[10] 0.28fF
C12897 a_14010_4138# col[11] 0.29fF
C12898 m2_6752_18014# m3_6884_18146# 2.78fF
C12899 a_1962_7190# a_13006_7150# 0.27fF
C12900 a_1962_12210# col[19] 0.11fF
C12901 a_15014_17190# VDD 0.55fF
C12902 a_2346_12212# a_31990_12170# 0.35fF
C12903 a_31078_13174# col_n[28] 0.28fF
C12904 a_22042_9158# vcm 0.62fF
C12905 a_5278_18234# vcm 0.22fF
C12906 a_25054_2130# VDD 0.55fF
C12907 a_22042_5142# a_22042_4138# 1.00fF
C12908 a_1962_4178# a_6282_4178# 0.14fF
C12909 a_2346_4180# a_7986_4138# 0.19fF
C12910 m3_1864_8106# m3_1864_7102# 0.22fF
C12911 a_18938_18194# m2_18800_18014# 0.16fF
C12912 a_1962_9198# a_26058_9158# 0.27fF
C12913 a_17022_11166# row_n[9] 0.17fF
C12914 a_15318_3174# vcm 0.22fF
C12915 a_23046_14178# a_24050_14178# 0.97fF
C12916 a_6982_10162# rowoff_n[8] 0.10fF
C12917 a_35094_13174# vcm 0.12fF
C12918 a_8990_13174# rowoff_n[11] 0.10fF
C12919 m2_1732_1950# VDD 1.04fF
C12920 m2_22816_946# col_n[20] 0.37fF
C12921 a_2346_1168# a_1962_1166# 2.55fF
C12922 a_4882_5142# VDD 0.23fF
C12923 a_2346_12212# col[3] 0.15fF
C12924 a_11910_6146# a_12002_6146# 0.26fF
C12925 a_1962_6186# a_19334_6186# 0.14fF
C12926 a_2346_6188# a_21038_6146# 0.19fF
C12927 a_17022_8154# rowoff_n[6] 0.10fF
C12928 a_14010_6146# col_n[11] 0.28fF
C12929 a_1962_1166# col_n[17] 0.12fF
C12930 a_28370_7190# vcm 0.22fF
C12931 a_1962_14218# col_n[19] 0.13fF
C12932 a_1962_1166# m2_5748_946# 0.18fF
C12933 a_3970_1126# m2_2736_946# 0.96fF
C12934 a_23046_17190# rowoff_n[15] 0.10fF
C12935 a_27062_6146# rowoff_n[4] 0.10fF
C12936 a_7986_2130# m3_7888_1078# 0.15fF
C12937 a_17934_9158# VDD 0.23fF
C12938 a_4974_9158# rowon_n[7] 0.14fF
C12939 a_32082_2130# col_n[29] 0.29fF
C12940 col[22] rowoff_n[14] 0.11fF
C12941 a_1962_8194# col[10] 0.11fF
C12942 a_2346_8196# a_34090_8154# 0.19fF
C12943 a_1962_8194# a_32386_8194# 0.14fF
C12944 m2_13780_946# ctop 0.18fF
C12945 a_1962_18234# a_8290_18234# 0.14fF
C12946 a_29070_16186# col[26] 0.29fF
C12947 m2_5748_946# m2_6176_1374# 0.16fF
C12948 a_1962_17230# a_2966_17190# 0.27fF
C12949 a_2346_7192# col[30] 0.15fF
C12950 a_1962_4178# m2_34864_3958# 0.17fF
C12951 m2_10768_18014# m2_11772_18014# 0.96fF
C12952 a_23046_5142# ctop 3.58fF
C12953 m2_30848_946# ctop 0.18fF
C12954 a_30986_13174# VDD 0.23fF
C12955 a_24962_10162# a_25054_10162# 0.26fF
C12956 a_7986_10162# a_7986_9158# 1.00fF
C12957 a_3970_4138# vcm 0.62fF
C12958 a_24050_12170# rowon_n[10] 0.14fF
C12959 a_2346_2172# a_23958_2130# 0.35fF
C12960 VDD col_n[22] 4.94fF
C12961 vcm col_n[18] 2.80fF
C12962 a_2346_8196# ctop 1.59fF
C12963 col[6] rowoff_n[15] 0.11fF
C12964 a_33086_15182# m2_33284_15430# 0.16fF
C12965 a_9994_16186# VDD 0.52fF
C12966 a_12002_9158# col[9] 0.29fF
C12967 a_1962_10202# col_n[10] 0.13fF
C12968 a_17022_8154# vcm 0.62fF
C12969 a_1962_16226# a_10998_16186# 0.27fF
C12970 a_20034_1126# VDD 0.58fF
C12971 a_19030_4138# a_20034_4138# 0.97fF
C12972 a_1962_4178# a_1962_3174# 0.16fF
C12973 a_1962_4178# col[1] 0.11fF
C12974 a_30074_5142# col[27] 0.29fF
C12975 a_1962_17230# col[3] 0.11fF
C12976 a_17022_2130# row_n[0] 0.17fF
C12977 a_10298_2170# vcm 0.22fF
C12978 a_1962_13214# a_4274_13214# 0.14fF
C12979 a_2346_13216# a_5978_13174# 0.19fF
C12980 a_21038_14178# a_21038_13174# 1.00fF
C12981 a_30074_12170# vcm 0.62fF
C12982 a_3878_12170# rowoff_n[10] 0.24fF
C12983 a_2346_3176# col[21] 0.15fF
C12984 a_2346_16228# col[23] 0.15fF
C12985 a_33086_5142# VDD 0.52fF
C12986 m3_31984_18146# VDD 0.29fF
C12987 a_21038_15182# row_n[13] 0.17fF
C12988 a_23350_6186# vcm 0.22fF
C12989 a_10906_15182# a_10998_15182# 0.26fF
C12990 a_2346_15224# a_19030_15182# 0.19fF
C12991 a_1962_15222# a_17326_15222# 0.14fF
C12992 a_12002_11166# col_n[9] 0.28fF
C12993 a_1962_12210# col[30] 0.11fF
C12994 a_3970_1126# m3_3872_1078# 2.44fF
C12995 a_12914_8154# VDD 0.23fF
C12996 a_32082_8154# a_33086_8154# 0.97fF
C12997 a_30074_16186# m2_30272_16434# 0.16fF
C12998 a_1962_6186# col_n[1] 0.13fF
C12999 a_30074_7150# col_n[27] 0.28fF
C13000 a_2346_17232# a_32082_17190# 0.19fF
C13001 a_1962_17230# a_30378_17230# 0.14fF
C13002 a_32082_4138# m2_32280_4386# 0.16fF
C13003 a_18026_4138# ctop 3.58fF
C13004 m2_6752_946# m3_7888_1078# 0.13fF
C13005 a_1962_13214# ctop 1.49fF
C13006 a_8990_13174# rowon_n[11] 0.14fF
C13007 a_25966_12170# VDD 0.23fF
C13008 m3_18932_18146# m3_19936_18146# 0.22fF
C13009 a_4974_9158# a_5978_9158# 0.97fF
C13010 a_2346_9200# a_8898_9158# 0.35fF
C13011 a_9994_3134# rowoff_n[1] 0.10fF
C13012 a_24050_3134# rowon_n[1] 0.14fF
C13013 a_25054_14178# rowoff_n[12] 0.10fF
C13014 a_2346_12212# col[14] 0.15fF
C13015 a_2966_6146# m2_3164_6394# 0.16fF
C13016 a_31078_8154# ctop 3.58fF
C13017 a_2346_6188# a_2966_6146# 0.21fF
C13018 a_1962_1166# col_n[28] 0.13fF
C13019 a_4974_15182# VDD 0.52fF
C13020 a_1962_14218# col_n[30] 0.13fF
C13021 a_2346_11208# a_21950_11166# 0.35fF
C13022 m2_11772_946# a_12002_2130# 0.99fF
C13023 a_12002_7150# vcm 0.62fF
C13024 a_9994_14178# col[7] 0.29fF
C13025 a_28066_16186# rowon_n[14] 0.14fF
C13026 a_1962_8194# col[21] 0.11fF
C13027 a_17022_4138# a_17022_3134# 1.00fF
C13028 a_33998_4138# a_34090_4138# 0.26fF
C13029 a_1962_8194# a_16018_8154# 0.27fF
C13030 a_27062_17190# m2_27260_17438# 0.16fF
C13031 a_28066_10162# col[25] 0.29fF
C13032 a_5278_1166# vcm 0.23fF
C13033 a_2346_13216# a_35002_13174# 0.35fF
C13034 a_18026_13174# a_19030_13174# 0.97fF
C13035 a_25054_11166# vcm 0.62fF
C13036 a_5978_16186# row_n[14] 0.17fF
C13037 a_29070_5142# m2_29268_5390# 0.16fF
C13038 a_28066_4138# VDD 0.52fF
C13039 a_1962_5182# a_9294_5182# 0.14fF
C13040 a_2346_5184# a_10998_5142# 0.19fF
C13041 a_6890_5142# a_6982_5142# 0.26fF
C13042 a_21038_6146# row_n[4] 0.17fF
C13043 a_1962_10202# a_29070_10162# 0.27fF
C13044 a_8898_9158# rowoff_n[7] 0.24fF
C13045 a_18330_5182# vcm 0.22fF
C13046 vcm col_n[29] 2.80fF
C13047 VDD row_n[15] 3.05fF
C13048 col[24] col[25] 0.20fF
C13049 col[17] rowoff_n[15] 0.11fF
C13050 a_2346_8196# col[5] 0.15fF
C13051 a_12914_15182# rowoff_n[13] 0.24fF
C13052 a_34090_8154# m2_34864_7974# 0.96fF
C13053 m2_20808_18014# m3_21944_18146# 0.13fF
C13054 vcm rowoff_n[11] 0.20fF
C13055 a_9994_16186# col_n[7] 0.28fF
C13056 a_7894_7150# VDD 0.23fF
C13057 a_18938_7150# rowoff_n[5] 0.24fF
C13058 a_2346_7192# a_24050_7150# 0.19fF
C13059 a_1962_7190# a_22346_7190# 0.14fF
C13060 a_30074_8154# a_30074_7150# 1.00fF
C13061 a_1962_10202# col_n[21] 0.13fF
C13062 a_10998_3134# col[8] 0.29fF
C13063 a_31382_9198# vcm 0.22fF
C13064 a_31078_17190# a_32082_17190# 0.97fF
C13065 a_28066_12170# col_n[25] 0.28fF
C13066 a_8990_4138# rowon_n[2] 0.14fF
C13067 a_28978_5142# rowoff_n[3] 0.24fF
C13068 a_1962_4178# col[12] 0.11fF
C13069 a_13006_3134# ctop 3.57fF
C13070 a_1962_17230# col[14] 0.11fF
C13071 a_20946_11166# VDD 0.23fF
C13072 m3_8892_1078# m3_9896_1078# 0.22fF
C13073 a_19942_9158# a_20034_9158# 0.26fF
C13074 m2_1732_13998# sample 0.19fF
C13075 m2_34864_7974# ctop 0.17fF
C13076 a_2346_1168# a_13918_1126# 0.35fF
C13077 a_26058_6146# m2_26256_6394# 0.16fF
C13078 a_26058_7150# ctop 3.58fF
C13079 a_13006_17190# rowon_n[15] 0.14fF
C13080 a_33998_15182# VDD 0.23fF
C13081 m2_1732_10986# rowon_n[9] 0.11fF
C13082 m2_21812_946# a_1962_1166# 0.18fF
C13083 a_22042_17190# m3_21944_18146# 0.15fF
C13084 a_2966_15182# row_n[13] 0.16fF
C13085 a_28066_7150# rowon_n[5] 0.14fF
C13086 a_6982_6146# vcm 0.62fF
C13087 a_10998_5142# col_n[8] 0.28fF
C13088 m2_34864_11990# m2_35292_12418# 0.16fF
C13089 a_2346_3176# a_26970_3134# 0.35fF
C13090 a_14010_3134# a_15014_3134# 0.97fF
C13091 m2_33860_946# col_n[31] 0.62fF
C13092 a_1962_6186# col_n[12] 0.13fF
C13093 m2_1732_18014# vcm 0.27fF
C13094 a_32994_13174# a_33086_13174# 0.26fF
C13095 a_16018_13174# a_16018_12170# 1.00fF
C13096 a_5978_7150# row_n[5] 0.17fF
C13097 a_2966_3134# col_n[0] 0.28fF
C13098 a_27062_11166# rowoff_n[9] 0.10fF
C13099 a_20034_10162# vcm 0.62fF
C13100 a_1962_17230# a_14010_17190# 0.27fF
C13101 a_26058_15182# col[23] 0.29fF
C13102 m2_21812_18014# m2_22240_18442# 0.16fF
C13103 a_1962_13214# col[5] 0.11fF
C13104 a_23046_3134# VDD 0.52fF
C13105 a_1962_11206# m2_1732_10986# 0.15fF
C13106 a_2346_12212# col[25] 0.15fF
C13107 a_13310_4178# vcm 0.22fF
C13108 a_2346_14220# a_8990_14178# 0.19fF
C13109 a_1962_14218# a_7286_14218# 0.14fF
C13110 a_5886_14178# a_5978_14178# 0.26fF
C13111 a_33086_14178# vcm 0.62fF
C13112 a_1962_2170# a_34090_2130# 0.27fF
C13113 a_23046_7150# m2_23244_7398# 0.16fF
C13114 a_2346_6188# VDD 32.63fF
C13115 a_27062_7150# a_28066_7150# 0.97fF
C13116 a_25054_10162# row_n[8] 0.17fF
C13117 a_2874_11166# a_2966_11166# 0.26fF
C13118 a_2346_11208# a_3878_11166# 0.35fF
C13119 a_8990_8154# col[6] 0.29fF
C13120 a_26362_8194# vcm 0.22fF
C13121 a_2346_16228# a_22042_16186# 0.19fF
C13122 a_29070_17190# a_29070_16186# 1.00fF
C13123 a_1962_16226# a_20338_16226# 0.14fF
C13124 a_7986_2130# ctop 3.39fF
C13125 a_1962_18234# m2_7756_18014# 0.18fF
C13126 a_1962_2170# col_n[3] 0.13fF
C13127 a_15926_10162# VDD 0.23fF
C13128 a_26058_17190# col_n[23] 0.28fF
C13129 a_1962_15222# col_n[5] 0.13fF
C13130 a_27062_4138# col[24] 0.29fF
C13131 a_14922_12170# rowoff_n[10] 0.24fF
C13132 a_13006_8154# rowon_n[6] 0.14fF
C13133 a_21038_6146# ctop 3.58fF
C13134 m3_7888_1078# VDD 0.14fF
C13135 a_2346_18236# m2_2736_18014# 0.20fF
C13136 a_28978_14178# VDD 0.23fF
C13137 a_2966_6146# row_n[4] 0.16fF
C13138 a_2346_10204# a_11910_10162# 0.35fF
C13139 a_11910_2130# rowoff_n[0] 0.24fF
C13140 VDD rowon_n[9] 2.61fF
C13141 vcm rowon_n[11] 0.50fF
C13142 col_n[0] row_n[11] 0.23fF
C13143 col_n[5] row_n[14] 0.23fF
C13144 col_n[1] row_n[12] 0.23fF
C13145 col_n[3] row_n[13] 0.23fF
C13146 col_n[7] row_n[15] 0.23fF
C13147 a_2346_8196# col[16] 0.15fF
C13148 col[28] rowoff_n[15] 0.11fF
C13149 a_34394_6186# vcm 0.22fF
C13150 a_28978_16186# rowoff_n[14] 0.24fF
C13151 m2_29844_18014# ctop 0.18fF
C13152 a_20034_8154# m2_20232_8402# 0.16fF
C13153 a_28978_3134# a_29070_3134# 0.26fF
C13154 a_12002_3134# a_12002_2130# 1.00fF
C13155 a_8990_10162# col_n[6] 0.28fF
C13156 a_34090_10162# ctop 3.42fF
C13157 a_1962_7190# a_5978_7150# 0.27fF
C13158 a_7986_17190# VDD 0.55fF
C13159 a_13006_12170# a_14010_12170# 0.97fF
C13160 a_2346_12212# a_24962_12170# 0.35fF
C13161 a_1962_4178# col[23] 0.11fF
C13162 m2_16792_946# m3_16924_1078# 2.79fF
C13163 a_32082_11166# rowon_n[9] 0.14fF
C13164 a_15014_9158# vcm 0.62fF
C13165 a_1962_17230# col[25] 0.11fF
C13166 a_27062_6146# col_n[24] 0.28fF
C13167 a_18026_2130# VDD 0.54fF
C13168 a_1962_11206# VDD 2.73fF
C13169 m2_27836_946# m3_28972_1078# 0.13fF
C13170 m3_1864_15134# m3_1864_14130# 0.22fF
C13171 a_1962_9198# a_19030_9158# 0.27fF
C13172 a_8290_3174# vcm 0.22fF
C13173 a_9994_11166# row_n[9] 0.17fF
C13174 a_2966_14178# a_2966_13174# 1.00fF
C13175 a_28066_13174# vcm 0.62fF
C13176 a_31078_6146# VDD 0.52fF
C13177 a_25054_7150# a_25054_6146# 1.00fF
C13178 a_1962_6186# a_12306_6186# 0.14fF
C13179 a_2346_6188# a_14010_6146# 0.19fF
C13180 a_9994_8154# rowoff_n[6] 0.10fF
C13181 a_1962_11206# a_32082_11166# 0.27fF
C13182 a_2346_4180# col[7] 0.15fF
C13183 a_2346_17232# col[9] 0.15fF
C13184 a_21342_7190# vcm 0.22fF
C13185 a_26058_16186# a_27062_16186# 0.97fF
C13186 a_16018_17190# rowoff_n[15] 0.10fF
C13187 a_1962_6186# col_n[23] 0.13fF
C13188 a_20034_6146# rowoff_n[4] 0.10fF
C13189 a_6982_13174# col[4] 0.29fF
C13190 a_17022_9158# m2_17220_9406# 0.16fF
C13191 a_10906_9158# VDD 0.23fF
C13192 a_14922_8154# a_15014_8154# 0.26fF
C13193 a_2346_8196# a_27062_8154# 0.19fF
C13194 a_1962_8194# a_25358_8194# 0.14fF
C13195 a_29070_14178# row_n[12] 0.17fF
C13196 a_1962_13214# col[16] 0.11fF
C13197 m2_6752_946# ctop 0.18fF
C13198 a_35398_11206# vcm 0.23fF
C13199 a_30074_4138# rowoff_n[2] 0.10fF
C13200 a_25054_9158# col[22] 0.29fF
C13201 m2_3740_18014# m2_4744_18014# 0.96fF
C13202 a_16018_5142# ctop 3.58fF
C13203 a_23958_13174# VDD 0.23fF
C13204 a_17022_12170# rowon_n[10] 0.14fF
C13205 a_8990_2130# a_9994_2130# 0.97fF
C13206 a_2346_2172# a_16930_2130# 0.35fF
C13207 m2_34864_18014# m3_34996_17142# 0.15fF
C13208 a_29070_9158# ctop 3.58fF
C13209 a_32082_2130# rowon_n[0] 0.14fF
C13210 a_2874_16186# VDD 0.24fF
C13211 a_6982_15182# col_n[4] 0.28fF
C13212 a_27974_12170# a_28066_12170# 0.26fF
C13213 a_10998_12170# a_10998_11166# 1.00fF
C13214 a_2346_13216# col[0] 0.15fF
C13215 a_7986_2130# col[5] 0.29fF
C13216 a_9994_8154# vcm 0.62fF
C13217 a_1962_16226# a_3970_16186# 0.27fF
C13218 a_1962_2170# col_n[14] 0.13fF
C13219 a_1962_15222# col_n[16] 0.13fF
C13220 a_2346_4180# a_29982_4138# 0.35fF
C13221 a_14010_10162# m2_14208_10410# 0.16fF
C13222 a_25054_11166# col_n[22] 0.28fF
C13223 a_9994_2130# row_n[0] 0.17fF
C13224 a_3270_2170# vcm 0.23fF
C13225 a_28978_10162# rowoff_n[8] 0.24fF
C13226 a_1962_9198# col[7] 0.11fF
C13227 a_23046_12170# vcm 0.62fF
C13228 a_30986_13174# rowoff_n[11] 0.24fF
C13229 a_35002_6146# m2_34864_5966# 0.16fF
C13230 a_2966_6146# ctop 3.42fF
C13231 a_26058_5142# VDD 0.52fF
C13232 m3_3872_18146# VDD 0.30fF
C13233 a_22042_6146# a_23046_6146# 0.97fF
C13234 col_n[10] row_n[11] 0.23fF
C13235 col_n[18] row_n[15] 0.23fF
C13236 col_n[8] row_n[10] 0.23fF
C13237 col_n[16] row_n[14] 0.23fF
C13238 sample row_n[5] 1.03fF
C13239 vcm row_n[6] 0.49fF
C13240 col_n[14] row_n[13] 0.23fF
C13241 col_n[2] row_n[7] 0.23fF
C13242 VDD row_n[4] 2.93fF
C13243 col_n[12] row_n[12] 0.23fF
C13244 col_n[4] row_n[8] 0.23fF
C13245 col_n[6] row_n[9] 0.23fF
C13246 col_n[25] col_n[26] 0.10fF
C13247 a_2346_8196# col[27] 0.15fF
C13248 a_14010_15182# row_n[13] 0.17fF
C13249 a_16322_6186# vcm 0.22fF
C13250 a_1962_15222# a_10298_15222# 0.14fF
C13251 a_24050_16186# a_24050_15182# 1.00fF
C13252 a_2346_15224# a_12002_15182# 0.19fF
C13253 a_2346_15224# vcm 0.40fF
C13254 m2_34864_13998# VDD 1.03fF
C13255 m2_21812_946# m2_22240_1374# 0.16fF
C13256 a_29070_5142# row_n[3] 0.17fF
C13257 a_7986_4138# col_n[5] 0.28fF
C13258 m2_2736_1950# col[0] 0.28fF
C13259 a_5886_8154# VDD 0.23fF
C13260 a_29374_10202# vcm 0.22fF
C13261 a_1962_17230# a_23350_17230# 0.14fF
C13262 a_2346_17232# a_25054_17190# 0.19fF
C13263 a_13918_17190# a_14010_17190# 0.26fF
C13264 a_1962_11206# col_n[7] 0.13fF
C13265 a_10998_4138# ctop 3.58fF
C13266 m3_10900_1078# ctop 0.23fF
C13267 m2_14784_18014# col_n[12] 0.25fF
C13268 a_10998_11166# m2_11196_11414# 0.16fF
C13269 a_23046_14178# col[20] 0.29fF
C13270 a_18938_12170# VDD 0.23fF
C13271 m3_4876_18146# m3_5880_18146# 0.22fF
C13272 a_3878_18194# VDD 0.33fF
C13273 a_17022_3134# rowon_n[1] 0.14fF
C13274 a_2874_3134# rowoff_n[1] 0.24fF
C13275 m2_1732_10986# ctop 0.17fF
C13276 a_18026_14178# rowoff_n[12] 0.10fF
C13277 a_23958_2130# a_24050_2130# 0.26fF
C13278 a_24050_8154# ctop 3.58fF
C13279 m2_34864_15002# m3_34996_14130# 0.15fF
C13280 a_2346_4180# col[18] 0.15fF
C13281 a_2346_17232# col[20] 0.15fF
C13282 a_31990_16186# VDD 0.23fF
C13283 a_2346_11208# a_14922_11166# 0.35fF
C13284 a_7986_11166# a_8990_11166# 0.97fF
C13285 a_4974_7150# vcm 0.62fF
C13286 a_18026_2130# m2_18224_2378# 0.16fF
C13287 a_21038_16186# rowon_n[14] 0.14fF
C13288 a_5978_7150# col[3] 0.29fF
C13289 a_2966_9158# m2_1732_8978# 0.96fF
C13290 m2_4744_946# col_n[2] 0.37fF
C13291 a_1962_8194# a_8990_8154# 0.27fF
C13292 a_1962_13214# col[27] 0.11fF
C13293 a_2346_13216# a_27974_13174# 0.35fF
C13294 rowon_n[2] rowoff_n[2] 20.27fF
C13295 a_23046_16186# col_n[20] 0.28fF
C13296 a_18026_11166# vcm 0.62fF
C13297 a_24050_3134# col[21] 0.29fF
C13298 a_1962_7190# sample 0.14fF
C13299 a_21038_4138# VDD 0.52fF
C13300 a_2346_5184# a_3970_5142# 0.19fF
C13301 a_20034_6146# a_20034_5142# 1.00fF
C13302 a_7986_12170# m2_8184_12418# 0.16fF
C13303 a_14010_6146# row_n[4] 0.17fF
C13304 a_1962_10202# a_22042_10162# 0.27fF
C13305 a_11302_5182# vcm 0.22fF
C13306 a_21038_15182# a_22042_15182# 0.97fF
C13307 a_5886_15182# rowoff_n[13] 0.24fF
C13308 a_31078_15182# vcm 0.62fF
C13309 m2_11772_18014# m3_11904_18146# 2.79fF
C13310 a_34090_8154# VDD 0.54fF
C13311 a_11910_7150# rowoff_n[5] 0.24fF
C13312 a_2346_13216# col[11] 0.15fF
C13313 a_1962_7190# a_15318_7190# 0.14fF
C13314 a_9902_7150# a_9994_7150# 0.26fF
C13315 a_2346_7192# a_17022_7150# 0.19fF
C13316 a_5978_9158# col_n[3] 0.28fF
C13317 a_1962_2170# col_n[25] 0.13fF
C13318 a_24354_9198# vcm 0.22fF
C13319 a_1962_15222# col_n[27] 0.13fF
C13320 a_21950_5142# rowoff_n[3] 0.24fF
C13321 a_5978_3134# ctop 3.57fF
C13322 a_33086_9158# row_n[7] 0.17fF
C13323 a_24050_5142# col_n[21] 0.28fF
C13324 a_13918_11166# VDD 0.23fF
C13325 a_1962_9198# col[18] 0.11fF
C13326 a_2346_9200# a_30074_9158# 0.19fF
C13327 a_33086_10162# a_33086_9158# 1.00fF
C13328 a_1962_9198# a_28370_9198# 0.14fF
C13329 a_31990_3134# rowoff_n[1] 0.24fF
C13330 VDD ctop 92.86fF
C13331 col_n[29] row_n[15] 0.23fF
C13332 col_n[15] row_n[8] 0.23fF
C13333 col_n[17] row_n[9] 0.23fF
C13334 col_n[11] row_n[6] 0.23fF
C13335 col_n[9] row_n[5] 0.23fF
C13336 vcm rowon_n[0] 0.50fF
C13337 col_n[23] row_n[12] 0.23fF
C13338 col_n[3] row_n[2] 0.23fF
C13339 col_n[27] row_n[14] 0.23fF
C13340 col_n[21] row_n[11] 0.23fF
C13341 col_n[5] row_n[3] 0.23fF
C13342 col_n[1] row_n[1] 0.23fF
C13343 col_n[19] row_n[10] 0.23fF
C13344 col_n[7] row_n[4] 0.23fF
C13345 col_n[0] row_n[0] 0.23fF
C13346 col_n[25] row_n[13] 0.23fF
C13347 a_2346_1168# a_6890_1126# 0.35fF
C13348 col_n[13] row_n[7] 0.23fF
C13349 m2_34864_11990# m3_34996_11118# 0.15fF
C13350 a_19030_7150# ctop 3.58fF
C13351 a_4974_13174# m2_5172_13422# 0.16fF
C13352 a_5978_17190# rowon_n[15] 0.14fF
C13353 a_26970_15182# VDD 0.23fF
C13354 a_22954_11166# a_23046_11166# 0.26fF
C13355 a_5978_11166# a_5978_10162# 1.00fF
C13356 a_21038_7150# rowon_n[5] 0.14fF
C13357 a_2346_3176# a_19942_3134# 0.35fF
C13358 a_32082_2130# m2_31852_946# 0.99fF
C13359 a_2346_1168# m2_23820_946# 0.19fF
C13360 a_32082_11166# ctop 3.58fF
C13361 a_10998_2130# m3_10900_1078# 0.15fF
C13362 a_2346_9200# col[2] 0.15fF
C13363 a_2966_11166# m3_1864_11118# 0.14fF
C13364 a_3970_12170# col[1] 0.29fF
C13365 a_1962_18234# col_n[1] 0.13fF
C13366 a_1962_11206# col_n[18] 0.13fF
C13367 a_20034_11166# rowoff_n[9] 0.10fF
C13368 a_13006_10162# vcm 0.62fF
C13369 a_1962_17230# a_6982_17190# 0.27fF
C13370 m2_14784_18014# m2_15212_18442# 0.16fF
C13371 a_16018_3134# VDD 0.52fF
C13372 m3_6884_18146# ctop 0.23fF
C13373 a_17022_5142# a_18026_5142# 0.97fF
C13374 a_2346_5184# a_32994_5142# 0.35fF
C13375 a_22042_8154# col[19] 0.29fF
C13376 a_1962_5182# col[9] 0.11fF
C13377 a_30074_9158# rowoff_n[7] 0.10fF
C13378 a_6282_4178# vcm 0.22fF
C13379 a_19030_15182# a_19030_14178# 1.00fF
C13380 a_26058_14178# vcm 0.62fF
C13381 a_34090_15182# rowoff_n[13] 0.10fF
C13382 a_2346_4180# col[29] 0.15fF
C13383 a_1962_2170# a_27062_2130# 0.27fF
C13384 a_2346_17232# col[31] 0.15fF
C13385 a_29070_7150# VDD 0.52fF
C13386 m2_33860_946# sw 0.32fF
C13387 a_18026_10162# row_n[8] 0.17fF
C13388 a_19334_8194# vcm 0.22fF
C13389 a_2346_16228# a_15014_16186# 0.19fF
C13390 a_8898_16186# a_8990_16186# 0.26fF
C13391 a_1962_16226# a_13310_16226# 0.14fF
C13392 a_3970_14178# col_n[1] 0.28fF
C13393 a_2966_16186# rowon_n[14] 0.13fF
C13394 a_8898_10162# VDD 0.23fF
C13395 col[0] rowoff_n[5] 0.11fF
C13396 col[1] rowoff_n[6] 0.11fF
C13397 col[4] rowoff_n[9] 0.11fF
C13398 col[3] rowoff_n[8] 0.11fF
C13399 col[2] rowoff_n[7] 0.11fF
C13400 a_30074_9158# a_31078_9158# 0.97fF
C13401 a_22042_10162# col_n[19] 0.28fF
C13402 a_1962_7190# col_n[9] 0.13fF
C13403 a_32386_12210# vcm 0.22fF
C13404 a_7894_12170# rowoff_n[10] 0.24fF
C13405 a_18938_1126# a_19030_1126# 0.27fF
C13406 a_1962_5182# m2_34864_4962# 0.17fF
C13407 a_5978_8154# rowon_n[6] 0.14fF
C13408 a_1962_1166# a_35398_1166# 0.14fF
C13409 m2_34864_8978# m3_34996_8106# 0.15fF
C13410 a_14010_6146# ctop 3.58fF
C13411 a_2966_4138# VDD 0.56fF
C13412 m3_34996_12122# VDD 0.26fF
C13413 a_1962_1166# col[0] 0.11fF
C13414 a_21950_14178# VDD 0.23fF
C13415 a_1962_14218# col[2] 0.11fF
C13416 m2_34864_3958# vcm 0.51fF
C13417 a_2346_10204# a_4882_10162# 0.35fF
C13418 a_4882_2130# rowoff_n[0] 0.24fF
C13419 a_21950_16186# rowoff_n[14] 0.24fF
C13420 m2_15788_18014# ctop 0.18fF
C13421 a_2346_13216# col[22] 0.15fF
C13422 a_27062_10162# ctop 3.58fF
C13423 a_28978_1126# m2_28840_946# 0.16fF
C13424 a_33086_16186# m2_33284_16434# 0.16fF
C13425 a_4974_3134# col_n[2] 0.28fF
C13426 a_35002_18194# VDD 0.40fF
C13427 a_2346_12212# a_17934_12170# 0.35fF
C13428 a_25054_11166# rowon_n[9] 0.14fF
C13429 a_7986_9158# vcm 0.62fF
C13430 a_1962_17230# a_34394_17230# 0.14fF
C13431 a_3878_5142# rowoff_n[3] 0.24fF
C13432 a_10998_2130# VDD 0.55fF
C13433 a_1962_9198# col[29] 0.11fF
C13434 a_31990_5142# a_32082_5142# 0.26fF
C13435 a_15014_5142# a_15014_4138# 1.00fF
C13436 a_1962_9198# a_12002_9158# 0.27fF
C13437 a_20034_13174# col[17] 0.29fF
C13438 a_1962_3174# vcm 6.95fF
C13439 a_16018_14178# a_17022_14178# 0.97fF
C13440 a_2346_14220# a_30986_14178# 0.35fF
C13441 col_n[30] row_n[10] 0.23fF
C13442 col_n[7] ctop 2.02fF
C13443 rowon_n[13] row_n[13] 19.75fF
C13444 VDD col[5] 4.19fF
C13445 col_n[24] row_n[7] 0.23fF
C13446 col_n[22] row_n[6] 0.23fF
C13447 col_n[18] row_n[4] 0.23fF
C13448 col_n[14] row_n[2] 0.23fF
C13449 a_1962_16226# col_n[2] 0.13fF
C13450 col_n[20] row_n[5] 0.23fF
C13451 col_n[28] row_n[9] 0.23fF
C13452 col_n[26] row_n[8] 0.23fF
C13453 col_n[10] row_n[0] 0.23fF
C13454 col_n[12] row_n[1] 0.23fF
C13455 vcm col[1] 5.84fF
C13456 col_n[16] row_n[3] 0.23fF
C13457 a_21038_13174# vcm 0.62fF
C13458 m2_29844_18014# col[27] 0.28fF
C13459 a_24050_6146# VDD 0.52fF
C13460 a_1962_6186# a_5278_6186# 0.14fF
C13461 a_2346_6188# a_6982_6146# 0.19fF
C13462 a_4882_6146# a_4974_6146# 0.26fF
C13463 a_2874_8154# rowoff_n[6] 0.24fF
C13464 a_1962_11206# a_25054_11166# 0.27fF
C13465 a_2966_7150# rowon_n[5] 0.13fF
C13466 a_14314_7190# vcm 0.22fF
C13467 m2_1732_5966# sample_n 0.15fF
C13468 a_2346_9200# col[13] 0.15fF
C13469 a_8990_17190# rowoff_n[15] 0.10fF
C13470 a_34090_17190# vcm 0.60fF
C13471 m2_1732_17010# VDD 1.04fF
C13472 a_13006_6146# rowoff_n[4] 0.10fF
C13473 a_1962_18234# col_n[12] 0.13fF
C13474 a_30074_17190# m2_30272_17438# 0.16fF
C13475 a_28066_9158# a_28066_8154# 1.00fF
C13476 a_2346_8196# a_20034_8154# 0.19fF
C13477 a_1962_8194# a_18330_8194# 0.14fF
C13478 a_22042_14178# row_n[12] 0.17fF
C13479 a_1962_11206# col_n[29] 0.13fF
C13480 m2_34864_2954# m2_34864_1950# 0.99fF
C13481 a_23046_4138# rowoff_n[2] 0.10fF
C13482 a_27366_11206# vcm 0.22fF
C13483 a_20034_15182# col_n[17] 0.28fF
C13484 a_32082_5142# m2_32280_5390# 0.16fF
C13485 a_1962_5182# col[20] 0.11fF
C13486 m2_34864_5966# m3_34996_5094# 0.15fF
C13487 a_8990_5142# ctop 3.58fF
C13488 m2_14784_946# vcm 0.42fF
C13489 a_21038_2130# col[18] 0.29fF
C13490 a_16930_13174# VDD 0.23fF
C13491 a_1962_10202# a_31382_10202# 0.14fF
C13492 a_17934_10162# a_18026_10162# 0.26fF
C13493 a_2346_10204# a_33086_10162# 0.19fF
C13494 a_33086_2130# rowoff_n[0] 0.10fF
C13495 m2_31852_946# vcm 0.42fF
C13496 a_9994_12170# rowon_n[10] 0.14fF
C13497 a_2966_7150# m2_3164_7398# 0.16fF
C13498 a_2346_2172# a_9902_2130# 0.35fF
C13499 m2_25828_18014# m3_26964_18146# 0.13fF
C13500 a_22042_9158# ctop 3.58fF
C13501 a_29982_17190# VDD 0.24fF
C13502 a_25054_2130# rowon_n[0] 0.14fF
C13503 a_2346_5184# col[4] 0.15fF
C13504 m2_1732_15002# m2_2160_15430# 0.16fF
C13505 col[10] rowoff_n[4] 0.11fF
C13506 col[9] rowoff_n[3] 0.11fF
C13507 col[14] rowoff_n[8] 0.11fF
C13508 col[13] rowoff_n[7] 0.11fF
C13509 col[15] rowoff_n[9] 0.11fF
C13510 col[8] rowoff_n[2] 0.11fF
C13511 col[7] rowoff_n[1] 0.11fF
C13512 col[6] rowoff_n[0] 0.11fF
C13513 col[11] rowoff_n[5] 0.11fF
C13514 col[12] rowoff_n[6] 0.11fF
C13515 a_2346_4180# a_22954_4138# 0.35fF
C13516 a_12002_4138# a_13006_4138# 0.97fF
C13517 m2_1732_1950# rowon_n[0] 0.11fF
C13518 a_5978_17190# m2_5748_18014# 1.00fF
C13519 a_1962_7190# col_n[20] 0.13fF
C13520 a_21038_4138# col_n[18] 0.28fF
C13521 a_30986_14178# a_31078_14178# 0.26fF
C13522 a_14010_14178# a_14010_13174# 1.00fF
C13523 a_21950_10162# rowoff_n[8] 0.24fF
C13524 a_29070_15182# rowon_n[13] 0.14fF
C13525 a_23958_13174# rowoff_n[11] 0.24fF
C13526 a_16018_12170# vcm 0.62fF
C13527 a_29070_6146# m2_29268_6394# 0.16fF
C13528 a_1962_1166# col[11] 0.11fF
C13529 a_1962_14218# col[13] 0.11fF
C13530 a_19030_5142# VDD 0.52fF
C13531 a_31990_8154# rowoff_n[6] 0.24fF
C13532 a_3878_14178# VDD 0.23fF
C13533 a_2966_11166# col[0] 0.29fF
C13534 a_25054_17190# m3_24956_18146# 0.15fF
C13535 VDD rowoff_n[14] 1.17fF
C13536 a_6982_15182# row_n[13] 0.17fF
C13537 a_9294_6186# vcm 0.22fF
C13538 a_2346_15224# a_4974_15182# 0.19fF
C13539 a_1962_15222# a_3270_15222# 0.14fF
C13540 a_29070_16186# vcm 0.62fF
C13541 a_3878_16186# rowoff_n[14] 0.24fF
C13542 a_22042_5142# row_n[3] 0.17fF
C13543 a_34090_9158# m2_34864_8978# 0.96fF
C13544 a_1962_3174# a_30074_3134# 0.27fF
C13545 a_32082_9158# VDD 0.52fF
C13546 a_25054_8154# a_26058_8154# 0.97fF
C13547 a_22346_10202# vcm 0.22fF
C13548 a_2346_17232# a_18026_17190# 0.19fF
C13549 a_1962_17230# a_16322_17230# 0.14fF
C13550 a_3970_4138# ctop 3.57fF
C13551 m3_1864_10114# ctop 0.23fF
C13552 a_11910_12170# VDD 0.23fF
C13553 a_1962_3174# col_n[11] 0.13fF
C13554 col_n[29] row_n[4] 0.23fF
C13555 col_n[21] row_n[0] 0.23fF
C13556 col_n[6] col[6] 0.72fF
C13557 VDD col[16] 4.16fF
C13558 vcm col[12] 5.84fF
C13559 col_n[31] row_n[5] 0.23fF
C13560 col_n[25] row_n[2] 0.23fF
C13561 col_n[18] ctop 2.02fF
C13562 col_n[23] row_n[1] 0.23fF
C13563 col_n[27] row_n[3] 0.23fF
C13564 a_1962_16226# col_n[13] 0.13fF
C13565 a_19030_7150# col[16] 0.29fF
C13566 a_9994_3134# rowon_n[1] 0.14fF
C13567 a_2966_13174# vcm 0.61fF
C13568 a_10998_14178# rowoff_n[12] 0.10fF
C13569 a_26058_7150# m2_26256_7398# 0.16fF
C13570 a_1962_10202# col[4] 0.11fF
C13571 a_17022_8154# ctop 3.58fF
C13572 a_24962_16186# VDD 0.23fF
C13573 a_2346_11208# a_7894_11166# 0.35fF
C13574 a_2346_9200# col[24] 0.15fF
C13575 a_4974_2130# m2_4744_946# 0.99fF
C13576 a_14010_16186# rowon_n[14] 0.14fF
C13577 a_1962_18234# col_n[23] 0.13fF
C13578 a_26970_4138# a_27062_4138# 0.26fF
C13579 a_9994_4138# a_9994_3134# 1.00fF
C13580 a_30074_12170# ctop 3.58fF
C13581 a_25054_17190# m2_24824_18014# 1.00fF
C13582 a_29070_6146# rowon_n[4] 0.14fF
C13583 a_10998_13174# a_12002_13174# 0.97fF
C13584 a_2346_13216# a_20946_13174# 0.35fF
C13585 a_1962_5182# col[31] 0.11fF
C13586 a_10998_11166# vcm 0.62fF
C13587 m2_27836_946# col_n[25] 0.32fF
C13588 a_19030_9158# col_n[16] 0.28fF
C13589 a_14010_4138# VDD 0.52fF
C13590 m2_16792_946# col[14] 0.39fF
C13591 m3_22948_1078# VDD 0.14fF
C13592 a_1962_12210# m2_1732_11990# 0.15fF
C13593 a_6982_6146# row_n[4] 0.17fF
C13594 a_1962_12210# col_n[4] 0.13fF
C13595 a_1962_10202# a_15014_10162# 0.27fF
C13596 a_4274_5182# vcm 0.22fF
C13597 a_2346_15224# a_33998_15182# 0.35fF
C13598 a_24050_15182# vcm 0.62fF
C13599 a_23046_8154# m2_23244_8402# 0.16fF
C13600 m2_2736_18014# m3_1864_18146# 0.13fF
C13601 a_27062_8154# VDD 0.52fF
C13602 a_4882_7150# rowoff_n[5] 0.24fF
C13603 a_1962_7190# a_8290_7190# 0.14fF
C13604 a_2346_7192# a_9994_7150# 0.19fF
C13605 a_23046_8154# a_23046_7150# 1.00fF
C13606 a_1962_12210# a_28066_12170# 0.27fF
C13607 a_2346_5184# col[15] 0.15fF
C13608 a_17326_9198# vcm 0.22fF
C13609 a_24050_17190# a_25054_17190# 0.97fF
C13610 col[17] rowoff_n[0] 0.11fF
C13611 col[20] rowoff_n[3] 0.11fF
C13612 col[23] rowoff_n[6] 0.11fF
C13613 col[26] rowoff_n[9] 0.11fF
C13614 col[25] rowoff_n[8] 0.11fF
C13615 col[18] rowoff_n[1] 0.11fF
C13616 col[19] rowoff_n[2] 0.11fF
C13617 col[24] rowoff_n[7] 0.11fF
C13618 col[22] rowoff_n[5] 0.11fF
C13619 col[21] rowoff_n[4] 0.11fF
C13620 a_14922_5142# rowoff_n[3] 0.24fF
C13621 a_26058_9158# row_n[7] 0.17fF
C13622 a_1962_7190# col_n[31] 0.13fF
C13623 a_2966_4138# a_3970_4138# 0.97fF
C13624 a_34090_5142# m3_34996_5094# 0.13fF
C13625 a_6890_11166# VDD 0.23fF
C13626 a_1962_9198# a_21342_9198# 0.14fF
C13627 a_2346_9200# a_23046_9158# 0.19fF
C13628 a_12914_9158# a_13006_9158# 0.26fF
C13629 a_24962_3134# rowoff_n[1] 0.24fF
C13630 a_3878_10162# rowoff_n[8] 0.24fF
C13631 a_1962_1166# col[22] 0.11fF
C13632 a_1962_14218# col[24] 0.11fF
C13633 a_30378_13214# vcm 0.22fF
C13634 a_17022_12170# col[14] 0.29fF
C13635 a_12002_7150# ctop 3.58fF
C13636 a_19942_15182# VDD 0.23fF
C13637 m2_1732_6970# vcm 0.45fF
C13638 a_2346_11208# a_2346_10204# 0.22fF
C13639 a_1962_11206# a_35398_11206# 0.14fF
C13640 col[10] rowoff_n[10] 0.11fF
C13641 a_14010_7150# rowon_n[5] 0.14fF
C13642 a_20034_9158# m2_20232_9406# 0.16fF
C13643 a_2346_3176# a_12914_3134# 0.35fF
C13644 a_6982_3134# a_7986_3134# 0.97fF
C13645 a_25054_11166# ctop 3.58fF
C13646 a_2346_1168# col[6] 0.14fF
C13647 a_8990_13174# a_8990_12170# 1.00fF
C13648 a_25966_13174# a_26058_13174# 0.26fF
C13649 a_2346_14220# col[8] 0.15fF
C13650 m2_1732_946# m2_2736_946# 0.96fF
C13651 a_5978_10162# vcm 0.62fF
C13652 a_13006_11166# rowoff_n[9] 0.10fF
C13653 m2_7756_18014# m2_8184_18442# 0.16fF
C13654 a_1962_3174# col_n[22] 0.13fF
C13655 a_8990_3134# VDD 0.52fF
C13656 col_n[29] ctop 2.02fF
C13657 col_n[11] col[12] 5.98fF
C13658 vcm col[23] 5.84fF
C13659 VDD col[27] 4.17fF
C13660 a_2346_5184# a_25966_5142# 0.35fF
C13661 a_1962_16226# col_n[24] 0.13fF
C13662 a_17022_14178# col_n[14] 0.28fF
C13663 a_33086_10162# rowon_n[8] 0.14fF
C13664 a_18026_1126# col[15] 0.38fF
C13665 ctop rowoff_n[11] 0.60fF
C13666 a_23046_9158# rowoff_n[7] 0.10fF
C13667 a_1962_10202# col[15] 0.11fF
C13668 a_19030_14178# vcm 0.62fF
C13669 a_27062_15182# rowoff_n[13] 0.10fF
C13670 a_1962_2170# a_20034_2130# 0.27fF
C13671 a_22042_7150# VDD 0.52fF
C13672 a_33086_7150# rowoff_n[5] 0.10fF
C13673 a_20034_7150# a_21038_7150# 0.97fF
C13674 a_10998_10162# row_n[8] 0.17fF
C13675 a_12306_8194# vcm 0.22fF
C13676 a_1962_16226# a_6282_16226# 0.14fF
C13677 a_2346_16228# a_7986_16186# 0.19fF
C13678 a_22042_17190# a_22042_16186# 1.00fF
C13679 a_32082_18194# vcm 0.12fF
C13680 a_17022_10162# m2_17220_10410# 0.16fF
C13681 a_1962_4178# a_33086_4138# 0.27fF
C13682 a_2346_13216# a_1962_13214# 2.62fF
C13683 a_25358_12210# vcm 0.22fF
C13684 a_18026_3134# col_n[15] 0.28fF
C13685 a_1962_1166# a_26362_1166# 0.14fF
C13686 a_6982_6146# ctop 3.58fF
C13687 a_1962_12210# col_n[15] 0.13fF
C13688 a_30074_13174# row_n[11] 0.17fF
C13689 m3_18932_18146# VDD 0.37fF
C13690 a_15014_17190# col[12] 0.29fF
C13691 a_14922_14178# VDD 0.23fF
C13692 a_33086_11166# a_34090_11166# 0.97fF
C13693 a_1962_6186# col[6] 0.11fF
C13694 a_14922_16186# rowoff_n[14] 0.24fF
C13695 a_21950_3134# a_22042_3134# 0.26fF
C13696 a_33086_13174# col[30] 0.29fF
C13697 a_4974_3134# a_4974_2130# 1.00fF
C13698 a_20034_10162# ctop 3.58fF
C13699 a_2346_5184# col[26] 0.15fF
C13700 a_27974_18194# VDD 0.33fF
C13701 col[28] rowoff_n[0] 0.11fF
C13702 col[30] rowoff_n[2] 0.11fF
C13703 col[29] rowoff_n[1] 0.11fF
C13704 col[31] rowoff_n[3] 0.11fF
C13705 m2_30848_18014# vcm 0.28fF
C13706 a_2346_12212# a_10906_12170# 0.35fF
C13707 a_5978_12170# a_6982_12170# 0.97fF
C13708 a_18026_11166# rowon_n[9] 0.14fF
C13709 m2_2736_946# m3_1864_1078# 0.13fF
C13710 a_3970_2130# VDD 0.54fF
C13711 m3_25960_1078# ctop 0.23fF
C13712 a_14010_11166# m2_14208_11414# 0.16fF
C13713 a_33086_14178# ctop 3.57fF
C13714 a_4882_18194# m2_4744_18014# 0.16fF
C13715 a_1962_9198# a_4974_9158# 0.27fF
C13716 a_3878_9158# a_3970_9158# 0.26fF
C13717 a_2346_14220# a_23958_14178# 0.35fF
C13718 a_2346_18236# a_32994_18194# 0.35fF
C13719 a_14010_13174# vcm 0.62fF
C13720 a_16018_6146# col[13] 0.29fF
C13721 a_35002_7150# m2_34864_6970# 0.16fF
C13722 a_1962_8194# col_n[6] 0.13fF
C13723 a_17022_6146# VDD 0.52fF
C13724 a_18026_7150# a_18026_6146# 1.00fF
C13725 col[21] rowoff_n[10] 0.11fF
C13726 a_35494_16548# VDD 0.11fF
C13727 a_33086_15182# col_n[30] 0.28fF
C13728 a_1962_11206# a_18026_11166# 0.27fF
C13729 a_34090_2130# col[31] 0.30fF
C13730 a_7286_7190# vcm 0.22fF
C13731 a_19030_16186# a_20034_16186# 0.97fF
C13732 a_1962_16226# a_1962_15222# 0.16fF
C13733 a_21038_2130# m2_21236_2378# 0.16fF
C13734 a_27062_17190# vcm 0.60fF
C13735 m2_21812_18014# VDD 0.93fF
C13736 a_5978_6146# rowoff_n[4] 0.10fF
C13737 a_30074_10162# VDD 0.52fF
C13738 a_2346_1168# col[17] 0.14fF
C13739 a_1962_8194# a_11302_8194# 0.14fF
C13740 a_7894_8154# a_7986_8154# 0.26fF
C13741 a_2346_8196# a_13006_8154# 0.19fF
C13742 a_2346_14220# col[19] 0.15fF
C13743 a_15014_14178# row_n[12] 0.17fF
C13744 a_1962_13214# a_31078_13174# 0.27fF
C13745 m2_2736_1950# m2_3164_2378# 0.16fF
C13746 a_16018_4138# rowoff_n[2] 0.10fF
C13747 a_30074_4138# row_n[2] 0.17fF
C13748 a_20338_11206# vcm 0.22fF
C13749 a_29070_12170# rowoff_n[10] 0.10fF
C13750 rowon_n[11] ctop 1.40fF
C13751 rowon_n[5] rowon_n[4] 0.15fF
C13752 col_n[17] col[17] 0.64fF
C13753 a_1962_16226# row_n[14] 25.57fF
C13754 a_10998_12170# m2_11196_12418# 0.16fF
C13755 a_16018_8154# col_n[13] 0.28fF
C13756 col[5] rowoff_n[11] 0.11fF
C13757 a_2346_18236# m2_31852_18014# 0.19fF
C13758 a_9902_13174# VDD 0.23fF
C13759 m2_7756_946# vcm 0.42fF
C13760 a_1962_10202# a_24354_10202# 0.14fF
C13761 a_31078_11166# a_31078_10162# 1.00fF
C13762 a_2346_10204# a_26058_10162# 0.19fF
C13763 a_1962_10202# col[26] 0.11fF
C13764 a_26058_2130# rowoff_n[0] 0.10fF
C13765 m2_8760_18014# col_n[6] 0.25fF
C13766 a_33390_15222# vcm 0.22fF
C13767 a_34090_4138# col_n[31] 0.28fF
C13768 a_1962_17230# col_n[0] 0.13fF
C13769 a_15014_9158# ctop 3.58fF
C13770 m2_16792_18014# m3_16924_18146# 2.78fF
C13771 a_34090_17190# row_n[15] 0.17fF
C13772 a_18026_2130# rowon_n[0] 0.14fF
C13773 a_22954_17190# VDD 0.24fF
C13774 a_20946_12170# a_21038_12170# 0.26fF
C13775 a_3970_12170# a_3970_11166# 1.00fF
C13776 a_32994_2130# VDD 0.23fF
C13777 a_2346_4180# a_15926_4138# 0.35fF
C13778 a_2966_10162# m2_1732_9982# 0.96fF
C13779 a_28066_13174# ctop 3.58fF
C13780 a_2346_10204# col[10] 0.15fF
C13781 a_23958_18194# m2_23820_18014# 0.16fF
C13782 a_34090_14178# m3_34996_14130# 0.13fF
C13783 a_14922_10162# rowoff_n[8] 0.24fF
C13784 m2_1732_4962# m2_1732_3958# 0.99fF
C13785 a_22042_15182# rowon_n[13] 0.14fF
C13786 a_1962_12210# col_n[26] 0.13fF
C13787 a_16930_13174# rowoff_n[11] 0.24fF
C13788 a_8990_12170# vcm 0.62fF
C13789 a_12002_5142# VDD 0.52fF
C13790 a_2346_6188# a_28978_6146# 0.35fF
C13791 a_7986_13174# m2_8184_13422# 0.16fF
C13792 a_14010_11166# col[11] 0.29fF
C13793 a_15014_6146# a_16018_6146# 0.97fF
C13794 a_24962_8154# rowoff_n[6] 0.24fF
C13795 a_1962_6186# col[17] 0.11fF
C13796 m2_13780_946# a_1962_1166# 0.18fF
C13797 a_17022_16186# a_17022_15182# 1.00fF
C13798 a_33998_16186# a_34090_16186# 0.26fF
C13799 a_22042_16186# vcm 0.62fF
C13800 a_30986_17190# rowoff_n[15] 0.24fF
C13801 a_32082_7150# col[29] 0.29fF
C13802 a_1962_3174# a_23046_3134# 0.27fF
C13803 a_15014_5142# row_n[3] 0.17fF
C13804 a_35002_6146# rowoff_n[4] 0.24fF
C13805 a_14010_2130# m3_13912_1078# 0.15fF
C13806 a_1962_1166# m2_30848_946# 0.18fF
C13807 a_25054_9158# VDD 0.52fF
C13808 a_32082_1126# vcm 0.12fF
C13809 a_1962_7190# row_n[5] 25.57fF
C13810 a_15318_10202# vcm 0.22fF
C13811 a_2346_17232# a_10998_17190# 0.19fF
C13812 a_1962_17230# a_9294_17230# 0.14fF
C13813 a_6890_17190# a_6982_17190# 0.26fF
C13814 m2_1732_18014# m2_1732_17010# 0.99fF
C13815 m3_21944_18146# ctop 0.23fF
C13816 a_2346_6188# col[1] 0.15fF
C13817 a_4882_12170# VDD 0.23fF
C13818 a_28066_10162# a_29070_10162# 0.97fF
C13819 a_14010_13174# col_n[11] 0.28fF
C13820 a_1962_8194# col_n[17] 0.13fF
C13821 a_34090_8154# row_n[6] 0.17fF
C13822 a_28370_14218# vcm 0.22fF
C13823 a_3970_14178# rowoff_n[12] 0.10fF
C13824 a_16930_2130# a_17022_2130# 0.26fF
C13825 a_1962_2170# a_29374_2170# 0.14fF
C13826 a_2346_2172# a_31078_2130# 0.19fF
C13827 a_9994_8154# ctop 3.58fF
C13828 a_4974_14178# m2_5172_14426# 0.16fF
C13829 a_1962_2170# col[8] 0.11fF
C13830 a_32082_9158# col_n[29] 0.28fF
C13831 a_17934_16186# VDD 0.23fF
C13832 a_1962_15222# col[10] 0.11fF
C13833 a_27974_1126# VDD 0.44fF
C13834 a_6982_16186# rowon_n[14] 0.14fF
C13835 a_2346_1168# col[28] 0.14fF
C13836 a_2346_14220# col[30] 0.15fF
C13837 a_23046_12170# ctop 3.58fF
C13838 a_2346_18236# col[2] 0.14fF
C13839 a_22042_6146# rowon_n[4] 0.14fF
C13840 a_2346_13216# a_13918_13174# 0.35fF
C13841 row_n[6] ctop 1.65fF
C13842 col_n[22] col[23] 5.98fF
C13843 rowon_n[2] row_n[2] 19.75fF
C13844 a_3970_11166# vcm 0.62fF
C13845 col[16] rowoff_n[11] 0.11fF
C13846 a_6982_4138# VDD 0.52fF
C13847 a_15014_2130# col_n[12] 0.28fF
C13848 m3_1864_4090# VDD 0.25fF
C13849 a_29982_6146# a_30074_6146# 0.26fF
C13850 a_13006_6146# a_13006_5142# 1.00fF
C13851 a_2346_15224# ctop 1.59fF
C13852 a_1962_10202# a_7986_10162# 0.27fF
C13853 a_12002_16186# col[9] 0.29fF
C13854 a_14010_15182# a_15014_15182# 0.97fF
C13855 a_2346_15224# a_26970_15182# 0.35fF
C13856 a_1962_4178# col_n[8] 0.13fF
C13857 a_1962_17230# col_n[10] 0.13fF
C13858 a_17022_15182# vcm 0.62fF
C13859 a_20034_8154# VDD 0.52fF
C13860 a_2346_7192# a_2874_7150# 0.35fF
C13861 a_30074_12170# col[27] 0.29fF
C13862 a_1962_11206# col[1] 0.11fF
C13863 a_1962_12210# a_21038_12170# 0.27fF
C13864 m2_12776_946# m3_11904_1078# 0.13fF
C13865 a_10298_9198# vcm 0.22fF
C13866 col[0] rowoff_n[12] 0.11fF
C13867 a_3970_3134# m2_4168_3382# 0.16fF
C13868 a_7894_5142# rowoff_n[3] 0.24fF
C13869 a_2346_10204# col[21] 0.15fF
C13870 a_19030_9158# row_n[7] 0.17fF
C13871 a_33086_12170# VDD 0.52fF
C13872 m3_33992_18146# m3_34996_18146# 0.22fF
C13873 m2_23820_946# m3_23952_1078# 2.79fF
C13874 a_2346_9200# a_16018_9158# 0.19fF
C13875 a_26058_10162# a_26058_9158# 1.00fF
C13876 a_1962_9198# a_14314_9198# 0.14fF
C13877 m2_34864_16006# row_n[14] 0.15fF
C13878 a_1962_14218# a_34090_14178# 0.27fF
C13879 a_17934_3134# rowoff_n[1] 0.24fF
C13880 a_32994_14178# rowoff_n[12] 0.24fF
C13881 a_23350_13214# vcm 0.22fF
C13882 a_1962_6186# m2_34864_5966# 0.17fF
C13883 a_4974_7150# ctop 3.58fF
C13884 a_1962_6186# col[28] 0.11fF
C13885 a_13006_5142# col[10] 0.29fF
C13886 a_12914_15182# VDD 0.23fF
C13887 a_15926_11166# a_16018_11166# 0.26fF
C13888 a_2346_11208# a_29070_11166# 0.19fF
C13889 a_1962_11206# a_27366_11206# 0.14fF
C13890 m2_16792_946# a_17022_2130# 0.99fF
C13891 a_6982_7150# rowon_n[5] 0.14fF
C13892 a_30074_14178# col_n[27] 0.28fF
C13893 a_1962_13214# col_n[1] 0.13fF
C13894 a_2346_3176# a_5886_3134# 0.35fF
C13895 a_18026_11166# ctop 3.58fF
C13896 a_33086_17190# m2_33284_17438# 0.16fF
C13897 a_5978_11166# rowoff_n[9] 0.10fF
C13898 a_2346_6188# col[12] 0.15fF
C13899 a_9994_5142# a_10998_5142# 0.97fF
C13900 a_2346_5184# a_18938_5142# 0.35fF
C13901 a_31078_15182# ctop 3.58fF
C13902 a_26058_10162# rowon_n[8] 0.14fF
C13903 a_16018_9158# rowoff_n[7] 0.10fF
C13904 a_1962_8194# col_n[28] 0.13fF
C13905 a_13006_7150# col_n[10] 0.28fF
C13906 a_12002_15182# a_12002_14178# 1.00fF
C13907 a_28978_15182# a_29070_15182# 0.26fF
C13908 a_20034_15182# rowoff_n[13] 0.10fF
C13909 a_12002_14178# vcm 0.62fF
C13910 a_1962_2170# a_13006_2130# 0.27fF
C13911 a_1962_2170# col[19] 0.11fF
C13912 m2_30848_18014# m3_31984_18146# 0.13fF
C13913 a_15014_7150# VDD 0.52fF
C13914 a_1962_15222# col[21] 0.11fF
C13915 a_26058_7150# rowoff_n[5] 0.10fF
C13916 a_2346_7192# a_31990_7150# 0.35fF
C13917 a_31078_3134# col_n[28] 0.28fF
C13918 a_3970_10162# row_n[8] 0.17fF
C13919 a_5278_8194# vcm 0.22fF
C13920 a_28066_17190# col[25] 0.29fF
C13921 m2_23820_18014# col[21] 0.28fF
C13922 a_25054_18194# vcm 0.12fF
C13923 a_2346_18236# col[13] 0.14fF
C13924 a_1962_4178# a_26058_4138# 0.27fF
C13925 a_28066_11166# VDD 0.52fF
C13926 m3_23952_1078# m3_24956_1078# 0.22fF
C13927 rowon_n[0] ctop 1.17fF
C13928 col_n[28] col[28] 0.77fF
C13929 a_23046_9158# a_24050_9158# 0.97fF
C13930 a_35094_3134# vcm 0.12fF
C13931 col[27] rowoff_n[11] 0.11fF
C13932 a_18330_12210# vcm 0.22fF
C13933 a_2346_2172# col[3] 0.15fF
C13934 a_32082_6146# m2_32280_6394# 0.16fF
C13935 a_1962_1166# a_19334_1166# 0.19fF
C13936 a_2346_15224# col[5] 0.15fF
C13937 a_23046_13174# row_n[11] 0.17fF
C13938 a_7894_14178# VDD 0.23fF
C13939 a_1962_4178# col_n[19] 0.13fF
C13940 m2_13780_946# a_13918_1126# 0.16fF
C13941 a_1962_17230# col_n[21] 0.13fF
C13942 a_28066_17190# m3_27968_18146# 0.15fF
C13943 a_10998_10162# col[8] 0.29fF
C13944 a_31382_16226# vcm 0.22fF
C13945 a_7894_16186# rowoff_n[14] 0.24fF
C13946 a_2346_3176# a_34090_3134# 0.19fF
C13947 a_2966_8154# m2_3164_8402# 0.16fF
C13948 a_1962_3174# a_32386_3174# 0.14fF
C13949 a_1962_11206# col[12] 0.11fF
C13950 a_13006_10162# ctop 3.58fF
C13951 a_29070_6146# col[26] 0.29fF
C13952 m2_1732_9982# rowoff_n[8] 0.12fF
C13953 a_20946_18194# VDD 0.33fF
C13954 m2_16792_18014# vcm 0.28fF
C13955 col[11] rowoff_n[12] 0.11fF
C13956 a_1962_12210# a_2966_12170# 0.27fF
C13957 a_10998_11166# rowon_n[9] 0.14fF
C13958 a_35002_11166# rowoff_n[9] 0.24fF
C13959 a_30986_3134# VDD 0.23fF
C13960 m3_34996_3086# ctop 0.23fF
C13961 a_24962_5142# a_25054_5142# 0.26fF
C13962 a_7986_5142# a_7986_4138# 1.00fF
C13963 a_26058_14178# ctop 3.58fF
C13964 a_2346_14220# a_16930_14178# 0.35fF
C13965 a_8990_14178# a_9994_14178# 0.97fF
C13966 a_2346_18236# a_25966_18194# 0.35fF
C13967 a_6982_13174# vcm 0.62fF
C13968 a_10998_12170# col_n[8] 0.28fF
C13969 a_29070_7150# m2_29268_7398# 0.16fF
C13970 a_9994_6146# VDD 0.52fF
C13971 a_30074_14178# rowon_n[12] 0.14fF
C13972 a_1962_13214# col_n[12] 0.13fF
C13973 a_1962_11206# a_10998_11166# 0.27fF
C13974 a_29070_8154# col_n[26] 0.28fF
C13975 a_2346_16228# a_29982_16186# 0.35fF
C13976 a_2966_10162# col_n[0] 0.28fF
C13977 a_20034_17190# vcm 0.60fF
C13978 m2_7756_18014# VDD 1.08fF
C13979 a_1962_7190# col[3] 0.11fF
C13980 a_34090_10162# m2_34864_9982# 0.96fF
C13981 a_1962_18234# m2_22816_18014# 0.18fF
C13982 a_23046_10162# VDD 0.52fF
C13983 a_1962_8194# a_4274_8194# 0.14fF
C13984 a_21038_9158# a_21038_8154# 1.00fF
C13985 a_2346_8196# a_5978_8154# 0.19fF
C13986 a_7986_14178# row_n[12] 0.17fF
C13987 a_30074_2130# vcm 0.62fF
C13988 a_1962_13214# a_24050_13174# 0.27fF
C13989 m2_1732_9982# sample 0.19fF
C13990 a_2346_6188# col[23] 0.15fF
C13991 a_22042_12170# rowoff_n[10] 0.10fF
C13992 a_8990_4138# rowoff_n[2] 0.10fF
C13993 m2_34864_3958# ctop 0.17fF
C13994 a_23046_4138# row_n[2] 0.17fF
C13995 a_13310_11206# vcm 0.22fF
C13996 a_2346_18236# m2_17796_18014# 0.19fF
C13997 a_2346_13216# VDD 32.63fF
C13998 a_2346_10204# a_19030_10162# 0.19fF
C13999 a_1962_10202# a_17326_10202# 0.14fF
C14000 a_10906_10162# a_10998_10162# 0.26fF
C14001 a_19030_2130# rowoff_n[0] 0.10fF
C14002 m2_34864_9982# m2_35292_10410# 0.16fF
C14003 a_1962_2170# col[30] 0.11fF
C14004 a_26362_15222# vcm 0.22fF
C14005 a_8990_15182# col[6] 0.29fF
C14006 a_26058_8154# m2_26256_8402# 0.16fF
C14007 a_32082_3134# a_33086_3134# 0.97fF
C14008 m2_7756_18014# m3_6884_18146# 0.13fF
C14009 a_27062_17190# row_n[15] 0.17fF
C14010 a_7986_9158# ctop 3.58fF
C14011 a_1962_9198# col_n[3] 0.13fF
C14012 a_15926_17190# VDD 0.24fF
C14013 a_10998_2130# rowon_n[0] 0.14fF
C14014 a_1962_12210# a_30378_12210# 0.14fF
C14015 a_34090_13174# a_34090_12170# 1.00fF
C14016 a_2346_12212# a_32082_12170# 0.19fF
C14017 a_27062_11166# col[24] 0.29fF
C14018 a_2346_18236# col[24] 0.14fF
C14019 a_1962_3174# ctop 1.47fF
C14020 a_25966_2130# VDD 0.23fF
C14021 ctop col[1] 1.93fF
C14022 a_4974_4138# a_5978_4138# 0.97fF
C14023 a_2346_4180# a_8898_4138# 0.35fF
C14024 a_21038_13174# ctop 3.58fF
C14025 m3_34996_8106# m3_34996_7102# 0.22fF
C14026 a_23958_14178# a_24050_14178# 0.26fF
C14027 a_6982_14178# a_6982_13174# 1.00fF
C14028 a_7894_10162# rowoff_n[8] 0.24fF
C14029 a_2346_2172# col[14] 0.15fF
C14030 a_15014_15182# rowon_n[13] 0.14fF
C14031 a_2346_15224# col[16] 0.15fF
C14032 a_34394_13214# vcm 0.22fF
C14033 a_9902_13174# rowoff_n[11] 0.24fF
C14034 m2_2736_1950# VDD 0.57fF
C14035 a_4974_5142# VDD 0.52fF
C14036 a_30074_5142# rowon_n[3] 0.14fF
C14037 a_1962_4178# col_n[30] 0.13fF
C14038 a_1962_13214# m2_1732_12994# 0.15fF
C14039 a_2346_6188# a_21950_6146# 0.35fF
C14040 a_1962_17230# rowon_n[15] 1.18fF
C14041 a_8990_17190# col_n[6] 0.28fF
C14042 a_34090_17190# ctop 3.24fF
C14043 a_17934_8154# rowoff_n[6] 0.24fF
C14044 a_9994_4138# col[7] 0.29fF
C14045 a_1962_18234# col[6] 0.11fF
C14046 a_1962_11206# col[23] 0.11fF
C14047 a_3970_1126# m2_4168_1374# 0.16fF
C14048 a_1962_1166# m2_6752_946# 0.18fF
C14049 a_15014_16186# vcm 0.62fF
C14050 a_23958_17190# rowoff_n[15] 0.24fF
C14051 a_7986_5142# row_n[3] 0.17fF
C14052 a_27974_6146# rowoff_n[4] 0.24fF
C14053 a_23046_9158# m2_23244_9406# 0.16fF
C14054 a_27062_13174# col_n[24] 0.28fF
C14055 a_1962_3174# a_16018_3134# 0.27fF
C14056 a_18026_9158# VDD 0.52fF
C14057 col[22] rowoff_n[12] 0.11fF
C14058 a_2346_8196# a_35002_8154# 0.35fF
C14059 a_18026_8154# a_19030_8154# 0.97fF
C14060 m2_14784_946# ctop 0.18fF
C14061 a_25054_1126# vcm 0.12fF
C14062 a_8290_10202# vcm 0.22fF
C14063 a_2346_17232# a_3970_17190# 0.19fF
C14064 m2_31852_946# ctop 0.19fF
C14065 a_1962_5182# a_29070_5142# 0.27fF
C14066 a_31078_13174# VDD 0.52fF
C14067 a_2346_11208# col[7] 0.15fF
C14068 a_27062_8154# row_n[6] 0.17fF
C14069 a_21342_14218# vcm 0.22fF
C14070 a_9994_6146# col_n[7] 0.28fF
C14071 a_30074_3134# a_30074_2130# 1.00fF
C14072 a_1962_2170# a_22346_2170# 0.14fF
C14073 a_2346_2172# a_24050_2130# 0.19fF
C14074 col[6] rowoff_n[13] 0.11fF
C14075 a_1962_13214# col_n[23] 0.13fF
C14076 a_10906_16186# VDD 0.23fF
C14077 a_31078_12170# a_32082_12170# 0.97fF
C14078 a_28066_2130# col_n[25] 0.29fF
C14079 a_1962_7190# col[14] 0.11fF
C14080 a_2346_12212# row_n[10] 0.35fF
C14081 a_35398_18234# vcm 0.22fF
C14082 a_20946_1126# VDD 0.44fF
C14083 a_25054_16186# col[22] 0.29fF
C14084 a_19942_4138# a_20034_4138# 0.26fF
C14085 a_20034_10162# m2_20232_10410# 0.16fF
C14086 a_16018_12170# ctop 3.58fF
C14087 a_15014_6146# rowon_n[4] 0.14fF
C14088 a_2346_13216# a_6890_13174# 0.35fF
C14089 a_3970_13174# a_4974_13174# 0.97fF
C14090 a_1962_8194# rowon_n[6] 1.18fF
C14091 a_33998_5142# VDD 0.23fF
C14092 m3_33992_18146# VDD 0.26fF
C14093 a_29070_16186# ctop 3.57fF
C14094 a_2346_15224# a_19942_15182# 0.35fF
C14095 a_7986_9158# col[5] 0.29fF
C14096 a_9994_15182# vcm 0.62fF
C14097 a_1962_9198# col_n[14] 0.13fF
C14098 a_34090_9158# rowon_n[7] 0.14fF
C14099 a_13006_8154# VDD 0.52fF
C14100 a_32994_8154# a_33086_8154# 0.26fF
C14101 a_16018_8154# a_16018_7150# 1.00fF
C14102 a_1962_12210# a_14010_12170# 0.27fF
C14103 a_26058_5142# col[23] 0.29fF
C14104 a_1962_3174# col[5] 0.11fF
C14105 a_3270_9198# vcm 0.22fF
C14106 a_17022_17190# a_18026_17190# 0.97fF
C14107 a_2346_17232# a_32994_17190# 0.35fF
C14108 ctop col[12] 1.98fF
C14109 a_1962_16226# col[7] 0.11fF
C14110 m2_7756_946# m3_7888_1078# 2.79fF
C14111 a_12002_9158# row_n[7] 0.17fF
C14112 a_17022_11166# m2_17220_11414# 0.16fF
C14113 a_2966_13174# ctop 3.42fF
C14114 a_26058_12170# VDD 0.52fF
C14115 m3_19936_18146# m3_20940_18146# 0.22fF
C14116 a_1962_9198# a_7286_9198# 0.14fF
C14117 a_5886_9158# a_5978_9158# 0.26fF
C14118 a_2346_9200# a_8990_9158# 0.19fF
C14119 a_2346_2172# col[25] 0.15fF
C14120 a_2346_15224# col[27] 0.15fF
C14121 a_33086_4138# vcm 0.62fF
C14122 a_1962_14218# a_27062_14178# 0.27fF
C14123 a_10906_3134# rowoff_n[1] 0.24fF
C14124 a_25966_14178# rowoff_n[12] 0.24fF
C14125 a_16322_13214# vcm 0.22fF
C14126 a_27062_2130# a_28066_2130# 0.97fF
C14127 a_2346_6188# a_3878_6146# 0.35fF
C14128 a_7986_11166# col_n[5] 0.28fF
C14129 a_2874_6146# a_2966_6146# 0.26fF
C14130 a_5886_15182# VDD 0.23fF
C14131 a_1962_18234# col[17] 0.11fF
C14132 a_29070_12170# a_29070_11166# 1.00fF
C14133 a_1962_11206# a_20338_11206# 0.14fF
C14134 a_2346_11208# a_22042_11166# 0.19fF
C14135 a_2346_3176# row_n[1] 0.35fF
C14136 a_24050_2130# m2_24248_2378# 0.16fF
C14137 a_31078_12170# row_n[10] 0.17fF
C14138 a_29374_17230# vcm 0.22fF
C14139 a_26058_7150# col_n[23] 0.28fF
C14140 a_1962_5182# col_n[5] 0.13fF
C14141 a_10998_11166# ctop 3.58fF
C14142 a_1962_13214# a_33390_13214# 0.14fF
C14143 a_18938_13174# a_19030_13174# 0.26fF
C14144 a_28978_4138# VDD 0.23fF
C14145 a_2346_5184# a_11910_5142# 0.35fF
C14146 a_14010_12170# m2_14208_12418# 0.16fF
C14147 a_24050_15182# ctop 3.58fF
C14148 a_2346_11208# col[18] 0.15fF
C14149 a_19030_10162# rowon_n[8] 0.14fF
C14150 a_8990_9158# rowoff_n[7] 0.10fF
C14151 col[17] rowoff_n[13] 0.11fF
C14152 a_13006_15182# rowoff_n[13] 0.10fF
C14153 a_4974_14178# vcm 0.62fF
C14154 m2_34864_9982# VDD 1.03fF
C14155 a_35002_8154# m2_34864_7974# 0.16fF
C14156 a_1962_2170# a_5978_2130# 0.27fF
C14157 sample_n rowoff_n[6] 0.38fF
C14158 vcm rowoff_n[9] 0.20fF
C14159 m2_21812_18014# m3_21944_18146# 2.78fF
C14160 VDD rowoff_n[5] 1.17fF
C14161 a_7986_7150# VDD 0.52fF
C14162 a_19030_7150# rowoff_n[5] 0.10fF
C14163 a_5978_14178# col[3] 0.29fF
C14164 a_13006_7150# a_14010_7150# 0.97fF
C14165 a_2346_7192# a_24962_7150# 0.35fF
C14166 a_1962_7190# col[25] 0.11fF
C14167 a_31990_17190# a_32082_17190# 0.26fF
C14168 a_15014_17190# a_15014_16186# 1.00fF
C14169 a_29070_5142# rowoff_n[3] 0.10fF
C14170 a_18026_18194# vcm 0.12fF
C14171 a_24050_10162# col[21] 0.29fF
C14172 a_1962_1166# VDD 27.52fF
C14173 a_1962_4178# a_19030_4138# 0.27fF
C14174 a_1962_14218# sample 0.14fF
C14175 a_21038_11166# VDD 0.52fF
C14176 m3_9896_1078# m3_10900_1078# 0.22fF
C14177 a_2966_9158# a_2966_8154# 1.00fF
C14178 a_28066_3134# vcm 0.62fF
C14179 col[1] rowoff_n[14] 0.11fF
C14180 m2_1732_6970# ctop 0.17fF
C14181 a_11302_12210# vcm 0.22fF
C14182 a_1962_1166# a_12306_1166# 0.14fF
C14183 a_16018_13174# row_n[11] 0.17fF
C14184 a_1962_6186# a_32082_6146# 0.27fF
C14185 a_10998_13174# m2_11196_13422# 0.16fF
C14186 a_2346_7192# col[9] 0.15fF
C14187 a_34090_15182# VDD 0.54fF
C14188 a_26058_11166# a_27062_11166# 0.97fF
C14189 a_31078_3134# row_n[1] 0.17fF
C14190 a_5978_16186# col_n[3] 0.28fF
C14191 a_6982_3134# col[4] 0.29fF
C14192 a_1962_9198# col_n[25] 0.13fF
C14193 a_24354_16226# vcm 0.22fF
C14194 a_1962_3174# a_25358_3174# 0.14fF
C14195 a_2346_3176# a_27062_3134# 0.19fF
C14196 a_14922_3134# a_15014_3134# 0.26fF
C14197 a_17022_2130# m3_16924_1078# 0.15fF
C14198 a_5978_10162# ctop 3.58fF
C14199 a_24050_12170# col_n[21] 0.28fF
C14200 a_1962_3174# col[16] 0.11fF
C14201 a_13918_18194# VDD 0.33fF
C14202 VDD col_n[1] 4.67fF
C14203 sample_n vcm 1.11fF
C14204 m2_2736_18014# vcm 0.27fF
C14205 col[8] col[9] 0.20fF
C14206 a_1962_16226# col[18] 0.11fF
C14207 ctop col[23] 1.98fF
C14208 a_3970_11166# rowon_n[9] 0.14fF
C14209 a_27974_11166# rowoff_n[9] 0.24fF
C14210 a_23958_3134# VDD 0.23fF
C14211 m3_34996_17142# ctop 0.23fF
C14212 a_2966_11166# m2_1732_10986# 0.96fF
C14213 a_19030_14178# ctop 3.58fF
C14214 m2_26832_946# m2_27836_946# 0.96fF
C14215 a_2346_14220# a_9902_14178# 0.35fF
C14216 m2_20808_946# col[18] 0.39fF
C14217 a_2346_18236# a_18938_18194# 0.35fF
C14218 a_2874_6146# VDD 0.24fF
C14219 a_1962_18234# col[28] 0.11fF
C14220 a_6982_5142# col_n[4] 0.28fF
C14221 a_27974_7150# a_28066_7150# 0.26fF
C14222 a_7986_14178# m2_8184_14426# 0.16fF
C14223 a_10998_7150# a_10998_6146# 1.00fF
C14224 a_2346_3176# col[0] 0.15fF
C14225 a_2346_16228# col[2] 0.15fF
C14226 a_1962_11206# a_3970_11166# 0.27fF
C14227 a_23046_14178# rowon_n[12] 0.14fF
C14228 a_12002_16186# a_13006_16186# 0.97fF
C14229 a_2346_16228# a_22954_16186# 0.35fF
C14230 a_1962_5182# col_n[16] 0.13fF
C14231 a_13006_17190# vcm 0.60fF
C14232 a_1962_18234# m2_8760_18014# 0.18fF
C14233 a_16018_10162# VDD 0.52fF
C14234 a_22042_15182# col[19] 0.29fF
C14235 a_1962_12210# col[9] 0.11fF
C14236 a_23046_2130# vcm 0.62fF
C14237 a_1962_13214# a_17022_13174# 0.27fF
C14238 a_16018_4138# row_n[2] 0.17fF
C14239 a_15014_12170# rowoff_n[10] 0.10fF
C14240 a_6282_11206# vcm 0.22fF
C14241 a_2346_11208# col[29] 0.15fF
C14242 m3_9896_1078# VDD 0.14fF
C14243 a_29070_14178# VDD 0.52fF
C14244 a_2346_18236# m2_3740_18014# 0.19fF
C14245 a_1962_10202# a_10298_10202# 0.14fF
C14246 a_24050_11166# a_24050_10162# 1.00fF
C14247 a_2346_10204# a_12002_10162# 0.19fF
C14248 a_12002_2130# rowoff_n[0] 0.10fF
C14249 col[28] rowoff_n[13] 0.11fF
C14250 a_2346_5184# vcm 0.40fF
C14251 a_1962_15222# a_30074_15182# 0.27fF
C14252 a_19334_15222# vcm 0.22fF
C14253 a_29070_16186# rowoff_n[14] 0.10fF
C14254 m2_30848_18014# ctop 0.18fF
C14255 a_20034_17190# row_n[15] 0.17fF
C14256 a_4974_8154# col[2] 0.29fF
C14257 a_4974_15182# m2_5172_15430# 0.16fF
C14258 m2_34864_6970# row_n[5] 0.15fF
C14259 a_3970_2130# rowon_n[0] 0.14fF
C14260 a_8898_17190# VDD 0.24fF
C14261 a_2346_12212# a_25054_12170# 0.19fF
C14262 a_1962_12210# a_23350_12210# 0.14fF
C14263 a_13918_12170# a_14010_12170# 0.26fF
C14264 a_22042_17190# col_n[19] 0.28fF
C14265 a_1962_1166# col_n[7] 0.13fF
C14266 a_1962_14218# col_n[9] 0.13fF
C14267 a_6982_3134# m2_7180_3382# 0.16fF
C14268 a_23046_4138# col[20] 0.29fF
C14269 a_18938_2130# VDD 0.23fF
C14270 a_14010_13174# ctop 3.58fF
C14271 a_2966_11166# VDD 0.56fF
C14272 m2_28840_946# m3_28972_1078# 2.79fF
C14273 m3_34996_15134# m3_34996_14130# 0.22fF
C14274 a_1962_8194# col[0] 0.11fF
C14275 col[12] rowoff_n[14] 0.11fF
C14276 a_7986_15182# rowon_n[13] 0.14fF
C14277 a_2346_13216# rowoff_n[11] 4.09fF
C14278 a_2346_7192# col[20] 0.15fF
C14279 a_31990_6146# VDD 0.23fF
C14280 a_23046_5142# rowon_n[3] 0.14fF
C14281 a_2346_6188# a_14922_6146# 0.35fF
C14282 a_7986_6146# a_8990_6146# 0.97fF
C14283 a_27062_17190# ctop 3.39fF
C14284 a_10906_8154# rowoff_n[6] 0.24fF
C14285 a_4974_10162# col_n[2] 0.28fF
C14286 a_9994_16186# a_9994_15182# 1.00fF
C14287 a_26970_16186# a_27062_16186# 0.26fF
C14288 a_7986_16186# vcm 0.62fF
C14289 a_16930_17190# rowoff_n[15] 0.24fF
C14290 a_20946_6146# rowoff_n[4] 0.24fF
C14291 a_1962_3174# a_8990_3134# 0.27fF
C14292 a_1962_3174# col[27] 0.11fF
C14293 vcm col_n[8] 2.80fF
C14294 VDD col_n[12] 4.98fF
C14295 a_10998_9158# VDD 0.52fF
C14296 a_1962_16226# col[29] 0.11fF
C14297 a_2346_8196# a_27974_8154# 0.35fF
C14298 a_23046_6146# col_n[20] 0.28fF
C14299 a_18026_1126# vcm 0.59fF
C14300 a_1962_10202# vcm 6.95fF
C14301 a_30986_4138# rowoff_n[2] 0.24fF
C14302 m2_7756_946# ctop 0.18fF
C14303 a_3970_4138# m2_4168_4386# 0.16fF
C14304 a_1962_5182# a_22042_5142# 0.27fF
C14305 a_24050_13174# VDD 0.52fF
C14306 a_21038_10162# a_22042_10162# 0.97fF
C14307 a_31078_5142# vcm 0.62fF
C14308 a_20034_8154# row_n[6] 0.17fF
C14309 a_14314_14218# vcm 0.22fF
C14310 a_9902_2130# a_9994_2130# 0.26fF
C14311 a_2346_2172# a_17022_2130# 0.19fF
C14312 a_1962_2170# a_15318_2170# 0.14fF
C14313 a_1962_7190# m2_34864_6970# 0.17fF
C14314 a_2346_3176# col[11] 0.15fF
C14315 a_2346_16228# col[13] 0.15fF
C14316 a_1962_5182# col_n[27] 0.13fF
C14317 a_2966_16186# a_3970_16186# 0.97fF
C14318 a_27366_18234# vcm 0.22fF
C14319 a_13918_1126# VDD 0.44fF
C14320 a_2346_4180# a_30074_4138# 0.19fF
C14321 a_1962_4178# a_28370_4178# 0.14fF
C14322 a_33086_5142# a_33086_4138# 1.00fF
C14323 a_1962_12210# col[20] 0.11fF
C14324 a_8990_12170# ctop 3.58fF
C14325 a_21038_9158# col[18] 0.29fF
C14326 a_10998_17190# m2_10768_18014# 1.00fF
C14327 a_7986_6146# rowon_n[4] 0.14fF
C14328 a_29070_10162# rowoff_n[8] 0.10fF
C14329 a_31078_13174# rowoff_n[11] 0.10fF
C14330 a_26970_5142# VDD 0.23fF
C14331 m3_5880_18146# VDD 0.24fF
C14332 a_22954_6146# a_23046_6146# 0.26fF
C14333 a_5978_6146# a_5978_5142# 1.00fF
C14334 a_22042_16186# ctop 3.57fF
C14335 a_31078_17190# m3_30980_18146# 0.15fF
C14336 a_2346_15224# a_12914_15182# 0.35fF
C14337 a_6982_15182# a_7986_15182# 0.97fF
C14338 m2_1732_1950# sample_n 0.15fF
C14339 m2_1732_12994# VDD 1.02fF
C14340 a_2346_12212# col[4] 0.15fF
C14341 a_3970_2130# col[1] 0.29fF
C14342 a_27062_9158# rowon_n[7] 0.14fF
C14343 a_5978_8154# VDD 0.52fF
C14344 a_1962_1166# col_n[18] 0.13fF
C14345 a_1962_18234# a_30378_18234# 0.14fF
C14346 a_1962_12210# a_6982_12170# 0.27fF
C14347 a_1962_14218# col_n[20] 0.13fF
C14348 a_21038_11166# col_n[18] 0.28fF
C14349 a_2346_17232# a_25966_17190# 0.35fF
C14350 m2_32856_18014# m2_33860_18014# 0.96fF
C14351 m3_12908_1078# ctop 0.23fF
C14352 a_4974_9158# row_n[7] 0.17fF
C14353 col[23] rowoff_n[14] 0.11fF
C14354 a_1962_8194# col[11] 0.11fF
C14355 a_2346_13216# rowon_n[11] 0.26fF
C14356 a_19030_12170# VDD 0.52fF
C14357 m3_5880_18146# m3_6884_18146# 0.22fF
C14358 a_19030_10162# a_19030_9158# 1.00fF
C14359 m2_17796_18014# col[15] 0.28fF
C14360 a_26058_4138# vcm 0.62fF
C14361 a_1962_14218# a_20034_14178# 0.27fF
C14362 a_2346_7192# col[31] 0.15fF
C14363 a_18938_14178# rowoff_n[12] 0.24fF
C14364 a_9294_13214# vcm 0.22fF
C14365 a_32082_7150# m2_32280_7398# 0.16fF
C14366 a_32082_16186# VDD 0.52fF
C14367 a_2346_11208# a_15014_11166# 0.19fF
C14368 a_1962_11206# a_13310_11206# 0.14fF
C14369 a_8898_11166# a_8990_11166# 0.26fF
C14370 a_3970_4138# col_n[1] 0.28fF
C14371 a_1962_16226# a_33086_16186# 0.27fF
C14372 a_24050_12170# row_n[10] 0.17fF
C14373 m2_1732_12994# m2_2160_13422# 0.16fF
C14374 a_9994_2130# m2_9764_946# 0.99fF
C14375 col_n[9] col_n[10] 0.10fF
C14376 VDD col_n[23] 4.95fF
C14377 a_22346_17230# vcm 0.22fF
C14378 vcm col_n[19] 2.80fF
C14379 col[7] rowoff_n[15] 0.11fF
C14380 col[19] col[20] 0.20fF
C14381 a_2966_9158# m2_3164_9406# 0.16fF
C14382 a_30074_4138# a_31078_4138# 0.97fF
C14383 a_3970_11166# ctop 3.57fF
C14384 a_30074_17190# m2_29844_18014# 1.00fF
C14385 m2_7756_946# col[5] 0.39fF
C14386 a_1962_10202# col_n[11] 0.13fF
C14387 a_32386_2170# vcm 0.22fF
C14388 a_1962_13214# a_26362_13214# 0.14fF
C14389 a_2346_13216# a_28066_13174# 0.19fF
C14390 a_32082_14178# a_32082_13174# 1.00fF
C14391 a_19030_14178# col[16] 0.29fF
C14392 m2_33860_18014# col_n[31] 0.25fF
C14393 a_21950_4138# VDD 0.23fF
C14394 a_1962_4178# col[2] 0.11fF
C14395 a_2346_5184# a_4882_5142# 0.35fF
C14396 a_1962_17230# col[4] 0.11fF
C14397 a_17022_15182# ctop 3.58fF
C14398 m2_34864_1950# vcm 0.51fF
C14399 a_12002_10162# rowon_n[8] 0.14fF
C14400 a_21950_15182# a_22042_15182# 0.26fF
C14401 a_4974_15182# a_4974_14178# 1.00fF
C14402 a_2346_3176# col[22] 0.15fF
C14403 a_2346_16228# col[24] 0.15fF
C14404 a_5978_15182# rowoff_n[13] 0.10fF
C14405 a_29070_8154# m2_29268_8402# 0.16fF
C14406 m2_12776_18014# m3_11904_18146# 0.13fF
C14407 a_35002_8154# VDD 0.29fF
C14408 a_12002_7150# rowoff_n[5] 0.10fF
C14409 a_2346_7192# a_17934_7150# 0.35fF
C14410 a_1962_12210# a_34394_12210# 0.14fF
C14411 m2_34864_17010# m2_34864_16006# 0.99fF
C14412 a_22042_5142# rowoff_n[3] 0.10fF
C14413 a_2346_4180# rowon_n[2] 0.26fF
C14414 a_1962_12210# col[31] 0.11fF
C14415 a_10998_18194# vcm 0.12fF
C14416 a_19030_16186# col_n[16] 0.28fF
C14417 a_34090_11166# m2_34864_10986# 0.96fF
C14418 a_1962_4178# a_12002_4138# 0.27fF
C14419 a_31078_13174# rowon_n[11] 0.14fF
C14420 a_14010_11166# VDD 0.52fF
C14421 a_20034_3134# col[17] 0.29fF
C14422 a_2346_9200# a_30986_9158# 0.35fF
C14423 a_16018_9158# a_17022_9158# 0.97fF
C14424 a_1962_6186# col_n[2] 0.13fF
C14425 a_21038_3134# vcm 0.62fF
C14426 a_32082_3134# rowoff_n[1] 0.10fF
C14427 a_4274_12210# vcm 0.22fF
C14428 a_1962_1166# a_5278_1166# 0.14fF
C14429 a_8990_13174# row_n[11] 0.17fF
C14430 a_1962_6186# a_25054_6146# 0.27fF
C14431 a_27062_15182# VDD 0.52fF
C14432 a_24050_3134# row_n[1] 0.17fF
C14433 a_34090_7150# vcm 0.62fF
C14434 a_2346_12212# col[15] 0.15fF
C14435 a_6890_1126# m2_6752_946# 0.16fF
C14436 a_17326_16226# vcm 0.22fF
C14437 a_28066_4138# a_28066_3134# 1.00fF
C14438 a_26058_9158# m2_26256_9406# 0.16fF
C14439 a_1962_3174# a_18330_3174# 0.14fF
C14440 a_2346_3176# a_20034_3134# 0.19fF
C14441 a_2346_1168# m2_24824_946# 0.19fF
C14442 a_1962_1166# col_n[29] 0.13fF
C14443 a_1962_14218# col_n[31] 0.13fF
C14444 a_6890_18194# VDD 0.34fF
C14445 a_27366_1166# vcm 0.23fF
C14446 a_29070_13174# a_30074_13174# 0.97fF
C14447 m2_9764_946# m2_10768_946# 0.96fF
C14448 a_20034_5142# col_n[17] 0.28fF
C14449 a_20946_11166# rowoff_n[9] 0.24fF
C14450 a_28066_16186# row_n[14] 0.17fF
C14451 a_1962_8194# col[22] 0.11fF
C14452 a_16930_3134# VDD 0.23fF
C14453 m3_8892_18146# ctop 0.23fF
C14454 a_1962_5182# a_31382_5182# 0.14fF
C14455 a_17934_5142# a_18026_5142# 0.26fF
C14456 a_2346_5184# a_33086_5142# 0.19fF
C14457 a_12002_14178# ctop 3.58fF
C14458 a_30986_9158# rowoff_n[7] 0.24fF
C14459 a_2346_18236# a_11910_18194# 0.35fF
C14460 a_35002_15182# rowoff_n[13] 0.24fF
C14461 m2_34864_8978# rowon_n[7] 0.13fF
C14462 a_29982_7150# VDD 0.23fF
C14463 a_1962_14218# m2_1732_13998# 0.15fF
C14464 a_16018_14178# rowon_n[12] 0.14fF
C14465 VDD rowon_n[14] 2.61fF
C14466 vcm col_n[30] 2.80fF
C14467 a_2346_8196# col[6] 0.15fF
C14468 col[18] rowoff_n[15] 0.11fF
C14469 a_2346_16228# a_15926_16186# 0.35fF
C14470 a_31078_4138# rowon_n[2] 0.14fF
C14471 a_5978_17190# vcm 0.60fF
C14472 a_23046_10162# m2_23244_10410# 0.16fF
C14473 a_8990_10162# VDD 0.52fF
C14474 a_1962_10202# col_n[22] 0.13fF
C14475 a_30986_9158# a_31078_9158# 0.26fF
C14476 a_14010_9158# a_14010_8154# 1.00fF
C14477 a_16018_2130# vcm 0.62fF
C14478 a_1962_13214# a_9994_13174# 0.27fF
C14479 a_18026_8154# col[15] 0.29fF
C14480 a_7986_12170# rowoff_n[10] 0.10fF
C14481 a_8990_4138# row_n[2] 0.17fF
C14482 a_1962_4178# col[13] 0.11fF
C14483 a_1962_17230# col[15] 0.11fF
C14484 a_3878_4138# VDD 0.23fF
C14485 m3_34996_11118# VDD 0.26fF
C14486 a_22042_14178# VDD 0.52fF
C14487 m2_1732_2954# vcm 0.45fF
C14488 a_2346_10204# a_4974_10162# 0.19fF
C14489 a_1962_10202# a_3270_10202# 0.14fF
C14490 a_4974_2130# rowoff_n[0] 0.10fF
C14491 a_29070_6146# vcm 0.62fF
C14492 a_1962_15222# a_23046_15182# 0.27fF
C14493 a_12306_15222# vcm 0.22fF
C14494 m2_16792_18014# ctop 0.18fF
C14495 a_22042_16186# rowoff_n[14] 0.10fF
C14496 a_25054_3134# a_26058_3134# 0.97fF
C14497 a_13006_17190# row_n[15] 0.17fF
C14498 m2_1732_10986# row_n[9] 0.13fF
C14499 a_2346_12212# a_18026_12170# 0.19fF
C14500 a_27062_13174# a_27062_12170# 1.00fF
C14501 a_1962_12210# a_16322_12210# 0.14fF
C14502 a_28066_7150# row_n[5] 0.17fF
C14503 m2_34864_1950# m3_34996_1078# 0.15fF
C14504 a_11910_2130# VDD 0.23fF
C14505 a_18026_10162# col_n[15] 0.28fF
C14506 a_20034_11166# m2_20232_11414# 0.16fF
C14507 a_1962_6186# col_n[13] 0.13fF
C14508 a_6982_13174# ctop 3.58fF
C14509 a_9902_18194# m2_9764_18014# 0.16fF
C14510 a_2966_3134# vcm 0.61fF
C14511 a_16930_14178# a_17022_14178# 0.26fF
C14512 a_2346_14220# a_31078_14178# 0.19fF
C14513 a_1962_14218# a_29374_14218# 0.14fF
C14514 a_1962_13214# col[6] 0.11fF
C14515 rowon_n[9] rowoff_n[9] 20.27fF
C14516 a_24962_6146# VDD 0.23fF
C14517 a_16018_5142# rowon_n[3] 0.14fF
C14518 a_2346_6188# a_7894_6146# 0.35fF
C14519 a_20034_17190# ctop 3.39fF
C14520 a_2346_12212# col[26] 0.15fF
C14521 a_27062_2130# m2_27260_2378# 0.16fF
C14522 a_9902_17190# rowoff_n[15] 0.24fF
C14523 a_30074_2130# ctop 3.39fF
C14524 a_13918_6146# rowoff_n[4] 0.24fF
C14525 a_3970_9158# VDD 0.52fF
C14526 a_2346_8196# a_20946_8154# 0.35fF
C14527 a_10998_8154# a_12002_8154# 0.97fF
C14528 a_10998_1126# vcm 0.12fF
C14529 a_23958_4138# rowoff_n[2] 0.24fF
C14530 a_16018_13174# col[13] 0.29fF
C14531 m2_15788_946# vcm 0.42fF
C14532 a_1962_2170# col_n[4] 0.13fF
C14533 a_17022_12170# m2_17220_12418# 0.16fF
C14534 a_1962_5182# a_15014_5142# 0.27fF
C14535 a_1962_15222# col_n[6] 0.13fF
C14536 a_17022_13174# VDD 0.52fF
C14537 a_2346_10204# a_33998_10162# 0.35fF
C14538 a_33998_2130# rowoff_n[0] 0.24fF
C14539 a_24050_5142# vcm 0.62fF
C14540 m2_32856_946# vcm 0.41fF
C14541 a_34090_9158# col[31] 0.29fF
C14542 a_13006_8154# row_n[6] 0.17fF
C14543 a_7286_14218# vcm 0.22fF
C14544 a_1962_2170# a_8290_2170# 0.14fF
C14545 a_2346_2172# a_9994_2130# 0.19fF
C14546 a_23046_3134# a_23046_2130# 1.00fF
C14547 m2_26832_18014# m3_26964_18146# 2.78fF
C14548 a_2874_18194# VDD 0.34fF
C14549 a_1962_7190# a_28066_7150# 0.27fF
C14550 col_n[2] row_n[12] 0.23fF
C14551 vcm row_n[11] 0.49fF
C14552 VDD row_n[9] 2.93fF
C14553 col_n[8] row_n[15] 0.23fF
C14554 sample row_n[10] 1.03fF
C14555 col_n[4] row_n[13] 0.23fF
C14556 col_n[6] row_n[14] 0.23fF
C14557 col_n[20] col_n[21] 0.10fF
C14558 a_30074_17190# VDD 0.55fF
C14559 a_2346_8196# col[17] 0.15fF
C14560 col[30] col[31] 0.20fF
C14561 col[29] rowoff_n[15] 0.11fF
C14562 a_24050_12170# a_25054_12170# 0.97fF
C14563 a_20338_18234# vcm 0.22fF
C14564 a_6890_1126# VDD 0.44fF
C14565 a_12914_4138# a_13006_4138# 0.26fF
C14566 a_2346_4180# a_23046_4138# 0.19fF
C14567 a_1962_4178# a_21342_4178# 0.14fF
C14568 m2_2736_1950# rowon_n[0] 0.13fF
C14569 a_28978_18194# m2_28840_18014# 0.16fF
C14570 a_16018_15182# col_n[13] 0.28fF
C14571 a_1962_4178# col[24] 0.11fF
C14572 a_30378_3174# vcm 0.22fF
C14573 a_32082_11166# row_n[9] 0.17fF
C14574 a_17022_2130# col[14] 0.29fF
C14575 a_22042_10162# rowoff_n[8] 0.10fF
C14576 a_1962_17230# col[26] 0.11fF
C14577 a_24050_13174# rowoff_n[11] 0.10fF
C14578 a_19942_5142# VDD 0.23fF
C14579 a_14010_13174# m2_14208_13422# 0.16fF
C14580 a_1962_6186# a_35398_6186# 0.14fF
C14581 m2_23820_946# VDD 0.62fF
C14582 a_2346_6188# a_2346_5184# 0.22fF
C14583 a_34090_11166# col_n[31] 0.28fF
C14584 a_15014_16186# ctop 3.57fF
C14585 a_32082_8154# rowoff_n[6] 0.10fF
C14586 VDD rowoff_n[12] 1.17fF
C14587 a_2346_15224# a_5886_15182# 0.35fF
C14588 m2_13780_946# m2_14208_1374# 0.16fF
C14589 a_35002_9158# m2_34864_8978# 0.16fF
C14590 a_20034_2130# m3_19936_1078# 0.12fF
C14591 a_20034_9158# rowon_n[7] 0.14fF
C14592 a_32994_9158# VDD 0.23fF
C14593 a_25966_8154# a_26058_8154# 0.26fF
C14594 a_8990_8154# a_8990_7150# 1.00fF
C14595 a_2346_4180# col[8] 0.15fF
C14596 a_2346_17232# col[10] 0.15fF
C14597 a_1962_18234# a_23350_18234# 0.14fF
C14598 a_9994_17190# a_10998_17190# 0.97fF
C14599 a_2346_17232# a_18938_17190# 0.35fF
C14600 a_1962_6186# col_n[24] 0.13fF
C14601 m2_25828_18014# m2_26832_18014# 0.96fF
C14602 a_17022_4138# col_n[14] 0.28fF
C14603 m2_1732_1950# m3_2868_2082# 0.13fF
C14604 m3_1864_9110# ctop 0.23fF
C14605 a_12002_12170# VDD 0.52fF
C14606 m2_30848_946# m2_31276_1374# 0.16fF
C14607 a_1962_13214# col[17] 0.11fF
C14608 a_19030_4138# vcm 0.62fF
C14609 a_1962_14218# a_13006_14178# 0.27fF
C14610 a_11910_14178# rowoff_n[12] 0.24fF
C14611 a_20034_2130# a_21038_2130# 0.97fF
C14612 a_32082_14178# col[29] 0.29fF
C14613 a_10998_14178# m2_11196_14426# 0.16fF
C14614 a_25054_16186# VDD 0.52fF
C14615 m2_1732_12994# rowoff_n[11] 0.12fF
C14616 a_22042_12170# a_22042_11166# 1.00fF
C14617 a_2346_11208# a_7986_11166# 0.19fF
C14618 a_1962_11206# a_6282_11206# 0.14fF
C14619 a_32082_8154# vcm 0.62fF
C14620 a_1962_16226# a_26058_16186# 0.27fF
C14621 a_17022_12170# row_n[10] 0.17fF
C14622 a_15318_17230# vcm 0.22fF
C14623 m2_1046_19620# VDD 0.57fF
C14624 a_32082_2130# row_n[0] 0.17fF
C14625 a_2346_8196# a_1962_8194# 2.62fF
C14626 a_2346_13216# col[1] 0.15fF
C14627 a_25358_2170# vcm 0.22fF
C14628 a_1962_13214# a_19334_13214# 0.14fF
C14629 a_2346_13216# a_21038_13174# 0.19fF
C14630 a_11910_13174# a_12002_13174# 0.26fF
C14631 m2_1732_2954# m2_1732_1950# 0.99fF
C14632 a_1962_2170# col_n[15] 0.13fF
C14633 a_1962_15222# col_n[17] 0.13fF
C14634 a_15014_7150# col[12] 0.29fF
C14635 a_14922_4138# VDD 0.23fF
C14636 m3_24956_1078# VDD 0.14fF
C14637 m2_30848_946# col[28] 0.39fF
C14638 a_2966_12170# m2_1732_11990# 0.96fF
C14639 a_33086_6146# a_34090_6146# 0.97fF
C14640 a_9994_15182# ctop 3.58fF
C14641 a_4974_10162# rowon_n[8] 0.14fF
C14642 a_1962_9198# col[8] 0.11fF
C14643 a_32082_16186# col_n[29] 0.28fF
C14644 a_2346_15224# a_34090_15182# 0.19fF
C14645 a_1962_15222# a_32386_15222# 0.14fF
C14646 a_33086_3134# col[30] 0.29fF
C14647 m2_2736_18014# m3_3872_18146# 0.13fF
C14648 col_n[5] row_n[8] 0.23fF
C14649 col_n[7] row_n[9] 0.23fF
C14650 col_n[9] row_n[10] 0.23fF
C14651 col_n[0] row_n[5] 0.23fF
C14652 col_n[17] row_n[14] 0.23fF
C14653 col_n[15] row_n[13] 0.23fF
C14654 col_n[11] row_n[11] 0.23fF
C14655 vcm rowon_n[5] 0.50fF
C14656 VDD rowon_n[3] 2.61fF
C14657 col_n[3] row_n[7] 0.23fF
C14658 col_n[13] row_n[12] 0.23fF
C14659 col_n[19] row_n[15] 0.23fF
C14660 col_n[1] row_n[6] 0.23fF
C14661 a_2346_8196# col[28] 0.15fF
C14662 a_27974_8154# VDD 0.23fF
C14663 a_4974_7150# rowoff_n[5] 0.10fF
C14664 a_7986_15182# m2_8184_15430# 0.16fF
C14665 a_5978_7150# a_6982_7150# 0.97fF
C14666 a_2346_7192# a_10906_7150# 0.35fF
C14667 a_7986_17190# a_7986_16186# 1.00fF
C14668 a_24962_17190# a_25054_17190# 0.26fF
C14669 a_9994_3134# m2_10192_3382# 0.16fF
C14670 a_15014_5142# rowoff_n[3] 0.10fF
C14671 a_33086_4138# ctop 3.57fF
C14672 a_1962_4178# a_4974_4138# 0.27fF
C14673 a_3878_4138# a_3970_4138# 0.26fF
C14674 a_24050_13174# rowon_n[11] 0.14fF
C14675 a_6982_11166# VDD 0.52fF
C14676 m2_33860_946# m3_33992_1078# 0.84fF
C14677 a_15014_9158# col_n[12] 0.28fF
C14678 a_2346_9200# a_23958_9158# 0.35fF
C14679 a_14010_3134# vcm 0.62fF
C14680 a_25054_3134# rowoff_n[1] 0.10fF
C14681 a_1962_11206# col_n[8] 0.13fF
C14682 a_18026_2130# a_18026_1126# 1.00fF
C14683 a_35494_6508# VDD 0.11fF
C14684 a_33086_5142# col_n[30] 0.28fF
C14685 a_1962_6186# a_18026_6146# 0.27fF
C14686 a_20034_15182# VDD 0.52fF
C14687 a_19030_11166# a_20034_11166# 0.97fF
C14688 a_1962_11206# a_1962_10202# 0.16fF
C14689 a_17022_3134# row_n[1] 0.17fF
C14690 a_27062_7150# vcm 0.62fF
C14691 a_10298_16226# vcm 0.22fF
C14692 a_2346_3176# a_13006_3134# 0.19fF
C14693 a_7894_3134# a_7986_3134# 0.26fF
C14694 a_1962_3174# a_11302_3174# 0.14fF
C14695 a_2346_4180# col[19] 0.15fF
C14696 a_2346_17232# col[21] 0.15fF
C14697 a_4974_16186# m2_5172_16434# 0.16fF
C14698 a_1962_8194# a_31078_8154# 0.27fF
C14699 a_20338_1166# vcm 0.22fF
C14700 a_13918_11166# rowoff_n[9] 0.24fF
C14701 a_21038_16186# row_n[14] 0.17fF
C14702 a_6982_4138# m2_7180_4386# 0.16fF
C14703 a_9902_3134# VDD 0.23fF
C14704 a_31078_6146# a_31078_5142# 1.00fF
C14705 a_2346_5184# a_26058_5142# 0.19fF
C14706 a_1962_5182# a_24354_5182# 0.14fF
C14707 a_4974_14178# ctop 3.58fF
C14708 a_1962_13214# col[28] 0.11fF
C14709 a_13006_12170# col[10] 0.29fF
C14710 a_23958_9158# rowoff_n[7] 0.24fF
C14711 ctop rowoff_n[9] 0.60fF
C14712 a_33390_5182# vcm 0.22fF
C14713 a_32082_15182# a_33086_15182# 0.97fF
C14714 a_2346_18236# a_4882_18194# 0.35fF
C14715 a_1962_7190# col_n[0] 0.13fF
C14716 m2_1732_12994# rowon_n[11] 0.11fF
C14717 a_27974_15182# rowoff_n[13] 0.24fF
C14718 a_31078_8154# col[28] 0.29fF
C14719 a_22954_7150# VDD 0.23fF
C14720 a_33998_7150# rowoff_n[5] 0.24fF
C14721 a_20946_7150# a_21038_7150# 0.26fF
C14722 a_3970_7150# a_3970_6146# 1.00fF
C14723 a_8990_14178# rowon_n[12] 0.14fF
C14724 a_2346_16228# a_8898_16186# 0.35fF
C14725 a_4974_16186# a_5978_16186# 0.97fF
C14726 a_24050_4138# rowon_n[2] 0.14fF
C14727 a_28066_3134# ctop 3.57fF
C14728 a_2346_13216# col[12] 0.15fF
C14729 a_1962_2170# col_n[26] 0.13fF
C14730 a_8990_2130# vcm 0.62fF
C14731 a_2346_13216# a_2966_13174# 0.21fF
C14732 a_1962_15222# col_n[28] 0.13fF
C14733 a_13006_14178# col_n[10] 0.28fF
C14734 a_2346_1168# a_28978_1126# 0.35fF
C14735 a_3970_5142# m2_4168_5390# 0.16fF
C14736 m3_20940_18146# VDD 0.24fF
C14737 a_1962_9198# col[19] 0.11fF
C14738 a_28066_17190# rowon_n[15] 0.14fF
C14739 a_15014_14178# VDD 0.52fF
C14740 a_33998_11166# a_34090_11166# 0.26fF
C14741 a_17022_11166# a_17022_10162# 1.00fF
C14742 a_31078_10162# col_n[28] 0.28fF
C14743 a_34090_17190# m3_33992_18146# 0.15fF
C14744 a_22042_6146# vcm 0.62fF
C14745 a_1962_15222# a_16018_15182# 0.27fF
C14746 VDD en_C0_n 0.15fF
C14747 col_n[6] row_n[3] 0.23fF
C14748 col_n[28] row_n[14] 0.23fF
C14749 col_n[26] row_n[13] 0.23fF
C14750 col_n[2] row_n[1] 0.23fF
C14751 col_n[16] row_n[8] 0.23fF
C14752 col_n[8] row_n[4] 0.23fF
C14753 col_n[10] row_n[5] 0.23fF
C14754 col_n[20] row_n[10] 0.23fF
C14755 col_n[24] row_n[12] 0.23fF
C14756 col_n[4] row_n[2] 0.23fF
C14757 col_n[12] row_n[6] 0.23fF
C14758 col_n[14] row_n[7] 0.23fF
C14759 col_n[18] row_n[9] 0.23fF
C14760 col_n[30] row_n[15] 0.23fF
C14761 vcm row_n[0] 0.49fF
C14762 col_n[22] row_n[11] 0.23fF
C14763 a_5278_15222# vcm 0.22fF
C14764 a_15014_16186# rowoff_n[14] 0.10fF
C14765 m2_2736_18014# ctop 0.18fF
C14766 a_1962_8194# m2_34864_7974# 0.17fF
C14767 a_5978_17190# row_n[15] 0.17fF
C14768 m2_31852_18014# vcm 0.28fF
C14769 a_1962_12210# a_9294_12210# 0.14fF
C14770 a_1962_18234# a_34394_18234# 0.14fF
C14771 a_2346_12212# a_10998_12170# 0.19fF
C14772 a_6890_12170# a_6982_12170# 0.26fF
C14773 a_21038_7150# row_n[5] 0.17fF
C14774 a_35094_10162# vcm 0.12fF
C14775 a_1962_17230# a_29070_17190# 0.27fF
C14776 m2_2736_946# m3_3872_1078# 0.10fF
C14777 a_4882_2130# VDD 0.23fF
C14778 m3_27968_1078# ctop 0.23fF
C14779 a_2346_9200# col[3] 0.15fF
C14780 a_28066_5142# a_29070_5142# 0.97fF
C14781 a_14010_3134# col_n[11] 0.28fF
C14782 a_1962_18234# col_n[2] 0.13fF
C14783 a_28370_4178# vcm 0.22fF
C14784 a_1962_11206# col_n[19] 0.13fF
C14785 a_30074_15182# a_30074_14178# 1.00fF
C14786 a_1962_14218# a_22346_14218# 0.14fF
C14787 a_2346_14220# a_24050_14178# 0.19fF
C14788 a_10998_17190# col[8] 0.29fF
C14789 a_17934_6146# VDD 0.23fF
C14790 a_8990_5142# rowon_n[3] 0.14fF
C14791 a_1962_5182# col[10] 0.11fF
C14792 a_13006_17190# ctop 3.39fF
C14793 a_29070_13174# col[26] 0.29fF
C14794 a_19942_16186# a_20034_16186# 0.26fF
C14795 a_2346_4180# col[30] 0.15fF
C14796 a_23046_2130# ctop 3.39fF
C14797 a_2346_17232# rowoff_n[15] 4.09fF
C14798 m2_22816_18014# VDD 1.31fF
C14799 a_6890_6146# rowoff_n[4] 0.24fF
C14800 a_30986_10162# VDD 0.23fF
C14801 m2_33860_946# sw_n 0.57fF
C14802 a_2346_8196# a_13918_8154# 0.35fF
C14803 a_3970_1126# vcm 0.59fF
C14804 a_16930_4138# rowoff_n[2] 0.24fF
C14805 a_29982_12170# rowoff_n[10] 0.24fF
C14806 a_2966_16186# row_n[14] 0.16fF
C14807 a_28066_8154# rowon_n[6] 0.14fF
C14808 a_2346_5184# ctop 1.59fF
C14809 a_1962_5182# a_7986_5142# 0.27fF
C14810 col[0] rowoff_n[4] 0.11fF
C14811 col[2] rowoff_n[6] 0.11fF
C14812 col[1] rowoff_n[5] 0.11fF
C14813 col[5] rowoff_n[9] 0.11fF
C14814 col[3] rowoff_n[7] 0.11fF
C14815 col[4] rowoff_n[8] 0.11fF
C14816 a_2346_18236# m2_32856_18014# 0.19fF
C14817 a_12002_6146# col[9] 0.29fF
C14818 a_9994_13174# VDD 0.52fF
C14819 m2_8760_946# vcm 0.42fF
C14820 a_2346_10204# a_26970_10162# 0.35fF
C14821 a_14010_10162# a_15014_10162# 0.97fF
C14822 a_26970_2130# rowoff_n[0] 0.24fF
C14823 a_1962_7190# col_n[10] 0.13fF
C14824 a_17022_5142# vcm 0.62fF
C14825 a_5978_8154# row_n[6] 0.17fF
C14826 a_29070_15182# col_n[26] 0.28fF
C14827 a_2346_2172# a_2874_2130# 0.35fF
C14828 a_32082_8154# m2_32280_8402# 0.16fF
C14829 a_2966_17190# col_n[0] 0.28fF
C14830 m2_17796_18014# m3_16924_18146# 0.13fF
C14831 a_30074_2130# col[27] 0.29fF
C14832 a_1962_1166# col[1] 0.11fF
C14833 m2_11772_18014# col[9] 0.28fF
C14834 a_1962_14218# col[3] 0.11fF
C14835 a_1962_7190# a_21038_7150# 0.27fF
C14836 a_23046_17190# VDD 0.55fF
C14837 m2_34864_15002# vcm 0.51fF
C14838 a_30074_9158# vcm 0.62fF
C14839 a_2346_13216# col[23] 0.15fF
C14840 a_13310_18234# vcm 0.22fF
C14841 a_33086_2130# VDD 0.55fF
C14842 a_2966_10162# m2_3164_10410# 0.16fF
C14843 a_26058_5142# a_26058_4138# 1.00fF
C14844 a_2346_4180# a_16018_4138# 0.19fF
C14845 a_1962_4178# a_14314_4178# 0.14fF
C14846 a_1962_9198# a_34090_9158# 0.27fF
C14847 a_23350_3174# vcm 0.22fF
C14848 a_25054_11166# row_n[9] 0.17fF
C14849 a_27062_14178# a_28066_14178# 0.97fF
C14850 a_15014_10162# rowoff_n[8] 0.10fF
C14851 a_12002_8154# col_n[9] 0.28fF
C14852 a_17022_13174# rowoff_n[11] 0.10fF
C14853 a_1962_9198# col[30] 0.11fF
C14854 a_12914_5142# VDD 0.23fF
C14855 a_1962_6186# a_27366_6186# 0.14fF
C14856 a_15926_6146# a_16018_6146# 0.26fF
C14857 a_2346_6188# a_29070_6146# 0.19fF
C14858 a_7986_16186# ctop 3.57fF
C14859 a_25054_8154# rowoff_n[6] 0.10fF
C14860 a_30074_4138# col_n[27] 0.28fF
C14861 a_1962_3174# col_n[1] 0.13fF
C14862 m2_14784_946# a_1962_1166# 0.18fF
C14863 col_n[15] row_n[2] 0.23fF
C14864 vcm col[2] 5.84fF
C14865 col_n[11] row_n[0] 0.23fF
C14866 col_n[31] row_n[10] 0.23fF
C14867 col_n[27] row_n[8] 0.23fF
C14868 col_n[1] col[1] 0.64fF
C14869 col_n[29] row_n[9] 0.23fF
C14870 col_n[8] ctop 2.02fF
C14871 a_1962_16226# col_n[3] 0.13fF
C14872 rowon_n[13] rowon_n[12] 0.15fF
C14873 col_n[13] row_n[1] 0.23fF
C14874 col_n[19] row_n[4] 0.23fF
C14875 col_n[25] row_n[7] 0.23fF
C14876 VDD col[6] 4.17fF
C14877 col_n[21] row_n[5] 0.23fF
C14878 col_n[17] row_n[3] 0.23fF
C14879 col_n[23] row_n[6] 0.23fF
C14880 m2_27836_18014# col_n[25] 0.25fF
C14881 a_18026_1126# ctop 1.01fF
C14882 a_31078_17190# rowoff_n[15] 0.10fF
C14883 a_29070_9158# m2_29268_9406# 0.16fF
C14884 a_1962_1166# m2_31852_946# 0.18fF
C14885 a_1962_10202# ctop 1.49fF
C14886 a_13006_9158# rowon_n[7] 0.14fF
C14887 a_25966_9158# VDD 0.23fF
C14888 a_1962_18234# a_16322_18234# 0.14fF
C14889 a_2966_7150# row_n[5] 0.16fF
C14890 m2_1732_5966# sample 0.19fF
C14891 a_2346_17232# a_11910_17190# 0.35fF
C14892 a_2346_9200# col[14] 0.15fF
C14893 m2_1732_17010# sample_n 0.15fF
C14894 m2_18800_18014# m2_19804_18014# 0.96fF
C14895 a_31078_5142# ctop 3.58fF
C14896 m3_23952_18146# ctop 0.23fF
C14897 a_34090_12170# m2_34864_11990# 0.96fF
C14898 a_1962_18234# col_n[13] 0.13fF
C14899 a_4974_12170# VDD 0.52fF
C14900 a_1962_11206# col_n[30] 0.13fF
C14901 m2_23820_946# m2_24248_1374# 0.16fF
C14902 a_28978_10162# a_29070_10162# 0.26fF
C14903 a_12002_10162# a_12002_9158# 1.00fF
C14904 a_12002_4138# vcm 0.62fF
C14905 a_1962_14218# a_5978_14178# 0.27fF
C14906 a_9994_11166# col[7] 0.29fF
C14907 m2_34864_7974# m2_35292_8402# 0.16fF
C14908 a_4882_14178# rowoff_n[12] 0.24fF
C14909 a_1962_5182# col[21] 0.11fF
C14910 a_32082_12170# rowon_n[10] 0.14fF
C14911 a_2346_2172# a_31990_2130# 0.35fF
C14912 a_18026_16186# VDD 0.52fF
C14913 a_28066_7150# col[25] 0.29fF
C14914 a_25054_8154# vcm 0.62fF
C14915 a_1962_16226# a_19030_16186# 0.27fF
C14916 a_9994_12170# row_n[10] 0.17fF
C14917 a_8290_17230# vcm 0.22fF
C14918 a_23046_4138# a_24050_4138# 0.97fF
C14919 a_26058_10162# m2_26256_10410# 0.16fF
C14920 a_25054_2130# row_n[0] 0.17fF
C14921 a_18330_2170# vcm 0.22fF
C14922 a_2346_13216# a_14010_13174# 0.19fF
C14923 a_1962_13214# a_12306_13214# 0.14fF
C14924 a_25054_14178# a_25054_13174# 1.00fF
C14925 a_2346_5184# col[5] 0.15fF
C14926 col[12] rowoff_n[5] 0.11fF
C14927 col[11] rowoff_n[4] 0.11fF
C14928 col[13] rowoff_n[6] 0.11fF
C14929 col[10] rowoff_n[3] 0.11fF
C14930 col[8] rowoff_n[1] 0.11fF
C14931 col[15] rowoff_n[8] 0.11fF
C14932 col[9] rowoff_n[2] 0.11fF
C14933 col[7] rowoff_n[0] 0.11fF
C14934 col[16] rowoff_n[9] 0.11fF
C14935 col[14] rowoff_n[7] 0.11fF
C14936 a_9994_13174# col_n[7] 0.28fF
C14937 a_7894_4138# VDD 0.23fF
C14938 m2_1732_1950# row_n[0] 0.13fF
C14939 m3_1864_3086# VDD 0.25fF
C14940 a_1962_7190# col_n[21] 0.13fF
C14941 a_29070_15182# row_n[13] 0.17fF
C14942 a_31382_6186# vcm 0.22fF
C14943 a_14922_15182# a_15014_15182# 0.26fF
C14944 a_1962_15222# a_25358_15222# 0.14fF
C14945 a_2346_15224# a_27062_15182# 0.19fF
C14946 a_1962_1166# col[12] 0.11fF
C14947 a_28066_9158# col_n[25] 0.28fF
C14948 a_1962_14218# col[14] 0.11fF
C14949 a_20946_8154# VDD 0.23fF
C14950 a_1962_7190# a_2966_7150# 0.27fF
C14951 a_1962_15222# m2_1732_15002# 0.15fF
C14952 sample_n rowoff_n[14] 0.38fF
C14953 m2_12776_946# m3_13912_1078# 0.13fF
C14954 col[0] rowoff_n[10] 0.11fF
C14955 a_7986_5142# rowoff_n[3] 0.10fF
C14956 a_26058_4138# ctop 3.58fF
C14957 a_23046_11166# m2_23244_11414# 0.16fF
C14958 a_17022_13174# rowon_n[11] 0.14fF
C14959 a_33998_12170# VDD 0.23fF
C14960 m2_24824_946# m3_23952_1078# 0.13fF
C14961 a_2346_9200# a_16930_9158# 0.35fF
C14962 a_8990_9158# a_9994_9158# 0.97fF
C14963 a_6982_3134# vcm 0.62fF
C14964 a_10998_2130# col_n[8] 0.28fF
C14965 a_32082_3134# rowon_n[1] 0.14fF
C14966 a_18026_3134# rowoff_n[1] 0.10fF
C14967 a_33086_14178# rowoff_n[12] 0.10fF
C14968 a_7986_16186# col[5] 0.29fF
C14969 a_1962_6186# a_10998_6146# 0.27fF
C14970 a_1962_3174# col_n[12] 0.13fF
C14971 col_n[6] col[7] 5.98fF
C14972 vcm col[13] 5.84fF
C14973 col_n[22] row_n[0] 0.23fF
C14974 col_n[28] row_n[3] 0.23fF
C14975 a_1962_16226# col_n[14] 0.13fF
C14976 col_n[16] en_bit_n[2] 0.17fF
C14977 col_n[19] ctop 2.02fF
C14978 col_n[30] row_n[4] 0.23fF
C14979 VDD col[17] 4.18fF
C14980 rowon_n[10] row_n[10] 19.75fF
C14981 col_n[26] row_n[2] 0.23fF
C14982 col_n[24] row_n[1] 0.23fF
C14983 a_13006_15182# VDD 0.52fF
C14984 a_2346_11208# a_29982_11166# 0.35fF
C14985 a_9994_3134# row_n[1] 0.17fF
C14986 a_20034_7150# vcm 0.62fF
C14987 a_30074_2130# m2_30272_2378# 0.16fF
C14988 a_26058_12170# col[23] 0.29fF
C14989 a_1962_10202# col[5] 0.11fF
C14990 a_3270_16226# vcm 0.22fF
C14991 a_21038_4138# a_21038_3134# 1.00fF
C14992 a_1962_3174# a_4274_3174# 0.14fF
C14993 a_2346_3176# a_5978_3134# 0.19fF
C14994 a_1962_8194# a_24050_8154# 0.27fF
C14995 a_13310_1166# vcm 0.23fF
C14996 a_22042_13174# a_23046_13174# 0.97fF
C14997 a_2346_9200# col[25] 0.15fF
C14998 a_33086_11166# vcm 0.62fF
C14999 m2_34864_1950# ctop 0.18fF
C15000 a_6890_11166# rowoff_n[9] 0.24fF
C15001 a_14010_16186# row_n[14] 0.17fF
C15002 a_1962_18234# col_n[24] 0.13fF
C15003 a_2346_3176# VDD 32.63fF
C15004 a_1962_5182# a_17326_5182# 0.14fF
C15005 a_20034_12170# m2_20232_12418# 0.16fF
C15006 a_10906_5142# a_10998_5142# 0.26fF
C15007 a_2346_5184# a_19030_5142# 0.19fF
C15008 a_29070_6146# row_n[4] 0.17fF
C15009 a_16930_9158# rowoff_n[7] 0.24fF
C15010 a_8990_5142# col[6] 0.29fF
C15011 a_26362_5182# vcm 0.22fF
C15012 m2_14784_946# col_n[12] 0.37fF
C15013 a_20946_15182# rowoff_n[13] 0.24fF
C15014 m2_1732_6970# rowoff_n[5] 0.12fF
C15015 m2_31852_18014# m3_31984_18146# 2.78fF
C15016 a_15926_7150# VDD 0.23fF
C15017 a_26970_7150# rowoff_n[5] 0.24fF
C15018 a_26058_14178# col_n[23] 0.28fF
C15019 a_34090_8154# a_34090_7150# 1.00fF
C15020 a_1962_12210# col_n[5] 0.13fF
C15021 a_2346_7192# a_32082_7150# 0.19fF
C15022 a_1962_7190# a_30378_7190# 0.14fF
C15023 a_17022_4138# rowon_n[2] 0.14fF
C15024 a_21038_3134# ctop 3.57fF
C15025 a_28978_11166# VDD 0.23fF
C15026 m3_24956_1078# m3_25960_1078# 0.22fF
C15027 a_23958_9158# a_24050_9158# 0.26fF
C15028 a_6982_9158# a_6982_8154# 1.00fF
C15029 a_2346_5184# col[16] 0.15fF
C15030 a_34394_3174# vcm 0.22fF
C15031 col[22] rowoff_n[4] 0.11fF
C15032 col[21] rowoff_n[3] 0.11fF
C15033 col[27] rowoff_n[9] 0.11fF
C15034 col[18] rowoff_n[0] 0.11fF
C15035 col[24] rowoff_n[6] 0.11fF
C15036 col[23] rowoff_n[5] 0.11fF
C15037 col[26] rowoff_n[8] 0.11fF
C15038 col[25] rowoff_n[7] 0.11fF
C15039 col[19] rowoff_n[1] 0.11fF
C15040 col[20] rowoff_n[2] 0.11fF
C15041 a_2346_1168# a_21950_1126# 0.35fF
C15042 a_8990_7150# col_n[6] 0.28fF
C15043 a_34090_7150# ctop 3.42fF
C15044 a_17022_13174# m2_17220_13422# 0.16fF
C15045 a_21038_17190# rowon_n[15] 0.14fF
C15046 a_2966_7150# m3_1864_7102# 0.14fF
C15047 a_7986_14178# VDD 0.52fF
C15048 a_1962_1166# col[23] 0.11fF
C15049 a_15014_6146# vcm 0.62fF
C15050 a_1962_14218# col[25] 0.11fF
C15051 a_1962_15222# a_8990_15182# 0.27fF
C15052 a_27062_3134# col_n[24] 0.28fF
C15053 a_7986_16186# rowoff_n[14] 0.10fF
C15054 a_2346_3176# a_35002_3134# 0.35fF
C15055 a_18026_3134# a_19030_3134# 0.97fF
C15056 a_23046_2130# m3_22948_1078# 0.15fF
C15057 a_24050_17190# col[21] 0.29fF
C15058 a_1962_8194# VDD 2.73fF
C15059 col[11] rowoff_n[10] 0.11fF
C15060 m2_17796_18014# vcm 0.28fF
C15061 a_2346_12212# a_3970_12170# 0.19fF
C15062 a_20034_13174# a_20034_12170# 1.00fF
C15063 a_14010_7150# row_n[5] 0.17fF
C15064 a_28066_10162# vcm 0.62fF
C15065 a_1962_17230# a_22042_17190# 0.27fF
C15066 m2_29844_18014# m2_30272_18442# 0.16fF
C15067 a_31078_3134# VDD 0.52fF
C15068 m3_2868_2082# ctop 0.46fF
C15069 a_2346_1168# col[7] 0.14fF
C15070 a_2346_14220# col[9] 0.15fF
C15071 a_21342_4178# vcm 0.22fF
C15072 a_1962_14218# a_15318_14218# 0.14fF
C15073 a_2346_14220# a_17022_14178# 0.19fF
C15074 a_9902_14178# a_9994_14178# 0.26fF
C15075 m2_34864_5966# VDD 1.03fF
C15076 a_1962_3174# col_n[23] 0.13fF
C15077 a_6982_10162# col[4] 0.29fF
C15078 col_n[30] ctop 2.00fF
C15079 VDD col[28] 4.17fF
C15080 vcm col[24] 5.84fF
C15081 col_n[31] sw_n 0.39fF
C15082 col_n[12] col[12] 0.72fF
C15083 a_1962_16226# col_n[25] 0.13fF
C15084 a_10906_6146# VDD 0.23fF
C15085 a_14010_14178# m2_14208_14426# 0.16fF
C15086 a_31078_7150# a_32082_7150# 0.97fF
C15087 a_33086_10162# row_n[8] 0.17fF
C15088 a_5978_17190# ctop 3.39fF
C15089 a_1962_10202# col[16] 0.11fF
C15090 a_35398_8194# vcm 0.23fF
C15091 a_1962_16226# a_28370_16226# 0.14fF
C15092 a_2346_16228# a_30074_16186# 0.19fF
C15093 a_33086_17190# a_33086_16186# 1.00fF
C15094 a_25054_6146# col[22] 0.29fF
C15095 a_16018_2130# ctop 3.39fF
C15096 m2_8760_18014# VDD 0.91fF
C15097 a_35002_10162# m2_34864_9982# 0.16fF
C15098 a_1962_18234# m2_23820_18014# 0.18fF
C15099 a_23958_10162# VDD 0.23fF
C15100 a_3970_8154# a_4974_8154# 0.97fF
C15101 a_2346_8196# a_6890_8154# 0.35fF
C15102 m2_1732_2954# ctop 0.17fF
C15103 a_9902_4138# rowoff_n[2] 0.24fF
C15104 a_22954_12170# rowoff_n[10] 0.24fF
C15105 a_21038_8154# rowon_n[6] 0.14fF
C15106 a_29070_6146# ctop 3.58fF
C15107 a_2874_13174# VDD 0.24fF
C15108 a_2346_18236# m2_18800_18014# 0.19fF
C15109 a_6982_12170# col_n[4] 0.28fF
C15110 a_2346_10204# a_19942_10162# 0.35fF
C15111 a_2346_10204# col[0] 0.15fF
C15112 a_19942_2130# rowoff_n[0] 0.24fF
C15113 a_9994_5142# vcm 0.62fF
C15114 a_1962_12210# col_n[16] 0.13fF
C15115 a_16018_3134# a_16018_2130# 1.00fF
C15116 a_32994_3134# a_33086_3134# 0.26fF
C15117 m2_7756_18014# m3_8892_18146# 0.13fF
C15118 a_19030_1126# m3_18932_1078# 1.39fF
C15119 a_25054_8154# col_n[22] 0.28fF
C15120 a_1962_7190# a_14010_7150# 0.27fF
C15121 a_10998_15182# m2_11196_15430# 0.16fF
C15122 a_16018_17190# VDD 0.55fF
C15123 a_2346_12212# a_32994_12170# 0.35fF
C15124 a_17022_12170# a_18026_12170# 0.97fF
C15125 a_1962_6186# col[7] 0.11fF
C15126 a_23046_9158# vcm 0.62fF
C15127 a_13006_3134# m2_13204_3382# 0.16fF
C15128 a_2966_3134# ctop 3.24fF
C15129 a_6282_18234# vcm 0.22fF
C15130 a_26058_2130# VDD 0.55fF
C15131 a_2346_4180# a_8990_4138# 0.19fF
C15132 a_1962_4178# a_7286_4178# 0.14fF
C15133 a_5886_4138# a_5978_4138# 0.26fF
C15134 a_2346_5184# col[27] 0.15fF
C15135 m3_1864_7102# m3_1864_6098# 0.22fF
C15136 a_1962_9198# a_27062_9158# 0.27fF
C15137 col[31] rowoff_n[2] 0.11fF
C15138 col[30] rowoff_n[1] 0.11fF
C15139 col[29] rowoff_n[0] 0.11fF
C15140 a_16322_3174# vcm 0.22fF
C15141 a_18026_11166# row_n[9] 0.17fF
C15142 a_7986_10162# rowoff_n[8] 0.10fF
C15143 a_9994_13174# rowoff_n[11] 0.10fF
C15144 a_2346_12212# vcm 0.40fF
C15145 a_2346_1168# a_3878_1126# 0.39fF
C15146 a_5886_5142# VDD 0.23fF
C15147 a_2966_13174# m2_1732_12994# 0.96fF
C15148 a_2346_6188# a_22042_6146# 0.19fF
C15149 a_1962_6186# a_20338_6186# 0.14fF
C15150 a_29070_7150# a_29070_6146# 1.00fF
C15151 a_2966_17190# rowon_n[15] 0.13fF
C15152 a_4974_15182# col[2] 0.29fF
C15153 a_18026_8154# rowoff_n[6] 0.10fF
C15154 a_29374_7190# vcm 0.22fF
C15155 a_30074_16186# a_31078_16186# 0.97fF
C15156 a_1962_1166# m2_7756_946# 0.18fF
C15157 m2_24824_946# col[22] 0.39fF
C15158 a_1962_8194# col_n[7] 0.13fF
C15159 a_24050_17190# rowoff_n[15] 0.10fF
C15160 a_28066_6146# rowoff_n[4] 0.10fF
C15161 a_23046_11166# col[20] 0.29fF
C15162 a_18938_9158# VDD 0.23fF
C15163 a_5978_9158# rowon_n[7] 0.14fF
C15164 col[22] rowoff_n[10] 0.11fF
C15165 a_1962_8194# a_33390_8194# 0.14fF
C15166 a_18938_8154# a_19030_8154# 0.26fF
C15167 a_7986_16186# m2_8184_16434# 0.16fF
C15168 m2_15788_946# ctop 0.18fF
C15169 a_1962_18234# a_9294_18234# 0.14fF
C15170 a_1962_15222# col[0] 0.11fF
C15171 m2_6752_946# m2_7180_1374# 0.16fF
C15172 m2_1732_3958# rowon_n[2] 0.11fF
C15173 a_2346_17232# a_4882_17190# 0.35fF
C15174 m2_11772_18014# m2_12776_18014# 0.96fF
C15175 a_9994_4138# m2_10192_4386# 0.16fF
C15176 a_24050_5142# ctop 3.58fF
C15177 m2_32856_946# ctop 0.28fF
C15178 a_2346_1168# col[18] 0.14fF
C15179 a_2346_14220# col[20] 0.15fF
C15180 a_31990_13174# VDD 0.23fF
C15181 a_4974_4138# vcm 0.62fF
C15182 a_4974_17190# col_n[2] 0.28fF
C15183 col_n[17] col[18] 6.01fF
C15184 row_n[11] ctop 1.65fF
C15185 a_25054_12170# rowon_n[10] 0.14fF
C15186 a_5978_4138# col[3] 0.29fF
C15187 a_13006_2130# a_14010_2130# 0.97fF
C15188 a_2346_2172# a_24962_2130# 0.35fF
C15189 col[6] rowoff_n[11] 0.11fF
C15190 a_1962_10202# col[27] 0.11fF
C15191 a_10998_16186# VDD 0.52fF
C15192 a_15014_12170# a_15014_11166# 1.00fF
C15193 a_31990_12170# a_32082_12170# 0.26fF
C15194 a_23046_13174# col_n[20] 0.28fF
C15195 a_18026_8154# vcm 0.62fF
C15196 a_1962_16226# a_12002_16186# 0.27fF
C15197 a_1962_4178# sample 0.14fF
C15198 a_1962_17230# vcm 6.95fF
C15199 a_2966_4138# a_2966_3134# 1.00fF
C15200 a_18026_2130# row_n[0] 0.17fF
C15201 a_4974_17190# m2_5172_17438# 0.16fF
C15202 a_16018_17190# m2_15788_18014# 1.00fF
C15203 m2_2736_946# col_n[0] 0.37fF
C15204 a_11302_2170# vcm 0.22fF
C15205 a_1962_13214# a_5278_13214# 0.14fF
C15206 a_4882_13174# a_4974_13174# 0.26fF
C15207 a_2346_13216# a_6982_13174# 0.19fF
C15208 a_31078_12170# vcm 0.62fF
C15209 a_2966_8154# rowon_n[6] 0.13fF
C15210 a_6982_5142# m2_7180_5390# 0.16fF
C15211 a_34090_5142# VDD 0.54fF
C15212 m3_1864_17142# VDD 0.26fF
C15213 a_26058_6146# a_27062_6146# 0.97fF
C15214 a_2346_10204# col[11] 0.15fF
C15215 a_5978_6146# col_n[3] 0.28fF
C15216 m2_21812_946# a_21950_1126# 0.16fF
C15217 a_2966_16186# m3_1864_16138# 0.14fF
C15218 a_22042_15182# row_n[13] 0.17fF
C15219 a_24354_6186# vcm 0.22fF
C15220 a_2346_15224# a_20034_15182# 0.19fF
C15221 a_28066_16186# a_28066_15182# 1.00fF
C15222 a_1962_15222# a_18330_15222# 0.14fF
C15223 a_1962_12210# col_n[27] 0.13fF
C15224 a_24050_2130# col_n[21] 0.28fF
C15225 a_13918_8154# VDD 0.23fF
C15226 a_1962_6186# col[18] 0.11fF
C15227 a_21038_16186# col[18] 0.29fF
C15228 a_2346_17232# a_33086_17190# 0.19fF
C15229 a_1962_17230# a_31382_17230# 0.14fF
C15230 a_17934_17190# a_18026_17190# 0.26fF
C15231 m2_8760_946# m3_7888_1078# 0.13fF
C15232 a_19030_4138# ctop 3.58fF
C15233 a_9994_13174# rowon_n[11] 0.14fF
C15234 a_26970_12170# VDD 0.23fF
C15235 m3_20940_18146# m3_21944_18146# 0.22fF
C15236 a_2346_9200# a_9902_9158# 0.35fF
C15237 a_25054_3134# rowon_n[1] 0.14fF
C15238 a_10998_3134# rowoff_n[1] 0.10fF
C15239 a_26058_14178# rowoff_n[12] 0.10fF
C15240 a_3970_6146# m2_4168_6394# 0.16fF
C15241 a_27974_2130# a_28066_2130# 0.26fF
C15242 a_32082_8154# ctop 3.58fF
C15243 a_2346_6188# col[2] 0.15fF
C15244 a_1962_6186# a_3970_6146# 0.27fF
C15245 a_3970_9158# col[1] 0.29fF
C15246 a_5978_15182# VDD 0.52fF
C15247 a_2346_11208# a_22954_11166# 0.35fF
C15248 a_12002_11166# a_13006_11166# 0.97fF
C15249 a_1962_8194# col_n[18] 0.13fF
C15250 a_13006_7150# vcm 0.62fF
C15251 a_29070_16186# rowon_n[14] 0.14fF
C15252 a_1962_9198# m2_34864_8978# 0.17fF
C15253 a_22042_5142# col[19] 0.29fF
C15254 a_1962_2170# col[9] 0.11fF
C15255 a_1962_15222# col[11] 0.11fF
C15256 a_1962_8194# a_17022_8154# 0.27fF
C15257 a_6282_1166# vcm 0.23fF
C15258 a_26058_11166# vcm 0.62fF
C15259 a_2346_1168# col[29] 0.14fF
C15260 a_6982_16186# row_n[14] 0.17fF
C15261 a_2346_14220# col[31] 0.15fF
C15262 a_29070_4138# VDD 0.52fF
C15263 a_1962_5182# a_10298_5182# 0.14fF
C15264 a_24050_6146# a_24050_5142# 1.00fF
C15265 a_2346_5184# a_12002_5142# 0.19fF
C15266 a_2346_18236# col[3] 0.14fF
C15267 a_22042_6146# row_n[4] 0.17fF
C15268 a_1962_10202# a_30074_10162# 0.27fF
C15269 rowon_n[5] ctop 1.40fF
C15270 rowon_n[2] rowon_n[1] 0.15fF
C15271 col_n[23] col[23] 0.72fF
C15272 a_9902_9158# rowoff_n[7] 0.24fF
C15273 a_19334_5182# vcm 0.22fF
C15274 a_25054_15182# a_26058_15182# 0.97fF
C15275 a_3970_11166# col_n[1] 0.28fF
C15276 col[17] rowoff_n[11] 0.11fF
C15277 a_13918_15182# rowoff_n[13] 0.24fF
C15278 m2_1732_8978# VDD 1.02fF
C15279 m2_22816_18014# m3_21944_18146# 0.13fF
C15280 a_8898_7150# VDD 0.23fF
C15281 a_19942_7150# rowoff_n[5] 0.24fF
C15282 a_13918_7150# a_14010_7150# 0.26fF
C15283 a_1962_7190# a_23350_7190# 0.14fF
C15284 a_2346_7192# a_25054_7150# 0.19fF
C15285 a_22042_7150# col_n[19] 0.28fF
C15286 a_1962_4178# col_n[9] 0.13fF
C15287 a_1962_17230# col_n[11] 0.13fF
C15288 a_32386_9198# vcm 0.22fF
C15289 a_9994_4138# rowon_n[2] 0.14fF
C15290 a_29982_5142# rowoff_n[3] 0.24fF
C15291 a_14010_3134# ctop 3.57fF
C15292 a_1962_11206# col[2] 0.11fF
C15293 a_21950_11166# VDD 0.23fF
C15294 m3_10900_1078# m3_11904_1078# 0.22fF
C15295 col[1] rowoff_n[12] 0.11fF
C15296 a_2346_10204# col[22] 0.15fF
C15297 a_2346_1168# a_14922_1126# 0.35fF
C15298 a_27062_7150# ctop 3.58fF
C15299 a_14010_17190# rowon_n[15] 0.14fF
C15300 a_35002_15182# VDD 0.29fF
C15301 a_9994_11166# a_9994_10162# 1.00fF
C15302 a_26970_11166# a_27062_11166# 0.26fF
C15303 a_7986_6146# vcm 0.62fF
C15304 a_29070_7150# rowon_n[5] 0.14fF
C15305 m2_1732_10986# m2_2160_11414# 0.16fF
C15306 a_1962_6186# col[29] 0.11fF
C15307 a_32082_9158# m2_32280_9406# 0.16fF
C15308 a_2346_3176# a_27974_3134# 0.35fF
C15309 a_20034_10162# col[17] 0.29fF
C15310 m2_3740_18014# vcm 0.28fF
C15311 a_6982_7150# row_n[5] 0.17fF
C15312 a_1962_13214# col_n[2] 0.13fF
C15313 a_21038_10162# vcm 0.62fF
C15314 a_28066_11166# rowoff_n[9] 0.10fF
C15315 a_1962_17230# a_15014_17190# 0.27fF
C15316 m2_5748_18014# col[3] 0.28fF
C15317 m2_22816_18014# m2_23244_18442# 0.16fF
C15318 a_24050_3134# VDD 0.52fF
C15319 m3_34996_16138# ctop 0.23fF
C15320 a_2966_11166# m2_3164_11414# 0.16fF
C15321 a_21038_5142# a_22042_5142# 0.97fF
C15322 a_14314_4178# vcm 0.22fF
C15323 a_1962_14218# a_8290_14218# 0.14fF
C15324 a_2346_14220# a_9994_14178# 0.19fF
C15325 a_23046_15182# a_23046_14178# 1.00fF
C15326 a_2346_6188# col[13] 0.15fF
C15327 a_34090_14178# vcm 0.62fF
C15328 m2_1732_15002# m3_1864_16138# 0.15fF
C15329 a_26058_10162# row_n[8] 0.17fF
C15330 a_1962_8194# col_n[29] 0.13fF
C15331 a_2966_11166# a_3970_11166# 0.97fF
C15332 a_27366_8194# vcm 0.22fF
C15333 a_1962_16226# a_21342_16226# 0.14fF
C15334 a_2346_16228# a_23046_16186# 0.19fF
C15335 a_12914_16186# a_13006_16186# 0.26fF
C15336 a_20034_12170# col_n[17] 0.28fF
C15337 m2_34864_15002# m2_34864_13998# 0.99fF
C15338 a_1962_2170# col[20] 0.11fF
C15339 a_8990_2130# ctop 3.39fF
C15340 a_1962_15222# col[22] 0.11fF
C15341 a_1962_18234# m2_9764_18014# 0.18fF
C15342 a_29070_10162# m2_29268_10410# 0.16fF
C15343 a_16930_10162# VDD 0.23fF
C15344 m2_21812_18014# col_n[19] 0.25fF
C15345 a_2346_4180# rowoff_n[2] 4.09fF
C15346 a_15926_12170# rowoff_n[10] 0.24fF
C15347 a_14010_8154# rowon_n[6] 0.14fF
C15348 a_2346_18236# col[14] 0.14fF
C15349 a_22042_6146# ctop 3.58fF
C15350 m3_11904_1078# VDD 0.14fF
C15351 a_34090_13174# m2_34864_12994# 0.96fF
C15352 sw sw_n 0.22fF
C15353 col_n[28] col[29] 5.91fF
C15354 row_n[0] ctop 1.39fF
C15355 a_2346_18236# m2_4744_18014# 0.19fF
C15356 a_29982_14178# VDD 0.23fF
C15357 a_2346_10204# a_12914_10162# 0.35fF
C15358 a_6982_10162# a_7986_10162# 0.97fF
C15359 a_12914_2130# rowoff_n[0] 0.24fF
C15360 col[28] rowoff_n[11] 0.11fF
C15361 a_2346_2172# col[4] 0.15fF
C15362 a_2346_15224# col[6] 0.15fF
C15363 a_29982_16186# rowoff_n[14] 0.24fF
C15364 m2_31852_18014# ctop 0.18fF
C15365 a_1962_7190# a_6982_7150# 0.27fF
C15366 a_1962_4178# col_n[20] 0.13fF
C15367 a_8990_17190# VDD 0.55fF
C15368 a_1962_17230# col_n[22] 0.13fF
C15369 a_2346_12212# a_25966_12170# 0.35fF
C15370 a_33086_11166# rowon_n[9] 0.14fF
C15371 a_16018_9158# vcm 0.62fF
C15372 a_18026_15182# col[15] 0.29fF
C15373 a_1962_11206# col[13] 0.11fF
C15374 a_19030_2130# VDD 0.54fF
C15375 a_26058_11166# m2_26256_11414# 0.16fF
C15376 a_19030_5142# a_19030_4138# 1.00fF
C15377 a_3878_11166# VDD 0.23fF
C15378 m2_29844_946# m3_28972_1078# 0.13fF
C15379 m3_1864_14130# m3_1864_13126# 0.22fF
C15380 a_1962_9198# a_20034_9158# 0.27fF
C15381 a_14922_18194# m2_14784_18014# 0.16fF
C15382 col[12] rowoff_n[12] 0.11fF
C15383 a_2966_8154# col[0] 0.29fF
C15384 a_9294_3174# vcm 0.22fF
C15385 a_10998_11166# row_n[9] 0.17fF
C15386 a_20034_14178# a_21038_14178# 0.97fF
C15387 a_29070_13174# vcm 0.62fF
C15388 a_2874_13174# rowoff_n[11] 0.24fF
C15389 m2_1732_11990# m3_1864_13126# 0.15fF
C15390 a_32082_6146# VDD 0.52fF
C15391 a_8898_6146# a_8990_6146# 0.26fF
C15392 a_2346_6188# a_15014_6146# 0.19fF
C15393 a_1962_6186# a_13310_6186# 0.14fF
C15394 a_10998_8154# rowoff_n[6] 0.10fF
C15395 a_1962_11206# a_33086_11166# 0.27fF
C15396 a_22346_7190# vcm 0.22fF
C15397 a_33086_2130# m2_33284_2378# 0.16fF
C15398 a_17022_17190# rowoff_n[15] 0.10fF
C15399 a_3970_1126# ctop 0.57fF
C15400 a_21038_6146# rowoff_n[4] 0.10fF
C15401 a_3970_2130# m3_2868_2082# 0.14fF
C15402 a_18026_17190# col_n[15] 0.28fF
C15403 a_11910_9158# VDD 0.23fF
C15404 a_32082_9158# a_32082_8154# 1.00fF
C15405 a_1962_8194# a_26362_8194# 0.14fF
C15406 a_2346_8196# a_28066_8154# 0.19fF
C15407 a_1962_16226# m2_1732_16006# 0.15fF
C15408 a_1962_13214# col_n[13] 0.13fF
C15409 a_30074_14178# row_n[12] 0.17fF
C15410 a_19030_4138# col[16] 0.29fF
C15411 a_2966_10162# vcm 0.61fF
C15412 a_31078_4138# rowoff_n[2] 0.10fF
C15413 m2_8760_946# ctop 0.18fF
C15414 m2_4744_18014# m2_5748_18014# 0.96fF
C15415 a_1962_7190# col[4] 0.11fF
C15416 a_17022_5142# ctop 3.58fF
C15417 a_23046_12170# m2_23244_12418# 0.16fF
C15418 a_24962_13174# VDD 0.23fF
C15419 a_21950_10162# a_22042_10162# 0.26fF
C15420 a_4974_10162# a_4974_9158# 1.00fF
C15421 a_2346_6188# col[24] 0.15fF
C15422 m2_34864_15002# ctop 0.17fF
C15423 a_18026_12170# rowon_n[10] 0.14fF
C15424 a_2346_2172# a_17934_2130# 0.35fF
C15425 a_30074_9158# ctop 3.58fF
C15426 a_1962_7190# a_34394_7190# 0.14fF
C15427 a_34090_10162# m3_34996_10114# 0.13fF
C15428 a_33086_2130# rowon_n[0] 0.14fF
C15429 a_3970_16186# VDD 0.52fF
C15430 a_1962_2170# col[31] 0.11fF
C15431 a_10998_8154# vcm 0.62fF
C15432 a_1962_16226# a_4974_16186# 0.27fF
C15433 a_3878_16186# a_3970_16186# 0.26fF
C15434 a_19030_6146# col_n[16] 0.28fF
C15435 a_2346_4180# a_30986_4138# 0.35fF
C15436 a_16018_4138# a_17022_4138# 0.97fF
C15437 a_1962_9198# col_n[4] 0.13fF
C15438 a_10998_2130# row_n[0] 0.17fF
C15439 a_33998_18194# m2_33860_18014# 0.16fF
C15440 a_4274_2170# vcm 0.22fF
C15441 a_18026_14178# a_18026_13174# 1.00fF
C15442 a_29982_10162# rowoff_n[8] 0.24fF
C15443 a_2346_18236# col[25] 0.14fF
C15444 a_24050_12170# vcm 0.62fF
C15445 a_31990_13174# rowoff_n[11] 0.24fF
C15446 ctop col[2] 1.98fF
C15447 en_C0_n col[1] 0.16fF
C15448 a_34090_16186# col[31] 0.29fF
C15449 m2_1732_8978# m3_1864_10114# 0.15fF
C15450 a_27062_5142# VDD 0.52fF
C15451 m3_7888_18146# VDD 0.30fF
C15452 a_20034_13174# m2_20232_13422# 0.16fF
C15453 a_2346_2172# col[15] 0.15fF
C15454 a_15014_15182# row_n[13] 0.17fF
C15455 a_2346_15224# col[17] 0.15fF
C15456 a_17326_6186# vcm 0.22fF
C15457 a_7894_15182# a_7986_15182# 0.26fF
C15458 a_1962_15222# a_11302_15222# 0.14fF
C15459 a_2346_15224# a_13006_15182# 0.19fF
C15460 a_1962_4178# col_n[31] 0.13fF
C15461 a_30074_5142# row_n[3] 0.17fF
C15462 a_26058_2130# m3_25960_1078# 0.15fF
C15463 a_1962_17230# row_n[15] 25.57fF
C15464 a_6890_8154# VDD 0.23fF
C15465 a_29070_8154# a_30074_8154# 0.97fF
C15466 a_1962_18234# col[7] 0.11fF
C15467 a_1962_11206# col[24] 0.11fF
C15468 a_30378_10202# vcm 0.22fF
C15469 a_1962_17230# a_24354_17230# 0.14fF
C15470 a_2346_17232# a_26058_17190# 0.19fF
C15471 a_17022_9158# col[14] 0.29fF
C15472 a_12002_4138# ctop 3.58fF
C15473 m3_14916_1078# ctop 0.23fF
C15474 col[23] rowoff_n[12] 0.11fF
C15475 a_19942_12170# VDD 0.23fF
C15476 m3_6884_18146# m3_7888_18146# 0.22fF
C15477 a_18026_3134# rowon_n[1] 0.14fF
C15478 a_3970_3134# rowoff_n[1] 0.10fF
C15479 a_19030_14178# rowoff_n[12] 0.10fF
C15480 a_25054_8154# ctop 3.58fF
C15481 a_17022_14178# m2_17220_14426# 0.16fF
C15482 a_32994_16186# VDD 0.23fF
C15483 a_2346_11208# a_15926_11166# 0.35fF
C15484 a_2346_11208# col[8] 0.15fF
C15485 a_5978_7150# vcm 0.62fF
C15486 col[7] rowoff_n[13] 0.11fF
C15487 a_22042_16186# rowon_n[14] 0.14fF
C15488 a_14010_4138# a_14010_3134# 1.00fF
C15489 a_30986_4138# a_31078_4138# 0.26fF
C15490 a_2966_6146# rowoff_n[4] 0.10fF
C15491 a_1962_13214# col_n[24] 0.13fF
C15492 a_17022_11166# col_n[14] 0.28fF
C15493 a_1962_8194# a_9994_8154# 0.27fF
C15494 a_2346_13216# a_28978_13174# 0.35fF
C15495 a_15014_13174# a_16018_13174# 0.97fF
C15496 a_1962_7190# col[15] 0.11fF
C15497 a_19030_11166# vcm 0.62fF
C15498 m2_1732_5966# m3_1864_7102# 0.15fF
C15499 a_22042_4138# VDD 0.52fF
C15500 a_2346_5184# a_4974_5142# 0.19fF
C15501 a_1962_5182# a_3270_5182# 0.14fF
C15502 a_15014_6146# row_n[4] 0.17fF
.ends

