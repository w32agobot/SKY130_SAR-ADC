* SPICE3 file created from adc_array_wafflecap_16x544aF_41um2.ext - technology: sky130A

.subckt adc_array_wafflecap_16x544aF_41um2 cbot ctop
C0 cbot ctop 4.73fF
C1 cbot VSUBS 2.16fF
.ends
