magic
tech sky130A
timestamp 1663256564
<< psubdiff >>
rect -957 9110 -750 9274
rect -957 9093 -943 9110
rect -768 9093 -750 9110
rect -957 9070 -750 9093
rect -957 9053 -943 9070
rect -768 9053 -750 9070
rect -957 9030 -750 9053
rect -957 9013 -943 9030
rect -768 9013 -750 9030
rect -957 8990 -750 9013
rect -957 8973 -943 8990
rect -768 8973 -750 8990
rect -957 8950 -750 8973
rect -957 8933 -943 8950
rect -768 8933 -750 8950
rect -957 8910 -750 8933
rect -957 8893 -943 8910
rect -768 8893 -750 8910
rect -957 8870 -750 8893
rect -957 8853 -943 8870
rect -768 8853 -750 8870
rect -957 8830 -750 8853
rect -957 8813 -943 8830
rect -768 8813 -750 8830
rect -957 8790 -750 8813
rect -957 8773 -943 8790
rect -768 8773 -750 8790
rect -957 8750 -750 8773
rect -957 8733 -943 8750
rect -768 8733 -750 8750
rect -957 8710 -750 8733
rect -957 8693 -943 8710
rect -768 8693 -750 8710
rect -957 8670 -750 8693
rect -957 8653 -943 8670
rect -768 8653 -750 8670
rect -957 8630 -750 8653
rect -957 8613 -943 8630
rect -768 8613 -750 8630
rect -957 8590 -750 8613
rect -957 8573 -943 8590
rect -768 8573 -750 8590
rect -957 8550 -750 8573
rect -957 8533 -943 8550
rect -768 8533 -750 8550
rect -957 8510 -750 8533
rect -957 8493 -943 8510
rect -768 8493 -750 8510
rect -957 8470 -750 8493
rect -957 8453 -943 8470
rect -768 8453 -750 8470
rect -957 8430 -750 8453
rect -957 8413 -943 8430
rect -768 8413 -750 8430
rect -957 8390 -750 8413
rect -957 8373 -943 8390
rect -768 8373 -750 8390
rect -957 8350 -750 8373
rect -957 8333 -943 8350
rect -768 8333 -750 8350
rect -957 8310 -750 8333
rect -957 8293 -943 8310
rect -768 8293 -750 8310
rect -957 8270 -750 8293
rect -957 8253 -943 8270
rect -768 8253 -750 8270
rect -957 8230 -750 8253
rect -957 8213 -943 8230
rect -768 8213 -750 8230
rect -957 8190 -750 8213
rect -957 8173 -943 8190
rect -768 8173 -750 8190
rect -957 8150 -750 8173
rect -957 8133 -943 8150
rect -768 8133 -750 8150
rect -957 8110 -750 8133
rect -957 8093 -943 8110
rect -768 8093 -750 8110
rect -957 8070 -750 8093
rect -957 8053 -943 8070
rect -768 8053 -750 8070
rect -957 8030 -750 8053
rect -957 8013 -943 8030
rect -768 8013 -750 8030
rect -957 7990 -750 8013
rect -957 7973 -943 7990
rect -768 7973 -750 7990
rect -957 7950 -750 7973
rect -957 7933 -943 7950
rect -768 7933 -750 7950
rect -957 7910 -750 7933
rect -957 7893 -943 7910
rect -768 7893 -750 7910
rect -957 7870 -750 7893
rect -957 7853 -943 7870
rect -768 7853 -750 7870
rect -957 7830 -750 7853
rect -957 7813 -943 7830
rect -768 7813 -750 7830
rect -957 7790 -750 7813
rect -957 7773 -943 7790
rect -768 7773 -750 7790
rect -957 7750 -750 7773
rect -957 7733 -943 7750
rect -768 7733 -750 7750
rect -957 7710 -750 7733
rect -957 7693 -943 7710
rect -768 7693 -750 7710
rect -957 7670 -750 7693
rect -957 7653 -943 7670
rect -768 7653 -750 7670
rect -957 7630 -750 7653
rect -957 7613 -943 7630
rect -768 7613 -750 7630
rect -957 7590 -750 7613
rect -957 7573 -943 7590
rect -768 7573 -750 7590
rect -957 7550 -750 7573
rect -957 7533 -943 7550
rect -768 7533 -750 7550
rect -957 7510 -750 7533
rect -957 7493 -943 7510
rect -768 7493 -750 7510
rect -957 7470 -750 7493
rect -957 7453 -943 7470
rect -768 7453 -750 7470
rect -957 7430 -750 7453
rect -957 7413 -943 7430
rect -768 7413 -750 7430
rect -957 7390 -750 7413
rect -957 7373 -943 7390
rect -768 7373 -750 7390
rect -957 7350 -750 7373
rect -957 7333 -943 7350
rect -768 7333 -750 7350
rect -957 7310 -750 7333
rect -957 7293 -943 7310
rect -768 7293 -750 7310
rect -957 7270 -750 7293
rect -957 7253 -943 7270
rect -768 7253 -750 7270
rect -957 7230 -750 7253
rect -957 7213 -943 7230
rect -768 7213 -750 7230
rect -957 7190 -750 7213
rect -957 7173 -943 7190
rect -768 7173 -750 7190
rect -957 7150 -750 7173
rect -957 7133 -943 7150
rect -768 7133 -750 7150
rect -957 7110 -750 7133
rect -957 7093 -943 7110
rect -768 7093 -750 7110
rect -957 7070 -750 7093
rect -957 7053 -943 7070
rect -768 7053 -750 7070
rect -957 7030 -750 7053
rect -957 7013 -943 7030
rect -768 7013 -750 7030
rect -957 6990 -750 7013
rect -957 6973 -943 6990
rect -768 6973 -750 6990
rect -957 6950 -750 6973
rect -957 6933 -943 6950
rect -768 6933 -750 6950
rect -957 6910 -750 6933
rect -957 6893 -943 6910
rect -768 6893 -750 6910
rect -957 6870 -750 6893
rect -957 6853 -943 6870
rect -768 6853 -750 6870
rect -957 6830 -750 6853
rect -957 6813 -943 6830
rect -768 6813 -750 6830
rect -957 6790 -750 6813
rect -957 6773 -943 6790
rect -768 6773 -750 6790
rect -957 6750 -750 6773
rect -957 6733 -943 6750
rect -768 6733 -750 6750
rect -957 6710 -750 6733
rect -957 6693 -943 6710
rect -768 6693 -750 6710
rect -957 6670 -750 6693
rect -957 6653 -943 6670
rect -768 6653 -750 6670
rect -957 6630 -750 6653
rect -957 6613 -943 6630
rect -768 6613 -750 6630
rect -957 6590 -750 6613
rect -957 6573 -943 6590
rect -768 6573 -750 6590
rect -957 6550 -750 6573
rect -957 6533 -943 6550
rect -768 6533 -750 6550
rect -957 6510 -750 6533
rect -957 6493 -943 6510
rect -768 6493 -750 6510
rect -957 6470 -750 6493
rect -957 6453 -943 6470
rect -768 6453 -750 6470
rect -957 6430 -750 6453
rect -957 6413 -943 6430
rect -768 6413 -750 6430
rect -957 6390 -750 6413
rect -957 6373 -943 6390
rect -768 6373 -750 6390
rect -957 6350 -750 6373
rect -957 6333 -943 6350
rect -768 6333 -750 6350
rect -957 6310 -750 6333
rect -957 6293 -943 6310
rect -768 6293 -750 6310
rect -957 6270 -750 6293
rect -957 6253 -943 6270
rect -768 6253 -750 6270
rect -957 6230 -750 6253
rect -957 6213 -943 6230
rect -768 6213 -750 6230
rect -957 6190 -750 6213
rect -957 6173 -943 6190
rect -768 6173 -750 6190
rect -957 6150 -750 6173
rect -957 6133 -943 6150
rect -768 6133 -750 6150
rect -957 6110 -750 6133
rect -957 6093 -943 6110
rect -768 6093 -750 6110
rect -957 6070 -750 6093
rect -957 6053 -943 6070
rect -768 6053 -750 6070
rect -957 6030 -750 6053
rect -957 6013 -943 6030
rect -768 6013 -750 6030
rect -957 5990 -750 6013
rect -957 5973 -943 5990
rect -768 5973 -750 5990
rect -957 5950 -750 5973
rect -957 5933 -943 5950
rect -768 5933 -750 5950
rect -957 5910 -750 5933
rect -957 5893 -943 5910
rect -768 5893 -750 5910
rect -957 5870 -750 5893
rect -957 5853 -943 5870
rect -768 5853 -750 5870
rect -957 5830 -750 5853
rect -957 5813 -943 5830
rect -768 5813 -750 5830
rect -957 5790 -750 5813
rect -957 5773 -943 5790
rect -768 5773 -750 5790
rect -957 5750 -750 5773
rect -957 5733 -943 5750
rect -768 5733 -750 5750
rect -957 5710 -750 5733
rect -957 5693 -943 5710
rect -768 5693 -750 5710
rect -957 5670 -750 5693
rect -957 5653 -943 5670
rect -768 5653 -750 5670
rect -957 5630 -750 5653
rect -957 5613 -943 5630
rect -768 5613 -750 5630
rect -957 5590 -750 5613
rect -957 5573 -943 5590
rect -768 5573 -750 5590
rect -957 5550 -750 5573
rect -957 5533 -943 5550
rect -768 5533 -750 5550
rect -957 5510 -750 5533
rect -957 5493 -943 5510
rect -768 5493 -750 5510
rect -957 5470 -750 5493
rect -957 5453 -943 5470
rect -768 5453 -750 5470
rect -957 5430 -750 5453
rect -957 5413 -943 5430
rect -768 5413 -750 5430
rect -957 5390 -750 5413
rect -957 5373 -943 5390
rect -768 5373 -750 5390
rect -957 5350 -750 5373
rect -957 5333 -943 5350
rect -768 5333 -750 5350
rect -957 5310 -750 5333
rect -957 5293 -943 5310
rect -768 5293 -750 5310
rect -957 5270 -750 5293
rect -957 5253 -943 5270
rect -768 5253 -750 5270
rect -957 5230 -750 5253
rect -957 5213 -943 5230
rect -768 5213 -750 5230
rect -957 5190 -750 5213
rect -957 5173 -943 5190
rect -768 5173 -750 5190
rect -957 5150 -750 5173
rect -957 5133 -943 5150
rect -768 5133 -750 5150
rect -957 5110 -750 5133
rect -957 5093 -943 5110
rect -768 5093 -750 5110
rect -957 5070 -750 5093
rect -957 5053 -943 5070
rect -768 5053 -750 5070
rect -957 5030 -750 5053
rect -957 5013 -943 5030
rect -768 5013 -750 5030
rect -957 4990 -750 5013
rect -957 4973 -943 4990
rect -768 4973 -750 4990
rect -957 4950 -750 4973
rect -957 4933 -943 4950
rect -768 4933 -750 4950
rect -957 4910 -750 4933
rect -957 4893 -943 4910
rect -768 4893 -750 4910
rect -957 4870 -750 4893
rect -957 4853 -943 4870
rect -768 4853 -750 4870
rect -957 4830 -750 4853
rect -957 4813 -943 4830
rect -768 4813 -750 4830
rect -957 4790 -750 4813
rect -957 4773 -943 4790
rect -768 4773 -750 4790
rect -957 4750 -750 4773
rect -957 4733 -943 4750
rect -768 4733 -750 4750
rect -957 4710 -750 4733
rect -957 4693 -943 4710
rect -768 4693 -750 4710
rect -957 4670 -750 4693
rect -957 4653 -943 4670
rect -768 4653 -750 4670
rect -957 4630 -750 4653
rect -957 4613 -943 4630
rect -768 4613 -750 4630
rect -957 4590 -750 4613
rect -957 4573 -943 4590
rect -768 4573 -750 4590
rect -957 4550 -750 4573
rect -957 4533 -943 4550
rect -768 4533 -750 4550
rect -957 4510 -750 4533
rect -957 4493 -943 4510
rect -768 4493 -750 4510
rect -957 4470 -750 4493
rect -957 4453 -943 4470
rect -768 4453 -750 4470
rect -957 4430 -750 4453
rect -957 4413 -943 4430
rect -768 4413 -750 4430
rect -957 4390 -750 4413
rect -957 4373 -943 4390
rect -768 4373 -750 4390
rect -957 4350 -750 4373
rect -957 4333 -943 4350
rect -768 4333 -750 4350
rect -957 4310 -750 4333
rect -957 4293 -943 4310
rect -768 4293 -750 4310
rect -957 4270 -750 4293
rect -957 4253 -943 4270
rect -768 4253 -750 4270
rect -957 4230 -750 4253
rect -957 4213 -943 4230
rect -768 4213 -750 4230
rect -957 4190 -750 4213
rect -957 4173 -943 4190
rect -768 4173 -750 4190
rect -957 4150 -750 4173
rect -957 4133 -943 4150
rect -768 4133 -750 4150
rect -957 4110 -750 4133
rect -957 4093 -943 4110
rect -768 4093 -750 4110
rect -957 4070 -750 4093
rect -957 4053 -943 4070
rect -768 4053 -750 4070
rect -957 4030 -750 4053
rect -957 4013 -943 4030
rect -768 4013 -750 4030
rect -957 3990 -750 4013
rect -957 3973 -943 3990
rect -768 3973 -750 3990
rect -957 3950 -750 3973
rect -957 3933 -943 3950
rect -768 3933 -750 3950
rect -957 3910 -750 3933
rect -957 3893 -943 3910
rect -768 3893 -750 3910
rect -957 3870 -750 3893
rect -957 3853 -943 3870
rect -768 3853 -750 3870
rect -957 3830 -750 3853
rect -957 3813 -943 3830
rect -768 3813 -750 3830
rect -957 3790 -750 3813
rect -957 3773 -943 3790
rect -768 3773 -750 3790
rect -957 3750 -750 3773
rect -957 3733 -943 3750
rect -768 3733 -750 3750
rect -957 3710 -750 3733
rect -957 3693 -943 3710
rect -768 3693 -750 3710
rect -957 3670 -750 3693
rect -957 3653 -943 3670
rect -768 3653 -750 3670
rect -957 3630 -750 3653
rect -957 3613 -943 3630
rect -768 3613 -750 3630
rect -957 3590 -750 3613
rect -957 3573 -943 3590
rect -768 3573 -750 3590
rect -957 3550 -750 3573
rect -957 3533 -943 3550
rect -768 3533 -750 3550
rect -957 3510 -750 3533
rect -957 3493 -943 3510
rect -768 3493 -750 3510
rect -957 3470 -750 3493
rect -957 3453 -943 3470
rect -768 3453 -750 3470
rect -957 3430 -750 3453
rect -957 3413 -943 3430
rect -768 3413 -750 3430
rect -957 3390 -750 3413
rect -957 3373 -943 3390
rect -768 3373 -750 3390
rect -957 3350 -750 3373
rect -957 3333 -943 3350
rect -768 3333 -750 3350
rect -957 3310 -750 3333
rect -957 3293 -943 3310
rect -768 3293 -750 3310
rect -957 3270 -750 3293
rect -957 3253 -943 3270
rect -768 3253 -750 3270
rect -957 3230 -750 3253
rect -957 3213 -943 3230
rect -768 3213 -750 3230
rect -957 3190 -750 3213
rect -957 3173 -943 3190
rect -768 3173 -750 3190
rect -957 3150 -750 3173
rect -957 3133 -943 3150
rect -768 3133 -750 3150
rect -957 3110 -750 3133
rect -957 3093 -943 3110
rect -768 3093 -750 3110
rect -957 3070 -750 3093
rect -957 3053 -943 3070
rect -768 3053 -750 3070
rect -957 3030 -750 3053
rect -957 3013 -943 3030
rect -768 3013 -750 3030
rect -957 2990 -750 3013
rect -957 2973 -943 2990
rect -768 2973 -750 2990
rect -957 2950 -750 2973
rect -957 2933 -943 2950
rect -768 2933 -750 2950
rect -957 2910 -750 2933
rect -957 2893 -943 2910
rect -768 2893 -750 2910
rect -957 2870 -750 2893
rect -957 2853 -943 2870
rect -768 2853 -750 2870
rect -957 2830 -750 2853
rect -957 2813 -943 2830
rect -768 2813 -750 2830
rect -957 2790 -750 2813
rect -957 2773 -943 2790
rect -768 2773 -750 2790
rect -957 2750 -750 2773
rect -957 2733 -943 2750
rect -768 2733 -750 2750
rect -957 2710 -750 2733
rect -957 2693 -943 2710
rect -768 2693 -750 2710
rect -957 2670 -750 2693
rect -957 2653 -943 2670
rect -768 2653 -750 2670
rect -957 2630 -750 2653
rect -957 2613 -943 2630
rect -768 2613 -750 2630
rect -957 2590 -750 2613
rect -957 2573 -943 2590
rect -768 2573 -750 2590
rect -957 2550 -750 2573
rect -957 2533 -943 2550
rect -768 2533 -750 2550
rect -957 2510 -750 2533
rect -957 2493 -943 2510
rect -768 2493 -750 2510
rect -957 2470 -750 2493
rect -957 2453 -943 2470
rect -768 2453 -750 2470
rect -957 2430 -750 2453
rect -957 2413 -943 2430
rect -768 2413 -750 2430
rect -957 2390 -750 2413
rect -957 2373 -943 2390
rect -768 2373 -750 2390
rect -957 2350 -750 2373
rect -957 2333 -943 2350
rect -768 2333 -750 2350
rect -957 2310 -750 2333
rect -957 2293 -943 2310
rect -768 2293 -750 2310
rect -957 2270 -750 2293
rect -957 2253 -943 2270
rect -768 2253 -750 2270
rect -957 2230 -750 2253
rect -957 2213 -943 2230
rect -768 2213 -750 2230
rect -957 2190 -750 2213
rect -957 2173 -943 2190
rect -768 2173 -750 2190
rect -957 2150 -750 2173
rect -957 2133 -943 2150
rect -768 2133 -750 2150
rect -957 2110 -750 2133
rect -957 2093 -943 2110
rect -768 2093 -750 2110
rect -957 2070 -750 2093
rect -957 2053 -943 2070
rect -768 2053 -750 2070
rect -957 2030 -750 2053
rect -957 2013 -943 2030
rect -768 2013 -750 2030
rect -957 1990 -750 2013
rect -957 1973 -943 1990
rect -768 1973 -750 1990
rect -957 1950 -750 1973
rect -957 1933 -943 1950
rect -768 1933 -750 1950
rect -957 1910 -750 1933
rect -957 1893 -943 1910
rect -768 1893 -750 1910
rect -957 1870 -750 1893
rect -957 1853 -943 1870
rect -768 1853 -750 1870
rect -957 1830 -750 1853
rect -957 1813 -943 1830
rect -768 1813 -750 1830
rect -957 1790 -750 1813
rect -957 1773 -943 1790
rect -768 1773 -750 1790
rect -957 1750 -750 1773
rect -957 1733 -943 1750
rect -768 1733 -750 1750
rect -957 1710 -750 1733
rect -957 1693 -943 1710
rect -768 1693 -750 1710
rect -957 1670 -750 1693
rect -957 1653 -943 1670
rect -768 1653 -750 1670
rect -957 1630 -750 1653
rect -957 1613 -943 1630
rect -768 1613 -750 1630
rect -957 1590 -750 1613
rect -957 1573 -943 1590
rect -768 1573 -750 1590
rect -957 1550 -750 1573
rect -957 1533 -943 1550
rect -768 1533 -750 1550
rect -957 1510 -750 1533
rect -957 1493 -943 1510
rect -768 1493 -750 1510
rect -957 1470 -750 1493
rect -957 1453 -943 1470
rect -768 1453 -750 1470
rect -957 1430 -750 1453
rect -957 1413 -943 1430
rect -768 1413 -750 1430
rect -957 1390 -750 1413
rect -957 1373 -943 1390
rect -768 1373 -750 1390
rect -957 1350 -750 1373
rect -957 1333 -943 1350
rect -768 1333 -750 1350
rect -957 1310 -750 1333
rect -957 1293 -943 1310
rect -768 1293 -750 1310
rect -957 1270 -750 1293
rect -957 1253 -943 1270
rect -768 1253 -750 1270
rect -957 1230 -750 1253
rect -957 1213 -943 1230
rect -768 1213 -750 1230
rect -957 1190 -750 1213
rect -957 1173 -943 1190
rect -768 1173 -750 1190
rect -957 1150 -750 1173
rect -957 1133 -943 1150
rect -768 1133 -750 1150
rect -957 1110 -750 1133
rect -957 1093 -943 1110
rect -768 1093 -750 1110
rect -957 1070 -750 1093
rect -957 1053 -943 1070
rect -768 1053 -750 1070
rect -957 1030 -750 1053
rect -957 1013 -943 1030
rect -768 1013 -750 1030
rect -957 990 -750 1013
rect -957 973 -943 990
rect -768 973 -750 990
rect -957 950 -750 973
rect -957 933 -943 950
rect -768 933 -750 950
rect -957 910 -750 933
rect -957 893 -943 910
rect -768 893 -750 910
rect -957 870 -750 893
rect -957 853 -943 870
rect -768 853 -750 870
rect -957 830 -750 853
rect 17632 9110 17839 9274
rect 17632 9093 17650 9110
rect 17825 9093 17839 9110
rect 17632 9070 17839 9093
rect 17632 9053 17650 9070
rect 17825 9053 17839 9070
rect 17632 9030 17839 9053
rect 17632 9013 17650 9030
rect 17825 9013 17839 9030
rect 17632 8990 17839 9013
rect 17632 8973 17650 8990
rect 17825 8973 17839 8990
rect 17632 8950 17839 8973
rect 17632 8933 17650 8950
rect 17825 8933 17839 8950
rect 17632 8910 17839 8933
rect 17632 8893 17650 8910
rect 17825 8893 17839 8910
rect 17632 8874 17839 8893
rect 17632 8870 17840 8874
rect 17632 8853 17650 8870
rect 17825 8853 17840 8870
rect 17632 8830 17840 8853
rect 17632 8813 17650 8830
rect 17825 8813 17840 8830
rect 17632 8790 17840 8813
rect 17632 8773 17650 8790
rect 17825 8773 17840 8790
rect 17632 8750 17840 8773
rect 17632 8733 17650 8750
rect 17825 8733 17840 8750
rect 17632 8710 17839 8733
rect 17632 8693 17650 8710
rect 17825 8693 17839 8710
rect 17632 8670 17839 8693
rect 17632 8653 17650 8670
rect 17825 8653 17839 8670
rect 17632 8630 17839 8653
rect 17632 8613 17650 8630
rect 17825 8613 17839 8630
rect 17632 8590 17839 8613
rect 17632 8573 17650 8590
rect 17825 8573 17839 8590
rect 17632 8550 17839 8573
rect 17632 8533 17650 8550
rect 17825 8533 17839 8550
rect 17632 8510 17839 8533
rect 17632 8493 17650 8510
rect 17825 8493 17839 8510
rect 17632 8470 17839 8493
rect 17632 8453 17650 8470
rect 17825 8453 17839 8470
rect 17632 8430 17839 8453
rect 17632 8413 17650 8430
rect 17825 8413 17839 8430
rect 17632 8390 17839 8413
rect 17632 8373 17650 8390
rect 17825 8373 17839 8390
rect 17632 8350 17839 8373
rect 17632 8333 17650 8350
rect 17825 8333 17839 8350
rect 17632 8310 17839 8333
rect 17632 8293 17650 8310
rect 17825 8293 17839 8310
rect 17632 8270 17839 8293
rect 17632 8253 17650 8270
rect 17825 8253 17839 8270
rect 17632 8230 17839 8253
rect 17632 8213 17650 8230
rect 17825 8213 17839 8230
rect 17632 8190 17839 8213
rect 17632 8173 17650 8190
rect 17825 8173 17839 8190
rect 17632 8150 17839 8173
rect 17632 8133 17650 8150
rect 17825 8133 17839 8150
rect 17632 8110 17839 8133
rect 17632 8093 17650 8110
rect 17825 8093 17839 8110
rect 17632 8070 17839 8093
rect 17632 8053 17650 8070
rect 17825 8053 17839 8070
rect 17632 8030 17839 8053
rect 17632 8013 17650 8030
rect 17825 8013 17839 8030
rect 17632 7990 17839 8013
rect 17632 7973 17650 7990
rect 17825 7973 17839 7990
rect 17632 7950 17839 7973
rect 17632 7933 17650 7950
rect 17825 7933 17839 7950
rect 17632 7910 17839 7933
rect 17632 7893 17650 7910
rect 17825 7893 17839 7910
rect 17632 7870 17839 7893
rect 17632 7853 17650 7870
rect 17825 7853 17839 7870
rect 17632 7830 17839 7853
rect 17632 7813 17650 7830
rect 17825 7813 17839 7830
rect 17632 7790 17839 7813
rect 17632 7773 17650 7790
rect 17825 7773 17839 7790
rect 17632 7750 17839 7773
rect 17632 7733 17650 7750
rect 17825 7733 17839 7750
rect 17632 7710 17839 7733
rect 17632 7693 17650 7710
rect 17825 7693 17839 7710
rect 17632 7670 17839 7693
rect 17632 7653 17650 7670
rect 17825 7653 17839 7670
rect 17632 7630 17839 7653
rect 17632 7613 17650 7630
rect 17825 7613 17839 7630
rect 17632 7590 17839 7613
rect 17632 7573 17650 7590
rect 17825 7573 17839 7590
rect 17632 7550 17839 7573
rect 17632 7533 17650 7550
rect 17825 7533 17839 7550
rect 17632 7510 17839 7533
rect 17632 7493 17650 7510
rect 17825 7493 17839 7510
rect 17632 7470 17839 7493
rect 17632 7453 17650 7470
rect 17825 7453 17839 7470
rect 17632 7430 17839 7453
rect 17632 7413 17650 7430
rect 17825 7413 17839 7430
rect 17632 7390 17839 7413
rect 17632 7373 17650 7390
rect 17825 7373 17839 7390
rect 17632 7350 17839 7373
rect 17632 7333 17650 7350
rect 17825 7333 17839 7350
rect 17632 7310 17839 7333
rect 17632 7293 17650 7310
rect 17825 7293 17839 7310
rect 17632 7270 17839 7293
rect 17632 7253 17650 7270
rect 17825 7253 17839 7270
rect 17632 7230 17839 7253
rect 17632 7213 17650 7230
rect 17825 7213 17839 7230
rect 17632 7190 17839 7213
rect 17632 7173 17650 7190
rect 17825 7173 17839 7190
rect 17632 7150 17839 7173
rect 17632 7133 17650 7150
rect 17825 7133 17839 7150
rect 17632 7110 17839 7133
rect 17632 7093 17650 7110
rect 17825 7093 17839 7110
rect 17632 7070 17839 7093
rect 17632 7053 17650 7070
rect 17825 7053 17839 7070
rect 17632 7030 17839 7053
rect 17632 7013 17650 7030
rect 17825 7013 17839 7030
rect 17632 6990 17839 7013
rect 17632 6973 17650 6990
rect 17825 6973 17839 6990
rect 17632 6950 17839 6973
rect 17632 6933 17650 6950
rect 17825 6933 17839 6950
rect 17632 6910 17839 6933
rect 17632 6893 17650 6910
rect 17825 6893 17839 6910
rect 17632 6870 17839 6893
rect 17632 6853 17650 6870
rect 17825 6853 17839 6870
rect 17632 6830 17839 6853
rect 17632 6813 17650 6830
rect 17825 6813 17839 6830
rect 17632 6790 17839 6813
rect 17632 6773 17650 6790
rect 17825 6773 17839 6790
rect 17632 6750 17839 6773
rect 17632 6733 17650 6750
rect 17825 6733 17839 6750
rect 17632 6710 17839 6733
rect 17632 6693 17650 6710
rect 17825 6693 17839 6710
rect 17632 6670 17839 6693
rect 17632 6653 17650 6670
rect 17825 6653 17839 6670
rect 17632 6630 17839 6653
rect 17632 6613 17650 6630
rect 17825 6613 17839 6630
rect 17632 6590 17839 6613
rect 17632 6573 17650 6590
rect 17825 6573 17839 6590
rect 17632 6550 17839 6573
rect 17632 6533 17650 6550
rect 17825 6533 17839 6550
rect 17632 6510 17839 6533
rect 17632 6493 17650 6510
rect 17825 6493 17839 6510
rect 17632 6470 17839 6493
rect 17632 6453 17650 6470
rect 17825 6453 17839 6470
rect 17632 6430 17839 6453
rect 17632 6413 17650 6430
rect 17825 6413 17839 6430
rect 17632 6390 17839 6413
rect 17632 6373 17650 6390
rect 17825 6373 17839 6390
rect 17632 6350 17839 6373
rect 17632 6333 17650 6350
rect 17825 6333 17839 6350
rect 17632 6310 17839 6333
rect 17632 6293 17650 6310
rect 17825 6293 17839 6310
rect 17632 6270 17839 6293
rect 17632 6253 17650 6270
rect 17825 6253 17839 6270
rect 17632 6229 17839 6253
rect 17632 6212 17651 6229
rect 17826 6212 17839 6229
rect 17632 6190 17839 6212
rect 17632 6173 17650 6190
rect 17825 6173 17839 6190
rect 17632 6150 17839 6173
rect 17632 6133 17650 6150
rect 17825 6133 17839 6150
rect 17632 6110 17839 6133
rect 17632 6093 17650 6110
rect 17825 6093 17839 6110
rect 17632 6070 17839 6093
rect 17632 6053 17650 6070
rect 17825 6053 17839 6070
rect 17632 6030 17839 6053
rect 17632 6013 17650 6030
rect 17825 6013 17839 6030
rect 17632 5990 17839 6013
rect 17632 5973 17650 5990
rect 17825 5973 17839 5990
rect 17632 5950 17839 5973
rect 17632 5933 17650 5950
rect 17825 5933 17839 5950
rect 17632 5910 17839 5933
rect 17632 5893 17650 5910
rect 17825 5904 17839 5910
rect 17825 5893 17840 5904
rect 17632 5870 17840 5893
rect 17632 5853 17650 5870
rect 17825 5853 17840 5870
rect 17632 5830 17840 5853
rect 17632 5813 17650 5830
rect 17825 5813 17840 5830
rect 17632 5790 17840 5813
rect 17632 5773 17650 5790
rect 17825 5773 17840 5790
rect 17632 5763 17840 5773
rect 17632 5750 17839 5763
rect 17632 5733 17650 5750
rect 17825 5733 17839 5750
rect 17632 5710 17839 5733
rect 17632 5693 17650 5710
rect 17825 5693 17839 5710
rect 17632 5670 17839 5693
rect 17632 5653 17650 5670
rect 17825 5653 17839 5670
rect 17632 5630 17839 5653
rect 17632 5613 17650 5630
rect 17825 5613 17839 5630
rect 17632 5590 17839 5613
rect 17632 5573 17650 5590
rect 17825 5573 17839 5590
rect 17632 5550 17839 5573
rect 17632 5533 17650 5550
rect 17825 5533 17839 5550
rect 17632 5510 17839 5533
rect 17632 5493 17650 5510
rect 17825 5493 17839 5510
rect 17632 5470 17839 5493
rect 17632 5453 17650 5470
rect 17825 5453 17839 5470
rect 17632 5430 17839 5453
rect 17632 5413 17650 5430
rect 17825 5413 17839 5430
rect 17632 5390 17839 5413
rect 17632 5373 17650 5390
rect 17825 5373 17839 5390
rect 17632 5349 17839 5373
rect 17632 5332 17649 5349
rect 17824 5332 17839 5349
rect 17632 5310 17839 5332
rect 17632 5293 17650 5310
rect 17825 5293 17839 5310
rect 17632 5270 17839 5293
rect 17632 5253 17650 5270
rect 17825 5253 17839 5270
rect 17632 5230 17839 5253
rect 17632 5213 17650 5230
rect 17825 5213 17839 5230
rect 17632 5190 17839 5213
rect 17632 5173 17650 5190
rect 17825 5173 17839 5190
rect 17632 5150 17839 5173
rect 17632 5133 17650 5150
rect 17825 5133 17839 5150
rect 17632 5110 17839 5133
rect 17632 5093 17650 5110
rect 17825 5093 17839 5110
rect 17632 5070 17839 5093
rect 17632 5053 17650 5070
rect 17825 5053 17839 5070
rect 17632 5030 17839 5053
rect 17632 5013 17650 5030
rect 17825 5013 17839 5030
rect 17632 4990 17839 5013
rect 17632 4973 17650 4990
rect 17825 4973 17839 4990
rect 17632 4950 17839 4973
rect 17632 4933 17650 4950
rect 17825 4933 17839 4950
rect 17632 4910 17839 4933
rect 17632 4893 17650 4910
rect 17825 4893 17839 4910
rect 17632 4870 17839 4893
rect 17632 4853 17650 4870
rect 17825 4853 17839 4870
rect 17632 4830 17839 4853
rect 17632 4813 17650 4830
rect 17825 4813 17839 4830
rect 17632 4790 17839 4813
rect 17632 4773 17650 4790
rect 17825 4773 17839 4790
rect 17632 4750 17839 4773
rect 17632 4733 17650 4750
rect 17825 4733 17839 4750
rect 17632 4710 17839 4733
rect 17632 4693 17650 4710
rect 17825 4693 17839 4710
rect 17632 4670 17839 4693
rect 17632 4653 17650 4670
rect 17825 4653 17839 4670
rect 17632 4630 17839 4653
rect 17632 4613 17650 4630
rect 17825 4613 17839 4630
rect 17632 4590 17839 4613
rect 17632 4573 17650 4590
rect 17825 4573 17839 4590
rect 17632 4550 17839 4573
rect 17632 4533 17650 4550
rect 17825 4533 17839 4550
rect 17632 4510 17839 4533
rect 17632 4493 17650 4510
rect 17825 4493 17839 4510
rect 17632 4470 17839 4493
rect 17632 4453 17650 4470
rect 17825 4453 17839 4470
rect 17632 4430 17839 4453
rect 17632 4413 17650 4430
rect 17825 4413 17839 4430
rect 17632 4390 17839 4413
rect 17632 4373 17650 4390
rect 17825 4373 17839 4390
rect 17632 4350 17839 4373
rect 17632 4333 17650 4350
rect 17825 4333 17839 4350
rect 17632 4310 17839 4333
rect 17632 4293 17650 4310
rect 17825 4293 17839 4310
rect 17632 4270 17839 4293
rect 17632 4253 17650 4270
rect 17825 4253 17839 4270
rect 17632 4230 17839 4253
rect 17632 4213 17650 4230
rect 17825 4213 17839 4230
rect 17632 4190 17839 4213
rect 17632 4173 17650 4190
rect 17825 4173 17839 4190
rect 17632 4150 17839 4173
rect 17632 4133 17650 4150
rect 17825 4133 17839 4150
rect 17632 4110 17839 4133
rect 17632 4093 17650 4110
rect 17825 4093 17839 4110
rect 17632 4070 17839 4093
rect 17632 4053 17650 4070
rect 17825 4053 17839 4070
rect 17632 4030 17839 4053
rect 17632 4013 17650 4030
rect 17825 4013 17839 4030
rect 17632 3990 17839 4013
rect 17632 3973 17650 3990
rect 17825 3973 17839 3990
rect 17632 3950 17839 3973
rect 17632 3933 17650 3950
rect 17825 3933 17839 3950
rect 17632 3910 17839 3933
rect 17632 3893 17650 3910
rect 17825 3893 17839 3910
rect 17632 3870 17839 3893
rect 17632 3853 17650 3870
rect 17825 3853 17839 3870
rect 17632 3830 17840 3853
rect 17632 3813 17650 3830
rect 17825 3813 17840 3830
rect 17632 3790 17840 3813
rect 17632 3773 17650 3790
rect 17825 3773 17840 3790
rect 17632 3750 17840 3773
rect 17632 3733 17650 3750
rect 17825 3733 17840 3750
rect 17632 3712 17840 3733
rect 17632 3710 17839 3712
rect 17632 3693 17650 3710
rect 17825 3693 17839 3710
rect 17632 3670 17839 3693
rect 17632 3653 17650 3670
rect 17825 3653 17839 3670
rect 17632 3630 17839 3653
rect 17632 3613 17650 3630
rect 17825 3613 17839 3630
rect 17632 3590 17839 3613
rect 17632 3573 17650 3590
rect 17825 3573 17839 3590
rect 17632 3550 17839 3573
rect 17632 3533 17650 3550
rect 17825 3533 17839 3550
rect 17632 3510 17839 3533
rect 17632 3493 17650 3510
rect 17825 3493 17839 3510
rect 17632 3470 17839 3493
rect 17632 3453 17650 3470
rect 17825 3453 17839 3470
rect 17632 3430 17839 3453
rect 17632 3413 17650 3430
rect 17825 3413 17839 3430
rect 17632 3390 17839 3413
rect 17632 3373 17650 3390
rect 17825 3373 17839 3390
rect 17632 3350 17839 3373
rect 17632 3333 17650 3350
rect 17825 3333 17839 3350
rect 17632 3310 17839 3333
rect 17632 3293 17650 3310
rect 17825 3293 17839 3310
rect 17632 3270 17839 3293
rect 17632 3253 17650 3270
rect 17825 3253 17839 3270
rect 17632 3230 17839 3253
rect 17632 3213 17650 3230
rect 17825 3213 17839 3230
rect 17632 3190 17839 3213
rect 17632 3173 17650 3190
rect 17825 3173 17839 3190
rect 17632 3150 17839 3173
rect 17632 3133 17650 3150
rect 17825 3133 17839 3150
rect 17632 3110 17839 3133
rect 17632 3093 17650 3110
rect 17825 3093 17839 3110
rect 17632 3070 17839 3093
rect 17632 3053 17650 3070
rect 17825 3053 17839 3070
rect 17632 3030 17839 3053
rect 17632 3013 17650 3030
rect 17825 3013 17839 3030
rect 17632 2990 17839 3013
rect 17632 2973 17650 2990
rect 17825 2973 17839 2990
rect 17632 2950 17839 2973
rect 17632 2933 17650 2950
rect 17825 2933 17839 2950
rect 17632 2910 17839 2933
rect 17632 2893 17650 2910
rect 17825 2893 17839 2910
rect 17632 2870 17839 2893
rect 17632 2853 17650 2870
rect 17825 2853 17839 2870
rect 17632 2831 17839 2853
rect 17632 2830 17840 2831
rect 17632 2813 17650 2830
rect 17825 2813 17840 2830
rect 17632 2790 17840 2813
rect 17632 2773 17650 2790
rect 17825 2773 17840 2790
rect 17632 2750 17840 2773
rect 17632 2733 17650 2750
rect 17825 2733 17840 2750
rect 17632 2710 17840 2733
rect 17632 2693 17650 2710
rect 17825 2693 17840 2710
rect 17632 2690 17840 2693
rect 17632 2670 17839 2690
rect 17632 2653 17650 2670
rect 17825 2653 17839 2670
rect 17632 2630 17839 2653
rect 17632 2613 17650 2630
rect 17825 2613 17839 2630
rect 17632 2590 17839 2613
rect 17632 2573 17650 2590
rect 17825 2573 17839 2590
rect 17632 2550 17839 2573
rect 17632 2533 17650 2550
rect 17825 2533 17839 2550
rect 17632 2510 17839 2533
rect 17632 2493 17650 2510
rect 17825 2493 17839 2510
rect 17632 2470 17839 2493
rect 17632 2453 17650 2470
rect 17825 2453 17839 2470
rect 17632 2430 17839 2453
rect 17632 2413 17650 2430
rect 17825 2413 17839 2430
rect 17632 2390 17839 2413
rect 17632 2373 17650 2390
rect 17825 2373 17839 2390
rect 17632 2350 17839 2373
rect 17632 2333 17650 2350
rect 17825 2333 17839 2350
rect 17632 2310 17839 2333
rect 17632 2293 17650 2310
rect 17825 2293 17839 2310
rect 17632 2267 17839 2293
rect 17632 2250 17650 2267
rect 17825 2250 17839 2267
rect 17632 2230 17839 2250
rect 17632 2213 17650 2230
rect 17825 2213 17839 2230
rect 17632 2190 17839 2213
rect 17632 2173 17650 2190
rect 17825 2173 17839 2190
rect 17632 2150 17839 2173
rect 17632 2133 17650 2150
rect 17825 2133 17839 2150
rect 17632 2110 17839 2133
rect 17632 2093 17650 2110
rect 17825 2093 17839 2110
rect 17632 2070 17839 2093
rect 17632 2053 17650 2070
rect 17825 2053 17839 2070
rect 17632 2030 17839 2053
rect 17632 2013 17650 2030
rect 17825 2013 17839 2030
rect 17632 1990 17839 2013
rect 17632 1973 17650 1990
rect 17825 1973 17839 1990
rect 17632 1950 17839 1973
rect 17632 1933 17650 1950
rect 17825 1933 17839 1950
rect 17632 1910 17839 1933
rect 17632 1893 17650 1910
rect 17825 1893 17839 1910
rect 17632 1870 17839 1893
rect 17632 1853 17650 1870
rect 17825 1853 17839 1870
rect 17632 1830 17839 1853
rect 17632 1813 17650 1830
rect 17825 1813 17839 1830
rect 17632 1790 17839 1813
rect 17632 1773 17650 1790
rect 17825 1773 17839 1790
rect 17632 1750 17839 1773
rect 17632 1733 17650 1750
rect 17825 1733 17839 1750
rect 17632 1710 17839 1733
rect 17632 1693 17650 1710
rect 17825 1693 17839 1710
rect 17632 1670 17839 1693
rect 17632 1653 17650 1670
rect 17825 1653 17839 1670
rect 17632 1630 17839 1653
rect 17632 1613 17650 1630
rect 17825 1613 17839 1630
rect 17632 1590 17839 1613
rect 17632 1573 17650 1590
rect 17825 1573 17839 1590
rect 17632 1550 17839 1573
rect 17632 1533 17650 1550
rect 17825 1533 17839 1550
rect 17632 1510 17839 1533
rect 17632 1493 17650 1510
rect 17825 1493 17839 1510
rect 17632 1470 17839 1493
rect 17632 1453 17650 1470
rect 17825 1453 17839 1470
rect 17632 1430 17839 1453
rect 17632 1413 17650 1430
rect 17825 1413 17839 1430
rect 17632 1390 17839 1413
rect 17632 1373 17650 1390
rect 17825 1373 17839 1390
rect 17632 1350 17839 1373
rect 17632 1333 17650 1350
rect 17825 1333 17839 1350
rect 17632 1310 17839 1333
rect 17632 1293 17650 1310
rect 17825 1293 17839 1310
rect 17632 1270 17839 1293
rect 17632 1253 17650 1270
rect 17825 1253 17839 1270
rect 17632 1230 17839 1253
rect 17632 1213 17650 1230
rect 17825 1213 17839 1230
rect 17632 1190 17839 1213
rect 17632 1173 17650 1190
rect 17825 1173 17839 1190
rect 17632 1150 17839 1173
rect 17632 1133 17650 1150
rect 17825 1133 17839 1150
rect 17632 1110 17839 1133
rect 17632 1093 17650 1110
rect 17825 1093 17839 1110
rect 17632 1070 17839 1093
rect 17632 1053 17650 1070
rect 17825 1053 17839 1070
rect 17632 1030 17839 1053
rect 17632 1013 17650 1030
rect 17825 1013 17839 1030
rect 17632 990 17839 1013
rect 17632 973 17650 990
rect 17825 973 17839 990
rect 17632 950 17839 973
rect 17632 933 17650 950
rect 17825 933 17839 950
rect 17632 910 17839 933
rect 17632 893 17650 910
rect 17825 893 17839 910
rect 17632 870 17839 893
rect 17632 853 17650 870
rect 17825 853 17839 870
rect 17632 834 17839 853
rect -957 813 -943 830
rect -768 813 -750 830
rect -957 790 -750 813
rect -957 773 -943 790
rect -768 773 -750 790
rect -957 750 -750 773
rect -957 733 -943 750
rect -768 733 -750 750
rect -957 710 -750 733
rect -957 693 -943 710
rect -768 693 -750 710
rect 17631 830 17839 834
rect 17631 813 17650 830
rect 17825 813 17839 830
rect 17631 790 17839 813
rect 17631 773 17650 790
rect 17825 773 17839 790
rect 17631 750 17839 773
rect 17631 733 17650 750
rect 17825 733 17839 750
rect 17631 710 17839 733
rect 17631 693 17650 710
rect 17825 693 17839 710
rect -957 670 -750 693
rect -957 653 -943 670
rect -768 653 -750 670
rect -957 630 -750 653
rect -957 613 -943 630
rect -768 613 -750 630
rect -957 590 -750 613
rect -957 573 -943 590
rect -768 573 -750 590
rect -957 550 -750 573
rect -957 533 -943 550
rect -768 533 -750 550
rect -957 510 -750 533
rect -957 493 -943 510
rect -768 493 -750 510
rect -957 470 -750 493
rect -957 453 -943 470
rect -768 453 -750 470
rect -957 430 -750 453
rect -957 413 -943 430
rect -768 413 -750 430
rect -957 390 -750 413
rect -957 373 -943 390
rect -768 373 -750 390
rect -957 350 -750 373
rect -957 333 -943 350
rect -768 333 -750 350
rect -957 310 -750 333
rect -957 293 -943 310
rect -768 293 -750 310
rect -957 270 -750 293
rect -957 253 -943 270
rect -768 253 -750 270
rect -957 230 -750 253
rect -957 213 -943 230
rect -768 213 -750 230
rect -957 190 -750 213
rect -957 173 -943 190
rect -768 173 -750 190
rect -957 150 -750 173
rect -957 133 -943 150
rect -768 133 -750 150
rect -957 110 -750 133
rect -957 93 -943 110
rect -768 93 -750 110
rect -957 70 -750 93
rect -957 53 -943 70
rect -768 53 -750 70
rect -957 30 -750 53
rect -957 13 -943 30
rect -768 13 -750 30
rect -957 -217 -750 13
rect 17632 670 17839 693
rect 17632 653 17650 670
rect 17825 653 17839 670
rect 17632 630 17839 653
rect 17632 613 17650 630
rect 17825 613 17839 630
rect 17632 590 17839 613
rect 17632 573 17650 590
rect 17825 573 17839 590
rect 17632 550 17839 573
rect 17632 533 17650 550
rect 17825 533 17839 550
rect 17632 510 17839 533
rect 17632 493 17650 510
rect 17825 493 17839 510
rect 17632 470 17839 493
rect 17632 453 17650 470
rect 17825 453 17839 470
rect 17632 430 17839 453
rect 17632 413 17650 430
rect 17825 413 17839 430
rect 17632 390 17839 413
rect 17632 373 17650 390
rect 17825 373 17839 390
rect 17632 350 17839 373
rect 17632 333 17650 350
rect 17825 333 17839 350
rect 17632 310 17839 333
rect 17632 293 17650 310
rect 17825 293 17839 310
rect 17632 270 17839 293
rect 17632 253 17650 270
rect 17825 253 17839 270
rect 17632 230 17839 253
rect 17632 213 17650 230
rect 17825 213 17839 230
rect 17632 190 17839 213
rect 17632 173 17650 190
rect 17825 173 17839 190
rect 17632 150 17839 173
rect 17632 133 17650 150
rect 17825 133 17839 150
rect 17632 110 17839 133
rect 17632 93 17650 110
rect 17825 93 17839 110
rect 17632 70 17839 93
rect 17632 53 17650 70
rect 17825 53 17839 70
rect 17632 30 17839 53
rect 17632 13 17650 30
rect 17825 13 17839 30
rect 17632 -152 17839 13
<< psubdiffcont >>
rect -943 9093 -768 9110
rect -943 9053 -768 9070
rect -943 9013 -768 9030
rect -943 8973 -768 8990
rect -943 8933 -768 8950
rect -943 8893 -768 8910
rect -943 8853 -768 8870
rect -943 8813 -768 8830
rect -943 8773 -768 8790
rect -943 8733 -768 8750
rect -943 8693 -768 8710
rect -943 8653 -768 8670
rect -943 8613 -768 8630
rect -943 8573 -768 8590
rect -943 8533 -768 8550
rect -943 8493 -768 8510
rect -943 8453 -768 8470
rect -943 8413 -768 8430
rect -943 8373 -768 8390
rect -943 8333 -768 8350
rect -943 8293 -768 8310
rect -943 8253 -768 8270
rect -943 8213 -768 8230
rect -943 8173 -768 8190
rect -943 8133 -768 8150
rect -943 8093 -768 8110
rect -943 8053 -768 8070
rect -943 8013 -768 8030
rect -943 7973 -768 7990
rect -943 7933 -768 7950
rect -943 7893 -768 7910
rect -943 7853 -768 7870
rect -943 7813 -768 7830
rect -943 7773 -768 7790
rect -943 7733 -768 7750
rect -943 7693 -768 7710
rect -943 7653 -768 7670
rect -943 7613 -768 7630
rect -943 7573 -768 7590
rect -943 7533 -768 7550
rect -943 7493 -768 7510
rect -943 7453 -768 7470
rect -943 7413 -768 7430
rect -943 7373 -768 7390
rect -943 7333 -768 7350
rect -943 7293 -768 7310
rect -943 7253 -768 7270
rect -943 7213 -768 7230
rect -943 7173 -768 7190
rect -943 7133 -768 7150
rect -943 7093 -768 7110
rect -943 7053 -768 7070
rect -943 7013 -768 7030
rect -943 6973 -768 6990
rect -943 6933 -768 6950
rect -943 6893 -768 6910
rect -943 6853 -768 6870
rect -943 6813 -768 6830
rect -943 6773 -768 6790
rect -943 6733 -768 6750
rect -943 6693 -768 6710
rect -943 6653 -768 6670
rect -943 6613 -768 6630
rect -943 6573 -768 6590
rect -943 6533 -768 6550
rect -943 6493 -768 6510
rect -943 6453 -768 6470
rect -943 6413 -768 6430
rect -943 6373 -768 6390
rect -943 6333 -768 6350
rect -943 6293 -768 6310
rect -943 6253 -768 6270
rect -943 6213 -768 6230
rect -943 6173 -768 6190
rect -943 6133 -768 6150
rect -943 6093 -768 6110
rect -943 6053 -768 6070
rect -943 6013 -768 6030
rect -943 5973 -768 5990
rect -943 5933 -768 5950
rect -943 5893 -768 5910
rect -943 5853 -768 5870
rect -943 5813 -768 5830
rect -943 5773 -768 5790
rect -943 5733 -768 5750
rect -943 5693 -768 5710
rect -943 5653 -768 5670
rect -943 5613 -768 5630
rect -943 5573 -768 5590
rect -943 5533 -768 5550
rect -943 5493 -768 5510
rect -943 5453 -768 5470
rect -943 5413 -768 5430
rect -943 5373 -768 5390
rect -943 5333 -768 5350
rect -943 5293 -768 5310
rect -943 5253 -768 5270
rect -943 5213 -768 5230
rect -943 5173 -768 5190
rect -943 5133 -768 5150
rect -943 5093 -768 5110
rect -943 5053 -768 5070
rect -943 5013 -768 5030
rect -943 4973 -768 4990
rect -943 4933 -768 4950
rect -943 4893 -768 4910
rect -943 4853 -768 4870
rect -943 4813 -768 4830
rect -943 4773 -768 4790
rect -943 4733 -768 4750
rect -943 4693 -768 4710
rect -943 4653 -768 4670
rect -943 4613 -768 4630
rect -943 4573 -768 4590
rect -943 4533 -768 4550
rect -943 4493 -768 4510
rect -943 4453 -768 4470
rect -943 4413 -768 4430
rect -943 4373 -768 4390
rect -943 4333 -768 4350
rect -943 4293 -768 4310
rect -943 4253 -768 4270
rect -943 4213 -768 4230
rect -943 4173 -768 4190
rect -943 4133 -768 4150
rect -943 4093 -768 4110
rect -943 4053 -768 4070
rect -943 4013 -768 4030
rect -943 3973 -768 3990
rect -943 3933 -768 3950
rect -943 3893 -768 3910
rect -943 3853 -768 3870
rect -943 3813 -768 3830
rect -943 3773 -768 3790
rect -943 3733 -768 3750
rect -943 3693 -768 3710
rect -943 3653 -768 3670
rect -943 3613 -768 3630
rect -943 3573 -768 3590
rect -943 3533 -768 3550
rect -943 3493 -768 3510
rect -943 3453 -768 3470
rect -943 3413 -768 3430
rect -943 3373 -768 3390
rect -943 3333 -768 3350
rect -943 3293 -768 3310
rect -943 3253 -768 3270
rect -943 3213 -768 3230
rect -943 3173 -768 3190
rect -943 3133 -768 3150
rect -943 3093 -768 3110
rect -943 3053 -768 3070
rect -943 3013 -768 3030
rect -943 2973 -768 2990
rect -943 2933 -768 2950
rect -943 2893 -768 2910
rect -943 2853 -768 2870
rect -943 2813 -768 2830
rect -943 2773 -768 2790
rect -943 2733 -768 2750
rect -943 2693 -768 2710
rect -943 2653 -768 2670
rect -943 2613 -768 2630
rect -943 2573 -768 2590
rect -943 2533 -768 2550
rect -943 2493 -768 2510
rect -943 2453 -768 2470
rect -943 2413 -768 2430
rect -943 2373 -768 2390
rect -943 2333 -768 2350
rect -943 2293 -768 2310
rect -943 2253 -768 2270
rect -943 2213 -768 2230
rect -943 2173 -768 2190
rect -943 2133 -768 2150
rect -943 2093 -768 2110
rect -943 2053 -768 2070
rect -943 2013 -768 2030
rect -943 1973 -768 1990
rect -943 1933 -768 1950
rect -943 1893 -768 1910
rect -943 1853 -768 1870
rect -943 1813 -768 1830
rect -943 1773 -768 1790
rect -943 1733 -768 1750
rect -943 1693 -768 1710
rect -943 1653 -768 1670
rect -943 1613 -768 1630
rect -943 1573 -768 1590
rect -943 1533 -768 1550
rect -943 1493 -768 1510
rect -943 1453 -768 1470
rect -943 1413 -768 1430
rect -943 1373 -768 1390
rect -943 1333 -768 1350
rect -943 1293 -768 1310
rect -943 1253 -768 1270
rect -943 1213 -768 1230
rect -943 1173 -768 1190
rect -943 1133 -768 1150
rect -943 1093 -768 1110
rect -943 1053 -768 1070
rect -943 1013 -768 1030
rect -943 973 -768 990
rect -943 933 -768 950
rect -943 893 -768 910
rect -943 853 -768 870
rect 17650 9093 17825 9110
rect 17650 9053 17825 9070
rect 17650 9013 17825 9030
rect 17650 8973 17825 8990
rect 17650 8933 17825 8950
rect 17650 8893 17825 8910
rect 17650 8853 17825 8870
rect 17650 8813 17825 8830
rect 17650 8773 17825 8790
rect 17650 8733 17825 8750
rect 17650 8693 17825 8710
rect 17650 8653 17825 8670
rect 17650 8613 17825 8630
rect 17650 8573 17825 8590
rect 17650 8533 17825 8550
rect 17650 8493 17825 8510
rect 17650 8453 17825 8470
rect 17650 8413 17825 8430
rect 17650 8373 17825 8390
rect 17650 8333 17825 8350
rect 17650 8293 17825 8310
rect 17650 8253 17825 8270
rect 17650 8213 17825 8230
rect 17650 8173 17825 8190
rect 17650 8133 17825 8150
rect 17650 8093 17825 8110
rect 17650 8053 17825 8070
rect 17650 8013 17825 8030
rect 17650 7973 17825 7990
rect 17650 7933 17825 7950
rect 17650 7893 17825 7910
rect 17650 7853 17825 7870
rect 17650 7813 17825 7830
rect 17650 7773 17825 7790
rect 17650 7733 17825 7750
rect 17650 7693 17825 7710
rect 17650 7653 17825 7670
rect 17650 7613 17825 7630
rect 17650 7573 17825 7590
rect 17650 7533 17825 7550
rect 17650 7493 17825 7510
rect 17650 7453 17825 7470
rect 17650 7413 17825 7430
rect 17650 7373 17825 7390
rect 17650 7333 17825 7350
rect 17650 7293 17825 7310
rect 17650 7253 17825 7270
rect 17650 7213 17825 7230
rect 17650 7173 17825 7190
rect 17650 7133 17825 7150
rect 17650 7093 17825 7110
rect 17650 7053 17825 7070
rect 17650 7013 17825 7030
rect 17650 6973 17825 6990
rect 17650 6933 17825 6950
rect 17650 6893 17825 6910
rect 17650 6853 17825 6870
rect 17650 6813 17825 6830
rect 17650 6773 17825 6790
rect 17650 6733 17825 6750
rect 17650 6693 17825 6710
rect 17650 6653 17825 6670
rect 17650 6613 17825 6630
rect 17650 6573 17825 6590
rect 17650 6533 17825 6550
rect 17650 6493 17825 6510
rect 17650 6453 17825 6470
rect 17650 6413 17825 6430
rect 17650 6373 17825 6390
rect 17650 6333 17825 6350
rect 17650 6293 17825 6310
rect 17650 6253 17825 6270
rect 17651 6212 17826 6229
rect 17650 6173 17825 6190
rect 17650 6133 17825 6150
rect 17650 6093 17825 6110
rect 17650 6053 17825 6070
rect 17650 6013 17825 6030
rect 17650 5973 17825 5990
rect 17650 5933 17825 5950
rect 17650 5893 17825 5910
rect 17650 5853 17825 5870
rect 17650 5813 17825 5830
rect 17650 5773 17825 5790
rect 17650 5733 17825 5750
rect 17650 5693 17825 5710
rect 17650 5653 17825 5670
rect 17650 5613 17825 5630
rect 17650 5573 17825 5590
rect 17650 5533 17825 5550
rect 17650 5493 17825 5510
rect 17650 5453 17825 5470
rect 17650 5413 17825 5430
rect 17650 5373 17825 5390
rect 17649 5332 17824 5349
rect 17650 5293 17825 5310
rect 17650 5253 17825 5270
rect 17650 5213 17825 5230
rect 17650 5173 17825 5190
rect 17650 5133 17825 5150
rect 17650 5093 17825 5110
rect 17650 5053 17825 5070
rect 17650 5013 17825 5030
rect 17650 4973 17825 4990
rect 17650 4933 17825 4950
rect 17650 4893 17825 4910
rect 17650 4853 17825 4870
rect 17650 4813 17825 4830
rect 17650 4773 17825 4790
rect 17650 4733 17825 4750
rect 17650 4693 17825 4710
rect 17650 4653 17825 4670
rect 17650 4613 17825 4630
rect 17650 4573 17825 4590
rect 17650 4533 17825 4550
rect 17650 4493 17825 4510
rect 17650 4453 17825 4470
rect 17650 4413 17825 4430
rect 17650 4373 17825 4390
rect 17650 4333 17825 4350
rect 17650 4293 17825 4310
rect 17650 4253 17825 4270
rect 17650 4213 17825 4230
rect 17650 4173 17825 4190
rect 17650 4133 17825 4150
rect 17650 4093 17825 4110
rect 17650 4053 17825 4070
rect 17650 4013 17825 4030
rect 17650 3973 17825 3990
rect 17650 3933 17825 3950
rect 17650 3893 17825 3910
rect 17650 3853 17825 3870
rect 17650 3813 17825 3830
rect 17650 3773 17825 3790
rect 17650 3733 17825 3750
rect 17650 3693 17825 3710
rect 17650 3653 17825 3670
rect 17650 3613 17825 3630
rect 17650 3573 17825 3590
rect 17650 3533 17825 3550
rect 17650 3493 17825 3510
rect 17650 3453 17825 3470
rect 17650 3413 17825 3430
rect 17650 3373 17825 3390
rect 17650 3333 17825 3350
rect 17650 3293 17825 3310
rect 17650 3253 17825 3270
rect 17650 3213 17825 3230
rect 17650 3173 17825 3190
rect 17650 3133 17825 3150
rect 17650 3093 17825 3110
rect 17650 3053 17825 3070
rect 17650 3013 17825 3030
rect 17650 2973 17825 2990
rect 17650 2933 17825 2950
rect 17650 2893 17825 2910
rect 17650 2853 17825 2870
rect 17650 2813 17825 2830
rect 17650 2773 17825 2790
rect 17650 2733 17825 2750
rect 17650 2693 17825 2710
rect 17650 2653 17825 2670
rect 17650 2613 17825 2630
rect 17650 2573 17825 2590
rect 17650 2533 17825 2550
rect 17650 2493 17825 2510
rect 17650 2453 17825 2470
rect 17650 2413 17825 2430
rect 17650 2373 17825 2390
rect 17650 2333 17825 2350
rect 17650 2293 17825 2310
rect 17650 2250 17825 2267
rect 17650 2213 17825 2230
rect 17650 2173 17825 2190
rect 17650 2133 17825 2150
rect 17650 2093 17825 2110
rect 17650 2053 17825 2070
rect 17650 2013 17825 2030
rect 17650 1973 17825 1990
rect 17650 1933 17825 1950
rect 17650 1893 17825 1910
rect 17650 1853 17825 1870
rect 17650 1813 17825 1830
rect 17650 1773 17825 1790
rect 17650 1733 17825 1750
rect 17650 1693 17825 1710
rect 17650 1653 17825 1670
rect 17650 1613 17825 1630
rect 17650 1573 17825 1590
rect 17650 1533 17825 1550
rect 17650 1493 17825 1510
rect 17650 1453 17825 1470
rect 17650 1413 17825 1430
rect 17650 1373 17825 1390
rect 17650 1333 17825 1350
rect 17650 1293 17825 1310
rect 17650 1253 17825 1270
rect 17650 1213 17825 1230
rect 17650 1173 17825 1190
rect 17650 1133 17825 1150
rect 17650 1093 17825 1110
rect 17650 1053 17825 1070
rect 17650 1013 17825 1030
rect 17650 973 17825 990
rect 17650 933 17825 950
rect 17650 893 17825 910
rect 17650 853 17825 870
rect -943 813 -768 830
rect -943 773 -768 790
rect -943 733 -768 750
rect -943 693 -768 710
rect 17650 813 17825 830
rect 17650 773 17825 790
rect 17650 733 17825 750
rect 17650 693 17825 710
rect -943 653 -768 670
rect -943 613 -768 630
rect -943 573 -768 590
rect -943 533 -768 550
rect -943 493 -768 510
rect -943 453 -768 470
rect -943 413 -768 430
rect -943 373 -768 390
rect -943 333 -768 350
rect -943 293 -768 310
rect -943 253 -768 270
rect -943 213 -768 230
rect -943 173 -768 190
rect -943 133 -768 150
rect -943 93 -768 110
rect -943 53 -768 70
rect -943 13 -768 30
rect 17650 653 17825 670
rect 17650 613 17825 630
rect 17650 573 17825 590
rect 17650 533 17825 550
rect 17650 493 17825 510
rect 17650 453 17825 470
rect 17650 413 17825 430
rect 17650 373 17825 390
rect 17650 333 17825 350
rect 17650 293 17825 310
rect 17650 253 17825 270
rect 17650 213 17825 230
rect 17650 173 17825 190
rect 17650 133 17825 150
rect 17650 93 17825 110
rect 17650 53 17825 70
rect 17650 13 17825 30
<< locali >>
rect 20151 11168 20567 11181
rect 20151 10962 20448 11168
rect 20554 10962 20567 11168
rect 20151 10950 20567 10962
rect 20151 10289 20567 10302
rect 20151 10083 20448 10289
rect 20554 10083 20567 10289
rect 20151 10071 20567 10083
rect 292 9595 438 9603
rect 292 9516 299 9595
rect 430 9516 438 9595
rect -1195 -436 -988 9493
rect -440 9483 -294 9514
rect -440 9455 -430 9483
rect -402 9455 -383 9483
rect -355 9455 -336 9483
rect -308 9455 -294 9483
rect -440 9436 -294 9455
rect -440 9408 -430 9436
rect -402 9408 -383 9436
rect -355 9408 -336 9436
rect -308 9408 -294 9436
rect -440 9389 -294 9408
rect -440 9361 -430 9389
rect -402 9361 -383 9389
rect -355 9361 -336 9389
rect -308 9361 -294 9389
rect -957 9110 -750 9274
rect -957 9093 -943 9110
rect -768 9093 -750 9110
rect -957 9070 -750 9093
rect -957 9053 -943 9070
rect -768 9053 -750 9070
rect -957 9030 -750 9053
rect -957 9013 -943 9030
rect -768 9013 -750 9030
rect -957 8990 -750 9013
rect -957 8973 -943 8990
rect -768 8973 -750 8990
rect -957 8950 -750 8973
rect -957 8933 -943 8950
rect -768 8933 -750 8950
rect -957 8910 -750 8933
rect -957 8893 -943 8910
rect -768 8893 -750 8910
rect -957 8870 -750 8893
rect -957 8853 -943 8870
rect -768 8853 -750 8870
rect -957 8830 -750 8853
rect -957 8813 -943 8830
rect -768 8813 -750 8830
rect -957 8790 -750 8813
rect -957 8773 -943 8790
rect -768 8773 -750 8790
rect -957 8750 -750 8773
rect -957 8733 -943 8750
rect -768 8733 -750 8750
rect -957 8710 -750 8733
rect -957 8693 -943 8710
rect -768 8693 -750 8710
rect -957 8670 -750 8693
rect -957 8653 -943 8670
rect -768 8653 -750 8670
rect -957 8630 -750 8653
rect -957 8613 -943 8630
rect -768 8613 -750 8630
rect -957 8590 -750 8613
rect -957 8573 -943 8590
rect -768 8573 -750 8590
rect -957 8550 -750 8573
rect -957 8533 -943 8550
rect -768 8533 -750 8550
rect -957 8510 -750 8533
rect -957 8493 -943 8510
rect -768 8493 -750 8510
rect -957 8470 -750 8493
rect -957 8453 -943 8470
rect -768 8453 -750 8470
rect -957 8430 -750 8453
rect -957 8413 -943 8430
rect -768 8413 -750 8430
rect -957 8390 -750 8413
rect -957 8373 -943 8390
rect -768 8373 -750 8390
rect -957 8350 -750 8373
rect -957 8333 -943 8350
rect -768 8333 -750 8350
rect -957 8310 -750 8333
rect -957 8293 -943 8310
rect -768 8293 -750 8310
rect -957 8270 -750 8293
rect -957 8253 -943 8270
rect -768 8253 -750 8270
rect -957 8230 -750 8253
rect -957 8213 -943 8230
rect -768 8213 -750 8230
rect -957 8190 -750 8213
rect -957 8173 -943 8190
rect -768 8173 -750 8190
rect -957 8150 -750 8173
rect -957 8133 -943 8150
rect -768 8133 -750 8150
rect -957 8110 -750 8133
rect -957 8093 -943 8110
rect -768 8093 -750 8110
rect -957 8070 -750 8093
rect -957 8053 -943 8070
rect -768 8053 -750 8070
rect -957 8030 -750 8053
rect -957 8013 -943 8030
rect -768 8013 -750 8030
rect -957 7990 -750 8013
rect -957 7973 -943 7990
rect -768 7973 -750 7990
rect -957 7950 -750 7973
rect -957 7933 -943 7950
rect -768 7933 -750 7950
rect -957 7910 -750 7933
rect -957 7893 -943 7910
rect -768 7893 -750 7910
rect -957 7870 -750 7893
rect -957 7853 -943 7870
rect -768 7853 -750 7870
rect -957 7830 -750 7853
rect -957 7813 -943 7830
rect -768 7813 -750 7830
rect -957 7790 -750 7813
rect -957 7773 -943 7790
rect -768 7773 -750 7790
rect -957 7750 -750 7773
rect -957 7733 -943 7750
rect -768 7733 -750 7750
rect -957 7710 -750 7733
rect -957 7693 -943 7710
rect -768 7693 -750 7710
rect -957 7670 -750 7693
rect -957 7653 -943 7670
rect -768 7653 -750 7670
rect -957 7630 -750 7653
rect -957 7613 -943 7630
rect -768 7613 -750 7630
rect -957 7590 -750 7613
rect -957 7573 -943 7590
rect -768 7573 -750 7590
rect -957 7550 -750 7573
rect -957 7533 -943 7550
rect -768 7533 -750 7550
rect -957 7510 -750 7533
rect -957 7493 -943 7510
rect -768 7493 -750 7510
rect -957 7470 -750 7493
rect -957 7453 -943 7470
rect -768 7453 -750 7470
rect -957 7430 -750 7453
rect -957 7413 -943 7430
rect -768 7413 -750 7430
rect -957 7390 -750 7413
rect -957 7373 -943 7390
rect -768 7373 -750 7390
rect -957 7350 -750 7373
rect -957 7333 -943 7350
rect -768 7333 -750 7350
rect -957 7310 -750 7333
rect -957 7293 -943 7310
rect -768 7293 -750 7310
rect -957 7270 -750 7293
rect -957 7253 -943 7270
rect -768 7253 -750 7270
rect -957 7230 -750 7253
rect -957 7213 -943 7230
rect -768 7213 -750 7230
rect -957 7190 -750 7213
rect -957 7173 -943 7190
rect -768 7173 -750 7190
rect -957 7150 -750 7173
rect -957 7133 -943 7150
rect -768 7133 -750 7150
rect -957 7110 -750 7133
rect -957 7093 -943 7110
rect -768 7093 -750 7110
rect -957 7070 -750 7093
rect -957 7053 -943 7070
rect -768 7053 -750 7070
rect -957 7030 -750 7053
rect -957 7013 -943 7030
rect -768 7013 -750 7030
rect -957 6990 -750 7013
rect -957 6973 -943 6990
rect -768 6973 -750 6990
rect -957 6950 -750 6973
rect -957 6933 -943 6950
rect -768 6933 -750 6950
rect -957 6910 -750 6933
rect -957 6893 -943 6910
rect -768 6893 -750 6910
rect -957 6870 -750 6893
rect -957 6853 -943 6870
rect -768 6853 -750 6870
rect -957 6830 -750 6853
rect -957 6813 -943 6830
rect -768 6813 -750 6830
rect -957 6790 -750 6813
rect -957 6773 -943 6790
rect -768 6773 -750 6790
rect -957 6750 -750 6773
rect -957 6733 -943 6750
rect -768 6733 -750 6750
rect -957 6710 -750 6733
rect -957 6693 -943 6710
rect -768 6693 -750 6710
rect -957 6670 -750 6693
rect -957 6653 -943 6670
rect -768 6653 -750 6670
rect -957 6630 -750 6653
rect -957 6613 -943 6630
rect -768 6613 -750 6630
rect -957 6590 -750 6613
rect -957 6573 -943 6590
rect -768 6573 -750 6590
rect -957 6550 -750 6573
rect -957 6533 -943 6550
rect -768 6533 -750 6550
rect -957 6510 -750 6533
rect -957 6493 -943 6510
rect -768 6493 -750 6510
rect -957 6470 -750 6493
rect -957 6453 -943 6470
rect -768 6453 -750 6470
rect -957 6430 -750 6453
rect -957 6413 -943 6430
rect -768 6413 -750 6430
rect -957 6390 -750 6413
rect -957 6373 -943 6390
rect -768 6373 -750 6390
rect -957 6350 -750 6373
rect -957 6333 -943 6350
rect -768 6333 -750 6350
rect -957 6310 -750 6333
rect -957 6293 -943 6310
rect -768 6293 -750 6310
rect -957 6270 -750 6293
rect -957 6253 -943 6270
rect -768 6253 -750 6270
rect -957 6230 -750 6253
rect -957 6213 -943 6230
rect -768 6213 -750 6230
rect -957 6190 -750 6213
rect -957 6173 -943 6190
rect -768 6173 -750 6190
rect -957 6150 -750 6173
rect -957 6133 -943 6150
rect -768 6133 -750 6150
rect -957 6110 -750 6133
rect -957 6093 -943 6110
rect -768 6093 -750 6110
rect -957 6070 -750 6093
rect -957 6053 -943 6070
rect -768 6053 -750 6070
rect -957 6030 -750 6053
rect -957 6013 -943 6030
rect -768 6013 -750 6030
rect -957 5990 -750 6013
rect -957 5973 -943 5990
rect -768 5973 -750 5990
rect -957 5950 -750 5973
rect -957 5933 -943 5950
rect -768 5933 -750 5950
rect -957 5910 -750 5933
rect -957 5893 -943 5910
rect -768 5893 -750 5910
rect -957 5870 -750 5893
rect -957 5853 -943 5870
rect -768 5853 -750 5870
rect -957 5830 -750 5853
rect -957 5813 -943 5830
rect -768 5813 -750 5830
rect -957 5790 -750 5813
rect -957 5773 -943 5790
rect -768 5773 -750 5790
rect -957 5750 -750 5773
rect -957 5733 -943 5750
rect -768 5733 -750 5750
rect -957 5710 -750 5733
rect -957 5693 -943 5710
rect -768 5693 -750 5710
rect -957 5670 -750 5693
rect -957 5653 -943 5670
rect -768 5653 -750 5670
rect -957 5630 -750 5653
rect -957 5613 -943 5630
rect -768 5613 -750 5630
rect -957 5590 -750 5613
rect -957 5573 -943 5590
rect -768 5573 -750 5590
rect -957 5550 -750 5573
rect -957 5533 -943 5550
rect -768 5533 -750 5550
rect -957 5510 -750 5533
rect -957 5493 -943 5510
rect -768 5493 -750 5510
rect -957 5470 -750 5493
rect -957 5453 -943 5470
rect -768 5453 -750 5470
rect -957 5430 -750 5453
rect -957 5413 -943 5430
rect -768 5413 -750 5430
rect -957 5390 -750 5413
rect -957 5373 -943 5390
rect -768 5373 -750 5390
rect -957 5350 -750 5373
rect -957 5333 -943 5350
rect -768 5333 -750 5350
rect -957 5310 -750 5333
rect -957 5293 -943 5310
rect -768 5293 -750 5310
rect -957 5270 -750 5293
rect -957 5253 -943 5270
rect -768 5253 -750 5270
rect -957 5230 -750 5253
rect -957 5213 -943 5230
rect -768 5213 -750 5230
rect -957 5190 -750 5213
rect -957 5173 -943 5190
rect -768 5173 -750 5190
rect -957 5150 -750 5173
rect -957 5133 -943 5150
rect -768 5133 -750 5150
rect -957 5110 -750 5133
rect -957 5093 -943 5110
rect -768 5093 -750 5110
rect -957 5070 -750 5093
rect -957 5053 -943 5070
rect -768 5053 -750 5070
rect -957 5030 -750 5053
rect -957 5013 -943 5030
rect -768 5013 -750 5030
rect -957 4990 -750 5013
rect -957 4973 -943 4990
rect -768 4973 -750 4990
rect -957 4950 -750 4973
rect -957 4933 -943 4950
rect -768 4933 -750 4950
rect -957 4910 -750 4933
rect -957 4893 -943 4910
rect -768 4893 -750 4910
rect -957 4870 -750 4893
rect -957 4853 -943 4870
rect -768 4853 -750 4870
rect -957 4830 -750 4853
rect -957 4813 -943 4830
rect -768 4813 -750 4830
rect -957 4790 -750 4813
rect -957 4773 -943 4790
rect -768 4773 -750 4790
rect -957 4750 -750 4773
rect -957 4733 -943 4750
rect -768 4733 -750 4750
rect -957 4710 -750 4733
rect -957 4693 -943 4710
rect -768 4693 -750 4710
rect -957 4670 -750 4693
rect -957 4653 -943 4670
rect -768 4653 -750 4670
rect -957 4630 -750 4653
rect -957 4613 -943 4630
rect -768 4613 -750 4630
rect -957 4590 -750 4613
rect -957 4573 -943 4590
rect -768 4573 -750 4590
rect -957 4550 -750 4573
rect -957 4533 -943 4550
rect -768 4533 -750 4550
rect -957 4510 -750 4533
rect -957 4493 -943 4510
rect -768 4493 -750 4510
rect -957 4470 -750 4493
rect -957 4453 -943 4470
rect -768 4453 -750 4470
rect -957 4430 -750 4453
rect -957 4413 -943 4430
rect -768 4413 -750 4430
rect -957 4390 -750 4413
rect -957 4373 -943 4390
rect -768 4373 -750 4390
rect -957 4350 -750 4373
rect -957 4333 -943 4350
rect -768 4333 -750 4350
rect -957 4310 -750 4333
rect -957 4293 -943 4310
rect -768 4293 -750 4310
rect -957 4270 -750 4293
rect -957 4253 -943 4270
rect -768 4253 -750 4270
rect -957 4230 -750 4253
rect -957 4213 -943 4230
rect -768 4213 -750 4230
rect -957 4190 -750 4213
rect -957 4173 -943 4190
rect -768 4173 -750 4190
rect -957 4150 -750 4173
rect -957 4133 -943 4150
rect -768 4133 -750 4150
rect -957 4110 -750 4133
rect -957 4093 -943 4110
rect -768 4093 -750 4110
rect -957 4070 -750 4093
rect -957 4053 -943 4070
rect -768 4053 -750 4070
rect -957 4030 -750 4053
rect -957 4013 -943 4030
rect -768 4013 -750 4030
rect -957 3990 -750 4013
rect -957 3973 -943 3990
rect -768 3973 -750 3990
rect -957 3950 -750 3973
rect -957 3933 -943 3950
rect -768 3933 -750 3950
rect -957 3910 -750 3933
rect -957 3893 -943 3910
rect -768 3893 -750 3910
rect -957 3870 -750 3893
rect -957 3853 -943 3870
rect -768 3853 -750 3870
rect -957 3830 -750 3853
rect -957 3813 -943 3830
rect -768 3813 -750 3830
rect -957 3790 -750 3813
rect -957 3773 -943 3790
rect -768 3773 -750 3790
rect -957 3750 -750 3773
rect -957 3733 -943 3750
rect -768 3733 -750 3750
rect -957 3710 -750 3733
rect -957 3693 -943 3710
rect -768 3693 -750 3710
rect -957 3670 -750 3693
rect -957 3653 -943 3670
rect -768 3653 -750 3670
rect -957 3630 -750 3653
rect -957 3613 -943 3630
rect -768 3613 -750 3630
rect -957 3590 -750 3613
rect -957 3573 -943 3590
rect -768 3573 -750 3590
rect -957 3550 -750 3573
rect -957 3533 -943 3550
rect -768 3533 -750 3550
rect -957 3510 -750 3533
rect -957 3493 -943 3510
rect -768 3493 -750 3510
rect -957 3470 -750 3493
rect -957 3453 -943 3470
rect -768 3453 -750 3470
rect -957 3430 -750 3453
rect -957 3413 -943 3430
rect -768 3413 -750 3430
rect -957 3390 -750 3413
rect -957 3373 -943 3390
rect -768 3373 -750 3390
rect -957 3350 -750 3373
rect -957 3333 -943 3350
rect -768 3333 -750 3350
rect -957 3310 -750 3333
rect -957 3293 -943 3310
rect -768 3293 -750 3310
rect -957 3270 -750 3293
rect -957 3253 -943 3270
rect -768 3253 -750 3270
rect -957 3230 -750 3253
rect -957 3213 -943 3230
rect -768 3213 -750 3230
rect -957 3190 -750 3213
rect -957 3173 -943 3190
rect -768 3173 -750 3190
rect -957 3150 -750 3173
rect -957 3133 -943 3150
rect -768 3133 -750 3150
rect -957 3110 -750 3133
rect -957 3093 -943 3110
rect -768 3093 -750 3110
rect -957 3070 -750 3093
rect -957 3053 -943 3070
rect -768 3053 -750 3070
rect -957 3030 -750 3053
rect -957 3013 -943 3030
rect -768 3013 -750 3030
rect -957 2990 -750 3013
rect -957 2973 -943 2990
rect -768 2973 -750 2990
rect -957 2950 -750 2973
rect -957 2933 -943 2950
rect -768 2933 -750 2950
rect -957 2910 -750 2933
rect -957 2893 -943 2910
rect -768 2893 -750 2910
rect -957 2870 -750 2893
rect -957 2853 -943 2870
rect -768 2853 -750 2870
rect -957 2830 -750 2853
rect -957 2813 -943 2830
rect -768 2813 -750 2830
rect -957 2790 -750 2813
rect -957 2773 -943 2790
rect -768 2773 -750 2790
rect -957 2750 -750 2773
rect -957 2733 -943 2750
rect -768 2733 -750 2750
rect -957 2710 -750 2733
rect -957 2693 -943 2710
rect -768 2693 -750 2710
rect -957 2670 -750 2693
rect -957 2653 -943 2670
rect -768 2653 -750 2670
rect -957 2630 -750 2653
rect -957 2613 -943 2630
rect -768 2613 -750 2630
rect -957 2590 -750 2613
rect -957 2573 -943 2590
rect -768 2573 -750 2590
rect -957 2550 -750 2573
rect -957 2533 -943 2550
rect -768 2533 -750 2550
rect -957 2510 -750 2533
rect -957 2493 -943 2510
rect -768 2493 -750 2510
rect -957 2470 -750 2493
rect -957 2453 -943 2470
rect -768 2453 -750 2470
rect -957 2430 -750 2453
rect -957 2413 -943 2430
rect -768 2413 -750 2430
rect -957 2390 -750 2413
rect -957 2373 -943 2390
rect -768 2373 -750 2390
rect -957 2350 -750 2373
rect -957 2333 -943 2350
rect -768 2333 -750 2350
rect -957 2310 -750 2333
rect -957 2293 -943 2310
rect -768 2293 -750 2310
rect -957 2270 -750 2293
rect -957 2253 -943 2270
rect -768 2253 -750 2270
rect -957 2230 -750 2253
rect -957 2213 -943 2230
rect -768 2213 -750 2230
rect -957 2190 -750 2213
rect -957 2173 -943 2190
rect -768 2173 -750 2190
rect -957 2150 -750 2173
rect -957 2133 -943 2150
rect -768 2133 -750 2150
rect -957 2110 -750 2133
rect -957 2093 -943 2110
rect -768 2093 -750 2110
rect -957 2070 -750 2093
rect -957 2053 -943 2070
rect -768 2053 -750 2070
rect -957 2030 -750 2053
rect -957 2013 -943 2030
rect -768 2013 -750 2030
rect -957 1990 -750 2013
rect -957 1973 -943 1990
rect -768 1973 -750 1990
rect -957 1950 -750 1973
rect -957 1933 -943 1950
rect -768 1933 -750 1950
rect -957 1910 -750 1933
rect -957 1893 -943 1910
rect -768 1893 -750 1910
rect -957 1870 -750 1893
rect -957 1853 -943 1870
rect -768 1853 -750 1870
rect -957 1830 -750 1853
rect -957 1813 -943 1830
rect -768 1813 -750 1830
rect -957 1790 -750 1813
rect -957 1773 -943 1790
rect -768 1773 -750 1790
rect -957 1750 -750 1773
rect -957 1733 -943 1750
rect -768 1733 -750 1750
rect -957 1710 -750 1733
rect -957 1693 -943 1710
rect -768 1693 -750 1710
rect -957 1670 -750 1693
rect -957 1653 -943 1670
rect -768 1653 -750 1670
rect -957 1630 -750 1653
rect -957 1613 -943 1630
rect -768 1613 -750 1630
rect -957 1590 -750 1613
rect -957 1573 -943 1590
rect -768 1573 -750 1590
rect -957 1550 -750 1573
rect -957 1533 -943 1550
rect -768 1533 -750 1550
rect -957 1510 -750 1533
rect -957 1493 -943 1510
rect -768 1493 -750 1510
rect -957 1470 -750 1493
rect -957 1453 -943 1470
rect -768 1453 -750 1470
rect -957 1430 -750 1453
rect -957 1413 -943 1430
rect -768 1413 -750 1430
rect -957 1390 -750 1413
rect -957 1373 -943 1390
rect -768 1373 -750 1390
rect -957 1350 -750 1373
rect -957 1333 -943 1350
rect -768 1333 -750 1350
rect -957 1310 -750 1333
rect -957 1293 -943 1310
rect -768 1293 -750 1310
rect -957 1270 -750 1293
rect -957 1253 -943 1270
rect -768 1253 -750 1270
rect -957 1230 -750 1253
rect -957 1213 -943 1230
rect -768 1213 -750 1230
rect -957 1190 -750 1213
rect -957 1173 -943 1190
rect -768 1173 -750 1190
rect -957 1150 -750 1173
rect -957 1133 -943 1150
rect -768 1133 -750 1150
rect -957 1110 -750 1133
rect -957 1093 -943 1110
rect -768 1093 -750 1110
rect -957 1070 -750 1093
rect -957 1053 -943 1070
rect -768 1053 -750 1070
rect -957 1030 -750 1053
rect -957 1013 -943 1030
rect -768 1013 -750 1030
rect -957 990 -750 1013
rect -957 973 -943 990
rect -768 973 -750 990
rect -957 950 -750 973
rect -957 933 -943 950
rect -768 933 -750 950
rect -957 910 -750 933
rect -957 893 -943 910
rect -768 893 -750 910
rect -957 870 -750 893
rect -957 853 -943 870
rect -768 853 -750 870
rect -957 830 -750 853
rect -957 813 -943 830
rect -768 813 -750 830
rect -957 790 -750 813
rect -957 773 -943 790
rect -768 773 -750 790
rect -957 750 -750 773
rect -957 733 -943 750
rect -768 733 -750 750
rect -957 710 -750 733
rect -957 693 -943 710
rect -768 693 -750 710
rect -957 670 -750 693
rect -957 653 -943 670
rect -768 653 -750 670
rect -957 630 -750 653
rect -957 613 -943 630
rect -768 613 -750 630
rect -957 590 -750 613
rect -957 573 -943 590
rect -768 573 -750 590
rect -957 550 -750 573
rect -957 533 -943 550
rect -768 533 -750 550
rect -957 510 -750 533
rect -957 493 -943 510
rect -768 493 -750 510
rect -957 470 -750 493
rect -957 453 -943 470
rect -768 453 -750 470
rect -957 430 -750 453
rect -957 413 -943 430
rect -768 413 -750 430
rect -957 390 -750 413
rect -957 373 -943 390
rect -768 373 -750 390
rect -957 350 -750 373
rect -957 333 -943 350
rect -768 333 -750 350
rect -957 310 -750 333
rect -957 293 -943 310
rect -768 293 -750 310
rect -957 270 -750 293
rect -957 253 -943 270
rect -768 253 -750 270
rect -957 230 -750 253
rect -957 213 -943 230
rect -768 213 -750 230
rect -957 190 -750 213
rect -957 173 -943 190
rect -768 173 -750 190
rect -957 150 -750 173
rect -957 133 -943 150
rect -768 133 -750 150
rect -957 110 -750 133
rect -957 93 -943 110
rect -768 93 -750 110
rect -957 70 -750 93
rect -957 53 -943 70
rect -768 53 -750 70
rect -957 30 -750 53
rect -957 13 -943 30
rect -768 13 -750 30
rect -957 -217 -750 13
rect -659 8424 -625 9036
rect -659 8407 -651 8424
rect -634 8407 -625 8424
rect -659 7922 -625 8407
rect -659 7905 -651 7922
rect -634 7905 -625 7922
rect -659 7420 -625 7905
rect -659 7403 -651 7420
rect -634 7403 -625 7420
rect -659 6918 -625 7403
rect -659 6901 -651 6918
rect -634 6901 -625 6918
rect -659 6416 -625 6901
rect -659 6399 -651 6416
rect -634 6399 -625 6416
rect -659 5914 -625 6399
rect -659 5897 -651 5914
rect -634 5897 -625 5914
rect -659 5412 -625 5897
rect -659 5395 -651 5412
rect -634 5395 -625 5412
rect -659 4910 -625 5395
rect -659 4893 -651 4910
rect -634 4893 -625 4910
rect -659 4408 -625 4893
rect -659 4391 -651 4408
rect -634 4391 -625 4408
rect -659 3906 -625 4391
rect -659 3889 -651 3906
rect -634 3889 -625 3906
rect -659 3404 -625 3889
rect -659 3387 -651 3404
rect -634 3387 -625 3404
rect -659 2902 -625 3387
rect -659 2885 -651 2902
rect -634 2885 -625 2902
rect -659 2400 -625 2885
rect -659 2383 -651 2400
rect -634 2383 -625 2400
rect -659 1898 -625 2383
rect -659 1881 -651 1898
rect -634 1881 -625 1898
rect -659 1396 -625 1881
rect -659 1379 -651 1396
rect -634 1379 -625 1396
rect -659 894 -625 1379
rect -659 877 -651 894
rect -634 877 -625 894
rect -659 -457 -625 877
rect -605 8230 -571 9036
rect -605 8213 -597 8230
rect -580 8213 -571 8230
rect -605 7728 -571 8213
rect -605 7711 -597 7728
rect -580 7711 -571 7728
rect -605 7226 -571 7711
rect -605 7209 -597 7226
rect -580 7209 -571 7226
rect -605 6724 -571 7209
rect -605 6707 -597 6724
rect -580 6707 -571 6724
rect -605 6222 -571 6707
rect -605 6205 -597 6222
rect -580 6205 -571 6222
rect -605 5720 -571 6205
rect -605 5703 -597 5720
rect -580 5703 -571 5720
rect -605 5218 -571 5703
rect -605 5201 -597 5218
rect -580 5201 -571 5218
rect -605 4716 -571 5201
rect -605 4699 -597 4716
rect -580 4699 -571 4716
rect -605 4214 -571 4699
rect -605 4197 -597 4214
rect -580 4197 -571 4214
rect -605 3712 -571 4197
rect -605 3695 -597 3712
rect -580 3695 -571 3712
rect -605 3210 -571 3695
rect -605 3193 -597 3210
rect -580 3193 -571 3210
rect -605 2708 -571 3193
rect -605 2691 -597 2708
rect -580 2691 -571 2708
rect -605 2206 -571 2691
rect -605 2189 -597 2206
rect -580 2189 -571 2206
rect -605 1704 -571 2189
rect -605 1687 -597 1704
rect -580 1687 -571 1704
rect -605 1202 -571 1687
rect -605 1185 -597 1202
rect -580 1185 -571 1202
rect -605 700 -571 1185
rect -605 683 -597 700
rect -580 683 -571 700
rect -605 -457 -571 683
rect -551 8661 -483 9036
rect -551 8641 -545 8661
rect -525 8641 -506 8661
rect -486 8641 -483 8661
rect -551 8159 -483 8641
rect -551 8139 -545 8159
rect -525 8139 -506 8159
rect -486 8139 -483 8159
rect -551 7657 -483 8139
rect -551 7637 -545 7657
rect -525 7637 -506 7657
rect -486 7637 -483 7657
rect -551 7155 -483 7637
rect -551 7135 -545 7155
rect -525 7135 -506 7155
rect -486 7135 -483 7155
rect -551 6653 -483 7135
rect -551 6633 -545 6653
rect -525 6633 -506 6653
rect -486 6633 -483 6653
rect -551 6151 -483 6633
rect -551 6131 -545 6151
rect -525 6131 -506 6151
rect -486 6131 -483 6151
rect -551 5649 -483 6131
rect -551 5629 -545 5649
rect -525 5629 -506 5649
rect -486 5629 -483 5649
rect -551 5147 -483 5629
rect -551 5127 -545 5147
rect -525 5127 -506 5147
rect -486 5127 -483 5147
rect -551 4645 -483 5127
rect -551 4625 -545 4645
rect -525 4625 -506 4645
rect -486 4625 -483 4645
rect -551 4143 -483 4625
rect -551 4123 -545 4143
rect -525 4123 -506 4143
rect -486 4123 -483 4143
rect -551 3641 -483 4123
rect -551 3621 -545 3641
rect -525 3621 -506 3641
rect -486 3621 -483 3641
rect -551 3139 -483 3621
rect -551 3119 -545 3139
rect -525 3119 -506 3139
rect -486 3119 -483 3139
rect -551 2637 -483 3119
rect -551 2617 -545 2637
rect -525 2617 -506 2637
rect -486 2617 -483 2637
rect -551 2135 -483 2617
rect -551 2115 -545 2135
rect -525 2115 -506 2135
rect -486 2115 -483 2135
rect -551 1633 -483 2115
rect -551 1613 -545 1633
rect -525 1613 -506 1633
rect -486 1613 -483 1633
rect -551 1131 -483 1613
rect -551 1111 -545 1131
rect -525 1111 -506 1131
rect -486 1111 -483 1131
rect -551 629 -483 1111
rect -551 609 -545 629
rect -525 609 -506 629
rect -486 609 -483 629
rect -551 127 -483 609
rect -551 107 -545 127
rect -525 107 -506 127
rect -486 107 -483 127
rect -551 -457 -483 107
rect -440 8957 -294 9361
rect -440 8937 -434 8957
rect -414 8937 -395 8957
rect -375 8937 -356 8957
rect -336 8937 -317 8957
rect -297 8937 -294 8957
rect -440 8915 -294 8937
rect -440 8895 -434 8915
rect -414 8895 -395 8915
rect -375 8895 -356 8915
rect -336 8895 -317 8915
rect -297 8895 -294 8915
rect -440 8787 -294 8895
rect -440 8767 -434 8787
rect -414 8767 -395 8787
rect -375 8767 -356 8787
rect -336 8767 -317 8787
rect -297 8767 -294 8787
rect -440 8455 -294 8767
rect -440 8435 -434 8455
rect -414 8435 -395 8455
rect -375 8435 -356 8455
rect -336 8435 -317 8455
rect -297 8435 -294 8455
rect -440 7953 -294 8435
rect -440 7933 -434 7953
rect -414 7933 -395 7953
rect -375 7933 -356 7953
rect -336 7933 -317 7953
rect -297 7933 -294 7953
rect -440 7451 -294 7933
rect -440 7431 -434 7451
rect -414 7431 -395 7451
rect -375 7431 -356 7451
rect -336 7431 -317 7451
rect -297 7431 -294 7451
rect -440 6949 -294 7431
rect -440 6929 -434 6949
rect -414 6929 -395 6949
rect -375 6929 -356 6949
rect -336 6929 -317 6949
rect -297 6929 -294 6949
rect -440 6447 -294 6929
rect -440 6427 -434 6447
rect -414 6427 -395 6447
rect -375 6427 -356 6447
rect -336 6427 -317 6447
rect -297 6427 -294 6447
rect -440 5945 -294 6427
rect -440 5925 -434 5945
rect -414 5925 -395 5945
rect -375 5925 -356 5945
rect -336 5925 -317 5945
rect -297 5925 -294 5945
rect -440 5443 -294 5925
rect -440 5423 -434 5443
rect -414 5423 -395 5443
rect -375 5423 -356 5443
rect -336 5423 -317 5443
rect -297 5423 -294 5443
rect -440 4941 -294 5423
rect -440 4921 -434 4941
rect -414 4921 -395 4941
rect -375 4921 -356 4941
rect -336 4921 -317 4941
rect -297 4921 -294 4941
rect -440 4439 -294 4921
rect -440 4419 -434 4439
rect -414 4419 -395 4439
rect -375 4419 -356 4439
rect -336 4419 -317 4439
rect -297 4419 -294 4439
rect -440 3937 -294 4419
rect -440 3917 -434 3937
rect -414 3917 -395 3937
rect -375 3917 -356 3937
rect -336 3917 -317 3937
rect -297 3917 -294 3937
rect -440 3435 -294 3917
rect -440 3415 -434 3435
rect -414 3415 -395 3435
rect -375 3415 -356 3435
rect -336 3415 -317 3435
rect -297 3415 -294 3435
rect -440 2933 -294 3415
rect -440 2913 -434 2933
rect -414 2913 -395 2933
rect -375 2913 -356 2933
rect -336 2913 -317 2933
rect -297 2913 -294 2933
rect -440 2431 -294 2913
rect -440 2411 -434 2431
rect -414 2411 -395 2431
rect -375 2411 -356 2431
rect -336 2411 -317 2431
rect -297 2411 -294 2431
rect -440 1929 -294 2411
rect -440 1909 -434 1929
rect -414 1909 -395 1929
rect -375 1909 -356 1929
rect -336 1909 -317 1929
rect -297 1909 -294 1929
rect -440 1427 -294 1909
rect -440 1407 -434 1427
rect -414 1407 -395 1427
rect -375 1407 -356 1427
rect -336 1407 -317 1427
rect -297 1407 -294 1427
rect -440 925 -294 1407
rect -440 905 -434 925
rect -414 905 -395 925
rect -375 905 -356 925
rect -336 905 -317 925
rect -297 905 -294 925
rect -440 423 -294 905
rect -440 403 -434 423
rect -414 403 -395 423
rect -375 403 -356 423
rect -336 403 -317 423
rect -297 403 -294 423
rect -440 381 -294 403
rect -440 361 -434 381
rect -414 361 -395 381
rect -375 361 -356 381
rect -336 361 -317 381
rect -297 361 -294 381
rect -440 -304 -294 361
rect -440 -332 -430 -304
rect -402 -332 -383 -304
rect -355 -332 -336 -304
rect -308 -332 -294 -304
rect -440 -351 -294 -332
rect -440 -379 -430 -351
rect -402 -379 -383 -351
rect -355 -379 -336 -351
rect -308 -379 -294 -351
rect -440 -398 -294 -379
rect -440 -426 -430 -398
rect -402 -426 -383 -398
rect -355 -426 -336 -398
rect -308 -426 -294 -398
rect -440 -457 -294 -426
rect -251 9264 -105 9514
rect -251 9236 -241 9264
rect -213 9236 -194 9264
rect -166 9236 -147 9264
rect -119 9236 -105 9264
rect -251 9217 -105 9236
rect -251 9189 -241 9217
rect -213 9189 -194 9217
rect -166 9189 -147 9217
rect -119 9189 -105 9217
rect -251 9170 -105 9189
rect -251 9142 -241 9170
rect -213 9142 -194 9170
rect -166 9142 -147 9170
rect -119 9142 -105 9170
rect -251 8731 -105 9142
rect 292 9264 438 9516
rect 292 9236 302 9264
rect 330 9236 349 9264
rect 377 9236 396 9264
rect 424 9236 438 9264
rect 292 9217 438 9236
rect 292 9189 302 9217
rect 330 9189 349 9217
rect 377 9189 396 9217
rect 424 9189 438 9217
rect 292 9170 438 9189
rect 292 9142 302 9170
rect 330 9142 349 9170
rect 377 9142 396 9170
rect 424 9142 438 9170
rect 292 9134 438 9142
rect 642 9264 788 9626
rect 642 9236 652 9264
rect 680 9236 699 9264
rect 727 9236 746 9264
rect 774 9236 788 9264
rect 642 9217 788 9236
rect 642 9189 652 9217
rect 680 9189 699 9217
rect 727 9189 746 9217
rect 774 9189 788 9217
rect 642 9170 788 9189
rect 642 9142 652 9170
rect 680 9142 699 9170
rect 727 9142 746 9170
rect 774 9142 788 9170
rect 642 9134 788 9142
rect 1856 9595 2002 9603
rect 1856 9516 1863 9595
rect 1994 9516 2002 9595
rect 1856 9264 2002 9516
rect 1856 9236 1866 9264
rect 1894 9236 1913 9264
rect 1941 9236 1960 9264
rect 1988 9236 2002 9264
rect 1856 9217 2002 9236
rect 1856 9189 1866 9217
rect 1894 9189 1913 9217
rect 1941 9189 1960 9217
rect 1988 9189 2002 9217
rect 1856 9170 2002 9189
rect 1856 9142 1866 9170
rect 1894 9142 1913 9170
rect 1941 9142 1960 9170
rect 1988 9142 2002 9170
rect 1856 9134 2002 9142
rect 2292 9595 2438 9603
rect 2292 9516 2299 9595
rect 2430 9516 2438 9595
rect 2292 9264 2438 9516
rect 2292 9236 2302 9264
rect 2330 9236 2349 9264
rect 2377 9236 2396 9264
rect 2424 9236 2438 9264
rect 2292 9217 2438 9236
rect 2292 9189 2302 9217
rect 2330 9189 2349 9217
rect 2377 9189 2396 9217
rect 2424 9189 2438 9217
rect 2292 9170 2438 9189
rect 2292 9142 2302 9170
rect 2330 9142 2349 9170
rect 2377 9142 2396 9170
rect 2424 9142 2438 9170
rect 2292 9134 2438 9142
rect 2642 9264 2788 9626
rect 2642 9236 2652 9264
rect 2680 9236 2699 9264
rect 2727 9236 2746 9264
rect 2774 9236 2788 9264
rect 2642 9217 2788 9236
rect 2642 9189 2652 9217
rect 2680 9189 2699 9217
rect 2727 9189 2746 9217
rect 2774 9189 2788 9217
rect 2642 9170 2788 9189
rect 2642 9142 2652 9170
rect 2680 9142 2699 9170
rect 2727 9142 2746 9170
rect 2774 9142 2788 9170
rect 2642 9134 2788 9142
rect 3856 9595 4002 9603
rect 3856 9516 3863 9595
rect 3994 9516 4002 9595
rect 3856 9264 4002 9516
rect 3856 9236 3866 9264
rect 3894 9236 3913 9264
rect 3941 9236 3960 9264
rect 3988 9236 4002 9264
rect 3856 9217 4002 9236
rect 3856 9189 3866 9217
rect 3894 9189 3913 9217
rect 3941 9189 3960 9217
rect 3988 9189 4002 9217
rect 3856 9170 4002 9189
rect 3856 9142 3866 9170
rect 3894 9142 3913 9170
rect 3941 9142 3960 9170
rect 3988 9142 4002 9170
rect 3856 9134 4002 9142
rect 4292 9595 4438 9603
rect 4292 9516 4299 9595
rect 4430 9516 4438 9595
rect 4292 9264 4438 9516
rect 4292 9236 4302 9264
rect 4330 9236 4349 9264
rect 4377 9236 4396 9264
rect 4424 9236 4438 9264
rect 4292 9217 4438 9236
rect 4292 9189 4302 9217
rect 4330 9189 4349 9217
rect 4377 9189 4396 9217
rect 4424 9189 4438 9217
rect 4292 9170 4438 9189
rect 4292 9142 4302 9170
rect 4330 9142 4349 9170
rect 4377 9142 4396 9170
rect 4424 9142 4438 9170
rect 4292 9134 4438 9142
rect 4642 9264 4788 9626
rect 4642 9236 4652 9264
rect 4680 9236 4699 9264
rect 4727 9236 4746 9264
rect 4774 9236 4788 9264
rect 4642 9217 4788 9236
rect 4642 9189 4652 9217
rect 4680 9189 4699 9217
rect 4727 9189 4746 9217
rect 4774 9189 4788 9217
rect 4642 9170 4788 9189
rect 4642 9142 4652 9170
rect 4680 9142 4699 9170
rect 4727 9142 4746 9170
rect 4774 9142 4788 9170
rect 4642 9134 4788 9142
rect 5856 9595 6002 9603
rect 5856 9516 5863 9595
rect 5994 9516 6002 9595
rect 5856 9264 6002 9516
rect 5856 9236 5866 9264
rect 5894 9236 5913 9264
rect 5941 9236 5960 9264
rect 5988 9236 6002 9264
rect 5856 9217 6002 9236
rect 5856 9189 5866 9217
rect 5894 9189 5913 9217
rect 5941 9189 5960 9217
rect 5988 9189 6002 9217
rect 5856 9170 6002 9189
rect 5856 9142 5866 9170
rect 5894 9142 5913 9170
rect 5941 9142 5960 9170
rect 5988 9142 6002 9170
rect 5856 9134 6002 9142
rect 6292 9595 6438 9603
rect 6292 9516 6299 9595
rect 6430 9516 6438 9595
rect 6292 9264 6438 9516
rect 6292 9236 6302 9264
rect 6330 9236 6349 9264
rect 6377 9236 6396 9264
rect 6424 9236 6438 9264
rect 6292 9217 6438 9236
rect 6292 9189 6302 9217
rect 6330 9189 6349 9217
rect 6377 9189 6396 9217
rect 6424 9189 6438 9217
rect 6292 9170 6438 9189
rect 6292 9142 6302 9170
rect 6330 9142 6349 9170
rect 6377 9142 6396 9170
rect 6424 9142 6438 9170
rect 6292 9134 6438 9142
rect 6642 9264 6788 9626
rect 6642 9236 6652 9264
rect 6680 9236 6699 9264
rect 6727 9236 6746 9264
rect 6774 9236 6788 9264
rect 6642 9217 6788 9236
rect 6642 9189 6652 9217
rect 6680 9189 6699 9217
rect 6727 9189 6746 9217
rect 6774 9189 6788 9217
rect 6642 9170 6788 9189
rect 6642 9142 6652 9170
rect 6680 9142 6699 9170
rect 6727 9142 6746 9170
rect 6774 9142 6788 9170
rect 6642 9134 6788 9142
rect 7856 9595 8002 9603
rect 7856 9516 7863 9595
rect 7994 9516 8002 9595
rect 7856 9264 8002 9516
rect 7856 9236 7866 9264
rect 7894 9236 7913 9264
rect 7941 9236 7960 9264
rect 7988 9236 8002 9264
rect 7856 9217 8002 9236
rect 7856 9189 7866 9217
rect 7894 9189 7913 9217
rect 7941 9189 7960 9217
rect 7988 9189 8002 9217
rect 7856 9170 8002 9189
rect 7856 9142 7866 9170
rect 7894 9142 7913 9170
rect 7941 9142 7960 9170
rect 7988 9142 8002 9170
rect 7856 9134 8002 9142
rect 8292 9595 8438 9603
rect 8292 9516 8299 9595
rect 8430 9516 8438 9595
rect 8292 9264 8438 9516
rect 8292 9236 8302 9264
rect 8330 9236 8349 9264
rect 8377 9236 8396 9264
rect 8424 9236 8438 9264
rect 8292 9217 8438 9236
rect 8292 9189 8302 9217
rect 8330 9189 8349 9217
rect 8377 9189 8396 9217
rect 8424 9189 8438 9217
rect 8292 9170 8438 9189
rect 8292 9142 8302 9170
rect 8330 9142 8349 9170
rect 8377 9142 8396 9170
rect 8424 9142 8438 9170
rect 8292 9134 8438 9142
rect 8642 9264 8788 9626
rect 8642 9236 8652 9264
rect 8680 9236 8699 9264
rect 8727 9236 8746 9264
rect 8774 9236 8788 9264
rect 8642 9217 8788 9236
rect 8642 9189 8652 9217
rect 8680 9189 8699 9217
rect 8727 9189 8746 9217
rect 8774 9189 8788 9217
rect 8642 9170 8788 9189
rect 8642 9142 8652 9170
rect 8680 9142 8699 9170
rect 8727 9142 8746 9170
rect 8774 9142 8788 9170
rect 8642 9134 8788 9142
rect 9856 9595 10002 9603
rect 9856 9516 9863 9595
rect 9994 9516 10002 9595
rect 9856 9264 10002 9516
rect 9856 9236 9866 9264
rect 9894 9236 9913 9264
rect 9941 9236 9960 9264
rect 9988 9236 10002 9264
rect 9856 9217 10002 9236
rect 9856 9189 9866 9217
rect 9894 9189 9913 9217
rect 9941 9189 9960 9217
rect 9988 9189 10002 9217
rect 9856 9170 10002 9189
rect 9856 9142 9866 9170
rect 9894 9142 9913 9170
rect 9941 9142 9960 9170
rect 9988 9142 10002 9170
rect 9856 9134 10002 9142
rect 10292 9595 10438 9603
rect 10292 9516 10299 9595
rect 10430 9516 10438 9595
rect 10292 9264 10438 9516
rect 10292 9236 10302 9264
rect 10330 9236 10349 9264
rect 10377 9236 10396 9264
rect 10424 9236 10438 9264
rect 10292 9217 10438 9236
rect 10292 9189 10302 9217
rect 10330 9189 10349 9217
rect 10377 9189 10396 9217
rect 10424 9189 10438 9217
rect 10292 9170 10438 9189
rect 10292 9142 10302 9170
rect 10330 9142 10349 9170
rect 10377 9142 10396 9170
rect 10424 9142 10438 9170
rect 10292 9134 10438 9142
rect 10642 9264 10788 9626
rect 10642 9236 10652 9264
rect 10680 9236 10699 9264
rect 10727 9236 10746 9264
rect 10774 9236 10788 9264
rect 10642 9217 10788 9236
rect 10642 9189 10652 9217
rect 10680 9189 10699 9217
rect 10727 9189 10746 9217
rect 10774 9189 10788 9217
rect 10642 9170 10788 9189
rect 10642 9142 10652 9170
rect 10680 9142 10699 9170
rect 10727 9142 10746 9170
rect 10774 9142 10788 9170
rect 10642 9134 10788 9142
rect 11856 9595 12002 9603
rect 11856 9516 11863 9595
rect 11994 9516 12002 9595
rect 11856 9264 12002 9516
rect 11856 9236 11866 9264
rect 11894 9236 11913 9264
rect 11941 9236 11960 9264
rect 11988 9236 12002 9264
rect 11856 9217 12002 9236
rect 11856 9189 11866 9217
rect 11894 9189 11913 9217
rect 11941 9189 11960 9217
rect 11988 9189 12002 9217
rect 11856 9170 12002 9189
rect 11856 9142 11866 9170
rect 11894 9142 11913 9170
rect 11941 9142 11960 9170
rect 11988 9142 12002 9170
rect 11856 9134 12002 9142
rect 12292 9595 12438 9603
rect 12292 9516 12299 9595
rect 12430 9516 12438 9595
rect 12292 9264 12438 9516
rect 12292 9236 12302 9264
rect 12330 9236 12349 9264
rect 12377 9236 12396 9264
rect 12424 9236 12438 9264
rect 12292 9217 12438 9236
rect 12292 9189 12302 9217
rect 12330 9189 12349 9217
rect 12377 9189 12396 9217
rect 12424 9189 12438 9217
rect 12292 9170 12438 9189
rect 12292 9142 12302 9170
rect 12330 9142 12349 9170
rect 12377 9142 12396 9170
rect 12424 9142 12438 9170
rect 12292 9134 12438 9142
rect 12642 9264 12788 9626
rect 12642 9236 12652 9264
rect 12680 9236 12699 9264
rect 12727 9236 12746 9264
rect 12774 9236 12788 9264
rect 12642 9217 12788 9236
rect 12642 9189 12652 9217
rect 12680 9189 12699 9217
rect 12727 9189 12746 9217
rect 12774 9189 12788 9217
rect 12642 9170 12788 9189
rect 12642 9142 12652 9170
rect 12680 9142 12699 9170
rect 12727 9142 12746 9170
rect 12774 9142 12788 9170
rect 12642 9134 12788 9142
rect 13856 9595 14002 9603
rect 13856 9516 13863 9595
rect 13994 9516 14002 9595
rect 13856 9264 14002 9516
rect 13856 9236 13866 9264
rect 13894 9236 13913 9264
rect 13941 9236 13960 9264
rect 13988 9236 14002 9264
rect 13856 9217 14002 9236
rect 13856 9189 13866 9217
rect 13894 9189 13913 9217
rect 13941 9189 13960 9217
rect 13988 9189 14002 9217
rect 13856 9170 14002 9189
rect 13856 9142 13866 9170
rect 13894 9142 13913 9170
rect 13941 9142 13960 9170
rect 13988 9142 14002 9170
rect 13856 9134 14002 9142
rect 14292 9595 14438 9603
rect 14292 9516 14299 9595
rect 14430 9516 14438 9595
rect 14292 9264 14438 9516
rect 14292 9236 14302 9264
rect 14330 9236 14349 9264
rect 14377 9236 14396 9264
rect 14424 9236 14438 9264
rect 14292 9217 14438 9236
rect 14292 9189 14302 9217
rect 14330 9189 14349 9217
rect 14377 9189 14396 9217
rect 14424 9189 14438 9217
rect 14292 9170 14438 9189
rect 14292 9142 14302 9170
rect 14330 9142 14349 9170
rect 14377 9142 14396 9170
rect 14424 9142 14438 9170
rect 14292 9134 14438 9142
rect 14642 9264 14788 9626
rect 14642 9236 14652 9264
rect 14680 9236 14699 9264
rect 14727 9236 14746 9264
rect 14774 9236 14788 9264
rect 14642 9217 14788 9236
rect 14642 9189 14652 9217
rect 14680 9189 14699 9217
rect 14727 9189 14746 9217
rect 14774 9189 14788 9217
rect 14642 9170 14788 9189
rect 14642 9142 14652 9170
rect 14680 9142 14699 9170
rect 14727 9142 14746 9170
rect 14774 9142 14788 9170
rect 14642 9134 14788 9142
rect 15856 9595 16002 9603
rect 15856 9516 15863 9595
rect 15994 9516 16002 9595
rect 15856 9264 16002 9516
rect 15856 9236 15866 9264
rect 15894 9236 15913 9264
rect 15941 9236 15960 9264
rect 15988 9236 16002 9264
rect 15856 9217 16002 9236
rect 15856 9189 15866 9217
rect 15894 9189 15913 9217
rect 15941 9189 15960 9217
rect 15988 9189 16002 9217
rect 15856 9170 16002 9189
rect 15856 9142 15866 9170
rect 15894 9142 15913 9170
rect 15941 9142 15960 9170
rect 15988 9142 16002 9170
rect 15856 9134 16002 9142
rect 16292 9595 16438 9603
rect 16292 9516 16299 9595
rect 16430 9516 16438 9595
rect 16292 9264 16438 9516
rect 16292 9236 16302 9264
rect 16330 9236 16349 9264
rect 16377 9236 16396 9264
rect 16424 9236 16438 9264
rect 16292 9217 16438 9236
rect 16292 9189 16302 9217
rect 16330 9189 16349 9217
rect 16377 9189 16396 9217
rect 16424 9189 16438 9217
rect 16292 9170 16438 9189
rect 16292 9142 16302 9170
rect 16330 9142 16349 9170
rect 16377 9142 16396 9170
rect 16424 9142 16438 9170
rect 16292 9134 16438 9142
rect 16642 9264 16788 9626
rect 17856 9595 18002 9603
rect 17856 9533 17863 9595
rect 17994 9533 18002 9595
rect 16642 9236 16652 9264
rect 16680 9236 16699 9264
rect 16727 9236 16746 9264
rect 16774 9236 16788 9264
rect 16642 9217 16788 9236
rect 16642 9189 16652 9217
rect 16680 9189 16699 9217
rect 16727 9189 16746 9217
rect 16774 9189 16788 9217
rect 16642 9170 16788 9189
rect 16642 9142 16652 9170
rect 16680 9142 16699 9170
rect 16727 9142 16746 9170
rect 16774 9142 16788 9170
rect 16642 9134 16788 9142
rect 17167 9259 17315 9509
rect 17167 9231 17181 9259
rect 17209 9231 17228 9259
rect 17256 9231 17275 9259
rect 17303 9231 17315 9259
rect 17167 9212 17315 9231
rect 17167 9184 17181 9212
rect 17209 9184 17228 9212
rect 17256 9184 17275 9212
rect 17303 9184 17315 9212
rect 17167 9165 17315 9184
rect 17167 9137 17181 9165
rect 17209 9137 17228 9165
rect 17256 9137 17275 9165
rect 17303 9137 17315 9165
rect -251 8711 -245 8731
rect -225 8711 -206 8731
rect -186 8711 -167 8731
rect -147 8711 -128 8731
rect -108 8711 -105 8731
rect -251 8626 -105 8711
rect -251 8606 -245 8626
rect -225 8606 -206 8626
rect -186 8606 -167 8626
rect -147 8606 -128 8626
rect -108 8606 -105 8626
rect -251 8124 -105 8606
rect -251 8104 -245 8124
rect -225 8104 -206 8124
rect -186 8104 -167 8124
rect -147 8104 -128 8124
rect -108 8104 -105 8124
rect -251 7622 -105 8104
rect -251 7602 -245 7622
rect -225 7602 -206 7622
rect -186 7602 -167 7622
rect -147 7602 -128 7622
rect -108 7602 -105 7622
rect -251 7120 -105 7602
rect -251 7100 -245 7120
rect -225 7100 -206 7120
rect -186 7100 -167 7120
rect -147 7100 -128 7120
rect -108 7100 -105 7120
rect -251 6618 -105 7100
rect -251 6598 -245 6618
rect -225 6598 -206 6618
rect -186 6598 -167 6618
rect -147 6598 -128 6618
rect -108 6598 -105 6618
rect -251 6116 -105 6598
rect -251 6096 -245 6116
rect -225 6096 -206 6116
rect -186 6096 -167 6116
rect -147 6096 -128 6116
rect -108 6096 -105 6116
rect -251 5614 -105 6096
rect -251 5594 -245 5614
rect -225 5594 -206 5614
rect -186 5594 -167 5614
rect -147 5594 -128 5614
rect -108 5594 -105 5614
rect -251 5112 -105 5594
rect -251 5092 -245 5112
rect -225 5092 -206 5112
rect -186 5092 -167 5112
rect -147 5092 -128 5112
rect -108 5092 -105 5112
rect -251 4610 -105 5092
rect -251 4590 -245 4610
rect -225 4590 -206 4610
rect -186 4590 -167 4610
rect -147 4590 -128 4610
rect -108 4590 -105 4610
rect -251 4108 -105 4590
rect -251 4088 -245 4108
rect -225 4088 -206 4108
rect -186 4088 -167 4108
rect -147 4088 -128 4108
rect -108 4088 -105 4108
rect -251 3606 -105 4088
rect -251 3586 -245 3606
rect -225 3586 -206 3606
rect -186 3586 -167 3606
rect -147 3586 -128 3606
rect -108 3586 -105 3606
rect -251 3104 -105 3586
rect -251 3084 -245 3104
rect -225 3084 -206 3104
rect -186 3084 -167 3104
rect -147 3084 -128 3104
rect -108 3084 -105 3104
rect -251 2602 -105 3084
rect -251 2582 -245 2602
rect -225 2582 -206 2602
rect -186 2582 -167 2602
rect -147 2582 -128 2602
rect -108 2582 -105 2602
rect -251 2100 -105 2582
rect -251 2080 -245 2100
rect -225 2080 -206 2100
rect -186 2080 -167 2100
rect -147 2080 -128 2100
rect -108 2080 -105 2100
rect -251 1598 -105 2080
rect -251 1578 -245 1598
rect -225 1578 -206 1598
rect -186 1578 -167 1598
rect -147 1578 -128 1598
rect -108 1578 -105 1598
rect -251 1096 -105 1578
rect -251 1076 -245 1096
rect -225 1076 -206 1096
rect -186 1076 -167 1096
rect -147 1076 -128 1096
rect -108 1076 -105 1096
rect -251 594 -105 1076
rect 17167 8865 17315 9137
rect 17167 8837 17182 8865
rect 17210 8837 17229 8865
rect 17257 8837 17276 8865
rect 17304 8837 17315 8865
rect 17167 8818 17315 8837
rect 17167 8790 17182 8818
rect 17210 8790 17229 8818
rect 17257 8790 17276 8818
rect 17304 8790 17315 8818
rect 17167 8771 17315 8790
rect 17167 8743 17182 8771
rect 17210 8743 17229 8771
rect 17257 8743 17276 8771
rect 17304 8743 17315 8771
rect 17167 8626 17315 8743
rect 17167 8606 17170 8626
rect 17190 8606 17209 8626
rect 17229 8606 17248 8626
rect 17268 8606 17287 8626
rect 17307 8606 17315 8626
rect 17167 8124 17315 8606
rect 17167 8104 17170 8124
rect 17190 8104 17209 8124
rect 17229 8104 17248 8124
rect 17268 8104 17287 8124
rect 17307 8104 17315 8124
rect 17167 7857 17315 8104
rect 17167 7829 17181 7857
rect 17209 7829 17228 7857
rect 17256 7829 17275 7857
rect 17303 7829 17315 7857
rect 17167 7810 17315 7829
rect 17167 7782 17181 7810
rect 17209 7782 17228 7810
rect 17256 7782 17275 7810
rect 17303 7782 17315 7810
rect 17167 7763 17315 7782
rect 17167 7735 17181 7763
rect 17209 7735 17228 7763
rect 17256 7735 17275 7763
rect 17303 7735 17315 7763
rect 17167 7622 17315 7735
rect 17167 7602 17170 7622
rect 17190 7602 17209 7622
rect 17229 7602 17248 7622
rect 17268 7602 17287 7622
rect 17307 7602 17315 7622
rect 17167 7120 17315 7602
rect 17167 7100 17170 7120
rect 17190 7100 17209 7120
rect 17229 7100 17248 7120
rect 17268 7100 17287 7120
rect 17307 7100 17315 7120
rect 17167 6857 17315 7100
rect 17167 6829 17181 6857
rect 17209 6829 17228 6857
rect 17256 6829 17275 6857
rect 17303 6829 17315 6857
rect 17167 6810 17315 6829
rect 17167 6782 17181 6810
rect 17209 6782 17228 6810
rect 17256 6782 17275 6810
rect 17303 6782 17315 6810
rect 17167 6763 17315 6782
rect 17167 6735 17181 6763
rect 17209 6735 17228 6763
rect 17256 6735 17275 6763
rect 17303 6735 17315 6763
rect 17167 6618 17315 6735
rect 17167 6598 17170 6618
rect 17190 6598 17209 6618
rect 17229 6598 17248 6618
rect 17268 6598 17287 6618
rect 17307 6598 17315 6618
rect 17167 6116 17315 6598
rect 17355 9478 17502 9509
rect 17355 9450 17370 9478
rect 17398 9450 17417 9478
rect 17445 9450 17464 9478
rect 17492 9450 17502 9478
rect 17355 9431 17502 9450
rect 17355 9403 17370 9431
rect 17398 9403 17417 9431
rect 17445 9403 17464 9431
rect 17492 9403 17502 9431
rect 17355 9384 17502 9403
rect 17355 9356 17370 9384
rect 17398 9356 17417 9384
rect 17445 9356 17464 9384
rect 17492 9356 17502 9384
rect 17355 9036 17502 9356
rect 17856 9493 18002 9533
rect 17632 9110 17839 9274
rect 17856 9264 18077 9493
rect 17856 9236 17866 9264
rect 17894 9236 17913 9264
rect 17941 9236 17960 9264
rect 17988 9236 18077 9264
rect 17856 9217 18077 9236
rect 17856 9189 17866 9217
rect 17894 9189 17913 9217
rect 17941 9189 17960 9217
rect 17988 9189 18077 9217
rect 17856 9170 18077 9189
rect 17856 9142 17866 9170
rect 17894 9142 17913 9170
rect 17941 9142 17960 9170
rect 17988 9142 18077 9170
rect 17856 9134 18077 9142
rect 17632 9093 17650 9110
rect 17825 9093 17839 9110
rect 17632 9070 17839 9093
rect 17632 9053 17650 9070
rect 17825 9053 17839 9070
rect 17355 8957 17503 9036
rect 17355 8937 17359 8957
rect 17379 8937 17398 8957
rect 17418 8937 17437 8957
rect 17457 8937 17476 8957
rect 17496 8937 17503 8957
rect 17355 8874 17503 8937
rect 17355 8733 17504 8874
rect 17355 8455 17503 8733
rect 17355 8435 17359 8455
rect 17379 8435 17398 8455
rect 17418 8435 17437 8455
rect 17457 8435 17476 8455
rect 17496 8435 17503 8455
rect 17355 8373 17503 8435
rect 17355 8345 17370 8373
rect 17398 8345 17417 8373
rect 17445 8345 17464 8373
rect 17492 8345 17503 8373
rect 17355 8326 17503 8345
rect 17355 8298 17370 8326
rect 17398 8298 17417 8326
rect 17445 8298 17464 8326
rect 17492 8298 17503 8326
rect 17355 8279 17503 8298
rect 17355 8251 17370 8279
rect 17398 8251 17417 8279
rect 17445 8251 17464 8279
rect 17492 8251 17503 8279
rect 17355 7953 17503 8251
rect 17355 7933 17359 7953
rect 17379 7933 17398 7953
rect 17418 7933 17437 7953
rect 17457 7933 17476 7953
rect 17496 7933 17503 7953
rect 17355 7451 17503 7933
rect 17355 7431 17359 7451
rect 17379 7431 17398 7451
rect 17418 7431 17437 7451
rect 17457 7431 17476 7451
rect 17496 7431 17503 7451
rect 17355 7319 17503 7431
rect 17355 7291 17370 7319
rect 17398 7291 17417 7319
rect 17445 7291 17464 7319
rect 17492 7291 17503 7319
rect 17355 7272 17503 7291
rect 17355 7244 17370 7272
rect 17398 7244 17417 7272
rect 17445 7244 17464 7272
rect 17492 7244 17503 7272
rect 17355 7225 17503 7244
rect 17355 7197 17370 7225
rect 17398 7197 17417 7225
rect 17445 7197 17464 7225
rect 17492 7197 17503 7225
rect 17355 6949 17503 7197
rect 17355 6929 17359 6949
rect 17379 6929 17398 6949
rect 17418 6929 17437 6949
rect 17457 6929 17476 6949
rect 17496 6929 17503 6949
rect 17355 6447 17503 6929
rect 17355 6427 17359 6447
rect 17379 6427 17398 6447
rect 17418 6427 17437 6447
rect 17457 6427 17476 6447
rect 17496 6427 17503 6447
rect 17355 6361 17503 6427
rect 17354 6354 17503 6361
rect 17354 6326 17369 6354
rect 17397 6326 17416 6354
rect 17444 6326 17463 6354
rect 17491 6326 17503 6354
rect 17354 6307 17503 6326
rect 17354 6279 17369 6307
rect 17397 6279 17416 6307
rect 17444 6279 17463 6307
rect 17491 6279 17503 6307
rect 17354 6260 17503 6279
rect 17354 6232 17369 6260
rect 17397 6232 17416 6260
rect 17444 6232 17463 6260
rect 17491 6232 17503 6260
rect 17354 6221 17503 6232
rect 17167 6096 17170 6116
rect 17190 6096 17209 6116
rect 17229 6096 17248 6116
rect 17268 6096 17287 6116
rect 17307 6096 17315 6116
rect 17167 5895 17315 6096
rect 17167 5867 17182 5895
rect 17210 5867 17229 5895
rect 17257 5867 17276 5895
rect 17304 5867 17315 5895
rect 17167 5848 17315 5867
rect 17167 5820 17182 5848
rect 17210 5820 17229 5848
rect 17257 5820 17276 5848
rect 17304 5820 17315 5848
rect 17167 5801 17315 5820
rect 17167 5773 17182 5801
rect 17210 5773 17229 5801
rect 17257 5773 17276 5801
rect 17304 5773 17315 5801
rect 17167 5614 17315 5773
rect 17167 5594 17170 5614
rect 17190 5594 17209 5614
rect 17229 5594 17248 5614
rect 17268 5594 17287 5614
rect 17307 5594 17315 5614
rect 17167 5112 17315 5594
rect 17167 5092 17170 5112
rect 17190 5092 17209 5112
rect 17229 5092 17248 5112
rect 17268 5092 17287 5112
rect 17307 5092 17315 5112
rect 17167 4832 17315 5092
rect 17167 4804 17181 4832
rect 17209 4804 17228 4832
rect 17256 4804 17275 4832
rect 17303 4804 17315 4832
rect 17167 4785 17315 4804
rect 17167 4757 17181 4785
rect 17209 4757 17228 4785
rect 17256 4757 17275 4785
rect 17303 4757 17315 4785
rect 17167 4738 17315 4757
rect 17167 4710 17181 4738
rect 17209 4710 17228 4738
rect 17256 4710 17275 4738
rect 17303 4710 17315 4738
rect 17167 4610 17315 4710
rect 17167 4590 17170 4610
rect 17190 4590 17209 4610
rect 17229 4590 17248 4610
rect 17268 4590 17287 4610
rect 17307 4590 17315 4610
rect 17167 4108 17315 4590
rect 17167 4088 17170 4108
rect 17190 4088 17209 4108
rect 17229 4088 17248 4108
rect 17268 4088 17287 4108
rect 17307 4088 17315 4108
rect 17167 3844 17315 4088
rect 17167 3816 17182 3844
rect 17210 3816 17229 3844
rect 17257 3816 17276 3844
rect 17304 3816 17315 3844
rect 17167 3797 17315 3816
rect 17167 3769 17182 3797
rect 17210 3769 17229 3797
rect 17257 3769 17276 3797
rect 17304 3769 17315 3797
rect 17167 3750 17315 3769
rect 17167 3722 17182 3750
rect 17210 3722 17229 3750
rect 17257 3722 17276 3750
rect 17304 3722 17315 3750
rect 17167 3606 17315 3722
rect 17167 3586 17170 3606
rect 17190 3586 17209 3606
rect 17229 3586 17248 3606
rect 17268 3586 17287 3606
rect 17307 3586 17315 3606
rect 17167 3104 17315 3586
rect 17355 5945 17503 6221
rect 17355 5925 17359 5945
rect 17379 5925 17398 5945
rect 17418 5925 17437 5945
rect 17457 5925 17476 5945
rect 17496 5925 17503 5945
rect 17355 5904 17503 5925
rect 17545 8661 17613 9036
rect 17545 8641 17548 8661
rect 17568 8641 17587 8661
rect 17607 8641 17613 8661
rect 17545 8159 17613 8641
rect 17545 8139 17548 8159
rect 17568 8139 17587 8159
rect 17607 8139 17613 8159
rect 17545 7657 17613 8139
rect 17545 7637 17548 7657
rect 17568 7637 17587 7657
rect 17607 7637 17613 7657
rect 17545 7155 17613 7637
rect 17545 7135 17548 7155
rect 17568 7135 17587 7155
rect 17607 7135 17613 7155
rect 17545 6653 17613 7135
rect 17545 6633 17548 6653
rect 17568 6633 17587 6653
rect 17607 6633 17613 6653
rect 17545 6151 17613 6633
rect 17545 6131 17548 6151
rect 17568 6131 17587 6151
rect 17607 6131 17613 6151
rect 17355 5763 17504 5904
rect 17355 5443 17503 5763
rect 17355 5423 17359 5443
rect 17379 5423 17398 5443
rect 17418 5423 17437 5443
rect 17457 5423 17476 5443
rect 17496 5423 17503 5443
rect 17355 5346 17503 5423
rect 17355 5318 17370 5346
rect 17398 5318 17417 5346
rect 17445 5318 17464 5346
rect 17492 5318 17503 5346
rect 17355 5299 17503 5318
rect 17355 5271 17370 5299
rect 17398 5271 17417 5299
rect 17445 5271 17464 5299
rect 17492 5271 17503 5299
rect 17355 5252 17503 5271
rect 17355 5224 17370 5252
rect 17398 5224 17417 5252
rect 17445 5224 17464 5252
rect 17492 5224 17503 5252
rect 17355 4941 17503 5224
rect 17355 4921 17359 4941
rect 17379 4921 17398 4941
rect 17418 4921 17437 4941
rect 17457 4921 17476 4941
rect 17496 4921 17503 4941
rect 17355 4439 17503 4921
rect 17355 4419 17359 4439
rect 17379 4419 17398 4439
rect 17418 4419 17437 4439
rect 17457 4419 17476 4439
rect 17496 4419 17503 4439
rect 17355 4345 17503 4419
rect 17355 4317 17370 4345
rect 17398 4317 17417 4345
rect 17445 4317 17464 4345
rect 17492 4317 17503 4345
rect 17355 4298 17503 4317
rect 17355 4270 17370 4298
rect 17398 4270 17417 4298
rect 17445 4270 17464 4298
rect 17492 4270 17503 4298
rect 17355 4251 17503 4270
rect 17355 4223 17370 4251
rect 17398 4223 17417 4251
rect 17445 4223 17464 4251
rect 17492 4223 17503 4251
rect 17355 3937 17503 4223
rect 17355 3917 17359 3937
rect 17379 3917 17398 3937
rect 17418 3917 17437 3937
rect 17457 3917 17476 3937
rect 17496 3917 17503 3937
rect 17355 3853 17503 3917
rect 17545 5649 17613 6131
rect 17545 5629 17548 5649
rect 17568 5629 17587 5649
rect 17607 5629 17613 5649
rect 17545 5147 17613 5629
rect 17545 5127 17548 5147
rect 17568 5127 17587 5147
rect 17607 5127 17613 5147
rect 17545 4645 17613 5127
rect 17545 4625 17548 4645
rect 17568 4625 17587 4645
rect 17607 4625 17613 4645
rect 17545 4143 17613 4625
rect 17545 4123 17548 4143
rect 17568 4123 17587 4143
rect 17607 4123 17613 4143
rect 17355 3712 17504 3853
rect 17355 3435 17503 3712
rect 17355 3415 17359 3435
rect 17379 3415 17398 3435
rect 17418 3415 17437 3435
rect 17457 3415 17476 3435
rect 17496 3415 17503 3435
rect 17355 3353 17503 3415
rect 17354 3346 17503 3353
rect 17354 3318 17369 3346
rect 17397 3318 17416 3346
rect 17444 3318 17463 3346
rect 17491 3318 17503 3346
rect 17354 3299 17503 3318
rect 17354 3271 17369 3299
rect 17397 3271 17416 3299
rect 17444 3271 17463 3299
rect 17491 3271 17503 3299
rect 17354 3252 17503 3271
rect 17354 3224 17369 3252
rect 17397 3224 17416 3252
rect 17444 3224 17463 3252
rect 17491 3224 17503 3252
rect 17354 3213 17503 3224
rect 17167 3084 17170 3104
rect 17190 3084 17209 3104
rect 17229 3084 17248 3104
rect 17268 3084 17287 3104
rect 17307 3084 17315 3104
rect 17167 2822 17315 3084
rect 17167 2794 17182 2822
rect 17210 2794 17229 2822
rect 17257 2794 17276 2822
rect 17304 2794 17315 2822
rect 17167 2775 17315 2794
rect 17167 2747 17182 2775
rect 17210 2747 17229 2775
rect 17257 2747 17276 2775
rect 17304 2747 17315 2775
rect 17167 2728 17315 2747
rect 17167 2700 17182 2728
rect 17210 2700 17229 2728
rect 17257 2700 17276 2728
rect 17304 2700 17315 2728
rect 17167 2602 17315 2700
rect 17167 2582 17170 2602
rect 17190 2582 17209 2602
rect 17229 2582 17248 2602
rect 17268 2582 17287 2602
rect 17307 2582 17315 2602
rect 17167 2100 17315 2582
rect 17167 2080 17170 2100
rect 17190 2080 17209 2100
rect 17229 2080 17248 2100
rect 17268 2080 17287 2100
rect 17307 2080 17315 2100
rect 17167 1825 17315 2080
rect 17167 1797 17182 1825
rect 17210 1797 17229 1825
rect 17257 1797 17276 1825
rect 17304 1797 17315 1825
rect 17167 1778 17315 1797
rect 17167 1750 17182 1778
rect 17210 1750 17229 1778
rect 17257 1750 17276 1778
rect 17304 1750 17315 1778
rect 17167 1731 17315 1750
rect 17167 1703 17182 1731
rect 17210 1703 17229 1731
rect 17257 1703 17276 1731
rect 17304 1703 17315 1731
rect 17167 1598 17315 1703
rect 17167 1578 17170 1598
rect 17190 1578 17209 1598
rect 17229 1578 17248 1598
rect 17268 1578 17287 1598
rect 17307 1578 17315 1598
rect 17167 1096 17315 1578
rect 17167 1076 17170 1096
rect 17190 1076 17209 1096
rect 17229 1076 17248 1096
rect 17268 1076 17287 1096
rect 17307 1076 17315 1096
rect 17167 834 17315 1076
rect 17355 2933 17503 3213
rect 17355 2913 17359 2933
rect 17379 2913 17398 2933
rect 17418 2913 17437 2933
rect 17457 2913 17476 2933
rect 17496 2913 17503 2933
rect 17355 2831 17503 2913
rect 17545 3641 17613 4123
rect 17545 3621 17548 3641
rect 17568 3621 17587 3641
rect 17607 3621 17613 3641
rect 17545 3139 17613 3621
rect 17545 3119 17548 3139
rect 17568 3119 17587 3139
rect 17607 3119 17613 3139
rect 17355 2690 17504 2831
rect 17355 2431 17503 2690
rect 17355 2411 17359 2431
rect 17379 2411 17398 2431
rect 17418 2411 17437 2431
rect 17457 2411 17476 2431
rect 17496 2411 17503 2431
rect 17355 2312 17503 2411
rect 17355 2284 17370 2312
rect 17398 2284 17417 2312
rect 17445 2284 17464 2312
rect 17492 2284 17503 2312
rect 17355 2265 17503 2284
rect 17355 2237 17370 2265
rect 17398 2237 17417 2265
rect 17445 2237 17464 2265
rect 17492 2237 17503 2265
rect 17355 2218 17503 2237
rect 17355 2190 17370 2218
rect 17398 2190 17417 2218
rect 17445 2190 17464 2218
rect 17492 2190 17503 2218
rect 17355 1929 17503 2190
rect 17355 1909 17359 1929
rect 17379 1909 17398 1929
rect 17418 1909 17437 1929
rect 17457 1909 17476 1929
rect 17496 1909 17503 1929
rect 17355 1833 17503 1909
rect 17545 2637 17613 3119
rect 17545 2617 17548 2637
rect 17568 2617 17587 2637
rect 17607 2617 17613 2637
rect 17545 2135 17613 2617
rect 17545 2115 17548 2135
rect 17568 2115 17587 2135
rect 17607 2115 17613 2135
rect 17355 1692 17504 1833
rect 17355 1427 17503 1692
rect 17355 1407 17359 1427
rect 17379 1407 17398 1427
rect 17418 1407 17437 1427
rect 17457 1407 17476 1427
rect 17496 1407 17503 1427
rect 17355 1310 17503 1407
rect 17355 1282 17370 1310
rect 17398 1282 17417 1310
rect 17445 1282 17464 1310
rect 17492 1282 17503 1310
rect 17355 1263 17503 1282
rect 17355 1235 17370 1263
rect 17398 1235 17417 1263
rect 17445 1235 17464 1263
rect 17492 1235 17503 1263
rect 17355 1216 17503 1235
rect 17355 1188 17370 1216
rect 17398 1188 17417 1216
rect 17445 1188 17464 1216
rect 17492 1188 17503 1216
rect 17355 925 17503 1188
rect 17355 905 17359 925
rect 17379 905 17398 925
rect 17418 905 17437 925
rect 17457 905 17476 925
rect 17496 905 17503 925
rect 17355 834 17503 905
rect 17166 825 17315 834
rect 17166 797 17180 825
rect 17208 797 17227 825
rect 17255 797 17274 825
rect 17302 797 17315 825
rect 17166 778 17315 797
rect 17166 750 17180 778
rect 17208 750 17227 778
rect 17255 750 17274 778
rect 17302 750 17315 778
rect 17166 731 17315 750
rect 17166 703 17180 731
rect 17208 703 17227 731
rect 17255 703 17274 731
rect 17302 703 17315 731
rect 17166 693 17315 703
rect 17354 693 17503 834
rect -251 574 -245 594
rect -225 574 -206 594
rect -186 574 -167 594
rect -147 574 -128 594
rect -108 574 -105 594
rect -251 253 -105 574
rect -251 233 -245 253
rect -225 233 -206 253
rect -186 233 -167 253
rect -147 233 -128 253
rect -108 233 -105 253
rect -251 197 -105 233
rect -251 177 -245 197
rect -225 177 -206 197
rect -186 177 -167 197
rect -147 177 -128 197
rect -108 177 -105 197
rect -251 92 -105 177
rect -251 72 -245 92
rect -225 72 -206 92
rect -186 72 -167 92
rect -147 72 -128 92
rect -108 72 -105 92
rect -251 -85 -105 72
rect 17167 594 17315 693
rect 17167 574 17170 594
rect 17190 574 17209 594
rect 17229 574 17248 594
rect 17268 574 17287 594
rect 17307 574 17315 594
rect 17167 92 17315 574
rect 17167 72 17170 92
rect 17190 72 17209 92
rect 17229 72 17248 92
rect 17268 72 17287 92
rect 17307 72 17315 92
rect -251 -113 -241 -85
rect -213 -113 -194 -85
rect -166 -113 -147 -85
rect -119 -113 -105 -85
rect -251 -132 -105 -113
rect -251 -160 -241 -132
rect -213 -160 -194 -132
rect -166 -160 -147 -132
rect -119 -160 -105 -132
rect -251 -179 -105 -160
rect -251 -207 -241 -179
rect -213 -207 -194 -179
rect -166 -207 -147 -179
rect -119 -207 -105 -179
rect -251 -457 -105 -207
rect 427 -292 444 0
rect 422 -295 444 -292
rect 422 -312 425 -295
rect 442 -312 444 -295
rect 422 -316 444 -312
rect 929 -457 946 0
rect 1431 -457 1448 0
rect 1933 -457 1950 0
rect 2435 -457 2452 0
rect 2937 -457 2954 0
rect 3439 -457 3456 0
rect 3941 -457 3958 0
rect 4443 -457 4460 0
rect 4779 -457 4796 0
rect 4945 -457 4962 0
rect 5447 -457 5464 0
rect 5949 -457 5966 0
rect 6451 -457 6468 0
rect 6953 -457 6970 0
rect 7455 -457 7472 0
rect 7957 -457 7974 0
rect 8459 -457 8476 0
rect 8795 -457 8812 0
rect 8961 -457 8978 0
rect 9463 -457 9480 0
rect 9965 -457 9982 0
rect 10467 -457 10484 0
rect 10969 -457 10986 0
rect 11471 -457 11488 0
rect 11973 -457 11990 0
rect 12475 -457 12492 0
rect 12811 -457 12828 0
rect 12977 -457 12994 0
rect 13479 -60 13496 0
rect 13079 -77 13496 -60
rect 13079 -457 13096 -77
rect 13981 -95 13998 0
rect 13181 -112 13998 -95
rect 13181 -457 13198 -112
rect 13283 -136 13300 -135
rect 13283 -457 13300 -153
rect 14483 -136 14500 0
rect 14483 -157 14500 -153
rect 13385 -175 13402 -174
rect 13385 -457 13402 -192
rect 14985 -175 15002 0
rect 14985 -196 15002 -192
rect 13487 -213 13504 -212
rect 13487 -457 13504 -230
rect 15487 -213 15504 0
rect 15487 -234 15504 -230
rect 13589 -251 13606 -250
rect 13589 -457 13606 -268
rect 15989 -251 16006 0
rect 16238 -26 16255 0
rect 15989 -272 16006 -268
rect 16043 -43 16255 -26
rect 13691 -289 13708 -288
rect 13691 -457 13708 -306
rect 16043 -456 16060 -43
rect 16104 -64 16121 -61
rect 16104 -456 16121 -81
rect 16274 -113 16291 0
rect 16348 -64 16365 0
rect 16348 -85 16365 -81
rect 16274 -135 16418 -113
rect 16401 -432 16418 -135
rect 16491 -289 16508 0
rect 16491 -310 16508 -306
rect 16993 -295 17010 0
rect 17167 -20 17315 72
rect 17167 -48 17181 -20
rect 17209 -48 17228 -20
rect 17256 -48 17275 -20
rect 17303 -48 17315 -20
rect 17167 -67 17315 -48
rect 17167 -95 17181 -67
rect 17209 -95 17228 -67
rect 17256 -95 17275 -67
rect 17303 -95 17315 -67
rect 17167 -114 17315 -95
rect 17167 -142 17181 -114
rect 17209 -142 17228 -114
rect 17256 -142 17275 -114
rect 17303 -142 17315 -114
rect 16993 -298 17014 -295
rect 16993 -315 16995 -298
rect 17012 -315 17014 -298
rect 16993 -318 17014 -315
rect 17167 -392 17315 -142
rect 17355 423 17503 693
rect 17355 403 17359 423
rect 17379 403 17398 423
rect 17418 403 17437 423
rect 17457 403 17476 423
rect 17496 403 17503 423
rect 17355 313 17503 403
rect 17355 285 17370 313
rect 17398 285 17417 313
rect 17445 285 17464 313
rect 17492 285 17503 313
rect 17355 266 17503 285
rect 17355 238 17370 266
rect 17398 238 17417 266
rect 17445 238 17464 266
rect 17492 238 17503 266
rect 17355 219 17503 238
rect 17355 191 17370 219
rect 17398 191 17417 219
rect 17445 191 17464 219
rect 17492 191 17503 219
rect 17355 -238 17503 191
rect 17545 1633 17613 2115
rect 17545 1613 17548 1633
rect 17568 1613 17587 1633
rect 17607 1613 17613 1633
rect 17545 1131 17613 1613
rect 17545 1111 17548 1131
rect 17568 1111 17587 1131
rect 17607 1111 17613 1131
rect 17545 629 17613 1111
rect 17632 9030 17839 9053
rect 17632 9013 17650 9030
rect 17825 9013 17839 9030
rect 17632 8990 17839 9013
rect 17632 8973 17650 8990
rect 17825 8973 17839 8990
rect 17632 8950 17839 8973
rect 17632 8933 17650 8950
rect 17825 8933 17839 8950
rect 17632 8910 17839 8933
rect 17632 8893 17650 8910
rect 17825 8893 17839 8910
rect 17632 8874 17839 8893
rect 17632 8870 17840 8874
rect 17632 8853 17650 8870
rect 17825 8853 17840 8870
rect 17632 8830 17840 8853
rect 17632 8813 17650 8830
rect 17825 8813 17840 8830
rect 17632 8790 17840 8813
rect 17632 8773 17650 8790
rect 17825 8773 17840 8790
rect 17632 8750 17840 8773
rect 17632 8733 17650 8750
rect 17825 8733 17840 8750
rect 17632 8710 17839 8733
rect 17632 8693 17650 8710
rect 17825 8693 17839 8710
rect 17632 8670 17839 8693
rect 17632 8653 17650 8670
rect 17825 8653 17839 8670
rect 17632 8630 17839 8653
rect 17632 8613 17650 8630
rect 17825 8613 17839 8630
rect 17632 8590 17839 8613
rect 17632 8573 17650 8590
rect 17825 8573 17839 8590
rect 17632 8550 17839 8573
rect 17632 8533 17650 8550
rect 17825 8533 17839 8550
rect 17632 8510 17839 8533
rect 17632 8493 17650 8510
rect 17825 8493 17839 8510
rect 17632 8470 17839 8493
rect 17632 8453 17650 8470
rect 17825 8453 17839 8470
rect 17632 8430 17839 8453
rect 17632 8413 17650 8430
rect 17825 8413 17839 8430
rect 17632 8390 17839 8413
rect 17632 8373 17650 8390
rect 17825 8373 17839 8390
rect 17632 8350 17839 8373
rect 17632 8333 17650 8350
rect 17825 8333 17839 8350
rect 17632 8310 17839 8333
rect 17632 8293 17650 8310
rect 17825 8293 17839 8310
rect 17632 8270 17839 8293
rect 17632 8253 17650 8270
rect 17825 8253 17839 8270
rect 17632 8230 17839 8253
rect 17632 8213 17650 8230
rect 17825 8213 17839 8230
rect 17632 8190 17839 8213
rect 17632 8173 17650 8190
rect 17825 8173 17839 8190
rect 17632 8150 17839 8173
rect 17632 8133 17650 8150
rect 17825 8133 17839 8150
rect 17632 8110 17839 8133
rect 17632 8093 17650 8110
rect 17825 8093 17839 8110
rect 17632 8070 17839 8093
rect 17632 8053 17650 8070
rect 17825 8053 17839 8070
rect 17632 8030 17839 8053
rect 17632 8013 17650 8030
rect 17825 8013 17839 8030
rect 17632 7990 17839 8013
rect 17632 7973 17650 7990
rect 17825 7973 17839 7990
rect 17632 7950 17839 7973
rect 17632 7933 17650 7950
rect 17825 7933 17839 7950
rect 17632 7910 17839 7933
rect 17632 7893 17650 7910
rect 17825 7893 17839 7910
rect 17632 7870 17839 7893
rect 17632 7853 17650 7870
rect 17825 7853 17839 7870
rect 17632 7830 17839 7853
rect 17632 7813 17650 7830
rect 17825 7813 17839 7830
rect 17632 7790 17839 7813
rect 17632 7773 17650 7790
rect 17825 7773 17839 7790
rect 17632 7750 17839 7773
rect 17632 7733 17650 7750
rect 17825 7733 17839 7750
rect 17632 7710 17839 7733
rect 17632 7693 17650 7710
rect 17825 7693 17839 7710
rect 17632 7670 17839 7693
rect 17632 7653 17650 7670
rect 17825 7653 17839 7670
rect 17632 7630 17839 7653
rect 17632 7613 17650 7630
rect 17825 7613 17839 7630
rect 17632 7590 17839 7613
rect 17632 7573 17650 7590
rect 17825 7573 17839 7590
rect 17632 7550 17839 7573
rect 17632 7533 17650 7550
rect 17825 7533 17839 7550
rect 17632 7510 17839 7533
rect 17632 7493 17650 7510
rect 17825 7493 17839 7510
rect 17632 7470 17839 7493
rect 17632 7453 17650 7470
rect 17825 7453 17839 7470
rect 17632 7430 17839 7453
rect 17632 7413 17650 7430
rect 17825 7413 17839 7430
rect 17632 7390 17839 7413
rect 17632 7373 17650 7390
rect 17825 7373 17839 7390
rect 17632 7350 17839 7373
rect 17632 7333 17650 7350
rect 17825 7333 17839 7350
rect 17632 7310 17839 7333
rect 17632 7293 17650 7310
rect 17825 7293 17839 7310
rect 17632 7270 17839 7293
rect 17632 7253 17650 7270
rect 17825 7253 17839 7270
rect 17632 7230 17839 7253
rect 17632 7213 17650 7230
rect 17825 7213 17839 7230
rect 17632 7190 17839 7213
rect 17632 7173 17650 7190
rect 17825 7173 17839 7190
rect 17632 7150 17839 7173
rect 17632 7133 17650 7150
rect 17825 7133 17839 7150
rect 17632 7110 17839 7133
rect 17632 7093 17650 7110
rect 17825 7093 17839 7110
rect 17632 7070 17839 7093
rect 17632 7053 17650 7070
rect 17825 7053 17839 7070
rect 17632 7030 17839 7053
rect 17632 7013 17650 7030
rect 17825 7013 17839 7030
rect 17632 6990 17839 7013
rect 17632 6973 17650 6990
rect 17825 6973 17839 6990
rect 17632 6950 17839 6973
rect 17632 6933 17650 6950
rect 17825 6933 17839 6950
rect 17632 6910 17839 6933
rect 17632 6893 17650 6910
rect 17825 6893 17839 6910
rect 17632 6870 17839 6893
rect 17632 6853 17650 6870
rect 17825 6853 17839 6870
rect 17632 6830 17839 6853
rect 17632 6813 17650 6830
rect 17825 6813 17839 6830
rect 17632 6790 17839 6813
rect 17632 6773 17650 6790
rect 17825 6773 17839 6790
rect 17632 6750 17839 6773
rect 17632 6733 17650 6750
rect 17825 6733 17839 6750
rect 17632 6710 17839 6733
rect 17632 6693 17650 6710
rect 17825 6693 17839 6710
rect 17632 6670 17839 6693
rect 17632 6653 17650 6670
rect 17825 6653 17839 6670
rect 17632 6630 17839 6653
rect 17632 6613 17650 6630
rect 17825 6613 17839 6630
rect 17632 6590 17839 6613
rect 17632 6573 17650 6590
rect 17825 6573 17839 6590
rect 17632 6550 17839 6573
rect 17632 6533 17650 6550
rect 17825 6533 17839 6550
rect 17632 6510 17839 6533
rect 17632 6493 17650 6510
rect 17825 6493 17839 6510
rect 17632 6470 17839 6493
rect 17632 6453 17650 6470
rect 17825 6453 17839 6470
rect 17632 6430 17839 6453
rect 17632 6413 17650 6430
rect 17825 6413 17839 6430
rect 17632 6390 17839 6413
rect 17632 6373 17650 6390
rect 17825 6373 17839 6390
rect 17632 6350 17839 6373
rect 17870 6361 18077 9134
rect 20151 9168 20567 9181
rect 20151 8962 20448 9168
rect 20554 8962 20567 9168
rect 20151 8950 20567 8962
rect 20151 8289 20567 8302
rect 20151 8083 20448 8289
rect 20554 8083 20567 8289
rect 20151 8071 20567 8083
rect 20151 7168 20567 7181
rect 20151 6962 20448 7168
rect 20554 6962 20567 7168
rect 20151 6950 20567 6962
rect 17632 6333 17650 6350
rect 17825 6333 17839 6350
rect 17632 6310 17839 6333
rect 17632 6293 17650 6310
rect 17825 6293 17839 6310
rect 17632 6270 17839 6293
rect 17632 6253 17650 6270
rect 17825 6253 17839 6270
rect 17632 6229 17839 6253
rect 17632 6212 17651 6229
rect 17826 6212 17839 6229
rect 17869 6221 18077 6361
rect 17632 6190 17839 6212
rect 17632 6173 17650 6190
rect 17825 6173 17839 6190
rect 17632 6150 17839 6173
rect 17632 6133 17650 6150
rect 17825 6133 17839 6150
rect 17632 6110 17839 6133
rect 17632 6093 17650 6110
rect 17825 6093 17839 6110
rect 17632 6070 17839 6093
rect 17632 6053 17650 6070
rect 17825 6053 17839 6070
rect 17632 6030 17839 6053
rect 17632 6013 17650 6030
rect 17825 6013 17839 6030
rect 17632 5990 17839 6013
rect 17632 5973 17650 5990
rect 17825 5973 17839 5990
rect 17632 5950 17839 5973
rect 17632 5933 17650 5950
rect 17825 5933 17839 5950
rect 17632 5910 17839 5933
rect 17632 5893 17650 5910
rect 17825 5904 17839 5910
rect 17825 5893 17840 5904
rect 17632 5870 17840 5893
rect 17632 5853 17650 5870
rect 17825 5853 17840 5870
rect 17632 5830 17840 5853
rect 17632 5813 17650 5830
rect 17825 5813 17840 5830
rect 17632 5790 17840 5813
rect 17632 5773 17650 5790
rect 17825 5773 17840 5790
rect 17632 5763 17840 5773
rect 17632 5750 17839 5763
rect 17632 5733 17650 5750
rect 17825 5733 17839 5750
rect 17632 5710 17839 5733
rect 17632 5693 17650 5710
rect 17825 5693 17839 5710
rect 17632 5670 17839 5693
rect 17632 5653 17650 5670
rect 17825 5653 17839 5670
rect 17632 5630 17839 5653
rect 17632 5613 17650 5630
rect 17825 5613 17839 5630
rect 17632 5590 17839 5613
rect 17632 5573 17650 5590
rect 17825 5573 17839 5590
rect 17632 5550 17839 5573
rect 17632 5533 17650 5550
rect 17825 5533 17839 5550
rect 17632 5510 17839 5533
rect 17632 5493 17650 5510
rect 17825 5493 17839 5510
rect 17632 5470 17839 5493
rect 17632 5453 17650 5470
rect 17825 5453 17839 5470
rect 17632 5430 17839 5453
rect 17632 5413 17650 5430
rect 17825 5413 17839 5430
rect 17632 5390 17839 5413
rect 17632 5373 17650 5390
rect 17825 5373 17839 5390
rect 17632 5349 17839 5373
rect 17632 5332 17649 5349
rect 17824 5332 17839 5349
rect 17632 5310 17839 5332
rect 17632 5293 17650 5310
rect 17825 5293 17839 5310
rect 17632 5270 17839 5293
rect 17632 5253 17650 5270
rect 17825 5253 17839 5270
rect 17632 5230 17839 5253
rect 17632 5213 17650 5230
rect 17825 5213 17839 5230
rect 17632 5190 17839 5213
rect 17632 5173 17650 5190
rect 17825 5173 17839 5190
rect 17632 5150 17839 5173
rect 17632 5133 17650 5150
rect 17825 5133 17839 5150
rect 17632 5110 17839 5133
rect 17632 5093 17650 5110
rect 17825 5093 17839 5110
rect 17632 5070 17839 5093
rect 17632 5053 17650 5070
rect 17825 5053 17839 5070
rect 17632 5030 17839 5053
rect 17632 5013 17650 5030
rect 17825 5013 17839 5030
rect 17632 4990 17839 5013
rect 17632 4973 17650 4990
rect 17825 4973 17839 4990
rect 17632 4950 17839 4973
rect 17632 4933 17650 4950
rect 17825 4933 17839 4950
rect 17632 4910 17839 4933
rect 17632 4893 17650 4910
rect 17825 4893 17839 4910
rect 17632 4870 17839 4893
rect 17632 4853 17650 4870
rect 17825 4853 17839 4870
rect 17632 4830 17839 4853
rect 17632 4813 17650 4830
rect 17825 4813 17839 4830
rect 17632 4790 17839 4813
rect 17632 4773 17650 4790
rect 17825 4773 17839 4790
rect 17632 4750 17839 4773
rect 17632 4733 17650 4750
rect 17825 4733 17839 4750
rect 17632 4710 17839 4733
rect 17632 4693 17650 4710
rect 17825 4693 17839 4710
rect 17632 4670 17839 4693
rect 17632 4653 17650 4670
rect 17825 4653 17839 4670
rect 17632 4630 17839 4653
rect 17632 4613 17650 4630
rect 17825 4613 17839 4630
rect 17632 4590 17839 4613
rect 17632 4573 17650 4590
rect 17825 4573 17839 4590
rect 17632 4550 17839 4573
rect 17632 4533 17650 4550
rect 17825 4533 17839 4550
rect 17632 4510 17839 4533
rect 17632 4493 17650 4510
rect 17825 4493 17839 4510
rect 17632 4470 17839 4493
rect 17632 4453 17650 4470
rect 17825 4453 17839 4470
rect 17632 4430 17839 4453
rect 17632 4413 17650 4430
rect 17825 4413 17839 4430
rect 17632 4390 17839 4413
rect 17632 4373 17650 4390
rect 17825 4373 17839 4390
rect 17632 4350 17839 4373
rect 17632 4333 17650 4350
rect 17825 4333 17839 4350
rect 17632 4310 17839 4333
rect 17632 4293 17650 4310
rect 17825 4293 17839 4310
rect 17632 4270 17839 4293
rect 17632 4253 17650 4270
rect 17825 4253 17839 4270
rect 17632 4230 17839 4253
rect 17632 4213 17650 4230
rect 17825 4213 17839 4230
rect 17632 4190 17839 4213
rect 17632 4173 17650 4190
rect 17825 4173 17839 4190
rect 17632 4150 17839 4173
rect 17632 4133 17650 4150
rect 17825 4133 17839 4150
rect 17632 4110 17839 4133
rect 17632 4093 17650 4110
rect 17825 4093 17839 4110
rect 17632 4070 17839 4093
rect 17632 4053 17650 4070
rect 17825 4053 17839 4070
rect 17632 4030 17839 4053
rect 17632 4013 17650 4030
rect 17825 4013 17839 4030
rect 17632 3990 17839 4013
rect 17632 3973 17650 3990
rect 17825 3973 17839 3990
rect 17632 3950 17839 3973
rect 17632 3933 17650 3950
rect 17825 3933 17839 3950
rect 17632 3910 17839 3933
rect 17632 3893 17650 3910
rect 17825 3893 17839 3910
rect 17632 3870 17839 3893
rect 17632 3853 17650 3870
rect 17825 3853 17839 3870
rect 17632 3830 17840 3853
rect 17632 3813 17650 3830
rect 17825 3813 17840 3830
rect 17632 3790 17840 3813
rect 17632 3773 17650 3790
rect 17825 3773 17840 3790
rect 17632 3750 17840 3773
rect 17632 3733 17650 3750
rect 17825 3733 17840 3750
rect 17632 3712 17840 3733
rect 17632 3710 17839 3712
rect 17632 3693 17650 3710
rect 17825 3693 17839 3710
rect 17632 3670 17839 3693
rect 17632 3653 17650 3670
rect 17825 3653 17839 3670
rect 17632 3630 17839 3653
rect 17632 3613 17650 3630
rect 17825 3613 17839 3630
rect 17632 3590 17839 3613
rect 17632 3573 17650 3590
rect 17825 3573 17839 3590
rect 17632 3550 17839 3573
rect 17632 3533 17650 3550
rect 17825 3533 17839 3550
rect 17632 3510 17839 3533
rect 17632 3493 17650 3510
rect 17825 3493 17839 3510
rect 17632 3470 17839 3493
rect 17632 3453 17650 3470
rect 17825 3453 17839 3470
rect 17632 3430 17839 3453
rect 17632 3413 17650 3430
rect 17825 3413 17839 3430
rect 17632 3390 17839 3413
rect 17632 3373 17650 3390
rect 17825 3373 17839 3390
rect 17632 3350 17839 3373
rect 17870 3353 18077 6221
rect 20151 6289 20567 6302
rect 20151 6083 20448 6289
rect 20554 6083 20567 6289
rect 20151 6071 20567 6083
rect 20151 5168 20567 5181
rect 20151 4962 20448 5168
rect 20554 4962 20567 5168
rect 20151 4950 20567 4962
rect 20151 4289 20567 4302
rect 20151 4083 20448 4289
rect 20554 4083 20567 4289
rect 20151 4071 20567 4083
rect 17632 3333 17650 3350
rect 17825 3333 17839 3350
rect 17632 3310 17839 3333
rect 17632 3293 17650 3310
rect 17825 3293 17839 3310
rect 17632 3270 17839 3293
rect 17632 3253 17650 3270
rect 17825 3253 17839 3270
rect 17632 3230 17839 3253
rect 17632 3213 17650 3230
rect 17825 3213 17839 3230
rect 17869 3213 18077 3353
rect 17632 3190 17839 3213
rect 17632 3173 17650 3190
rect 17825 3173 17839 3190
rect 17632 3150 17839 3173
rect 17632 3133 17650 3150
rect 17825 3133 17839 3150
rect 17632 3110 17839 3133
rect 17632 3093 17650 3110
rect 17825 3093 17839 3110
rect 17632 3070 17839 3093
rect 17632 3053 17650 3070
rect 17825 3053 17839 3070
rect 17632 3030 17839 3053
rect 17632 3013 17650 3030
rect 17825 3013 17839 3030
rect 17632 2990 17839 3013
rect 17632 2973 17650 2990
rect 17825 2973 17839 2990
rect 17632 2950 17839 2973
rect 17632 2933 17650 2950
rect 17825 2933 17839 2950
rect 17632 2910 17839 2933
rect 17632 2893 17650 2910
rect 17825 2893 17839 2910
rect 17632 2870 17839 2893
rect 17632 2853 17650 2870
rect 17825 2853 17839 2870
rect 17632 2831 17839 2853
rect 17632 2830 17840 2831
rect 17632 2813 17650 2830
rect 17825 2813 17840 2830
rect 17632 2790 17840 2813
rect 17632 2773 17650 2790
rect 17825 2773 17840 2790
rect 17632 2750 17840 2773
rect 17632 2733 17650 2750
rect 17825 2733 17840 2750
rect 17632 2710 17840 2733
rect 17632 2693 17650 2710
rect 17825 2693 17840 2710
rect 17632 2690 17840 2693
rect 17632 2670 17839 2690
rect 17632 2653 17650 2670
rect 17825 2653 17839 2670
rect 17632 2630 17839 2653
rect 17632 2613 17650 2630
rect 17825 2613 17839 2630
rect 17632 2590 17839 2613
rect 17632 2573 17650 2590
rect 17825 2573 17839 2590
rect 17632 2550 17839 2573
rect 17632 2533 17650 2550
rect 17825 2533 17839 2550
rect 17632 2510 17839 2533
rect 17632 2493 17650 2510
rect 17825 2493 17839 2510
rect 17632 2470 17839 2493
rect 17632 2453 17650 2470
rect 17825 2453 17839 2470
rect 17632 2430 17839 2453
rect 17632 2413 17650 2430
rect 17825 2413 17839 2430
rect 17632 2390 17839 2413
rect 17632 2373 17650 2390
rect 17825 2373 17839 2390
rect 17632 2350 17839 2373
rect 17632 2333 17650 2350
rect 17825 2333 17839 2350
rect 17632 2310 17839 2333
rect 17632 2293 17650 2310
rect 17825 2293 17839 2310
rect 17632 2267 17839 2293
rect 17632 2250 17650 2267
rect 17825 2250 17839 2267
rect 17632 2230 17839 2250
rect 17632 2213 17650 2230
rect 17825 2213 17839 2230
rect 17632 2190 17839 2213
rect 17632 2173 17650 2190
rect 17825 2173 17839 2190
rect 17632 2150 17839 2173
rect 17632 2133 17650 2150
rect 17825 2133 17839 2150
rect 17632 2110 17839 2133
rect 17632 2093 17650 2110
rect 17825 2093 17839 2110
rect 17632 2070 17839 2093
rect 17632 2053 17650 2070
rect 17825 2053 17839 2070
rect 17632 2030 17839 2053
rect 17632 2013 17650 2030
rect 17825 2013 17839 2030
rect 17632 1990 17839 2013
rect 17632 1973 17650 1990
rect 17825 1973 17839 1990
rect 17632 1950 17839 1973
rect 17632 1933 17650 1950
rect 17825 1933 17839 1950
rect 17632 1910 17839 1933
rect 17632 1893 17650 1910
rect 17825 1893 17839 1910
rect 17632 1870 17839 1893
rect 17632 1853 17650 1870
rect 17825 1853 17839 1870
rect 17632 1830 17839 1853
rect 17632 1813 17650 1830
rect 17825 1813 17839 1830
rect 17632 1790 17839 1813
rect 17632 1773 17650 1790
rect 17825 1773 17839 1790
rect 17632 1750 17839 1773
rect 17632 1733 17650 1750
rect 17825 1733 17839 1750
rect 17632 1710 17839 1733
rect 17632 1693 17650 1710
rect 17825 1693 17839 1710
rect 17632 1670 17839 1693
rect 17632 1653 17650 1670
rect 17825 1653 17839 1670
rect 17632 1630 17839 1653
rect 17632 1613 17650 1630
rect 17825 1613 17839 1630
rect 17632 1590 17839 1613
rect 17632 1573 17650 1590
rect 17825 1573 17839 1590
rect 17632 1550 17839 1573
rect 17632 1533 17650 1550
rect 17825 1533 17839 1550
rect 17632 1510 17839 1533
rect 17632 1493 17650 1510
rect 17825 1493 17839 1510
rect 17632 1470 17839 1493
rect 17632 1453 17650 1470
rect 17825 1453 17839 1470
rect 17632 1430 17839 1453
rect 17632 1413 17650 1430
rect 17825 1413 17839 1430
rect 17632 1390 17839 1413
rect 17632 1373 17650 1390
rect 17825 1373 17839 1390
rect 17632 1350 17839 1373
rect 17632 1333 17650 1350
rect 17825 1333 17839 1350
rect 17632 1310 17839 1333
rect 17632 1293 17650 1310
rect 17825 1293 17839 1310
rect 17632 1270 17839 1293
rect 17632 1253 17650 1270
rect 17825 1253 17839 1270
rect 17632 1230 17839 1253
rect 17632 1213 17650 1230
rect 17825 1213 17839 1230
rect 17632 1190 17839 1213
rect 17632 1173 17650 1190
rect 17825 1173 17839 1190
rect 17632 1150 17839 1173
rect 17632 1133 17650 1150
rect 17825 1133 17839 1150
rect 17632 1110 17839 1133
rect 17632 1093 17650 1110
rect 17825 1093 17839 1110
rect 17632 1070 17839 1093
rect 17632 1053 17650 1070
rect 17825 1053 17839 1070
rect 17632 1030 17839 1053
rect 17632 1013 17650 1030
rect 17825 1013 17839 1030
rect 17632 990 17839 1013
rect 17632 973 17650 990
rect 17825 973 17839 990
rect 17632 950 17839 973
rect 17632 933 17650 950
rect 17825 933 17839 950
rect 17632 910 17839 933
rect 17632 893 17650 910
rect 17825 893 17839 910
rect 17632 870 17839 893
rect 17632 853 17650 870
rect 17825 853 17839 870
rect 17632 834 17839 853
rect 17631 830 17839 834
rect 17631 813 17650 830
rect 17825 813 17839 830
rect 17631 790 17839 813
rect 17631 773 17650 790
rect 17825 773 17839 790
rect 17631 750 17839 773
rect 17631 733 17650 750
rect 17825 733 17839 750
rect 17631 710 17839 733
rect 17631 693 17650 710
rect 17825 693 17839 710
rect 17545 609 17548 629
rect 17568 609 17587 629
rect 17607 609 17613 629
rect 17545 127 17613 609
rect 17545 107 17548 127
rect 17568 107 17587 127
rect 17607 107 17613 127
rect 17545 0 17613 107
rect 17632 670 17839 693
rect 17632 653 17650 670
rect 17825 653 17839 670
rect 17632 630 17839 653
rect 17632 613 17650 630
rect 17825 613 17839 630
rect 17632 590 17839 613
rect 17632 573 17650 590
rect 17825 573 17839 590
rect 17632 550 17839 573
rect 17632 533 17650 550
rect 17825 533 17839 550
rect 17632 510 17839 533
rect 17632 493 17650 510
rect 17825 493 17839 510
rect 17632 470 17839 493
rect 17632 453 17650 470
rect 17825 453 17839 470
rect 17632 430 17839 453
rect 17632 413 17650 430
rect 17825 413 17839 430
rect 17632 390 17839 413
rect 17632 373 17650 390
rect 17825 373 17839 390
rect 17632 350 17839 373
rect 17632 333 17650 350
rect 17825 333 17839 350
rect 17632 310 17839 333
rect 17632 293 17650 310
rect 17825 293 17839 310
rect 17632 270 17839 293
rect 17632 253 17650 270
rect 17825 253 17839 270
rect 17632 230 17839 253
rect 17632 213 17650 230
rect 17825 213 17839 230
rect 17632 190 17839 213
rect 17632 173 17650 190
rect 17825 173 17839 190
rect 17632 150 17839 173
rect 17632 133 17650 150
rect 17825 133 17839 150
rect 17632 110 17839 133
rect 17632 93 17650 110
rect 17825 93 17839 110
rect 17632 70 17839 93
rect 17632 53 17650 70
rect 17825 53 17839 70
rect 17632 30 17839 53
rect 17632 13 17650 30
rect 17825 13 17839 30
rect 17632 -152 17839 13
rect 17355 -266 17370 -238
rect 17398 -266 17417 -238
rect 17445 -266 17464 -238
rect 17492 -266 17503 -238
rect 17355 -285 17503 -266
rect 17355 -313 17370 -285
rect 17398 -313 17417 -285
rect 17445 -313 17464 -285
rect 17492 -313 17503 -285
rect 17355 -332 17503 -313
rect 17355 -360 17370 -332
rect 17398 -360 17417 -332
rect 17445 -360 17464 -332
rect 17492 -360 17503 -332
rect 17355 -392 17503 -360
rect 17870 -371 18077 3213
rect 20151 3168 20567 3181
rect 20151 2962 20448 3168
rect 20554 2962 20567 3168
rect 20151 2950 20567 2962
rect 20151 2289 20567 2302
rect 20151 2083 20448 2289
rect 20554 2083 20567 2289
rect 20151 2071 20567 2083
rect 20151 1168 20567 1181
rect 20151 962 20448 1168
rect 20554 962 20567 1168
rect 20151 950 20567 962
rect 20151 289 20567 302
rect 20151 83 20448 289
rect 20554 83 20567 289
rect 20151 71 20567 83
rect 16437 -432 16454 -429
rect 16395 -449 16401 -432
rect 16418 -449 16437 -432
rect 16454 -449 16460 -432
rect 16401 -456 16418 -449
rect 16437 -453 16454 -449
<< viali >>
rect 20448 10962 20554 11168
rect 20448 10083 20554 10289
rect 299 9516 430 9595
rect -430 9455 -402 9483
rect -383 9455 -355 9483
rect -336 9455 -308 9483
rect -430 9408 -402 9436
rect -383 9408 -355 9436
rect -336 9408 -308 9436
rect -430 9361 -402 9389
rect -383 9361 -355 9389
rect -336 9361 -308 9389
rect -943 8853 -768 8870
rect -943 8413 -768 8430
rect -943 7973 -768 7990
rect -943 7533 -768 7550
rect -943 7093 -768 7110
rect -943 6653 -768 6670
rect -943 6213 -768 6230
rect -943 5773 -768 5790
rect -943 5333 -768 5350
rect -943 4893 -768 4910
rect -943 4453 -768 4470
rect -943 4013 -768 4030
rect -943 3573 -768 3590
rect -943 3133 -768 3150
rect -943 2693 -768 2710
rect -943 2253 -768 2270
rect -943 1813 -768 1830
rect -943 1373 -768 1390
rect -943 933 -768 950
rect -943 493 -768 510
rect -943 53 -768 70
rect -651 8407 -634 8424
rect -651 7905 -634 7922
rect -651 7403 -634 7420
rect -651 6901 -634 6918
rect -651 6399 -634 6416
rect -651 5897 -634 5914
rect -651 5395 -634 5412
rect -651 4893 -634 4910
rect -651 4391 -634 4408
rect -651 3889 -634 3906
rect -651 3387 -634 3404
rect -651 2885 -634 2902
rect -651 2383 -634 2400
rect -651 1881 -634 1898
rect -651 1379 -634 1396
rect -651 877 -634 894
rect -597 8213 -580 8230
rect -597 7711 -580 7728
rect -597 7209 -580 7226
rect -597 6707 -580 6724
rect -597 6205 -580 6222
rect -597 5703 -580 5720
rect -597 5201 -580 5218
rect -597 4699 -580 4716
rect -597 4197 -580 4214
rect -597 3695 -580 3712
rect -597 3193 -580 3210
rect -597 2691 -580 2708
rect -597 2189 -580 2206
rect -597 1687 -580 1704
rect -597 1185 -580 1202
rect -597 683 -580 700
rect -545 8641 -525 8661
rect -506 8641 -486 8661
rect -545 8139 -525 8159
rect -506 8139 -486 8159
rect -545 7637 -525 7657
rect -506 7637 -486 7657
rect -545 7135 -525 7155
rect -506 7135 -486 7155
rect -545 6633 -525 6653
rect -506 6633 -486 6653
rect -545 6131 -525 6151
rect -506 6131 -486 6151
rect -545 5629 -525 5649
rect -506 5629 -486 5649
rect -545 5127 -525 5147
rect -506 5127 -486 5147
rect -545 4625 -525 4645
rect -506 4625 -486 4645
rect -545 4123 -525 4143
rect -506 4123 -486 4143
rect -545 3621 -525 3641
rect -506 3621 -486 3641
rect -545 3119 -525 3139
rect -506 3119 -486 3139
rect -545 2617 -525 2637
rect -506 2617 -486 2637
rect -545 2115 -525 2135
rect -506 2115 -486 2135
rect -545 1613 -525 1633
rect -506 1613 -486 1633
rect -545 1111 -525 1131
rect -506 1111 -486 1131
rect -545 609 -525 629
rect -506 609 -486 629
rect -545 107 -525 127
rect -506 107 -486 127
rect -434 8937 -414 8957
rect -395 8937 -375 8957
rect -356 8937 -336 8957
rect -317 8937 -297 8957
rect -434 8895 -414 8915
rect -395 8895 -375 8915
rect -356 8895 -336 8915
rect -317 8895 -297 8915
rect -434 8767 -414 8787
rect -395 8767 -375 8787
rect -356 8767 -336 8787
rect -317 8767 -297 8787
rect -434 8435 -414 8455
rect -395 8435 -375 8455
rect -356 8435 -336 8455
rect -317 8435 -297 8455
rect -434 7933 -414 7953
rect -395 7933 -375 7953
rect -356 7933 -336 7953
rect -317 7933 -297 7953
rect -434 7431 -414 7451
rect -395 7431 -375 7451
rect -356 7431 -336 7451
rect -317 7431 -297 7451
rect -434 6929 -414 6949
rect -395 6929 -375 6949
rect -356 6929 -336 6949
rect -317 6929 -297 6949
rect -434 6427 -414 6447
rect -395 6427 -375 6447
rect -356 6427 -336 6447
rect -317 6427 -297 6447
rect -434 5925 -414 5945
rect -395 5925 -375 5945
rect -356 5925 -336 5945
rect -317 5925 -297 5945
rect -434 5423 -414 5443
rect -395 5423 -375 5443
rect -356 5423 -336 5443
rect -317 5423 -297 5443
rect -434 4921 -414 4941
rect -395 4921 -375 4941
rect -356 4921 -336 4941
rect -317 4921 -297 4941
rect -434 4419 -414 4439
rect -395 4419 -375 4439
rect -356 4419 -336 4439
rect -317 4419 -297 4439
rect -434 3917 -414 3937
rect -395 3917 -375 3937
rect -356 3917 -336 3937
rect -317 3917 -297 3937
rect -434 3415 -414 3435
rect -395 3415 -375 3435
rect -356 3415 -336 3435
rect -317 3415 -297 3435
rect -434 2913 -414 2933
rect -395 2913 -375 2933
rect -356 2913 -336 2933
rect -317 2913 -297 2933
rect -434 2411 -414 2431
rect -395 2411 -375 2431
rect -356 2411 -336 2431
rect -317 2411 -297 2431
rect -434 1909 -414 1929
rect -395 1909 -375 1929
rect -356 1909 -336 1929
rect -317 1909 -297 1929
rect -434 1407 -414 1427
rect -395 1407 -375 1427
rect -356 1407 -336 1427
rect -317 1407 -297 1427
rect -434 905 -414 925
rect -395 905 -375 925
rect -356 905 -336 925
rect -317 905 -297 925
rect -434 403 -414 423
rect -395 403 -375 423
rect -356 403 -336 423
rect -317 403 -297 423
rect -434 361 -414 381
rect -395 361 -375 381
rect -356 361 -336 381
rect -317 361 -297 381
rect -430 -332 -402 -304
rect -383 -332 -355 -304
rect -336 -332 -308 -304
rect -430 -379 -402 -351
rect -383 -379 -355 -351
rect -336 -379 -308 -351
rect -430 -426 -402 -398
rect -383 -426 -355 -398
rect -336 -426 -308 -398
rect -241 9236 -213 9264
rect -194 9236 -166 9264
rect -147 9236 -119 9264
rect -241 9189 -213 9217
rect -194 9189 -166 9217
rect -147 9189 -119 9217
rect -241 9142 -213 9170
rect -194 9142 -166 9170
rect -147 9142 -119 9170
rect 302 9236 330 9264
rect 349 9236 377 9264
rect 396 9236 424 9264
rect 302 9189 330 9217
rect 349 9189 377 9217
rect 396 9189 424 9217
rect 302 9142 330 9170
rect 349 9142 377 9170
rect 396 9142 424 9170
rect 652 9236 680 9264
rect 699 9236 727 9264
rect 746 9236 774 9264
rect 652 9189 680 9217
rect 699 9189 727 9217
rect 746 9189 774 9217
rect 652 9142 680 9170
rect 699 9142 727 9170
rect 746 9142 774 9170
rect 1863 9516 1994 9595
rect 1866 9236 1894 9264
rect 1913 9236 1941 9264
rect 1960 9236 1988 9264
rect 1866 9189 1894 9217
rect 1913 9189 1941 9217
rect 1960 9189 1988 9217
rect 1866 9142 1894 9170
rect 1913 9142 1941 9170
rect 1960 9142 1988 9170
rect 2299 9516 2430 9595
rect 2302 9236 2330 9264
rect 2349 9236 2377 9264
rect 2396 9236 2424 9264
rect 2302 9189 2330 9217
rect 2349 9189 2377 9217
rect 2396 9189 2424 9217
rect 2302 9142 2330 9170
rect 2349 9142 2377 9170
rect 2396 9142 2424 9170
rect 2652 9236 2680 9264
rect 2699 9236 2727 9264
rect 2746 9236 2774 9264
rect 2652 9189 2680 9217
rect 2699 9189 2727 9217
rect 2746 9189 2774 9217
rect 2652 9142 2680 9170
rect 2699 9142 2727 9170
rect 2746 9142 2774 9170
rect 3863 9516 3994 9595
rect 3866 9236 3894 9264
rect 3913 9236 3941 9264
rect 3960 9236 3988 9264
rect 3866 9189 3894 9217
rect 3913 9189 3941 9217
rect 3960 9189 3988 9217
rect 3866 9142 3894 9170
rect 3913 9142 3941 9170
rect 3960 9142 3988 9170
rect 4299 9516 4430 9595
rect 4302 9236 4330 9264
rect 4349 9236 4377 9264
rect 4396 9236 4424 9264
rect 4302 9189 4330 9217
rect 4349 9189 4377 9217
rect 4396 9189 4424 9217
rect 4302 9142 4330 9170
rect 4349 9142 4377 9170
rect 4396 9142 4424 9170
rect 4652 9236 4680 9264
rect 4699 9236 4727 9264
rect 4746 9236 4774 9264
rect 4652 9189 4680 9217
rect 4699 9189 4727 9217
rect 4746 9189 4774 9217
rect 4652 9142 4680 9170
rect 4699 9142 4727 9170
rect 4746 9142 4774 9170
rect 5863 9516 5994 9595
rect 5866 9236 5894 9264
rect 5913 9236 5941 9264
rect 5960 9236 5988 9264
rect 5866 9189 5894 9217
rect 5913 9189 5941 9217
rect 5960 9189 5988 9217
rect 5866 9142 5894 9170
rect 5913 9142 5941 9170
rect 5960 9142 5988 9170
rect 6299 9516 6430 9595
rect 6302 9236 6330 9264
rect 6349 9236 6377 9264
rect 6396 9236 6424 9264
rect 6302 9189 6330 9217
rect 6349 9189 6377 9217
rect 6396 9189 6424 9217
rect 6302 9142 6330 9170
rect 6349 9142 6377 9170
rect 6396 9142 6424 9170
rect 6652 9236 6680 9264
rect 6699 9236 6727 9264
rect 6746 9236 6774 9264
rect 6652 9189 6680 9217
rect 6699 9189 6727 9217
rect 6746 9189 6774 9217
rect 6652 9142 6680 9170
rect 6699 9142 6727 9170
rect 6746 9142 6774 9170
rect 7863 9516 7994 9595
rect 7866 9236 7894 9264
rect 7913 9236 7941 9264
rect 7960 9236 7988 9264
rect 7866 9189 7894 9217
rect 7913 9189 7941 9217
rect 7960 9189 7988 9217
rect 7866 9142 7894 9170
rect 7913 9142 7941 9170
rect 7960 9142 7988 9170
rect 8299 9516 8430 9595
rect 8302 9236 8330 9264
rect 8349 9236 8377 9264
rect 8396 9236 8424 9264
rect 8302 9189 8330 9217
rect 8349 9189 8377 9217
rect 8396 9189 8424 9217
rect 8302 9142 8330 9170
rect 8349 9142 8377 9170
rect 8396 9142 8424 9170
rect 8652 9236 8680 9264
rect 8699 9236 8727 9264
rect 8746 9236 8774 9264
rect 8652 9189 8680 9217
rect 8699 9189 8727 9217
rect 8746 9189 8774 9217
rect 8652 9142 8680 9170
rect 8699 9142 8727 9170
rect 8746 9142 8774 9170
rect 9863 9516 9994 9595
rect 9866 9236 9894 9264
rect 9913 9236 9941 9264
rect 9960 9236 9988 9264
rect 9866 9189 9894 9217
rect 9913 9189 9941 9217
rect 9960 9189 9988 9217
rect 9866 9142 9894 9170
rect 9913 9142 9941 9170
rect 9960 9142 9988 9170
rect 10299 9516 10430 9595
rect 10302 9236 10330 9264
rect 10349 9236 10377 9264
rect 10396 9236 10424 9264
rect 10302 9189 10330 9217
rect 10349 9189 10377 9217
rect 10396 9189 10424 9217
rect 10302 9142 10330 9170
rect 10349 9142 10377 9170
rect 10396 9142 10424 9170
rect 10652 9236 10680 9264
rect 10699 9236 10727 9264
rect 10746 9236 10774 9264
rect 10652 9189 10680 9217
rect 10699 9189 10727 9217
rect 10746 9189 10774 9217
rect 10652 9142 10680 9170
rect 10699 9142 10727 9170
rect 10746 9142 10774 9170
rect 11863 9516 11994 9595
rect 11866 9236 11894 9264
rect 11913 9236 11941 9264
rect 11960 9236 11988 9264
rect 11866 9189 11894 9217
rect 11913 9189 11941 9217
rect 11960 9189 11988 9217
rect 11866 9142 11894 9170
rect 11913 9142 11941 9170
rect 11960 9142 11988 9170
rect 12299 9516 12430 9595
rect 12302 9236 12330 9264
rect 12349 9236 12377 9264
rect 12396 9236 12424 9264
rect 12302 9189 12330 9217
rect 12349 9189 12377 9217
rect 12396 9189 12424 9217
rect 12302 9142 12330 9170
rect 12349 9142 12377 9170
rect 12396 9142 12424 9170
rect 12652 9236 12680 9264
rect 12699 9236 12727 9264
rect 12746 9236 12774 9264
rect 12652 9189 12680 9217
rect 12699 9189 12727 9217
rect 12746 9189 12774 9217
rect 12652 9142 12680 9170
rect 12699 9142 12727 9170
rect 12746 9142 12774 9170
rect 13863 9516 13994 9595
rect 13866 9236 13894 9264
rect 13913 9236 13941 9264
rect 13960 9236 13988 9264
rect 13866 9189 13894 9217
rect 13913 9189 13941 9217
rect 13960 9189 13988 9217
rect 13866 9142 13894 9170
rect 13913 9142 13941 9170
rect 13960 9142 13988 9170
rect 14299 9516 14430 9595
rect 14302 9236 14330 9264
rect 14349 9236 14377 9264
rect 14396 9236 14424 9264
rect 14302 9189 14330 9217
rect 14349 9189 14377 9217
rect 14396 9189 14424 9217
rect 14302 9142 14330 9170
rect 14349 9142 14377 9170
rect 14396 9142 14424 9170
rect 14652 9236 14680 9264
rect 14699 9236 14727 9264
rect 14746 9236 14774 9264
rect 14652 9189 14680 9217
rect 14699 9189 14727 9217
rect 14746 9189 14774 9217
rect 14652 9142 14680 9170
rect 14699 9142 14727 9170
rect 14746 9142 14774 9170
rect 15863 9516 15994 9595
rect 15866 9236 15894 9264
rect 15913 9236 15941 9264
rect 15960 9236 15988 9264
rect 15866 9189 15894 9217
rect 15913 9189 15941 9217
rect 15960 9189 15988 9217
rect 15866 9142 15894 9170
rect 15913 9142 15941 9170
rect 15960 9142 15988 9170
rect 16299 9516 16430 9595
rect 16302 9236 16330 9264
rect 16349 9236 16377 9264
rect 16396 9236 16424 9264
rect 16302 9189 16330 9217
rect 16349 9189 16377 9217
rect 16396 9189 16424 9217
rect 16302 9142 16330 9170
rect 16349 9142 16377 9170
rect 16396 9142 16424 9170
rect 17863 9533 17994 9595
rect 16652 9236 16680 9264
rect 16699 9236 16727 9264
rect 16746 9236 16774 9264
rect 16652 9189 16680 9217
rect 16699 9189 16727 9217
rect 16746 9189 16774 9217
rect 16652 9142 16680 9170
rect 16699 9142 16727 9170
rect 16746 9142 16774 9170
rect 17181 9231 17209 9259
rect 17228 9231 17256 9259
rect 17275 9231 17303 9259
rect 17181 9184 17209 9212
rect 17228 9184 17256 9212
rect 17275 9184 17303 9212
rect 17181 9137 17209 9165
rect 17228 9137 17256 9165
rect 17275 9137 17303 9165
rect -245 8711 -225 8731
rect -206 8711 -186 8731
rect -167 8711 -147 8731
rect -128 8711 -108 8731
rect -245 8606 -225 8626
rect -206 8606 -186 8626
rect -167 8606 -147 8626
rect -128 8606 -108 8626
rect -245 8104 -225 8124
rect -206 8104 -186 8124
rect -167 8104 -147 8124
rect -128 8104 -108 8124
rect -245 7602 -225 7622
rect -206 7602 -186 7622
rect -167 7602 -147 7622
rect -128 7602 -108 7622
rect -245 7100 -225 7120
rect -206 7100 -186 7120
rect -167 7100 -147 7120
rect -128 7100 -108 7120
rect -245 6598 -225 6618
rect -206 6598 -186 6618
rect -167 6598 -147 6618
rect -128 6598 -108 6618
rect -245 6096 -225 6116
rect -206 6096 -186 6116
rect -167 6096 -147 6116
rect -128 6096 -108 6116
rect -245 5594 -225 5614
rect -206 5594 -186 5614
rect -167 5594 -147 5614
rect -128 5594 -108 5614
rect -245 5092 -225 5112
rect -206 5092 -186 5112
rect -167 5092 -147 5112
rect -128 5092 -108 5112
rect -245 4590 -225 4610
rect -206 4590 -186 4610
rect -167 4590 -147 4610
rect -128 4590 -108 4610
rect -245 4088 -225 4108
rect -206 4088 -186 4108
rect -167 4088 -147 4108
rect -128 4088 -108 4108
rect -245 3586 -225 3606
rect -206 3586 -186 3606
rect -167 3586 -147 3606
rect -128 3586 -108 3606
rect -245 3084 -225 3104
rect -206 3084 -186 3104
rect -167 3084 -147 3104
rect -128 3084 -108 3104
rect -245 2582 -225 2602
rect -206 2582 -186 2602
rect -167 2582 -147 2602
rect -128 2582 -108 2602
rect -245 2080 -225 2100
rect -206 2080 -186 2100
rect -167 2080 -147 2100
rect -128 2080 -108 2100
rect -245 1578 -225 1598
rect -206 1578 -186 1598
rect -167 1578 -147 1598
rect -128 1578 -108 1598
rect -245 1076 -225 1096
rect -206 1076 -186 1096
rect -167 1076 -147 1096
rect -128 1076 -108 1096
rect 17182 8837 17210 8865
rect 17229 8837 17257 8865
rect 17276 8837 17304 8865
rect 17182 8790 17210 8818
rect 17229 8790 17257 8818
rect 17276 8790 17304 8818
rect 17182 8743 17210 8771
rect 17229 8743 17257 8771
rect 17276 8743 17304 8771
rect 17170 8606 17190 8626
rect 17209 8606 17229 8626
rect 17248 8606 17268 8626
rect 17287 8606 17307 8626
rect 17170 8104 17190 8124
rect 17209 8104 17229 8124
rect 17248 8104 17268 8124
rect 17287 8104 17307 8124
rect 17181 7829 17209 7857
rect 17228 7829 17256 7857
rect 17275 7829 17303 7857
rect 17181 7782 17209 7810
rect 17228 7782 17256 7810
rect 17275 7782 17303 7810
rect 17181 7735 17209 7763
rect 17228 7735 17256 7763
rect 17275 7735 17303 7763
rect 17170 7602 17190 7622
rect 17209 7602 17229 7622
rect 17248 7602 17268 7622
rect 17287 7602 17307 7622
rect 17170 7100 17190 7120
rect 17209 7100 17229 7120
rect 17248 7100 17268 7120
rect 17287 7100 17307 7120
rect 17181 6829 17209 6857
rect 17228 6829 17256 6857
rect 17275 6829 17303 6857
rect 17181 6782 17209 6810
rect 17228 6782 17256 6810
rect 17275 6782 17303 6810
rect 17181 6735 17209 6763
rect 17228 6735 17256 6763
rect 17275 6735 17303 6763
rect 17170 6598 17190 6618
rect 17209 6598 17229 6618
rect 17248 6598 17268 6618
rect 17287 6598 17307 6618
rect 17370 9450 17398 9478
rect 17417 9450 17445 9478
rect 17464 9450 17492 9478
rect 17370 9403 17398 9431
rect 17417 9403 17445 9431
rect 17464 9403 17492 9431
rect 17370 9356 17398 9384
rect 17417 9356 17445 9384
rect 17464 9356 17492 9384
rect 17866 9236 17894 9264
rect 17913 9236 17941 9264
rect 17960 9236 17988 9264
rect 17866 9189 17894 9217
rect 17913 9189 17941 9217
rect 17960 9189 17988 9217
rect 17866 9142 17894 9170
rect 17913 9142 17941 9170
rect 17960 9142 17988 9170
rect 17359 8937 17379 8957
rect 17398 8937 17418 8957
rect 17437 8937 17457 8957
rect 17476 8937 17496 8957
rect 17359 8435 17379 8455
rect 17398 8435 17418 8455
rect 17437 8435 17457 8455
rect 17476 8435 17496 8455
rect 17370 8345 17398 8373
rect 17417 8345 17445 8373
rect 17464 8345 17492 8373
rect 17370 8298 17398 8326
rect 17417 8298 17445 8326
rect 17464 8298 17492 8326
rect 17370 8251 17398 8279
rect 17417 8251 17445 8279
rect 17464 8251 17492 8279
rect 17359 7933 17379 7953
rect 17398 7933 17418 7953
rect 17437 7933 17457 7953
rect 17476 7933 17496 7953
rect 17359 7431 17379 7451
rect 17398 7431 17418 7451
rect 17437 7431 17457 7451
rect 17476 7431 17496 7451
rect 17370 7291 17398 7319
rect 17417 7291 17445 7319
rect 17464 7291 17492 7319
rect 17370 7244 17398 7272
rect 17417 7244 17445 7272
rect 17464 7244 17492 7272
rect 17370 7197 17398 7225
rect 17417 7197 17445 7225
rect 17464 7197 17492 7225
rect 17359 6929 17379 6949
rect 17398 6929 17418 6949
rect 17437 6929 17457 6949
rect 17476 6929 17496 6949
rect 17359 6427 17379 6447
rect 17398 6427 17418 6447
rect 17437 6427 17457 6447
rect 17476 6427 17496 6447
rect 17369 6326 17397 6354
rect 17416 6326 17444 6354
rect 17463 6326 17491 6354
rect 17369 6279 17397 6307
rect 17416 6279 17444 6307
rect 17463 6279 17491 6307
rect 17369 6232 17397 6260
rect 17416 6232 17444 6260
rect 17463 6232 17491 6260
rect 17170 6096 17190 6116
rect 17209 6096 17229 6116
rect 17248 6096 17268 6116
rect 17287 6096 17307 6116
rect 17182 5867 17210 5895
rect 17229 5867 17257 5895
rect 17276 5867 17304 5895
rect 17182 5820 17210 5848
rect 17229 5820 17257 5848
rect 17276 5820 17304 5848
rect 17182 5773 17210 5801
rect 17229 5773 17257 5801
rect 17276 5773 17304 5801
rect 17170 5594 17190 5614
rect 17209 5594 17229 5614
rect 17248 5594 17268 5614
rect 17287 5594 17307 5614
rect 17170 5092 17190 5112
rect 17209 5092 17229 5112
rect 17248 5092 17268 5112
rect 17287 5092 17307 5112
rect 17181 4804 17209 4832
rect 17228 4804 17256 4832
rect 17275 4804 17303 4832
rect 17181 4757 17209 4785
rect 17228 4757 17256 4785
rect 17275 4757 17303 4785
rect 17181 4710 17209 4738
rect 17228 4710 17256 4738
rect 17275 4710 17303 4738
rect 17170 4590 17190 4610
rect 17209 4590 17229 4610
rect 17248 4590 17268 4610
rect 17287 4590 17307 4610
rect 17170 4088 17190 4108
rect 17209 4088 17229 4108
rect 17248 4088 17268 4108
rect 17287 4088 17307 4108
rect 17182 3816 17210 3844
rect 17229 3816 17257 3844
rect 17276 3816 17304 3844
rect 17182 3769 17210 3797
rect 17229 3769 17257 3797
rect 17276 3769 17304 3797
rect 17182 3722 17210 3750
rect 17229 3722 17257 3750
rect 17276 3722 17304 3750
rect 17170 3586 17190 3606
rect 17209 3586 17229 3606
rect 17248 3586 17268 3606
rect 17287 3586 17307 3606
rect 17359 5925 17379 5945
rect 17398 5925 17418 5945
rect 17437 5925 17457 5945
rect 17476 5925 17496 5945
rect 17548 8641 17568 8661
rect 17587 8641 17607 8661
rect 17548 8139 17568 8159
rect 17587 8139 17607 8159
rect 17548 7637 17568 7657
rect 17587 7637 17607 7657
rect 17548 7135 17568 7155
rect 17587 7135 17607 7155
rect 17548 6633 17568 6653
rect 17587 6633 17607 6653
rect 17548 6131 17568 6151
rect 17587 6131 17607 6151
rect 17359 5423 17379 5443
rect 17398 5423 17418 5443
rect 17437 5423 17457 5443
rect 17476 5423 17496 5443
rect 17370 5318 17398 5346
rect 17417 5318 17445 5346
rect 17464 5318 17492 5346
rect 17370 5271 17398 5299
rect 17417 5271 17445 5299
rect 17464 5271 17492 5299
rect 17370 5224 17398 5252
rect 17417 5224 17445 5252
rect 17464 5224 17492 5252
rect 17359 4921 17379 4941
rect 17398 4921 17418 4941
rect 17437 4921 17457 4941
rect 17476 4921 17496 4941
rect 17359 4419 17379 4439
rect 17398 4419 17418 4439
rect 17437 4419 17457 4439
rect 17476 4419 17496 4439
rect 17370 4317 17398 4345
rect 17417 4317 17445 4345
rect 17464 4317 17492 4345
rect 17370 4270 17398 4298
rect 17417 4270 17445 4298
rect 17464 4270 17492 4298
rect 17370 4223 17398 4251
rect 17417 4223 17445 4251
rect 17464 4223 17492 4251
rect 17359 3917 17379 3937
rect 17398 3917 17418 3937
rect 17437 3917 17457 3937
rect 17476 3917 17496 3937
rect 17548 5629 17568 5649
rect 17587 5629 17607 5649
rect 17548 5127 17568 5147
rect 17587 5127 17607 5147
rect 17548 4625 17568 4645
rect 17587 4625 17607 4645
rect 17548 4123 17568 4143
rect 17587 4123 17607 4143
rect 17359 3415 17379 3435
rect 17398 3415 17418 3435
rect 17437 3415 17457 3435
rect 17476 3415 17496 3435
rect 17369 3318 17397 3346
rect 17416 3318 17444 3346
rect 17463 3318 17491 3346
rect 17369 3271 17397 3299
rect 17416 3271 17444 3299
rect 17463 3271 17491 3299
rect 17369 3224 17397 3252
rect 17416 3224 17444 3252
rect 17463 3224 17491 3252
rect 17170 3084 17190 3104
rect 17209 3084 17229 3104
rect 17248 3084 17268 3104
rect 17287 3084 17307 3104
rect 17182 2794 17210 2822
rect 17229 2794 17257 2822
rect 17276 2794 17304 2822
rect 17182 2747 17210 2775
rect 17229 2747 17257 2775
rect 17276 2747 17304 2775
rect 17182 2700 17210 2728
rect 17229 2700 17257 2728
rect 17276 2700 17304 2728
rect 17170 2582 17190 2602
rect 17209 2582 17229 2602
rect 17248 2582 17268 2602
rect 17287 2582 17307 2602
rect 17170 2080 17190 2100
rect 17209 2080 17229 2100
rect 17248 2080 17268 2100
rect 17287 2080 17307 2100
rect 17182 1797 17210 1825
rect 17229 1797 17257 1825
rect 17276 1797 17304 1825
rect 17182 1750 17210 1778
rect 17229 1750 17257 1778
rect 17276 1750 17304 1778
rect 17182 1703 17210 1731
rect 17229 1703 17257 1731
rect 17276 1703 17304 1731
rect 17170 1578 17190 1598
rect 17209 1578 17229 1598
rect 17248 1578 17268 1598
rect 17287 1578 17307 1598
rect 17170 1076 17190 1096
rect 17209 1076 17229 1096
rect 17248 1076 17268 1096
rect 17287 1076 17307 1096
rect 17359 2913 17379 2933
rect 17398 2913 17418 2933
rect 17437 2913 17457 2933
rect 17476 2913 17496 2933
rect 17548 3621 17568 3641
rect 17587 3621 17607 3641
rect 17548 3119 17568 3139
rect 17587 3119 17607 3139
rect 17359 2411 17379 2431
rect 17398 2411 17418 2431
rect 17437 2411 17457 2431
rect 17476 2411 17496 2431
rect 17370 2284 17398 2312
rect 17417 2284 17445 2312
rect 17464 2284 17492 2312
rect 17370 2237 17398 2265
rect 17417 2237 17445 2265
rect 17464 2237 17492 2265
rect 17370 2190 17398 2218
rect 17417 2190 17445 2218
rect 17464 2190 17492 2218
rect 17359 1909 17379 1929
rect 17398 1909 17418 1929
rect 17437 1909 17457 1929
rect 17476 1909 17496 1929
rect 17548 2617 17568 2637
rect 17587 2617 17607 2637
rect 17548 2115 17568 2135
rect 17587 2115 17607 2135
rect 17359 1407 17379 1427
rect 17398 1407 17418 1427
rect 17437 1407 17457 1427
rect 17476 1407 17496 1427
rect 17370 1282 17398 1310
rect 17417 1282 17445 1310
rect 17464 1282 17492 1310
rect 17370 1235 17398 1263
rect 17417 1235 17445 1263
rect 17464 1235 17492 1263
rect 17370 1188 17398 1216
rect 17417 1188 17445 1216
rect 17464 1188 17492 1216
rect 17359 905 17379 925
rect 17398 905 17418 925
rect 17437 905 17457 925
rect 17476 905 17496 925
rect 17180 797 17208 825
rect 17227 797 17255 825
rect 17274 797 17302 825
rect 17180 750 17208 778
rect 17227 750 17255 778
rect 17274 750 17302 778
rect 17180 703 17208 731
rect 17227 703 17255 731
rect 17274 703 17302 731
rect -245 574 -225 594
rect -206 574 -186 594
rect -167 574 -147 594
rect -128 574 -108 594
rect -245 233 -225 253
rect -206 233 -186 253
rect -167 233 -147 253
rect -128 233 -108 253
rect -245 177 -225 197
rect -206 177 -186 197
rect -167 177 -147 197
rect -128 177 -108 197
rect -245 72 -225 92
rect -206 72 -186 92
rect -167 72 -147 92
rect -128 72 -108 92
rect 17170 574 17190 594
rect 17209 574 17229 594
rect 17248 574 17268 594
rect 17287 574 17307 594
rect 17170 72 17190 92
rect 17209 72 17229 92
rect 17248 72 17268 92
rect 17287 72 17307 92
rect -241 -113 -213 -85
rect -194 -113 -166 -85
rect -147 -113 -119 -85
rect -241 -160 -213 -132
rect -194 -160 -166 -132
rect -147 -160 -119 -132
rect -241 -207 -213 -179
rect -194 -207 -166 -179
rect -147 -207 -119 -179
rect 425 -312 442 -295
rect 13283 -153 13300 -136
rect 14483 -153 14500 -136
rect 13385 -192 13402 -175
rect 14985 -192 15002 -175
rect 13487 -230 13504 -213
rect 15487 -230 15504 -213
rect 13589 -268 13606 -251
rect 15989 -268 16006 -251
rect 13691 -306 13708 -289
rect 16104 -81 16121 -64
rect 16348 -81 16365 -64
rect 16491 -306 16508 -289
rect 17181 -48 17209 -20
rect 17228 -48 17256 -20
rect 17275 -48 17303 -20
rect 17181 -95 17209 -67
rect 17228 -95 17256 -67
rect 17275 -95 17303 -67
rect 17181 -142 17209 -114
rect 17228 -142 17256 -114
rect 17275 -142 17303 -114
rect 16995 -315 17012 -298
rect 17359 403 17379 423
rect 17398 403 17418 423
rect 17437 403 17457 423
rect 17476 403 17496 423
rect 17370 285 17398 313
rect 17417 285 17445 313
rect 17464 285 17492 313
rect 17370 238 17398 266
rect 17417 238 17445 266
rect 17464 238 17492 266
rect 17370 191 17398 219
rect 17417 191 17445 219
rect 17464 191 17492 219
rect 17548 1613 17568 1633
rect 17587 1613 17607 1633
rect 17548 1111 17568 1131
rect 17587 1111 17607 1131
rect 17650 8853 17825 8870
rect 17650 8413 17825 8430
rect 17650 7973 17825 7990
rect 17650 7533 17825 7550
rect 17650 7093 17825 7110
rect 17650 6653 17825 6670
rect 20448 8962 20554 9168
rect 20448 8083 20554 8289
rect 20448 6962 20554 7168
rect 17650 5773 17825 5790
rect 17650 4893 17825 4910
rect 17650 4453 17825 4470
rect 17650 4013 17825 4030
rect 17650 3573 17825 3590
rect 20448 6083 20554 6289
rect 20448 4962 20554 5168
rect 20448 4083 20554 4289
rect 17650 3133 17825 3150
rect 17650 2693 17825 2710
rect 17650 1813 17825 1830
rect 17650 1373 17825 1390
rect 17650 933 17825 950
rect 17548 609 17568 629
rect 17587 609 17607 629
rect 17548 107 17568 127
rect 17587 107 17607 127
rect 17650 493 17825 510
rect 17650 53 17825 70
rect 17370 -266 17398 -238
rect 17417 -266 17445 -238
rect 17464 -266 17492 -238
rect 17370 -313 17398 -285
rect 17417 -313 17445 -285
rect 17464 -313 17492 -285
rect 17370 -360 17398 -332
rect 17417 -360 17445 -332
rect 17464 -360 17492 -332
rect 20448 2962 20554 3168
rect 20448 2083 20554 2289
rect 20448 962 20554 1168
rect 20448 83 20554 289
rect 16401 -449 16418 -432
rect 16437 -449 16454 -432
<< metal1 >>
rect 20151 11371 20567 11377
rect 20151 11290 20442 11371
rect 20561 11290 20567 11371
rect 20151 11285 20567 11290
rect 20435 11168 20567 11181
rect 20435 10962 20448 11168
rect 20554 10962 20567 11168
rect 20435 10950 20567 10962
rect 20151 10937 20319 10946
rect 20151 10862 20202 10937
rect 20308 10862 20319 10937
rect 20151 10855 20319 10862
rect 20151 10666 20319 10675
rect 20151 10591 20202 10666
rect 20308 10591 20319 10666
rect 20151 10584 20319 10591
rect 20151 10388 20319 10397
rect 20151 10313 20202 10388
rect 20308 10313 20319 10388
rect 20151 10306 20319 10313
rect 20435 10289 20567 10302
rect 20435 10083 20448 10289
rect 20554 10083 20567 10289
rect 20435 10071 20567 10083
rect 20151 9816 20567 9822
rect 20151 9735 20442 9816
rect 20561 9735 20567 9816
rect 20151 9730 20567 9735
rect 292 9595 438 9626
rect 292 9516 299 9595
rect 430 9516 438 9595
rect 292 9510 438 9516
rect 1060 9493 1245 9626
rect 1856 9595 2002 9626
rect 1856 9516 1863 9595
rect 1994 9516 2002 9595
rect 1856 9510 2002 9516
rect 2292 9595 2438 9626
rect 2292 9516 2299 9595
rect 2430 9516 2438 9595
rect 2292 9510 2438 9516
rect 3060 9493 3245 9626
rect 3856 9595 4002 9626
rect 3856 9516 3863 9595
rect 3994 9516 4002 9595
rect 3856 9510 4002 9516
rect 4292 9595 4438 9626
rect 4292 9516 4299 9595
rect 4430 9516 4438 9595
rect 4292 9510 4438 9516
rect 5060 9493 5245 9626
rect 5856 9595 6002 9626
rect 5856 9516 5863 9595
rect 5994 9516 6002 9595
rect 5856 9510 6002 9516
rect 6292 9595 6438 9626
rect 6292 9516 6299 9595
rect 6430 9516 6438 9595
rect 6292 9510 6438 9516
rect 7060 9493 7245 9626
rect 7856 9595 8002 9626
rect 7856 9516 7863 9595
rect 7994 9516 8002 9595
rect 7856 9510 8002 9516
rect 8292 9595 8438 9626
rect 8292 9516 8299 9595
rect 8430 9516 8438 9595
rect 8292 9510 8438 9516
rect 9060 9493 9245 9626
rect 9856 9595 10002 9626
rect 9856 9516 9863 9595
rect 9994 9516 10002 9595
rect 9856 9510 10002 9516
rect 10292 9595 10438 9626
rect 10292 9516 10299 9595
rect 10430 9516 10438 9595
rect 10292 9510 10438 9516
rect 11060 9493 11245 9626
rect 11856 9595 12002 9626
rect 11856 9516 11863 9595
rect 11994 9516 12002 9595
rect 11856 9510 12002 9516
rect 12292 9595 12438 9626
rect 12292 9516 12299 9595
rect 12430 9516 12438 9595
rect 12292 9510 12438 9516
rect 13060 9493 13245 9626
rect 13856 9595 14002 9626
rect 13856 9516 13863 9595
rect 13994 9516 14002 9595
rect 13856 9510 14002 9516
rect 14292 9595 14438 9626
rect 14292 9516 14299 9595
rect 14430 9516 14438 9595
rect 14292 9510 14438 9516
rect 15060 9493 15245 9626
rect 15856 9595 16002 9626
rect 15856 9516 15863 9595
rect 15994 9516 16002 9595
rect 15856 9510 16002 9516
rect 16292 9595 16438 9626
rect 16292 9516 16299 9595
rect 16430 9516 16438 9595
rect 16292 9510 16438 9516
rect 17060 9493 17245 9626
rect 17856 9595 18002 9626
rect 17856 9533 17863 9595
rect 17994 9533 18002 9595
rect 17856 9527 18002 9533
rect -1195 9489 18077 9493
rect -1195 9457 -1180 9489
rect -1148 9457 -1136 9489
rect -1104 9457 -1092 9489
rect -1060 9457 -1048 9489
rect -1016 9484 17898 9489
rect -1016 9483 1072 9484
rect -1016 9457 -430 9483
rect -1195 9455 -430 9457
rect -402 9455 -383 9483
rect -355 9455 -336 9483
rect -308 9455 1072 9483
rect -1195 9444 1072 9455
rect -1195 9412 -1180 9444
rect -1148 9412 -1136 9444
rect -1104 9412 -1092 9444
rect -1060 9412 -1048 9444
rect -1016 9436 1072 9444
rect -1016 9412 -430 9436
rect -1195 9408 -430 9412
rect -402 9408 -383 9436
rect -355 9408 -336 9436
rect -308 9408 1072 9436
rect -1195 9399 1072 9408
rect -1195 9367 -1180 9399
rect -1148 9367 -1136 9399
rect -1104 9367 -1092 9399
rect -1060 9367 -1048 9399
rect -1016 9389 1072 9399
rect -1016 9367 -430 9389
rect -1195 9361 -430 9367
rect -402 9361 -383 9389
rect -355 9361 -336 9389
rect -308 9362 1072 9389
rect 1235 9362 3072 9484
rect 3235 9362 5072 9484
rect 5235 9362 7072 9484
rect 7235 9362 9072 9484
rect 9235 9362 11072 9484
rect 11235 9362 13072 9484
rect 13235 9362 15072 9484
rect 15235 9362 17072 9484
rect 17235 9478 17898 9484
rect 17235 9450 17370 9478
rect 17398 9450 17417 9478
rect 17445 9450 17464 9478
rect 17492 9457 17898 9478
rect 17930 9457 17942 9489
rect 17974 9457 17986 9489
rect 18018 9457 18030 9489
rect 18062 9457 18077 9489
rect 17492 9450 18077 9457
rect 17235 9444 18077 9450
rect 17235 9431 17898 9444
rect 17235 9403 17370 9431
rect 17398 9403 17417 9431
rect 17445 9403 17464 9431
rect 17492 9412 17898 9431
rect 17930 9412 17942 9444
rect 17974 9412 17986 9444
rect 18018 9412 18030 9444
rect 18062 9412 18077 9444
rect 17492 9403 18077 9412
rect 17235 9399 18077 9403
rect 17235 9384 17898 9399
rect 17235 9362 17370 9384
rect -308 9361 17370 9362
rect -1195 9356 17370 9361
rect 17398 9356 17417 9384
rect 17445 9356 17464 9384
rect 17492 9367 17898 9384
rect 17930 9367 17942 9399
rect 17974 9367 17986 9399
rect 18018 9367 18030 9399
rect 18062 9367 18077 9399
rect 17492 9356 18077 9367
rect -1195 9353 18077 9356
rect 20151 9371 20567 9377
rect 17166 9348 17502 9353
rect 20151 9290 20442 9371
rect 20561 9290 20567 9371
rect 20151 9285 20567 9290
rect -957 9270 18077 9274
rect -957 9238 -942 9270
rect -910 9238 -898 9270
rect -866 9238 -854 9270
rect -822 9238 -810 9270
rect -778 9264 17660 9270
rect -778 9238 -241 9264
rect -957 9236 -241 9238
rect -213 9236 -194 9264
rect -166 9236 -147 9264
rect -119 9236 302 9264
rect 330 9236 349 9264
rect 377 9236 396 9264
rect 424 9236 652 9264
rect 680 9236 699 9264
rect 727 9236 746 9264
rect 774 9236 1866 9264
rect 1894 9236 1913 9264
rect 1941 9236 1960 9264
rect 1988 9236 2302 9264
rect 2330 9236 2349 9264
rect 2377 9236 2396 9264
rect 2424 9236 2652 9264
rect 2680 9236 2699 9264
rect 2727 9236 2746 9264
rect 2774 9236 3866 9264
rect 3894 9236 3913 9264
rect 3941 9236 3960 9264
rect 3988 9236 4302 9264
rect 4330 9236 4349 9264
rect 4377 9236 4396 9264
rect 4424 9236 4652 9264
rect 4680 9236 4699 9264
rect 4727 9236 4746 9264
rect 4774 9236 5866 9264
rect 5894 9236 5913 9264
rect 5941 9236 5960 9264
rect 5988 9236 6302 9264
rect 6330 9236 6349 9264
rect 6377 9236 6396 9264
rect 6424 9236 6652 9264
rect 6680 9236 6699 9264
rect 6727 9236 6746 9264
rect 6774 9236 7866 9264
rect 7894 9236 7913 9264
rect 7941 9236 7960 9264
rect 7988 9236 8302 9264
rect 8330 9236 8349 9264
rect 8377 9236 8396 9264
rect 8424 9236 8652 9264
rect 8680 9236 8699 9264
rect 8727 9236 8746 9264
rect 8774 9236 9866 9264
rect 9894 9236 9913 9264
rect 9941 9236 9960 9264
rect 9988 9236 10302 9264
rect 10330 9236 10349 9264
rect 10377 9236 10396 9264
rect 10424 9236 10652 9264
rect 10680 9236 10699 9264
rect 10727 9236 10746 9264
rect 10774 9236 11866 9264
rect 11894 9236 11913 9264
rect 11941 9236 11960 9264
rect 11988 9236 12302 9264
rect 12330 9236 12349 9264
rect 12377 9236 12396 9264
rect 12424 9236 12652 9264
rect 12680 9236 12699 9264
rect 12727 9236 12746 9264
rect 12774 9236 13866 9264
rect 13894 9236 13913 9264
rect 13941 9236 13960 9264
rect 13988 9236 14302 9264
rect 14330 9236 14349 9264
rect 14377 9236 14396 9264
rect 14424 9236 14652 9264
rect 14680 9236 14699 9264
rect 14727 9236 14746 9264
rect 14774 9236 15866 9264
rect 15894 9236 15913 9264
rect 15941 9236 15960 9264
rect 15988 9236 16302 9264
rect 16330 9236 16349 9264
rect 16377 9236 16396 9264
rect 16424 9236 16652 9264
rect 16680 9236 16699 9264
rect 16727 9236 16746 9264
rect 16774 9259 17660 9264
rect 16774 9236 17181 9259
rect -957 9231 17181 9236
rect 17209 9231 17228 9259
rect 17256 9231 17275 9259
rect 17303 9238 17660 9259
rect 17692 9238 17704 9270
rect 17736 9238 17748 9270
rect 17780 9238 17792 9270
rect 17824 9264 18077 9270
rect 17824 9238 17866 9264
rect 17303 9236 17866 9238
rect 17894 9236 17913 9264
rect 17941 9236 17960 9264
rect 17988 9236 18077 9264
rect 17303 9231 18077 9236
rect -957 9225 18077 9231
rect -957 9193 -942 9225
rect -910 9193 -898 9225
rect -866 9193 -854 9225
rect -822 9193 -810 9225
rect -778 9217 17660 9225
rect -778 9193 -241 9217
rect -957 9189 -241 9193
rect -213 9189 -194 9217
rect -166 9189 -147 9217
rect -119 9189 302 9217
rect 330 9189 349 9217
rect 377 9189 396 9217
rect 424 9189 652 9217
rect 680 9189 699 9217
rect 727 9189 746 9217
rect 774 9189 1866 9217
rect 1894 9189 1913 9217
rect 1941 9189 1960 9217
rect 1988 9189 2302 9217
rect 2330 9189 2349 9217
rect 2377 9189 2396 9217
rect 2424 9189 2652 9217
rect 2680 9189 2699 9217
rect 2727 9189 2746 9217
rect 2774 9189 3866 9217
rect 3894 9189 3913 9217
rect 3941 9189 3960 9217
rect 3988 9189 4302 9217
rect 4330 9189 4349 9217
rect 4377 9189 4396 9217
rect 4424 9189 4652 9217
rect 4680 9189 4699 9217
rect 4727 9189 4746 9217
rect 4774 9189 5866 9217
rect 5894 9189 5913 9217
rect 5941 9189 5960 9217
rect 5988 9189 6302 9217
rect 6330 9189 6349 9217
rect 6377 9189 6396 9217
rect 6424 9189 6652 9217
rect 6680 9189 6699 9217
rect 6727 9189 6746 9217
rect 6774 9189 7866 9217
rect 7894 9189 7913 9217
rect 7941 9189 7960 9217
rect 7988 9189 8302 9217
rect 8330 9189 8349 9217
rect 8377 9189 8396 9217
rect 8424 9189 8652 9217
rect 8680 9189 8699 9217
rect 8727 9189 8746 9217
rect 8774 9189 9866 9217
rect 9894 9189 9913 9217
rect 9941 9189 9960 9217
rect 9988 9189 10302 9217
rect 10330 9189 10349 9217
rect 10377 9189 10396 9217
rect 10424 9189 10652 9217
rect 10680 9189 10699 9217
rect 10727 9189 10746 9217
rect 10774 9189 11866 9217
rect 11894 9189 11913 9217
rect 11941 9189 11960 9217
rect 11988 9189 12302 9217
rect 12330 9189 12349 9217
rect 12377 9189 12396 9217
rect 12424 9189 12652 9217
rect 12680 9189 12699 9217
rect 12727 9189 12746 9217
rect 12774 9189 13866 9217
rect 13894 9189 13913 9217
rect 13941 9189 13960 9217
rect 13988 9189 14302 9217
rect 14330 9189 14349 9217
rect 14377 9189 14396 9217
rect 14424 9189 14652 9217
rect 14680 9189 14699 9217
rect 14727 9189 14746 9217
rect 14774 9189 15866 9217
rect 15894 9189 15913 9217
rect 15941 9189 15960 9217
rect 15988 9189 16302 9217
rect 16330 9189 16349 9217
rect 16377 9189 16396 9217
rect 16424 9189 16652 9217
rect 16680 9189 16699 9217
rect 16727 9189 16746 9217
rect 16774 9212 17660 9217
rect 16774 9189 17181 9212
rect -957 9184 17181 9189
rect 17209 9184 17228 9212
rect 17256 9184 17275 9212
rect 17303 9193 17660 9212
rect 17692 9193 17704 9225
rect 17736 9193 17748 9225
rect 17780 9193 17792 9225
rect 17824 9217 18077 9225
rect 17824 9193 17866 9217
rect 17303 9189 17866 9193
rect 17894 9189 17913 9217
rect 17941 9189 17960 9217
rect 17988 9189 18077 9217
rect 17303 9184 18077 9189
rect -957 9180 18077 9184
rect -957 9148 -942 9180
rect -910 9148 -898 9180
rect -866 9148 -854 9180
rect -822 9148 -810 9180
rect -778 9170 17660 9180
rect -778 9148 -241 9170
rect -957 9142 -241 9148
rect -213 9142 -194 9170
rect -166 9142 -147 9170
rect -119 9142 302 9170
rect 330 9142 349 9170
rect 377 9142 396 9170
rect 424 9142 652 9170
rect 680 9142 699 9170
rect 727 9142 746 9170
rect 774 9142 1866 9170
rect 1894 9142 1913 9170
rect 1941 9142 1960 9170
rect 1988 9142 2302 9170
rect 2330 9142 2349 9170
rect 2377 9142 2396 9170
rect 2424 9142 2652 9170
rect 2680 9142 2699 9170
rect 2727 9142 2746 9170
rect 2774 9142 3866 9170
rect 3894 9142 3913 9170
rect 3941 9142 3960 9170
rect 3988 9142 4302 9170
rect 4330 9142 4349 9170
rect 4377 9142 4396 9170
rect 4424 9142 4652 9170
rect 4680 9142 4699 9170
rect 4727 9142 4746 9170
rect 4774 9142 5866 9170
rect 5894 9142 5913 9170
rect 5941 9142 5960 9170
rect 5988 9142 6302 9170
rect 6330 9142 6349 9170
rect 6377 9142 6396 9170
rect 6424 9142 6652 9170
rect 6680 9142 6699 9170
rect 6727 9142 6746 9170
rect 6774 9142 7866 9170
rect 7894 9142 7913 9170
rect 7941 9142 7960 9170
rect 7988 9142 8302 9170
rect 8330 9142 8349 9170
rect 8377 9142 8396 9170
rect 8424 9142 8652 9170
rect 8680 9142 8699 9170
rect 8727 9142 8746 9170
rect 8774 9142 9866 9170
rect 9894 9142 9913 9170
rect 9941 9142 9960 9170
rect 9988 9142 10302 9170
rect 10330 9142 10349 9170
rect 10377 9142 10396 9170
rect 10424 9142 10652 9170
rect 10680 9142 10699 9170
rect 10727 9142 10746 9170
rect 10774 9142 11866 9170
rect 11894 9142 11913 9170
rect 11941 9142 11960 9170
rect 11988 9142 12302 9170
rect 12330 9142 12349 9170
rect 12377 9142 12396 9170
rect 12424 9142 12652 9170
rect 12680 9142 12699 9170
rect 12727 9142 12746 9170
rect 12774 9142 13866 9170
rect 13894 9142 13913 9170
rect 13941 9142 13960 9170
rect 13988 9142 14302 9170
rect 14330 9142 14349 9170
rect 14377 9142 14396 9170
rect 14424 9142 14652 9170
rect 14680 9142 14699 9170
rect 14727 9142 14746 9170
rect 14774 9142 15866 9170
rect 15894 9142 15913 9170
rect 15941 9142 15960 9170
rect 15988 9142 16302 9170
rect 16330 9142 16349 9170
rect 16377 9142 16396 9170
rect 16424 9142 16652 9170
rect 16680 9142 16699 9170
rect 16727 9142 16746 9170
rect 16774 9165 17660 9170
rect 16774 9142 17181 9165
rect -957 9137 17181 9142
rect 17209 9137 17228 9165
rect 17256 9137 17275 9165
rect 17303 9148 17660 9165
rect 17692 9148 17704 9180
rect 17736 9148 17748 9180
rect 17780 9148 17792 9180
rect 17824 9170 18077 9180
rect 17824 9148 17866 9170
rect 17303 9142 17866 9148
rect 17894 9142 17913 9170
rect 17941 9142 17960 9170
rect 17988 9142 18077 9170
rect 17303 9137 18077 9142
rect -957 9135 18077 9137
rect -956 9134 18077 9135
rect 20435 9168 20567 9181
rect 17166 9129 17502 9134
rect 20435 8962 20448 9168
rect 20554 8962 20567 9168
rect -440 8957 0 8961
rect -440 8937 -434 8957
rect -414 8937 -395 8957
rect -375 8937 -356 8957
rect -336 8937 -317 8957
rect -297 8937 0 8957
rect -440 8933 0 8937
rect 17068 8957 17503 8961
rect 17068 8937 17359 8957
rect 17379 8937 17398 8957
rect 17418 8937 17437 8957
rect 17457 8937 17476 8957
rect 17496 8937 17503 8957
rect 20435 8950 20567 8962
rect 17068 8933 17503 8937
rect 20151 8937 20319 8946
rect -440 8915 0 8919
rect -440 8895 -434 8915
rect -414 8895 -395 8915
rect -375 8895 -356 8915
rect -336 8895 -317 8915
rect -297 8905 0 8915
rect -297 8895 -291 8905
rect -440 8891 -291 8895
rect -949 8848 -943 8874
rect -768 8848 -762 8874
rect 17644 8873 17650 8874
rect 17168 8865 17650 8873
rect 17825 8873 17831 8874
rect 17825 8872 17839 8873
rect 17168 8837 17182 8865
rect 17210 8837 17229 8865
rect 17257 8837 17276 8865
rect 17304 8848 17650 8865
rect 17304 8837 17661 8848
rect 17168 8827 17661 8837
rect 17693 8827 17705 8848
rect 17737 8827 17749 8848
rect 17781 8827 17793 8848
rect 17825 8827 17840 8872
rect 20151 8862 20202 8937
rect 20308 8862 20319 8937
rect 20151 8855 20319 8862
rect 17168 8818 17840 8827
rect -440 8790 0 8804
rect 17168 8790 17182 8818
rect 17210 8790 17229 8818
rect 17257 8790 17276 8818
rect 17304 8814 17840 8818
rect 17304 8790 17661 8814
rect -440 8787 -291 8790
rect -440 8767 -434 8787
rect -414 8767 -395 8787
rect -375 8767 -356 8787
rect -336 8767 -317 8787
rect -297 8767 -291 8787
rect -440 8763 -291 8767
rect 17168 8782 17661 8790
rect 17693 8782 17705 8814
rect 17737 8782 17749 8814
rect 17781 8782 17793 8814
rect 17825 8782 17840 8814
rect 17168 8771 17840 8782
rect -440 8749 0 8763
rect 17168 8743 17182 8771
rect 17210 8743 17229 8771
rect 17257 8743 17276 8771
rect 17304 8769 17840 8771
rect 17304 8743 17661 8769
rect 17168 8737 17661 8743
rect 17693 8737 17705 8769
rect 17737 8737 17749 8769
rect 17781 8737 17793 8769
rect 17825 8737 17840 8769
rect -251 8731 0 8735
rect 17168 8733 17840 8737
rect -251 8711 -245 8731
rect -225 8711 -206 8731
rect -186 8711 -167 8731
rect -147 8711 -128 8731
rect -108 8721 0 8731
rect -108 8711 -102 8721
rect -251 8707 -102 8711
rect 20151 8666 20319 8675
rect -551 8661 -465 8664
rect -551 8641 -545 8661
rect -525 8641 -506 8661
rect -486 8658 -465 8661
rect 17527 8661 17613 8664
rect 17527 8658 17548 8661
rect -486 8644 0 8658
rect 17068 8644 17548 8658
rect -486 8641 -465 8644
rect -551 8638 -465 8641
rect 17527 8641 17548 8644
rect 17568 8641 17587 8661
rect 17607 8641 17613 8661
rect 17527 8638 17613 8641
rect -251 8626 0 8630
rect -251 8606 -245 8626
rect -225 8606 -206 8626
rect -186 8606 -167 8626
rect -147 8606 -128 8626
rect -108 8606 0 8626
rect -251 8602 0 8606
rect 17068 8626 17313 8630
rect 17068 8606 17170 8626
rect 17190 8606 17209 8626
rect 17229 8606 17248 8626
rect 17268 8606 17287 8626
rect 17307 8606 17313 8626
rect 17068 8602 17313 8606
rect 20151 8591 20202 8666
rect 20308 8591 20319 8666
rect 20151 8584 20319 8591
rect -440 8455 0 8459
rect -440 8435 -434 8455
rect -414 8435 -395 8455
rect -375 8435 -356 8455
rect -336 8435 -317 8455
rect -297 8435 0 8455
rect -949 8408 -943 8434
rect -768 8408 -762 8434
rect -440 8431 0 8435
rect 17068 8455 17503 8459
rect 17068 8435 17359 8455
rect 17379 8435 17398 8455
rect 17418 8435 17437 8455
rect 17457 8435 17476 8455
rect 17496 8435 17503 8455
rect 17068 8431 17503 8435
rect -659 8424 -625 8427
rect -659 8407 -651 8424
rect -634 8417 -625 8424
rect -634 8407 0 8417
rect 17644 8408 17650 8434
rect 17825 8408 17831 8434
rect -659 8403 0 8407
rect 20151 8388 20319 8397
rect 17355 8380 17503 8381
rect 17355 8373 18077 8380
rect 17355 8345 17370 8373
rect 17398 8345 17417 8373
rect 17445 8345 17464 8373
rect 17492 8366 18077 8373
rect 17492 8345 17898 8366
rect 17355 8334 17898 8345
rect 17930 8334 17942 8366
rect 17974 8334 17986 8366
rect 18018 8334 18030 8366
rect 18062 8334 18077 8366
rect 17355 8326 18077 8334
rect -673 8288 0 8302
rect 17355 8298 17370 8326
rect 17398 8298 17417 8326
rect 17445 8298 17464 8326
rect 17492 8321 18077 8326
rect 17492 8298 17898 8321
rect 17355 8289 17898 8298
rect 17930 8289 17942 8321
rect 17974 8289 17986 8321
rect 18018 8289 18030 8321
rect 18062 8289 18077 8321
rect 20151 8313 20202 8388
rect 20308 8313 20319 8388
rect 20151 8306 20319 8313
rect 17355 8279 18077 8289
rect -673 8247 0 8261
rect 17355 8251 17370 8279
rect 17398 8251 17417 8279
rect 17445 8251 17464 8279
rect 17492 8276 18077 8279
rect 17492 8251 17898 8276
rect 17355 8244 17898 8251
rect 17930 8244 17942 8276
rect 17974 8244 17986 8276
rect 18018 8244 18030 8276
rect 18062 8244 18077 8276
rect 17355 8240 18077 8244
rect 20435 8289 20567 8302
rect -605 8230 0 8233
rect -605 8213 -597 8230
rect -580 8219 0 8230
rect -580 8213 -571 8219
rect -605 8209 -571 8213
rect -551 8159 -465 8162
rect -551 8139 -545 8159
rect -525 8139 -506 8159
rect -486 8156 -465 8159
rect 17527 8159 17613 8162
rect 17527 8156 17548 8159
rect -486 8142 0 8156
rect 17068 8142 17548 8156
rect -486 8139 -465 8142
rect -551 8136 -465 8139
rect 17527 8139 17548 8142
rect 17568 8139 17587 8159
rect 17607 8139 17613 8159
rect 17527 8136 17613 8139
rect -251 8124 0 8128
rect -251 8104 -245 8124
rect -225 8104 -206 8124
rect -186 8104 -167 8124
rect -147 8104 -128 8124
rect -108 8104 0 8124
rect -251 8100 0 8104
rect 17068 8124 17313 8128
rect 17068 8104 17170 8124
rect 17190 8104 17209 8124
rect 17229 8104 17248 8124
rect 17268 8104 17287 8124
rect 17307 8104 17313 8124
rect 17068 8100 17313 8104
rect 20435 8083 20448 8289
rect 20554 8083 20567 8289
rect 20435 8071 20567 8083
rect -949 7968 -943 7994
rect -768 7968 -762 7994
rect 17644 7968 17650 7994
rect 17825 7968 17831 7994
rect -440 7953 0 7957
rect -440 7933 -434 7953
rect -414 7933 -395 7953
rect -375 7933 -356 7953
rect -336 7933 -317 7953
rect -297 7933 0 7953
rect -440 7929 0 7933
rect 17068 7953 17503 7957
rect 17068 7933 17359 7953
rect 17379 7933 17398 7953
rect 17418 7933 17437 7953
rect 17457 7933 17476 7953
rect 17496 7933 17503 7953
rect 17068 7929 17503 7933
rect -659 7922 -625 7925
rect -659 7905 -651 7922
rect -634 7915 -625 7922
rect -634 7905 0 7915
rect -659 7901 0 7905
rect 17167 7864 17838 7865
rect 17167 7857 17839 7864
rect 17167 7829 17181 7857
rect 17209 7829 17228 7857
rect 17256 7829 17275 7857
rect 17303 7851 17839 7857
rect 17303 7829 17660 7851
rect 17167 7819 17660 7829
rect 17692 7819 17704 7851
rect 17736 7819 17748 7851
rect 17780 7819 17792 7851
rect 17824 7819 17839 7851
rect 17167 7810 17839 7819
rect -673 7786 0 7800
rect 17167 7782 17181 7810
rect 17209 7782 17228 7810
rect 17256 7782 17275 7810
rect 17303 7806 17839 7810
rect 17303 7782 17660 7806
rect 17167 7774 17660 7782
rect 17692 7774 17704 7806
rect 17736 7774 17748 7806
rect 17780 7774 17792 7806
rect 17824 7774 17839 7806
rect 17167 7763 17839 7774
rect -673 7745 0 7759
rect 17167 7735 17181 7763
rect 17209 7735 17228 7763
rect 17256 7735 17275 7763
rect 17303 7761 17839 7763
rect 17303 7735 17660 7761
rect -605 7728 0 7731
rect -605 7711 -597 7728
rect -580 7717 0 7728
rect 17167 7729 17660 7735
rect 17692 7729 17704 7761
rect 17736 7729 17748 7761
rect 17780 7729 17792 7761
rect 17824 7729 17839 7761
rect 20151 7816 20567 7822
rect 20151 7735 20442 7816
rect 20561 7735 20567 7816
rect 20151 7730 20567 7735
rect 17167 7725 17839 7729
rect -580 7711 -571 7717
rect -605 7707 -571 7711
rect -551 7657 -465 7660
rect -551 7637 -545 7657
rect -525 7637 -506 7657
rect -486 7654 -465 7657
rect 17527 7657 17613 7660
rect 17527 7654 17548 7657
rect -486 7640 0 7654
rect 17068 7640 17548 7654
rect -486 7637 -465 7640
rect -551 7634 -465 7637
rect 17527 7637 17548 7640
rect 17568 7637 17587 7657
rect 17607 7637 17613 7657
rect 17527 7634 17613 7637
rect -251 7622 0 7626
rect -251 7602 -245 7622
rect -225 7602 -206 7622
rect -186 7602 -167 7622
rect -147 7602 -128 7622
rect -108 7602 0 7622
rect -251 7598 0 7602
rect 17068 7622 17313 7626
rect 17068 7602 17170 7622
rect 17190 7602 17209 7622
rect 17229 7602 17248 7622
rect 17268 7602 17287 7622
rect 17307 7602 17313 7622
rect 17068 7598 17313 7602
rect -949 7528 -943 7554
rect -768 7528 -762 7554
rect 17644 7528 17650 7554
rect 17825 7528 17831 7554
rect -440 7451 0 7455
rect -440 7431 -434 7451
rect -414 7431 -395 7451
rect -375 7431 -356 7451
rect -336 7431 -317 7451
rect -297 7431 0 7451
rect -440 7427 0 7431
rect 17068 7451 17503 7455
rect 17068 7431 17359 7451
rect 17379 7431 17398 7451
rect 17418 7431 17437 7451
rect 17457 7431 17476 7451
rect 17496 7431 17503 7451
rect 17068 7427 17503 7431
rect -659 7420 -625 7423
rect -659 7403 -651 7420
rect -634 7413 -625 7420
rect -634 7403 0 7413
rect -659 7399 0 7403
rect 20151 7371 20567 7377
rect 17355 7319 18077 7326
rect -673 7284 0 7298
rect 17355 7291 17370 7319
rect 17398 7291 17417 7319
rect 17445 7291 17464 7319
rect 17492 7312 18077 7319
rect 17492 7291 17898 7312
rect 17355 7280 17898 7291
rect 17930 7280 17942 7312
rect 17974 7280 17986 7312
rect 18018 7280 18030 7312
rect 18062 7280 18077 7312
rect 20151 7290 20442 7371
rect 20561 7290 20567 7371
rect 20151 7285 20567 7290
rect 17355 7272 18077 7280
rect -673 7243 0 7257
rect 17355 7244 17370 7272
rect 17398 7244 17417 7272
rect 17445 7244 17464 7272
rect 17492 7267 18077 7272
rect 17492 7244 17898 7267
rect 17355 7235 17898 7244
rect 17930 7235 17942 7267
rect 17974 7235 17986 7267
rect 18018 7235 18030 7267
rect 18062 7235 18077 7267
rect -605 7226 0 7229
rect -605 7209 -597 7226
rect -580 7215 0 7226
rect 17355 7225 18077 7235
rect -580 7209 -571 7215
rect -605 7205 -571 7209
rect 17355 7197 17370 7225
rect 17398 7197 17417 7225
rect 17445 7197 17464 7225
rect 17492 7222 18077 7225
rect 17492 7197 17898 7222
rect 17355 7190 17898 7197
rect 17930 7190 17942 7222
rect 17974 7190 17986 7222
rect 18018 7190 18030 7222
rect 18062 7190 18077 7222
rect 17355 7186 18077 7190
rect 20435 7168 20567 7181
rect -551 7155 -465 7158
rect -551 7135 -545 7155
rect -525 7135 -506 7155
rect -486 7152 -465 7155
rect 17527 7155 17613 7158
rect 17527 7152 17548 7155
rect -486 7138 0 7152
rect 17068 7138 17548 7152
rect -486 7135 -465 7138
rect -551 7132 -465 7135
rect 17527 7135 17548 7138
rect 17568 7135 17587 7155
rect 17607 7135 17613 7155
rect 17527 7132 17613 7135
rect -251 7120 0 7124
rect -949 7088 -943 7114
rect -768 7088 -762 7114
rect -251 7100 -245 7120
rect -225 7100 -206 7120
rect -186 7100 -167 7120
rect -147 7100 -128 7120
rect -108 7100 0 7120
rect -251 7096 0 7100
rect 17068 7120 17313 7124
rect 17068 7100 17170 7120
rect 17190 7100 17209 7120
rect 17229 7100 17248 7120
rect 17268 7100 17287 7120
rect 17307 7100 17313 7120
rect 17068 7096 17313 7100
rect 17644 7088 17650 7114
rect 17825 7088 17831 7114
rect 20435 6962 20448 7168
rect 20554 6962 20567 7168
rect -440 6949 0 6953
rect -440 6929 -434 6949
rect -414 6929 -395 6949
rect -375 6929 -356 6949
rect -336 6929 -317 6949
rect -297 6929 0 6949
rect -440 6925 0 6929
rect 17068 6949 17503 6953
rect 20435 6950 20567 6962
rect 17068 6929 17359 6949
rect 17379 6929 17398 6949
rect 17418 6929 17437 6949
rect 17457 6929 17476 6949
rect 17496 6929 17503 6949
rect 17068 6925 17503 6929
rect 20151 6937 20319 6946
rect -659 6918 -625 6921
rect -659 6901 -651 6918
rect -634 6911 -625 6918
rect -634 6901 0 6911
rect -659 6897 0 6901
rect 17167 6864 17838 6865
rect 17167 6857 17839 6864
rect 17167 6829 17181 6857
rect 17209 6829 17228 6857
rect 17256 6829 17275 6857
rect 17303 6851 17839 6857
rect 20151 6862 20202 6937
rect 20308 6862 20319 6937
rect 20151 6855 20319 6862
rect 17303 6829 17660 6851
rect 17167 6819 17660 6829
rect 17692 6819 17704 6851
rect 17736 6819 17748 6851
rect 17780 6819 17792 6851
rect 17824 6819 17839 6851
rect 17167 6810 17839 6819
rect -673 6782 0 6796
rect 17167 6782 17181 6810
rect 17209 6782 17228 6810
rect 17256 6782 17275 6810
rect 17303 6806 17839 6810
rect 17303 6782 17660 6806
rect 17167 6774 17660 6782
rect 17692 6774 17704 6806
rect 17736 6774 17748 6806
rect 17780 6774 17792 6806
rect 17824 6774 17839 6806
rect 17167 6763 17839 6774
rect -673 6741 0 6755
rect 17167 6735 17181 6763
rect 17209 6735 17228 6763
rect 17256 6735 17275 6763
rect 17303 6761 17839 6763
rect 17303 6735 17660 6761
rect 17167 6729 17660 6735
rect 17692 6729 17704 6761
rect 17736 6729 17748 6761
rect 17780 6729 17792 6761
rect 17824 6729 17839 6761
rect -605 6724 0 6727
rect 17167 6726 17839 6729
rect -605 6707 -597 6724
rect -580 6713 0 6724
rect -580 6707 -571 6713
rect -605 6703 -571 6707
rect -949 6648 -943 6674
rect -768 6648 -762 6674
rect -551 6653 -465 6656
rect -551 6633 -545 6653
rect -525 6633 -506 6653
rect -486 6650 -465 6653
rect 17527 6653 17613 6656
rect 17527 6650 17548 6653
rect -486 6636 0 6650
rect 17068 6636 17548 6650
rect -486 6633 -465 6636
rect -551 6630 -465 6633
rect 17527 6633 17548 6636
rect 17568 6633 17587 6653
rect 17607 6633 17613 6653
rect 17644 6648 17650 6674
rect 17825 6648 17831 6674
rect 20151 6666 20319 6675
rect 17527 6630 17613 6633
rect -251 6618 0 6622
rect -251 6598 -245 6618
rect -225 6598 -206 6618
rect -186 6598 -167 6618
rect -147 6598 -128 6618
rect -108 6598 0 6618
rect -251 6594 0 6598
rect 17068 6618 17313 6622
rect 17068 6598 17170 6618
rect 17190 6598 17209 6618
rect 17229 6598 17248 6618
rect 17268 6598 17287 6618
rect 17307 6598 17313 6618
rect 17068 6594 17313 6598
rect 20151 6591 20202 6666
rect 20308 6591 20319 6666
rect 20151 6584 20319 6591
rect -440 6447 0 6451
rect -440 6427 -434 6447
rect -414 6427 -395 6447
rect -375 6427 -356 6447
rect -336 6427 -317 6447
rect -297 6427 0 6447
rect -440 6423 0 6427
rect 17068 6447 17503 6451
rect 17068 6427 17359 6447
rect 17379 6427 17398 6447
rect 17418 6427 17437 6447
rect 17457 6427 17476 6447
rect 17496 6427 17503 6447
rect 17068 6423 17503 6427
rect -659 6416 -625 6419
rect -659 6399 -651 6416
rect -634 6409 -625 6416
rect -634 6399 0 6409
rect -659 6395 0 6399
rect 20151 6388 20319 6397
rect 17354 6354 18076 6361
rect 17354 6326 17369 6354
rect 17397 6326 17416 6354
rect 17444 6326 17463 6354
rect 17491 6347 18076 6354
rect 17491 6326 17897 6347
rect 17354 6315 17897 6326
rect 17929 6315 17941 6347
rect 17973 6315 17985 6347
rect 18017 6315 18029 6347
rect 18061 6315 18076 6347
rect 17354 6307 18076 6315
rect -673 6280 0 6294
rect 17354 6279 17369 6307
rect 17397 6279 17416 6307
rect 17444 6279 17463 6307
rect 17491 6302 18076 6307
rect 20151 6313 20202 6388
rect 20308 6313 20319 6388
rect 20151 6306 20319 6313
rect 17491 6279 17897 6302
rect 17354 6270 17897 6279
rect 17929 6270 17941 6302
rect 17973 6270 17985 6302
rect 18017 6270 18029 6302
rect 18061 6270 18076 6302
rect 17354 6260 18076 6270
rect -673 6239 0 6253
rect -949 6208 -943 6234
rect -768 6208 -762 6234
rect 17354 6232 17369 6260
rect 17397 6232 17416 6260
rect 17444 6232 17463 6260
rect 17491 6257 18076 6260
rect 17491 6232 17897 6257
rect 17354 6225 17897 6232
rect 17929 6225 17941 6257
rect 17973 6225 17985 6257
rect 18017 6225 18029 6257
rect 18061 6225 18076 6257
rect -605 6222 0 6225
rect -605 6205 -597 6222
rect -580 6211 0 6222
rect 17354 6221 18076 6225
rect 20435 6289 20567 6302
rect -580 6205 -571 6211
rect -605 6201 -571 6205
rect -551 6151 -465 6154
rect -551 6131 -545 6151
rect -525 6131 -506 6151
rect -486 6148 -465 6151
rect 17527 6151 17613 6154
rect 17527 6148 17548 6151
rect -486 6134 0 6148
rect 17068 6134 17548 6148
rect -486 6131 -465 6134
rect -551 6128 -465 6131
rect 17527 6131 17548 6134
rect 17568 6131 17587 6151
rect 17607 6131 17613 6151
rect 17527 6128 17613 6131
rect -251 6116 0 6120
rect -251 6096 -245 6116
rect -225 6096 -206 6116
rect -186 6096 -167 6116
rect -147 6096 -128 6116
rect -108 6096 0 6116
rect -251 6092 0 6096
rect 17068 6116 17313 6120
rect 17068 6096 17170 6116
rect 17190 6096 17209 6116
rect 17229 6096 17248 6116
rect 17268 6096 17287 6116
rect 17307 6096 17313 6116
rect 17068 6092 17313 6096
rect 20435 6083 20448 6289
rect 20554 6083 20567 6289
rect 20435 6071 20567 6083
rect -440 5945 0 5949
rect -440 5925 -434 5945
rect -414 5925 -395 5945
rect -375 5925 -356 5945
rect -336 5925 -317 5945
rect -297 5925 0 5945
rect -440 5921 0 5925
rect 17068 5945 17503 5949
rect 17068 5925 17359 5945
rect 17379 5925 17398 5945
rect 17418 5925 17437 5945
rect 17457 5925 17476 5945
rect 17496 5925 17503 5945
rect 17068 5921 17503 5925
rect -659 5914 -625 5917
rect -659 5897 -651 5914
rect -634 5907 -625 5914
rect -634 5897 0 5907
rect -659 5893 0 5897
rect 17168 5902 17839 5903
rect 17168 5895 17840 5902
rect 17168 5867 17182 5895
rect 17210 5867 17229 5895
rect 17257 5867 17276 5895
rect 17304 5889 17840 5895
rect 17304 5867 17661 5889
rect 17168 5857 17661 5867
rect 17693 5857 17705 5889
rect 17737 5857 17749 5889
rect 17781 5857 17793 5889
rect 17825 5857 17840 5889
rect 17168 5848 17840 5857
rect 17168 5820 17182 5848
rect 17210 5820 17229 5848
rect 17257 5820 17276 5848
rect 17304 5844 17840 5848
rect 17304 5820 17661 5844
rect 17168 5812 17661 5820
rect 17693 5812 17705 5844
rect 17737 5812 17749 5844
rect 17781 5812 17793 5844
rect 17825 5812 17840 5844
rect 17168 5801 17840 5812
rect -949 5768 -943 5794
rect -768 5768 -762 5794
rect -673 5778 0 5792
rect 17168 5773 17182 5801
rect 17210 5773 17229 5801
rect 17257 5773 17276 5801
rect 17304 5799 17840 5801
rect 17304 5794 17661 5799
rect 17693 5794 17705 5799
rect 17737 5794 17749 5799
rect 17781 5794 17793 5799
rect 17304 5773 17650 5794
rect 17168 5768 17650 5773
rect 17168 5767 17661 5768
rect 17693 5767 17705 5768
rect 17737 5767 17749 5768
rect 17781 5767 17793 5768
rect 17825 5767 17840 5799
rect 17168 5763 17840 5767
rect 20151 5816 20567 5822
rect -673 5737 0 5751
rect 20151 5735 20442 5816
rect 20561 5735 20567 5816
rect 20151 5730 20567 5735
rect -605 5720 0 5723
rect -605 5703 -597 5720
rect -580 5709 0 5720
rect -580 5703 -571 5709
rect -605 5699 -571 5703
rect -551 5649 -465 5652
rect -551 5629 -545 5649
rect -525 5629 -506 5649
rect -486 5646 -465 5649
rect 17527 5649 17613 5652
rect 17527 5646 17548 5649
rect -486 5632 0 5646
rect 17068 5632 17548 5646
rect -486 5629 -465 5632
rect -551 5626 -465 5629
rect 17527 5629 17548 5632
rect 17568 5629 17587 5649
rect 17607 5629 17613 5649
rect 17527 5626 17613 5629
rect -251 5614 0 5618
rect -251 5594 -245 5614
rect -225 5594 -206 5614
rect -186 5594 -167 5614
rect -147 5594 -128 5614
rect -108 5594 0 5614
rect -251 5590 0 5594
rect 17068 5614 17313 5618
rect 17068 5594 17170 5614
rect 17190 5594 17209 5614
rect 17229 5594 17248 5614
rect 17268 5594 17287 5614
rect 17307 5594 17313 5614
rect 17068 5590 17313 5594
rect -440 5443 0 5447
rect -440 5423 -434 5443
rect -414 5423 -395 5443
rect -375 5423 -356 5443
rect -336 5423 -317 5443
rect -297 5423 0 5443
rect -440 5419 0 5423
rect 17068 5443 17503 5447
rect 17068 5423 17359 5443
rect 17379 5423 17398 5443
rect 17418 5423 17437 5443
rect 17457 5423 17476 5443
rect 17496 5423 17503 5443
rect 17068 5419 17503 5423
rect -659 5412 -625 5415
rect -659 5395 -651 5412
rect -634 5405 -625 5412
rect -634 5395 0 5405
rect -659 5391 0 5395
rect 20151 5371 20567 5377
rect -949 5328 -943 5354
rect -768 5328 -762 5354
rect 17355 5346 18077 5353
rect 17355 5318 17370 5346
rect 17398 5318 17417 5346
rect 17445 5318 17464 5346
rect 17492 5339 18077 5346
rect 17492 5318 17898 5339
rect 17355 5307 17898 5318
rect 17930 5307 17942 5339
rect 17974 5307 17986 5339
rect 18018 5307 18030 5339
rect 18062 5307 18077 5339
rect 17355 5299 18077 5307
rect -673 5276 0 5290
rect 17355 5271 17370 5299
rect 17398 5271 17417 5299
rect 17445 5271 17464 5299
rect 17492 5294 18077 5299
rect 17492 5271 17898 5294
rect 17355 5262 17898 5271
rect 17930 5262 17942 5294
rect 17974 5262 17986 5294
rect 18018 5262 18030 5294
rect 18062 5262 18077 5294
rect 20151 5290 20442 5371
rect 20561 5290 20567 5371
rect 20151 5285 20567 5290
rect 17355 5252 18077 5262
rect -673 5235 0 5249
rect 17355 5224 17370 5252
rect 17398 5224 17417 5252
rect 17445 5224 17464 5252
rect 17492 5249 18077 5252
rect 17492 5224 17898 5249
rect -605 5218 0 5221
rect -605 5201 -597 5218
rect -580 5207 0 5218
rect 17355 5217 17898 5224
rect 17930 5217 17942 5249
rect 17974 5217 17986 5249
rect 18018 5217 18030 5249
rect 18062 5217 18077 5249
rect 17355 5213 18077 5217
rect -580 5201 -571 5207
rect -605 5197 -571 5201
rect 20435 5168 20567 5181
rect -551 5147 -465 5150
rect -551 5127 -545 5147
rect -525 5127 -506 5147
rect -486 5144 -465 5147
rect 17527 5147 17613 5150
rect 17527 5144 17548 5147
rect -486 5130 0 5144
rect 17068 5130 17548 5144
rect -486 5127 -465 5130
rect -551 5124 -465 5127
rect 17527 5127 17548 5130
rect 17568 5127 17587 5147
rect 17607 5127 17613 5147
rect 17527 5124 17613 5127
rect -251 5112 0 5116
rect -251 5092 -245 5112
rect -225 5092 -206 5112
rect -186 5092 -167 5112
rect -147 5092 -128 5112
rect -108 5092 0 5112
rect -251 5088 0 5092
rect 17068 5112 17313 5116
rect 17068 5092 17170 5112
rect 17190 5092 17209 5112
rect 17229 5092 17248 5112
rect 17268 5092 17287 5112
rect 17307 5092 17313 5112
rect 17068 5088 17313 5092
rect 20435 4962 20448 5168
rect 20554 4962 20567 5168
rect 20435 4950 20567 4962
rect -440 4941 0 4945
rect -440 4921 -434 4941
rect -414 4921 -395 4941
rect -375 4921 -356 4941
rect -336 4921 -317 4941
rect -297 4921 0 4941
rect -440 4917 0 4921
rect 17068 4941 17503 4945
rect 17068 4921 17359 4941
rect 17379 4921 17398 4941
rect 17418 4921 17437 4941
rect 17457 4921 17476 4941
rect 17496 4921 17503 4941
rect 17068 4917 17503 4921
rect 20151 4937 20319 4946
rect -949 4888 -943 4914
rect -768 4888 -762 4914
rect -659 4910 -625 4913
rect -659 4893 -651 4910
rect -634 4903 -625 4910
rect -634 4893 0 4903
rect -659 4889 0 4893
rect 17644 4888 17650 4914
rect 17825 4888 17831 4914
rect 20151 4862 20202 4937
rect 20308 4862 20319 4937
rect 20151 4855 20319 4862
rect 17167 4839 17838 4840
rect 17167 4832 17839 4839
rect 17167 4804 17181 4832
rect 17209 4804 17228 4832
rect 17256 4804 17275 4832
rect 17303 4826 17839 4832
rect 17303 4804 17660 4826
rect 17167 4794 17660 4804
rect 17692 4794 17704 4826
rect 17736 4794 17748 4826
rect 17780 4794 17792 4826
rect 17824 4794 17839 4826
rect -673 4774 0 4788
rect 17167 4785 17839 4794
rect 17167 4757 17181 4785
rect 17209 4757 17228 4785
rect 17256 4757 17275 4785
rect 17303 4781 17839 4785
rect 17303 4757 17660 4781
rect 17167 4749 17660 4757
rect 17692 4749 17704 4781
rect 17736 4749 17748 4781
rect 17780 4749 17792 4781
rect 17824 4749 17839 4781
rect -673 4733 0 4747
rect 17167 4738 17839 4749
rect -605 4716 0 4719
rect -605 4699 -597 4716
rect -580 4705 0 4716
rect 17167 4710 17181 4738
rect 17209 4710 17228 4738
rect 17256 4710 17275 4738
rect 17303 4736 17839 4738
rect 17303 4710 17660 4736
rect -580 4699 -571 4705
rect 17167 4704 17660 4710
rect 17692 4704 17704 4736
rect 17736 4704 17748 4736
rect 17780 4704 17792 4736
rect 17824 4704 17839 4736
rect 17167 4700 17839 4704
rect -605 4695 -571 4699
rect 20151 4666 20319 4675
rect -551 4645 -465 4648
rect -551 4625 -545 4645
rect -525 4625 -506 4645
rect -486 4642 -465 4645
rect 17527 4645 17613 4648
rect 17527 4642 17548 4645
rect -486 4628 0 4642
rect 17068 4628 17548 4642
rect -486 4625 -465 4628
rect -551 4622 -465 4625
rect 17527 4625 17548 4628
rect 17568 4625 17587 4645
rect 17607 4625 17613 4645
rect 17527 4622 17613 4625
rect -251 4610 0 4614
rect -251 4590 -245 4610
rect -225 4590 -206 4610
rect -186 4590 -167 4610
rect -147 4590 -128 4610
rect -108 4590 0 4610
rect -251 4586 0 4590
rect 17068 4610 17313 4614
rect 17068 4590 17170 4610
rect 17190 4590 17209 4610
rect 17229 4590 17248 4610
rect 17268 4590 17287 4610
rect 17307 4590 17313 4610
rect 17068 4586 17313 4590
rect 20151 4591 20202 4666
rect 20308 4591 20319 4666
rect 20151 4584 20319 4591
rect -949 4448 -943 4474
rect -768 4448 -762 4474
rect 17644 4448 17650 4474
rect 17825 4448 17831 4474
rect -440 4439 0 4443
rect -440 4419 -434 4439
rect -414 4419 -395 4439
rect -375 4419 -356 4439
rect -336 4419 -317 4439
rect -297 4419 0 4439
rect -440 4415 0 4419
rect 17068 4439 17503 4443
rect 17068 4419 17359 4439
rect 17379 4419 17398 4439
rect 17418 4419 17437 4439
rect 17457 4419 17476 4439
rect 17496 4419 17503 4439
rect 17068 4415 17503 4419
rect -659 4408 -625 4411
rect -659 4391 -651 4408
rect -634 4401 -625 4408
rect -634 4391 0 4401
rect -659 4387 0 4391
rect 20151 4388 20319 4397
rect 17355 4345 18077 4352
rect 17355 4317 17370 4345
rect 17398 4317 17417 4345
rect 17445 4317 17464 4345
rect 17492 4338 18077 4345
rect 17492 4317 17898 4338
rect 17355 4306 17898 4317
rect 17930 4306 17942 4338
rect 17974 4306 17986 4338
rect 18018 4306 18030 4338
rect 18062 4306 18077 4338
rect 20151 4313 20202 4388
rect 20308 4313 20319 4388
rect 20151 4306 20319 4313
rect 17355 4298 18077 4306
rect -673 4272 0 4286
rect 17355 4270 17370 4298
rect 17398 4270 17417 4298
rect 17445 4270 17464 4298
rect 17492 4293 18077 4298
rect 17492 4270 17898 4293
rect 17355 4261 17898 4270
rect 17930 4261 17942 4293
rect 17974 4261 17986 4293
rect 18018 4261 18030 4293
rect 18062 4261 18077 4293
rect 17355 4251 18077 4261
rect -673 4231 0 4245
rect 17355 4223 17370 4251
rect 17398 4223 17417 4251
rect 17445 4223 17464 4251
rect 17492 4248 18077 4251
rect 17492 4223 17898 4248
rect -605 4214 0 4217
rect -605 4197 -597 4214
rect -580 4203 0 4214
rect 17355 4216 17898 4223
rect 17930 4216 17942 4248
rect 17974 4216 17986 4248
rect 18018 4216 18030 4248
rect 18062 4216 18077 4248
rect 17355 4212 18077 4216
rect 20435 4289 20567 4302
rect -580 4197 -571 4203
rect -605 4193 -571 4197
rect -551 4143 -465 4146
rect -551 4123 -545 4143
rect -525 4123 -506 4143
rect -486 4140 -465 4143
rect 17527 4143 17613 4146
rect 17527 4140 17548 4143
rect -486 4126 0 4140
rect 17068 4126 17548 4140
rect -486 4123 -465 4126
rect -551 4120 -465 4123
rect 17527 4123 17548 4126
rect 17568 4123 17587 4143
rect 17607 4123 17613 4143
rect 17527 4120 17613 4123
rect -251 4108 0 4112
rect -251 4088 -245 4108
rect -225 4088 -206 4108
rect -186 4088 -167 4108
rect -147 4088 -128 4108
rect -108 4088 0 4108
rect -251 4084 0 4088
rect 17068 4108 17313 4112
rect 17068 4088 17170 4108
rect 17190 4088 17209 4108
rect 17229 4088 17248 4108
rect 17268 4088 17287 4108
rect 17307 4088 17313 4108
rect 17068 4084 17313 4088
rect 20435 4083 20448 4289
rect 20554 4083 20567 4289
rect 20435 4071 20567 4083
rect -949 4008 -943 4034
rect -768 4008 -762 4034
rect 17644 4008 17650 4034
rect 17825 4008 17831 4034
rect -440 3937 0 3941
rect -440 3917 -434 3937
rect -414 3917 -395 3937
rect -375 3917 -356 3937
rect -336 3917 -317 3937
rect -297 3917 0 3937
rect -440 3913 0 3917
rect 17068 3937 17503 3941
rect 17068 3917 17359 3937
rect 17379 3917 17398 3937
rect 17418 3917 17437 3937
rect 17457 3917 17476 3937
rect 17496 3917 17503 3937
rect 17068 3913 17503 3917
rect -659 3906 -625 3909
rect -659 3889 -651 3906
rect -634 3899 -625 3906
rect -634 3889 0 3899
rect -659 3885 0 3889
rect 17168 3851 17839 3852
rect 17168 3844 17840 3851
rect 17168 3816 17182 3844
rect 17210 3816 17229 3844
rect 17257 3816 17276 3844
rect 17304 3838 17840 3844
rect 17304 3816 17661 3838
rect 17168 3806 17661 3816
rect 17693 3806 17705 3838
rect 17737 3806 17749 3838
rect 17781 3806 17793 3838
rect 17825 3806 17840 3838
rect 17168 3797 17840 3806
rect -673 3770 0 3784
rect 17168 3769 17182 3797
rect 17210 3769 17229 3797
rect 17257 3769 17276 3797
rect 17304 3793 17840 3797
rect 17304 3769 17661 3793
rect 17168 3761 17661 3769
rect 17693 3761 17705 3793
rect 17737 3761 17749 3793
rect 17781 3761 17793 3793
rect 17825 3761 17840 3793
rect 17168 3750 17840 3761
rect -673 3729 0 3743
rect 17168 3722 17182 3750
rect 17210 3722 17229 3750
rect 17257 3722 17276 3750
rect 17304 3748 17840 3750
rect 17304 3722 17661 3748
rect 17168 3716 17661 3722
rect 17693 3716 17705 3748
rect 17737 3716 17749 3748
rect 17781 3716 17793 3748
rect 17825 3716 17840 3748
rect 20151 3816 20567 3822
rect 20151 3735 20442 3816
rect 20561 3735 20567 3816
rect 20151 3730 20567 3735
rect -605 3712 0 3715
rect 17168 3712 17840 3716
rect -605 3695 -597 3712
rect -580 3701 0 3712
rect -580 3695 -571 3701
rect -605 3691 -571 3695
rect -551 3641 -465 3644
rect -551 3621 -545 3641
rect -525 3621 -506 3641
rect -486 3638 -465 3641
rect 17527 3641 17613 3644
rect 17527 3638 17548 3641
rect -486 3624 0 3638
rect 17068 3624 17548 3638
rect -486 3621 -465 3624
rect -551 3618 -465 3621
rect 17527 3621 17548 3624
rect 17568 3621 17587 3641
rect 17607 3621 17613 3641
rect 17527 3618 17613 3621
rect -251 3606 0 3610
rect -949 3568 -943 3594
rect -768 3568 -762 3594
rect -251 3586 -245 3606
rect -225 3586 -206 3606
rect -186 3586 -167 3606
rect -147 3586 -128 3606
rect -108 3586 0 3606
rect -251 3582 0 3586
rect 17068 3606 17313 3610
rect 17068 3586 17170 3606
rect 17190 3586 17209 3606
rect 17229 3586 17248 3606
rect 17268 3586 17287 3606
rect 17307 3586 17313 3606
rect 17068 3582 17313 3586
rect 17644 3568 17650 3594
rect 17825 3568 17831 3594
rect -440 3435 0 3439
rect -440 3415 -434 3435
rect -414 3415 -395 3435
rect -375 3415 -356 3435
rect -336 3415 -317 3435
rect -297 3415 0 3435
rect -440 3411 0 3415
rect 17068 3435 17503 3439
rect 17068 3415 17359 3435
rect 17379 3415 17398 3435
rect 17418 3415 17437 3435
rect 17457 3415 17476 3435
rect 17496 3415 17503 3435
rect 17068 3411 17503 3415
rect -659 3404 -625 3407
rect -659 3387 -651 3404
rect -634 3397 -625 3404
rect -634 3387 0 3397
rect -659 3383 0 3387
rect 20151 3371 20567 3377
rect 17354 3346 18076 3353
rect 17354 3318 17369 3346
rect 17397 3318 17416 3346
rect 17444 3318 17463 3346
rect 17491 3339 18076 3346
rect 17491 3318 17897 3339
rect 17354 3307 17897 3318
rect 17929 3307 17941 3339
rect 17973 3307 17985 3339
rect 18017 3307 18029 3339
rect 18061 3307 18076 3339
rect 17354 3299 18076 3307
rect -673 3268 0 3282
rect 17354 3271 17369 3299
rect 17397 3271 17416 3299
rect 17444 3271 17463 3299
rect 17491 3294 18076 3299
rect 17491 3271 17897 3294
rect 17354 3262 17897 3271
rect 17929 3262 17941 3294
rect 17973 3262 17985 3294
rect 18017 3262 18029 3294
rect 18061 3262 18076 3294
rect 20151 3290 20442 3371
rect 20561 3290 20567 3371
rect 20151 3285 20567 3290
rect 17354 3252 18076 3262
rect -673 3227 0 3241
rect 17354 3224 17369 3252
rect 17397 3224 17416 3252
rect 17444 3224 17463 3252
rect 17491 3249 18076 3252
rect 17491 3224 17897 3249
rect 17354 3217 17897 3224
rect 17929 3217 17941 3249
rect 17973 3217 17985 3249
rect 18017 3217 18029 3249
rect 18061 3217 18076 3249
rect 17354 3213 18076 3217
rect -605 3210 0 3213
rect -605 3193 -597 3210
rect -580 3199 0 3210
rect -580 3193 -571 3199
rect -605 3189 -571 3193
rect 20435 3168 20567 3181
rect -949 3128 -943 3154
rect -768 3128 -762 3154
rect -551 3139 -465 3142
rect -551 3119 -545 3139
rect -525 3119 -506 3139
rect -486 3136 -465 3139
rect 17527 3139 17613 3142
rect 17527 3136 17548 3139
rect -486 3122 0 3136
rect 17068 3122 17548 3136
rect -486 3119 -465 3122
rect -551 3116 -465 3119
rect 17527 3119 17548 3122
rect 17568 3119 17587 3139
rect 17607 3119 17613 3139
rect 17644 3128 17650 3154
rect 17825 3128 17831 3154
rect 17527 3116 17613 3119
rect -251 3104 0 3108
rect -251 3084 -245 3104
rect -225 3084 -206 3104
rect -186 3084 -167 3104
rect -147 3084 -128 3104
rect -108 3084 0 3104
rect -251 3080 0 3084
rect 17068 3104 17313 3108
rect 17068 3084 17170 3104
rect 17190 3084 17209 3104
rect 17229 3084 17248 3104
rect 17268 3084 17287 3104
rect 17307 3084 17313 3104
rect 17068 3080 17313 3084
rect 20435 2962 20448 3168
rect 20554 2962 20567 3168
rect 20435 2950 20567 2962
rect 20151 2937 20319 2946
rect -440 2933 0 2937
rect -440 2913 -434 2933
rect -414 2913 -395 2933
rect -375 2913 -356 2933
rect -336 2913 -317 2933
rect -297 2913 0 2933
rect -440 2909 0 2913
rect 17068 2933 17503 2937
rect 17068 2913 17359 2933
rect 17379 2913 17398 2933
rect 17418 2913 17437 2933
rect 17457 2913 17476 2933
rect 17496 2913 17503 2933
rect 17068 2909 17503 2913
rect -659 2902 -625 2905
rect -659 2885 -651 2902
rect -634 2895 -625 2902
rect -634 2885 0 2895
rect -659 2881 0 2885
rect 20151 2862 20202 2937
rect 20308 2862 20319 2937
rect 20151 2855 20319 2862
rect 17168 2829 17839 2830
rect 17168 2822 17840 2829
rect 17168 2794 17182 2822
rect 17210 2794 17229 2822
rect 17257 2794 17276 2822
rect 17304 2816 17840 2822
rect 17304 2794 17661 2816
rect 17168 2784 17661 2794
rect 17693 2784 17705 2816
rect 17737 2784 17749 2816
rect 17781 2784 17793 2816
rect 17825 2784 17840 2816
rect -673 2766 0 2780
rect 17168 2775 17840 2784
rect 17168 2747 17182 2775
rect 17210 2747 17229 2775
rect 17257 2747 17276 2775
rect 17304 2771 17840 2775
rect 17304 2747 17661 2771
rect 17168 2739 17661 2747
rect 17693 2739 17705 2771
rect 17737 2739 17749 2771
rect 17781 2739 17793 2771
rect 17825 2739 17840 2771
rect -673 2725 0 2739
rect 17168 2728 17840 2739
rect -949 2688 -943 2714
rect -768 2688 -762 2714
rect -605 2708 0 2711
rect -605 2691 -597 2708
rect -580 2697 0 2708
rect 17168 2700 17182 2728
rect 17210 2700 17229 2728
rect 17257 2700 17276 2728
rect 17304 2726 17840 2728
rect 17304 2714 17661 2726
rect 17693 2714 17705 2726
rect 17737 2714 17749 2726
rect 17781 2714 17793 2726
rect 17304 2700 17650 2714
rect -580 2691 -571 2697
rect -605 2687 -571 2691
rect 17168 2690 17650 2700
rect 17644 2688 17650 2690
rect 17825 2690 17840 2726
rect 17825 2688 17831 2690
rect 20151 2666 20319 2675
rect -551 2637 -465 2640
rect -551 2617 -545 2637
rect -525 2617 -506 2637
rect -486 2634 -465 2637
rect 17527 2637 17613 2640
rect 17527 2634 17548 2637
rect -486 2620 0 2634
rect 17068 2620 17548 2634
rect -486 2617 -465 2620
rect -551 2614 -465 2617
rect 17527 2617 17548 2620
rect 17568 2617 17587 2637
rect 17607 2617 17613 2637
rect 17527 2614 17613 2617
rect -251 2602 0 2606
rect -251 2582 -245 2602
rect -225 2582 -206 2602
rect -186 2582 -167 2602
rect -147 2582 -128 2602
rect -108 2582 0 2602
rect -251 2578 0 2582
rect 17068 2602 17313 2606
rect 17068 2582 17170 2602
rect 17190 2582 17209 2602
rect 17229 2582 17248 2602
rect 17268 2582 17287 2602
rect 17307 2582 17313 2602
rect 20151 2591 20202 2666
rect 20308 2591 20319 2666
rect 20151 2584 20319 2591
rect 17068 2578 17313 2582
rect -440 2431 0 2435
rect -440 2411 -434 2431
rect -414 2411 -395 2431
rect -375 2411 -356 2431
rect -336 2411 -317 2431
rect -297 2411 0 2431
rect -440 2407 0 2411
rect 17068 2431 17503 2435
rect 17068 2411 17359 2431
rect 17379 2411 17398 2431
rect 17418 2411 17437 2431
rect 17457 2411 17476 2431
rect 17496 2411 17503 2431
rect 17068 2407 17503 2411
rect -659 2400 -625 2403
rect -659 2383 -651 2400
rect -634 2393 -625 2400
rect -634 2383 0 2393
rect -659 2379 0 2383
rect 20151 2388 20319 2397
rect 17355 2312 18077 2319
rect 17355 2284 17370 2312
rect 17398 2284 17417 2312
rect 17445 2284 17464 2312
rect 17492 2305 18077 2312
rect 20151 2313 20202 2388
rect 20308 2313 20319 2388
rect 20151 2306 20319 2313
rect 17492 2284 17898 2305
rect -949 2248 -943 2274
rect -768 2248 -762 2274
rect -673 2264 0 2278
rect 17355 2273 17898 2284
rect 17930 2273 17942 2305
rect 17974 2273 17986 2305
rect 18018 2273 18030 2305
rect 18062 2273 18077 2305
rect 17355 2265 18077 2273
rect 17355 2237 17370 2265
rect 17398 2237 17417 2265
rect 17445 2237 17464 2265
rect 17492 2260 18077 2265
rect 17492 2237 17898 2260
rect -673 2223 0 2237
rect 17355 2228 17898 2237
rect 17930 2228 17942 2260
rect 17974 2228 17986 2260
rect 18018 2228 18030 2260
rect 18062 2228 18077 2260
rect 17355 2218 18077 2228
rect -605 2206 0 2209
rect -605 2189 -597 2206
rect -580 2195 0 2206
rect -580 2189 -571 2195
rect -605 2185 -571 2189
rect 17355 2190 17370 2218
rect 17398 2190 17417 2218
rect 17445 2190 17464 2218
rect 17492 2215 18077 2218
rect 17492 2190 17898 2215
rect 17355 2183 17898 2190
rect 17930 2183 17942 2215
rect 17974 2183 17986 2215
rect 18018 2183 18030 2215
rect 18062 2183 18077 2215
rect 17355 2179 18077 2183
rect 20435 2289 20567 2302
rect -551 2135 -465 2138
rect -551 2115 -545 2135
rect -525 2115 -506 2135
rect -486 2132 -465 2135
rect 17527 2135 17613 2138
rect 17527 2132 17548 2135
rect -486 2118 0 2132
rect 17068 2118 17548 2132
rect -486 2115 -465 2118
rect -551 2112 -465 2115
rect 17527 2115 17548 2118
rect 17568 2115 17587 2135
rect 17607 2115 17613 2135
rect 17527 2112 17613 2115
rect -251 2100 0 2104
rect -251 2080 -245 2100
rect -225 2080 -206 2100
rect -186 2080 -167 2100
rect -147 2080 -128 2100
rect -108 2080 0 2100
rect -251 2076 0 2080
rect 17068 2100 17313 2104
rect 17068 2080 17170 2100
rect 17190 2080 17209 2100
rect 17229 2080 17248 2100
rect 17268 2080 17287 2100
rect 17307 2080 17313 2100
rect 17068 2076 17313 2080
rect 20435 2083 20448 2289
rect 20554 2083 20567 2289
rect 20435 2071 20567 2083
rect -440 1929 0 1933
rect -440 1909 -434 1929
rect -414 1909 -395 1929
rect -375 1909 -356 1929
rect -336 1909 -317 1929
rect -297 1909 0 1929
rect -440 1905 0 1909
rect 17068 1929 17503 1933
rect 17068 1909 17359 1929
rect 17379 1909 17398 1929
rect 17418 1909 17437 1929
rect 17457 1909 17476 1929
rect 17496 1909 17503 1929
rect 17068 1905 17503 1909
rect -659 1898 -625 1901
rect -659 1881 -651 1898
rect -634 1891 -625 1898
rect -634 1881 0 1891
rect -659 1877 0 1881
rect -949 1808 -943 1834
rect -768 1808 -762 1834
rect 17644 1833 17650 1834
rect 17167 1825 17650 1833
rect 17825 1833 17831 1834
rect 17167 1797 17182 1825
rect 17210 1797 17229 1825
rect 17257 1797 17276 1825
rect 17304 1808 17650 1825
rect 17304 1797 17661 1808
rect 17167 1787 17661 1797
rect 17693 1787 17705 1808
rect 17737 1787 17749 1808
rect 17781 1787 17793 1808
rect 17825 1787 17839 1833
rect 17167 1778 17839 1787
rect -673 1762 0 1776
rect 17167 1750 17182 1778
rect 17210 1750 17229 1778
rect 17257 1750 17276 1778
rect 17304 1774 17839 1778
rect 17304 1750 17661 1774
rect 17167 1742 17661 1750
rect 17693 1742 17705 1774
rect 17737 1742 17749 1774
rect 17781 1742 17793 1774
rect 17825 1742 17839 1774
rect -673 1721 0 1735
rect 17167 1731 17839 1742
rect -605 1704 0 1707
rect -605 1687 -597 1704
rect -580 1693 0 1704
rect 17167 1703 17182 1731
rect 17210 1703 17229 1731
rect 17257 1703 17276 1731
rect 17304 1729 17839 1731
rect 20151 1816 20567 1822
rect 20151 1735 20442 1816
rect 20561 1735 20567 1816
rect 20151 1730 20567 1735
rect 17304 1703 17661 1729
rect 17167 1697 17661 1703
rect 17693 1697 17705 1729
rect 17737 1697 17749 1729
rect 17781 1697 17793 1729
rect 17825 1697 17839 1729
rect 17167 1693 17839 1697
rect -580 1687 -571 1693
rect -605 1683 -571 1687
rect -551 1633 -465 1636
rect -551 1613 -545 1633
rect -525 1613 -506 1633
rect -486 1630 -465 1633
rect 17527 1633 17613 1636
rect 17527 1630 17548 1633
rect -486 1616 0 1630
rect 17068 1616 17548 1630
rect -486 1613 -465 1616
rect -551 1610 -465 1613
rect 17527 1613 17548 1616
rect 17568 1613 17587 1633
rect 17607 1613 17613 1633
rect 17527 1610 17613 1613
rect -251 1598 0 1602
rect -251 1578 -245 1598
rect -225 1578 -206 1598
rect -186 1578 -167 1598
rect -147 1578 -128 1598
rect -108 1578 0 1598
rect -251 1574 0 1578
rect 17068 1598 17313 1602
rect 17068 1578 17170 1598
rect 17190 1578 17209 1598
rect 17229 1578 17248 1598
rect 17268 1578 17287 1598
rect 17307 1578 17313 1598
rect 17068 1574 17313 1578
rect -440 1427 0 1431
rect -440 1407 -434 1427
rect -414 1407 -395 1427
rect -375 1407 -356 1427
rect -336 1407 -317 1427
rect -297 1407 0 1427
rect -440 1403 0 1407
rect 17068 1427 17503 1431
rect 17068 1407 17359 1427
rect 17379 1407 17398 1427
rect 17418 1407 17437 1427
rect 17457 1407 17476 1427
rect 17496 1407 17503 1427
rect 17068 1403 17503 1407
rect -659 1396 -625 1399
rect -949 1368 -943 1394
rect -768 1368 -762 1394
rect -659 1379 -651 1396
rect -634 1389 -625 1396
rect -634 1379 0 1389
rect -659 1375 0 1379
rect 17644 1368 17650 1394
rect 17825 1368 17831 1394
rect 20151 1371 20567 1377
rect 17355 1310 18077 1317
rect 17355 1282 17370 1310
rect 17398 1282 17417 1310
rect 17445 1282 17464 1310
rect 17492 1303 18077 1310
rect 17492 1282 17898 1303
rect -673 1260 0 1274
rect 17355 1271 17898 1282
rect 17930 1271 17942 1303
rect 17974 1271 17986 1303
rect 18018 1271 18030 1303
rect 18062 1271 18077 1303
rect 20151 1290 20442 1371
rect 20561 1290 20567 1371
rect 20151 1285 20567 1290
rect 17355 1263 18077 1271
rect 17355 1235 17370 1263
rect 17398 1235 17417 1263
rect 17445 1235 17464 1263
rect 17492 1258 18077 1263
rect 17492 1235 17898 1258
rect -673 1219 0 1233
rect 17355 1226 17898 1235
rect 17930 1226 17942 1258
rect 17974 1226 17986 1258
rect 18018 1226 18030 1258
rect 18062 1226 18077 1258
rect 17355 1216 18077 1226
rect -605 1202 0 1205
rect -605 1185 -597 1202
rect -580 1191 0 1202
rect -580 1185 -571 1191
rect -605 1181 -571 1185
rect 17355 1188 17370 1216
rect 17398 1188 17417 1216
rect 17445 1188 17464 1216
rect 17492 1213 18077 1216
rect 17492 1188 17898 1213
rect 17355 1181 17898 1188
rect 17930 1181 17942 1213
rect 17974 1181 17986 1213
rect 18018 1181 18030 1213
rect 18062 1181 18077 1213
rect 17355 1177 18077 1181
rect 20435 1168 20567 1181
rect -551 1131 -465 1134
rect -551 1111 -545 1131
rect -525 1111 -506 1131
rect -486 1128 -465 1131
rect 17527 1131 17613 1134
rect 17527 1128 17548 1131
rect -486 1114 0 1128
rect 17068 1114 17548 1128
rect -486 1111 -465 1114
rect -551 1108 -465 1111
rect 17527 1111 17548 1114
rect 17568 1111 17587 1131
rect 17607 1111 17613 1131
rect 17527 1108 17613 1111
rect -251 1096 0 1100
rect -251 1076 -245 1096
rect -225 1076 -206 1096
rect -186 1076 -167 1096
rect -147 1076 -128 1096
rect -108 1076 0 1096
rect -251 1072 0 1076
rect 17068 1096 17313 1100
rect 17068 1076 17170 1096
rect 17190 1076 17209 1096
rect 17229 1076 17248 1096
rect 17268 1076 17287 1096
rect 17307 1076 17313 1096
rect 17068 1072 17313 1076
rect 20435 962 20448 1168
rect 20554 962 20567 1168
rect -949 928 -943 954
rect -768 928 -762 954
rect -440 925 0 929
rect -440 905 -434 925
rect -414 905 -395 925
rect -375 905 -356 925
rect -336 905 -317 925
rect -297 905 0 925
rect -440 901 0 905
rect 17068 925 17503 929
rect 17644 928 17650 954
rect 17825 928 17831 954
rect 20435 950 20567 962
rect 20151 937 20319 946
rect 17068 905 17359 925
rect 17379 905 17398 925
rect 17418 905 17437 925
rect 17457 905 17476 925
rect 17496 905 17503 925
rect 17068 901 17503 905
rect -659 894 -625 897
rect -659 877 -651 894
rect -634 887 -625 894
rect -634 877 0 887
rect -659 873 0 877
rect 20151 862 20202 937
rect 20308 862 20319 937
rect 20151 855 20319 862
rect 17166 832 17837 833
rect 17166 825 17838 832
rect 17166 797 17180 825
rect 17208 797 17227 825
rect 17255 797 17274 825
rect 17302 819 17838 825
rect 17302 797 17659 819
rect 17166 787 17659 797
rect 17691 787 17703 819
rect 17735 787 17747 819
rect 17779 787 17791 819
rect 17823 787 17838 819
rect 17166 778 17838 787
rect -673 758 0 772
rect 17166 750 17180 778
rect 17208 750 17227 778
rect 17255 750 17274 778
rect 17302 774 17838 778
rect 17302 750 17659 774
rect 17166 742 17659 750
rect 17691 742 17703 774
rect 17735 742 17747 774
rect 17779 742 17791 774
rect 17823 742 17838 774
rect 17166 731 17838 742
rect -673 717 0 731
rect 17166 703 17180 731
rect 17208 703 17227 731
rect 17255 703 17274 731
rect 17302 729 17838 731
rect 17302 703 17659 729
rect -605 700 0 703
rect -605 683 -597 700
rect -580 689 0 700
rect 17166 697 17659 703
rect 17691 697 17703 729
rect 17735 697 17747 729
rect 17779 697 17791 729
rect 17823 697 17838 729
rect 17166 693 17838 697
rect -580 683 -571 689
rect -605 679 -571 683
rect 20151 666 20319 675
rect -551 629 -465 632
rect -551 609 -545 629
rect -525 609 -506 629
rect -486 626 -465 629
rect 17527 629 17613 632
rect 17527 626 17548 629
rect -486 612 0 626
rect 17068 612 17548 626
rect -486 609 -465 612
rect -551 606 -465 609
rect 17527 609 17548 612
rect 17568 609 17587 629
rect 17607 609 17613 629
rect 17527 606 17613 609
rect -251 594 0 598
rect -251 574 -245 594
rect -225 574 -206 594
rect -186 574 -167 594
rect -147 574 -128 594
rect -108 574 0 594
rect -251 570 0 574
rect 17068 594 17313 598
rect 17068 574 17170 594
rect 17190 574 17209 594
rect 17229 574 17248 594
rect 17268 574 17287 594
rect 17307 574 17313 594
rect 20151 591 20202 666
rect 20308 591 20319 666
rect 20151 584 20319 591
rect 17068 570 17313 574
rect -949 488 -943 514
rect -768 488 -762 514
rect 17644 488 17650 514
rect 17825 488 17831 514
rect -440 423 0 427
rect -440 403 -434 423
rect -414 403 -395 423
rect -375 403 -356 423
rect -336 403 -317 423
rect -297 403 0 423
rect -440 399 0 403
rect 17068 423 17503 427
rect 17068 403 17359 423
rect 17379 403 17398 423
rect 17418 403 17437 423
rect 17457 403 17476 423
rect 17496 403 17503 423
rect 17068 399 17503 403
rect 20151 388 20319 397
rect -440 381 0 385
rect -440 361 -434 381
rect -414 361 -395 381
rect -375 361 -356 381
rect -336 361 -317 381
rect -297 371 0 381
rect -297 361 -291 371
rect -440 357 -291 361
rect 17355 313 18077 320
rect 17355 285 17370 313
rect 17398 285 17417 313
rect 17445 285 17464 313
rect 17492 306 18077 313
rect 20151 313 20202 388
rect 20308 313 20319 388
rect 20151 306 20319 313
rect 17492 285 17898 306
rect 17355 274 17898 285
rect 17930 274 17942 306
rect 17974 274 17986 306
rect 18018 274 18030 306
rect 18062 274 18077 306
rect -251 256 0 270
rect 17355 266 18077 274
rect -251 253 -102 256
rect -251 233 -245 253
rect -225 233 -206 253
rect -186 233 -167 253
rect -147 233 -128 253
rect -108 233 -102 253
rect -251 229 -102 233
rect 17355 238 17370 266
rect 17398 238 17417 266
rect 17445 238 17464 266
rect 17492 261 18077 266
rect 17492 238 17898 261
rect 17355 229 17898 238
rect 17930 229 17942 261
rect 17974 229 17986 261
rect 18018 229 18030 261
rect 18062 229 18077 261
rect -251 215 0 229
rect 17355 219 18077 229
rect -251 197 0 201
rect -251 177 -245 197
rect -225 177 -206 197
rect -186 177 -167 197
rect -147 177 -128 197
rect -108 187 0 197
rect 17355 191 17370 219
rect 17398 191 17417 219
rect 17445 191 17464 219
rect 17492 216 18077 219
rect 17492 191 17898 216
rect -108 177 -102 187
rect 17355 184 17898 191
rect 17930 184 17942 216
rect 17974 184 17986 216
rect 18018 184 18030 216
rect 18062 184 18077 216
rect 17355 180 18077 184
rect 20435 289 20567 302
rect -251 173 -102 177
rect -551 127 -465 130
rect -551 107 -545 127
rect -525 107 -506 127
rect -486 124 -465 127
rect 17527 127 17613 130
rect 17527 124 17548 127
rect -486 110 0 124
rect 17068 110 17548 124
rect -486 107 -465 110
rect -551 104 -465 107
rect 17527 107 17548 110
rect 17568 107 17587 127
rect 17607 107 17613 127
rect 17527 104 17613 107
rect -251 92 0 96
rect -949 48 -943 74
rect -768 48 -762 74
rect -251 72 -245 92
rect -225 72 -206 92
rect -186 72 -167 92
rect -147 72 -128 92
rect -108 72 0 92
rect -251 68 0 72
rect 17068 92 17313 96
rect 17068 72 17170 92
rect 17190 72 17209 92
rect 17229 72 17248 92
rect 17268 72 17287 92
rect 17307 72 17313 92
rect 20435 83 20448 289
rect 20554 83 20567 289
rect 17068 68 17313 72
rect 17644 48 17650 74
rect 17825 48 17831 74
rect 20435 71 20567 83
rect 17146 -13 17838 -12
rect 17146 -20 17839 -13
rect 17146 -48 17181 -20
rect 17209 -48 17228 -20
rect 17256 -48 17275 -20
rect 17303 -26 17839 -20
rect 17303 -48 17660 -26
rect 17146 -58 17660 -48
rect 17692 -58 17704 -26
rect 17736 -58 17748 -26
rect 17780 -58 17792 -26
rect 17824 -58 17839 -26
rect 16098 -64 16371 -61
rect -956 -78 -750 -77
rect -957 -91 -750 -78
rect -957 -123 -942 -91
rect -910 -123 -898 -91
rect -866 -123 -854 -91
rect -822 -123 -810 -91
rect -778 -123 -750 -91
rect -957 -136 -750 -123
rect -957 -168 -942 -136
rect -910 -168 -898 -136
rect -866 -168 -854 -136
rect -822 -168 -810 -136
rect -778 -168 -750 -136
rect -957 -181 -750 -168
rect -957 -213 -942 -181
rect -910 -213 -898 -181
rect -866 -213 -854 -181
rect -822 -213 -810 -181
rect -778 -213 -750 -181
rect -957 -217 -750 -213
rect -273 -85 -91 -77
rect 16098 -81 16104 -64
rect 16121 -81 16348 -64
rect 16365 -81 16371 -64
rect 16098 -85 16371 -81
rect 17146 -67 17839 -58
rect -273 -113 -241 -85
rect -213 -113 -194 -85
rect -166 -113 -147 -85
rect -119 -113 -91 -85
rect -273 -132 -91 -113
rect -273 -160 -241 -132
rect -213 -160 -194 -132
rect -166 -160 -147 -132
rect -119 -160 -91 -132
rect 17146 -95 17181 -67
rect 17209 -95 17228 -67
rect 17256 -95 17275 -67
rect 17303 -71 17839 -67
rect 17303 -95 17660 -71
rect 17146 -103 17660 -95
rect 17692 -103 17704 -71
rect 17736 -103 17748 -71
rect 17780 -103 17792 -71
rect 17824 -103 17839 -71
rect 17146 -114 17839 -103
rect 13277 -136 14506 -133
rect 13277 -153 13283 -136
rect 13300 -153 14483 -136
rect 14500 -153 14506 -136
rect 17146 -142 17181 -114
rect 17209 -142 17228 -114
rect 17256 -142 17275 -114
rect 17303 -116 17839 -114
rect 17303 -142 17660 -116
rect 17146 -148 17660 -142
rect 17692 -148 17704 -116
rect 17736 -148 17748 -116
rect 17780 -148 17792 -116
rect 17824 -148 17839 -116
rect 17146 -152 17839 -148
rect 13277 -157 14506 -153
rect -273 -179 -91 -160
rect -273 -207 -241 -179
rect -213 -207 -194 -179
rect -166 -207 -147 -179
rect -119 -207 -91 -179
rect 13379 -175 15008 -172
rect 13379 -192 13385 -175
rect 13402 -192 14985 -175
rect 15002 -192 15008 -175
rect 13379 -196 15008 -192
rect 20151 -184 20567 -178
rect -273 -217 -91 -207
rect 13481 -213 15510 -210
rect 13481 -230 13487 -213
rect 13504 -230 15487 -213
rect 15504 -230 15510 -213
rect 13481 -234 15510 -230
rect 17146 -231 17503 -230
rect 17146 -238 18077 -231
rect 13583 -251 16012 -248
rect 13583 -268 13589 -251
rect 13606 -268 15989 -251
rect 16006 -268 16012 -251
rect 13583 -272 16012 -268
rect 17146 -266 17370 -238
rect 17398 -266 17417 -238
rect 17445 -266 17464 -238
rect 17492 -245 18077 -238
rect 17492 -266 17898 -245
rect 17146 -277 17898 -266
rect 17930 -277 17942 -245
rect 17974 -277 17986 -245
rect 18018 -277 18030 -245
rect 18062 -277 18077 -245
rect 20151 -265 20442 -184
rect 20561 -265 20567 -184
rect 20151 -270 20567 -265
rect 17146 -285 18077 -277
rect 13685 -289 16514 -286
rect 422 -295 448 -292
rect -385 -296 425 -295
rect -1195 -310 -988 -296
rect -1195 -342 -1180 -310
rect -1148 -342 -1136 -310
rect -1104 -342 -1092 -310
rect -1060 -342 -1048 -310
rect -1016 -342 -988 -310
rect -1195 -355 -988 -342
rect -1195 -387 -1180 -355
rect -1148 -387 -1136 -355
rect -1104 -387 -1092 -355
rect -1060 -387 -1048 -355
rect -1016 -387 -988 -355
rect -1195 -400 -988 -387
rect -1195 -432 -1180 -400
rect -1148 -432 -1136 -400
rect -1104 -432 -1092 -400
rect -1060 -432 -1048 -400
rect -1016 -432 -988 -400
rect -1195 -436 -988 -432
rect -462 -304 425 -296
rect -462 -332 -430 -304
rect -402 -332 -383 -304
rect -355 -332 -336 -304
rect -308 -312 425 -304
rect 442 -312 448 -295
rect 13685 -306 13691 -289
rect 13708 -306 16491 -289
rect 16508 -306 16514 -289
rect 17146 -295 17370 -285
rect 13685 -310 16514 -306
rect 16989 -298 17370 -295
rect -308 -316 448 -312
rect 16989 -315 16995 -298
rect 17012 -313 17370 -298
rect 17398 -313 17417 -285
rect 17445 -313 17464 -285
rect 17492 -290 18077 -285
rect 17492 -313 17898 -290
rect 17012 -315 17898 -313
rect -308 -332 -91 -316
rect 16989 -319 17898 -315
rect -462 -351 -91 -332
rect -462 -379 -430 -351
rect -402 -379 -383 -351
rect -355 -379 -336 -351
rect -308 -379 -91 -351
rect 17146 -322 17898 -319
rect 17930 -322 17942 -290
rect 17974 -322 17986 -290
rect 18018 -322 18030 -290
rect 18062 -322 18077 -290
rect 17146 -332 18077 -322
rect 17146 -360 17370 -332
rect 17398 -360 17417 -332
rect 17445 -360 17464 -332
rect 17492 -335 18077 -332
rect 17492 -360 17898 -335
rect 17146 -367 17898 -360
rect 17930 -367 17942 -335
rect 17974 -367 17986 -335
rect 18018 -367 18030 -335
rect 18062 -367 18077 -335
rect 17146 -371 18077 -367
rect -462 -398 -91 -379
rect -462 -426 -430 -398
rect -402 -426 -383 -398
rect -355 -426 -336 -398
rect -308 -426 -91 -398
rect -462 -435 -91 -426
rect 16395 -432 18196 -429
rect -462 -436 -280 -435
rect 16395 -449 16401 -432
rect 16418 -449 16437 -432
rect 16454 -449 18196 -432
rect 16395 -453 18196 -449
<< via1 >>
rect 20442 11290 20561 11371
rect 20448 10962 20554 11168
rect 20202 10862 20308 10937
rect 20202 10591 20308 10666
rect 20202 10313 20308 10388
rect 20448 10083 20554 10289
rect 20442 9735 20561 9816
rect 299 9516 430 9595
rect 1863 9516 1994 9595
rect 2299 9516 2430 9595
rect 3863 9516 3994 9595
rect 4299 9516 4430 9595
rect 5863 9516 5994 9595
rect 6299 9516 6430 9595
rect 7863 9516 7994 9595
rect 8299 9516 8430 9595
rect 9863 9516 9994 9595
rect 10299 9516 10430 9595
rect 11863 9516 11994 9595
rect 12299 9516 12430 9595
rect 13863 9516 13994 9595
rect 14299 9516 14430 9595
rect 15863 9516 15994 9595
rect 16299 9516 16430 9595
rect 17863 9533 17994 9595
rect -1180 9457 -1148 9489
rect -1136 9457 -1104 9489
rect -1092 9457 -1060 9489
rect -1048 9457 -1016 9489
rect -1180 9412 -1148 9444
rect -1136 9412 -1104 9444
rect -1092 9412 -1060 9444
rect -1048 9412 -1016 9444
rect -1180 9367 -1148 9399
rect -1136 9367 -1104 9399
rect -1092 9367 -1060 9399
rect -1048 9367 -1016 9399
rect 1072 9362 1235 9484
rect 3072 9362 3235 9484
rect 5072 9362 5235 9484
rect 7072 9362 7235 9484
rect 9072 9362 9235 9484
rect 11072 9362 11235 9484
rect 13072 9362 13235 9484
rect 15072 9362 15235 9484
rect 17072 9362 17235 9484
rect 17898 9457 17930 9489
rect 17942 9457 17974 9489
rect 17986 9457 18018 9489
rect 18030 9457 18062 9489
rect 17898 9412 17930 9444
rect 17942 9412 17974 9444
rect 17986 9412 18018 9444
rect 18030 9412 18062 9444
rect 17898 9367 17930 9399
rect 17942 9367 17974 9399
rect 17986 9367 18018 9399
rect 18030 9367 18062 9399
rect 20442 9290 20561 9371
rect -942 9238 -910 9270
rect -898 9238 -866 9270
rect -854 9238 -822 9270
rect -810 9238 -778 9270
rect 17660 9238 17692 9270
rect 17704 9238 17736 9270
rect 17748 9238 17780 9270
rect 17792 9238 17824 9270
rect -942 9193 -910 9225
rect -898 9193 -866 9225
rect -854 9193 -822 9225
rect -810 9193 -778 9225
rect 17660 9193 17692 9225
rect 17704 9193 17736 9225
rect 17748 9193 17780 9225
rect 17792 9193 17824 9225
rect -942 9148 -910 9180
rect -898 9148 -866 9180
rect -854 9148 -822 9180
rect -810 9148 -778 9180
rect 17660 9148 17692 9180
rect 17704 9148 17736 9180
rect 17748 9148 17780 9180
rect 17792 9148 17824 9180
rect 20448 8962 20554 9168
rect -943 8870 -768 8874
rect -943 8853 -768 8870
rect -943 8848 -768 8853
rect 17650 8870 17825 8874
rect 17650 8853 17825 8870
rect 17650 8848 17825 8853
rect 17661 8827 17693 8848
rect 17705 8827 17737 8848
rect 17749 8827 17781 8848
rect 17793 8827 17825 8848
rect 20202 8862 20308 8937
rect 17661 8782 17693 8814
rect 17705 8782 17737 8814
rect 17749 8782 17781 8814
rect 17793 8782 17825 8814
rect 17661 8737 17693 8769
rect 17705 8737 17737 8769
rect 17749 8737 17781 8769
rect 17793 8737 17825 8769
rect 20202 8591 20308 8666
rect -943 8430 -768 8434
rect -943 8413 -768 8430
rect -943 8408 -768 8413
rect 17650 8430 17825 8434
rect 17650 8413 17825 8430
rect 17650 8408 17825 8413
rect 17898 8334 17930 8366
rect 17942 8334 17974 8366
rect 17986 8334 18018 8366
rect 18030 8334 18062 8366
rect 17898 8289 17930 8321
rect 17942 8289 17974 8321
rect 17986 8289 18018 8321
rect 18030 8289 18062 8321
rect 20202 8313 20308 8388
rect 17898 8244 17930 8276
rect 17942 8244 17974 8276
rect 17986 8244 18018 8276
rect 18030 8244 18062 8276
rect 20448 8083 20554 8289
rect -943 7990 -768 7994
rect -943 7973 -768 7990
rect -943 7968 -768 7973
rect 17650 7990 17825 7994
rect 17650 7973 17825 7990
rect 17650 7968 17825 7973
rect 17660 7819 17692 7851
rect 17704 7819 17736 7851
rect 17748 7819 17780 7851
rect 17792 7819 17824 7851
rect 17660 7774 17692 7806
rect 17704 7774 17736 7806
rect 17748 7774 17780 7806
rect 17792 7774 17824 7806
rect 17660 7729 17692 7761
rect 17704 7729 17736 7761
rect 17748 7729 17780 7761
rect 17792 7729 17824 7761
rect 20442 7735 20561 7816
rect -943 7550 -768 7554
rect -943 7533 -768 7550
rect -943 7528 -768 7533
rect 17650 7550 17825 7554
rect 17650 7533 17825 7550
rect 17650 7528 17825 7533
rect 17898 7280 17930 7312
rect 17942 7280 17974 7312
rect 17986 7280 18018 7312
rect 18030 7280 18062 7312
rect 20442 7290 20561 7371
rect 17898 7235 17930 7267
rect 17942 7235 17974 7267
rect 17986 7235 18018 7267
rect 18030 7235 18062 7267
rect 17898 7190 17930 7222
rect 17942 7190 17974 7222
rect 17986 7190 18018 7222
rect 18030 7190 18062 7222
rect -943 7110 -768 7114
rect -943 7093 -768 7110
rect -943 7088 -768 7093
rect 17650 7110 17825 7114
rect 17650 7093 17825 7110
rect 17650 7088 17825 7093
rect 20448 6962 20554 7168
rect 20202 6862 20308 6937
rect 17660 6819 17692 6851
rect 17704 6819 17736 6851
rect 17748 6819 17780 6851
rect 17792 6819 17824 6851
rect 17660 6774 17692 6806
rect 17704 6774 17736 6806
rect 17748 6774 17780 6806
rect 17792 6774 17824 6806
rect 17660 6729 17692 6761
rect 17704 6729 17736 6761
rect 17748 6729 17780 6761
rect 17792 6729 17824 6761
rect -943 6670 -768 6674
rect -943 6653 -768 6670
rect -943 6648 -768 6653
rect 17650 6670 17825 6674
rect 17650 6653 17825 6670
rect 17650 6648 17825 6653
rect 20202 6591 20308 6666
rect 17897 6315 17929 6347
rect 17941 6315 17973 6347
rect 17985 6315 18017 6347
rect 18029 6315 18061 6347
rect 20202 6313 20308 6388
rect 17897 6270 17929 6302
rect 17941 6270 17973 6302
rect 17985 6270 18017 6302
rect 18029 6270 18061 6302
rect -943 6230 -768 6234
rect -943 6213 -768 6230
rect -943 6208 -768 6213
rect 17897 6225 17929 6257
rect 17941 6225 17973 6257
rect 17985 6225 18017 6257
rect 18029 6225 18061 6257
rect 20448 6083 20554 6289
rect 17661 5857 17693 5889
rect 17705 5857 17737 5889
rect 17749 5857 17781 5889
rect 17793 5857 17825 5889
rect 17661 5812 17693 5844
rect 17705 5812 17737 5844
rect 17749 5812 17781 5844
rect 17793 5812 17825 5844
rect -943 5790 -768 5794
rect -943 5773 -768 5790
rect -943 5768 -768 5773
rect 17661 5794 17693 5799
rect 17705 5794 17737 5799
rect 17749 5794 17781 5799
rect 17793 5794 17825 5799
rect 17650 5790 17825 5794
rect 17650 5773 17825 5790
rect 17650 5768 17825 5773
rect 17661 5767 17693 5768
rect 17705 5767 17737 5768
rect 17749 5767 17781 5768
rect 17793 5767 17825 5768
rect 20442 5735 20561 5816
rect -943 5350 -768 5354
rect -943 5333 -768 5350
rect -943 5328 -768 5333
rect 17898 5307 17930 5339
rect 17942 5307 17974 5339
rect 17986 5307 18018 5339
rect 18030 5307 18062 5339
rect 17898 5262 17930 5294
rect 17942 5262 17974 5294
rect 17986 5262 18018 5294
rect 18030 5262 18062 5294
rect 20442 5290 20561 5371
rect 17898 5217 17930 5249
rect 17942 5217 17974 5249
rect 17986 5217 18018 5249
rect 18030 5217 18062 5249
rect 20448 4962 20554 5168
rect -943 4910 -768 4914
rect -943 4893 -768 4910
rect -943 4888 -768 4893
rect 17650 4910 17825 4914
rect 17650 4893 17825 4910
rect 17650 4888 17825 4893
rect 20202 4862 20308 4937
rect 17660 4794 17692 4826
rect 17704 4794 17736 4826
rect 17748 4794 17780 4826
rect 17792 4794 17824 4826
rect 17660 4749 17692 4781
rect 17704 4749 17736 4781
rect 17748 4749 17780 4781
rect 17792 4749 17824 4781
rect 17660 4704 17692 4736
rect 17704 4704 17736 4736
rect 17748 4704 17780 4736
rect 17792 4704 17824 4736
rect 20202 4591 20308 4666
rect -943 4470 -768 4474
rect -943 4453 -768 4470
rect -943 4448 -768 4453
rect 17650 4470 17825 4474
rect 17650 4453 17825 4470
rect 17650 4448 17825 4453
rect 17898 4306 17930 4338
rect 17942 4306 17974 4338
rect 17986 4306 18018 4338
rect 18030 4306 18062 4338
rect 20202 4313 20308 4388
rect 17898 4261 17930 4293
rect 17942 4261 17974 4293
rect 17986 4261 18018 4293
rect 18030 4261 18062 4293
rect 17898 4216 17930 4248
rect 17942 4216 17974 4248
rect 17986 4216 18018 4248
rect 18030 4216 18062 4248
rect 20448 4083 20554 4289
rect -943 4030 -768 4034
rect -943 4013 -768 4030
rect -943 4008 -768 4013
rect 17650 4030 17825 4034
rect 17650 4013 17825 4030
rect 17650 4008 17825 4013
rect 17661 3806 17693 3838
rect 17705 3806 17737 3838
rect 17749 3806 17781 3838
rect 17793 3806 17825 3838
rect 17661 3761 17693 3793
rect 17705 3761 17737 3793
rect 17749 3761 17781 3793
rect 17793 3761 17825 3793
rect 17661 3716 17693 3748
rect 17705 3716 17737 3748
rect 17749 3716 17781 3748
rect 17793 3716 17825 3748
rect 20442 3735 20561 3816
rect -943 3590 -768 3594
rect -943 3573 -768 3590
rect -943 3568 -768 3573
rect 17650 3590 17825 3594
rect 17650 3573 17825 3590
rect 17650 3568 17825 3573
rect 17897 3307 17929 3339
rect 17941 3307 17973 3339
rect 17985 3307 18017 3339
rect 18029 3307 18061 3339
rect 17897 3262 17929 3294
rect 17941 3262 17973 3294
rect 17985 3262 18017 3294
rect 18029 3262 18061 3294
rect 20442 3290 20561 3371
rect 17897 3217 17929 3249
rect 17941 3217 17973 3249
rect 17985 3217 18017 3249
rect 18029 3217 18061 3249
rect -943 3150 -768 3154
rect -943 3133 -768 3150
rect -943 3128 -768 3133
rect 17650 3150 17825 3154
rect 17650 3133 17825 3150
rect 17650 3128 17825 3133
rect 20448 2962 20554 3168
rect 20202 2862 20308 2937
rect 17661 2784 17693 2816
rect 17705 2784 17737 2816
rect 17749 2784 17781 2816
rect 17793 2784 17825 2816
rect 17661 2739 17693 2771
rect 17705 2739 17737 2771
rect 17749 2739 17781 2771
rect 17793 2739 17825 2771
rect -943 2710 -768 2714
rect -943 2693 -768 2710
rect -943 2688 -768 2693
rect 17661 2714 17693 2726
rect 17705 2714 17737 2726
rect 17749 2714 17781 2726
rect 17793 2714 17825 2726
rect 17650 2710 17825 2714
rect 17650 2693 17825 2710
rect 17650 2688 17825 2693
rect 20202 2591 20308 2666
rect 20202 2313 20308 2388
rect -943 2270 -768 2274
rect -943 2253 -768 2270
rect -943 2248 -768 2253
rect 17898 2273 17930 2305
rect 17942 2273 17974 2305
rect 17986 2273 18018 2305
rect 18030 2273 18062 2305
rect 17898 2228 17930 2260
rect 17942 2228 17974 2260
rect 17986 2228 18018 2260
rect 18030 2228 18062 2260
rect 17898 2183 17930 2215
rect 17942 2183 17974 2215
rect 17986 2183 18018 2215
rect 18030 2183 18062 2215
rect 20448 2083 20554 2289
rect -943 1830 -768 1834
rect -943 1813 -768 1830
rect -943 1808 -768 1813
rect 17650 1830 17825 1834
rect 17650 1813 17825 1830
rect 17650 1808 17825 1813
rect 17661 1787 17693 1808
rect 17705 1787 17737 1808
rect 17749 1787 17781 1808
rect 17793 1787 17825 1808
rect 17661 1742 17693 1774
rect 17705 1742 17737 1774
rect 17749 1742 17781 1774
rect 17793 1742 17825 1774
rect 20442 1735 20561 1816
rect 17661 1697 17693 1729
rect 17705 1697 17737 1729
rect 17749 1697 17781 1729
rect 17793 1697 17825 1729
rect -943 1390 -768 1394
rect -943 1373 -768 1390
rect -943 1368 -768 1373
rect 17650 1390 17825 1394
rect 17650 1373 17825 1390
rect 17650 1368 17825 1373
rect 17898 1271 17930 1303
rect 17942 1271 17974 1303
rect 17986 1271 18018 1303
rect 18030 1271 18062 1303
rect 20442 1290 20561 1371
rect 17898 1226 17930 1258
rect 17942 1226 17974 1258
rect 17986 1226 18018 1258
rect 18030 1226 18062 1258
rect 17898 1181 17930 1213
rect 17942 1181 17974 1213
rect 17986 1181 18018 1213
rect 18030 1181 18062 1213
rect 20448 962 20554 1168
rect -943 950 -768 954
rect -943 933 -768 950
rect -943 928 -768 933
rect 17650 950 17825 954
rect 17650 933 17825 950
rect 17650 928 17825 933
rect 20202 862 20308 937
rect 17659 787 17691 819
rect 17703 787 17735 819
rect 17747 787 17779 819
rect 17791 787 17823 819
rect 17659 742 17691 774
rect 17703 742 17735 774
rect 17747 742 17779 774
rect 17791 742 17823 774
rect 17659 697 17691 729
rect 17703 697 17735 729
rect 17747 697 17779 729
rect 17791 697 17823 729
rect 20202 591 20308 666
rect -943 510 -768 514
rect -943 493 -768 510
rect -943 488 -768 493
rect 17650 510 17825 514
rect 17650 493 17825 510
rect 17650 488 17825 493
rect 20202 313 20308 388
rect 17898 274 17930 306
rect 17942 274 17974 306
rect 17986 274 18018 306
rect 18030 274 18062 306
rect 17898 229 17930 261
rect 17942 229 17974 261
rect 17986 229 18018 261
rect 18030 229 18062 261
rect 17898 184 17930 216
rect 17942 184 17974 216
rect 17986 184 18018 216
rect 18030 184 18062 216
rect -943 70 -768 74
rect -943 53 -768 70
rect -943 48 -768 53
rect 20448 83 20554 289
rect 17650 70 17825 74
rect 17650 53 17825 70
rect 17650 48 17825 53
rect 17660 -58 17692 -26
rect 17704 -58 17736 -26
rect 17748 -58 17780 -26
rect 17792 -58 17824 -26
rect -942 -123 -910 -91
rect -898 -123 -866 -91
rect -854 -123 -822 -91
rect -810 -123 -778 -91
rect -942 -168 -910 -136
rect -898 -168 -866 -136
rect -854 -168 -822 -136
rect -810 -168 -778 -136
rect -942 -213 -910 -181
rect -898 -213 -866 -181
rect -854 -213 -822 -181
rect -810 -213 -778 -181
rect -241 -113 -213 -85
rect -194 -113 -166 -85
rect -147 -113 -119 -85
rect -241 -160 -213 -132
rect -194 -160 -166 -132
rect -147 -160 -119 -132
rect 17660 -103 17692 -71
rect 17704 -103 17736 -71
rect 17748 -103 17780 -71
rect 17792 -103 17824 -71
rect 17660 -148 17692 -116
rect 17704 -148 17736 -116
rect 17748 -148 17780 -116
rect 17792 -148 17824 -116
rect -241 -207 -213 -179
rect -194 -207 -166 -179
rect -147 -207 -119 -179
rect 17898 -277 17930 -245
rect 17942 -277 17974 -245
rect 17986 -277 18018 -245
rect 18030 -277 18062 -245
rect 20442 -265 20561 -184
rect -1180 -342 -1148 -310
rect -1136 -342 -1104 -310
rect -1092 -342 -1060 -310
rect -1048 -342 -1016 -310
rect -1180 -387 -1148 -355
rect -1136 -387 -1104 -355
rect -1092 -387 -1060 -355
rect -1048 -387 -1016 -355
rect -1180 -432 -1148 -400
rect -1136 -432 -1104 -400
rect -1092 -432 -1060 -400
rect -1048 -432 -1016 -400
rect -430 -332 -402 -304
rect -383 -332 -355 -304
rect -336 -332 -308 -304
rect -430 -379 -402 -351
rect -383 -379 -355 -351
rect -336 -379 -308 -351
rect 17898 -322 17930 -290
rect 17942 -322 17974 -290
rect 17986 -322 18018 -290
rect 18030 -322 18062 -290
rect 17898 -367 17930 -335
rect 17942 -367 17974 -335
rect 17986 -367 18018 -335
rect 18030 -367 18062 -335
rect -430 -426 -402 -398
rect -383 -426 -355 -398
rect -336 -426 -308 -398
<< metal2 >>
rect 20151 11371 20567 11377
rect 20151 11290 20442 11371
rect 20561 11290 20567 11371
rect 20151 11285 20567 11290
rect 20435 11168 20567 11181
rect 20435 10962 20448 11168
rect 20554 10962 20567 11168
rect 20435 10950 20567 10962
rect 20151 10937 20319 10946
rect 20151 10862 20202 10937
rect 20308 10862 20319 10937
rect 20151 10855 20319 10862
rect 20151 10666 20319 10675
rect 20151 10591 20202 10666
rect 20308 10591 20319 10666
rect 20151 10584 20319 10591
rect 20151 10388 20319 10397
rect 20151 10313 20202 10388
rect 20308 10313 20319 10388
rect 20151 10306 20319 10313
rect 20435 10289 20567 10302
rect 20435 10083 20448 10289
rect 20554 10083 20567 10289
rect 20435 10071 20567 10083
rect 20151 9816 20567 9822
rect 20151 9735 20442 9816
rect 20561 9735 20567 9816
rect 20151 9730 20567 9735
rect 292 9595 438 9603
rect 292 9516 299 9595
rect 430 9516 438 9595
rect 292 9510 438 9516
rect 1856 9595 2002 9603
rect 1856 9516 1863 9595
rect 1994 9516 2002 9595
rect 1856 9510 2002 9516
rect 2292 9595 2438 9603
rect 2292 9516 2299 9595
rect 2430 9516 2438 9595
rect 2292 9510 2438 9516
rect 3856 9595 4002 9603
rect 3856 9516 3863 9595
rect 3994 9516 4002 9595
rect 3856 9510 4002 9516
rect 4292 9595 4438 9603
rect 4292 9516 4299 9595
rect 4430 9516 4438 9595
rect 4292 9510 4438 9516
rect 5856 9595 6002 9603
rect 5856 9516 5863 9595
rect 5994 9516 6002 9595
rect 5856 9510 6002 9516
rect 6292 9595 6438 9603
rect 6292 9516 6299 9595
rect 6430 9516 6438 9595
rect 6292 9510 6438 9516
rect 7856 9595 8002 9603
rect 7856 9516 7863 9595
rect 7994 9516 8002 9595
rect 7856 9510 8002 9516
rect 8292 9595 8438 9603
rect 8292 9516 8299 9595
rect 8430 9516 8438 9595
rect 8292 9510 8438 9516
rect 9856 9595 10002 9603
rect 9856 9516 9863 9595
rect 9994 9516 10002 9595
rect 9856 9510 10002 9516
rect 10292 9595 10438 9603
rect 10292 9516 10299 9595
rect 10430 9516 10438 9595
rect 10292 9510 10438 9516
rect 11856 9595 12002 9603
rect 11856 9516 11863 9595
rect 11994 9516 12002 9595
rect 11856 9510 12002 9516
rect 12292 9595 12438 9603
rect 12292 9516 12299 9595
rect 12430 9516 12438 9595
rect 12292 9510 12438 9516
rect 13856 9595 14002 9603
rect 13856 9516 13863 9595
rect 13994 9516 14002 9595
rect 13856 9510 14002 9516
rect 14292 9595 14438 9603
rect 14292 9516 14299 9595
rect 14430 9516 14438 9595
rect 14292 9510 14438 9516
rect 15856 9595 16002 9603
rect 15856 9516 15863 9595
rect 15994 9516 16002 9595
rect 15856 9510 16002 9516
rect 16292 9595 16438 9603
rect 16292 9516 16299 9595
rect 16430 9516 16438 9595
rect 17856 9595 18002 9603
rect 17856 9533 17863 9595
rect 17994 9533 18002 9595
rect 17856 9527 18002 9533
rect 16292 9510 16438 9516
rect -1195 9489 -988 9493
rect -1195 9457 -1180 9489
rect -1148 9457 -1136 9489
rect -1104 9457 -1092 9489
rect -1060 9457 -1048 9489
rect -1016 9457 -988 9489
rect -1195 9444 -988 9457
rect -1195 9412 -1180 9444
rect -1148 9412 -1136 9444
rect -1104 9412 -1092 9444
rect -1060 9412 -1048 9444
rect -1016 9412 -988 9444
rect -1195 9399 -988 9412
rect -1195 9367 -1180 9399
rect -1148 9367 -1136 9399
rect -1104 9367 -1092 9399
rect -1060 9367 -1048 9399
rect -1016 9367 -988 9399
rect -1195 9353 -988 9367
rect 1060 9484 1245 9493
rect 1060 9362 1072 9484
rect 1235 9362 1245 9484
rect 1060 9353 1245 9362
rect 3060 9484 3245 9493
rect 3060 9362 3072 9484
rect 3235 9362 3245 9484
rect 3060 9353 3245 9362
rect 5060 9484 5245 9493
rect 5060 9362 5072 9484
rect 5235 9362 5245 9484
rect 5060 9353 5245 9362
rect 7060 9484 7245 9493
rect 7060 9362 7072 9484
rect 7235 9362 7245 9484
rect 7060 9353 7245 9362
rect 9060 9484 9245 9493
rect 9060 9362 9072 9484
rect 9235 9362 9245 9484
rect 9060 9353 9245 9362
rect 11060 9484 11245 9493
rect 11060 9362 11072 9484
rect 11235 9362 11245 9484
rect 11060 9353 11245 9362
rect 13060 9484 13245 9493
rect 13060 9362 13072 9484
rect 13235 9362 13245 9484
rect 13060 9353 13245 9362
rect 15060 9484 15245 9493
rect 15060 9362 15072 9484
rect 15235 9362 15245 9484
rect 15060 9353 15245 9362
rect 17060 9484 17245 9493
rect 17060 9362 17072 9484
rect 17235 9362 17245 9484
rect 17060 9353 17245 9362
rect 17870 9489 18077 9493
rect 17870 9457 17898 9489
rect 17930 9457 17942 9489
rect 17974 9457 17986 9489
rect 18018 9457 18030 9489
rect 18062 9457 18077 9489
rect 17870 9444 18077 9457
rect 17870 9412 17898 9444
rect 17930 9412 17942 9444
rect 17974 9412 17986 9444
rect 18018 9412 18030 9444
rect 18062 9412 18077 9444
rect 17870 9399 18077 9412
rect 17870 9367 17898 9399
rect 17930 9367 17942 9399
rect 17974 9367 17986 9399
rect 18018 9367 18030 9399
rect 18062 9367 18077 9399
rect 17870 9353 18077 9367
rect 20151 9371 20567 9377
rect 20151 9290 20442 9371
rect 20561 9290 20567 9371
rect 20151 9285 20567 9290
rect -957 9270 -750 9274
rect -957 9238 -942 9270
rect -910 9238 -898 9270
rect -866 9238 -854 9270
rect -822 9238 -810 9270
rect -778 9238 -750 9270
rect -957 9225 -750 9238
rect -957 9193 -942 9225
rect -910 9193 -898 9225
rect -866 9193 -854 9225
rect -822 9193 -810 9225
rect -778 9193 -750 9225
rect -957 9180 -750 9193
rect -957 9148 -942 9180
rect -910 9148 -898 9180
rect -866 9148 -854 9180
rect -822 9148 -810 9180
rect -778 9148 -750 9180
rect -957 9134 -750 9148
rect 17632 9270 18151 9274
rect 17632 9238 17660 9270
rect 17692 9238 17704 9270
rect 17736 9238 17748 9270
rect 17780 9238 17792 9270
rect 17824 9238 18151 9270
rect 17632 9225 18151 9238
rect 17632 9193 17660 9225
rect 17692 9193 17704 9225
rect 17736 9193 17748 9225
rect 17780 9193 17792 9225
rect 17824 9193 18151 9225
rect 17632 9180 18151 9193
rect 17632 9148 17660 9180
rect 17692 9148 17704 9180
rect 17736 9148 17748 9180
rect 17780 9148 17792 9180
rect 17824 9148 18151 9180
rect 17632 9134 18151 9148
rect 20435 9168 20567 9181
rect 20435 8962 20448 9168
rect 20554 8962 20567 9168
rect 20435 8950 20567 8962
rect 20151 8937 20319 8946
rect -949 8847 -943 8875
rect -768 8847 -762 8875
rect 17644 8873 17650 8875
rect 17633 8847 17650 8873
rect 17825 8873 17831 8875
rect 17633 8827 17661 8847
rect 17693 8827 17705 8847
rect 17737 8827 17749 8847
rect 17781 8827 17793 8847
rect 17825 8827 17840 8873
rect 20151 8862 20202 8937
rect 20308 8862 20319 8937
rect 20151 8855 20319 8862
rect 17633 8814 17840 8827
rect 17633 8782 17661 8814
rect 17693 8782 17705 8814
rect 17737 8782 17749 8814
rect 17781 8782 17793 8814
rect 17825 8782 17840 8814
rect 17633 8769 17840 8782
rect 17633 8737 17661 8769
rect 17693 8737 17705 8769
rect 17737 8737 17749 8769
rect 17781 8737 17793 8769
rect 17825 8737 17840 8769
rect 17633 8733 17840 8737
rect 20151 8666 20319 8675
rect 20151 8591 20202 8666
rect 20308 8591 20319 8666
rect 20151 8584 20319 8591
rect -949 8407 -943 8435
rect -768 8407 -762 8435
rect 17644 8407 17650 8435
rect 17825 8407 17831 8435
rect 17870 8380 18151 8520
rect 20151 8388 20319 8397
rect 17870 8366 18077 8380
rect 17870 8334 17898 8366
rect 17930 8334 17942 8366
rect 17974 8334 17986 8366
rect 18018 8334 18030 8366
rect 18062 8334 18077 8366
rect 17870 8321 18077 8334
rect 17870 8289 17898 8321
rect 17930 8289 17942 8321
rect 17974 8289 17986 8321
rect 18018 8289 18030 8321
rect 18062 8289 18077 8321
rect 20151 8313 20202 8388
rect 20308 8313 20319 8388
rect 20151 8306 20319 8313
rect 17870 8276 18077 8289
rect 17870 8244 17898 8276
rect 17930 8244 17942 8276
rect 17974 8244 17986 8276
rect 18018 8244 18030 8276
rect 18062 8244 18077 8276
rect 17870 8240 18077 8244
rect 20435 8289 20567 8302
rect 20435 8083 20448 8289
rect 20554 8083 20567 8289
rect 20435 8071 20567 8083
rect -949 7967 -943 7995
rect -768 7967 -762 7995
rect 17644 7967 17650 7995
rect 17825 7967 17831 7995
rect 17632 7851 18151 7865
rect 17632 7819 17660 7851
rect 17692 7819 17704 7851
rect 17736 7819 17748 7851
rect 17780 7819 17792 7851
rect 17824 7819 18151 7851
rect 17632 7806 18151 7819
rect 17632 7774 17660 7806
rect 17692 7774 17704 7806
rect 17736 7774 17748 7806
rect 17780 7774 17792 7806
rect 17824 7774 18151 7806
rect 17632 7761 18151 7774
rect 17632 7729 17660 7761
rect 17692 7729 17704 7761
rect 17736 7729 17748 7761
rect 17780 7729 17792 7761
rect 17824 7729 18151 7761
rect 20151 7816 20567 7822
rect 20151 7735 20442 7816
rect 20561 7735 20567 7816
rect 20151 7730 20567 7735
rect 17632 7725 18151 7729
rect -949 7527 -943 7555
rect -768 7527 -762 7555
rect 17644 7527 17650 7555
rect 17825 7527 17831 7555
rect 20151 7371 20567 7377
rect 17870 7312 18077 7326
rect 17870 7280 17898 7312
rect 17930 7280 17942 7312
rect 17974 7280 17986 7312
rect 18018 7280 18030 7312
rect 18062 7280 18077 7312
rect 20151 7290 20442 7371
rect 20561 7290 20567 7371
rect 20151 7285 20567 7290
rect 17870 7267 18077 7280
rect 17870 7235 17898 7267
rect 17930 7235 17942 7267
rect 17974 7235 17986 7267
rect 18018 7235 18030 7267
rect 18062 7235 18077 7267
rect 17870 7222 18077 7235
rect 17870 7190 17898 7222
rect 17930 7190 17942 7222
rect 17974 7190 17986 7222
rect 18018 7190 18030 7222
rect 18062 7190 18077 7222
rect 17870 7186 18077 7190
rect 20435 7168 20567 7181
rect -949 7087 -943 7115
rect -768 7087 -762 7115
rect 17644 7087 17650 7115
rect 17825 7087 17831 7115
rect 20435 6962 20448 7168
rect 20554 6962 20567 7168
rect 20435 6950 20567 6962
rect 20151 6937 20319 6946
rect 17632 6851 17839 6865
rect 20151 6862 20202 6937
rect 20308 6862 20319 6937
rect 20151 6855 20319 6862
rect 17632 6819 17660 6851
rect 17692 6819 17704 6851
rect 17736 6819 17748 6851
rect 17780 6819 17792 6851
rect 17824 6819 17839 6851
rect 17632 6806 17839 6819
rect 17632 6774 17660 6806
rect 17692 6774 17704 6806
rect 17736 6774 17748 6806
rect 17780 6774 17792 6806
rect 17824 6774 17839 6806
rect 17632 6761 17839 6774
rect 17632 6729 17660 6761
rect 17692 6729 17704 6761
rect 17736 6729 17748 6761
rect 17780 6729 17792 6761
rect 17824 6729 17839 6761
rect 17632 6726 17839 6729
rect -949 6647 -943 6675
rect -768 6647 -762 6675
rect 17644 6647 17650 6675
rect 17825 6647 17831 6675
rect 20151 6666 20319 6675
rect 20151 6591 20202 6666
rect 20308 6591 20319 6666
rect 20151 6584 20319 6591
rect 17869 6361 18151 6502
rect 20151 6388 20319 6397
rect 17869 6347 18076 6361
rect 17869 6315 17897 6347
rect 17929 6315 17941 6347
rect 17973 6315 17985 6347
rect 18017 6315 18029 6347
rect 18061 6315 18076 6347
rect 17869 6302 18076 6315
rect 20151 6313 20202 6388
rect 20308 6313 20319 6388
rect 20151 6306 20319 6313
rect 17869 6270 17897 6302
rect 17929 6270 17941 6302
rect 17973 6270 17985 6302
rect 18017 6270 18029 6302
rect 18061 6270 18076 6302
rect 17869 6257 18076 6270
rect -949 6207 -943 6235
rect -768 6207 -762 6235
rect 17869 6225 17897 6257
rect 17929 6225 17941 6257
rect 17973 6225 17985 6257
rect 18017 6225 18029 6257
rect 18061 6225 18076 6257
rect 17869 6221 18076 6225
rect 20435 6289 20567 6302
rect 20435 6083 20448 6289
rect 20554 6083 20567 6289
rect 20435 6071 20567 6083
rect 17838 5903 18151 5904
rect 17633 5889 18151 5903
rect 17633 5857 17661 5889
rect 17693 5857 17705 5889
rect 17737 5857 17749 5889
rect 17781 5857 17793 5889
rect 17825 5857 18151 5889
rect 17633 5844 18151 5857
rect 17633 5812 17661 5844
rect 17693 5812 17705 5844
rect 17737 5812 17749 5844
rect 17781 5812 17793 5844
rect 17825 5812 18151 5844
rect 17633 5799 18151 5812
rect 17633 5795 17661 5799
rect -949 5767 -943 5795
rect -768 5767 -762 5795
rect 17633 5767 17650 5795
rect 17693 5795 17705 5799
rect 17737 5795 17749 5799
rect 17781 5795 17793 5799
rect 17825 5767 18151 5799
rect 17633 5763 18151 5767
rect 20151 5816 20567 5822
rect 20151 5735 20442 5816
rect 20561 5735 20567 5816
rect 20151 5730 20567 5735
rect 20151 5371 20567 5377
rect -949 5327 -943 5355
rect -768 5327 -762 5355
rect 17870 5339 18077 5353
rect 17870 5307 17898 5339
rect 17930 5307 17942 5339
rect 17974 5307 17986 5339
rect 18018 5307 18030 5339
rect 18062 5307 18077 5339
rect 17870 5294 18077 5307
rect 17870 5262 17898 5294
rect 17930 5262 17942 5294
rect 17974 5262 17986 5294
rect 18018 5262 18030 5294
rect 18062 5262 18077 5294
rect 20151 5290 20442 5371
rect 20561 5290 20567 5371
rect 20151 5285 20567 5290
rect 17870 5249 18077 5262
rect 17870 5217 17898 5249
rect 17930 5217 17942 5249
rect 17974 5217 17986 5249
rect 18018 5217 18030 5249
rect 18062 5217 18077 5249
rect 17870 5213 18077 5217
rect 20435 5168 20567 5181
rect 20435 4962 20448 5168
rect 20554 4962 20567 5168
rect 20435 4950 20567 4962
rect 20151 4937 20319 4946
rect -949 4887 -943 4915
rect -768 4887 -762 4915
rect 17644 4887 17650 4915
rect 17825 4887 17831 4915
rect 20151 4862 20202 4937
rect 20308 4862 20319 4937
rect 20151 4855 20319 4862
rect 17632 4826 17839 4840
rect 17632 4794 17660 4826
rect 17692 4794 17704 4826
rect 17736 4794 17748 4826
rect 17780 4794 17792 4826
rect 17824 4794 17839 4826
rect 17632 4781 17839 4794
rect 17632 4749 17660 4781
rect 17692 4749 17704 4781
rect 17736 4749 17748 4781
rect 17780 4749 17792 4781
rect 17824 4749 17839 4781
rect 17632 4736 17839 4749
rect 17632 4704 17660 4736
rect 17692 4704 17704 4736
rect 17736 4704 17748 4736
rect 17780 4704 17792 4736
rect 17824 4704 17839 4736
rect 17632 4700 17839 4704
rect 20151 4666 20319 4675
rect 20151 4591 20202 4666
rect 20308 4591 20319 4666
rect 20151 4584 20319 4591
rect -949 4447 -943 4475
rect -768 4447 -762 4475
rect 17644 4447 17650 4475
rect 17825 4447 17831 4475
rect 17870 4352 18151 4491
rect 20151 4388 20319 4397
rect 17870 4338 18077 4352
rect 17870 4306 17898 4338
rect 17930 4306 17942 4338
rect 17974 4306 17986 4338
rect 18018 4306 18030 4338
rect 18062 4306 18077 4338
rect 20151 4313 20202 4388
rect 20308 4313 20319 4388
rect 20151 4306 20319 4313
rect 17870 4293 18077 4306
rect 17870 4261 17898 4293
rect 17930 4261 17942 4293
rect 17974 4261 17986 4293
rect 18018 4261 18030 4293
rect 18062 4261 18077 4293
rect 17870 4248 18077 4261
rect 17870 4216 17898 4248
rect 17930 4216 17942 4248
rect 17974 4216 17986 4248
rect 18018 4216 18030 4248
rect 18062 4216 18077 4248
rect 17870 4212 18077 4216
rect 20435 4289 20567 4302
rect 20435 4083 20448 4289
rect 20554 4083 20567 4289
rect 20435 4071 20567 4083
rect -949 4007 -943 4035
rect -768 4007 -762 4035
rect 17644 4007 17650 4035
rect 17825 4007 17831 4035
rect 17633 3838 18151 3852
rect 17633 3806 17661 3838
rect 17693 3806 17705 3838
rect 17737 3806 17749 3838
rect 17781 3806 17793 3838
rect 17825 3806 18151 3838
rect 17633 3793 18151 3806
rect 17633 3761 17661 3793
rect 17693 3761 17705 3793
rect 17737 3761 17749 3793
rect 17781 3761 17793 3793
rect 17825 3761 18151 3793
rect 17633 3748 18151 3761
rect 17633 3716 17661 3748
rect 17693 3716 17705 3748
rect 17737 3716 17749 3748
rect 17781 3716 17793 3748
rect 17825 3716 18151 3748
rect 20151 3816 20567 3822
rect 20151 3735 20442 3816
rect 20561 3735 20567 3816
rect 20151 3730 20567 3735
rect 17633 3712 18151 3716
rect -949 3567 -943 3595
rect -768 3567 -762 3595
rect 17644 3567 17650 3595
rect 17825 3567 17831 3595
rect 20151 3371 20567 3377
rect 17869 3339 18076 3353
rect 17869 3307 17897 3339
rect 17929 3307 17941 3339
rect 17973 3307 17985 3339
rect 18017 3307 18029 3339
rect 18061 3307 18076 3339
rect 17869 3294 18076 3307
rect 17869 3262 17897 3294
rect 17929 3262 17941 3294
rect 17973 3262 17985 3294
rect 18017 3262 18029 3294
rect 18061 3262 18076 3294
rect 20151 3290 20442 3371
rect 20561 3290 20567 3371
rect 20151 3285 20567 3290
rect 17869 3249 18076 3262
rect 17869 3217 17897 3249
rect 17929 3217 17941 3249
rect 17973 3217 17985 3249
rect 18017 3217 18029 3249
rect 18061 3217 18076 3249
rect 17869 3213 18076 3217
rect 20435 3168 20567 3181
rect -949 3127 -943 3155
rect -768 3127 -762 3155
rect 17644 3127 17650 3155
rect 17825 3127 17831 3155
rect 20435 2962 20448 3168
rect 20554 2962 20567 3168
rect 20435 2950 20567 2962
rect 20151 2937 20319 2946
rect 20151 2862 20202 2937
rect 20308 2862 20319 2937
rect 20151 2855 20319 2862
rect 17633 2816 17840 2830
rect 17633 2784 17661 2816
rect 17693 2784 17705 2816
rect 17737 2784 17749 2816
rect 17781 2784 17793 2816
rect 17825 2784 17840 2816
rect 17633 2771 17840 2784
rect 17633 2739 17661 2771
rect 17693 2739 17705 2771
rect 17737 2739 17749 2771
rect 17781 2739 17793 2771
rect 17825 2739 17840 2771
rect 17633 2726 17840 2739
rect 17633 2715 17661 2726
rect -949 2687 -943 2715
rect -768 2687 -762 2715
rect 17633 2690 17650 2715
rect 17693 2715 17705 2726
rect 17737 2715 17749 2726
rect 17781 2715 17793 2726
rect 17644 2687 17650 2690
rect 17825 2690 17840 2726
rect 17825 2687 17831 2690
rect 20151 2666 20319 2675
rect 20151 2591 20202 2666
rect 20308 2591 20319 2666
rect 20151 2584 20319 2591
rect 17870 2319 18151 2458
rect 20151 2388 20319 2397
rect 17870 2305 18077 2319
rect 20151 2313 20202 2388
rect 20308 2313 20319 2388
rect 20151 2306 20319 2313
rect -949 2247 -943 2275
rect -768 2247 -762 2275
rect 17870 2273 17898 2305
rect 17930 2273 17942 2305
rect 17974 2273 17986 2305
rect 18018 2273 18030 2305
rect 18062 2273 18077 2305
rect 17870 2260 18077 2273
rect 17870 2228 17898 2260
rect 17930 2228 17942 2260
rect 17974 2228 17986 2260
rect 18018 2228 18030 2260
rect 18062 2228 18077 2260
rect 17870 2215 18077 2228
rect 17870 2183 17898 2215
rect 17930 2183 17942 2215
rect 17974 2183 17986 2215
rect 18018 2183 18030 2215
rect 18062 2183 18077 2215
rect 17870 2179 18077 2183
rect 20435 2289 20567 2302
rect 20435 2083 20448 2289
rect 20554 2083 20567 2289
rect 20435 2071 20567 2083
rect -949 1807 -943 1835
rect -768 1807 -762 1835
rect 17644 1833 17650 1835
rect 17633 1807 17650 1833
rect 17825 1833 17831 1835
rect 17633 1787 17661 1807
rect 17693 1787 17705 1807
rect 17737 1787 17749 1807
rect 17781 1787 17793 1807
rect 17825 1787 18151 1833
rect 17633 1774 18151 1787
rect 17633 1742 17661 1774
rect 17693 1742 17705 1774
rect 17737 1742 17749 1774
rect 17781 1742 17793 1774
rect 17825 1742 18151 1774
rect 17633 1729 18151 1742
rect 20151 1816 20567 1822
rect 20151 1735 20442 1816
rect 20561 1735 20567 1816
rect 20151 1730 20567 1735
rect 17633 1697 17661 1729
rect 17693 1697 17705 1729
rect 17737 1697 17749 1729
rect 17781 1697 17793 1729
rect 17825 1697 18151 1729
rect 17633 1693 18151 1697
rect -949 1367 -943 1395
rect -768 1367 -762 1395
rect 17644 1367 17650 1395
rect 17825 1367 17831 1395
rect 20151 1371 20567 1377
rect 17870 1303 18077 1317
rect 17870 1271 17898 1303
rect 17930 1271 17942 1303
rect 17974 1271 17986 1303
rect 18018 1271 18030 1303
rect 18062 1271 18077 1303
rect 20151 1290 20442 1371
rect 20561 1290 20567 1371
rect 20151 1285 20567 1290
rect 17870 1258 18077 1271
rect 17870 1226 17898 1258
rect 17930 1226 17942 1258
rect 17974 1226 17986 1258
rect 18018 1226 18030 1258
rect 18062 1226 18077 1258
rect 17870 1213 18077 1226
rect 17870 1181 17898 1213
rect 17930 1181 17942 1213
rect 17974 1181 17986 1213
rect 18018 1181 18030 1213
rect 18062 1181 18077 1213
rect 17870 1177 18077 1181
rect 20435 1168 20567 1181
rect 20435 962 20448 1168
rect 20554 962 20567 1168
rect -949 927 -943 955
rect -768 927 -762 955
rect 17644 927 17650 955
rect 17825 927 17831 955
rect 20435 950 20567 962
rect 20151 937 20319 946
rect 20151 862 20202 937
rect 20308 862 20319 937
rect 20151 855 20319 862
rect 17631 819 17838 833
rect 17631 787 17659 819
rect 17691 787 17703 819
rect 17735 787 17747 819
rect 17779 787 17791 819
rect 17823 787 17838 819
rect 17631 774 17838 787
rect 17631 742 17659 774
rect 17691 742 17703 774
rect 17735 742 17747 774
rect 17779 742 17791 774
rect 17823 742 17838 774
rect 17631 729 17838 742
rect 17631 697 17659 729
rect 17691 697 17703 729
rect 17735 697 17747 729
rect 17779 697 17791 729
rect 17823 697 17838 729
rect 17631 693 17838 697
rect 20151 666 20319 675
rect 20151 591 20202 666
rect 20308 591 20319 666
rect 20151 584 20319 591
rect -949 487 -943 515
rect -768 487 -762 515
rect 17644 487 17650 515
rect 17825 487 17831 515
rect 17870 319 18151 440
rect 20151 388 20319 397
rect 17870 306 18077 319
rect 20151 313 20202 388
rect 20308 313 20319 388
rect 20151 306 20319 313
rect 17870 274 17898 306
rect 17930 274 17942 306
rect 17974 274 17986 306
rect 18018 274 18030 306
rect 18062 274 18077 306
rect 17870 261 18077 274
rect 17870 229 17898 261
rect 17930 229 17942 261
rect 17974 229 17986 261
rect 18018 229 18030 261
rect 18062 229 18077 261
rect 17870 216 18077 229
rect 17870 184 17898 216
rect 17930 184 17942 216
rect 17974 184 17986 216
rect 18018 184 18030 216
rect 18062 184 18077 216
rect 17870 180 18077 184
rect 20435 289 20567 302
rect 20435 83 20448 289
rect 20554 83 20567 289
rect -949 47 -943 75
rect -768 47 -762 75
rect 17644 47 17650 75
rect 17825 47 17831 75
rect 20435 71 20567 83
rect 17632 -26 18151 -12
rect 17632 -58 17660 -26
rect 17692 -58 17704 -26
rect 17736 -58 17748 -26
rect 17780 -58 17792 -26
rect 17824 -58 18151 -26
rect 17632 -71 18151 -58
rect -957 -91 -750 -77
rect -957 -123 -942 -91
rect -910 -123 -898 -91
rect -866 -123 -854 -91
rect -822 -123 -810 -91
rect -778 -123 -750 -91
rect -957 -136 -750 -123
rect -957 -168 -942 -136
rect -910 -168 -898 -136
rect -866 -168 -854 -136
rect -822 -168 -810 -136
rect -778 -168 -750 -136
rect -957 -181 -750 -168
rect -957 -213 -942 -181
rect -910 -213 -898 -181
rect -866 -213 -854 -181
rect -822 -213 -810 -181
rect -778 -213 -750 -181
rect -957 -217 -750 -213
rect -273 -85 -91 -76
rect -273 -113 -241 -85
rect -213 -113 -194 -85
rect -166 -113 -147 -85
rect -119 -113 -91 -85
rect -273 -132 -91 -113
rect -273 -160 -241 -132
rect -213 -160 -194 -132
rect -166 -160 -147 -132
rect -119 -160 -91 -132
rect 17632 -103 17660 -71
rect 17692 -103 17704 -71
rect 17736 -103 17748 -71
rect 17780 -103 17792 -71
rect 17824 -103 18151 -71
rect 17632 -116 18151 -103
rect 17632 -148 17660 -116
rect 17692 -148 17704 -116
rect 17736 -148 17748 -116
rect 17780 -148 17792 -116
rect 17824 -148 18151 -116
rect 17632 -152 18151 -148
rect -273 -179 -91 -160
rect -273 -207 -241 -179
rect -213 -207 -194 -179
rect -166 -207 -147 -179
rect -119 -207 -91 -179
rect -273 -217 -91 -207
rect 20151 -184 20567 -178
rect 17870 -245 18077 -231
rect 17870 -277 17898 -245
rect 17930 -277 17942 -245
rect 17974 -277 17986 -245
rect 18018 -277 18030 -245
rect 18062 -277 18077 -245
rect 20151 -265 20442 -184
rect 20561 -265 20567 -184
rect 20151 -270 20567 -265
rect 17870 -290 18077 -277
rect -1195 -310 -988 -296
rect -1195 -342 -1180 -310
rect -1148 -342 -1136 -310
rect -1104 -342 -1092 -310
rect -1060 -342 -1048 -310
rect -1016 -342 -988 -310
rect -1195 -355 -988 -342
rect -1195 -387 -1180 -355
rect -1148 -387 -1136 -355
rect -1104 -387 -1092 -355
rect -1060 -387 -1048 -355
rect -1016 -387 -988 -355
rect -1195 -400 -988 -387
rect -1195 -432 -1180 -400
rect -1148 -432 -1136 -400
rect -1104 -432 -1092 -400
rect -1060 -432 -1048 -400
rect -1016 -432 -988 -400
rect -1195 -436 -988 -432
rect -462 -304 -280 -295
rect -462 -332 -430 -304
rect -402 -332 -383 -304
rect -355 -332 -336 -304
rect -308 -332 -280 -304
rect -462 -351 -280 -332
rect -462 -379 -430 -351
rect -402 -379 -383 -351
rect -355 -379 -336 -351
rect -308 -379 -280 -351
rect 17870 -322 17898 -290
rect 17930 -322 17942 -290
rect 17974 -322 17986 -290
rect 18018 -322 18030 -290
rect 18062 -322 18077 -290
rect 17870 -335 18077 -322
rect 17870 -367 17898 -335
rect 17930 -367 17942 -335
rect 17974 -367 17986 -335
rect 18018 -367 18030 -335
rect 18062 -367 18077 -335
rect 17870 -371 18077 -367
rect -462 -398 -280 -379
rect -462 -426 -430 -398
rect -402 -426 -383 -398
rect -355 -426 -336 -398
rect -308 -426 -280 -398
rect -462 -436 -280 -426
<< via2 >>
rect 20442 11290 20561 11371
rect 20448 10962 20554 11168
rect 20202 10862 20308 10937
rect 20202 10591 20308 10666
rect 20202 10313 20308 10388
rect 20448 10083 20554 10289
rect 20442 9735 20561 9816
rect 299 9516 430 9595
rect 1863 9516 1994 9595
rect 2299 9516 2430 9595
rect 3863 9516 3994 9595
rect 4299 9516 4430 9595
rect 5863 9516 5994 9595
rect 6299 9516 6430 9595
rect 7863 9516 7994 9595
rect 8299 9516 8430 9595
rect 9863 9516 9994 9595
rect 10299 9516 10430 9595
rect 11863 9516 11994 9595
rect 12299 9516 12430 9595
rect 13863 9516 13994 9595
rect 14299 9516 14430 9595
rect 15863 9516 15994 9595
rect 16299 9516 16430 9595
rect 17863 9533 17994 9595
rect -1180 9457 -1148 9489
rect -1136 9457 -1104 9489
rect -1092 9457 -1060 9489
rect -1048 9457 -1016 9489
rect -1180 9412 -1148 9444
rect -1136 9412 -1104 9444
rect -1092 9412 -1060 9444
rect -1048 9412 -1016 9444
rect -1180 9367 -1148 9399
rect -1136 9367 -1104 9399
rect -1092 9367 -1060 9399
rect -1048 9367 -1016 9399
rect 1072 9362 1235 9484
rect 3072 9362 3235 9484
rect 5072 9362 5235 9484
rect 7072 9362 7235 9484
rect 9072 9362 9235 9484
rect 11072 9362 11235 9484
rect 13072 9362 13235 9484
rect 15072 9362 15235 9484
rect 17072 9362 17235 9484
rect 17898 9457 17930 9489
rect 17942 9457 17974 9489
rect 17986 9457 18018 9489
rect 18030 9457 18062 9489
rect 17898 9412 17930 9444
rect 17942 9412 17974 9444
rect 17986 9412 18018 9444
rect 18030 9412 18062 9444
rect 17898 9367 17930 9399
rect 17942 9367 17974 9399
rect 17986 9367 18018 9399
rect 18030 9367 18062 9399
rect 20442 9290 20561 9371
rect -942 9238 -910 9270
rect -898 9238 -866 9270
rect -854 9238 -822 9270
rect -810 9238 -778 9270
rect -942 9193 -910 9225
rect -898 9193 -866 9225
rect -854 9193 -822 9225
rect -810 9193 -778 9225
rect -942 9148 -910 9180
rect -898 9148 -866 9180
rect -854 9148 -822 9180
rect -810 9148 -778 9180
rect 17660 9238 17692 9270
rect 17704 9238 17736 9270
rect 17748 9238 17780 9270
rect 17792 9238 17824 9270
rect 17660 9193 17692 9225
rect 17704 9193 17736 9225
rect 17748 9193 17780 9225
rect 17792 9193 17824 9225
rect 17660 9148 17692 9180
rect 17704 9148 17736 9180
rect 17748 9148 17780 9180
rect 17792 9148 17824 9180
rect 20448 8962 20554 9168
rect -943 8874 -768 8875
rect -943 8848 -768 8874
rect -943 8847 -768 8848
rect 17650 8874 17825 8875
rect 17650 8848 17825 8874
rect 17650 8847 17661 8848
rect 17661 8827 17693 8848
rect 17693 8847 17705 8848
rect 17705 8827 17737 8848
rect 17737 8847 17749 8848
rect 17749 8827 17781 8848
rect 17781 8847 17793 8848
rect 17793 8827 17825 8848
rect 20202 8862 20308 8937
rect 17661 8782 17693 8814
rect 17705 8782 17737 8814
rect 17749 8782 17781 8814
rect 17793 8782 17825 8814
rect 17661 8737 17693 8769
rect 17705 8737 17737 8769
rect 17749 8737 17781 8769
rect 17793 8737 17825 8769
rect 20202 8591 20308 8666
rect -943 8434 -768 8435
rect -943 8408 -768 8434
rect -943 8407 -768 8408
rect 17650 8434 17825 8435
rect 17650 8408 17825 8434
rect 17650 8407 17825 8408
rect 17898 8334 17930 8366
rect 17942 8334 17974 8366
rect 17986 8334 18018 8366
rect 18030 8334 18062 8366
rect 17898 8289 17930 8321
rect 17942 8289 17974 8321
rect 17986 8289 18018 8321
rect 18030 8289 18062 8321
rect 20202 8313 20308 8388
rect 17898 8244 17930 8276
rect 17942 8244 17974 8276
rect 17986 8244 18018 8276
rect 18030 8244 18062 8276
rect 20448 8083 20554 8289
rect -943 7994 -768 7995
rect -943 7968 -768 7994
rect -943 7967 -768 7968
rect 17650 7994 17825 7995
rect 17650 7968 17825 7994
rect 17650 7967 17825 7968
rect 17660 7819 17692 7851
rect 17704 7819 17736 7851
rect 17748 7819 17780 7851
rect 17792 7819 17824 7851
rect 17660 7774 17692 7806
rect 17704 7774 17736 7806
rect 17748 7774 17780 7806
rect 17792 7774 17824 7806
rect 17660 7729 17692 7761
rect 17704 7729 17736 7761
rect 17748 7729 17780 7761
rect 17792 7729 17824 7761
rect 20442 7735 20561 7816
rect -943 7554 -768 7555
rect -943 7528 -768 7554
rect -943 7527 -768 7528
rect 17650 7554 17825 7555
rect 17650 7528 17825 7554
rect 17650 7527 17825 7528
rect 17898 7280 17930 7312
rect 17942 7280 17974 7312
rect 17986 7280 18018 7312
rect 18030 7280 18062 7312
rect 20442 7290 20561 7371
rect 17898 7235 17930 7267
rect 17942 7235 17974 7267
rect 17986 7235 18018 7267
rect 18030 7235 18062 7267
rect 17898 7190 17930 7222
rect 17942 7190 17974 7222
rect 17986 7190 18018 7222
rect 18030 7190 18062 7222
rect -943 7114 -768 7115
rect -943 7088 -768 7114
rect -943 7087 -768 7088
rect 17650 7114 17825 7115
rect 17650 7088 17825 7114
rect 17650 7087 17825 7088
rect 20448 6962 20554 7168
rect 20202 6862 20308 6937
rect 17660 6819 17692 6851
rect 17704 6819 17736 6851
rect 17748 6819 17780 6851
rect 17792 6819 17824 6851
rect 17660 6774 17692 6806
rect 17704 6774 17736 6806
rect 17748 6774 17780 6806
rect 17792 6774 17824 6806
rect 17660 6729 17692 6761
rect 17704 6729 17736 6761
rect 17748 6729 17780 6761
rect 17792 6729 17824 6761
rect -943 6674 -768 6675
rect -943 6648 -768 6674
rect -943 6647 -768 6648
rect 17650 6674 17825 6675
rect 17650 6648 17825 6674
rect 17650 6647 17825 6648
rect 20202 6591 20308 6666
rect 17897 6315 17929 6347
rect 17941 6315 17973 6347
rect 17985 6315 18017 6347
rect 18029 6315 18061 6347
rect 20202 6313 20308 6388
rect 17897 6270 17929 6302
rect 17941 6270 17973 6302
rect 17985 6270 18017 6302
rect 18029 6270 18061 6302
rect -943 6234 -768 6235
rect -943 6208 -768 6234
rect -943 6207 -768 6208
rect 17897 6225 17929 6257
rect 17941 6225 17973 6257
rect 17985 6225 18017 6257
rect 18029 6225 18061 6257
rect 20448 6083 20554 6289
rect 17661 5857 17693 5889
rect 17705 5857 17737 5889
rect 17749 5857 17781 5889
rect 17793 5857 17825 5889
rect 17661 5812 17693 5844
rect 17705 5812 17737 5844
rect 17749 5812 17781 5844
rect 17793 5812 17825 5844
rect -943 5794 -768 5795
rect -943 5768 -768 5794
rect -943 5767 -768 5768
rect 17650 5794 17661 5795
rect 17661 5794 17693 5799
rect 17693 5794 17705 5795
rect 17705 5794 17737 5799
rect 17737 5794 17749 5795
rect 17749 5794 17781 5799
rect 17781 5794 17793 5795
rect 17793 5794 17825 5799
rect 17650 5768 17825 5794
rect 17650 5767 17661 5768
rect 17661 5767 17693 5768
rect 17693 5767 17705 5768
rect 17705 5767 17737 5768
rect 17737 5767 17749 5768
rect 17749 5767 17781 5768
rect 17781 5767 17793 5768
rect 17793 5767 17825 5768
rect 20442 5735 20561 5816
rect -943 5354 -768 5355
rect -943 5328 -768 5354
rect -943 5327 -768 5328
rect 17898 5307 17930 5339
rect 17942 5307 17974 5339
rect 17986 5307 18018 5339
rect 18030 5307 18062 5339
rect 17898 5262 17930 5294
rect 17942 5262 17974 5294
rect 17986 5262 18018 5294
rect 18030 5262 18062 5294
rect 20442 5290 20561 5371
rect 17898 5217 17930 5249
rect 17942 5217 17974 5249
rect 17986 5217 18018 5249
rect 18030 5217 18062 5249
rect 20448 4962 20554 5168
rect -943 4914 -768 4915
rect -943 4888 -768 4914
rect -943 4887 -768 4888
rect 17650 4914 17825 4915
rect 17650 4888 17825 4914
rect 17650 4887 17825 4888
rect 20202 4862 20308 4937
rect 17660 4794 17692 4826
rect 17704 4794 17736 4826
rect 17748 4794 17780 4826
rect 17792 4794 17824 4826
rect 17660 4749 17692 4781
rect 17704 4749 17736 4781
rect 17748 4749 17780 4781
rect 17792 4749 17824 4781
rect 17660 4704 17692 4736
rect 17704 4704 17736 4736
rect 17748 4704 17780 4736
rect 17792 4704 17824 4736
rect 20202 4591 20308 4666
rect -943 4474 -768 4475
rect -943 4448 -768 4474
rect -943 4447 -768 4448
rect 17650 4474 17825 4475
rect 17650 4448 17825 4474
rect 17650 4447 17825 4448
rect 17898 4306 17930 4338
rect 17942 4306 17974 4338
rect 17986 4306 18018 4338
rect 18030 4306 18062 4338
rect 20202 4313 20308 4388
rect 17898 4261 17930 4293
rect 17942 4261 17974 4293
rect 17986 4261 18018 4293
rect 18030 4261 18062 4293
rect 17898 4216 17930 4248
rect 17942 4216 17974 4248
rect 17986 4216 18018 4248
rect 18030 4216 18062 4248
rect 20448 4083 20554 4289
rect -943 4034 -768 4035
rect -943 4008 -768 4034
rect -943 4007 -768 4008
rect 17650 4034 17825 4035
rect 17650 4008 17825 4034
rect 17650 4007 17825 4008
rect 17661 3806 17693 3838
rect 17705 3806 17737 3838
rect 17749 3806 17781 3838
rect 17793 3806 17825 3838
rect 17661 3761 17693 3793
rect 17705 3761 17737 3793
rect 17749 3761 17781 3793
rect 17793 3761 17825 3793
rect 17661 3716 17693 3748
rect 17705 3716 17737 3748
rect 17749 3716 17781 3748
rect 17793 3716 17825 3748
rect 20442 3735 20561 3816
rect -943 3594 -768 3595
rect -943 3568 -768 3594
rect -943 3567 -768 3568
rect 17650 3594 17825 3595
rect 17650 3568 17825 3594
rect 17650 3567 17825 3568
rect 17897 3307 17929 3339
rect 17941 3307 17973 3339
rect 17985 3307 18017 3339
rect 18029 3307 18061 3339
rect 17897 3262 17929 3294
rect 17941 3262 17973 3294
rect 17985 3262 18017 3294
rect 18029 3262 18061 3294
rect 20442 3290 20561 3371
rect 17897 3217 17929 3249
rect 17941 3217 17973 3249
rect 17985 3217 18017 3249
rect 18029 3217 18061 3249
rect -943 3154 -768 3155
rect -943 3128 -768 3154
rect -943 3127 -768 3128
rect 17650 3154 17825 3155
rect 17650 3128 17825 3154
rect 17650 3127 17825 3128
rect 20448 2962 20554 3168
rect 20202 2862 20308 2937
rect 17661 2784 17693 2816
rect 17705 2784 17737 2816
rect 17749 2784 17781 2816
rect 17793 2784 17825 2816
rect 17661 2739 17693 2771
rect 17705 2739 17737 2771
rect 17749 2739 17781 2771
rect 17793 2739 17825 2771
rect -943 2714 -768 2715
rect -943 2688 -768 2714
rect -943 2687 -768 2688
rect 17650 2714 17661 2715
rect 17661 2714 17693 2726
rect 17693 2714 17705 2715
rect 17705 2714 17737 2726
rect 17737 2714 17749 2715
rect 17749 2714 17781 2726
rect 17781 2714 17793 2715
rect 17793 2714 17825 2726
rect 17650 2688 17825 2714
rect 17650 2687 17825 2688
rect 20202 2591 20308 2666
rect 20202 2313 20308 2388
rect -943 2274 -768 2275
rect -943 2248 -768 2274
rect -943 2247 -768 2248
rect 17898 2273 17930 2305
rect 17942 2273 17974 2305
rect 17986 2273 18018 2305
rect 18030 2273 18062 2305
rect 17898 2228 17930 2260
rect 17942 2228 17974 2260
rect 17986 2228 18018 2260
rect 18030 2228 18062 2260
rect 17898 2183 17930 2215
rect 17942 2183 17974 2215
rect 17986 2183 18018 2215
rect 18030 2183 18062 2215
rect 20448 2083 20554 2289
rect -943 1834 -768 1835
rect -943 1808 -768 1834
rect -943 1807 -768 1808
rect 17650 1834 17825 1835
rect 17650 1808 17825 1834
rect 17650 1807 17661 1808
rect 17661 1787 17693 1808
rect 17693 1807 17705 1808
rect 17705 1787 17737 1808
rect 17737 1807 17749 1808
rect 17749 1787 17781 1808
rect 17781 1807 17793 1808
rect 17793 1787 17825 1808
rect 17661 1742 17693 1774
rect 17705 1742 17737 1774
rect 17749 1742 17781 1774
rect 17793 1742 17825 1774
rect 20442 1735 20561 1816
rect 17661 1697 17693 1729
rect 17705 1697 17737 1729
rect 17749 1697 17781 1729
rect 17793 1697 17825 1729
rect -943 1394 -768 1395
rect -943 1368 -768 1394
rect -943 1367 -768 1368
rect 17650 1394 17825 1395
rect 17650 1368 17825 1394
rect 17650 1367 17825 1368
rect 17898 1271 17930 1303
rect 17942 1271 17974 1303
rect 17986 1271 18018 1303
rect 18030 1271 18062 1303
rect 20442 1290 20561 1371
rect 17898 1226 17930 1258
rect 17942 1226 17974 1258
rect 17986 1226 18018 1258
rect 18030 1226 18062 1258
rect 17898 1181 17930 1213
rect 17942 1181 17974 1213
rect 17986 1181 18018 1213
rect 18030 1181 18062 1213
rect 20448 962 20554 1168
rect -943 954 -768 955
rect -943 928 -768 954
rect -943 927 -768 928
rect 17650 954 17825 955
rect 17650 928 17825 954
rect 17650 927 17825 928
rect 20202 862 20308 937
rect 17659 787 17691 819
rect 17703 787 17735 819
rect 17747 787 17779 819
rect 17791 787 17823 819
rect 17659 742 17691 774
rect 17703 742 17735 774
rect 17747 742 17779 774
rect 17791 742 17823 774
rect 17659 697 17691 729
rect 17703 697 17735 729
rect 17747 697 17779 729
rect 17791 697 17823 729
rect 20202 591 20308 666
rect -943 514 -768 515
rect -943 488 -768 514
rect -943 487 -768 488
rect 17650 514 17825 515
rect 17650 488 17825 514
rect 17650 487 17825 488
rect 20202 313 20308 388
rect 17898 274 17930 306
rect 17942 274 17974 306
rect 17986 274 18018 306
rect 18030 274 18062 306
rect 17898 229 17930 261
rect 17942 229 17974 261
rect 17986 229 18018 261
rect 18030 229 18062 261
rect 17898 184 17930 216
rect 17942 184 17974 216
rect 17986 184 18018 216
rect 18030 184 18062 216
rect 20448 83 20554 289
rect -943 74 -768 75
rect -943 48 -768 74
rect -943 47 -768 48
rect 17650 74 17825 75
rect 17650 48 17825 74
rect 17650 47 17825 48
rect 17660 -58 17692 -26
rect 17704 -58 17736 -26
rect 17748 -58 17780 -26
rect 17792 -58 17824 -26
rect -942 -123 -910 -91
rect -898 -123 -866 -91
rect -854 -123 -822 -91
rect -810 -123 -778 -91
rect -942 -168 -910 -136
rect -898 -168 -866 -136
rect -854 -168 -822 -136
rect -810 -168 -778 -136
rect -942 -213 -910 -181
rect -898 -213 -866 -181
rect -854 -213 -822 -181
rect -810 -213 -778 -181
rect -241 -113 -213 -85
rect -194 -113 -166 -85
rect -147 -113 -119 -85
rect -241 -160 -213 -132
rect -194 -160 -166 -132
rect -147 -160 -119 -132
rect 17660 -103 17692 -71
rect 17704 -103 17736 -71
rect 17748 -103 17780 -71
rect 17792 -103 17824 -71
rect 17660 -148 17692 -116
rect 17704 -148 17736 -116
rect 17748 -148 17780 -116
rect 17792 -148 17824 -116
rect -241 -207 -213 -179
rect -194 -207 -166 -179
rect -147 -207 -119 -179
rect 17898 -277 17930 -245
rect 17942 -277 17974 -245
rect 17986 -277 18018 -245
rect 18030 -277 18062 -245
rect 20442 -265 20561 -184
rect -1180 -342 -1148 -310
rect -1136 -342 -1104 -310
rect -1092 -342 -1060 -310
rect -1048 -342 -1016 -310
rect -1180 -387 -1148 -355
rect -1136 -387 -1104 -355
rect -1092 -387 -1060 -355
rect -1048 -387 -1016 -355
rect -1180 -432 -1148 -400
rect -1136 -432 -1104 -400
rect -1092 -432 -1060 -400
rect -1048 -432 -1016 -400
rect -430 -332 -402 -304
rect -383 -332 -355 -304
rect -336 -332 -308 -304
rect -430 -379 -402 -351
rect -383 -379 -355 -351
rect -336 -379 -308 -351
rect 17898 -322 17930 -290
rect 17942 -322 17974 -290
rect 17986 -322 18018 -290
rect 18030 -322 18062 -290
rect 17898 -367 17930 -335
rect 17942 -367 17974 -335
rect 17986 -367 18018 -335
rect 18030 -367 18062 -335
rect -430 -426 -402 -398
rect -383 -426 -355 -398
rect -336 -426 -308 -398
<< metal3 >>
rect 20151 11371 20567 11377
rect 20151 11290 20442 11371
rect 20561 11290 20567 11371
rect 20151 11285 20567 11290
rect 20435 11168 20567 11181
rect 20435 10962 20448 11168
rect 20554 10962 20567 11168
rect 20435 10950 20567 10962
rect 20151 10937 20319 10946
rect 20151 10862 20202 10937
rect 20308 10862 20319 10937
rect 20151 10855 20319 10862
rect 20151 10666 20319 10675
rect 20151 10591 20202 10666
rect 20308 10591 20319 10666
rect 20151 10584 20319 10591
rect 20151 10388 20319 10397
rect 20151 10313 20202 10388
rect 20308 10313 20319 10388
rect 20151 10306 20319 10313
rect 20435 10289 20567 10302
rect 20435 10083 20448 10289
rect 20554 10083 20567 10289
rect 20435 10071 20567 10083
rect 20151 9816 20567 9822
rect 20151 9735 20442 9816
rect 20561 9735 20567 9816
rect 20151 9730 20567 9735
rect 292 9595 438 9627
rect 292 9516 299 9595
rect 430 9516 438 9595
rect 292 9510 438 9516
rect 1856 9595 2002 9626
rect 1856 9516 1863 9595
rect 1994 9516 2002 9595
rect 1856 9510 2002 9516
rect 2292 9595 2438 9626
rect 2292 9516 2299 9595
rect 2430 9516 2438 9595
rect 2292 9510 2438 9516
rect 3856 9595 4002 9626
rect 3856 9516 3863 9595
rect 3994 9516 4002 9595
rect 3856 9510 4002 9516
rect 4292 9595 4438 9626
rect 4292 9516 4299 9595
rect 4430 9516 4438 9595
rect 4292 9510 4438 9516
rect 5856 9595 6002 9626
rect 5856 9516 5863 9595
rect 5994 9516 6002 9595
rect 5856 9510 6002 9516
rect 6292 9595 6438 9626
rect 6292 9516 6299 9595
rect 6430 9516 6438 9595
rect 6292 9510 6438 9516
rect 7856 9595 8002 9626
rect 7856 9516 7863 9595
rect 7994 9516 8002 9595
rect 7856 9510 8002 9516
rect 8292 9595 8438 9626
rect 8292 9516 8299 9595
rect 8430 9516 8438 9595
rect 8292 9510 8438 9516
rect 9856 9595 10002 9626
rect 9856 9516 9863 9595
rect 9994 9516 10002 9595
rect 9856 9510 10002 9516
rect 10292 9595 10438 9626
rect 10292 9516 10299 9595
rect 10430 9516 10438 9595
rect 10292 9510 10438 9516
rect 11856 9595 12002 9626
rect 11856 9516 11863 9595
rect 11994 9516 12002 9595
rect 11856 9510 12002 9516
rect 12292 9595 12438 9626
rect 12292 9516 12299 9595
rect 12430 9516 12438 9595
rect 12292 9510 12438 9516
rect 13856 9595 14002 9626
rect 13856 9516 13863 9595
rect 13994 9516 14002 9595
rect 13856 9510 14002 9516
rect 14292 9595 14438 9626
rect 14292 9516 14299 9595
rect 14430 9516 14438 9595
rect 14292 9510 14438 9516
rect 15856 9595 16002 9626
rect 15856 9516 15863 9595
rect 15994 9516 16002 9595
rect 15856 9510 16002 9516
rect 16292 9595 16438 9626
rect 16292 9516 16299 9595
rect 16430 9516 16438 9595
rect 17856 9595 18002 9626
rect 17856 9533 17863 9595
rect 17994 9533 18002 9595
rect 17856 9527 18002 9533
rect 16292 9510 16438 9516
rect -1195 9489 -988 9493
rect -1195 9457 -1180 9489
rect -1148 9457 -1136 9489
rect -1104 9457 -1092 9489
rect -1060 9457 -1048 9489
rect -1016 9457 -988 9489
rect -1195 9444 -988 9457
rect -1195 9412 -1180 9444
rect -1148 9412 -1136 9444
rect -1104 9412 -1092 9444
rect -1060 9412 -1048 9444
rect -1016 9412 -988 9444
rect -1195 9399 -988 9412
rect -1195 9367 -1180 9399
rect -1148 9367 -1136 9399
rect -1104 9367 -1092 9399
rect -1060 9367 -1048 9399
rect -1016 9367 -988 9399
rect -1195 9353 -988 9367
rect 1060 9484 1245 9493
rect 1060 9362 1072 9484
rect 1235 9362 1245 9484
rect 1060 9353 1245 9362
rect 3060 9484 3245 9493
rect 3060 9362 3072 9484
rect 3235 9362 3245 9484
rect 3060 9353 3245 9362
rect 5060 9484 5245 9493
rect 5060 9362 5072 9484
rect 5235 9362 5245 9484
rect 5060 9353 5245 9362
rect 7060 9484 7245 9493
rect 7060 9362 7072 9484
rect 7235 9362 7245 9484
rect 7060 9353 7245 9362
rect 9060 9484 9245 9493
rect 9060 9362 9072 9484
rect 9235 9362 9245 9484
rect 9060 9353 9245 9362
rect 11060 9484 11245 9493
rect 11060 9362 11072 9484
rect 11235 9362 11245 9484
rect 11060 9353 11245 9362
rect 13060 9484 13245 9493
rect 13060 9362 13072 9484
rect 13235 9362 13245 9484
rect 13060 9353 13245 9362
rect 15060 9484 15245 9493
rect 15060 9362 15072 9484
rect 15235 9362 15245 9484
rect 15060 9353 15245 9362
rect 17060 9484 17245 9493
rect 17060 9362 17072 9484
rect 17235 9362 17245 9484
rect 17060 9353 17245 9362
rect 17870 9489 18077 9493
rect 17870 9457 17898 9489
rect 17930 9457 17942 9489
rect 17974 9457 17986 9489
rect 18018 9457 18030 9489
rect 18062 9457 18077 9489
rect 17870 9444 18077 9457
rect 17870 9412 17898 9444
rect 17930 9412 17942 9444
rect 17974 9412 17986 9444
rect 18018 9412 18030 9444
rect 18062 9412 18077 9444
rect 17870 9399 18077 9412
rect 17870 9367 17898 9399
rect 17930 9367 17942 9399
rect 17974 9367 17986 9399
rect 18018 9367 18030 9399
rect 18062 9367 18077 9399
rect 17870 9353 18077 9367
rect 20151 9371 20567 9377
rect 20151 9290 20442 9371
rect 20561 9290 20567 9371
rect 20151 9285 20567 9290
rect -957 9270 -750 9274
rect -957 9238 -942 9270
rect -910 9238 -898 9270
rect -866 9238 -854 9270
rect -822 9238 -810 9270
rect -778 9238 -750 9270
rect -957 9225 -750 9238
rect -957 9193 -942 9225
rect -910 9193 -898 9225
rect -866 9193 -854 9225
rect -822 9193 -810 9225
rect -778 9193 -750 9225
rect -957 9180 -750 9193
rect -957 9148 -942 9180
rect -910 9148 -898 9180
rect -866 9148 -854 9180
rect -822 9148 -810 9180
rect -778 9148 -750 9180
rect -957 9134 -750 9148
rect 17632 9270 17839 9274
rect 17632 9238 17660 9270
rect 17692 9238 17704 9270
rect 17736 9238 17748 9270
rect 17780 9238 17792 9270
rect 17824 9238 17839 9270
rect 17632 9225 17839 9238
rect 17632 9193 17660 9225
rect 17692 9193 17704 9225
rect 17736 9193 17748 9225
rect 17780 9193 17792 9225
rect 17824 9193 17839 9225
rect 17632 9180 17839 9193
rect 17632 9148 17660 9180
rect 17692 9148 17704 9180
rect 17736 9148 17748 9180
rect 17780 9148 17792 9180
rect 17824 9148 17839 9180
rect 17632 9134 17839 9148
rect 20435 9168 20567 9181
rect 20435 8962 20448 9168
rect 20554 8962 20567 9168
rect 20435 8950 20567 8962
rect 20151 8937 20319 8946
rect -949 8877 -762 8878
rect -949 8845 -943 8877
rect -768 8845 -762 8877
rect 17644 8877 17831 8878
rect 17644 8873 17650 8877
rect -949 8844 -762 8845
rect 17633 8845 17650 8873
rect 17825 8873 17831 8877
rect 17633 8827 17661 8845
rect 17693 8827 17705 8845
rect 17737 8827 17749 8845
rect 17781 8827 17793 8845
rect 17825 8827 17840 8873
rect 20151 8862 20202 8937
rect 20308 8862 20319 8937
rect 20151 8855 20319 8862
rect 17633 8814 17840 8827
rect 17633 8782 17661 8814
rect 17693 8782 17705 8814
rect 17737 8782 17749 8814
rect 17781 8782 17793 8814
rect 17825 8782 17840 8814
rect 17633 8769 17840 8782
rect 17633 8737 17661 8769
rect 17693 8737 17705 8769
rect 17737 8737 17749 8769
rect 17781 8737 17793 8769
rect 17825 8737 17840 8769
rect 17633 8733 17840 8737
rect 20151 8666 20319 8675
rect 20151 8591 20202 8666
rect 20308 8591 20319 8666
rect 20151 8584 20319 8591
rect -949 8437 -762 8438
rect -949 8405 -943 8437
rect -768 8405 -762 8437
rect -949 8404 -762 8405
rect 17644 8437 17831 8438
rect 17644 8405 17650 8437
rect 17825 8405 17831 8437
rect 17644 8404 17831 8405
rect 20151 8388 20319 8397
rect 17870 8366 18077 8380
rect 17870 8334 17898 8366
rect 17930 8334 17942 8366
rect 17974 8334 17986 8366
rect 18018 8334 18030 8366
rect 18062 8334 18077 8366
rect 17870 8321 18077 8334
rect 17870 8289 17898 8321
rect 17930 8289 17942 8321
rect 17974 8289 17986 8321
rect 18018 8289 18030 8321
rect 18062 8289 18077 8321
rect 20151 8313 20202 8388
rect 20308 8313 20319 8388
rect 20151 8306 20319 8313
rect 17870 8276 18077 8289
rect 17870 8244 17898 8276
rect 17930 8244 17942 8276
rect 17974 8244 17986 8276
rect 18018 8244 18030 8276
rect 18062 8244 18077 8276
rect 17870 8240 18077 8244
rect 20435 8289 20567 8302
rect 20435 8083 20448 8289
rect 20554 8083 20567 8289
rect 20435 8071 20567 8083
rect -949 7997 -762 7998
rect -949 7965 -943 7997
rect -768 7965 -762 7997
rect -949 7964 -762 7965
rect 17644 7997 17831 7998
rect 17644 7965 17650 7997
rect 17825 7965 17831 7997
rect 17644 7964 17831 7965
rect 17632 7851 18151 7865
rect 17632 7819 17660 7851
rect 17692 7819 17704 7851
rect 17736 7819 17748 7851
rect 17780 7819 17792 7851
rect 17824 7819 18151 7851
rect 17632 7806 18151 7819
rect 17632 7774 17660 7806
rect 17692 7774 17704 7806
rect 17736 7774 17748 7806
rect 17780 7774 17792 7806
rect 17824 7774 18151 7806
rect 17632 7761 18151 7774
rect 17632 7729 17660 7761
rect 17692 7729 17704 7761
rect 17736 7729 17748 7761
rect 17780 7729 17792 7761
rect 17824 7729 18151 7761
rect 20151 7816 20567 7822
rect 20151 7735 20442 7816
rect 20561 7735 20567 7816
rect 20151 7730 20567 7735
rect 17632 7726 18151 7729
rect 17632 7725 17839 7726
rect -949 7557 -762 7558
rect -949 7525 -943 7557
rect -768 7525 -762 7557
rect -949 7524 -762 7525
rect 17644 7557 17831 7558
rect 17644 7525 17650 7557
rect 17825 7525 17831 7557
rect 17644 7524 17831 7525
rect 20151 7371 20567 7377
rect 17870 7312 18077 7326
rect 17870 7280 17898 7312
rect 17930 7280 17942 7312
rect 17974 7280 17986 7312
rect 18018 7280 18030 7312
rect 18062 7280 18077 7312
rect 20151 7290 20442 7371
rect 20561 7290 20567 7371
rect 20151 7285 20567 7290
rect 17870 7267 18077 7280
rect 17870 7235 17898 7267
rect 17930 7235 17942 7267
rect 17974 7235 17986 7267
rect 18018 7235 18030 7267
rect 18062 7235 18077 7267
rect 17870 7222 18077 7235
rect 17870 7190 17898 7222
rect 17930 7190 17942 7222
rect 17974 7190 17986 7222
rect 18018 7190 18030 7222
rect 18062 7190 18077 7222
rect 17870 7186 18077 7190
rect 20435 7168 20567 7181
rect -949 7117 -762 7118
rect -949 7085 -943 7117
rect -768 7085 -762 7117
rect -949 7084 -762 7085
rect 17644 7117 17831 7118
rect 17644 7085 17650 7117
rect 17825 7085 17831 7117
rect 17644 7084 17831 7085
rect 20435 6962 20448 7168
rect 20554 6962 20567 7168
rect 20435 6950 20567 6962
rect 20151 6937 20319 6946
rect 17632 6851 17839 6865
rect 20151 6862 20202 6937
rect 20308 6862 20319 6937
rect 20151 6855 20319 6862
rect 17632 6819 17660 6851
rect 17692 6819 17704 6851
rect 17736 6819 17748 6851
rect 17780 6819 17792 6851
rect 17824 6819 17839 6851
rect 17632 6806 17839 6819
rect 17632 6774 17660 6806
rect 17692 6774 17704 6806
rect 17736 6774 17748 6806
rect 17780 6774 17792 6806
rect 17824 6774 17839 6806
rect 17632 6761 17839 6774
rect 17632 6729 17660 6761
rect 17692 6729 17704 6761
rect 17736 6729 17748 6761
rect 17780 6729 17792 6761
rect 17824 6729 17839 6761
rect 17632 6726 17839 6729
rect -949 6677 -762 6678
rect -949 6645 -943 6677
rect -768 6645 -762 6677
rect -949 6644 -762 6645
rect 17644 6677 17831 6678
rect 17644 6645 17650 6677
rect 17825 6645 17831 6677
rect 17644 6644 17831 6645
rect 20151 6666 20319 6675
rect 20151 6591 20202 6666
rect 20308 6591 20319 6666
rect 20151 6584 20319 6591
rect 20151 6388 20319 6397
rect 17869 6347 18076 6361
rect 17869 6315 17897 6347
rect 17929 6315 17941 6347
rect 17973 6315 17985 6347
rect 18017 6315 18029 6347
rect 18061 6315 18076 6347
rect 17869 6302 18076 6315
rect 20151 6313 20202 6388
rect 20308 6313 20319 6388
rect 20151 6306 20319 6313
rect 17869 6270 17897 6302
rect 17929 6270 17941 6302
rect 17973 6270 17985 6302
rect 18017 6270 18029 6302
rect 18061 6270 18076 6302
rect 17869 6257 18076 6270
rect -949 6237 -762 6238
rect -949 6205 -943 6237
rect -768 6205 -762 6237
rect 17869 6225 17897 6257
rect 17929 6225 17941 6257
rect 17973 6225 17985 6257
rect 18017 6225 18029 6257
rect 18061 6225 18076 6257
rect 17869 6221 18076 6225
rect 20435 6289 20567 6302
rect -949 6204 -762 6205
rect 20435 6083 20448 6289
rect 20554 6083 20567 6289
rect 20435 6071 20567 6083
rect 17633 5902 17840 5903
rect 17633 5889 18151 5902
rect 17633 5857 17661 5889
rect 17693 5857 17705 5889
rect 17737 5857 17749 5889
rect 17781 5857 17793 5889
rect 17825 5857 18151 5889
rect 17633 5844 18151 5857
rect 17633 5812 17661 5844
rect 17693 5812 17705 5844
rect 17737 5812 17749 5844
rect 17781 5812 17793 5844
rect 17825 5812 18151 5844
rect 17633 5799 18151 5812
rect -949 5797 -762 5798
rect -949 5765 -943 5797
rect -768 5765 -762 5797
rect -949 5764 -762 5765
rect 17633 5797 17661 5799
rect 17633 5765 17650 5797
rect 17693 5797 17705 5799
rect 17737 5797 17749 5799
rect 17781 5797 17793 5799
rect 17825 5765 18151 5799
rect 17633 5763 18151 5765
rect 20151 5816 20567 5822
rect 20151 5735 20442 5816
rect 20561 5735 20567 5816
rect 20151 5730 20567 5735
rect 20151 5371 20567 5377
rect -949 5357 -762 5358
rect -949 5325 -943 5357
rect -768 5325 -762 5357
rect -949 5324 -762 5325
rect 17870 5339 18077 5353
rect 17870 5307 17898 5339
rect 17930 5307 17942 5339
rect 17974 5307 17986 5339
rect 18018 5307 18030 5339
rect 18062 5307 18077 5339
rect 17870 5294 18077 5307
rect 17870 5262 17898 5294
rect 17930 5262 17942 5294
rect 17974 5262 17986 5294
rect 18018 5262 18030 5294
rect 18062 5262 18077 5294
rect 20151 5290 20442 5371
rect 20561 5290 20567 5371
rect 20151 5285 20567 5290
rect 17870 5249 18077 5262
rect 17870 5217 17898 5249
rect 17930 5217 17942 5249
rect 17974 5217 17986 5249
rect 18018 5217 18030 5249
rect 18062 5217 18077 5249
rect 17870 5213 18077 5217
rect 20435 5168 20567 5181
rect 20435 4962 20448 5168
rect 20554 4962 20567 5168
rect 20435 4950 20567 4962
rect 20151 4937 20319 4946
rect -949 4917 -762 4918
rect -949 4885 -943 4917
rect -768 4885 -762 4917
rect -949 4884 -762 4885
rect 17644 4917 17831 4918
rect 17644 4885 17650 4917
rect 17825 4885 17831 4917
rect 17644 4884 17831 4885
rect 20151 4862 20202 4937
rect 20308 4862 20319 4937
rect 20151 4855 20319 4862
rect 17632 4826 17839 4840
rect 17632 4794 17660 4826
rect 17692 4794 17704 4826
rect 17736 4794 17748 4826
rect 17780 4794 17792 4826
rect 17824 4794 17839 4826
rect 17632 4781 17839 4794
rect 17632 4749 17660 4781
rect 17692 4749 17704 4781
rect 17736 4749 17748 4781
rect 17780 4749 17792 4781
rect 17824 4749 17839 4781
rect 17632 4736 17839 4749
rect 17632 4704 17660 4736
rect 17692 4704 17704 4736
rect 17736 4704 17748 4736
rect 17780 4704 17792 4736
rect 17824 4704 17839 4736
rect 17632 4700 17839 4704
rect 20151 4666 20319 4675
rect 20151 4591 20202 4666
rect 20308 4591 20319 4666
rect 20151 4584 20319 4591
rect -949 4477 -762 4478
rect -949 4445 -943 4477
rect -768 4445 -762 4477
rect -949 4444 -762 4445
rect 17644 4477 17831 4478
rect 17644 4445 17650 4477
rect 17825 4445 17831 4477
rect 17644 4444 17831 4445
rect 20151 4388 20319 4397
rect 17870 4338 18077 4352
rect 17870 4306 17898 4338
rect 17930 4306 17942 4338
rect 17974 4306 17986 4338
rect 18018 4306 18030 4338
rect 18062 4306 18077 4338
rect 20151 4313 20202 4388
rect 20308 4313 20319 4388
rect 20151 4306 20319 4313
rect 17870 4293 18077 4306
rect 17870 4261 17898 4293
rect 17930 4261 17942 4293
rect 17974 4261 17986 4293
rect 18018 4261 18030 4293
rect 18062 4261 18077 4293
rect 17870 4248 18077 4261
rect 17870 4216 17898 4248
rect 17930 4216 17942 4248
rect 17974 4216 17986 4248
rect 18018 4216 18030 4248
rect 18062 4216 18077 4248
rect 17870 4212 18077 4216
rect 20435 4289 20567 4302
rect 20435 4083 20448 4289
rect 20554 4083 20567 4289
rect 20435 4071 20567 4083
rect -949 4037 -762 4038
rect -949 4005 -943 4037
rect -768 4005 -762 4037
rect -949 4004 -762 4005
rect 17644 4037 17831 4038
rect 17644 4005 17650 4037
rect 17825 4005 17831 4037
rect 17644 4004 17831 4005
rect 17633 3851 17840 3852
rect 17633 3838 18151 3851
rect 17633 3806 17661 3838
rect 17693 3806 17705 3838
rect 17737 3806 17749 3838
rect 17781 3806 17793 3838
rect 17825 3806 18151 3838
rect 17633 3793 18151 3806
rect 17633 3761 17661 3793
rect 17693 3761 17705 3793
rect 17737 3761 17749 3793
rect 17781 3761 17793 3793
rect 17825 3761 18151 3793
rect 17633 3748 18151 3761
rect 17633 3716 17661 3748
rect 17693 3716 17705 3748
rect 17737 3716 17749 3748
rect 17781 3716 17793 3748
rect 17825 3716 18151 3748
rect 20151 3816 20567 3822
rect 20151 3735 20442 3816
rect 20561 3735 20567 3816
rect 20151 3730 20567 3735
rect 17633 3712 18151 3716
rect -949 3597 -762 3598
rect -949 3565 -943 3597
rect -768 3565 -762 3597
rect -949 3564 -762 3565
rect 17644 3597 17831 3598
rect 17644 3565 17650 3597
rect 17825 3565 17831 3597
rect 17644 3564 17831 3565
rect 20151 3371 20567 3377
rect 17869 3339 18076 3353
rect 17869 3307 17897 3339
rect 17929 3307 17941 3339
rect 17973 3307 17985 3339
rect 18017 3307 18029 3339
rect 18061 3307 18076 3339
rect 17869 3294 18076 3307
rect 17869 3262 17897 3294
rect 17929 3262 17941 3294
rect 17973 3262 17985 3294
rect 18017 3262 18029 3294
rect 18061 3262 18076 3294
rect 20151 3290 20442 3371
rect 20561 3290 20567 3371
rect 20151 3285 20567 3290
rect 17869 3249 18076 3262
rect 17869 3217 17897 3249
rect 17929 3217 17941 3249
rect 17973 3217 17985 3249
rect 18017 3217 18029 3249
rect 18061 3217 18076 3249
rect 17869 3213 18076 3217
rect 20435 3168 20567 3181
rect -949 3157 -762 3158
rect -949 3125 -943 3157
rect -768 3125 -762 3157
rect -949 3124 -762 3125
rect 17644 3157 17831 3158
rect 17644 3125 17650 3157
rect 17825 3125 17831 3157
rect 17644 3124 17831 3125
rect 20435 2962 20448 3168
rect 20554 2962 20567 3168
rect 20435 2950 20567 2962
rect 20151 2937 20319 2946
rect 20151 2862 20202 2937
rect 20308 2862 20319 2937
rect 20151 2855 20319 2862
rect 17633 2816 17840 2830
rect 17633 2784 17661 2816
rect 17693 2784 17705 2816
rect 17737 2784 17749 2816
rect 17781 2784 17793 2816
rect 17825 2784 17840 2816
rect 17633 2771 17840 2784
rect 17633 2739 17661 2771
rect 17693 2739 17705 2771
rect 17737 2739 17749 2771
rect 17781 2739 17793 2771
rect 17825 2739 17840 2771
rect 17633 2726 17840 2739
rect -949 2717 -762 2718
rect -949 2685 -943 2717
rect -768 2685 -762 2717
rect 17633 2717 17661 2726
rect 17633 2690 17650 2717
rect 17693 2717 17705 2726
rect 17737 2717 17749 2726
rect 17781 2717 17793 2726
rect -949 2684 -762 2685
rect 17644 2685 17650 2690
rect 17825 2690 17840 2726
rect 17825 2685 17831 2690
rect 17644 2684 17831 2685
rect 20151 2666 20319 2675
rect 20151 2591 20202 2666
rect 20308 2591 20319 2666
rect 20151 2584 20319 2591
rect 20151 2388 20319 2397
rect 17870 2305 18077 2319
rect 20151 2313 20202 2388
rect 20308 2313 20319 2388
rect 20151 2306 20319 2313
rect -949 2277 -762 2278
rect -949 2245 -943 2277
rect -768 2245 -762 2277
rect -949 2244 -762 2245
rect 17870 2273 17898 2305
rect 17930 2273 17942 2305
rect 17974 2273 17986 2305
rect 18018 2273 18030 2305
rect 18062 2273 18077 2305
rect 17870 2260 18077 2273
rect 17870 2228 17898 2260
rect 17930 2228 17942 2260
rect 17974 2228 17986 2260
rect 18018 2228 18030 2260
rect 18062 2228 18077 2260
rect 17870 2215 18077 2228
rect 17870 2183 17898 2215
rect 17930 2183 17942 2215
rect 17974 2183 17986 2215
rect 18018 2183 18030 2215
rect 18062 2183 18077 2215
rect 17870 2179 18077 2183
rect 20435 2289 20567 2302
rect 20435 2083 20448 2289
rect 20554 2083 20567 2289
rect 20435 2071 20567 2083
rect -949 1837 -762 1838
rect -949 1805 -943 1837
rect -768 1805 -762 1837
rect 17644 1837 17831 1838
rect 17644 1833 17650 1837
rect -949 1804 -762 1805
rect 17633 1805 17650 1833
rect 17825 1833 17831 1837
rect 17633 1787 17661 1805
rect 17693 1787 17705 1805
rect 17737 1787 17749 1805
rect 17781 1787 17793 1805
rect 17825 1787 18151 1833
rect 17633 1774 18151 1787
rect 17633 1742 17661 1774
rect 17693 1742 17705 1774
rect 17737 1742 17749 1774
rect 17781 1742 17793 1774
rect 17825 1742 18151 1774
rect 17633 1729 18151 1742
rect 20151 1816 20567 1822
rect 20151 1735 20442 1816
rect 20561 1735 20567 1816
rect 20151 1730 20567 1735
rect 17633 1697 17661 1729
rect 17693 1697 17705 1729
rect 17737 1697 17749 1729
rect 17781 1697 17793 1729
rect 17825 1697 18151 1729
rect 17633 1694 18151 1697
rect 17633 1693 17839 1694
rect -949 1397 -762 1398
rect -949 1365 -943 1397
rect -768 1365 -762 1397
rect -949 1364 -762 1365
rect 17644 1397 17831 1398
rect 17644 1365 17650 1397
rect 17825 1365 17831 1397
rect 17644 1364 17831 1365
rect 20151 1371 20567 1377
rect 17870 1303 18077 1317
rect 17870 1271 17898 1303
rect 17930 1271 17942 1303
rect 17974 1271 17986 1303
rect 18018 1271 18030 1303
rect 18062 1271 18077 1303
rect 20151 1290 20442 1371
rect 20561 1290 20567 1371
rect 20151 1285 20567 1290
rect 17870 1258 18077 1271
rect 17870 1226 17898 1258
rect 17930 1226 17942 1258
rect 17974 1226 17986 1258
rect 18018 1226 18030 1258
rect 18062 1226 18077 1258
rect 17870 1213 18077 1226
rect 17870 1181 17898 1213
rect 17930 1181 17942 1213
rect 17974 1181 17986 1213
rect 18018 1181 18030 1213
rect 18062 1181 18077 1213
rect 17870 1177 18077 1181
rect 20435 1168 20567 1181
rect 20435 962 20448 1168
rect 20554 962 20567 1168
rect -949 957 -762 958
rect -949 925 -943 957
rect -768 925 -762 957
rect -949 924 -762 925
rect 17644 957 17831 958
rect 17644 925 17650 957
rect 17825 925 17831 957
rect 20435 950 20567 962
rect 17644 924 17831 925
rect 20151 937 20319 946
rect 20151 862 20202 937
rect 20308 862 20319 937
rect 20151 855 20319 862
rect 17631 819 17838 833
rect 17631 787 17659 819
rect 17691 787 17703 819
rect 17735 787 17747 819
rect 17779 787 17791 819
rect 17823 787 17838 819
rect 17631 774 17838 787
rect 17631 742 17659 774
rect 17691 742 17703 774
rect 17735 742 17747 774
rect 17779 742 17791 774
rect 17823 742 17838 774
rect 17631 729 17838 742
rect 17631 697 17659 729
rect 17691 697 17703 729
rect 17735 697 17747 729
rect 17779 697 17791 729
rect 17823 697 17838 729
rect 17631 693 17838 697
rect 20151 666 20319 675
rect 20151 591 20202 666
rect 20308 591 20319 666
rect 20151 584 20319 591
rect -949 517 -762 518
rect -949 485 -943 517
rect -768 485 -762 517
rect -949 484 -762 485
rect 17644 517 17831 518
rect 17644 485 17650 517
rect 17825 485 17831 517
rect 17644 484 17831 485
rect 20151 388 20319 397
rect 17870 306 18077 320
rect 20151 313 20202 388
rect 20308 313 20319 388
rect 20151 306 20319 313
rect 17870 274 17898 306
rect 17930 274 17942 306
rect 17974 274 17986 306
rect 18018 274 18030 306
rect 18062 274 18077 306
rect 17870 261 18077 274
rect 17870 229 17898 261
rect 17930 229 17942 261
rect 17974 229 17986 261
rect 18018 229 18030 261
rect 18062 229 18077 261
rect 17870 216 18077 229
rect 17870 184 17898 216
rect 17930 184 17942 216
rect 17974 184 17986 216
rect 18018 184 18030 216
rect 18062 184 18077 216
rect 17870 180 18077 184
rect 20435 289 20567 302
rect 20435 83 20448 289
rect 20554 83 20567 289
rect -949 77 -762 78
rect -949 45 -943 77
rect -768 45 -762 77
rect -949 44 -762 45
rect 17644 77 17831 78
rect 17644 45 17650 77
rect 17825 45 17831 77
rect 20435 71 20567 83
rect 17644 44 17831 45
rect 17632 -13 17839 -12
rect 17632 -26 18151 -13
rect 17632 -58 17660 -26
rect 17692 -58 17704 -26
rect 17736 -58 17748 -26
rect 17780 -58 17792 -26
rect 17824 -58 18151 -26
rect 17632 -71 18151 -58
rect -958 -85 -91 -76
rect -958 -91 -241 -85
rect -958 -123 -942 -91
rect -910 -123 -898 -91
rect -866 -123 -854 -91
rect -822 -123 -810 -91
rect -778 -113 -241 -91
rect -213 -113 -194 -85
rect -166 -113 -147 -85
rect -119 -113 -91 -85
rect -778 -123 -91 -113
rect -958 -132 -91 -123
rect -958 -136 -241 -132
rect -958 -168 -942 -136
rect -910 -168 -898 -136
rect -866 -168 -854 -136
rect -822 -168 -810 -136
rect -778 -160 -241 -136
rect -213 -160 -194 -132
rect -166 -160 -147 -132
rect -119 -160 -91 -132
rect 17632 -103 17660 -71
rect 17692 -103 17704 -71
rect 17736 -103 17748 -71
rect 17780 -103 17792 -71
rect 17824 -103 18151 -71
rect 17632 -116 18151 -103
rect 17632 -148 17660 -116
rect 17692 -148 17704 -116
rect 17736 -148 17748 -116
rect 17780 -148 17792 -116
rect 17824 -148 18151 -116
rect 17632 -152 18151 -148
rect -778 -168 -91 -160
rect -958 -179 -91 -168
rect -958 -181 -241 -179
rect -958 -213 -942 -181
rect -910 -213 -898 -181
rect -866 -213 -854 -181
rect -822 -213 -810 -181
rect -778 -207 -241 -181
rect -213 -207 -194 -179
rect -166 -207 -147 -179
rect -119 -207 -91 -179
rect -778 -213 -91 -207
rect -958 -217 -91 -213
rect 20151 -184 20567 -178
rect 17870 -245 18077 -231
rect 17870 -277 17898 -245
rect 17930 -277 17942 -245
rect 17974 -277 17986 -245
rect 18018 -277 18030 -245
rect 18062 -277 18077 -245
rect 20151 -265 20442 -184
rect 20561 -265 20567 -184
rect 20151 -270 20567 -265
rect 17870 -290 18077 -277
rect -988 -296 -280 -295
rect -1195 -304 -280 -296
rect -1195 -310 -430 -304
rect -1195 -342 -1180 -310
rect -1148 -342 -1136 -310
rect -1104 -342 -1092 -310
rect -1060 -342 -1048 -310
rect -1016 -332 -430 -310
rect -402 -332 -383 -304
rect -355 -332 -336 -304
rect -308 -332 -280 -304
rect -1016 -342 -280 -332
rect -1195 -351 -280 -342
rect -1195 -355 -430 -351
rect -1195 -387 -1180 -355
rect -1148 -387 -1136 -355
rect -1104 -387 -1092 -355
rect -1060 -387 -1048 -355
rect -1016 -379 -430 -355
rect -402 -379 -383 -351
rect -355 -379 -336 -351
rect -308 -379 -280 -351
rect 17870 -322 17898 -290
rect 17930 -322 17942 -290
rect 17974 -322 17986 -290
rect 18018 -322 18030 -290
rect 18062 -322 18077 -290
rect 17870 -335 18077 -322
rect 17870 -367 17898 -335
rect 17930 -367 17942 -335
rect 17974 -367 17986 -335
rect 18018 -367 18030 -335
rect 18062 -367 18077 -335
rect 17870 -371 18077 -367
rect -1016 -387 -280 -379
rect -1195 -398 -280 -387
rect -1195 -400 -430 -398
rect -1195 -432 -1180 -400
rect -1148 -432 -1136 -400
rect -1104 -432 -1092 -400
rect -1060 -432 -1048 -400
rect -1016 -426 -430 -400
rect -402 -426 -383 -398
rect -355 -426 -336 -398
rect -308 -426 -280 -398
rect -1016 -432 -280 -426
rect -1195 -436 -280 -432
<< via3 >>
rect 20442 11290 20561 11371
rect 20448 10962 20554 11168
rect 20202 10862 20308 10937
rect 20202 10591 20308 10666
rect 20202 10313 20308 10388
rect 20448 10083 20554 10289
rect 20442 9735 20561 9816
rect -1180 9457 -1148 9489
rect -1136 9457 -1104 9489
rect -1092 9457 -1060 9489
rect -1048 9457 -1016 9489
rect -1180 9412 -1148 9444
rect -1136 9412 -1104 9444
rect -1092 9412 -1060 9444
rect -1048 9412 -1016 9444
rect -1180 9367 -1148 9399
rect -1136 9367 -1104 9399
rect -1092 9367 -1060 9399
rect -1048 9367 -1016 9399
rect 1072 9362 1235 9484
rect 3072 9362 3235 9484
rect 5072 9362 5235 9484
rect 7072 9362 7235 9484
rect 9072 9362 9235 9484
rect 11072 9362 11235 9484
rect 13072 9362 13235 9484
rect 15072 9362 15235 9484
rect 17072 9362 17235 9484
rect 17898 9457 17930 9489
rect 17942 9457 17974 9489
rect 17986 9457 18018 9489
rect 18030 9457 18062 9489
rect 17898 9412 17930 9444
rect 17942 9412 17974 9444
rect 17986 9412 18018 9444
rect 18030 9412 18062 9444
rect 17898 9367 17930 9399
rect 17942 9367 17974 9399
rect 17986 9367 18018 9399
rect 18030 9367 18062 9399
rect 20442 9290 20561 9371
rect -942 9238 -910 9270
rect -898 9238 -866 9270
rect -854 9238 -822 9270
rect -810 9238 -778 9270
rect -942 9193 -910 9225
rect -898 9193 -866 9225
rect -854 9193 -822 9225
rect -810 9193 -778 9225
rect -942 9148 -910 9180
rect -898 9148 -866 9180
rect -854 9148 -822 9180
rect -810 9148 -778 9180
rect 17660 9238 17692 9270
rect 17704 9238 17736 9270
rect 17748 9238 17780 9270
rect 17792 9238 17824 9270
rect 17660 9193 17692 9225
rect 17704 9193 17736 9225
rect 17748 9193 17780 9225
rect 17792 9193 17824 9225
rect 17660 9148 17692 9180
rect 17704 9148 17736 9180
rect 17748 9148 17780 9180
rect 17792 9148 17824 9180
rect 20448 8962 20554 9168
rect -943 8875 -768 8877
rect -943 8847 -768 8875
rect -943 8845 -768 8847
rect 17650 8875 17825 8877
rect 17650 8847 17825 8875
rect 17650 8845 17661 8847
rect 17661 8827 17693 8847
rect 17693 8845 17705 8847
rect 17705 8827 17737 8847
rect 17737 8845 17749 8847
rect 17749 8827 17781 8847
rect 17781 8845 17793 8847
rect 17793 8827 17825 8847
rect 20202 8862 20308 8937
rect 17661 8782 17693 8814
rect 17705 8782 17737 8814
rect 17749 8782 17781 8814
rect 17793 8782 17825 8814
rect 17661 8737 17693 8769
rect 17705 8737 17737 8769
rect 17749 8737 17781 8769
rect 17793 8737 17825 8769
rect 20202 8591 20308 8666
rect -943 8435 -768 8437
rect -943 8407 -768 8435
rect -943 8405 -768 8407
rect 17650 8435 17825 8437
rect 17650 8407 17825 8435
rect 17650 8405 17825 8407
rect 17898 8334 17930 8366
rect 17942 8334 17974 8366
rect 17986 8334 18018 8366
rect 18030 8334 18062 8366
rect 17898 8289 17930 8321
rect 17942 8289 17974 8321
rect 17986 8289 18018 8321
rect 18030 8289 18062 8321
rect 20202 8313 20308 8388
rect 17898 8244 17930 8276
rect 17942 8244 17974 8276
rect 17986 8244 18018 8276
rect 18030 8244 18062 8276
rect 20448 8083 20554 8289
rect -943 7995 -768 7997
rect -943 7967 -768 7995
rect -943 7965 -768 7967
rect 17650 7995 17825 7997
rect 17650 7967 17825 7995
rect 17650 7965 17825 7967
rect 17660 7819 17692 7851
rect 17704 7819 17736 7851
rect 17748 7819 17780 7851
rect 17792 7819 17824 7851
rect 17660 7774 17692 7806
rect 17704 7774 17736 7806
rect 17748 7774 17780 7806
rect 17792 7774 17824 7806
rect 17660 7729 17692 7761
rect 17704 7729 17736 7761
rect 17748 7729 17780 7761
rect 17792 7729 17824 7761
rect 20442 7735 20561 7816
rect -943 7555 -768 7557
rect -943 7527 -768 7555
rect -943 7525 -768 7527
rect 17650 7555 17825 7557
rect 17650 7527 17825 7555
rect 17650 7525 17825 7527
rect 17898 7280 17930 7312
rect 17942 7280 17974 7312
rect 17986 7280 18018 7312
rect 18030 7280 18062 7312
rect 20442 7290 20561 7371
rect 17898 7235 17930 7267
rect 17942 7235 17974 7267
rect 17986 7235 18018 7267
rect 18030 7235 18062 7267
rect 17898 7190 17930 7222
rect 17942 7190 17974 7222
rect 17986 7190 18018 7222
rect 18030 7190 18062 7222
rect -943 7115 -768 7117
rect -943 7087 -768 7115
rect -943 7085 -768 7087
rect 17650 7115 17825 7117
rect 17650 7087 17825 7115
rect 17650 7085 17825 7087
rect 20448 6962 20554 7168
rect 20202 6862 20308 6937
rect 17660 6819 17692 6851
rect 17704 6819 17736 6851
rect 17748 6819 17780 6851
rect 17792 6819 17824 6851
rect 17660 6774 17692 6806
rect 17704 6774 17736 6806
rect 17748 6774 17780 6806
rect 17792 6774 17824 6806
rect 17660 6729 17692 6761
rect 17704 6729 17736 6761
rect 17748 6729 17780 6761
rect 17792 6729 17824 6761
rect -943 6675 -768 6677
rect -943 6647 -768 6675
rect -943 6645 -768 6647
rect 17650 6675 17825 6677
rect 17650 6647 17825 6675
rect 17650 6645 17825 6647
rect 20202 6591 20308 6666
rect 17897 6315 17929 6347
rect 17941 6315 17973 6347
rect 17985 6315 18017 6347
rect 18029 6315 18061 6347
rect 20202 6313 20308 6388
rect 17897 6270 17929 6302
rect 17941 6270 17973 6302
rect 17985 6270 18017 6302
rect 18029 6270 18061 6302
rect -943 6235 -768 6237
rect -943 6207 -768 6235
rect -943 6205 -768 6207
rect 17897 6225 17929 6257
rect 17941 6225 17973 6257
rect 17985 6225 18017 6257
rect 18029 6225 18061 6257
rect 20448 6083 20554 6289
rect 17661 5857 17693 5889
rect 17705 5857 17737 5889
rect 17749 5857 17781 5889
rect 17793 5857 17825 5889
rect 17661 5812 17693 5844
rect 17705 5812 17737 5844
rect 17749 5812 17781 5844
rect 17793 5812 17825 5844
rect -943 5795 -768 5797
rect -943 5767 -768 5795
rect -943 5765 -768 5767
rect 17650 5795 17661 5797
rect 17661 5795 17693 5799
rect 17693 5795 17705 5797
rect 17705 5795 17737 5799
rect 17737 5795 17749 5797
rect 17749 5795 17781 5799
rect 17781 5795 17793 5797
rect 17793 5795 17825 5799
rect 17650 5767 17825 5795
rect 17650 5765 17825 5767
rect 20442 5735 20561 5816
rect -943 5355 -768 5357
rect -943 5327 -768 5355
rect -943 5325 -768 5327
rect 17898 5307 17930 5339
rect 17942 5307 17974 5339
rect 17986 5307 18018 5339
rect 18030 5307 18062 5339
rect 17898 5262 17930 5294
rect 17942 5262 17974 5294
rect 17986 5262 18018 5294
rect 18030 5262 18062 5294
rect 20442 5290 20561 5371
rect 17898 5217 17930 5249
rect 17942 5217 17974 5249
rect 17986 5217 18018 5249
rect 18030 5217 18062 5249
rect 20448 4962 20554 5168
rect -943 4915 -768 4917
rect -943 4887 -768 4915
rect -943 4885 -768 4887
rect 17650 4915 17825 4917
rect 17650 4887 17825 4915
rect 17650 4885 17825 4887
rect 20202 4862 20308 4937
rect 17660 4794 17692 4826
rect 17704 4794 17736 4826
rect 17748 4794 17780 4826
rect 17792 4794 17824 4826
rect 17660 4749 17692 4781
rect 17704 4749 17736 4781
rect 17748 4749 17780 4781
rect 17792 4749 17824 4781
rect 17660 4704 17692 4736
rect 17704 4704 17736 4736
rect 17748 4704 17780 4736
rect 17792 4704 17824 4736
rect 20202 4591 20308 4666
rect -943 4475 -768 4477
rect -943 4447 -768 4475
rect -943 4445 -768 4447
rect 17650 4475 17825 4477
rect 17650 4447 17825 4475
rect 17650 4445 17825 4447
rect 17898 4306 17930 4338
rect 17942 4306 17974 4338
rect 17986 4306 18018 4338
rect 18030 4306 18062 4338
rect 20202 4313 20308 4388
rect 17898 4261 17930 4293
rect 17942 4261 17974 4293
rect 17986 4261 18018 4293
rect 18030 4261 18062 4293
rect 17898 4216 17930 4248
rect 17942 4216 17974 4248
rect 17986 4216 18018 4248
rect 18030 4216 18062 4248
rect 20448 4083 20554 4289
rect -943 4035 -768 4037
rect -943 4007 -768 4035
rect -943 4005 -768 4007
rect 17650 4035 17825 4037
rect 17650 4007 17825 4035
rect 17650 4005 17825 4007
rect 17661 3806 17693 3838
rect 17705 3806 17737 3838
rect 17749 3806 17781 3838
rect 17793 3806 17825 3838
rect 17661 3761 17693 3793
rect 17705 3761 17737 3793
rect 17749 3761 17781 3793
rect 17793 3761 17825 3793
rect 17661 3716 17693 3748
rect 17705 3716 17737 3748
rect 17749 3716 17781 3748
rect 17793 3716 17825 3748
rect 20442 3735 20561 3816
rect -943 3595 -768 3597
rect -943 3567 -768 3595
rect -943 3565 -768 3567
rect 17650 3595 17825 3597
rect 17650 3567 17825 3595
rect 17650 3565 17825 3567
rect 17897 3307 17929 3339
rect 17941 3307 17973 3339
rect 17985 3307 18017 3339
rect 18029 3307 18061 3339
rect 17897 3262 17929 3294
rect 17941 3262 17973 3294
rect 17985 3262 18017 3294
rect 18029 3262 18061 3294
rect 20442 3290 20561 3371
rect 17897 3217 17929 3249
rect 17941 3217 17973 3249
rect 17985 3217 18017 3249
rect 18029 3217 18061 3249
rect -943 3155 -768 3157
rect -943 3127 -768 3155
rect -943 3125 -768 3127
rect 17650 3155 17825 3157
rect 17650 3127 17825 3155
rect 17650 3125 17825 3127
rect 20448 2962 20554 3168
rect 20202 2862 20308 2937
rect 17661 2784 17693 2816
rect 17705 2784 17737 2816
rect 17749 2784 17781 2816
rect 17793 2784 17825 2816
rect 17661 2739 17693 2771
rect 17705 2739 17737 2771
rect 17749 2739 17781 2771
rect 17793 2739 17825 2771
rect -943 2715 -768 2717
rect -943 2687 -768 2715
rect -943 2685 -768 2687
rect 17650 2715 17661 2717
rect 17661 2715 17693 2726
rect 17693 2715 17705 2717
rect 17705 2715 17737 2726
rect 17737 2715 17749 2717
rect 17749 2715 17781 2726
rect 17781 2715 17793 2717
rect 17793 2715 17825 2726
rect 17650 2687 17825 2715
rect 17650 2685 17825 2687
rect 20202 2591 20308 2666
rect 20202 2313 20308 2388
rect -943 2275 -768 2277
rect -943 2247 -768 2275
rect -943 2245 -768 2247
rect 17898 2273 17930 2305
rect 17942 2273 17974 2305
rect 17986 2273 18018 2305
rect 18030 2273 18062 2305
rect 17898 2228 17930 2260
rect 17942 2228 17974 2260
rect 17986 2228 18018 2260
rect 18030 2228 18062 2260
rect 17898 2183 17930 2215
rect 17942 2183 17974 2215
rect 17986 2183 18018 2215
rect 18030 2183 18062 2215
rect 20448 2083 20554 2289
rect -943 1835 -768 1837
rect -943 1807 -768 1835
rect -943 1805 -768 1807
rect 17650 1835 17825 1837
rect 17650 1807 17825 1835
rect 17650 1805 17661 1807
rect 17661 1787 17693 1807
rect 17693 1805 17705 1807
rect 17705 1787 17737 1807
rect 17737 1805 17749 1807
rect 17749 1787 17781 1807
rect 17781 1805 17793 1807
rect 17793 1787 17825 1807
rect 17661 1742 17693 1774
rect 17705 1742 17737 1774
rect 17749 1742 17781 1774
rect 17793 1742 17825 1774
rect 20442 1735 20561 1816
rect 17661 1697 17693 1729
rect 17705 1697 17737 1729
rect 17749 1697 17781 1729
rect 17793 1697 17825 1729
rect -943 1395 -768 1397
rect -943 1367 -768 1395
rect -943 1365 -768 1367
rect 17650 1395 17825 1397
rect 17650 1367 17825 1395
rect 17650 1365 17825 1367
rect 17898 1271 17930 1303
rect 17942 1271 17974 1303
rect 17986 1271 18018 1303
rect 18030 1271 18062 1303
rect 20442 1290 20561 1371
rect 17898 1226 17930 1258
rect 17942 1226 17974 1258
rect 17986 1226 18018 1258
rect 18030 1226 18062 1258
rect 17898 1181 17930 1213
rect 17942 1181 17974 1213
rect 17986 1181 18018 1213
rect 18030 1181 18062 1213
rect 20448 962 20554 1168
rect -943 955 -768 957
rect -943 927 -768 955
rect -943 925 -768 927
rect 17650 955 17825 957
rect 17650 927 17825 955
rect 17650 925 17825 927
rect 20202 862 20308 937
rect 17659 787 17691 819
rect 17703 787 17735 819
rect 17747 787 17779 819
rect 17791 787 17823 819
rect 17659 742 17691 774
rect 17703 742 17735 774
rect 17747 742 17779 774
rect 17791 742 17823 774
rect 17659 697 17691 729
rect 17703 697 17735 729
rect 17747 697 17779 729
rect 17791 697 17823 729
rect 20202 591 20308 666
rect -943 515 -768 517
rect -943 487 -768 515
rect -943 485 -768 487
rect 17650 515 17825 517
rect 17650 487 17825 515
rect 17650 485 17825 487
rect 20202 313 20308 388
rect 17898 274 17930 306
rect 17942 274 17974 306
rect 17986 274 18018 306
rect 18030 274 18062 306
rect 17898 229 17930 261
rect 17942 229 17974 261
rect 17986 229 18018 261
rect 18030 229 18062 261
rect 17898 184 17930 216
rect 17942 184 17974 216
rect 17986 184 18018 216
rect 18030 184 18062 216
rect 20448 83 20554 289
rect -943 75 -768 77
rect -943 47 -768 75
rect -943 45 -768 47
rect 17650 75 17825 77
rect 17650 47 17825 75
rect 17650 45 17825 47
rect 17660 -58 17692 -26
rect 17704 -58 17736 -26
rect 17748 -58 17780 -26
rect 17792 -58 17824 -26
rect -942 -123 -910 -91
rect -898 -123 -866 -91
rect -854 -123 -822 -91
rect -810 -123 -778 -91
rect -942 -168 -910 -136
rect -898 -168 -866 -136
rect -854 -168 -822 -136
rect -810 -168 -778 -136
rect 17660 -103 17692 -71
rect 17704 -103 17736 -71
rect 17748 -103 17780 -71
rect 17792 -103 17824 -71
rect 17660 -148 17692 -116
rect 17704 -148 17736 -116
rect 17748 -148 17780 -116
rect 17792 -148 17824 -116
rect -942 -213 -910 -181
rect -898 -213 -866 -181
rect -854 -213 -822 -181
rect -810 -213 -778 -181
rect 17898 -277 17930 -245
rect 17942 -277 17974 -245
rect 17986 -277 18018 -245
rect 18030 -277 18062 -245
rect 20442 -265 20561 -184
rect -1180 -342 -1148 -310
rect -1136 -342 -1104 -310
rect -1092 -342 -1060 -310
rect -1048 -342 -1016 -310
rect -1180 -387 -1148 -355
rect -1136 -387 -1104 -355
rect -1092 -387 -1060 -355
rect -1048 -387 -1016 -355
rect 17898 -322 17930 -290
rect 17942 -322 17974 -290
rect 17986 -322 18018 -290
rect 18030 -322 18062 -290
rect 17898 -367 17930 -335
rect 17942 -367 17974 -335
rect 17986 -367 18018 -335
rect 18030 -367 18062 -335
rect -1180 -432 -1148 -400
rect -1136 -432 -1104 -400
rect -1092 -432 -1060 -400
rect -1048 -432 -1016 -400
<< metal4 >>
rect -1195 9489 -988 11626
rect -1195 9457 -1180 9489
rect -1148 9457 -1136 9489
rect -1104 9457 -1092 9489
rect -1060 9457 -1048 9489
rect -1016 9457 -988 9489
rect -1195 9444 -988 9457
rect -1195 9412 -1180 9444
rect -1148 9412 -1136 9444
rect -1104 9412 -1092 9444
rect -1060 9412 -1048 9444
rect -1016 9412 -988 9444
rect -1195 9399 -988 9412
rect -1195 9367 -1180 9399
rect -1148 9367 -1136 9399
rect -1104 9367 -1092 9399
rect -1060 9367 -1048 9399
rect -1016 9367 -988 9399
rect -1195 -310 -988 9367
rect -957 9270 -750 11626
rect 20191 10946 20398 11626
rect 20151 10937 20398 10946
rect 20151 10862 20202 10937
rect 20308 10862 20398 10937
rect 20151 10855 20398 10862
rect 20191 10675 20398 10855
rect 20151 10666 20398 10675
rect 20151 10591 20202 10666
rect 20308 10591 20398 10666
rect 20151 10584 20398 10591
rect 20191 10397 20398 10584
rect 20151 10388 20398 10397
rect 20151 10313 20202 10388
rect 20308 10313 20398 10388
rect 20151 10306 20398 10313
rect 1060 9484 1245 9626
rect 1060 9362 1072 9484
rect 1235 9362 1245 9484
rect 1060 9353 1245 9362
rect 3060 9484 3245 9626
rect 3060 9362 3072 9484
rect 3235 9362 3245 9484
rect 3060 9353 3245 9362
rect 5060 9484 5245 9626
rect 5060 9362 5072 9484
rect 5235 9362 5245 9484
rect 5060 9353 5245 9362
rect 7060 9484 7245 9626
rect 7060 9362 7072 9484
rect 7235 9362 7245 9484
rect 7060 9353 7245 9362
rect 9060 9484 9245 9626
rect 9060 9362 9072 9484
rect 9235 9362 9245 9484
rect 9060 9353 9245 9362
rect 11060 9484 11245 9626
rect 11060 9362 11072 9484
rect 11235 9362 11245 9484
rect 11060 9353 11245 9362
rect 13060 9484 13245 9626
rect 13060 9362 13072 9484
rect 13235 9362 13245 9484
rect 13060 9353 13245 9362
rect 15060 9484 15245 9626
rect 15060 9362 15072 9484
rect 15235 9362 15245 9484
rect 15060 9353 15245 9362
rect 17060 9484 17245 9626
rect 17060 9362 17072 9484
rect 17235 9362 17245 9484
rect 17060 9353 17245 9362
rect -957 9238 -942 9270
rect -910 9238 -898 9270
rect -866 9238 -854 9270
rect -822 9238 -810 9270
rect -778 9238 -750 9270
rect -957 9225 -750 9238
rect -957 9193 -942 9225
rect -910 9193 -898 9225
rect -866 9193 -854 9225
rect -822 9193 -810 9225
rect -778 9193 -750 9225
rect -957 9180 -750 9193
rect -957 9148 -942 9180
rect -910 9148 -898 9180
rect -866 9148 -854 9180
rect -822 9148 -810 9180
rect -778 9148 -750 9180
rect -957 8877 -750 9148
rect -957 8845 -943 8877
rect -768 8845 -750 8877
rect -957 8437 -750 8845
rect 17632 9270 17839 9494
rect 17632 9238 17660 9270
rect 17692 9238 17704 9270
rect 17736 9238 17748 9270
rect 17780 9238 17792 9270
rect 17824 9238 17839 9270
rect 17632 9225 17839 9238
rect 17632 9193 17660 9225
rect 17692 9193 17704 9225
rect 17736 9193 17748 9225
rect 17780 9193 17792 9225
rect 17824 9193 17839 9225
rect 17632 9180 17839 9193
rect 17632 9148 17660 9180
rect 17692 9148 17704 9180
rect 17736 9148 17748 9180
rect 17780 9148 17792 9180
rect 17824 9148 17839 9180
rect 17632 8877 17839 9148
rect 17632 8845 17650 8877
rect 17825 8874 17839 8877
rect 17870 9489 18077 9494
rect 17870 9457 17898 9489
rect 17930 9457 17942 9489
rect 17974 9457 17986 9489
rect 18018 9457 18030 9489
rect 18062 9457 18077 9489
rect 17870 9444 18077 9457
rect 17870 9412 17898 9444
rect 17930 9412 17942 9444
rect 17974 9412 17986 9444
rect 18018 9412 18030 9444
rect 18062 9412 18077 9444
rect 17870 9399 18077 9412
rect 17870 9367 17898 9399
rect 17930 9367 17942 9399
rect 17974 9367 17986 9399
rect 18018 9367 18030 9399
rect 18062 9367 18077 9399
rect 17632 8827 17661 8845
rect 17693 8827 17705 8845
rect 17737 8827 17749 8845
rect 17781 8827 17793 8845
rect 17825 8827 17840 8874
rect 17632 8814 17840 8827
rect 17632 8782 17661 8814
rect 17693 8782 17705 8814
rect 17737 8782 17749 8814
rect 17781 8782 17793 8814
rect 17825 8782 17840 8814
rect 17632 8769 17840 8782
rect 17632 8737 17661 8769
rect 17693 8737 17705 8769
rect 17737 8737 17749 8769
rect 17781 8737 17793 8769
rect 17825 8737 17840 8769
rect 17632 8733 17840 8737
rect -957 8405 -943 8437
rect -768 8405 -750 8437
rect 969 8412 1039 8442
rect 1471 8412 1541 8442
rect 1973 8412 2043 8442
rect 2475 8412 2545 8442
rect 2977 8412 3047 8442
rect 3479 8412 3549 8442
rect 3981 8412 4051 8442
rect 4483 8412 4553 8442
rect 4985 8412 5055 8442
rect 5487 8412 5557 8442
rect 5989 8412 6059 8442
rect 6491 8412 6561 8442
rect 6993 8412 7063 8442
rect 7495 8412 7565 8442
rect 7997 8412 8067 8442
rect 8499 8412 8569 8442
rect 9001 8412 9071 8442
rect 9503 8412 9573 8442
rect 10005 8412 10075 8442
rect 10507 8412 10577 8442
rect 11009 8412 11079 8442
rect 11511 8412 11581 8442
rect 12013 8412 12083 8442
rect 12515 8412 12585 8442
rect 13017 8412 13087 8442
rect 13519 8412 13589 8442
rect 14021 8412 14091 8442
rect 14523 8412 14593 8442
rect 15025 8412 15095 8442
rect 15527 8412 15597 8442
rect 16029 8412 16099 8442
rect 17632 8437 17839 8733
rect -957 7997 -750 8405
rect 17632 8405 17650 8437
rect 17825 8405 17839 8437
rect 969 8124 1039 8154
rect 1471 8124 1541 8154
rect 1973 8124 2043 8154
rect 2475 8124 2545 8154
rect 2977 8124 3047 8154
rect 3479 8124 3549 8154
rect 3981 8124 4051 8154
rect 4483 8124 4553 8154
rect 4985 8124 5055 8154
rect 5487 8124 5557 8154
rect 5989 8124 6059 8154
rect 6491 8124 6561 8154
rect 6993 8124 7063 8154
rect 7495 8124 7565 8154
rect 7997 8124 8067 8154
rect 8499 8124 8569 8154
rect 9001 8124 9071 8154
rect 9503 8124 9573 8154
rect 10005 8124 10075 8154
rect 10507 8124 10577 8154
rect 11009 8124 11079 8154
rect 11511 8124 11581 8154
rect 12013 8124 12083 8154
rect 12515 8124 12585 8154
rect 13017 8124 13087 8154
rect 13519 8124 13589 8154
rect 14021 8124 14091 8154
rect 14523 8124 14593 8154
rect 15025 8124 15095 8154
rect 15527 8124 15597 8154
rect 16029 8124 16099 8154
rect 594 7997 624 8067
rect 882 7997 912 8067
rect 1096 7997 1126 8067
rect 1384 7997 1414 8067
rect 1598 7997 1628 8067
rect 1886 7997 1916 8067
rect 2100 7997 2130 8067
rect 2388 7997 2418 8067
rect 2602 7997 2632 8067
rect 2890 7997 2920 8067
rect 3104 7997 3134 8067
rect 3392 7997 3422 8067
rect 3606 7997 3636 8067
rect 3894 7997 3924 8067
rect 4108 7997 4138 8067
rect 4396 7997 4426 8067
rect 4610 7997 4640 8067
rect 4898 7997 4928 8067
rect 5112 7997 5142 8067
rect 5400 7997 5430 8067
rect 5614 7997 5644 8067
rect 5902 7997 5932 8067
rect 6116 7997 6146 8067
rect 6404 7997 6434 8067
rect 6618 7997 6648 8067
rect 6906 7997 6936 8067
rect 7120 7997 7150 8067
rect 7408 7997 7438 8067
rect 7622 7997 7652 8067
rect 7910 7997 7940 8067
rect 8124 7997 8154 8067
rect 8412 7997 8442 8067
rect 8626 7997 8656 8067
rect 8914 7997 8944 8067
rect 9128 7997 9158 8067
rect 9416 7997 9446 8067
rect 9630 7997 9660 8067
rect 9918 7997 9948 8067
rect 10132 7997 10162 8067
rect 10420 7997 10450 8067
rect 10634 7997 10664 8067
rect 10922 7997 10952 8067
rect 11136 7997 11166 8067
rect 11424 7997 11454 8067
rect 11638 7997 11668 8067
rect 11926 7997 11956 8067
rect 12140 7997 12170 8067
rect 12428 7997 12458 8067
rect 12642 7997 12672 8067
rect 12930 7997 12960 8067
rect 13144 7997 13174 8067
rect 13432 7997 13462 8067
rect 13646 7997 13676 8067
rect 13934 7997 13964 8067
rect 14148 7997 14178 8067
rect 14436 7997 14466 8067
rect 14650 7997 14680 8067
rect 14938 7997 14968 8067
rect 15152 7997 15182 8067
rect 15440 7997 15470 8067
rect 15654 7997 15684 8067
rect 15942 7997 15972 8067
rect 16156 7997 16186 8067
rect 16444 7997 16474 8067
rect 17632 7997 17839 8405
rect -957 7965 -943 7997
rect -768 7965 -750 7997
rect -957 7557 -750 7965
rect 17632 7965 17650 7997
rect 17825 7965 17839 7997
rect 969 7910 1039 7940
rect 1471 7910 1541 7940
rect 1973 7910 2043 7940
rect 2475 7910 2545 7940
rect 2977 7910 3047 7940
rect 3479 7910 3549 7940
rect 3981 7910 4051 7940
rect 4483 7910 4553 7940
rect 4985 7910 5055 7940
rect 5487 7910 5557 7940
rect 5989 7910 6059 7940
rect 6491 7910 6561 7940
rect 6993 7910 7063 7940
rect 7495 7910 7565 7940
rect 7997 7910 8067 7940
rect 8499 7910 8569 7940
rect 9001 7910 9071 7940
rect 9503 7910 9573 7940
rect 10005 7910 10075 7940
rect 10507 7910 10577 7940
rect 11009 7910 11079 7940
rect 11511 7910 11581 7940
rect 12013 7910 12083 7940
rect 12515 7910 12585 7940
rect 13017 7910 13087 7940
rect 13519 7910 13589 7940
rect 14021 7910 14091 7940
rect 14523 7910 14593 7940
rect 15025 7910 15095 7940
rect 15527 7910 15597 7940
rect 16029 7910 16099 7940
rect 17632 7851 17839 7965
rect 17632 7819 17660 7851
rect 17692 7819 17704 7851
rect 17736 7819 17748 7851
rect 17780 7819 17792 7851
rect 17824 7819 17839 7851
rect 17632 7806 17839 7819
rect 17632 7774 17660 7806
rect 17692 7774 17704 7806
rect 17736 7774 17748 7806
rect 17780 7774 17792 7806
rect 17824 7774 17839 7806
rect 17632 7761 17839 7774
rect 17632 7729 17660 7761
rect 17692 7729 17704 7761
rect 17736 7729 17748 7761
rect 17780 7729 17792 7761
rect 17824 7729 17839 7761
rect 969 7622 1039 7652
rect 1471 7622 1541 7652
rect 1973 7622 2043 7652
rect 2475 7622 2545 7652
rect 2977 7622 3047 7652
rect 3479 7622 3549 7652
rect 3981 7622 4051 7652
rect 4483 7622 4553 7652
rect 4985 7622 5055 7652
rect 5487 7622 5557 7652
rect 5989 7622 6059 7652
rect 6491 7622 6561 7652
rect 6993 7622 7063 7652
rect 7495 7622 7565 7652
rect 7997 7622 8067 7652
rect 8499 7622 8569 7652
rect 9001 7622 9071 7652
rect 9503 7622 9573 7652
rect 10005 7622 10075 7652
rect 10507 7622 10577 7652
rect 11009 7622 11079 7652
rect 11511 7622 11581 7652
rect 12013 7622 12083 7652
rect 12515 7622 12585 7652
rect 13017 7622 13087 7652
rect 13519 7622 13589 7652
rect 14021 7622 14091 7652
rect 14523 7622 14593 7652
rect 15025 7622 15095 7652
rect 15527 7622 15597 7652
rect 16029 7622 16099 7652
rect -957 7525 -943 7557
rect -768 7525 -750 7557
rect -957 7117 -750 7525
rect 594 7495 624 7565
rect 882 7495 912 7565
rect 1096 7495 1126 7565
rect 1384 7495 1414 7565
rect 1598 7495 1628 7565
rect 1886 7495 1916 7565
rect 2100 7495 2130 7565
rect 2388 7495 2418 7565
rect 2602 7495 2632 7565
rect 2890 7495 2920 7565
rect 3104 7495 3134 7565
rect 3392 7495 3422 7565
rect 3606 7495 3636 7565
rect 3894 7495 3924 7565
rect 4108 7495 4138 7565
rect 4396 7495 4426 7565
rect 4610 7495 4640 7565
rect 4898 7495 4928 7565
rect 5112 7495 5142 7565
rect 5400 7495 5430 7565
rect 5614 7495 5644 7565
rect 5902 7495 5932 7565
rect 6116 7495 6146 7565
rect 6404 7495 6434 7565
rect 6618 7495 6648 7565
rect 6906 7495 6936 7565
rect 7120 7495 7150 7565
rect 7408 7495 7438 7565
rect 7622 7495 7652 7565
rect 7910 7495 7940 7565
rect 8124 7495 8154 7565
rect 8412 7495 8442 7565
rect 8626 7495 8656 7565
rect 8914 7495 8944 7565
rect 9128 7495 9158 7565
rect 9416 7495 9446 7565
rect 9630 7495 9660 7565
rect 9918 7495 9948 7565
rect 10132 7495 10162 7565
rect 10420 7495 10450 7565
rect 10634 7495 10664 7565
rect 10922 7495 10952 7565
rect 11136 7495 11166 7565
rect 11424 7495 11454 7565
rect 11638 7495 11668 7565
rect 11926 7495 11956 7565
rect 12140 7495 12170 7565
rect 12428 7495 12458 7565
rect 12642 7495 12672 7565
rect 12930 7495 12960 7565
rect 13144 7495 13174 7565
rect 13432 7495 13462 7565
rect 13646 7495 13676 7565
rect 13934 7495 13964 7565
rect 14148 7495 14178 7565
rect 14436 7495 14466 7565
rect 14650 7495 14680 7565
rect 14938 7495 14968 7565
rect 15152 7495 15182 7565
rect 15440 7495 15470 7565
rect 15654 7495 15684 7565
rect 15942 7495 15972 7565
rect 16156 7495 16186 7565
rect 16444 7495 16474 7565
rect 17632 7557 17839 7729
rect 17632 7525 17650 7557
rect 17825 7525 17839 7557
rect 969 7408 1039 7438
rect 1471 7408 1541 7438
rect 1973 7408 2043 7438
rect 2475 7408 2545 7438
rect 2977 7408 3047 7438
rect 3479 7408 3549 7438
rect 3981 7408 4051 7438
rect 4483 7408 4553 7438
rect 4985 7408 5055 7438
rect 5487 7408 5557 7438
rect 5989 7408 6059 7438
rect 6491 7408 6561 7438
rect 6993 7408 7063 7438
rect 7495 7408 7565 7438
rect 7997 7408 8067 7438
rect 8499 7408 8569 7438
rect 9001 7408 9071 7438
rect 9503 7408 9573 7438
rect 10005 7408 10075 7438
rect 10507 7408 10577 7438
rect 11009 7408 11079 7438
rect 11511 7408 11581 7438
rect 12013 7408 12083 7438
rect 12515 7408 12585 7438
rect 13017 7408 13087 7438
rect 13519 7408 13589 7438
rect 14021 7408 14091 7438
rect 14523 7408 14593 7438
rect 15025 7408 15095 7438
rect 15527 7408 15597 7438
rect 16029 7408 16099 7438
rect 969 7120 1039 7150
rect 1471 7120 1541 7150
rect 1973 7120 2043 7150
rect 2475 7120 2545 7150
rect 2977 7120 3047 7150
rect 3479 7120 3549 7150
rect 3981 7120 4051 7150
rect 4483 7120 4553 7150
rect 4985 7120 5055 7150
rect 5487 7120 5557 7150
rect 5989 7120 6059 7150
rect 6491 7120 6561 7150
rect 6993 7120 7063 7150
rect 7495 7120 7565 7150
rect 7997 7120 8067 7150
rect 8499 7120 8569 7150
rect 9001 7120 9071 7150
rect 9503 7120 9573 7150
rect 10005 7120 10075 7150
rect 10507 7120 10577 7150
rect 11009 7120 11079 7150
rect 11511 7120 11581 7150
rect 12013 7120 12083 7150
rect 12515 7120 12585 7150
rect 13017 7120 13087 7150
rect 13519 7120 13589 7150
rect 14021 7120 14091 7150
rect 14523 7120 14593 7150
rect 15025 7120 15095 7150
rect 15527 7120 15597 7150
rect 16029 7120 16099 7150
rect -957 7085 -943 7117
rect -768 7085 -750 7117
rect -957 6677 -750 7085
rect 17632 7117 17839 7525
rect 17632 7085 17650 7117
rect 17825 7085 17839 7117
rect 594 6993 624 7063
rect 882 6993 912 7063
rect 1096 6993 1126 7063
rect 1384 6993 1414 7063
rect 1598 6993 1628 7063
rect 1886 6993 1916 7063
rect 2100 6993 2130 7063
rect 2388 6993 2418 7063
rect 2602 6993 2632 7063
rect 2890 6993 2920 7063
rect 3104 6993 3134 7063
rect 3392 6993 3422 7063
rect 3606 6993 3636 7063
rect 3894 6993 3924 7063
rect 4108 6993 4138 7063
rect 4396 6993 4426 7063
rect 4610 6993 4640 7063
rect 4898 6993 4928 7063
rect 5112 6993 5142 7063
rect 5400 6993 5430 7063
rect 5614 6993 5644 7063
rect 5902 6993 5932 7063
rect 6116 6993 6146 7063
rect 6404 6993 6434 7063
rect 6618 6993 6648 7063
rect 6906 6993 6936 7063
rect 7120 6993 7150 7063
rect 7408 6993 7438 7063
rect 7622 6993 7652 7063
rect 7910 6993 7940 7063
rect 8124 6993 8154 7063
rect 8412 6993 8442 7063
rect 8626 6993 8656 7063
rect 8914 6993 8944 7063
rect 9128 6993 9158 7063
rect 9416 6993 9446 7063
rect 9630 6993 9660 7063
rect 9918 6993 9948 7063
rect 10132 6993 10162 7063
rect 10420 6993 10450 7063
rect 10634 6993 10664 7063
rect 10922 6993 10952 7063
rect 11136 6993 11166 7063
rect 11424 6993 11454 7063
rect 11638 6993 11668 7063
rect 11926 6993 11956 7063
rect 12140 6993 12170 7063
rect 12428 6993 12458 7063
rect 12642 6993 12672 7063
rect 12930 6993 12960 7063
rect 13144 6993 13174 7063
rect 13432 6993 13462 7063
rect 13646 6993 13676 7063
rect 13934 6993 13964 7063
rect 14148 6993 14178 7063
rect 14436 6993 14466 7063
rect 14650 6993 14680 7063
rect 14938 6993 14968 7063
rect 15152 6993 15182 7063
rect 15440 6993 15470 7063
rect 15654 6993 15684 7063
rect 15942 6993 15972 7063
rect 16156 6993 16186 7063
rect 16444 6993 16474 7063
rect 969 6906 1039 6936
rect 1471 6906 1541 6936
rect 1973 6906 2043 6936
rect 2475 6906 2545 6936
rect 2977 6906 3047 6936
rect 3479 6906 3549 6936
rect 3981 6906 4051 6936
rect 4483 6906 4553 6936
rect 4985 6906 5055 6936
rect 5487 6906 5557 6936
rect 5989 6906 6059 6936
rect 6491 6906 6561 6936
rect 6993 6906 7063 6936
rect 7495 6906 7565 6936
rect 7997 6906 8067 6936
rect 8499 6906 8569 6936
rect 9001 6906 9071 6936
rect 9503 6906 9573 6936
rect 10005 6906 10075 6936
rect 10507 6906 10577 6936
rect 11009 6906 11079 6936
rect 11511 6906 11581 6936
rect 12013 6906 12083 6936
rect 12515 6906 12585 6936
rect 13017 6906 13087 6936
rect 13519 6906 13589 6936
rect 14021 6906 14091 6936
rect 14523 6906 14593 6936
rect 15025 6906 15095 6936
rect 15527 6906 15597 6936
rect 16029 6906 16099 6936
rect -957 6645 -943 6677
rect -768 6645 -750 6677
rect 17632 6851 17839 7085
rect 17632 6819 17660 6851
rect 17692 6819 17704 6851
rect 17736 6819 17748 6851
rect 17780 6819 17792 6851
rect 17824 6819 17839 6851
rect 17632 6806 17839 6819
rect 17632 6774 17660 6806
rect 17692 6774 17704 6806
rect 17736 6774 17748 6806
rect 17780 6774 17792 6806
rect 17824 6774 17839 6806
rect 17632 6761 17839 6774
rect 17632 6729 17660 6761
rect 17692 6729 17704 6761
rect 17736 6729 17748 6761
rect 17780 6729 17792 6761
rect 17824 6729 17839 6761
rect 17632 6677 17839 6729
rect -957 6237 -750 6645
rect 969 6618 1039 6648
rect 1471 6618 1541 6648
rect 1973 6618 2043 6648
rect 2475 6618 2545 6648
rect 2977 6618 3047 6648
rect 3479 6618 3549 6648
rect 3981 6618 4051 6648
rect 4483 6618 4553 6648
rect 4985 6618 5055 6648
rect 5487 6618 5557 6648
rect 5989 6618 6059 6648
rect 6491 6618 6561 6648
rect 6993 6618 7063 6648
rect 7495 6618 7565 6648
rect 7997 6618 8067 6648
rect 8499 6618 8569 6648
rect 9001 6618 9071 6648
rect 9503 6618 9573 6648
rect 10005 6618 10075 6648
rect 10507 6618 10577 6648
rect 11009 6618 11079 6648
rect 11511 6618 11581 6648
rect 12013 6618 12083 6648
rect 12515 6618 12585 6648
rect 13017 6618 13087 6648
rect 13519 6618 13589 6648
rect 14021 6618 14091 6648
rect 14523 6618 14593 6648
rect 15025 6618 15095 6648
rect 15527 6618 15597 6648
rect 16029 6618 16099 6648
rect 17632 6645 17650 6677
rect 17825 6645 17839 6677
rect 594 6491 624 6561
rect 882 6491 912 6561
rect 1096 6491 1126 6561
rect 1384 6491 1414 6561
rect 1598 6491 1628 6561
rect 1886 6491 1916 6561
rect 2100 6491 2130 6561
rect 2388 6491 2418 6561
rect 2602 6491 2632 6561
rect 2890 6491 2920 6561
rect 3104 6491 3134 6561
rect 3392 6491 3422 6561
rect 3606 6491 3636 6561
rect 3894 6491 3924 6561
rect 4108 6491 4138 6561
rect 4396 6491 4426 6561
rect 4610 6491 4640 6561
rect 4898 6491 4928 6561
rect 5112 6491 5142 6561
rect 5400 6491 5430 6561
rect 5614 6491 5644 6561
rect 5902 6491 5932 6561
rect 6116 6491 6146 6561
rect 6404 6491 6434 6561
rect 6618 6491 6648 6561
rect 6906 6491 6936 6561
rect 7120 6491 7150 6561
rect 7408 6491 7438 6561
rect 7622 6491 7652 6561
rect 7910 6491 7940 6561
rect 8124 6491 8154 6561
rect 8412 6491 8442 6561
rect 8626 6491 8656 6561
rect 8914 6491 8944 6561
rect 9128 6491 9158 6561
rect 9416 6491 9446 6561
rect 9630 6491 9660 6561
rect 9918 6491 9948 6561
rect 10132 6491 10162 6561
rect 10420 6491 10450 6561
rect 10634 6491 10664 6561
rect 10922 6491 10952 6561
rect 11136 6491 11166 6561
rect 11424 6491 11454 6561
rect 11638 6491 11668 6561
rect 11926 6491 11956 6561
rect 12140 6491 12170 6561
rect 12428 6491 12458 6561
rect 12642 6491 12672 6561
rect 12930 6491 12960 6561
rect 13144 6491 13174 6561
rect 13432 6491 13462 6561
rect 13646 6491 13676 6561
rect 13934 6491 13964 6561
rect 14148 6491 14178 6561
rect 14436 6491 14466 6561
rect 14650 6491 14680 6561
rect 14938 6491 14968 6561
rect 15152 6491 15182 6561
rect 15440 6491 15470 6561
rect 15654 6491 15684 6561
rect 15942 6491 15972 6561
rect 16156 6491 16186 6561
rect 16444 6491 16474 6561
rect 969 6404 1039 6434
rect 1471 6404 1541 6434
rect 1973 6404 2043 6434
rect 2475 6404 2545 6434
rect 2977 6404 3047 6434
rect 3479 6404 3549 6434
rect 3981 6404 4051 6434
rect 4483 6404 4553 6434
rect 4985 6404 5055 6434
rect 5487 6404 5557 6434
rect 5989 6404 6059 6434
rect 6491 6404 6561 6434
rect 6993 6404 7063 6434
rect 7495 6404 7565 6434
rect 7997 6404 8067 6434
rect 8499 6404 8569 6434
rect 9001 6404 9071 6434
rect 9503 6404 9573 6434
rect 10005 6404 10075 6434
rect 10507 6404 10577 6434
rect 11009 6404 11079 6434
rect 11511 6404 11581 6434
rect 12013 6404 12083 6434
rect 12515 6404 12585 6434
rect 13017 6404 13087 6434
rect 13519 6404 13589 6434
rect 14021 6404 14091 6434
rect 14523 6404 14593 6434
rect 15025 6404 15095 6434
rect 15527 6404 15597 6434
rect 16029 6404 16099 6434
rect -957 6205 -943 6237
rect -768 6205 -750 6237
rect -957 5797 -750 6205
rect 969 6116 1039 6146
rect 1471 6116 1541 6146
rect 1973 6116 2043 6146
rect 2475 6116 2545 6146
rect 2977 6116 3047 6146
rect 3479 6116 3549 6146
rect 3981 6116 4051 6146
rect 4483 6116 4553 6146
rect 4985 6116 5055 6146
rect 5487 6116 5557 6146
rect 5989 6116 6059 6146
rect 6491 6116 6561 6146
rect 6993 6116 7063 6146
rect 7495 6116 7565 6146
rect 7997 6116 8067 6146
rect 8499 6116 8569 6146
rect 9001 6116 9071 6146
rect 9503 6116 9573 6146
rect 10005 6116 10075 6146
rect 10507 6116 10577 6146
rect 11009 6116 11079 6146
rect 11511 6116 11581 6146
rect 12013 6116 12083 6146
rect 12515 6116 12585 6146
rect 13017 6116 13087 6146
rect 13519 6116 13589 6146
rect 14021 6116 14091 6146
rect 14523 6116 14593 6146
rect 15025 6116 15095 6146
rect 15527 6116 15597 6146
rect 16029 6116 16099 6146
rect 594 5989 624 6059
rect 882 5989 912 6059
rect 1096 5989 1126 6059
rect 1384 5989 1414 6059
rect 1598 5989 1628 6059
rect 1886 5989 1916 6059
rect 2100 5989 2130 6059
rect 2388 5989 2418 6059
rect 2602 5989 2632 6059
rect 2890 5989 2920 6059
rect 3104 5989 3134 6059
rect 3392 5989 3422 6059
rect 3606 5989 3636 6059
rect 3894 5989 3924 6059
rect 4108 5989 4138 6059
rect 4396 5989 4426 6059
rect 4610 5989 4640 6059
rect 4898 5989 4928 6059
rect 5112 5989 5142 6059
rect 5400 5989 5430 6059
rect 5614 5989 5644 6059
rect 5902 5989 5932 6059
rect 6116 5989 6146 6059
rect 6404 5989 6434 6059
rect 6618 5989 6648 6059
rect 6906 5989 6936 6059
rect 7120 5989 7150 6059
rect 7408 5989 7438 6059
rect 7622 5989 7652 6059
rect 7910 5989 7940 6059
rect 8124 5989 8154 6059
rect 8412 5989 8442 6059
rect 8626 5989 8656 6059
rect 8914 5989 8944 6059
rect 9128 5989 9158 6059
rect 9416 5989 9446 6059
rect 9630 5989 9660 6059
rect 9918 5989 9948 6059
rect 10132 5989 10162 6059
rect 10420 5989 10450 6059
rect 10634 5989 10664 6059
rect 10922 5989 10952 6059
rect 11136 5989 11166 6059
rect 11424 5989 11454 6059
rect 11638 5989 11668 6059
rect 11926 5989 11956 6059
rect 12140 5989 12170 6059
rect 12428 5989 12458 6059
rect 12642 5989 12672 6059
rect 12930 5989 12960 6059
rect 13144 5989 13174 6059
rect 13432 5989 13462 6059
rect 13646 5989 13676 6059
rect 13934 5989 13964 6059
rect 14148 5989 14178 6059
rect 14436 5989 14466 6059
rect 14650 5989 14680 6059
rect 14938 5989 14968 6059
rect 15152 5989 15182 6059
rect 15440 5989 15470 6059
rect 15654 5989 15684 6059
rect 15942 5989 15972 6059
rect 16156 5989 16186 6059
rect 16444 5989 16474 6059
rect 969 5902 1039 5932
rect 1471 5902 1541 5932
rect 1973 5902 2043 5932
rect 2475 5902 2545 5932
rect 2977 5902 3047 5932
rect 3479 5902 3549 5932
rect 3981 5902 4051 5932
rect 4483 5902 4553 5932
rect 4985 5902 5055 5932
rect 5487 5902 5557 5932
rect 5989 5902 6059 5932
rect 6491 5902 6561 5932
rect 6993 5902 7063 5932
rect 7495 5902 7565 5932
rect 7997 5902 8067 5932
rect 8499 5902 8569 5932
rect 9001 5902 9071 5932
rect 9503 5902 9573 5932
rect 10005 5902 10075 5932
rect 10507 5902 10577 5932
rect 11009 5902 11079 5932
rect 11511 5902 11581 5932
rect 12013 5902 12083 5932
rect 12515 5902 12585 5932
rect 13017 5902 13087 5932
rect 13519 5902 13589 5932
rect 14021 5902 14091 5932
rect 14523 5902 14593 5932
rect 15025 5902 15095 5932
rect 15527 5902 15597 5932
rect 16029 5902 16099 5932
rect 17632 5904 17839 6645
rect 17870 8709 18077 9367
rect 20191 8946 20398 10306
rect 20151 8937 20398 8946
rect 20151 8862 20202 8937
rect 20308 8862 20398 8937
rect 20151 8855 20398 8862
rect 17870 8537 18151 8709
rect 20191 8675 20398 8855
rect 20151 8666 20398 8675
rect 20151 8591 20202 8666
rect 20308 8591 20398 8666
rect 20151 8584 20398 8591
rect 17870 8366 18077 8537
rect 20191 8397 20398 8584
rect 17870 8334 17898 8366
rect 17930 8334 17942 8366
rect 17974 8334 17986 8366
rect 18018 8334 18030 8366
rect 18062 8334 18077 8366
rect 17870 8321 18077 8334
rect 17870 8289 17898 8321
rect 17930 8289 17942 8321
rect 17974 8289 17986 8321
rect 18018 8289 18030 8321
rect 18062 8289 18077 8321
rect 20151 8388 20398 8397
rect 20151 8313 20202 8388
rect 20308 8313 20398 8388
rect 20151 8306 20398 8313
rect 17870 8276 18077 8289
rect 17870 8244 17898 8276
rect 17930 8244 17942 8276
rect 17974 8244 17986 8276
rect 18018 8244 18030 8276
rect 18062 8244 18077 8276
rect 17870 7312 18077 8244
rect 17870 7280 17898 7312
rect 17930 7280 17942 7312
rect 17974 7280 17986 7312
rect 18018 7280 18030 7312
rect 18062 7280 18077 7312
rect 17870 7267 18077 7280
rect 17870 7235 17898 7267
rect 17930 7235 17942 7267
rect 17974 7235 17986 7267
rect 18018 7235 18030 7267
rect 18062 7235 18077 7267
rect 17870 7222 18077 7235
rect 17870 7190 17898 7222
rect 17930 7190 17942 7222
rect 17974 7190 17986 7222
rect 18018 7190 18030 7222
rect 18062 7190 18077 7222
rect 17870 6709 18077 7190
rect 20191 6946 20398 8306
rect 20151 6937 20398 6946
rect 20151 6862 20202 6937
rect 20308 6862 20398 6937
rect 20151 6855 20398 6862
rect 17870 6537 18151 6709
rect 20191 6675 20398 6855
rect 20151 6666 20398 6675
rect 20151 6591 20202 6666
rect 20308 6591 20398 6666
rect 20151 6584 20398 6591
rect 17870 6361 18077 6537
rect 20191 6397 20398 6584
rect 17869 6347 18077 6361
rect 17869 6315 17897 6347
rect 17929 6315 17941 6347
rect 17973 6315 17985 6347
rect 18017 6315 18029 6347
rect 18061 6315 18077 6347
rect 17869 6302 18077 6315
rect 20151 6388 20398 6397
rect 20151 6313 20202 6388
rect 20308 6313 20398 6388
rect 20151 6306 20398 6313
rect 17869 6270 17897 6302
rect 17929 6270 17941 6302
rect 17973 6270 17985 6302
rect 18017 6270 18029 6302
rect 18061 6270 18077 6302
rect 17869 6257 18077 6270
rect 17869 6225 17897 6257
rect 17929 6225 17941 6257
rect 17973 6225 17985 6257
rect 18017 6225 18029 6257
rect 18061 6225 18077 6257
rect 17869 6221 18077 6225
rect -957 5765 -943 5797
rect -768 5765 -750 5797
rect -957 5357 -750 5765
rect 17632 5889 17840 5904
rect 17632 5857 17661 5889
rect 17693 5857 17705 5889
rect 17737 5857 17749 5889
rect 17781 5857 17793 5889
rect 17825 5857 17840 5889
rect 17632 5844 17840 5857
rect 17632 5812 17661 5844
rect 17693 5812 17705 5844
rect 17737 5812 17749 5844
rect 17781 5812 17793 5844
rect 17825 5812 17840 5844
rect 17632 5799 17840 5812
rect 17632 5797 17661 5799
rect 17693 5797 17705 5799
rect 17737 5797 17749 5799
rect 17781 5797 17793 5799
rect 17632 5765 17650 5797
rect 17825 5765 17840 5799
rect 17632 5763 17840 5765
rect 969 5614 1039 5644
rect 1471 5614 1541 5644
rect 1973 5614 2043 5644
rect 2475 5614 2545 5644
rect 2977 5614 3047 5644
rect 3479 5614 3549 5644
rect 3981 5614 4051 5644
rect 4483 5614 4553 5644
rect 4985 5614 5055 5644
rect 5487 5614 5557 5644
rect 5989 5614 6059 5644
rect 6491 5614 6561 5644
rect 6993 5614 7063 5644
rect 7495 5614 7565 5644
rect 7997 5614 8067 5644
rect 8499 5614 8569 5644
rect 9001 5614 9071 5644
rect 9503 5614 9573 5644
rect 10005 5614 10075 5644
rect 10507 5614 10577 5644
rect 11009 5614 11079 5644
rect 11511 5614 11581 5644
rect 12013 5614 12083 5644
rect 12515 5614 12585 5644
rect 13017 5614 13087 5644
rect 13519 5614 13589 5644
rect 14021 5614 14091 5644
rect 14523 5614 14593 5644
rect 15025 5614 15095 5644
rect 15527 5614 15597 5644
rect 16029 5614 16099 5644
rect 594 5487 624 5557
rect 882 5487 912 5557
rect 1096 5487 1126 5557
rect 1384 5487 1414 5557
rect 1598 5487 1628 5557
rect 1886 5487 1916 5557
rect 2100 5487 2130 5557
rect 2388 5487 2418 5557
rect 2602 5487 2632 5557
rect 2890 5487 2920 5557
rect 3104 5487 3134 5557
rect 3392 5487 3422 5557
rect 3606 5487 3636 5557
rect 3894 5487 3924 5557
rect 4108 5487 4138 5557
rect 4396 5487 4426 5557
rect 4610 5487 4640 5557
rect 4898 5487 4928 5557
rect 5112 5487 5142 5557
rect 5400 5487 5430 5557
rect 5614 5487 5644 5557
rect 5902 5487 5932 5557
rect 6116 5487 6146 5557
rect 6404 5487 6434 5557
rect 6618 5487 6648 5557
rect 6906 5487 6936 5557
rect 7120 5487 7150 5557
rect 7408 5487 7438 5557
rect 7622 5487 7652 5557
rect 7910 5487 7940 5557
rect 8124 5487 8154 5557
rect 8412 5487 8442 5557
rect 8626 5487 8656 5557
rect 8914 5487 8944 5557
rect 9128 5487 9158 5557
rect 9416 5487 9446 5557
rect 9630 5487 9660 5557
rect 9918 5487 9948 5557
rect 10132 5487 10162 5557
rect 10420 5487 10450 5557
rect 10634 5487 10664 5557
rect 10922 5487 10952 5557
rect 11136 5487 11166 5557
rect 11424 5487 11454 5557
rect 11638 5487 11668 5557
rect 11926 5487 11956 5557
rect 12140 5487 12170 5557
rect 12428 5487 12458 5557
rect 12642 5487 12672 5557
rect 12930 5487 12960 5557
rect 13144 5487 13174 5557
rect 13432 5487 13462 5557
rect 13646 5487 13676 5557
rect 13934 5487 13964 5557
rect 14148 5487 14178 5557
rect 14436 5487 14466 5557
rect 14650 5487 14680 5557
rect 14938 5487 14968 5557
rect 15152 5487 15182 5557
rect 15440 5487 15470 5557
rect 15654 5487 15684 5557
rect 15942 5487 15972 5557
rect 16156 5487 16186 5557
rect 16444 5487 16474 5557
rect 969 5400 1039 5430
rect 1471 5400 1541 5430
rect 1973 5400 2043 5430
rect 2475 5400 2545 5430
rect 2977 5400 3047 5430
rect 3479 5400 3549 5430
rect 3981 5400 4051 5430
rect 4483 5400 4553 5430
rect 4985 5400 5055 5430
rect 5487 5400 5557 5430
rect 5989 5400 6059 5430
rect 6491 5400 6561 5430
rect 6993 5400 7063 5430
rect 7495 5400 7565 5430
rect 7997 5400 8067 5430
rect 8499 5400 8569 5430
rect 9001 5400 9071 5430
rect 9503 5400 9573 5430
rect 10005 5400 10075 5430
rect 10507 5400 10577 5430
rect 11009 5400 11079 5430
rect 11511 5400 11581 5430
rect 12013 5400 12083 5430
rect 12515 5400 12585 5430
rect 13017 5400 13087 5430
rect 13519 5400 13589 5430
rect 14021 5400 14091 5430
rect 14523 5400 14593 5430
rect 15025 5400 15095 5430
rect 15527 5400 15597 5430
rect 16029 5400 16099 5430
rect -957 5325 -943 5357
rect -768 5325 -750 5357
rect -957 4917 -750 5325
rect 969 5112 1039 5142
rect 1471 5112 1541 5142
rect 1973 5112 2043 5142
rect 2475 5112 2545 5142
rect 2977 5112 3047 5142
rect 3479 5112 3549 5142
rect 3981 5112 4051 5142
rect 4483 5112 4553 5142
rect 4985 5112 5055 5142
rect 5487 5112 5557 5142
rect 5989 5112 6059 5142
rect 6491 5112 6561 5142
rect 6993 5112 7063 5142
rect 7495 5112 7565 5142
rect 7997 5112 8067 5142
rect 8499 5112 8569 5142
rect 9001 5112 9071 5142
rect 9503 5112 9573 5142
rect 10005 5112 10075 5142
rect 10507 5112 10577 5142
rect 11009 5112 11079 5142
rect 11511 5112 11581 5142
rect 12013 5112 12083 5142
rect 12515 5112 12585 5142
rect 13017 5112 13087 5142
rect 13519 5112 13589 5142
rect 14021 5112 14091 5142
rect 14523 5112 14593 5142
rect 15025 5112 15095 5142
rect 15527 5112 15597 5142
rect 16029 5112 16099 5142
rect 594 4985 624 5055
rect 882 4985 912 5055
rect 1096 4985 1126 5055
rect 1384 4985 1414 5055
rect 1598 4985 1628 5055
rect 1886 4985 1916 5055
rect 2100 4985 2130 5055
rect 2388 4985 2418 5055
rect 2602 4985 2632 5055
rect 2890 4985 2920 5055
rect 3104 4985 3134 5055
rect 3392 4985 3422 5055
rect 3606 4985 3636 5055
rect 3894 4985 3924 5055
rect 4108 4985 4138 5055
rect 4396 4985 4426 5055
rect 4610 4985 4640 5055
rect 4898 4985 4928 5055
rect 5112 4985 5142 5055
rect 5400 4985 5430 5055
rect 5614 4985 5644 5055
rect 5902 4985 5932 5055
rect 6116 4985 6146 5055
rect 6404 4985 6434 5055
rect 6618 4985 6648 5055
rect 6906 4985 6936 5055
rect 7120 4985 7150 5055
rect 7408 4985 7438 5055
rect 7622 4985 7652 5055
rect 7910 4985 7940 5055
rect 8124 4985 8154 5055
rect 8412 4985 8442 5055
rect 8626 4985 8656 5055
rect 8914 4985 8944 5055
rect 9128 4985 9158 5055
rect 9416 4985 9446 5055
rect 9630 4985 9660 5055
rect 9918 4985 9948 5055
rect 10132 4985 10162 5055
rect 10420 4985 10450 5055
rect 10634 4985 10664 5055
rect 10922 4985 10952 5055
rect 11136 4985 11166 5055
rect 11424 4985 11454 5055
rect 11638 4985 11668 5055
rect 11926 4985 11956 5055
rect 12140 4985 12170 5055
rect 12428 4985 12458 5055
rect 12642 4985 12672 5055
rect 12930 4985 12960 5055
rect 13144 4985 13174 5055
rect 13432 4985 13462 5055
rect 13646 4985 13676 5055
rect 13934 4985 13964 5055
rect 14148 4985 14178 5055
rect 14436 4985 14466 5055
rect 14650 4985 14680 5055
rect 14938 4985 14968 5055
rect 15152 4985 15182 5055
rect 15440 4985 15470 5055
rect 15654 4985 15684 5055
rect 15942 4985 15972 5055
rect 16156 4985 16186 5055
rect 16444 4985 16474 5055
rect -957 4885 -943 4917
rect -768 4885 -750 4917
rect 969 4898 1039 4928
rect 1471 4898 1541 4928
rect 1973 4898 2043 4928
rect 2475 4898 2545 4928
rect 2977 4898 3047 4928
rect 3479 4898 3549 4928
rect 3981 4898 4051 4928
rect 4483 4898 4553 4928
rect 4985 4898 5055 4928
rect 5487 4898 5557 4928
rect 5989 4898 6059 4928
rect 6491 4898 6561 4928
rect 6993 4898 7063 4928
rect 7495 4898 7565 4928
rect 7997 4898 8067 4928
rect 8499 4898 8569 4928
rect 9001 4898 9071 4928
rect 9503 4898 9573 4928
rect 10005 4898 10075 4928
rect 10507 4898 10577 4928
rect 11009 4898 11079 4928
rect 11511 4898 11581 4928
rect 12013 4898 12083 4928
rect 12515 4898 12585 4928
rect 13017 4898 13087 4928
rect 13519 4898 13589 4928
rect 14021 4898 14091 4928
rect 14523 4898 14593 4928
rect 15025 4898 15095 4928
rect 15527 4898 15597 4928
rect 16029 4898 16099 4928
rect 17632 4917 17839 5763
rect -957 4477 -750 4885
rect 17632 4885 17650 4917
rect 17825 4885 17839 4917
rect 17632 4826 17839 4885
rect 17632 4794 17660 4826
rect 17692 4794 17704 4826
rect 17736 4794 17748 4826
rect 17780 4794 17792 4826
rect 17824 4794 17839 4826
rect 17632 4781 17839 4794
rect 17632 4749 17660 4781
rect 17692 4749 17704 4781
rect 17736 4749 17748 4781
rect 17780 4749 17792 4781
rect 17824 4749 17839 4781
rect 17632 4736 17839 4749
rect 17632 4704 17660 4736
rect 17692 4704 17704 4736
rect 17736 4704 17748 4736
rect 17780 4704 17792 4736
rect 17824 4704 17839 4736
rect 969 4610 1039 4640
rect 1471 4610 1541 4640
rect 1973 4610 2043 4640
rect 2475 4610 2545 4640
rect 2977 4610 3047 4640
rect 3479 4610 3549 4640
rect 3981 4610 4051 4640
rect 4483 4610 4553 4640
rect 4985 4610 5055 4640
rect 5487 4610 5557 4640
rect 5989 4610 6059 4640
rect 6491 4610 6561 4640
rect 6993 4610 7063 4640
rect 7495 4610 7565 4640
rect 7997 4610 8067 4640
rect 8499 4610 8569 4640
rect 9001 4610 9071 4640
rect 9503 4610 9573 4640
rect 10005 4610 10075 4640
rect 10507 4610 10577 4640
rect 11009 4610 11079 4640
rect 11511 4610 11581 4640
rect 12013 4610 12083 4640
rect 12515 4610 12585 4640
rect 13017 4610 13087 4640
rect 13519 4610 13589 4640
rect 14021 4610 14091 4640
rect 14523 4610 14593 4640
rect 15025 4610 15095 4640
rect 15527 4610 15597 4640
rect 16029 4610 16099 4640
rect 594 4483 624 4553
rect 882 4483 912 4553
rect 1096 4483 1126 4553
rect 1384 4483 1414 4553
rect 1598 4483 1628 4553
rect 1886 4483 1916 4553
rect 2100 4483 2130 4553
rect 2388 4483 2418 4553
rect 2602 4483 2632 4553
rect 2890 4483 2920 4553
rect 3104 4483 3134 4553
rect 3392 4483 3422 4553
rect 3606 4483 3636 4553
rect 3894 4483 3924 4553
rect 4108 4483 4138 4553
rect 4396 4483 4426 4553
rect 4610 4483 4640 4553
rect 4898 4483 4928 4553
rect 5112 4483 5142 4553
rect 5400 4483 5430 4553
rect 5614 4483 5644 4553
rect 5902 4483 5932 4553
rect 6116 4483 6146 4553
rect 6404 4483 6434 4553
rect 6618 4483 6648 4553
rect 6906 4483 6936 4553
rect 7120 4483 7150 4553
rect 7408 4483 7438 4553
rect 7622 4483 7652 4553
rect 7910 4483 7940 4553
rect 8124 4483 8154 4553
rect 8412 4483 8442 4553
rect 8626 4483 8656 4553
rect 8914 4483 8944 4553
rect 9128 4483 9158 4553
rect 9416 4483 9446 4553
rect 9630 4483 9660 4553
rect 9918 4483 9948 4553
rect 10132 4483 10162 4553
rect 10420 4483 10450 4553
rect 10634 4483 10664 4553
rect 10922 4483 10952 4553
rect 11136 4483 11166 4553
rect 11424 4483 11454 4553
rect 11638 4483 11668 4553
rect 11926 4483 11956 4553
rect 12140 4483 12170 4553
rect 12428 4483 12458 4553
rect 12642 4483 12672 4553
rect 12930 4483 12960 4553
rect 13144 4483 13174 4553
rect 13432 4483 13462 4553
rect 13646 4483 13676 4553
rect 13934 4483 13964 4553
rect 14148 4483 14178 4553
rect 14436 4483 14466 4553
rect 14650 4483 14680 4553
rect 14938 4483 14968 4553
rect 15152 4483 15182 4553
rect 15440 4483 15470 4553
rect 15654 4483 15684 4553
rect 15942 4483 15972 4553
rect 16156 4483 16186 4553
rect 16444 4483 16474 4553
rect -957 4445 -943 4477
rect -768 4445 -750 4477
rect -957 4037 -750 4445
rect 17632 4477 17839 4704
rect 17632 4445 17650 4477
rect 17825 4445 17839 4477
rect 969 4396 1039 4426
rect 1471 4396 1541 4426
rect 1973 4396 2043 4426
rect 2475 4396 2545 4426
rect 2977 4396 3047 4426
rect 3479 4396 3549 4426
rect 3981 4396 4051 4426
rect 4483 4396 4553 4426
rect 4985 4396 5055 4426
rect 5487 4396 5557 4426
rect 5989 4396 6059 4426
rect 6491 4396 6561 4426
rect 6993 4396 7063 4426
rect 7495 4396 7565 4426
rect 7997 4396 8067 4426
rect 8499 4396 8569 4426
rect 9001 4396 9071 4426
rect 9503 4396 9573 4426
rect 10005 4396 10075 4426
rect 10507 4396 10577 4426
rect 11009 4396 11079 4426
rect 11511 4396 11581 4426
rect 12013 4396 12083 4426
rect 12515 4396 12585 4426
rect 13017 4396 13087 4426
rect 13519 4396 13589 4426
rect 14021 4396 14091 4426
rect 14523 4396 14593 4426
rect 15025 4396 15095 4426
rect 15527 4396 15597 4426
rect 16029 4396 16099 4426
rect 969 4108 1039 4138
rect 1471 4108 1541 4138
rect 1973 4108 2043 4138
rect 2475 4108 2545 4138
rect 2977 4108 3047 4138
rect 3479 4108 3549 4138
rect 3981 4108 4051 4138
rect 4483 4108 4553 4138
rect 4985 4108 5055 4138
rect 5487 4108 5557 4138
rect 5989 4108 6059 4138
rect 6491 4108 6561 4138
rect 6993 4108 7063 4138
rect 7495 4108 7565 4138
rect 7997 4108 8067 4138
rect 8499 4108 8569 4138
rect 9001 4108 9071 4138
rect 9503 4108 9573 4138
rect 10005 4108 10075 4138
rect 10507 4108 10577 4138
rect 11009 4108 11079 4138
rect 11511 4108 11581 4138
rect 12013 4108 12083 4138
rect 12515 4108 12585 4138
rect 13017 4108 13087 4138
rect 13519 4108 13589 4138
rect 14021 4108 14091 4138
rect 14523 4108 14593 4138
rect 15025 4108 15095 4138
rect 15527 4108 15597 4138
rect 16029 4108 16099 4138
rect -957 4005 -943 4037
rect -768 4005 -750 4037
rect -957 3597 -750 4005
rect 594 3981 624 4051
rect 882 3981 912 4051
rect 1096 3981 1126 4051
rect 1384 3981 1414 4051
rect 1598 3981 1628 4051
rect 1886 3981 1916 4051
rect 2100 3981 2130 4051
rect 2388 3981 2418 4051
rect 2602 3981 2632 4051
rect 2890 3981 2920 4051
rect 3104 3981 3134 4051
rect 3392 3981 3422 4051
rect 3606 3981 3636 4051
rect 3894 3981 3924 4051
rect 4108 3981 4138 4051
rect 4396 3981 4426 4051
rect 4610 3981 4640 4051
rect 4898 3981 4928 4051
rect 5112 3981 5142 4051
rect 5400 3981 5430 4051
rect 5614 3981 5644 4051
rect 5902 3981 5932 4051
rect 6116 3981 6146 4051
rect 6404 3981 6434 4051
rect 6618 3981 6648 4051
rect 6906 3981 6936 4051
rect 7120 3981 7150 4051
rect 7408 3981 7438 4051
rect 7622 3981 7652 4051
rect 7910 3981 7940 4051
rect 8124 3981 8154 4051
rect 8412 3981 8442 4051
rect 8626 3981 8656 4051
rect 8914 3981 8944 4051
rect 9128 3981 9158 4051
rect 9416 3981 9446 4051
rect 9630 3981 9660 4051
rect 9918 3981 9948 4051
rect 10132 3981 10162 4051
rect 10420 3981 10450 4051
rect 10634 3981 10664 4051
rect 10922 3981 10952 4051
rect 11136 3981 11166 4051
rect 11424 3981 11454 4051
rect 11638 3981 11668 4051
rect 11926 3981 11956 4051
rect 12140 3981 12170 4051
rect 12428 3981 12458 4051
rect 12642 3981 12672 4051
rect 12930 3981 12960 4051
rect 13144 3981 13174 4051
rect 13432 3981 13462 4051
rect 13646 3981 13676 4051
rect 13934 3981 13964 4051
rect 14148 3981 14178 4051
rect 14436 3981 14466 4051
rect 14650 3981 14680 4051
rect 14938 3981 14968 4051
rect 15152 3981 15182 4051
rect 15440 3981 15470 4051
rect 15654 3981 15684 4051
rect 15942 3981 15972 4051
rect 16156 3981 16186 4051
rect 16444 3981 16474 4051
rect 17632 4037 17839 4445
rect 17632 4005 17650 4037
rect 17825 4005 17839 4037
rect 969 3894 1039 3924
rect 1471 3894 1541 3924
rect 1973 3894 2043 3924
rect 2475 3894 2545 3924
rect 2977 3894 3047 3924
rect 3479 3894 3549 3924
rect 3981 3894 4051 3924
rect 4483 3894 4553 3924
rect 4985 3894 5055 3924
rect 5487 3894 5557 3924
rect 5989 3894 6059 3924
rect 6491 3894 6561 3924
rect 6993 3894 7063 3924
rect 7495 3894 7565 3924
rect 7997 3894 8067 3924
rect 8499 3894 8569 3924
rect 9001 3894 9071 3924
rect 9503 3894 9573 3924
rect 10005 3894 10075 3924
rect 10507 3894 10577 3924
rect 11009 3894 11079 3924
rect 11511 3894 11581 3924
rect 12013 3894 12083 3924
rect 12515 3894 12585 3924
rect 13017 3894 13087 3924
rect 13519 3894 13589 3924
rect 14021 3894 14091 3924
rect 14523 3894 14593 3924
rect 15025 3894 15095 3924
rect 15527 3894 15597 3924
rect 16029 3894 16099 3924
rect 17632 3853 17839 4005
rect 17870 5339 18077 6221
rect 17870 5307 17898 5339
rect 17930 5307 17942 5339
rect 17974 5307 17986 5339
rect 18018 5307 18030 5339
rect 18062 5307 18077 5339
rect 17870 5294 18077 5307
rect 17870 5262 17898 5294
rect 17930 5262 17942 5294
rect 17974 5262 17986 5294
rect 18018 5262 18030 5294
rect 18062 5262 18077 5294
rect 17870 5249 18077 5262
rect 17870 5217 17898 5249
rect 17930 5217 17942 5249
rect 17974 5217 17986 5249
rect 18018 5217 18030 5249
rect 18062 5217 18077 5249
rect 17870 4709 18077 5217
rect 20191 4946 20398 6306
rect 20151 4937 20398 4946
rect 20151 4862 20202 4937
rect 20308 4862 20398 4937
rect 20151 4855 20398 4862
rect 17870 4537 18151 4709
rect 20191 4675 20398 4855
rect 20151 4666 20398 4675
rect 20151 4591 20202 4666
rect 20308 4591 20398 4666
rect 20151 4584 20398 4591
rect 17870 4338 18077 4537
rect 20191 4397 20398 4584
rect 17870 4306 17898 4338
rect 17930 4306 17942 4338
rect 17974 4306 17986 4338
rect 18018 4306 18030 4338
rect 18062 4306 18077 4338
rect 20151 4388 20398 4397
rect 20151 4313 20202 4388
rect 20308 4313 20398 4388
rect 20151 4306 20398 4313
rect 17870 4293 18077 4306
rect 17870 4261 17898 4293
rect 17930 4261 17942 4293
rect 17974 4261 17986 4293
rect 18018 4261 18030 4293
rect 18062 4261 18077 4293
rect 17870 4248 18077 4261
rect 17870 4216 17898 4248
rect 17930 4216 17942 4248
rect 17974 4216 17986 4248
rect 18018 4216 18030 4248
rect 18062 4216 18077 4248
rect 17632 3838 17840 3853
rect 17632 3806 17661 3838
rect 17693 3806 17705 3838
rect 17737 3806 17749 3838
rect 17781 3806 17793 3838
rect 17825 3806 17840 3838
rect 17632 3793 17840 3806
rect 17632 3761 17661 3793
rect 17693 3761 17705 3793
rect 17737 3761 17749 3793
rect 17781 3761 17793 3793
rect 17825 3761 17840 3793
rect 17632 3748 17840 3761
rect 17632 3716 17661 3748
rect 17693 3716 17705 3748
rect 17737 3716 17749 3748
rect 17781 3716 17793 3748
rect 17825 3716 17840 3748
rect 17632 3712 17840 3716
rect 969 3606 1039 3636
rect 1471 3606 1541 3636
rect 1973 3606 2043 3636
rect 2475 3606 2545 3636
rect 2977 3606 3047 3636
rect 3479 3606 3549 3636
rect 3981 3606 4051 3636
rect 4483 3606 4553 3636
rect 4985 3606 5055 3636
rect 5487 3606 5557 3636
rect 5989 3606 6059 3636
rect 6491 3606 6561 3636
rect 6993 3606 7063 3636
rect 7495 3606 7565 3636
rect 7997 3606 8067 3636
rect 8499 3606 8569 3636
rect 9001 3606 9071 3636
rect 9503 3606 9573 3636
rect 10005 3606 10075 3636
rect 10507 3606 10577 3636
rect 11009 3606 11079 3636
rect 11511 3606 11581 3636
rect 12013 3606 12083 3636
rect 12515 3606 12585 3636
rect 13017 3606 13087 3636
rect 13519 3606 13589 3636
rect 14021 3606 14091 3636
rect 14523 3606 14593 3636
rect 15025 3606 15095 3636
rect 15527 3606 15597 3636
rect 16029 3606 16099 3636
rect -957 3565 -943 3597
rect -768 3565 -750 3597
rect -957 3157 -750 3565
rect 17632 3597 17839 3712
rect 17632 3565 17650 3597
rect 17825 3565 17839 3597
rect 594 3479 624 3549
rect 882 3479 912 3549
rect 1096 3479 1126 3549
rect 1384 3479 1414 3549
rect 1598 3479 1628 3549
rect 1886 3479 1916 3549
rect 2100 3479 2130 3549
rect 2388 3479 2418 3549
rect 2602 3479 2632 3549
rect 2890 3479 2920 3549
rect 3104 3479 3134 3549
rect 3392 3479 3422 3549
rect 3606 3479 3636 3549
rect 3894 3479 3924 3549
rect 4108 3479 4138 3549
rect 4396 3479 4426 3549
rect 4610 3479 4640 3549
rect 4898 3479 4928 3549
rect 5112 3479 5142 3549
rect 5400 3479 5430 3549
rect 5614 3479 5644 3549
rect 5902 3479 5932 3549
rect 6116 3479 6146 3549
rect 6404 3479 6434 3549
rect 6618 3479 6648 3549
rect 6906 3479 6936 3549
rect 7120 3479 7150 3549
rect 7408 3479 7438 3549
rect 7622 3479 7652 3549
rect 7910 3479 7940 3549
rect 8124 3479 8154 3549
rect 8412 3479 8442 3549
rect 8626 3479 8656 3549
rect 8914 3479 8944 3549
rect 9128 3479 9158 3549
rect 9416 3479 9446 3549
rect 9630 3479 9660 3549
rect 9918 3479 9948 3549
rect 10132 3479 10162 3549
rect 10420 3479 10450 3549
rect 10634 3479 10664 3549
rect 10922 3479 10952 3549
rect 11136 3479 11166 3549
rect 11424 3479 11454 3549
rect 11638 3479 11668 3549
rect 11926 3479 11956 3549
rect 12140 3479 12170 3549
rect 12428 3479 12458 3549
rect 12642 3479 12672 3549
rect 12930 3479 12960 3549
rect 13144 3479 13174 3549
rect 13432 3479 13462 3549
rect 13646 3479 13676 3549
rect 13934 3479 13964 3549
rect 14148 3479 14178 3549
rect 14436 3479 14466 3549
rect 14650 3479 14680 3549
rect 14938 3479 14968 3549
rect 15152 3479 15182 3549
rect 15440 3479 15470 3549
rect 15654 3479 15684 3549
rect 15942 3479 15972 3549
rect 16156 3479 16186 3549
rect 16444 3479 16474 3549
rect 969 3392 1039 3422
rect 1471 3392 1541 3422
rect 1973 3392 2043 3422
rect 2475 3392 2545 3422
rect 2977 3392 3047 3422
rect 3479 3392 3549 3422
rect 3981 3392 4051 3422
rect 4483 3392 4553 3422
rect 4985 3392 5055 3422
rect 5487 3392 5557 3422
rect 5989 3392 6059 3422
rect 6491 3392 6561 3422
rect 6993 3392 7063 3422
rect 7495 3392 7565 3422
rect 7997 3392 8067 3422
rect 8499 3392 8569 3422
rect 9001 3392 9071 3422
rect 9503 3392 9573 3422
rect 10005 3392 10075 3422
rect 10507 3392 10577 3422
rect 11009 3392 11079 3422
rect 11511 3392 11581 3422
rect 12013 3392 12083 3422
rect 12515 3392 12585 3422
rect 13017 3392 13087 3422
rect 13519 3392 13589 3422
rect 14021 3392 14091 3422
rect 14523 3392 14593 3422
rect 15025 3392 15095 3422
rect 15527 3392 15597 3422
rect 16029 3392 16099 3422
rect -957 3125 -943 3157
rect -768 3125 -750 3157
rect 17632 3157 17839 3565
rect 17870 3353 18077 4216
rect 17869 3339 18077 3353
rect 17869 3307 17897 3339
rect 17929 3307 17941 3339
rect 17973 3307 17985 3339
rect 18017 3307 18029 3339
rect 18061 3307 18077 3339
rect 17869 3294 18077 3307
rect 17869 3262 17897 3294
rect 17929 3262 17941 3294
rect 17973 3262 17985 3294
rect 18017 3262 18029 3294
rect 18061 3262 18077 3294
rect 17869 3249 18077 3262
rect 17869 3217 17897 3249
rect 17929 3217 17941 3249
rect 17973 3217 17985 3249
rect 18017 3217 18029 3249
rect 18061 3217 18077 3249
rect 17869 3213 18077 3217
rect -957 2717 -750 3125
rect 969 3104 1039 3134
rect 1471 3104 1541 3134
rect 1973 3104 2043 3134
rect 2475 3104 2545 3134
rect 2977 3104 3047 3134
rect 3479 3104 3549 3134
rect 3981 3104 4051 3134
rect 4483 3104 4553 3134
rect 4985 3104 5055 3134
rect 5487 3104 5557 3134
rect 5989 3104 6059 3134
rect 6491 3104 6561 3134
rect 6993 3104 7063 3134
rect 7495 3104 7565 3134
rect 7997 3104 8067 3134
rect 8499 3104 8569 3134
rect 9001 3104 9071 3134
rect 9503 3104 9573 3134
rect 10005 3104 10075 3134
rect 10507 3104 10577 3134
rect 11009 3104 11079 3134
rect 11511 3104 11581 3134
rect 12013 3104 12083 3134
rect 12515 3104 12585 3134
rect 13017 3104 13087 3134
rect 13519 3104 13589 3134
rect 14021 3104 14091 3134
rect 14523 3104 14593 3134
rect 15025 3104 15095 3134
rect 15527 3104 15597 3134
rect 16029 3104 16099 3134
rect 17632 3125 17650 3157
rect 17825 3125 17839 3157
rect 594 2977 624 3047
rect 882 2977 912 3047
rect 1096 2977 1126 3047
rect 1384 2977 1414 3047
rect 1598 2977 1628 3047
rect 1886 2977 1916 3047
rect 2100 2977 2130 3047
rect 2388 2977 2418 3047
rect 2602 2977 2632 3047
rect 2890 2977 2920 3047
rect 3104 2977 3134 3047
rect 3392 2977 3422 3047
rect 3606 2977 3636 3047
rect 3894 2977 3924 3047
rect 4108 2977 4138 3047
rect 4396 2977 4426 3047
rect 4610 2977 4640 3047
rect 4898 2977 4928 3047
rect 5112 2977 5142 3047
rect 5400 2977 5430 3047
rect 5614 2977 5644 3047
rect 5902 2977 5932 3047
rect 6116 2977 6146 3047
rect 6404 2977 6434 3047
rect 6618 2977 6648 3047
rect 6906 2977 6936 3047
rect 7120 2977 7150 3047
rect 7408 2977 7438 3047
rect 7622 2977 7652 3047
rect 7910 2977 7940 3047
rect 8124 2977 8154 3047
rect 8412 2977 8442 3047
rect 8626 2977 8656 3047
rect 8914 2977 8944 3047
rect 9128 2977 9158 3047
rect 9416 2977 9446 3047
rect 9630 2977 9660 3047
rect 9918 2977 9948 3047
rect 10132 2977 10162 3047
rect 10420 2977 10450 3047
rect 10634 2977 10664 3047
rect 10922 2977 10952 3047
rect 11136 2977 11166 3047
rect 11424 2977 11454 3047
rect 11638 2977 11668 3047
rect 11926 2977 11956 3047
rect 12140 2977 12170 3047
rect 12428 2977 12458 3047
rect 12642 2977 12672 3047
rect 12930 2977 12960 3047
rect 13144 2977 13174 3047
rect 13432 2977 13462 3047
rect 13646 2977 13676 3047
rect 13934 2977 13964 3047
rect 14148 2977 14178 3047
rect 14436 2977 14466 3047
rect 14650 2977 14680 3047
rect 14938 2977 14968 3047
rect 15152 2977 15182 3047
rect 15440 2977 15470 3047
rect 15654 2977 15684 3047
rect 15942 2977 15972 3047
rect 16156 2977 16186 3047
rect 16444 2977 16474 3047
rect 969 2890 1039 2920
rect 1471 2890 1541 2920
rect 1973 2890 2043 2920
rect 2475 2890 2545 2920
rect 2977 2890 3047 2920
rect 3479 2890 3549 2920
rect 3981 2890 4051 2920
rect 4483 2890 4553 2920
rect 4985 2890 5055 2920
rect 5487 2890 5557 2920
rect 5989 2890 6059 2920
rect 6491 2890 6561 2920
rect 6993 2890 7063 2920
rect 7495 2890 7565 2920
rect 7997 2890 8067 2920
rect 8499 2890 8569 2920
rect 9001 2890 9071 2920
rect 9503 2890 9573 2920
rect 10005 2890 10075 2920
rect 10507 2890 10577 2920
rect 11009 2890 11079 2920
rect 11511 2890 11581 2920
rect 12013 2890 12083 2920
rect 12515 2890 12585 2920
rect 13017 2890 13087 2920
rect 13519 2890 13589 2920
rect 14021 2890 14091 2920
rect 14523 2890 14593 2920
rect 15025 2890 15095 2920
rect 15527 2890 15597 2920
rect 16029 2890 16099 2920
rect -957 2685 -943 2717
rect -768 2685 -750 2717
rect -957 2277 -750 2685
rect 17632 2831 17839 3125
rect 17632 2816 17840 2831
rect 17632 2784 17661 2816
rect 17693 2784 17705 2816
rect 17737 2784 17749 2816
rect 17781 2784 17793 2816
rect 17825 2784 17840 2816
rect 17632 2771 17840 2784
rect 17632 2739 17661 2771
rect 17693 2739 17705 2771
rect 17737 2739 17749 2771
rect 17781 2739 17793 2771
rect 17825 2739 17840 2771
rect 17632 2726 17840 2739
rect 17632 2717 17661 2726
rect 17693 2717 17705 2726
rect 17737 2717 17749 2726
rect 17781 2717 17793 2726
rect 17632 2685 17650 2717
rect 17825 2690 17840 2726
rect 17870 2708 18077 3213
rect 20191 2946 20398 4306
rect 20151 2937 20398 2946
rect 20151 2862 20202 2937
rect 20308 2862 20398 2937
rect 20151 2855 20398 2862
rect 17825 2685 17839 2690
rect 969 2602 1039 2632
rect 1471 2602 1541 2632
rect 1973 2602 2043 2632
rect 2475 2602 2545 2632
rect 2977 2602 3047 2632
rect 3479 2602 3549 2632
rect 3981 2602 4051 2632
rect 4483 2602 4553 2632
rect 4985 2602 5055 2632
rect 5487 2602 5557 2632
rect 5989 2602 6059 2632
rect 6491 2602 6561 2632
rect 6993 2602 7063 2632
rect 7495 2602 7565 2632
rect 7997 2602 8067 2632
rect 8499 2602 8569 2632
rect 9001 2602 9071 2632
rect 9503 2602 9573 2632
rect 10005 2602 10075 2632
rect 10507 2602 10577 2632
rect 11009 2602 11079 2632
rect 11511 2602 11581 2632
rect 12013 2602 12083 2632
rect 12515 2602 12585 2632
rect 13017 2602 13087 2632
rect 13519 2602 13589 2632
rect 14021 2602 14091 2632
rect 14523 2602 14593 2632
rect 15025 2602 15095 2632
rect 15527 2602 15597 2632
rect 16029 2602 16099 2632
rect 594 2475 624 2545
rect 882 2475 912 2545
rect 1096 2475 1126 2545
rect 1384 2475 1414 2545
rect 1598 2475 1628 2545
rect 1886 2475 1916 2545
rect 2100 2475 2130 2545
rect 2388 2475 2418 2545
rect 2602 2475 2632 2545
rect 2890 2475 2920 2545
rect 3104 2475 3134 2545
rect 3392 2475 3422 2545
rect 3606 2475 3636 2545
rect 3894 2475 3924 2545
rect 4108 2475 4138 2545
rect 4396 2475 4426 2545
rect 4610 2475 4640 2545
rect 4898 2475 4928 2545
rect 5112 2475 5142 2545
rect 5400 2475 5430 2545
rect 5614 2475 5644 2545
rect 5902 2475 5932 2545
rect 6116 2475 6146 2545
rect 6404 2475 6434 2545
rect 6618 2475 6648 2545
rect 6906 2475 6936 2545
rect 7120 2475 7150 2545
rect 7408 2475 7438 2545
rect 7622 2475 7652 2545
rect 7910 2475 7940 2545
rect 8124 2475 8154 2545
rect 8412 2475 8442 2545
rect 8626 2475 8656 2545
rect 8914 2475 8944 2545
rect 9128 2475 9158 2545
rect 9416 2475 9446 2545
rect 9630 2475 9660 2545
rect 9918 2475 9948 2545
rect 10132 2475 10162 2545
rect 10420 2475 10450 2545
rect 10634 2475 10664 2545
rect 10922 2475 10952 2545
rect 11136 2475 11166 2545
rect 11424 2475 11454 2545
rect 11638 2475 11668 2545
rect 11926 2475 11956 2545
rect 12140 2475 12170 2545
rect 12428 2475 12458 2545
rect 12642 2475 12672 2545
rect 12930 2475 12960 2545
rect 13144 2475 13174 2545
rect 13432 2475 13462 2545
rect 13646 2475 13676 2545
rect 13934 2475 13964 2545
rect 14148 2475 14178 2545
rect 14436 2475 14466 2545
rect 14650 2475 14680 2545
rect 14938 2475 14968 2545
rect 15152 2475 15182 2545
rect 15440 2475 15470 2545
rect 15654 2475 15684 2545
rect 15942 2475 15972 2545
rect 16156 2475 16186 2545
rect 16444 2475 16474 2545
rect 969 2388 1039 2418
rect 1471 2388 1541 2418
rect 1973 2388 2043 2418
rect 2475 2388 2545 2418
rect 2977 2388 3047 2418
rect 3479 2388 3549 2418
rect 3981 2388 4051 2418
rect 4483 2388 4553 2418
rect 4985 2388 5055 2418
rect 5487 2388 5557 2418
rect 5989 2388 6059 2418
rect 6491 2388 6561 2418
rect 6993 2388 7063 2418
rect 7495 2388 7565 2418
rect 7997 2388 8067 2418
rect 8499 2388 8569 2418
rect 9001 2388 9071 2418
rect 9503 2388 9573 2418
rect 10005 2388 10075 2418
rect 10507 2388 10577 2418
rect 11009 2388 11079 2418
rect 11511 2388 11581 2418
rect 12013 2388 12083 2418
rect 12515 2388 12585 2418
rect 13017 2388 13087 2418
rect 13519 2388 13589 2418
rect 14021 2388 14091 2418
rect 14523 2388 14593 2418
rect 15025 2388 15095 2418
rect 15527 2388 15597 2418
rect 16029 2388 16099 2418
rect -957 2245 -943 2277
rect -768 2245 -750 2277
rect -957 1837 -750 2245
rect 969 2100 1039 2130
rect 1471 2100 1541 2130
rect 1973 2100 2043 2130
rect 2475 2100 2545 2130
rect 2977 2100 3047 2130
rect 3479 2100 3549 2130
rect 3981 2100 4051 2130
rect 4483 2100 4553 2130
rect 4985 2100 5055 2130
rect 5487 2100 5557 2130
rect 5989 2100 6059 2130
rect 6491 2100 6561 2130
rect 6993 2100 7063 2130
rect 7495 2100 7565 2130
rect 7997 2100 8067 2130
rect 8499 2100 8569 2130
rect 9001 2100 9071 2130
rect 9503 2100 9573 2130
rect 10005 2100 10075 2130
rect 10507 2100 10577 2130
rect 11009 2100 11079 2130
rect 11511 2100 11581 2130
rect 12013 2100 12083 2130
rect 12515 2100 12585 2130
rect 13017 2100 13087 2130
rect 13519 2100 13589 2130
rect 14021 2100 14091 2130
rect 14523 2100 14593 2130
rect 15025 2100 15095 2130
rect 15527 2100 15597 2130
rect 16029 2100 16099 2130
rect 594 1973 624 2043
rect 882 1973 912 2043
rect 1096 1973 1126 2043
rect 1384 1973 1414 2043
rect 1598 1973 1628 2043
rect 1886 1973 1916 2043
rect 2100 1973 2130 2043
rect 2388 1973 2418 2043
rect 2602 1973 2632 2043
rect 2890 1973 2920 2043
rect 3104 1973 3134 2043
rect 3392 1973 3422 2043
rect 3606 1973 3636 2043
rect 3894 1973 3924 2043
rect 4108 1973 4138 2043
rect 4396 1973 4426 2043
rect 4610 1973 4640 2043
rect 4898 1973 4928 2043
rect 5112 1973 5142 2043
rect 5400 1973 5430 2043
rect 5614 1973 5644 2043
rect 5902 1973 5932 2043
rect 6116 1973 6146 2043
rect 6404 1973 6434 2043
rect 6618 1973 6648 2043
rect 6906 1973 6936 2043
rect 7120 1973 7150 2043
rect 7408 1973 7438 2043
rect 7622 1973 7652 2043
rect 7910 1973 7940 2043
rect 8124 1973 8154 2043
rect 8412 1973 8442 2043
rect 8626 1973 8656 2043
rect 8914 1973 8944 2043
rect 9128 1973 9158 2043
rect 9416 1973 9446 2043
rect 9630 1973 9660 2043
rect 9918 1973 9948 2043
rect 10132 1973 10162 2043
rect 10420 1973 10450 2043
rect 10634 1973 10664 2043
rect 10922 1973 10952 2043
rect 11136 1973 11166 2043
rect 11424 1973 11454 2043
rect 11638 1973 11668 2043
rect 11926 1973 11956 2043
rect 12140 1973 12170 2043
rect 12428 1973 12458 2043
rect 12642 1973 12672 2043
rect 12930 1973 12960 2043
rect 13144 1973 13174 2043
rect 13432 1973 13462 2043
rect 13646 1973 13676 2043
rect 13934 1973 13964 2043
rect 14148 1973 14178 2043
rect 14436 1973 14466 2043
rect 14650 1973 14680 2043
rect 14938 1973 14968 2043
rect 15152 1973 15182 2043
rect 15440 1973 15470 2043
rect 15654 1973 15684 2043
rect 15942 1973 15972 2043
rect 16156 1973 16186 2043
rect 16444 1973 16474 2043
rect 969 1886 1039 1916
rect 1471 1886 1541 1916
rect 1973 1886 2043 1916
rect 2475 1886 2545 1916
rect 2977 1886 3047 1916
rect 3479 1886 3549 1916
rect 3981 1886 4051 1916
rect 4483 1886 4553 1916
rect 4985 1886 5055 1916
rect 5487 1886 5557 1916
rect 5989 1886 6059 1916
rect 6491 1886 6561 1916
rect 6993 1886 7063 1916
rect 7495 1886 7565 1916
rect 7997 1886 8067 1916
rect 8499 1886 8569 1916
rect 9001 1886 9071 1916
rect 9503 1886 9573 1916
rect 10005 1886 10075 1916
rect 10507 1886 10577 1916
rect 11009 1886 11079 1916
rect 11511 1886 11581 1916
rect 12013 1886 12083 1916
rect 12515 1886 12585 1916
rect 13017 1886 13087 1916
rect 13519 1886 13589 1916
rect 14021 1886 14091 1916
rect 14523 1886 14593 1916
rect 15025 1886 15095 1916
rect 15527 1886 15597 1916
rect 16029 1886 16099 1916
rect -957 1805 -943 1837
rect -768 1805 -750 1837
rect -957 1397 -750 1805
rect 17632 1837 17839 2685
rect 17632 1805 17650 1837
rect 17632 1787 17661 1805
rect 17693 1787 17705 1805
rect 17737 1787 17749 1805
rect 17781 1787 17793 1805
rect 17825 1787 17839 1837
rect 17632 1774 17839 1787
rect 17632 1742 17661 1774
rect 17693 1742 17705 1774
rect 17737 1742 17749 1774
rect 17781 1742 17793 1774
rect 17825 1742 17839 1774
rect 17632 1729 17839 1742
rect 17632 1697 17661 1729
rect 17693 1697 17705 1729
rect 17737 1697 17749 1729
rect 17781 1697 17793 1729
rect 17825 1697 17839 1729
rect 969 1598 1039 1628
rect 1471 1598 1541 1628
rect 1973 1598 2043 1628
rect 2475 1598 2545 1628
rect 2977 1598 3047 1628
rect 3479 1598 3549 1628
rect 3981 1598 4051 1628
rect 4483 1598 4553 1628
rect 4985 1598 5055 1628
rect 5487 1598 5557 1628
rect 5989 1598 6059 1628
rect 6491 1598 6561 1628
rect 6993 1598 7063 1628
rect 7495 1598 7565 1628
rect 7997 1598 8067 1628
rect 8499 1598 8569 1628
rect 9001 1598 9071 1628
rect 9503 1598 9573 1628
rect 10005 1598 10075 1628
rect 10507 1598 10577 1628
rect 11009 1598 11079 1628
rect 11511 1598 11581 1628
rect 12013 1598 12083 1628
rect 12515 1598 12585 1628
rect 13017 1598 13087 1628
rect 13519 1598 13589 1628
rect 14021 1598 14091 1628
rect 14523 1598 14593 1628
rect 15025 1598 15095 1628
rect 15527 1598 15597 1628
rect 16029 1598 16099 1628
rect 594 1471 624 1541
rect 882 1471 912 1541
rect 1096 1471 1126 1541
rect 1384 1471 1414 1541
rect 1598 1471 1628 1541
rect 1886 1471 1916 1541
rect 2100 1471 2130 1541
rect 2388 1471 2418 1541
rect 2602 1471 2632 1541
rect 2890 1471 2920 1541
rect 3104 1471 3134 1541
rect 3392 1471 3422 1541
rect 3606 1471 3636 1541
rect 3894 1471 3924 1541
rect 4108 1471 4138 1541
rect 4396 1471 4426 1541
rect 4610 1471 4640 1541
rect 4898 1471 4928 1541
rect 5112 1471 5142 1541
rect 5400 1471 5430 1541
rect 5614 1471 5644 1541
rect 5902 1471 5932 1541
rect 6116 1471 6146 1541
rect 6404 1471 6434 1541
rect 6618 1471 6648 1541
rect 6906 1471 6936 1541
rect 7120 1471 7150 1541
rect 7408 1471 7438 1541
rect 7622 1471 7652 1541
rect 7910 1471 7940 1541
rect 8124 1471 8154 1541
rect 8412 1471 8442 1541
rect 8626 1471 8656 1541
rect 8914 1471 8944 1541
rect 9128 1471 9158 1541
rect 9416 1471 9446 1541
rect 9630 1471 9660 1541
rect 9918 1471 9948 1541
rect 10132 1471 10162 1541
rect 10420 1471 10450 1541
rect 10634 1471 10664 1541
rect 10922 1471 10952 1541
rect 11136 1471 11166 1541
rect 11424 1471 11454 1541
rect 11638 1471 11668 1541
rect 11926 1471 11956 1541
rect 12140 1471 12170 1541
rect 12428 1471 12458 1541
rect 12642 1471 12672 1541
rect 12930 1471 12960 1541
rect 13144 1471 13174 1541
rect 13432 1471 13462 1541
rect 13646 1471 13676 1541
rect 13934 1471 13964 1541
rect 14148 1471 14178 1541
rect 14436 1471 14466 1541
rect 14650 1471 14680 1541
rect 14938 1471 14968 1541
rect 15152 1471 15182 1541
rect 15440 1471 15470 1541
rect 15654 1471 15684 1541
rect 15942 1471 15972 1541
rect 16156 1471 16186 1541
rect 16444 1471 16474 1541
rect -957 1365 -943 1397
rect -768 1365 -750 1397
rect 969 1384 1039 1414
rect 1471 1384 1541 1414
rect 1973 1384 2043 1414
rect 2475 1384 2545 1414
rect 2977 1384 3047 1414
rect 3479 1384 3549 1414
rect 3981 1384 4051 1414
rect 4483 1384 4553 1414
rect 4985 1384 5055 1414
rect 5487 1384 5557 1414
rect 5989 1384 6059 1414
rect 6491 1384 6561 1414
rect 6993 1384 7063 1414
rect 7495 1384 7565 1414
rect 7997 1384 8067 1414
rect 8499 1384 8569 1414
rect 9001 1384 9071 1414
rect 9503 1384 9573 1414
rect 10005 1384 10075 1414
rect 10507 1384 10577 1414
rect 11009 1384 11079 1414
rect 11511 1384 11581 1414
rect 12013 1384 12083 1414
rect 12515 1384 12585 1414
rect 13017 1384 13087 1414
rect 13519 1384 13589 1414
rect 14021 1384 14091 1414
rect 14523 1384 14593 1414
rect 15025 1384 15095 1414
rect 15527 1384 15597 1414
rect 16029 1384 16099 1414
rect 17632 1397 17839 1697
rect -957 957 -750 1365
rect 17632 1365 17650 1397
rect 17825 1365 17839 1397
rect 969 1096 1039 1126
rect 1471 1096 1541 1126
rect 1973 1096 2043 1126
rect 2475 1096 2545 1126
rect 2977 1096 3047 1126
rect 3479 1096 3549 1126
rect 3981 1096 4051 1126
rect 4483 1096 4553 1126
rect 4985 1096 5055 1126
rect 5487 1096 5557 1126
rect 5989 1096 6059 1126
rect 6491 1096 6561 1126
rect 6993 1096 7063 1126
rect 7495 1096 7565 1126
rect 7997 1096 8067 1126
rect 8499 1096 8569 1126
rect 9001 1096 9071 1126
rect 9503 1096 9573 1126
rect 10005 1096 10075 1126
rect 10507 1096 10577 1126
rect 11009 1096 11079 1126
rect 11511 1096 11581 1126
rect 12013 1096 12083 1126
rect 12515 1096 12585 1126
rect 13017 1096 13087 1126
rect 13519 1096 13589 1126
rect 14021 1096 14091 1126
rect 14523 1096 14593 1126
rect 15025 1096 15095 1126
rect 15527 1096 15597 1126
rect 16029 1096 16099 1126
rect 594 969 624 1039
rect 882 969 912 1039
rect 1096 969 1126 1039
rect 1384 969 1414 1039
rect 1598 969 1628 1039
rect 1886 969 1916 1039
rect 2100 969 2130 1039
rect 2388 969 2418 1039
rect 2602 969 2632 1039
rect 2890 969 2920 1039
rect 3104 969 3134 1039
rect 3392 969 3422 1039
rect 3606 969 3636 1039
rect 3894 969 3924 1039
rect 4108 969 4138 1039
rect 4396 969 4426 1039
rect 4610 969 4640 1039
rect 4898 969 4928 1039
rect 5112 969 5142 1039
rect 5400 969 5430 1039
rect 5614 969 5644 1039
rect 5902 969 5932 1039
rect 6116 969 6146 1039
rect 6404 969 6434 1039
rect 6618 969 6648 1039
rect 6906 969 6936 1039
rect 7120 969 7150 1039
rect 7408 969 7438 1039
rect 7622 969 7652 1039
rect 7910 969 7940 1039
rect 8124 969 8154 1039
rect 8412 969 8442 1039
rect 8626 969 8656 1039
rect 8914 969 8944 1039
rect 9128 969 9158 1039
rect 9416 969 9446 1039
rect 9630 969 9660 1039
rect 9918 969 9948 1039
rect 10132 969 10162 1039
rect 10420 969 10450 1039
rect 10634 969 10664 1039
rect 10922 969 10952 1039
rect 11136 969 11166 1039
rect 11424 969 11454 1039
rect 11638 969 11668 1039
rect 11926 969 11956 1039
rect 12140 969 12170 1039
rect 12428 969 12458 1039
rect 12642 969 12672 1039
rect 12930 969 12960 1039
rect 13144 969 13174 1039
rect 13432 969 13462 1039
rect 13646 969 13676 1039
rect 13934 969 13964 1039
rect 14148 969 14178 1039
rect 14436 969 14466 1039
rect 14650 969 14680 1039
rect 14938 969 14968 1039
rect 15152 969 15182 1039
rect 15440 969 15470 1039
rect 15654 969 15684 1039
rect 15942 969 15972 1039
rect 16156 969 16186 1039
rect 16444 969 16474 1039
rect -957 925 -943 957
rect -768 925 -750 957
rect -957 517 -750 925
rect 17632 957 17839 1365
rect 17632 925 17650 957
rect 17825 925 17839 957
rect 969 882 1039 912
rect 1471 882 1541 912
rect 1973 882 2043 912
rect 2475 882 2545 912
rect 2977 882 3047 912
rect 3479 882 3549 912
rect 3981 882 4051 912
rect 4483 882 4553 912
rect 4985 882 5055 912
rect 5487 882 5557 912
rect 5989 882 6059 912
rect 6491 882 6561 912
rect 6993 882 7063 912
rect 7495 882 7565 912
rect 7997 882 8067 912
rect 8499 882 8569 912
rect 9001 882 9071 912
rect 9503 882 9573 912
rect 10005 882 10075 912
rect 10507 882 10577 912
rect 11009 882 11079 912
rect 11511 882 11581 912
rect 12013 882 12083 912
rect 12515 882 12585 912
rect 13017 882 13087 912
rect 13519 882 13589 912
rect 14021 882 14091 912
rect 14523 882 14593 912
rect 15025 882 15095 912
rect 15527 882 15597 912
rect 16029 882 16099 912
rect 17632 834 17839 925
rect 17631 819 17839 834
rect 17631 787 17659 819
rect 17691 787 17703 819
rect 17735 787 17747 819
rect 17779 787 17791 819
rect 17823 787 17839 819
rect 17631 774 17839 787
rect 17631 742 17659 774
rect 17691 742 17703 774
rect 17735 742 17747 774
rect 17779 742 17791 774
rect 17823 742 17839 774
rect 17631 729 17839 742
rect 17631 697 17659 729
rect 17691 697 17703 729
rect 17735 697 17747 729
rect 17779 697 17791 729
rect 17823 697 17839 729
rect 17631 693 17839 697
rect 969 594 1039 624
rect 1471 594 1541 624
rect 1973 594 2043 624
rect 2475 594 2545 624
rect 2977 594 3047 624
rect 3479 594 3549 624
rect 3981 594 4051 624
rect 4483 594 4553 624
rect 4985 594 5055 624
rect 5487 594 5557 624
rect 5989 594 6059 624
rect 6491 594 6561 624
rect 6993 594 7063 624
rect 7495 594 7565 624
rect 7997 594 8067 624
rect 8499 594 8569 624
rect 9001 594 9071 624
rect 9503 594 9573 624
rect 10005 594 10075 624
rect 10507 594 10577 624
rect 11009 594 11079 624
rect 11511 594 11581 624
rect 12013 594 12083 624
rect 12515 594 12585 624
rect 13017 594 13087 624
rect 13519 594 13589 624
rect 14021 594 14091 624
rect 14523 594 14593 624
rect 15025 594 15095 624
rect 15527 594 15597 624
rect 16029 594 16099 624
rect -957 485 -943 517
rect -768 485 -750 517
rect -957 77 -750 485
rect 4610 467 4640 537
rect 4898 467 4928 537
rect 6762 467 6792 537
rect 8626 467 8656 537
rect 8770 467 8800 537
rect 12642 467 12672 537
rect 14292 467 14322 537
rect 17632 517 17839 693
rect 17632 485 17650 517
rect 17825 485 17839 517
rect 4518 380 4553 410
rect 4985 380 5020 410
rect -957 45 -943 77
rect -768 45 -750 77
rect -957 -91 -750 45
rect 17632 77 17839 485
rect 17632 45 17650 77
rect 17825 45 17839 77
rect -957 -123 -942 -91
rect -910 -123 -898 -91
rect -866 -123 -854 -91
rect -822 -123 -810 -91
rect -778 -123 -750 -91
rect -957 -136 -750 -123
rect -957 -168 -942 -136
rect -910 -168 -898 -136
rect -866 -168 -854 -136
rect -822 -168 -810 -136
rect -778 -168 -750 -136
rect -957 -181 -750 -168
rect -957 -213 -942 -181
rect -910 -213 -898 -181
rect -866 -213 -854 -181
rect -822 -213 -810 -181
rect -778 -213 -750 -181
rect -957 -217 -750 -213
rect -1195 -342 -1180 -310
rect -1148 -342 -1136 -310
rect -1104 -342 -1092 -310
rect -1060 -342 -1048 -310
rect -1016 -342 -988 -310
rect -1195 -355 -988 -342
rect -1195 -387 -1180 -355
rect -1148 -387 -1136 -355
rect -1104 -387 -1092 -355
rect -1060 -387 -1048 -355
rect -1016 -387 -988 -355
rect -1195 -400 -988 -387
rect -1195 -432 -1180 -400
rect -1148 -432 -1136 -400
rect -1104 -432 -1092 -400
rect -1060 -432 -1048 -400
rect -1016 -432 -988 -400
rect -1195 -436 -988 -432
rect 16300 -456 16330 0
rect 17632 -26 17839 45
rect 17632 -58 17660 -26
rect 17692 -58 17704 -26
rect 17736 -58 17748 -26
rect 17780 -58 17792 -26
rect 17824 -58 17839 -26
rect 17632 -71 17839 -58
rect 17632 -103 17660 -71
rect 17692 -103 17704 -71
rect 17736 -103 17748 -71
rect 17780 -103 17792 -71
rect 17824 -103 17839 -71
rect 17632 -116 17839 -103
rect 17632 -148 17660 -116
rect 17692 -148 17704 -116
rect 17736 -148 17748 -116
rect 17780 -148 17792 -116
rect 17824 -148 17839 -116
rect 17632 -371 17839 -148
rect 17870 2536 18151 2708
rect 20191 2675 20398 2855
rect 20151 2666 20398 2675
rect 20151 2591 20202 2666
rect 20308 2591 20398 2666
rect 20151 2584 20398 2591
rect 17870 2305 18077 2536
rect 20191 2397 20398 2584
rect 20151 2388 20398 2397
rect 20151 2313 20202 2388
rect 20308 2313 20398 2388
rect 20151 2306 20398 2313
rect 17870 2273 17898 2305
rect 17930 2273 17942 2305
rect 17974 2273 17986 2305
rect 18018 2273 18030 2305
rect 18062 2273 18077 2305
rect 17870 2260 18077 2273
rect 17870 2228 17898 2260
rect 17930 2228 17942 2260
rect 17974 2228 17986 2260
rect 18018 2228 18030 2260
rect 18062 2228 18077 2260
rect 17870 2215 18077 2228
rect 17870 2183 17898 2215
rect 17930 2183 17942 2215
rect 17974 2183 17986 2215
rect 18018 2183 18030 2215
rect 18062 2183 18077 2215
rect 17870 1303 18077 2183
rect 17870 1271 17898 1303
rect 17930 1271 17942 1303
rect 17974 1271 17986 1303
rect 18018 1271 18030 1303
rect 18062 1271 18077 1303
rect 17870 1258 18077 1271
rect 17870 1226 17898 1258
rect 17930 1226 17942 1258
rect 17974 1226 17986 1258
rect 18018 1226 18030 1258
rect 18062 1226 18077 1258
rect 17870 1213 18077 1226
rect 17870 1181 17898 1213
rect 17930 1181 17942 1213
rect 17974 1181 17986 1213
rect 18018 1181 18030 1213
rect 18062 1181 18077 1213
rect 17870 711 18077 1181
rect 20191 946 20398 2306
rect 20151 937 20398 946
rect 20151 862 20202 937
rect 20308 862 20398 937
rect 20151 855 20398 862
rect 17870 539 18151 711
rect 20191 675 20398 855
rect 20151 666 20398 675
rect 20151 591 20202 666
rect 20308 591 20398 666
rect 20151 584 20398 591
rect 17870 306 18077 539
rect 20191 397 20398 584
rect 20151 388 20398 397
rect 20151 313 20202 388
rect 20308 313 20398 388
rect 20151 306 20398 313
rect 17870 274 17898 306
rect 17930 274 17942 306
rect 17974 274 17986 306
rect 18018 274 18030 306
rect 18062 274 18077 306
rect 17870 261 18077 274
rect 17870 229 17898 261
rect 17930 229 17942 261
rect 17974 229 17986 261
rect 18018 229 18030 261
rect 18062 229 18077 261
rect 17870 216 18077 229
rect 17870 184 17898 216
rect 17930 184 17942 216
rect 17974 184 17986 216
rect 18018 184 18030 216
rect 18062 184 18077 216
rect 17870 -245 18077 184
rect 17870 -277 17898 -245
rect 17930 -277 17942 -245
rect 17974 -277 17986 -245
rect 18018 -277 18030 -245
rect 18062 -277 18077 -245
rect 17870 -290 18077 -277
rect 17870 -322 17898 -290
rect 17930 -322 17942 -290
rect 17974 -322 17986 -290
rect 18018 -322 18030 -290
rect 18062 -322 18077 -290
rect 17870 -335 18077 -322
rect 17870 -367 17898 -335
rect 17930 -367 17942 -335
rect 17974 -367 17986 -335
rect 18018 -367 18030 -335
rect 18062 -367 18077 -335
rect 17870 -371 18077 -367
rect 20191 -374 20398 306
rect 20435 11371 20642 11627
rect 20435 11290 20442 11371
rect 20561 11290 20642 11371
rect 20435 11168 20642 11290
rect 20435 10962 20448 11168
rect 20554 10962 20642 11168
rect 20435 10289 20642 10962
rect 20435 10083 20448 10289
rect 20554 10083 20642 10289
rect 20435 9816 20642 10083
rect 20435 9735 20442 9816
rect 20561 9735 20642 9816
rect 20435 9371 20642 9735
rect 20435 9290 20442 9371
rect 20561 9290 20642 9371
rect 20435 9168 20642 9290
rect 20435 8962 20448 9168
rect 20554 8962 20642 9168
rect 20435 8289 20642 8962
rect 20435 8083 20448 8289
rect 20554 8083 20642 8289
rect 20435 7816 20642 8083
rect 20435 7735 20442 7816
rect 20561 7735 20642 7816
rect 20435 7371 20642 7735
rect 20435 7290 20442 7371
rect 20561 7290 20642 7371
rect 20435 7168 20642 7290
rect 20435 6962 20448 7168
rect 20554 6962 20642 7168
rect 20435 6289 20642 6962
rect 20435 6083 20448 6289
rect 20554 6083 20642 6289
rect 20435 5816 20642 6083
rect 20435 5735 20442 5816
rect 20561 5735 20642 5816
rect 20435 5371 20642 5735
rect 20435 5290 20442 5371
rect 20561 5290 20642 5371
rect 20435 5168 20642 5290
rect 20435 4962 20448 5168
rect 20554 4962 20642 5168
rect 20435 4289 20642 4962
rect 20435 4083 20448 4289
rect 20554 4083 20642 4289
rect 20435 3816 20642 4083
rect 20435 3735 20442 3816
rect 20561 3735 20642 3816
rect 20435 3371 20642 3735
rect 20435 3290 20442 3371
rect 20561 3290 20642 3371
rect 20435 3168 20642 3290
rect 20435 2962 20448 3168
rect 20554 2962 20642 3168
rect 20435 2289 20642 2962
rect 20435 2083 20448 2289
rect 20554 2083 20642 2289
rect 20435 1816 20642 2083
rect 20435 1735 20442 1816
rect 20561 1735 20642 1816
rect 20435 1371 20642 1735
rect 20435 1290 20442 1371
rect 20561 1290 20642 1371
rect 20435 1168 20642 1290
rect 20435 962 20448 1168
rect 20554 962 20642 1168
rect 20435 289 20642 962
rect 20435 83 20448 289
rect 20554 83 20642 289
rect 20435 -184 20642 83
rect 20435 -265 20442 -184
rect 20561 -265 20642 -184
rect 20435 -373 20642 -265
use adc_array_wafflecap_8_1  adc_array_wafflecap_8_1_0 ../adc_array_cap
timestamp 1662987872
transform 1 0 12550 0 1 0
box 0 0 502 502
use adc_array_wafflecap_8_2  adc_array_wafflecap_8_2_0 ../adc_array_cap
timestamp 1662983799
transform 1 0 8534 0 1 0
box 0 0 502 502
use adc_array_wafflecap_8_4  adc_array_wafflecap_8_4_0 ../adc_array_cap
timestamp 1662985026
transform 1 0 4518 0 1 0
box 0 0 502 502
use adc_array_wafflecap_8_8  adc_array_wafflecap_8_8_0 ../adc_array_cap
array 0 31 502 0 15 502
timestamp 1662984960
transform 1 0 502 0 1 502
box 0 0 502 502
use adc_array_wafflecap_8_Drv  adc_array_wafflecap_8_Drv_0 ../adc_array_cap
array 0 0 502 0 15 502
timestamp 1663255439
transform 1 0 0 0 1 502
box 0 0 502 502
use adc_array_wafflecap_8_Dummy  adc_array_wafflecap_8_Dummy_0 ../adc_array_cap
array 0 8 502 0 0 502
timestamp 1663073688
transform 1 0 0 0 1 0
box 0 0 502 502
use adc_array_wafflecap_8_Dummy  adc_array_wafflecap_8_Dummy_1
array 0 6 502 0 0 502
timestamp 1663073688
transform 1 0 5020 0 1 0
box 0 0 502 502
use adc_array_wafflecap_8_Dummy  adc_array_wafflecap_8_Dummy_2
array 0 6 502 0 0 502
timestamp 1663073688
transform 1 0 9036 0 1 0
box 0 0 502 502
use adc_array_wafflecap_8_Dummy  adc_array_wafflecap_8_Dummy_3
array 0 5 502 0 0 502
timestamp 1663073688
transform 1 0 13052 0 1 0
box 0 0 502 502
use adc_array_wafflecap_8_Dummy  adc_array_wafflecap_8_Dummy_4
array 0 33 502 0 0 502
timestamp 1663073688
transform 1 0 0 0 1 8534
box 0 0 502 502
use adc_array_wafflecap_8_Dummy  adc_array_wafflecap_8_Dummy_5
array 0 0 502 0 15 502
timestamp 1663073688
transform 1 0 16566 0 1 502
box 0 0 502 502
use adc_array_wafflecap_8_Dummy  adc_array_wafflecap_8_Dummy_6
timestamp 1663073688
transform 1 0 16566 0 1 0
box 0 0 502 502
use adc_array_wafflecap_8_Gate  adc_array_wafflecap_8_Gate_0 ../adc_array_cap
timestamp 1663061126
transform 1 0 16064 0 1 0
box 0 0 502 502
use adc_noise_decoup_cell1  adc_noise_decoup_cell1_0 ../adc_noise_decoup_cell
array 0 0 2000 0 5 2000
timestamp 1663254830
transform 1 0 18151 0 1 -374
box 0 0 2000 2000
use adc_noise_decoup_cell1  adc_noise_decoup_cell1_1
array 0 8 2000 0 0 2000
timestamp 1663254830
transform 1 0 151 0 1 9626
box 0 0 2000 2000
<< labels >>
flabel locali s -659 -457 -625 -436 5 FreeSans 40 0 0 0 sample_n
port 44 s
flabel locali s -605 -457 -571 -436 5 FreeSans 40 0 0 0 sample
port 45 s
flabel locali s -551 -457 -483 -436 5 FreeSans 40 0 0 0 vcom
port 46 s
flabel locali s -440 -457 -294 -436 5 FreeSans 40 0 0 0 VDD
port 61 s
flabel locali s -251 -457 -105 -436 5 FreeSans 40 0 0 0 VSS
port 62 s
flabel locali s 929 -457 946 -436 5 FreeSans 80 0 0 0 row_n[0]
port 70 s
flabel locali s 1431 -457 1448 -436 5 FreeSans 80 0 0 0 row_n[1]
port 71 s
flabel locali s 1933 -457 1950 -436 5 FreeSans 80 0 0 0 row_n[2]
port 72 s
flabel locali s 2435 -457 2452 -436 5 FreeSans 80 0 0 0 row_n[3]
port 73 s
flabel locali s 2937 -457 2954 -436 5 FreeSans 80 0 0 0 row_n[4]
port 74 s
flabel locali s 3439 -457 3456 -436 5 FreeSans 80 0 0 0 row_n[5]
port 75 s
flabel locali s 3941 -457 3958 -436 5 FreeSans 80 0 0 0 row_n[6]
port 76 s
flabel locali s 4443 -457 4460 -436 5 FreeSans 80 0 0 0 row_n[7]
port 77 s
flabel locali s 4945 -457 4962 -436 5 FreeSans 80 0 0 0 row_n[8]
port 78 s
flabel locali s 5447 -457 5464 -436 5 FreeSans 80 0 0 0 row_n[9]
port 79 s
flabel locali s 5949 -457 5966 -436 5 FreeSans 80 0 0 0 row_n[10]
port 80 s
flabel locali s 6451 -457 6468 -436 5 FreeSans 80 0 0 0 row_n[11]
port 81 s
flabel locali s 6953 -457 6970 -436 5 FreeSans 80 0 0 0 row_n[12]
port 82 s
flabel locali s 7455 -457 7472 -436 5 FreeSans 80 0 0 0 row_n[13]
port 83 s
flabel locali s 7957 -457 7974 -436 5 FreeSans 80 0 0 0 row_n[14]
port 84 s
flabel locali s 8459 -457 8476 -436 5 FreeSans 80 0 0 0 row_n[15]
port 85 s
flabel locali s 8961 -457 8978 -436 5 FreeSans 80 0 0 0 row_n[16]
port 86 s
flabel locali s 9463 -457 9480 -436 5 FreeSans 80 0 0 0 row_n[17]
port 87 s
flabel locali s 9965 -457 9982 -436 5 FreeSans 80 0 0 0 row_n[18]
port 88 s
flabel locali s 10467 -457 10484 -436 5 FreeSans 80 0 0 0 row_n[19]
port 89 s
flabel locali s 10969 -457 10986 -436 5 FreeSans 80 0 0 0 row_n[20]
port 90 s
flabel locali s 11471 -457 11488 -436 5 FreeSans 80 0 0 0 row_n[21]
port 91 s
flabel locali s 11973 -457 11990 -436 5 FreeSans 80 0 0 0 row_n[22]
port 92 s
flabel locali s 12475 -457 12492 -436 5 FreeSans 80 0 0 0 row_n[23]
port 93 s
flabel locali s 12977 -457 12994 -436 5 FreeSans 80 0 0 0 row_n[24]
port 94 s
flabel locali s 4779 -457 4796 -436 5 FreeSans 80 0 0 0 en_n_bit[2]
port 102 s
flabel locali s 8795 -457 8812 -436 5 FreeSans 80 0 0 0 en_n_bit[1]
port 103 s
flabel locali s 12811 -457 12828 -436 5 FreeSans 80 0 0 0 en_n_bit[0]
port 104 s
flabel locali s 13079 -457 13096 -436 5 FreeSans 80 0 0 0 row_n[25]
port 95 s
flabel locali s 13181 -457 13198 -436 5 FreeSans 80 0 0 0 row_n[26]
port 96 s
flabel locali s 13283 -457 13300 -436 5 FreeSans 80 0 0 0 row_n[27]
port 97 s
flabel locali s 13385 -457 13402 -436 5 FreeSans 80 0 0 0 row_n[28]
port 98 s
flabel locali s 13487 -457 13504 -436 5 FreeSans 80 0 0 0 row_n[29]
port 99 s
flabel locali s 13589 -457 13606 -436 5 FreeSans 80 0 0 0 row_n[30]
port 100 s
flabel locali s 13691 -457 13708 -436 5 FreeSans 80 0 0 0 row_n[31]
port 101 s
flabel locali s 16043 -456 16060 -435 5 FreeSans 80 90 0 0 sw_n
port 110 s
flabel locali s 16104 -456 16121 -435 5 FreeSans 80 90 0 0 sw
port 111 s
flabel metal4 s 16300 -456 16330 -427 5 FreeSans 80 0 0 0 ctop
port 115 s
flabel locali s 17167 -392 17315 -370 0 FreeSans 160 0 0 0 VSS
port 62 nsew
flabel locali s 17355 -392 17503 -370 0 FreeSans 160 0 0 0 VDD
port 61 nsew
flabel metal1 s 18102 -453 18196 -429 0 FreeSans 80 0 0 0 analog_in
port 122 nsew
flabel metal4 s -957 -217 -750 9494 0 FreeSans 800 90 0 0 VSS
port 62 nsew
flabel metal4 s -1195 -436 -988 9494 0 FreeSans 800 90 0 0 VDD
port 61 nsew
flabel metal1 s -673 717 -620 731 7 FreeSans 80 0 0 0 col_n[0]
port 123 w
flabel metal1 s -673 1219 -620 1233 7 FreeSans 80 0 0 0 col_n[1]
port 124 w
flabel metal1 s -673 1721 -620 1735 7 FreeSans 80 0 0 0 col_n[2]
port 125 w
flabel metal1 s -673 2223 -620 2237 7 FreeSans 80 0 0 0 col_n[3]
port 126 w
flabel metal1 s -673 2725 -620 2739 7 FreeSans 80 0 0 0 col_n[4]
port 127 w
flabel metal1 s -673 3227 -620 3241 7 FreeSans 80 0 0 0 col_n[5]
port 128 w
flabel metal1 s -673 3729 -620 3743 7 FreeSans 80 0 0 0 col_n[6]
port 129 w
flabel metal1 s -673 4231 -620 4245 7 FreeSans 80 0 0 0 col_n[7]
port 130 w
flabel metal1 s -673 4733 -620 4747 7 FreeSans 80 0 0 0 col_n[8]
port 131 w
flabel metal1 s -673 5235 -620 5249 7 FreeSans 80 0 0 0 col_n[9]
port 132 w
flabel metal1 s -673 5737 -620 5751 7 FreeSans 80 0 0 0 col_n[10]
port 133 w
flabel metal1 s -673 6239 -620 6253 7 FreeSans 80 0 0 0 col_n[11]
port 134 w
flabel metal1 s -673 6741 -620 6755 7 FreeSans 80 0 0 0 col_n[12]
port 135 w
flabel metal1 s -673 7243 -620 7257 7 FreeSans 80 0 0 0 col_n[13]
port 136 w
flabel metal1 s -673 7745 -620 7759 7 FreeSans 80 0 0 0 col_n[14]
port 137 w
flabel metal1 s -673 8247 -620 8261 7 FreeSans 80 0 0 0 col_n[15]
port 138 w
flabel metal1 s -673 758 -620 772 7 FreeSans 80 0 0 0 colon_n[0]
port 139 w
flabel metal1 s -673 1260 -620 1274 7 FreeSans 80 0 0 0 colon_n[1]
port 140 w
flabel metal1 s -673 1762 -620 1776 7 FreeSans 80 0 0 0 colon_n[2]
port 141 w
flabel metal1 s -673 2264 -620 2278 7 FreeSans 80 0 0 0 colon_n[3]
port 142 w
flabel metal1 s -674 2766 -621 2780 7 FreeSans 80 0 0 0 colon_n[4]
port 143 w
flabel metal1 s -673 3268 -620 3282 7 FreeSans 80 0 0 0 colon_n[5]
port 144 w
flabel metal1 s -673 3770 -620 3784 7 FreeSans 80 0 0 0 colon_n[6]
port 145 w
flabel metal1 s -673 4272 -620 4286 7 FreeSans 80 0 0 0 colon_n[7]
port 146 w
flabel metal1 s -673 4774 -620 4788 7 FreeSans 80 0 0 0 colon_n[8]
port 147 w
flabel metal1 s -673 5276 -620 5290 7 FreeSans 80 0 0 0 colon_n[9]
port 148 w
flabel metal1 s -673 5778 -620 5792 7 FreeSans 80 0 0 0 colon_n[10]
port 149 w
flabel metal1 s -673 6280 -620 6294 7 FreeSans 80 0 0 0 colon_n[11]
port 150 w
flabel metal1 s -673 6782 -620 6796 7 FreeSans 80 0 0 0 colon_n[12]
port 151 w
flabel metal1 s -673 7284 -620 7298 7 FreeSans 80 0 0 0 colon_n[13]
port 152 w
flabel metal1 s -673 7786 -620 7800 7 FreeSans 80 0 0 0 colon_n[14]
port 153 w
flabel metal1 s -673 8288 -620 8302 7 FreeSans 80 0 0 0 colon_n[15]
port 154 w
flabel metal4 s 17870 -371 18077 9495 0 FreeSans 800 90 0 0 VDD
port 117 nsew
flabel metal4 s 17632 -152 17839 9494 0 FreeSans 800 90 0 0 VSS
port 119 nsew
flabel metal4 s 20191 -374 20398 11626 0 FreeSans 800 90 0 0 VDD
port 158 nsew
flabel metal4 s 20435 -373 20642 11627 0 FreeSans 800 90 0 0 VSS
port 160 nsew
<< end >>
