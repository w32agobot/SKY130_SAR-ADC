magic
tech sky130A
timestamp 1660635965
<< checkpaint >>
rect -632 -690 1099 1040
<< metal2 >>
rect 42 306 412 351
rect 42 278 87 306
rect 115 278 173 306
rect 201 278 259 306
rect 287 278 345 306
rect 373 278 412 306
rect 42 220 412 278
rect 42 192 87 220
rect 115 192 173 220
rect 201 192 259 220
rect 287 192 345 220
rect 373 192 412 220
rect 42 134 412 192
rect 42 106 87 134
rect 115 106 173 134
rect 201 106 259 134
rect 287 106 345 134
rect 373 106 412 134
rect 42 48 412 106
rect 42 20 87 48
rect 115 20 173 48
rect 201 20 259 48
rect 287 20 345 48
rect 373 20 412 48
rect 42 -19 412 20
<< via2 >>
rect 87 278 115 306
rect 173 278 201 306
rect 259 278 287 306
rect 345 278 373 306
rect 87 192 115 220
rect 173 192 201 220
rect 259 192 287 220
rect 345 192 373 220
rect 87 106 115 134
rect 173 106 201 134
rect 259 106 287 134
rect 345 106 373 134
rect 87 20 115 48
rect 173 20 201 48
rect 259 20 287 48
rect 345 20 373 48
<< metal3 >>
rect 50 306 404 309
rect 50 278 87 306
rect 115 278 173 306
rect 201 278 259 306
rect 287 278 345 306
rect 373 278 404 306
rect 50 275 404 278
rect 50 220 404 223
rect 50 192 87 220
rect 115 192 173 220
rect 201 192 259 220
rect 287 192 345 220
rect 373 192 404 220
rect 50 189 404 192
rect 50 134 404 137
rect 50 106 87 134
rect 115 106 173 134
rect 201 106 259 134
rect 287 106 345 134
rect 373 106 404 134
rect 50 103 404 106
rect 50 48 404 51
rect 50 20 87 48
rect 115 20 173 48
rect 201 20 259 48
rect 287 20 345 48
rect 373 20 404 48
rect 50 17 404 20
<< metal4 >>
rect 28 368 426 383
rect 84 309 118 368
rect 170 309 204 368
rect 256 309 290 368
rect 342 309 376 368
rect 73 275 129 309
rect 159 275 215 309
rect 245 275 301 309
rect 331 275 387 309
rect 84 223 118 275
rect 170 223 204 275
rect 256 223 290 275
rect 342 223 376 275
rect 73 189 129 223
rect 159 189 215 223
rect 245 189 301 223
rect 331 189 387 223
rect 84 137 118 189
rect 170 137 204 189
rect 256 137 290 189
rect 342 137 376 189
rect 73 103 129 137
rect 159 103 215 137
rect 245 103 301 137
rect 331 103 387 137
rect 84 51 118 103
rect 170 51 204 103
rect 256 51 290 103
rect 342 51 376 103
rect 73 17 129 51
rect 159 17 215 51
rect 245 17 301 51
rect 331 17 387 51
rect 84 -36 118 17
rect 170 -36 204 17
rect 256 -36 290 17
rect 342 -36 376 17
rect 28 -51 426 -36
<< comment >>
rect 28 351 42 358
rect 412 351 426 358
rect 28 -26 42 -19
rect 412 -26 426 -19
<< end >>
