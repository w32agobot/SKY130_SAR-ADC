* SPICE3 file created from adc_array_wafflecap_16(2)x300aF_28um2.ext - technology: sky130A

.subckt adc_array_wafflecap_16(2)x300aF_28um2 cbot ctop
C0 cfloating cbot 4.10fF
C1 ctop cbot 0.60fF
C2 cfloating ctop 0.65fF
C3 cbot VSUBS 2.16fF
C4 cfloating VSUBS 0.62fF
.ends
