magic
tech sky130A
magscale 1 2
timestamp 1662625284
<< nwell >>
rect -38 247 1878 582
<< pwell >>
rect 1 -17 1839 214
<< nmos >>
rect 152 95 952 179
rect 1146 80 1176 164
rect 1242 80 1272 164
rect 1446 80 1476 164
rect 1542 80 1572 164
<< pmos >>
rect 1124 296 1154 456
rect 1220 296 1250 456
rect 1540 296 1570 456
rect 1636 296 1666 456
<< pmoslvt >>
rect 152 283 952 443
<< ndiff >>
rect 94 167 152 179
rect 94 107 106 167
rect 140 107 152 167
rect 94 95 152 107
rect 952 167 1010 179
rect 952 107 964 167
rect 998 107 1010 167
rect 952 95 1010 107
rect 1086 152 1146 164
rect 1086 92 1096 152
rect 1130 92 1146 152
rect 1086 80 1146 92
rect 1176 152 1242 164
rect 1176 92 1192 152
rect 1226 92 1242 152
rect 1176 80 1242 92
rect 1272 152 1330 164
rect 1272 92 1288 152
rect 1322 92 1330 152
rect 1272 80 1330 92
rect 1384 152 1446 164
rect 1384 92 1396 152
rect 1430 92 1446 152
rect 1384 80 1446 92
rect 1476 152 1542 164
rect 1476 92 1492 152
rect 1526 92 1542 152
rect 1476 80 1542 92
rect 1572 152 1634 164
rect 1572 92 1588 152
rect 1622 92 1634 152
rect 1572 80 1634 92
<< pdiff >>
rect 1064 444 1124 456
rect 94 431 152 443
rect 94 295 106 431
rect 140 295 152 431
rect 94 283 152 295
rect 952 431 1010 443
rect 952 295 964 431
rect 998 295 1010 431
rect 1064 308 1074 444
rect 1108 308 1124 444
rect 1064 296 1124 308
rect 1154 444 1220 456
rect 1154 308 1170 444
rect 1204 308 1220 444
rect 1154 296 1220 308
rect 1250 444 1310 456
rect 1250 308 1266 444
rect 1300 308 1310 444
rect 1250 296 1310 308
rect 1478 444 1540 456
rect 1478 308 1490 444
rect 1524 308 1540 444
rect 1478 296 1540 308
rect 1570 444 1636 456
rect 1570 308 1586 444
rect 1620 308 1636 444
rect 1570 296 1636 308
rect 1666 444 1726 456
rect 1666 308 1682 444
rect 1716 308 1726 444
rect 1666 296 1726 308
rect 952 283 1010 295
<< ndiffc >>
rect 106 107 140 167
rect 964 107 998 167
rect 1096 92 1130 152
rect 1192 92 1226 152
rect 1288 92 1322 152
rect 1396 92 1430 152
rect 1492 92 1526 152
rect 1588 92 1622 152
<< pdiffc >>
rect 106 295 140 431
rect 964 295 998 431
rect 1074 308 1108 444
rect 1170 308 1204 444
rect 1266 308 1300 444
rect 1490 308 1524 444
rect 1586 308 1620 444
rect 1682 308 1716 444
<< poly >>
rect 152 443 952 479
rect 1124 456 1154 490
rect 1220 456 1250 490
rect 1540 456 1570 490
rect 1636 456 1666 490
rect 152 264 952 283
rect 17 254 952 264
rect 1124 280 1154 296
rect 1220 280 1250 296
rect 1124 258 1272 280
rect 17 248 278 254
rect 17 214 27 248
rect 62 214 278 248
rect 17 208 278 214
rect 1066 250 1272 258
rect 1066 248 1176 250
rect 1066 214 1104 248
rect 1138 214 1176 248
rect 17 198 952 208
rect 1066 202 1176 214
rect 152 179 952 198
rect 1146 164 1176 202
rect 1242 164 1272 250
rect 1332 252 1398 262
rect 1332 218 1348 252
rect 1382 220 1398 252
rect 1540 220 1570 296
rect 1636 220 1666 296
rect 1382 218 1666 220
rect 1332 190 1666 218
rect 1446 164 1476 190
rect 1542 164 1572 190
rect 152 69 952 95
rect 1146 54 1176 80
rect 1242 54 1272 80
rect 1446 54 1476 80
rect 1542 54 1572 80
<< polycont >>
rect 27 214 62 248
rect 1104 214 1138 248
rect 1348 218 1382 252
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1840 561
rect 106 431 140 447
rect 106 279 140 295
rect 964 431 998 447
rect 17 248 65 264
rect 17 214 27 248
rect 62 214 65 248
rect 17 198 65 214
rect 964 236 998 295
rect 1074 444 1108 527
rect 1074 292 1108 308
rect 1170 444 1204 460
rect 1170 292 1204 308
rect 1266 444 1300 460
rect 1266 292 1300 308
rect 1082 248 1154 258
rect 964 214 1082 236
rect 1138 214 1154 248
rect 964 202 1154 214
rect 1348 252 1382 268
rect 1416 258 1450 527
rect 1484 444 1524 460
rect 1484 308 1490 444
rect 1484 292 1524 308
rect 1586 444 1620 460
rect 1416 224 1526 258
rect 1348 202 1382 218
rect 106 167 140 183
rect 106 91 140 107
rect 964 167 998 202
rect 964 73 998 107
rect 1096 152 1130 168
rect 1096 17 1130 92
rect 1192 152 1226 168
rect 1192 76 1226 92
rect 1288 76 1322 92
rect 1396 152 1430 168
rect 1396 76 1430 92
rect 1492 152 1526 224
rect 1586 236 1620 308
rect 1682 444 1722 460
rect 1716 308 1722 444
rect 1682 292 1722 308
rect 1724 254 1770 258
rect 1586 202 1690 236
rect 1492 76 1526 92
rect 1588 152 1622 168
rect 1588 76 1622 92
rect 1656 17 1690 202
rect 1724 220 1730 254
rect 1764 220 1770 254
rect 1724 196 1770 220
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1840 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 106 295 140 431
rect 964 295 998 417
rect 1170 308 1204 444
rect 1266 308 1300 364
rect 1082 214 1104 248
rect 1104 214 1138 248
rect 1348 218 1382 252
rect 1490 328 1524 444
rect 106 107 140 167
rect 1192 92 1226 152
rect 1288 152 1322 178
rect 1288 144 1322 152
rect 1396 92 1430 132
rect 1682 328 1716 444
rect 1588 92 1622 132
rect 1730 220 1764 254
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
<< metal1 >>
rect 0 561 1840 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1840 561
rect 0 496 1840 527
rect 100 431 146 496
rect 1164 444 1722 456
rect 100 295 106 431
rect 140 295 146 431
rect 100 283 146 295
rect 958 417 1004 439
rect 958 295 964 417
rect 998 295 1004 417
rect 1164 308 1170 444
rect 1204 422 1490 444
rect 1204 308 1210 422
rect 1164 296 1210 308
rect 1260 364 1306 394
rect 1260 308 1266 364
rect 1300 308 1306 364
rect 1484 328 1490 422
rect 1524 422 1682 444
rect 1524 328 1530 422
rect 1484 316 1530 328
rect 1676 328 1682 422
rect 1716 328 1722 444
rect 1676 316 1722 328
rect 958 258 1004 295
rect 958 256 1154 258
rect 958 204 1082 256
rect 1138 204 1154 256
rect 1260 248 1306 308
rect 1342 252 1388 264
rect 1342 248 1348 252
rect 1260 220 1348 248
rect 958 202 1154 204
rect 1282 218 1348 220
rect 1382 248 1388 252
rect 1718 254 1776 260
rect 1718 248 1730 254
rect 1382 220 1730 248
rect 1764 220 1776 254
rect 1382 218 1388 220
rect 1282 206 1388 218
rect 1718 214 1776 220
rect 100 167 146 182
rect 100 107 106 167
rect 140 107 146 167
rect 1282 178 1328 206
rect 1186 152 1232 164
rect 100 48 146 107
rect 960 128 1064 136
rect 960 58 980 128
rect 1044 58 1064 128
rect 1186 92 1192 152
rect 1226 104 1232 152
rect 1282 144 1288 178
rect 1322 144 1328 178
rect 1282 132 1328 144
rect 1390 132 1436 144
rect 1390 104 1396 132
rect 1226 92 1396 104
rect 1430 104 1436 132
rect 1582 132 1628 144
rect 1582 104 1588 132
rect 1430 92 1588 104
rect 1622 92 1628 132
rect 1186 76 1628 92
rect 960 48 1064 58
rect 0 17 1840 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1840 17
rect 0 -48 1840 -17
<< via1 >>
rect 1082 248 1138 256
rect 1082 214 1138 248
rect 1082 204 1138 214
rect 980 58 1044 128
<< metal2 >>
rect 1008 270 1154 286
rect 1008 214 1018 270
rect 1076 256 1154 270
rect 1076 214 1082 256
rect 1008 204 1082 214
rect 1138 204 1154 256
rect 1008 168 1154 204
rect 960 134 1064 136
rect 960 58 980 134
rect 1044 58 1064 134
rect 960 48 1064 58
<< via2 >>
rect 1018 214 1076 270
rect 980 128 1044 134
rect 980 60 1044 128
<< metal3 >>
rect 139 140 934 496
rect 1006 274 1088 320
rect 1006 210 1016 274
rect 1080 210 1088 274
rect 1006 200 1088 210
rect 1174 140 1706 496
rect 139 134 1706 140
rect 139 60 980 134
rect 1044 60 1706 134
rect 139 54 1706 60
<< via3 >>
rect 1016 270 1080 274
rect 1016 214 1018 270
rect 1018 214 1076 270
rect 1076 214 1080 270
rect 1016 210 1080 214
<< mimcap >>
rect 167 264 906 468
rect 167 200 826 264
rect 890 200 906 264
rect 167 82 906 200
rect 1202 264 1678 468
rect 1202 200 1220 264
rect 1284 200 1678 264
rect 1202 82 1678 200
<< mimcapcontact >>
rect 826 200 890 264
rect 1220 200 1284 264
<< metal4 >>
rect 1006 274 1088 286
rect 1006 268 1016 274
rect 822 264 1016 268
rect 822 200 826 264
rect 890 210 1016 264
rect 1080 268 1088 274
rect 1080 264 1294 268
rect 1080 210 1220 264
rect 890 200 1220 210
rect 1284 200 1294 264
rect 822 194 1294 200
rect 1006 168 1088 194
<< labels >>
flabel locali s 30 221 64 255 7 FreeSans 160 0 0 0 in
port 1 nsew signal input
flabel metal1 s 0 496 1840 592 0 FreeSans 160 0 0 0 VPWR
port 3 nsew power bidirectional abutment
flabel metal1 s 213 527 247 561 0 FreeSans 160 0 0 0 VPWR
port 3 nsew power bidirectional abutment
flabel metal1 s 213 -17 247 17 0 FreeSans 160 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 0 -48 1840 48 0 FreeSans 160 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel nwell s 213 527 247 561 0 FreeSans 160 0 0 0 VPB
port 5 nsew power bidirectional
flabel pwell s 213 -17 247 17 0 FreeSans 160 0 0 0 VNB
port 6 nsew ground bidirectional
rlabel locali 964 169 998 169 1 cap_top
flabel metal1 s 1730 220 1764 254 0 FreeSans 160 0 0 0 out
port 2 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1840 544
string LEFclass CORE
string LEForigin 0 0
string LEFsite unithd
string LEFsource USER
<< end >>
