magic
tech sky130A
magscale 1 2
timestamp 1661518820
<< nwell >>
rect 2402 226 2858 230
rect 44 16 2858 226
rect 44 -178 2570 16
rect 44 -196 2336 -178
rect 570 -198 812 -196
rect 1178 -546 2336 -196
<< nmos >>
rect 144 -910 174 -510
rect 240 -910 270 -510
rect 336 -910 366 -510
rect 432 -910 462 -510
rect 528 -910 558 -510
rect 624 -910 654 -510
rect 720 -910 750 -510
rect 816 -910 846 -510
rect 144 -1170 174 -1070
rect 240 -1170 270 -1070
rect 336 -1170 366 -1070
rect 432 -1170 462 -1070
rect 528 -1170 558 -1070
rect 624 -1170 654 -1070
rect 720 -1170 750 -1070
rect 816 -1170 846 -1070
rect 1598 -1176 1628 -776
rect 1694 -1176 1724 -776
rect 1790 -1176 1820 -776
rect 1886 -1176 1916 -776
<< pmos >>
rect 144 -96 174 4
rect 240 -96 270 4
rect 336 -96 366 4
rect 432 -96 462 4
rect 528 -96 558 4
rect 624 -96 654 4
rect 720 -96 750 4
rect 816 -96 846 4
rect 1276 -446 1306 -46
rect 1372 -446 1402 -46
rect 1598 -446 1628 -46
rect 1694 -446 1724 -46
rect 1790 -446 1820 -46
rect 1886 -446 1916 -46
rect 2112 -446 2142 -46
rect 2208 -446 2238 -46
<< ndiff >>
rect 82 -522 144 -510
rect 82 -898 94 -522
rect 128 -898 144 -522
rect 82 -910 144 -898
rect 174 -522 240 -510
rect 174 -898 190 -522
rect 224 -898 240 -522
rect 174 -910 240 -898
rect 270 -522 336 -510
rect 270 -898 286 -522
rect 320 -898 336 -522
rect 270 -910 336 -898
rect 366 -522 432 -510
rect 366 -898 382 -522
rect 416 -898 432 -522
rect 366 -910 432 -898
rect 462 -522 528 -510
rect 462 -898 478 -522
rect 512 -898 528 -522
rect 462 -910 528 -898
rect 558 -522 624 -510
rect 558 -898 574 -522
rect 608 -898 624 -522
rect 558 -910 624 -898
rect 654 -522 720 -510
rect 654 -898 670 -522
rect 704 -898 720 -522
rect 654 -910 720 -898
rect 750 -522 816 -510
rect 750 -898 766 -522
rect 800 -898 816 -522
rect 750 -910 816 -898
rect 846 -522 908 -510
rect 846 -898 862 -522
rect 896 -898 908 -522
rect 846 -910 908 -898
rect 1536 -788 1598 -776
rect 82 -1082 144 -1070
rect 82 -1158 94 -1082
rect 128 -1158 144 -1082
rect 82 -1170 144 -1158
rect 174 -1082 240 -1070
rect 174 -1158 190 -1082
rect 224 -1158 240 -1082
rect 174 -1170 240 -1158
rect 270 -1082 336 -1070
rect 270 -1158 286 -1082
rect 320 -1158 336 -1082
rect 270 -1170 336 -1158
rect 366 -1082 432 -1070
rect 366 -1158 382 -1082
rect 416 -1158 432 -1082
rect 366 -1170 432 -1158
rect 462 -1082 528 -1070
rect 462 -1158 478 -1082
rect 512 -1158 528 -1082
rect 462 -1170 528 -1158
rect 558 -1082 624 -1070
rect 558 -1158 574 -1082
rect 608 -1158 624 -1082
rect 558 -1170 624 -1158
rect 654 -1082 720 -1070
rect 654 -1158 670 -1082
rect 704 -1158 720 -1082
rect 654 -1170 720 -1158
rect 750 -1082 816 -1070
rect 750 -1158 766 -1082
rect 800 -1158 816 -1082
rect 750 -1170 816 -1158
rect 846 -1082 908 -1070
rect 846 -1158 862 -1082
rect 896 -1158 908 -1082
rect 846 -1170 908 -1158
rect 1536 -1164 1548 -788
rect 1582 -1164 1598 -788
rect 1536 -1176 1598 -1164
rect 1628 -788 1694 -776
rect 1628 -1164 1644 -788
rect 1678 -1164 1694 -788
rect 1628 -1176 1694 -1164
rect 1724 -788 1790 -776
rect 1724 -1164 1740 -788
rect 1774 -1164 1790 -788
rect 1724 -1176 1790 -1164
rect 1820 -788 1886 -776
rect 1820 -1164 1836 -788
rect 1870 -1164 1886 -788
rect 1820 -1176 1886 -1164
rect 1916 -788 1978 -776
rect 1916 -1164 1932 -788
rect 1966 -1164 1978 -788
rect 1916 -1176 1978 -1164
<< pdiff >>
rect 82 -8 144 4
rect 82 -84 94 -8
rect 128 -84 144 -8
rect 82 -96 144 -84
rect 174 -8 240 4
rect 174 -84 190 -8
rect 224 -84 240 -8
rect 174 -96 240 -84
rect 270 -8 336 4
rect 270 -84 286 -8
rect 320 -84 336 -8
rect 270 -96 336 -84
rect 366 -8 432 4
rect 366 -84 382 -8
rect 416 -84 432 -8
rect 366 -96 432 -84
rect 462 -8 528 4
rect 462 -84 478 -8
rect 512 -84 528 -8
rect 462 -96 528 -84
rect 558 -8 624 4
rect 558 -84 574 -8
rect 608 -84 624 -8
rect 558 -96 624 -84
rect 654 -8 720 4
rect 654 -84 670 -8
rect 704 -84 720 -8
rect 654 -96 720 -84
rect 750 -8 816 4
rect 750 -84 766 -8
rect 800 -84 816 -8
rect 750 -96 816 -84
rect 846 -8 908 4
rect 846 -84 862 -8
rect 896 -84 908 -8
rect 846 -96 908 -84
rect 1214 -58 1276 -46
rect 1214 -434 1226 -58
rect 1260 -434 1276 -58
rect 1214 -446 1276 -434
rect 1306 -58 1372 -46
rect 1306 -434 1322 -58
rect 1356 -434 1372 -58
rect 1306 -446 1372 -434
rect 1402 -58 1464 -46
rect 1402 -434 1418 -58
rect 1452 -434 1464 -58
rect 1402 -446 1464 -434
rect 1536 -58 1598 -46
rect 1536 -434 1548 -58
rect 1582 -434 1598 -58
rect 1536 -446 1598 -434
rect 1628 -58 1694 -46
rect 1628 -434 1644 -58
rect 1678 -434 1694 -58
rect 1628 -446 1694 -434
rect 1724 -58 1790 -46
rect 1724 -434 1740 -58
rect 1774 -434 1790 -58
rect 1724 -446 1790 -434
rect 1820 -58 1886 -46
rect 1820 -434 1836 -58
rect 1870 -434 1886 -58
rect 1820 -446 1886 -434
rect 1916 -58 1978 -46
rect 1916 -434 1932 -58
rect 1966 -434 1978 -58
rect 1916 -446 1978 -434
rect 2050 -58 2112 -46
rect 2050 -434 2062 -58
rect 2096 -434 2112 -58
rect 2050 -446 2112 -434
rect 2142 -58 2208 -46
rect 2142 -434 2158 -58
rect 2192 -434 2208 -58
rect 2142 -446 2208 -434
rect 2238 -58 2300 -46
rect 2238 -434 2254 -58
rect 2288 -434 2300 -58
rect 2238 -446 2300 -434
<< ndiffc >>
rect 94 -898 128 -522
rect 190 -898 224 -522
rect 286 -898 320 -522
rect 382 -898 416 -522
rect 478 -898 512 -522
rect 574 -898 608 -522
rect 670 -898 704 -522
rect 766 -898 800 -522
rect 862 -898 896 -522
rect 94 -1158 128 -1082
rect 190 -1158 224 -1082
rect 286 -1158 320 -1082
rect 382 -1158 416 -1082
rect 478 -1158 512 -1082
rect 574 -1158 608 -1082
rect 670 -1158 704 -1082
rect 766 -1158 800 -1082
rect 862 -1158 896 -1082
rect 1548 -1164 1582 -788
rect 1644 -1164 1678 -788
rect 1740 -1164 1774 -788
rect 1836 -1164 1870 -788
rect 1932 -1164 1966 -788
<< pdiffc >>
rect 94 -84 128 -8
rect 190 -84 224 -8
rect 286 -84 320 -8
rect 382 -84 416 -8
rect 478 -84 512 -8
rect 574 -84 608 -8
rect 670 -84 704 -8
rect 766 -84 800 -8
rect 862 -84 896 -8
rect 1226 -434 1260 -58
rect 1322 -434 1356 -58
rect 1418 -434 1452 -58
rect 1548 -434 1582 -58
rect 1644 -434 1678 -58
rect 1740 -434 1774 -58
rect 1836 -434 1870 -58
rect 1932 -434 1966 -58
rect 2062 -434 2096 -58
rect 2158 -434 2192 -58
rect 2254 -434 2288 -58
<< psubdiff >>
rect -286 3826 -164 3852
rect -286 3752 -262 3826
rect -188 3752 -164 3826
rect -286 3728 -164 3752
rect 262 3826 384 3852
rect 262 3752 286 3826
rect 360 3752 384 3826
rect 262 3728 384 3752
rect 810 3826 932 3852
rect 810 3752 834 3826
rect 908 3752 932 3826
rect 810 3728 932 3752
rect 1358 3826 1480 3852
rect 1358 3752 1382 3826
rect 1456 3752 1480 3826
rect 1358 3728 1480 3752
rect 1906 3826 2028 3852
rect 1906 3752 1930 3826
rect 2004 3752 2028 3826
rect 1906 3728 2028 3752
rect 2436 3826 2558 3852
rect 2436 3752 2460 3826
rect 2534 3752 2558 3826
rect 2436 3728 2558 3752
rect 2984 3826 3106 3852
rect 2984 3752 3008 3826
rect 3082 3752 3106 3826
rect 2984 3728 3106 3752
rect 3534 3826 3656 3852
rect 3534 3752 3558 3826
rect 3632 3752 3656 3826
rect 3534 3728 3656 3752
rect -652 3350 -530 3376
rect -652 3276 -628 3350
rect -554 3276 -530 3350
rect -652 3252 -530 3276
rect 4030 3282 4152 3308
rect 4030 3208 4054 3282
rect 4128 3208 4152 3282
rect 4030 3184 4152 3208
rect -652 2876 -530 2902
rect -652 2802 -628 2876
rect -554 2802 -530 2876
rect -652 2778 -530 2802
rect 4030 2808 4152 2834
rect 4030 2734 4054 2808
rect 4128 2734 4152 2808
rect 4030 2710 4152 2734
rect -652 2402 -530 2428
rect -652 2328 -628 2402
rect -554 2328 -530 2402
rect -652 2304 -530 2328
rect 4030 2334 4152 2360
rect 4030 2260 4054 2334
rect 4128 2260 4152 2334
rect 4030 2236 4152 2260
rect -652 1928 -530 1954
rect -652 1854 -628 1928
rect -554 1854 -530 1928
rect -652 1830 -530 1854
rect 4030 1858 4152 1884
rect 4030 1784 4054 1858
rect 4128 1784 4152 1858
rect 4030 1760 4152 1784
rect -652 1454 -530 1480
rect -652 1380 -628 1454
rect -554 1380 -530 1454
rect -652 1356 -530 1380
rect 4030 1382 4152 1408
rect 4030 1308 4054 1382
rect 4128 1308 4152 1382
rect 4030 1284 4152 1308
rect -652 980 -530 1006
rect -652 906 -628 980
rect -554 906 -530 980
rect -652 882 -530 906
rect 4030 908 4152 934
rect 4030 834 4054 908
rect 4128 834 4152 908
rect 4030 810 4152 834
rect -652 506 -530 532
rect -652 432 -628 506
rect -554 432 -530 506
rect -652 408 -530 432
rect 4028 434 4150 460
rect 4028 360 4052 434
rect 4126 360 4150 434
rect 4028 288 4150 360
rect -652 -88 -530 -62
rect -652 -162 -628 -88
rect -554 -162 -530 -88
rect -652 -186 -530 -162
rect 4028 -86 4150 -60
rect 4028 -160 4052 -86
rect 4126 -160 4150 -86
rect 4028 -184 4150 -160
rect -660 -614 -538 -588
rect -660 -688 -636 -614
rect -562 -688 -538 -614
rect -660 -712 -538 -688
rect 2474 -530 2826 -514
rect 2474 -564 2508 -530
rect 2542 -564 2594 -530
rect 2628 -564 2680 -530
rect 2714 -564 2766 -530
rect 2800 -564 2826 -530
rect 2474 -582 2826 -564
rect 4028 -560 4150 -534
rect 4028 -634 4052 -560
rect 4126 -634 4150 -560
rect 4028 -658 4150 -634
rect -660 -1088 -538 -1062
rect -660 -1162 -636 -1088
rect -562 -1162 -538 -1088
rect -660 -1186 -538 -1162
rect 4028 -1034 4150 -1008
rect 4028 -1108 4052 -1034
rect 4126 -1108 4150 -1034
rect 4028 -1132 4150 -1108
rect 1542 -1324 1566 -1288
rect 1602 -1324 1658 -1288
rect 1694 -1324 1750 -1288
rect 1786 -1324 1842 -1288
rect 1878 -1324 1934 -1288
rect 1970 -1324 1994 -1288
rect 1542 -1326 1994 -1324
rect 76 -1332 894 -1330
rect 76 -1368 100 -1332
rect 136 -1368 218 -1332
rect 254 -1368 336 -1332
rect 372 -1368 454 -1332
rect 490 -1368 572 -1332
rect 608 -1368 690 -1332
rect 726 -1368 808 -1332
rect 844 -1368 894 -1332
rect 76 -1372 894 -1368
rect -646 -1740 -524 -1714
rect -646 -1814 -622 -1740
rect -548 -1814 -524 -1740
rect -646 -1838 -524 -1814
rect 4028 -1770 4150 -1744
rect 4028 -1844 4052 -1770
rect 4126 -1844 4150 -1770
rect 4028 -1868 4150 -1844
rect -646 -2214 -524 -2188
rect -646 -2288 -622 -2214
rect -548 -2288 -524 -2214
rect -646 -2312 -524 -2288
rect 4028 -2244 4150 -2218
rect 4028 -2318 4052 -2244
rect 4126 -2318 4150 -2244
rect 4028 -2342 4150 -2318
rect -646 -2688 -524 -2662
rect -646 -2762 -622 -2688
rect -548 -2762 -524 -2688
rect -646 -2786 -524 -2762
rect 4028 -2718 4150 -2692
rect 4028 -2792 4052 -2718
rect 4126 -2792 4150 -2718
rect 4028 -2816 4150 -2792
rect -646 -3164 -524 -3138
rect -646 -3238 -622 -3164
rect -548 -3238 -524 -3164
rect -646 -3262 -524 -3238
rect 4028 -3192 4150 -3166
rect 4028 -3266 4052 -3192
rect 4126 -3266 4150 -3192
rect 4028 -3290 4150 -3266
rect -646 -3638 -524 -3612
rect -646 -3712 -622 -3638
rect -548 -3712 -524 -3638
rect -646 -3736 -524 -3712
rect 4028 -3666 4150 -3640
rect 4028 -3740 4052 -3666
rect 4126 -3740 4150 -3666
rect 4028 -3764 4150 -3740
rect -646 -4112 -524 -4086
rect -646 -4186 -622 -4112
rect -548 -4186 -524 -4112
rect -646 -4210 -524 -4186
rect 4028 -4140 4150 -4114
rect 4028 -4214 4052 -4140
rect 4126 -4214 4150 -4140
rect 4028 -4238 4150 -4214
rect -646 -4586 -524 -4560
rect -646 -4660 -622 -4586
rect -548 -4660 -524 -4586
rect -646 -4684 -524 -4660
rect 4030 -4614 4152 -4588
rect 4030 -4688 4054 -4614
rect 4128 -4688 4152 -4614
rect 4030 -4712 4152 -4688
rect -116 -5000 6 -4974
rect -116 -5074 -92 -5000
rect -18 -5074 6 -5000
rect -116 -5098 6 -5074
rect 432 -5000 554 -4974
rect 432 -5074 456 -5000
rect 530 -5074 554 -5000
rect 432 -5098 554 -5074
rect 980 -5000 1102 -4974
rect 980 -5074 1004 -5000
rect 1078 -5074 1102 -5000
rect 980 -5098 1102 -5074
rect 1528 -5000 1650 -4974
rect 1528 -5074 1552 -5000
rect 1626 -5074 1650 -5000
rect 1528 -5098 1650 -5074
rect 2076 -5000 2198 -4974
rect 2076 -5074 2100 -5000
rect 2174 -5074 2198 -5000
rect 2076 -5098 2198 -5074
rect 2624 -5000 2746 -4974
rect 2624 -5074 2648 -5000
rect 2722 -5074 2746 -5000
rect 2624 -5098 2746 -5074
rect 3174 -5000 3296 -4974
rect 3174 -5074 3198 -5000
rect 3272 -5074 3296 -5000
rect 3174 -5098 3296 -5074
<< nsubdiff >>
rect 1382 110 2106 118
rect 82 100 938 108
rect 82 66 112 100
rect 146 66 196 100
rect 230 66 280 100
rect 314 66 364 100
rect 398 66 448 100
rect 482 66 532 100
rect 566 66 616 100
rect 650 66 700 100
rect 734 66 784 100
rect 818 66 874 100
rect 908 66 938 100
rect 1382 76 1420 110
rect 1454 76 1504 110
rect 1538 76 1588 110
rect 1622 76 1672 110
rect 1706 76 1756 110
rect 1790 76 1840 110
rect 1874 76 1924 110
rect 1958 76 2008 110
rect 2042 76 2106 110
rect 1382 70 2106 76
rect 82 60 938 66
<< psubdiffcont >>
rect -262 3752 -188 3826
rect 286 3752 360 3826
rect 834 3752 908 3826
rect 1382 3752 1456 3826
rect 1930 3752 2004 3826
rect 2460 3752 2534 3826
rect 3008 3752 3082 3826
rect 3558 3752 3632 3826
rect -628 3276 -554 3350
rect 4054 3208 4128 3282
rect -628 2802 -554 2876
rect 4054 2734 4128 2808
rect -628 2328 -554 2402
rect 4054 2260 4128 2334
rect -628 1854 -554 1928
rect 4054 1784 4128 1858
rect -628 1380 -554 1454
rect 4054 1308 4128 1382
rect -628 906 -554 980
rect 4054 834 4128 908
rect -628 432 -554 506
rect 4052 360 4126 434
rect -628 -162 -554 -88
rect 4052 -160 4126 -86
rect -636 -688 -562 -614
rect 2508 -564 2542 -530
rect 2594 -564 2628 -530
rect 2680 -564 2714 -530
rect 2766 -564 2800 -530
rect 4052 -634 4126 -560
rect -636 -1162 -562 -1088
rect 4052 -1108 4126 -1034
rect 1566 -1324 1602 -1288
rect 1658 -1324 1694 -1288
rect 1750 -1324 1786 -1288
rect 1842 -1324 1878 -1288
rect 1934 -1324 1970 -1288
rect 100 -1368 136 -1332
rect 218 -1368 254 -1332
rect 336 -1368 372 -1332
rect 454 -1368 490 -1332
rect 572 -1368 608 -1332
rect 690 -1368 726 -1332
rect 808 -1368 844 -1332
rect -622 -1814 -548 -1740
rect 4052 -1844 4126 -1770
rect -622 -2288 -548 -2214
rect 4052 -2318 4126 -2244
rect -622 -2762 -548 -2688
rect 4052 -2792 4126 -2718
rect -622 -3238 -548 -3164
rect 4052 -3266 4126 -3192
rect -622 -3712 -548 -3638
rect 4052 -3740 4126 -3666
rect -622 -4186 -548 -4112
rect 4052 -4214 4126 -4140
rect -622 -4660 -548 -4586
rect 4054 -4688 4128 -4614
rect -92 -5074 -18 -5000
rect 456 -5074 530 -5000
rect 1004 -5074 1078 -5000
rect 1552 -5074 1626 -5000
rect 2100 -5074 2174 -5000
rect 2648 -5074 2722 -5000
rect 3198 -5074 3272 -5000
<< nsubdiffcont >>
rect 112 66 146 100
rect 196 66 230 100
rect 280 66 314 100
rect 364 66 398 100
rect 448 66 482 100
rect 532 66 566 100
rect 616 66 650 100
rect 700 66 734 100
rect 784 66 818 100
rect 874 66 908 100
rect 1420 76 1454 110
rect 1504 76 1538 110
rect 1588 76 1622 110
rect 1672 76 1706 110
rect 1756 76 1790 110
rect 1840 76 1874 110
rect 1924 76 1958 110
rect 2008 76 2042 110
<< poly >>
rect 144 4 174 30
rect 240 4 270 30
rect 336 4 366 30
rect 432 4 462 30
rect 528 4 558 30
rect 624 4 654 30
rect 720 4 750 30
rect 816 4 846 30
rect 1276 -46 1306 -20
rect 1372 -46 1402 -20
rect 1598 -46 1628 -20
rect 1694 -46 1724 -20
rect 1790 -46 1820 -20
rect 1886 -46 1916 -20
rect 2112 -46 2142 -20
rect 2208 -46 2238 -20
rect 144 -122 174 -96
rect 240 -122 270 -96
rect 336 -122 366 -96
rect 432 -122 462 -96
rect 528 -122 558 -96
rect 624 -122 654 -96
rect 720 -122 750 -96
rect 816 -122 846 -96
rect 144 -154 846 -122
rect 466 -196 524 -154
rect -14 -206 524 -196
rect -14 -240 2 -206
rect 36 -232 524 -206
rect 36 -240 52 -232
rect -14 -254 52 -240
rect 652 -284 724 -274
rect 652 -324 668 -284
rect 708 -324 724 -284
rect 260 -334 332 -324
rect 652 -334 724 -324
rect 260 -374 276 -334
rect 316 -374 332 -334
rect 260 -384 332 -374
rect 284 -454 322 -384
rect 668 -454 706 -334
rect 1100 -368 1168 -358
rect 1100 -404 1116 -368
rect 1152 -404 1168 -368
rect 1100 -442 1168 -404
rect 144 -484 462 -454
rect 144 -510 174 -484
rect 240 -510 270 -484
rect 336 -510 366 -484
rect 432 -510 462 -484
rect 528 -484 846 -454
rect 528 -510 558 -484
rect 624 -510 654 -484
rect 720 -510 750 -484
rect 816 -510 846 -484
rect 1100 -478 1116 -442
rect 1152 -462 1168 -442
rect 2396 -206 2470 -190
rect 2396 -240 2410 -206
rect 2446 -240 2470 -206
rect 2396 -278 2470 -240
rect 2396 -312 2410 -278
rect 2446 -312 2470 -278
rect 2396 -328 2470 -312
rect 1276 -462 1306 -446
rect 1372 -462 1402 -446
rect 1152 -478 1402 -462
rect 1100 -492 1402 -478
rect 1598 -462 1628 -446
rect 1694 -462 1724 -446
rect 1598 -492 1724 -462
rect 1690 -558 1724 -492
rect 1658 -568 1724 -558
rect 1658 -602 1674 -568
rect 1708 -602 1724 -568
rect 1658 -612 1724 -602
rect 1598 -776 1628 -750
rect 1694 -776 1724 -612
rect 1790 -462 1820 -446
rect 1886 -462 1916 -446
rect 1790 -492 1916 -462
rect 2112 -462 2142 -446
rect 2208 -462 2238 -446
rect 2112 -492 2238 -462
rect 1790 -626 1824 -492
rect 1790 -636 2050 -626
rect 1790 -670 1808 -636
rect 1842 -670 2050 -636
rect 2204 -668 2238 -492
rect 1790 -680 2050 -670
rect 1790 -776 1820 -680
rect 1886 -776 1916 -750
rect 144 -938 174 -910
rect 240 -938 270 -910
rect 336 -938 366 -910
rect 432 -938 462 -910
rect 528 -938 558 -910
rect 624 -938 654 -910
rect 720 -938 750 -910
rect 816 -938 846 -910
rect -6 -1004 60 -994
rect -6 -1038 10 -1004
rect 44 -1014 60 -1004
rect 44 -1038 846 -1014
rect -6 -1044 846 -1038
rect -6 -1048 60 -1044
rect 144 -1070 174 -1044
rect 240 -1070 270 -1044
rect 336 -1070 366 -1044
rect 432 -1070 462 -1044
rect 528 -1070 558 -1044
rect 624 -1070 654 -1044
rect 720 -1070 750 -1044
rect 816 -1070 846 -1044
rect 144 -1196 174 -1170
rect 240 -1196 270 -1170
rect 336 -1196 366 -1170
rect 432 -1196 462 -1170
rect 528 -1196 558 -1170
rect 624 -1196 654 -1170
rect 720 -1196 750 -1170
rect 816 -1196 846 -1170
rect 1994 -796 2050 -680
rect 2108 -684 2238 -668
rect 2108 -720 2118 -684
rect 2154 -720 2192 -684
rect 2228 -720 2238 -684
rect 2108 -736 2238 -720
rect 1994 -852 2466 -796
rect 1598 -1244 1628 -1176
rect 1694 -1202 1724 -1176
rect 1790 -1202 1820 -1176
rect 1886 -1244 1916 -1176
rect 1440 -1254 1916 -1244
rect 1440 -1288 1456 -1254
rect 1490 -1274 1916 -1254
rect 1490 -1288 1506 -1274
rect 1440 -1298 1506 -1288
<< polycont >>
rect 2 -240 36 -206
rect 668 -324 708 -284
rect 276 -374 316 -334
rect 1116 -404 1152 -368
rect 1116 -478 1152 -442
rect 2410 -240 2446 -206
rect 2410 -312 2446 -278
rect 1674 -602 1708 -568
rect 1808 -670 1842 -636
rect 10 -1038 44 -1004
rect 2118 -720 2154 -684
rect 2192 -720 2228 -684
rect 1456 -1288 1490 -1254
<< locali >>
rect -686 3826 4192 3882
rect -686 3752 -262 3826
rect -188 3752 286 3826
rect 360 3752 834 3826
rect 908 3752 1382 3826
rect 1456 3752 1930 3826
rect 2004 3752 2460 3826
rect 2534 3752 3008 3826
rect 3082 3752 3558 3826
rect 3632 3752 4192 3826
rect -686 3684 4192 3752
rect -686 3350 -488 3684
rect -686 3276 -628 3350
rect -554 3276 -488 3350
rect -686 2876 -488 3276
rect -686 2802 -628 2876
rect -554 2802 -488 2876
rect -686 2402 -488 2802
rect -686 2328 -628 2402
rect -554 2328 -488 2402
rect -686 1928 -488 2328
rect -686 1854 -628 1928
rect -554 1854 -488 1928
rect -686 1454 -488 1854
rect -686 1380 -628 1454
rect -554 1380 -488 1454
rect -686 980 -488 1380
rect -686 906 -628 980
rect -554 906 -488 980
rect -686 512 -488 906
rect 3994 3282 4192 3684
rect 3994 3208 4054 3282
rect 4128 3208 4192 3282
rect 3994 2808 4192 3208
rect 3994 2734 4054 2808
rect 4128 2734 4192 2808
rect 3994 2334 4192 2734
rect 3994 2260 4054 2334
rect 4128 2260 4192 2334
rect 3994 1858 4192 2260
rect 3994 1784 4054 1858
rect 4128 1784 4192 1858
rect 3994 1382 4192 1784
rect 3994 1308 4054 1382
rect 4128 1308 4192 1382
rect 3994 908 4192 1308
rect 3994 834 4054 908
rect 4128 834 4192 908
rect 3994 512 4192 834
rect -686 506 788 512
rect -686 432 -628 506
rect -554 472 788 506
rect -554 432 -156 472
rect -686 406 -156 432
rect -92 406 -48 472
rect 16 406 60 472
rect 124 406 168 472
rect 232 406 276 472
rect 340 406 384 472
rect 448 406 492 472
rect 556 406 600 472
rect 664 406 708 472
rect 772 406 788 472
rect 2016 474 4192 512
rect 2016 472 2258 474
rect -686 384 788 406
rect 938 414 1050 430
rect -686 -88 -488 384
rect 938 348 950 414
rect 1032 348 1050 414
rect 938 328 1050 348
rect 82 100 938 108
rect 82 66 112 100
rect 146 66 196 100
rect 230 66 280 100
rect 314 66 364 100
rect 398 66 448 100
rect 482 66 532 100
rect 566 66 616 100
rect 650 66 700 100
rect 734 66 784 100
rect 818 66 874 100
rect 908 66 938 100
rect 82 60 938 66
rect -686 -162 -628 -88
rect -554 -162 -488 -88
rect 94 42 896 60
rect 94 -8 128 42
rect 94 -100 128 -84
rect 190 -8 224 8
rect -686 -614 -488 -162
rect 190 -160 224 -84
rect 286 -8 320 42
rect 286 -100 320 -84
rect 382 -8 416 8
rect 382 -160 416 -84
rect 478 -8 512 42
rect 478 -100 512 -84
rect 574 -8 608 8
rect 190 -194 416 -160
rect 574 -160 608 -84
rect 670 -8 704 42
rect 670 -100 704 -84
rect 766 -8 800 8
rect 766 -160 800 -84
rect 862 -8 896 42
rect 862 -100 896 -84
rect 574 -194 800 -160
rect -14 -206 52 -196
rect -14 -240 2 -206
rect 36 -240 52 -206
rect -14 -254 52 -240
rect -686 -688 -636 -614
rect -562 -688 -488 -614
rect -686 -1088 -488 -688
rect 6 -994 52 -254
rect 190 -418 224 -194
rect 260 -334 332 -324
rect 260 -374 276 -334
rect 316 -374 332 -334
rect 260 -384 332 -374
rect 368 -364 416 -358
rect 368 -400 374 -364
rect 410 -400 416 -364
rect 368 -418 416 -400
rect 190 -452 416 -418
rect 94 -522 128 -506
rect 94 -948 128 -898
rect 190 -522 224 -452
rect 190 -914 224 -898
rect 286 -522 320 -506
rect 286 -948 320 -898
rect 382 -522 416 -452
rect 574 -416 608 -194
rect 652 -284 724 -274
rect 652 -324 668 -284
rect 708 -324 724 -284
rect 652 -334 724 -324
rect 974 -416 1050 328
rect 574 -450 1050 -416
rect 382 -914 416 -898
rect 478 -522 512 -506
rect 478 -948 512 -898
rect 574 -522 608 -450
rect 574 -914 608 -898
rect 670 -522 704 -506
rect 670 -948 704 -898
rect 766 -522 800 -450
rect 766 -914 800 -898
rect 862 -522 896 -506
rect 862 -948 896 -898
rect 94 -984 896 -948
rect -6 -1004 60 -994
rect -6 -1038 10 -1004
rect 44 -1038 60 -1004
rect -6 -1048 60 -1038
rect -686 -1162 -636 -1088
rect -562 -1162 -488 -1088
rect -686 -1222 -488 -1162
rect 94 -1082 128 -984
rect 94 -1174 128 -1158
rect 190 -1082 224 -1064
rect -686 -1256 -670 -1222
rect -636 -1256 -598 -1222
rect -564 -1256 -526 -1222
rect -492 -1256 -488 -1222
rect -686 -1294 -488 -1256
rect -686 -1328 -670 -1294
rect -636 -1328 -598 -1294
rect -564 -1328 -526 -1294
rect -492 -1328 -488 -1294
rect -686 -1366 -488 -1328
rect 190 -1316 224 -1158
rect 286 -1082 320 -984
rect 286 -1174 320 -1158
rect 382 -1082 416 -1066
rect 382 -1316 416 -1158
rect 478 -1082 512 -984
rect 478 -1174 512 -1158
rect 574 -1082 608 -1066
rect 574 -1316 608 -1158
rect 670 -1082 704 -984
rect 670 -1174 704 -1158
rect 766 -1082 800 -1066
rect 766 -1316 800 -1158
rect 862 -1082 896 -984
rect 862 -1174 896 -1158
rect 974 -620 1050 -450
rect 974 -656 994 -620
rect 1030 -656 1050 -620
rect 974 -694 1050 -656
rect 974 -730 994 -694
rect 1030 -730 1050 -694
rect 190 -1330 800 -1316
rect -686 -1400 -670 -1366
rect -636 -1400 -598 -1366
rect -564 -1400 -526 -1366
rect -492 -1400 -488 -1366
rect 76 -1332 894 -1330
rect 76 -1368 100 -1332
rect 136 -1368 218 -1332
rect 254 -1368 336 -1332
rect 372 -1368 454 -1332
rect 490 -1368 572 -1332
rect 608 -1368 690 -1332
rect 726 -1368 808 -1332
rect 844 -1368 894 -1332
rect 76 -1372 894 -1368
rect -686 -1438 -488 -1400
rect -686 -1472 -670 -1438
rect -636 -1472 -598 -1438
rect -564 -1472 -526 -1438
rect -492 -1472 -488 -1438
rect -686 -1700 -488 -1472
rect 974 -1586 1050 -730
rect 954 -1602 1050 -1586
rect 954 -1668 968 -1602
rect 1042 -1668 1050 -1602
rect 954 -1680 1050 -1668
rect 1096 416 1222 432
rect 1096 350 1134 416
rect 1204 350 1222 416
rect 2016 406 2042 472
rect 2106 406 2150 472
rect 2214 408 2258 472
rect 2318 472 4192 474
rect 2318 408 2358 472
rect 2214 406 2358 408
rect 2422 406 2468 472
rect 2532 406 2576 472
rect 2640 406 2682 472
rect 2746 406 2792 472
rect 2856 406 2900 472
rect 2964 406 3008 472
rect 3072 406 3116 472
rect 3180 406 3224 472
rect 3288 406 3336 472
rect 3400 406 3444 472
rect 3508 406 3552 472
rect 3616 434 4192 472
rect 3616 406 4052 434
rect 2016 382 4052 406
rect 1096 328 1222 350
rect 3994 360 4052 382
rect 4126 360 4192 434
rect 1096 -368 1172 328
rect 2404 230 2952 250
rect 2404 194 2498 230
rect 2534 194 2574 230
rect 2610 194 2650 230
rect 2686 194 2726 230
rect 2762 194 2802 230
rect 2838 194 2878 230
rect 2914 194 2952 230
rect 2404 152 2952 194
rect 1382 110 2106 118
rect 1382 76 1420 110
rect 1454 76 1504 110
rect 1538 76 1588 110
rect 1622 76 1672 110
rect 1706 76 1756 110
rect 1790 76 1840 110
rect 1874 76 1924 110
rect 1958 76 2008 110
rect 2042 76 2106 110
rect 1382 70 2106 76
rect 1718 36 1808 70
rect 1096 -404 1116 -368
rect 1152 -404 1172 -368
rect 1096 -442 1172 -404
rect 1096 -478 1116 -442
rect 1152 -478 1172 -442
rect 1096 -1586 1172 -478
rect 1226 -8 1452 26
rect 1226 -58 1260 -8
rect 1226 -568 1260 -434
rect 1322 -58 1356 -42
rect 1322 -500 1356 -434
rect 1418 -58 1452 -8
rect 1418 -450 1452 -434
rect 1548 2 1966 36
rect 1548 -58 1582 2
rect 1548 -450 1582 -434
rect 1644 -58 1678 -42
rect 1644 -500 1678 -434
rect 1740 -58 1774 2
rect 1740 -450 1774 -434
rect 1836 -58 1870 -42
rect 1322 -534 1678 -500
rect 1836 -500 1870 -434
rect 1932 -58 1966 2
rect 1932 -450 1966 -434
rect 2062 -8 2288 26
rect 2062 -58 2096 -8
rect 2062 -450 2096 -434
rect 2158 -58 2192 -42
rect 2158 -500 2192 -434
rect 1836 -534 2192 -500
rect 2254 -58 2288 -8
rect 2288 -206 2452 -190
rect 2288 -240 2410 -206
rect 2446 -240 2452 -206
rect 2288 -278 2452 -240
rect 2288 -312 2410 -278
rect 2446 -312 2452 -278
rect 2786 -234 2846 -224
rect 2786 -236 2860 -234
rect 2786 -272 2792 -236
rect 2828 -272 2860 -236
rect 2786 -284 2846 -272
rect 2288 -328 2452 -312
rect 2254 -568 2288 -434
rect 2338 -530 2856 -514
rect 2338 -564 2508 -530
rect 2542 -564 2594 -530
rect 2628 -564 2680 -530
rect 2714 -564 2766 -530
rect 2800 -564 2856 -530
rect 1210 -602 1622 -568
rect 1658 -602 1674 -568
rect 1708 -602 2300 -568
rect 2338 -582 2856 -564
rect 1588 -636 1622 -602
rect 1588 -670 1808 -636
rect 1842 -670 1858 -636
rect 1548 -788 1582 -772
rect 1440 -1254 1506 -1244
rect 1440 -1288 1456 -1254
rect 1490 -1288 1506 -1254
rect 1548 -1288 1582 -1164
rect 1644 -788 1678 -670
rect 1902 -704 1936 -602
rect 1836 -738 1936 -704
rect 2112 -684 2234 -668
rect 2112 -720 2118 -684
rect 2154 -720 2192 -684
rect 2228 -720 2234 -684
rect 2112 -736 2234 -720
rect 1644 -1180 1678 -1164
rect 1740 -788 1774 -772
rect 1740 -1288 1774 -1164
rect 1836 -788 1870 -738
rect 1836 -1180 1870 -1164
rect 1932 -788 1966 -772
rect 2338 -908 2406 -582
rect 2790 -824 2850 -814
rect 2790 -826 2862 -824
rect 2790 -862 2796 -826
rect 2832 -862 2862 -826
rect 2790 -874 2850 -862
rect 1932 -1288 1966 -1164
rect 2268 -976 2406 -908
rect 1440 -1298 1506 -1288
rect 1542 -1324 1566 -1288
rect 1602 -1324 1658 -1288
rect 1694 -1324 1750 -1288
rect 1786 -1324 1842 -1288
rect 1878 -1324 1934 -1288
rect 1970 -1324 1994 -1288
rect 1542 -1326 1994 -1324
rect 2268 -1326 2348 -976
rect 2896 -1248 2952 152
rect 2406 -1286 2952 -1248
rect 3994 -86 4192 360
rect 3994 -160 4052 -86
rect 4126 -160 4192 -86
rect 3994 -560 4192 -160
rect 3994 -634 4052 -560
rect 4126 -634 4192 -560
rect 3994 -1034 4192 -634
rect 3994 -1108 4052 -1034
rect 4126 -1108 4192 -1034
rect 3994 -1222 4192 -1108
rect 3994 -1256 4008 -1222
rect 4042 -1256 4080 -1222
rect 4114 -1256 4152 -1222
rect 4186 -1256 4192 -1222
rect 3994 -1294 4192 -1256
rect 2268 -1344 2632 -1326
rect 2268 -1346 2350 -1344
rect 2268 -1382 2276 -1346
rect 2312 -1380 2350 -1346
rect 2386 -1380 2430 -1344
rect 2466 -1380 2510 -1344
rect 2546 -1380 2590 -1344
rect 2626 -1380 2632 -1344
rect 2312 -1382 2632 -1380
rect 2268 -1396 2632 -1382
rect 3994 -1328 4008 -1294
rect 4042 -1328 4080 -1294
rect 4114 -1328 4152 -1294
rect 4186 -1328 4192 -1294
rect 3994 -1366 4192 -1328
rect 3994 -1400 4008 -1366
rect 4042 -1400 4080 -1366
rect 4114 -1400 4152 -1366
rect 4186 -1400 4192 -1366
rect 3994 -1438 4192 -1400
rect 3994 -1472 4008 -1438
rect 4042 -1472 4080 -1438
rect 4114 -1472 4152 -1438
rect 4186 -1472 4192 -1438
rect 1096 -1602 1214 -1586
rect 1096 -1668 1120 -1602
rect 1196 -1668 1214 -1602
rect 1096 -1680 1214 -1668
rect 3994 -1698 4192 -1472
rect -686 -1740 864 -1700
rect -686 -1814 -622 -1740
rect -548 -1806 -354 -1740
rect -290 -1806 -220 -1740
rect -156 -1806 -86 -1740
rect -22 -1806 22 -1740
rect 86 -1806 130 -1740
rect 194 -1806 238 -1740
rect 302 -1806 346 -1740
rect 410 -1806 454 -1740
rect 518 -1806 562 -1740
rect 626 -1806 670 -1740
rect 734 -1806 778 -1740
rect 842 -1806 864 -1740
rect -548 -1814 864 -1806
rect -686 -1828 864 -1814
rect 2028 -1738 4192 -1698
rect 2028 -1804 2056 -1738
rect 2120 -1804 2164 -1738
rect 2228 -1804 2272 -1738
rect 2336 -1804 2380 -1738
rect 2444 -1804 2488 -1738
rect 2552 -1804 2596 -1738
rect 2660 -1804 2704 -1738
rect 2768 -1804 2812 -1738
rect 2876 -1804 2920 -1738
rect 2984 -1804 3028 -1738
rect 3092 -1804 3136 -1738
rect 3200 -1804 3244 -1738
rect 3308 -1804 3356 -1738
rect 3420 -1804 3464 -1738
rect 3528 -1804 3572 -1738
rect 3642 -1770 4192 -1738
rect 3642 -1804 4052 -1770
rect 2028 -1826 4052 -1804
rect -686 -2214 -488 -1828
rect -686 -2288 -622 -2214
rect -548 -2288 -488 -2214
rect -686 -2688 -488 -2288
rect -686 -2762 -622 -2688
rect -548 -2762 -488 -2688
rect -686 -3164 -488 -2762
rect -686 -3238 -622 -3164
rect -548 -3238 -488 -3164
rect -686 -3638 -488 -3238
rect -686 -3712 -622 -3638
rect -548 -3712 -488 -3638
rect -686 -4112 -488 -3712
rect -686 -4186 -622 -4112
rect -548 -4186 -488 -4112
rect -686 -4586 -488 -4186
rect -686 -4660 -622 -4586
rect -548 -4660 -488 -4586
rect -686 -4932 -488 -4660
rect 3994 -1844 4052 -1826
rect 4126 -1844 4192 -1770
rect 3994 -2244 4192 -1844
rect 3994 -2318 4052 -2244
rect 4126 -2318 4192 -2244
rect 3994 -2718 4192 -2318
rect 3994 -2792 4052 -2718
rect 4126 -2792 4192 -2718
rect 3994 -3192 4192 -2792
rect 3994 -3266 4052 -3192
rect 4126 -3266 4192 -3192
rect 3994 -3666 4192 -3266
rect 3994 -3740 4052 -3666
rect 4126 -3740 4192 -3666
rect 3994 -4140 4192 -3740
rect 3994 -4214 4052 -4140
rect 4126 -4214 4192 -4140
rect 3994 -4614 4192 -4214
rect 3994 -4688 4054 -4614
rect 4128 -4688 4192 -4614
rect 3994 -4932 4192 -4688
rect -686 -5000 4192 -4932
rect -686 -5074 -92 -5000
rect -18 -5074 456 -5000
rect 530 -5074 1004 -5000
rect 1078 -5074 1552 -5000
rect 1626 -5074 2100 -5000
rect 2174 -5074 2648 -5000
rect 2722 -5074 3198 -5000
rect 3272 -5074 4192 -5000
rect -686 -5130 4192 -5074
<< viali >>
rect -156 406 -92 472
rect -48 406 16 472
rect 60 406 124 472
rect 168 406 232 472
rect 276 406 340 472
rect 384 406 448 472
rect 492 406 556 472
rect 600 406 664 472
rect 708 406 772 472
rect 950 348 1032 414
rect 112 66 146 100
rect 196 66 230 100
rect 280 66 314 100
rect 364 66 398 100
rect 448 66 482 100
rect 532 66 566 100
rect 616 66 650 100
rect 700 66 734 100
rect 784 66 818 100
rect 874 66 908 100
rect 276 -374 316 -334
rect 374 -400 410 -364
rect 668 -324 708 -284
rect -670 -1256 -636 -1222
rect -598 -1256 -564 -1222
rect -526 -1256 -492 -1222
rect -670 -1328 -636 -1294
rect -598 -1328 -564 -1294
rect -526 -1328 -492 -1294
rect 994 -656 1030 -620
rect 994 -730 1030 -694
rect -670 -1400 -636 -1366
rect -598 -1400 -564 -1366
rect -526 -1400 -492 -1366
rect 100 -1368 136 -1332
rect 218 -1368 254 -1332
rect 336 -1368 372 -1332
rect 454 -1368 490 -1332
rect 572 -1368 608 -1332
rect 690 -1368 726 -1332
rect 808 -1368 844 -1332
rect -670 -1472 -636 -1438
rect -598 -1472 -564 -1438
rect -526 -1472 -492 -1438
rect 968 -1668 1042 -1602
rect 1134 350 1204 416
rect 2042 406 2106 472
rect 2150 406 2214 472
rect 2258 408 2318 474
rect 2358 406 2422 472
rect 2468 406 2532 472
rect 2576 406 2640 472
rect 2682 406 2746 472
rect 2792 406 2856 472
rect 2900 406 2964 472
rect 3008 406 3072 472
rect 3116 406 3180 472
rect 3224 406 3288 472
rect 3336 406 3400 472
rect 3444 406 3508 472
rect 3552 406 3616 472
rect 2498 194 2534 230
rect 2574 194 2610 230
rect 2650 194 2686 230
rect 2726 194 2762 230
rect 2802 194 2838 230
rect 2878 194 2914 230
rect 1420 76 1454 110
rect 1504 76 1538 110
rect 1588 76 1622 110
rect 1672 76 1706 110
rect 1756 76 1790 110
rect 1840 76 1874 110
rect 1924 76 1958 110
rect 2008 76 2042 110
rect 1116 -404 1152 -368
rect 1116 -478 1152 -442
rect 2410 -240 2446 -206
rect 2410 -312 2446 -278
rect 2792 -272 2828 -236
rect 2118 -720 2154 -684
rect 2192 -720 2228 -684
rect 2796 -862 2832 -826
rect 1566 -1324 1602 -1288
rect 1658 -1324 1694 -1288
rect 1750 -1324 1786 -1288
rect 1842 -1324 1878 -1288
rect 1934 -1324 1970 -1288
rect 4008 -1256 4042 -1222
rect 4080 -1256 4114 -1222
rect 4152 -1256 4186 -1222
rect 2276 -1382 2312 -1346
rect 2350 -1380 2386 -1344
rect 2430 -1380 2466 -1344
rect 2510 -1380 2546 -1344
rect 2590 -1380 2626 -1344
rect 4008 -1328 4042 -1294
rect 4080 -1328 4114 -1294
rect 4152 -1328 4186 -1294
rect 4008 -1400 4042 -1366
rect 4080 -1400 4114 -1366
rect 4152 -1400 4186 -1366
rect 4008 -1472 4042 -1438
rect 4080 -1472 4114 -1438
rect 4152 -1472 4186 -1438
rect 1120 -1668 1196 -1602
rect -354 -1806 -290 -1740
rect -220 -1806 -156 -1740
rect -86 -1806 -22 -1740
rect 22 -1806 86 -1740
rect 130 -1806 194 -1740
rect 238 -1806 302 -1740
rect 346 -1806 410 -1740
rect 454 -1806 518 -1740
rect 562 -1806 626 -1740
rect 670 -1806 734 -1740
rect 778 -1806 842 -1740
rect 2056 -1804 2120 -1738
rect 2164 -1804 2228 -1738
rect 2272 -1804 2336 -1738
rect 2380 -1804 2444 -1738
rect 2488 -1804 2552 -1738
rect 2596 -1804 2660 -1738
rect 2704 -1804 2768 -1738
rect 2812 -1804 2876 -1738
rect 2920 -1804 2984 -1738
rect 3028 -1804 3092 -1738
rect 3136 -1804 3200 -1738
rect 3244 -1804 3308 -1738
rect 3356 -1804 3420 -1738
rect 3464 -1804 3528 -1738
rect 3572 -1804 3642 -1738
<< metal1 >>
rect -488 472 788 512
rect -488 406 -156 472
rect -92 406 -48 472
rect 16 406 60 472
rect 124 406 168 472
rect 232 406 276 472
rect 340 406 384 472
rect 448 406 492 472
rect 556 406 600 472
rect 664 406 708 472
rect 772 406 788 472
rect 2016 474 3974 512
rect 2016 472 2258 474
rect 2318 472 3974 474
rect -488 384 788 406
rect 938 414 1050 430
rect 938 348 950 414
rect 1032 348 1050 414
rect 938 328 1050 348
rect 1110 416 1222 432
rect 1110 350 1134 416
rect 1204 350 1222 416
rect 2016 406 2042 472
rect 2106 406 2150 472
rect 2214 406 2258 472
rect 2318 406 2358 472
rect 2424 406 2468 472
rect 2532 406 2576 472
rect 2640 406 2682 472
rect 2748 406 2792 472
rect 2856 406 2900 472
rect 2964 406 3008 472
rect 3076 406 3116 472
rect 3184 406 3224 472
rect 3292 406 3336 472
rect 3400 406 3444 472
rect 3508 406 3552 472
rect 3616 406 3974 472
rect 2016 384 3974 406
rect 1110 338 1222 350
rect -838 230 4360 300
rect -838 194 2498 230
rect 2534 194 2574 230
rect 2610 194 2650 230
rect 2686 194 2726 230
rect 2762 194 2802 230
rect 2838 194 2878 230
rect 2914 194 4360 230
rect -838 162 4360 194
rect 82 100 938 162
rect 82 66 112 100
rect 146 66 196 100
rect 230 66 280 100
rect 314 66 364 100
rect 398 66 448 100
rect 482 66 532 100
rect 566 66 616 100
rect 650 66 700 100
rect 734 66 784 100
rect 818 66 874 100
rect 908 66 938 100
rect 1382 110 2106 162
rect 1382 76 1420 110
rect 1454 76 1504 110
rect 1538 76 1588 110
rect 1622 76 1672 110
rect 1706 76 1756 110
rect 1790 76 1840 110
rect 1874 76 1924 110
rect 1958 76 2008 110
rect 2042 76 2106 110
rect 1382 70 2106 76
rect 82 60 938 66
rect 2396 -206 2452 -190
rect 2396 -240 2410 -206
rect 2446 -240 2452 -206
rect -838 -284 724 -268
rect -838 -296 668 -284
rect 652 -324 668 -296
rect 708 -324 724 -284
rect -838 -334 332 -324
rect 652 -334 724 -324
rect 2396 -278 2452 -240
rect 2396 -312 2410 -278
rect 2446 -312 2452 -278
rect 2786 -236 2846 -224
rect 2786 -272 2792 -236
rect 2828 -272 2846 -236
rect 2786 -284 2846 -272
rect 2396 -328 2452 -312
rect -838 -352 276 -334
rect 260 -374 276 -352
rect 316 -374 332 -334
rect 260 -384 332 -374
rect 362 -362 416 -358
rect 362 -364 1164 -362
rect 362 -400 374 -364
rect 410 -368 1164 -364
rect 410 -400 1116 -368
rect 362 -402 1116 -400
rect 362 -406 416 -402
rect 1104 -404 1116 -402
rect 1152 -404 1164 -368
rect 1104 -442 1164 -404
rect 1104 -478 1116 -442
rect 1152 -478 1164 -442
rect 1104 -484 1164 -478
rect 982 -620 1042 -614
rect 982 -656 994 -620
rect 1030 -656 1042 -620
rect 982 -694 1042 -656
rect 982 -730 994 -694
rect 1030 -700 1042 -694
rect 2108 -684 2238 -668
rect 2108 -700 2118 -684
rect 1030 -720 2118 -700
rect 2154 -720 2192 -684
rect 2228 -720 2238 -684
rect 1030 -730 2238 -720
rect 982 -736 2238 -730
rect 2790 -826 2850 -814
rect 2790 -862 2796 -826
rect 2832 -862 2850 -826
rect 2790 -874 2850 -862
rect -686 -1222 -486 -1202
rect -686 -1256 -670 -1222
rect -636 -1256 -598 -1222
rect -564 -1256 -526 -1222
rect -492 -1256 -486 -1222
rect -686 -1294 -486 -1256
rect 3994 -1222 4192 -1202
rect 3994 -1256 4008 -1222
rect 4042 -1256 4080 -1222
rect 4114 -1256 4152 -1222
rect 4186 -1256 4192 -1222
rect -686 -1326 -670 -1294
rect -838 -1328 -670 -1326
rect -636 -1328 -598 -1294
rect -564 -1328 -526 -1294
rect -492 -1326 -486 -1294
rect 1542 -1288 1994 -1282
rect 1542 -1324 1566 -1288
rect 1602 -1324 1658 -1288
rect 1694 -1324 1750 -1288
rect 1786 -1324 1842 -1288
rect 1878 -1324 1934 -1288
rect 1970 -1324 1994 -1288
rect 1542 -1326 1994 -1324
rect 3994 -1294 4192 -1256
rect 3994 -1326 4008 -1294
rect -492 -1328 4008 -1326
rect 4042 -1328 4080 -1294
rect 4114 -1328 4152 -1294
rect 4186 -1326 4192 -1294
rect 4186 -1328 4360 -1326
rect -838 -1332 4360 -1328
rect -838 -1366 100 -1332
rect -838 -1400 -670 -1366
rect -636 -1400 -598 -1366
rect -564 -1400 -526 -1366
rect -492 -1368 100 -1366
rect 136 -1368 218 -1332
rect 254 -1368 336 -1332
rect 372 -1368 454 -1332
rect 490 -1368 572 -1332
rect 608 -1368 690 -1332
rect 726 -1368 808 -1332
rect 844 -1344 4360 -1332
rect 844 -1346 2350 -1344
rect 844 -1368 2276 -1346
rect -492 -1382 2276 -1368
rect 2312 -1380 2350 -1346
rect 2386 -1380 2430 -1344
rect 2466 -1380 2510 -1344
rect 2546 -1380 2590 -1344
rect 2626 -1366 4360 -1344
rect 2626 -1380 4008 -1366
rect 2312 -1382 4008 -1380
rect -492 -1400 4008 -1382
rect 4042 -1400 4080 -1366
rect 4114 -1400 4152 -1366
rect 4186 -1400 4360 -1366
rect -838 -1438 4360 -1400
rect -838 -1472 -670 -1438
rect -636 -1472 -598 -1438
rect -564 -1472 -526 -1438
rect -492 -1472 4008 -1438
rect 4042 -1472 4080 -1438
rect 4114 -1472 4152 -1438
rect 4186 -1472 4360 -1438
rect -838 -1484 4360 -1472
rect 3994 -1498 4192 -1484
rect 942 -1602 1050 -1586
rect 942 -1668 968 -1602
rect 1042 -1668 1050 -1602
rect 942 -1680 1050 -1668
rect 1110 -1602 1214 -1586
rect 1110 -1668 1120 -1602
rect 1196 -1668 1214 -1602
rect 1110 -1680 1214 -1668
rect -380 -1740 864 -1700
rect -380 -1806 -354 -1740
rect -290 -1806 -220 -1740
rect -156 -1806 -86 -1740
rect -22 -1806 22 -1740
rect 86 -1806 130 -1740
rect 194 -1806 238 -1740
rect 302 -1806 346 -1740
rect 410 -1806 454 -1740
rect 518 -1806 562 -1740
rect 626 -1806 670 -1740
rect 734 -1806 778 -1740
rect 842 -1806 864 -1740
rect -380 -1828 864 -1806
rect 2030 -1738 3994 -1698
rect 2030 -1804 2056 -1738
rect 2120 -1804 2164 -1738
rect 2228 -1804 2272 -1738
rect 2336 -1804 2380 -1738
rect 2444 -1804 2488 -1738
rect 2552 -1804 2596 -1738
rect 2660 -1804 2704 -1738
rect 2768 -1804 2812 -1738
rect 2876 -1804 2920 -1738
rect 2984 -1804 3028 -1738
rect 3096 -1804 3136 -1738
rect 3204 -1804 3244 -1738
rect 3312 -1804 3356 -1738
rect 3420 -1804 3464 -1738
rect 3528 -1804 3572 -1738
rect 3642 -1804 3994 -1738
rect 2030 -1826 3994 -1804
<< via1 >>
rect -156 406 -92 472
rect -48 406 16 472
rect 60 406 124 472
rect 168 406 232 472
rect 276 406 340 472
rect 384 406 448 472
rect 492 406 556 472
rect 600 406 664 472
rect 708 406 772 472
rect 950 348 1032 414
rect 1134 350 1204 416
rect 2042 406 2106 472
rect 2150 406 2214 472
rect 2258 408 2318 472
rect 2258 406 2318 408
rect 2360 406 2422 472
rect 2422 406 2424 472
rect 2468 406 2532 472
rect 2576 406 2640 472
rect 2684 406 2746 472
rect 2746 406 2748 472
rect 2792 406 2856 472
rect 2900 406 2964 472
rect 3008 406 3072 472
rect 3072 406 3076 472
rect 3116 406 3180 472
rect 3180 406 3184 472
rect 3224 406 3288 472
rect 3288 406 3292 472
rect 3336 406 3400 472
rect 3444 406 3508 472
rect 3552 406 3616 472
rect 968 -1668 1042 -1602
rect 1120 -1668 1196 -1602
rect -354 -1806 -290 -1740
rect -220 -1806 -156 -1740
rect -86 -1806 -22 -1740
rect 22 -1806 86 -1740
rect 130 -1806 194 -1740
rect 238 -1806 302 -1740
rect 346 -1806 410 -1740
rect 454 -1806 518 -1740
rect 562 -1806 626 -1740
rect 670 -1806 734 -1740
rect 778 -1806 842 -1740
rect 2056 -1804 2120 -1738
rect 2164 -1804 2228 -1738
rect 2272 -1804 2336 -1738
rect 2380 -1804 2444 -1738
rect 2488 -1804 2552 -1738
rect 2596 -1804 2660 -1738
rect 2704 -1804 2768 -1738
rect 2812 -1804 2876 -1738
rect 2920 -1804 2984 -1738
rect 3028 -1804 3092 -1738
rect 3092 -1804 3096 -1738
rect 3136 -1804 3200 -1738
rect 3200 -1804 3204 -1738
rect 3244 -1804 3308 -1738
rect 3308 -1804 3312 -1738
rect 3356 -1804 3420 -1738
rect 3464 -1804 3528 -1738
rect 3572 -1804 3642 -1738
<< metal2 >>
rect -488 472 788 512
rect -488 406 -156 472
rect -92 406 -48 472
rect 16 406 60 472
rect 124 406 168 472
rect 232 406 276 472
rect 340 406 384 472
rect 448 406 492 472
rect 556 406 600 472
rect 664 406 708 472
rect 772 406 788 472
rect 2016 472 3974 512
rect -488 384 788 406
rect 938 414 1050 430
rect 938 348 950 414
rect 1032 348 1050 414
rect 938 328 1050 348
rect 1110 416 1222 432
rect 1110 350 1134 416
rect 1204 350 1222 416
rect 2016 406 2042 472
rect 2106 406 2150 472
rect 2214 406 2258 472
rect 2318 406 2360 472
rect 2424 406 2468 472
rect 2532 406 2576 472
rect 2640 406 2684 472
rect 2748 406 2792 472
rect 2856 406 2900 472
rect 2964 406 3008 472
rect 3076 406 3116 472
rect 3184 406 3224 472
rect 3292 406 3336 472
rect 3400 406 3444 472
rect 3508 406 3552 472
rect 3616 406 3974 472
rect 2016 384 3974 406
rect 1110 338 1222 350
rect 942 -1602 1050 -1586
rect 942 -1668 968 -1602
rect 1042 -1668 1050 -1602
rect 942 -1680 1050 -1668
rect 1110 -1602 1214 -1586
rect 1110 -1668 1120 -1602
rect 1196 -1668 1214 -1602
rect 1110 -1680 1214 -1668
rect -380 -1740 864 -1700
rect -380 -1806 -354 -1740
rect -290 -1806 -220 -1740
rect -156 -1806 -86 -1740
rect -22 -1806 22 -1740
rect 86 -1806 130 -1740
rect 194 -1806 238 -1740
rect 302 -1806 346 -1740
rect 410 -1806 454 -1740
rect 518 -1806 562 -1740
rect 626 -1806 670 -1740
rect 734 -1806 778 -1740
rect 842 -1806 864 -1740
rect -380 -1828 864 -1806
rect 2030 -1738 3994 -1698
rect 2030 -1804 2056 -1738
rect 2120 -1804 2164 -1738
rect 2228 -1804 2272 -1738
rect 2336 -1804 2380 -1738
rect 2444 -1804 2488 -1738
rect 2552 -1804 2596 -1738
rect 2660 -1804 2704 -1738
rect 2768 -1804 2812 -1738
rect 2876 -1804 2920 -1738
rect 2984 -1804 3028 -1738
rect 3096 -1804 3136 -1738
rect 3204 -1804 3244 -1738
rect 3312 -1804 3356 -1738
rect 3420 -1804 3464 -1738
rect 3528 -1804 3572 -1738
rect 3642 -1804 3994 -1738
rect 2030 -1826 3994 -1804
<< via2 >>
rect -156 406 -92 472
rect -48 406 16 472
rect 60 406 124 472
rect 168 406 232 472
rect 276 406 340 472
rect 384 406 448 472
rect 492 406 556 472
rect 600 406 664 472
rect 708 406 772 472
rect 950 348 1032 414
rect 1134 350 1204 416
rect 2042 406 2106 472
rect 2150 406 2214 472
rect 2258 406 2318 472
rect 2360 406 2424 472
rect 2468 406 2532 472
rect 2576 406 2640 472
rect 2684 406 2748 472
rect 2792 406 2856 472
rect 2900 406 2964 472
rect 3008 406 3076 472
rect 3116 406 3184 472
rect 3224 406 3292 472
rect 3336 406 3400 472
rect 3444 406 3508 472
rect 3552 406 3616 472
rect 968 -1668 1042 -1602
rect 1120 -1668 1196 -1602
rect -354 -1806 -290 -1740
rect -220 -1806 -156 -1740
rect -86 -1806 -22 -1740
rect 22 -1806 86 -1740
rect 130 -1806 194 -1740
rect 238 -1806 302 -1740
rect 346 -1806 410 -1740
rect 454 -1806 518 -1740
rect 562 -1806 626 -1740
rect 670 -1806 734 -1740
rect 778 -1806 842 -1740
rect 2056 -1804 2120 -1738
rect 2164 -1804 2228 -1738
rect 2272 -1804 2336 -1738
rect 2380 -1804 2444 -1738
rect 2488 -1804 2552 -1738
rect 2596 -1804 2660 -1738
rect 2704 -1804 2768 -1738
rect 2812 -1804 2876 -1738
rect 2920 -1804 2984 -1738
rect 3028 -1804 3096 -1738
rect 3136 -1804 3204 -1738
rect 3244 -1804 3312 -1738
rect 3356 -1804 3420 -1738
rect 3464 -1804 3528 -1738
rect 3572 -1804 3642 -1738
<< metal3 >>
rect -488 472 788 512
rect -488 406 -156 472
rect -92 406 -48 472
rect 16 406 60 472
rect 124 406 168 472
rect 232 406 276 472
rect 340 406 384 472
rect 448 406 492 472
rect 556 406 600 472
rect 664 406 708 472
rect 772 406 788 472
rect 2016 472 3974 512
rect -488 382 788 406
rect 938 414 1050 430
rect 938 348 950 414
rect 1032 348 1050 414
rect 938 328 1050 348
rect 1110 416 1222 432
rect 1110 350 1134 416
rect 1204 350 1222 416
rect 2016 406 2042 472
rect 2106 406 2150 472
rect 2214 406 2258 472
rect 2318 406 2360 472
rect 2424 406 2468 472
rect 2532 406 2576 472
rect 2640 406 2684 472
rect 2748 406 2792 472
rect 2856 406 2900 472
rect 2964 406 3008 472
rect 3076 406 3116 472
rect 3184 406 3224 472
rect 3292 406 3336 472
rect 3400 406 3444 472
rect 3508 406 3552 472
rect 3616 406 3974 472
rect 2016 382 3974 406
rect 1110 338 1222 350
rect 942 -1602 1050 -1586
rect 942 -1668 968 -1602
rect 1042 -1668 1050 -1602
rect 942 -1680 1050 -1668
rect 1110 -1602 1214 -1586
rect 1110 -1668 1120 -1602
rect 1196 -1668 1214 -1602
rect 1110 -1680 1214 -1668
rect -380 -1740 864 -1700
rect -380 -1806 -354 -1740
rect -290 -1806 -220 -1740
rect -156 -1806 -86 -1740
rect -22 -1806 22 -1740
rect 86 -1806 130 -1740
rect 194 -1806 238 -1740
rect 302 -1806 346 -1740
rect 410 -1806 454 -1740
rect 518 -1806 562 -1740
rect 626 -1806 670 -1740
rect 734 -1806 778 -1740
rect 842 -1806 864 -1740
rect -380 -1828 864 -1806
rect 2030 -1738 3994 -1698
rect 2030 -1804 2056 -1738
rect 2120 -1804 2164 -1738
rect 2228 -1804 2272 -1738
rect 2336 -1804 2380 -1738
rect 2444 -1804 2488 -1738
rect 2552 -1804 2596 -1738
rect 2660 -1804 2704 -1738
rect 2768 -1804 2812 -1738
rect 2876 -1804 2920 -1738
rect 2984 -1804 3028 -1738
rect 3096 -1804 3136 -1738
rect 3204 -1804 3244 -1738
rect 3312 -1804 3356 -1738
rect 3420 -1804 3464 -1738
rect 3528 -1804 3572 -1738
rect 3642 -1804 3994 -1738
rect 2030 -1826 3994 -1804
rect 2029 -1828 3994 -1826
<< via3 >>
rect 950 348 1032 414
rect 1134 350 1204 416
rect 968 -1668 1042 -1602
rect 1120 -1668 1196 -1602
<< metal4 >>
rect 568 430 674 512
rect 2888 432 2992 548
rect 568 414 1050 430
rect 568 348 950 414
rect 1032 348 1050 414
rect 568 328 1050 348
rect 1110 416 2992 432
rect 1110 350 1134 416
rect 1204 350 2992 416
rect 1110 328 2992 350
rect 942 -1596 1050 -1586
rect 534 -1602 1050 -1596
rect 534 -1668 968 -1602
rect 1042 -1668 1050 -1602
rect 534 -1680 1050 -1668
rect 1110 -1596 1214 -1586
rect 1110 -1602 2960 -1596
rect 1110 -1668 1120 -1602
rect 1196 -1668 2960 -1602
rect 1110 -1680 2960 -1668
rect 534 -1832 640 -1680
rect 2854 -1834 2960 -1680
<< comment >>
rect 94 -58 126 -16
rect 290 -62 322 -20
rect 480 -64 512 -22
rect 672 -64 704 -22
rect 864 -62 896 -20
rect 1332 -350 1350 -146
rect 1554 -338 1574 -118
rect 1748 -366 1768 -146
rect 1942 -308 1962 -88
rect 2168 -350 2186 -146
rect 100 -752 132 -710
rect 288 -738 320 -696
rect 476 -736 508 -694
rect 680 -732 712 -690
rect 868 -724 900 -682
rect 1548 -1056 1576 -888
rect 1742 -1058 1770 -890
rect 1934 -1072 1962 -904
rect 192 -1140 224 -1098
rect 390 -1142 422 -1100
rect 578 -1140 610 -1098
rect 766 -1140 798 -1098
use adc_comp_buffer  adc_comp_buffer_0 ../adc_comp_buffer
timestamp 1661502601
transform 1 0 2448 0 1 -226
box -42 -326 408 452
use adc_comp_buffer  adc_comp_buffer_1
timestamp 1661502601
transform 1 0 2448 0 -1 -870
box -42 -326 408 452
use cap_64_92  cap_64_92_0
timestamp 1661518684
transform 1 0 1750 0 1 2042
box -2149 -1580 2210 1580
use cap_64_92  cap_64_92_1
timestamp 1661518684
transform 1 0 1717 0 -1 -3358
box -2149 -1580 2210 1580
<< labels >>
rlabel locali 1210 -602 1210 -568 7 bn
rlabel locali 2300 -602 2300 -568 3 bp
rlabel locali 2862 -862 2862 -824 3 outn
port 7 e
rlabel locali 2860 -272 2860 -234 3 outp
port 8 e
rlabel locali 574 -450 574 -418 7 on
rlabel locali 190 -450 190 -418 7 op
rlabel metal1 -838 -296 -838 -268 7 inp
port 5 w
rlabel metal1 -838 -352 -838 -324 7 inn
port 6 w
rlabel metal1 -838 -1484 -838 -1326 7 VSS
port 2 w
rlabel metal1 -838 162 -838 300 7 VDD
port 1 w
rlabel locali 1440 -1298 1440 -1244 7 nclk
port 10 w
rlabel locali -6 -1044 -6 -1014 7 clk
port 9 w
<< end >>
