* NGSPICE file created from adc_top.ext - technology: sky130A

.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VPWR VPB VNB
D0 VNB DIODE sky130_fd_pr__diode_pw2nd_05v5 pj=2.64e+06 area=4.347e+11
.ends

.subckt sky130_fd_sc_hd__decap_6 VPWR VGND VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=4.524e+11p pd=4.52e+06u as=0p ps=0u w=870000u l=1.97e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=2.86e+11p pd=3.24e+06u as=0p ps=0u w=550000u l=1.97e+06u
.ends

.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=4.524e+11p pd=4.52e+06u as=0p ps=0u w=870000u l=4.73e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=2.86e+11p pd=3.24e+06u as=0p ps=0u w=550000u l=4.73e+06u
.ends

.subckt sky130_fd_sc_hd__decap_8 VPWR VGND VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=4.524e+11p pd=4.52e+06u as=0p ps=0u w=870000u l=2.89e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=2.86e+11p pd=3.24e+06u as=0p ps=0u w=550000u l=2.89e+06u
.ends

.subckt sky130_fd_sc_hd__decap_4 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=4.524e+11p pd=4.52e+06u as=0p ps=0u w=870000u l=1.05e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=2.86e+11p pd=3.24e+06u as=0p ps=0u w=550000u l=1.05e+06u
.ends

.subckt sky130_fd_sc_hd__and3_1 VGND VPWR X B A C VNB VPB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=3.9785e+11p pd=4.05e+06u as=2.415e+11p ps=2.83e+06u w=420000u l=150000u
X1 VPWR C a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_181_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X3 VGND C a_181_47# VNB sky130_fd_pr__nfet_01v8 ad=2.633e+11p pd=2.28e+06u as=0p ps=0u w=420000u l=150000u
X4 a_27_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X6 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X7 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__and2_1 VPWR VGND X B A VNB VPB
X0 VPWR B a_59_75# VPB sky130_fd_pr__pfet_01v8_hvt ad=4.507e+11p pd=4.18e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X1 X a_59_75# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=4.75e+11p pd=2.95e+06u as=0p ps=0u w=1e+06u l=150000u
X2 VGND B a_145_75# VNB sky130_fd_pr__nfet_01v8 ad=2.236e+11p pd=2.08e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X3 a_59_75# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 X a_59_75# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X5 a_145_75# A a_59_75# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nor3_1 C Y A B VGND VPWR VNB VPB
X0 VPWR A a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1 a_193_297# B a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X2 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=3.445e+11p pd=3.66e+06u as=3.445e+11p ps=3.66e+06u w=650000u l=150000u
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_109_297# C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X5 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand2_1 Y B A VGND VPWR VNB VPB
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=5.2e+11p pd=5.04e+06u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1 Y A a_113_47# VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X2 a_113_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X3 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__o211a_1 C1 B1 A2 A1 X VGND VPWR VNB VPB
X0 VGND A1 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=3.8025e+11p pd=3.77e+06u as=4.55e+11p ps=4e+06u w=650000u l=150000u
X1 a_510_47# B1 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=2.275e+11p pd=2e+06u as=0p ps=0u w=650000u l=150000u
X2 a_79_21# C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=7.4e+11p pd=5.48e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=150000u
X3 VPWR B1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_79_21# A2 a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.25e+11p ps=2.65e+06u w=1e+06u l=150000u
X5 a_297_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_79_21# C1 a_510_47# VNB sky130_fd_pr__nfet_01v8 ad=1.95e+11p pd=1.9e+06u as=0p ps=0u w=650000u l=150000u
X7 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X8 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X9 a_215_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkbuf_1 VGND VPWR X A VNB VPB
X0 VPWR a_75_212# X VPB sky130_fd_pr__pfet_01v8_hvt ad=2.291e+11p pd=2.16e+06u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X1 a_75_212# A VGND VNB sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=1.508e+11p ps=1.62e+06u w=520000u l=150000u
X2 a_75_212# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X3 VGND a_75_212# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
.ends

.subckt sky130_fd_sc_hd__decap_3 VPWR VGND VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=4.524e+11p pd=4.52e+06u as=0p ps=0u w=870000u l=590000u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=2.86e+11p pd=3.24e+06u as=0p ps=0u w=550000u l=590000u
.ends

.subckt sky130_fd_sc_hd__inv_2 A Y VPWR VGND VNB VPB
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=5.2e+11p ps=5.04e+06u w=1e+06u l=150000u
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=3.38e+11p pd=3.64e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__a21o_4 A2 A1 X B1 VGND VPWR VNB VPB
X0 VGND B1 a_84_21# VNB sky130_fd_pr__nfet_01v8 ad=1.2675e+12p pd=1.04e+07u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u
X1 a_741_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=1.495e+11p pd=1.76e+06u as=0p ps=0u w=650000u l=150000u
X2 a_84_21# A1 a_741_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VGND A2 a_901_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X4 VPWR a_84_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=1.39e+12p pd=1.278e+07u as=5.6e+11p ps=5.12e+06u w=1e+06u l=150000u
X5 VPWR A2 a_483_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.195e+12p ps=1.039e+07u w=1e+06u l=150000u
X6 a_483_297# B1 a_84_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X7 X a_84_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=3.64e+11p pd=3.72e+06u as=0p ps=0u w=650000u l=150000u
X8 a_84_21# B1 a_483_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND a_84_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VPWR a_84_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_483_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VPWR A1 a_483_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VGND a_84_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 X a_84_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_84_21# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_483_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 X a_84_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 a_901_47# A1 a_84_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 X a_84_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__xnor2_4 Y B A VGND VPWR VNB VPB
X0 VGND A a_902_47# VNB sky130_fd_pr__nfet_01v8 ad=1.2155e+12p pd=1.284e+07u as=1.2285e+12p ps=1.288e+07u w=650000u l=150000u
X1 Y a_38_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1.37e+12p pd=1.274e+07u as=2.16e+12p ps=2.032e+07u w=1e+06u l=150000u
X2 a_38_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1.35e+12p pd=1.27e+07u as=0p ps=0u w=1e+06u l=150000u
X3 a_820_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=1.33e+12p pd=1.266e+07u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR a_38_297# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND A a_902_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND B a_902_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND B a_902_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 Y B a_820_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_38_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_38_297# B a_38_47# VNB sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=8.775e+11p ps=9.2e+06u w=650000u l=150000u
X11 VGND A a_38_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_902_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_820_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_902_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 VPWR A a_38_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 Y a_38_297# a_902_47# VNB sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u
X17 Y a_38_297# a_902_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 a_38_47# B a_38_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_38_47# B a_38_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 a_38_297# B a_38_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 a_38_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 VPWR B a_38_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 a_38_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 a_902_47# a_38_297# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 a_902_47# a_38_297# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 Y B a_820_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 a_38_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 a_820_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 VPWR A a_38_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 VGND A a_38_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X31 VPWR A a_820_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 a_902_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X33 a_820_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X34 Y a_38_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X35 a_902_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X36 a_38_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X37 VPWR A a_820_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X38 VPWR a_38_297# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X39 VPWR B a_38_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__a211o_2 X A2 A1 B1 C1 VGND VPWR VNB VPB
X0 a_79_21# A1 a_348_47# VNB sky130_fd_pr__nfet_01v8 ad=3.9975e+11p pd=3.83e+06u as=2.665e+11p ps=2.12e+06u w=650000u l=150000u
X1 a_79_21# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=7.8325e+11p ps=6.31e+06u w=650000u l=150000u
X2 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X3 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=9.1e+11p pd=7.82e+06u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X4 a_79_21# C1 a_585_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X5 VPWR A2 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.9e+11p ps=5.18e+06u w=1e+06u l=150000u
X6 a_299_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_585_297# B1 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_348_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__xnor2_1 VGND VPWR B Y A VNB VPB
X0 a_377_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=1.39e+12p ps=8.78e+06u w=1e+06u l=150000u
X1 a_47_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X2 a_129_47# B a_47_47# VNB sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.72e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X3 a_285_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=3.445e+11p pd=3.66e+06u as=3.445e+11p ps=3.66e+06u w=650000u l=150000u
X4 Y a_47_47# a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=1.95e+11p pd=1.9e+06u as=0p ps=0u w=650000u l=150000u
X5 VGND A a_129_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR A a_47_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR a_47_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X8 Y B a_377_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_285_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__xor2_1 B X A VPWR VGND VNB VPB
X0 X a_35_297# a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=3e+11p pd=2.6e+06u as=5.3e+11p ps=5.06e+06u w=1e+06u l=150000u
X1 X B a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=5.005e+11p pd=2.84e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X2 a_35_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=5.525e+11p ps=5.6e+06u w=650000u l=150000u
X3 a_117_297# B a_35_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X4 VPWR B a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=5.3e+11p pd=5.06e+06u as=0p ps=0u w=1e+06u l=150000u
X5 VGND A a_35_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND a_35_297# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_285_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VPWR A a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_285_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nor4b_1 C B A D_N Y VGND VPWR VNB VPB
X0 Y a_91_199# VGND VNB sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=5.97e+11p ps=5.79e+06u w=650000u l=150000u
X1 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_91_199# D_N VGND VNB sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VPWR A a_341_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=2.915e+11p pd=2.67e+06u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X6 a_245_297# C a_161_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=3.3e+11p pd=2.66e+06u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X7 a_341_297# B a_245_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_91_199# D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X9 a_161_297# a_91_199# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.2e+11p ps=3.04e+06u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand2_2 Y A B VGND VPWR VNB VPB
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=7.9e+11p pd=7.58e+06u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=5.135e+11p pd=5.48e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X4 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X5 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__conb_1 LO HI VPB VNB VGND VPWR
R0 HI VPWR sky130_fd_pr__res_generic_po w=480000u l=45000u
R1 VGND LO sky130_fd_pr__res_generic_po w=480000u l=45000u
.ends

.subckt sky130_fd_sc_hd__a311o_1 A1 A2 X B1 C1 A3 VGND VPWR VNB VPB
X0 a_75_199# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=3.8025e+11p pd=3.77e+06u as=4.94e+11p ps=4.12e+06u w=650000u l=150000u
X1 a_208_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=2.5025e+11p pd=2.07e+06u as=0p ps=0u w=650000u l=150000u
X2 a_315_47# A2 a_208_47# VNB sky130_fd_pr__nfet_01v8 ad=3.38e+11p pd=2.34e+06u as=0p ps=0u w=650000u l=150000u
X3 VGND B1 a_75_199# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_75_199# A1 a_315_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_75_199# C1 a_544_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=4.15e+11p ps=2.83e+06u w=1e+06u l=150000u
X6 a_544_297# B1 a_201_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6.55e+11p ps=5.31e+06u w=1e+06u l=150000u
X7 VPWR a_75_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=8.95e+11p pd=5.79e+06u as=2.85e+11p ps=2.57e+06u w=1e+06u l=150000u
X8 a_201_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR A2 a_201_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_201_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VGND a_75_199# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand2b_2 B Y A_N VGND VPWR VNB VPB
X0 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=1.2386e+12p ps=8.57e+06u w=1e+06u l=150000u
X1 VGND A_N a_27_93# VNB sky130_fd_pr__nfet_01v8 ad=3.695e+11p pd=3.79e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X2 VGND B a_229_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.135e+11p ps=5.48e+06u w=650000u l=150000u
X3 Y a_27_93# a_229_47# VNB sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X4 a_229_47# a_27_93# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y a_27_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR a_27_93# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_229_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR A_N a_27_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__dfrtp_1 Q RESET_B D CLK VGND VPWR VNB VPB
X0 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X1 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X2 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.998e+11p ps=1.97e+06u w=360000u l=150000u
X3 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X4 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=1.449e+11p ps=1.53e+06u w=420000u l=150000u
X5 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=1.0617e+12p pd=9.62e+06u as=0p ps=0u w=420000u l=150000u
X6 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=1.2195e+12p ps=1.255e+07u w=1e+06u l=150000u
X7 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X8 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X9 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X10 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X11 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=2.583e+11p ps=2.37e+06u w=420000u l=150000u
X12 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X13 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X17 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X18 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X20 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X23 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X24 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X27 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nor2_1 B Y A VGND VPWR VNB VPB
X0 VPWR A a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=3.38e+11p pd=3.64e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X2 a_109_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X3 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__buf_2 VPWR VGND X A VNB VPB
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=5.63e+11p pd=5.18e+06u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X3 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=3.6625e+11p ps=3.78e+06u w=650000u l=150000u
X4 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__or3b_1 A C_N X B VGND VPWR VNB VPB
X0 a_109_93# C_N VGND VNB sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=4.231e+11p ps=4.71e+06u w=420000u l=150000u
X1 a_215_53# B VGND VNB sky130_fd_pr__nfet_01v8 ad=2.226e+11p pd=2.74e+06u as=0p ps=0u w=420000u l=150000u
X2 VGND a_109_93# a_215_53# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VGND A a_215_53# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VPWR A a_369_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=4.057e+11p pd=4.04e+06u as=1.365e+11p ps=1.49e+06u w=420000u l=150000u
X5 a_369_297# B a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X6 X a_215_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.75e+11p pd=2.55e+06u as=0p ps=0u w=1e+06u l=150000u
X7 a_297_297# a_109_93# a_215_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X8 a_109_93# C_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X9 X a_215_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.7875e+11p pd=1.85e+06u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__mux2_1 VGND VPWR S A1 A0 X VNB VPB
X0 VPWR a_505_21# a_535_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=4.553e+11p pd=4.29e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X1 a_505_21# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X2 a_218_374# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X3 VGND a_505_21# a_439_47# VNB sky130_fd_pr__nfet_01v8 ad=5.155e+11p pd=4.31e+06u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4 a_76_199# A0 a_218_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X5 a_505_21# S VGND VNB sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X6 a_439_47# A0 a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X7 a_535_374# A1 a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_76_199# A1 a_218_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X9 a_218_47# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkinv_2 Y A VPWR VGND VNB VPB
X0 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=2.205e+11p ps=2.73e+06u w=420000u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=5.45e+11p pd=5.09e+06u as=5.45e+11p ps=5.09e+06u w=1e+06u l=150000u
X2 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__a211oi_1 A1 C1 B1 Y A2 VPWR VGND VNB VPB
X0 a_56_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=5.45e+11p pd=5.09e+06u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X1 VPWR A2 a_56_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=3.5425e+11p pd=3.69e+06u as=4.68e+11p ps=4.04e+06u w=650000u l=150000u
X3 a_139_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X4 a_311_297# B1 a_56_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=3.1e+11p pd=2.62e+06u as=0p ps=0u w=1e+06u l=150000u
X5 Y C1 a_311_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=0p ps=0u w=1e+06u l=150000u
X6 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Y A1 a_139_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o21a_1 X A1 B1 A2 VGND VPWR VNB VPB
X0 VPWR A1 a_382_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=9.15e+11p pd=5.83e+06u as=3.05e+11p ps=2.61e+06u w=1e+06u l=150000u
X1 a_297_47# B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=3.705e+11p pd=3.74e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X2 a_297_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.445e+11p ps=3.66e+06u w=650000u l=150000u
X3 VGND A2 a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X5 a_79_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=3.9e+11p pd=2.78e+06u as=0p ps=0u w=1e+06u l=150000u
X6 a_382_297# A2 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o2111a_1 X D1 C1 B1 A2 A1 VPWR VGND VNB VPB
X0 a_676_297# A2 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=8.6e+11p ps=5.72e+06u w=1e+06u l=150000u
X1 a_512_47# B1 a_409_47# VNB sky130_fd_pr__nfet_01v8 ad=5.6875e+11p pd=4.35e+06u as=2.3725e+11p ps=2.03e+06u w=650000u l=150000u
X2 a_306_47# D1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=2.3725e+11p pd=2.03e+06u as=1.9825e+11p ps=1.91e+06u w=650000u l=150000u
X3 VGND A2 a_512_47# VNB sky130_fd_pr__nfet_01v8 ad=3.445e+11p pd=3.66e+06u as=0p ps=0u w=650000u l=150000u
X4 VPWR C1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=1.64e+12p pd=9.28e+06u as=0p ps=0u w=1e+06u l=150000u
X5 a_79_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR A1 a_676_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_512_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_409_47# C1 a_306_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X10 a_79_21# D1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__or4_1 C A X B D VPWR VGND VNB VPB
X0 a_27_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=2.52e+11p pd=2.88e+06u as=4.2635e+11p ps=4.72e+06u w=420000u l=150000u
X1 a_27_297# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_277_297# B a_205_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X3 VPWR A a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=2.965e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X4 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X5 a_205_297# C a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X6 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X7 VGND C a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_109_297# D a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X9 VGND A a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a21bo_1 X A1 B1_N A2 VGND VPWR VNB VPB
X0 a_298_297# a_27_413# a_215_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=5.35e+11p pd=5.07e+06u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X1 a_215_297# a_27_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=7.8855e+11p ps=5.09e+06u w=650000u l=150000u
X2 a_298_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6.492e+11p ps=6.44e+06u w=1e+06u l=150000u
X3 X a_215_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X4 VPWR B1_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X5 X a_215_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X6 a_382_47# A1 a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X7 VGND B1_N a_27_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.113e+11p ps=1.37e+06u w=420000u l=150000u
X8 VPWR A1 a_298_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND A2 a_382_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o221a_1 A2 X B1 C1 A1 B2 VGND VPWR VNB VPB
X0 a_240_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=3.445e+11p ps=3.66e+06u w=650000u l=150000u
X1 X a_51_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X2 VGND A1 a_240_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_51_297# B2 a_245_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=1.165e+12p pd=6.33e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X4 a_149_47# C1 a_51_297# VNB sky130_fd_pr__nfet_01v8 ad=3.6725e+11p pd=3.73e+06u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X5 a_240_47# B1 a_149_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR A1 a_512_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X7 X a_51_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u
X8 a_149_47# B2 a_240_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_245_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VPWR C1 a_51_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_512_297# A2 a_51_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__or3_1 A X B C VPWR VGND VNB VPB
X0 X a_29_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=2.965e+11p ps=2.68e+06u w=1e+06u l=150000u
X1 a_111_297# C a_29_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X2 X a_29_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=3.1715e+11p ps=3.36e+06u w=650000u l=150000u
X3 a_183_297# B a_111_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4 VPWR A a_183_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_29_53# B VGND VNB sky130_fd_pr__nfet_01v8 ad=2.226e+11p pd=2.74e+06u as=0p ps=0u w=420000u l=150000u
X6 VGND C a_29_53# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VGND A a_29_53# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nor2_2 B Y A VGND VPWR VNB VPB
X0 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=8.1e+11p ps=7.62e+06u w=1e+06u l=150000u
X1 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=5.265e+11p ps=5.52e+06u w=650000u l=150000u
X2 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__a31o_1 A2 B1 A1 A3 X VGND VPWR VNB VPB
X0 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=6.75e+11p pd=5.35e+06u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X1 a_209_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=6.5e+11p pd=5.3e+06u as=0p ps=0u w=1e+06u l=150000u
X2 a_303_47# A2 a_209_47# VNB sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=2.08e+11p ps=1.94e+06u w=650000u l=150000u
X3 a_209_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.3225e+11p ps=3.93e+06u w=650000u l=150000u
X4 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=150000u
X5 VGND B1 a_80_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.145e+11p ps=1.96e+06u w=650000u l=150000u
X6 a_80_21# A1 a_303_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR A2 a_209_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_80_21# B1 a_209_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=3.2e+11p pd=2.64e+06u as=0p ps=0u w=1e+06u l=150000u
X9 a_209_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 Y C1 B1 VGND VPWR VNB VPB
X0 a_110_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=6.55e+11p ps=5.31e+06u w=1e+06u l=150000u
X1 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=2.535e+11p pd=2.08e+06u as=4.2575e+11p ps=3.91e+06u w=650000u l=150000u
X2 Y A2 a_110_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=1.025e+12p pd=6.05e+06u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_326_47# B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.72e+06u as=0p ps=0u w=650000u l=150000u
X6 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 Y C1 a_326_47# VNB sky130_fd_pr__nfet_01v8 ad=3.9325e+11p pd=2.51e+06u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o22a_1 A2 X B1 A1 B2 VGND VPWR VNB VPB
X0 a_78_199# B1 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=150000u
X1 VPWR A1 a_493_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=1.005e+12p pd=6.01e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X2 a_493_297# A2 a_78_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.7e+11p ps=2.94e+06u w=1e+06u l=150000u
X3 VPWR a_78_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X4 VGND A2 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=3.445e+11p pd=3.66e+06u as=0p ps=0u w=650000u l=150000u
X5 a_78_199# B2 a_292_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.35e+11p ps=2.47e+06u w=1e+06u l=150000u
X6 a_215_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_215_47# B2 a_78_199# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_292_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND a_78_199# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a41o_1 VGND VPWR A3 A4 A2 X B1 A1 VNB VPB
X0 a_465_47# A2 a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X1 VGND A4 a_561_47# VNB sky130_fd_pr__nfet_01v8 ad=4.9075e+11p pd=4.11e+06u as=2.145e+11p ps=1.96e+06u w=650000u l=150000u
X2 VPWR A3 a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=8.6e+11p pd=7.72e+06u as=8.6e+11p ps=7.72e+06u w=1e+06u l=150000u
X3 a_297_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_297_297# A4 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR A1 a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_381_47# A1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.6725e+11p ps=2.43e+06u w=650000u l=150000u
X7 a_297_297# B1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X8 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X9 a_79_21# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X11 a_561_47# A3 a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a21o_1 A2 A1 B1 X VPWR VGND VNB VPB
X0 a_81_21# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=1.7875e+11p pd=1.85e+06u as=6.8575e+11p ps=4.71e+06u w=650000u l=150000u
X1 a_299_297# B1 a_81_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X2 VPWR a_81_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X3 VPWR A1 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND a_81_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X5 VGND A2 a_384_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X6 a_299_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_384_47# A1 a_81_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o21bai_1 A1 Y B1_N A2 VPWR VGND VNB VPB
X0 a_388_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=2.55e+11p pd=2.51e+06u as=3.05e+11p ps=2.61e+06u w=1e+06u l=150000u
X1 a_105_352# B1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=2.847e+11p ps=3.2e+06u w=420000u l=150000u
X2 a_297_47# a_105_352# Y VNB sky130_fd_pr__nfet_01v8 ad=3.705e+11p pd=3.74e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X3 a_297_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR A1 a_388_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=6.365e+11p pd=5.36e+06u as=0p ps=0u w=1e+06u l=150000u
X5 VGND A2 a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR B1_N a_105_352# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X7 Y a_105_352# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__o311a_1 X A1 A2 A3 B1 C1 VGND VPWR VNB VPB
X0 a_585_47# B1 a_266_47# VNB sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.72e+06u as=4.7125e+11p ps=4.05e+06u w=650000u l=150000u
X1 VGND A2 a_266_47# VNB sky130_fd_pr__nfet_01v8 ad=6.7925e+11p pd=4.69e+06u as=0p ps=0u w=650000u l=150000u
X2 VPWR a_81_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=9.25e+11p pd=5.85e+06u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X3 a_81_21# C1 a_585_47# VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X4 VGND a_81_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X5 a_266_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=3.6e+11p pd=2.72e+06u as=0p ps=0u w=1e+06u l=150000u
X6 a_368_297# A2 a_266_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=4.2e+11p pd=2.84e+06u as=0p ps=0u w=1e+06u l=150000u
X7 a_266_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_266_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_81_21# A3 a_368_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=5.35e+11p pd=5.07e+06u as=0p ps=0u w=1e+06u l=150000u
X10 a_81_21# C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VPWR B1 a_81_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__o21a_2 A1 B1 A2 X VGND VPWR VNB VPB
X0 VPWR A1 a_470_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=1.325e+12p pd=8.65e+06u as=3.2e+11p ps=2.64e+06u w=1e+06u l=150000u
X1 a_79_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u
X2 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=5.4925e+11p pd=5.59e+06u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X3 VGND A2 a_384_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.5425e+11p ps=3.69e+06u w=650000u l=150000u
X4 a_470_297# A2 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.75e+11p ps=2.55e+06u w=1e+06u l=150000u
X6 a_384_47# B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=150000u
X7 a_384_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a21oi_1 A1 B1 Y A2 VPWR VGND VNB VPB
X0 a_199_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=1.9175e+11p pd=1.89e+06u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X1 a_113_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=5.45e+11p pd=5.09e+06u as=2.95e+11p ps=2.59e+06u w=1e+06u l=150000u
X2 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.445e+11p ps=3.66e+06u w=650000u l=150000u
X3 VPWR A1 a_113_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_113_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X5 VGND A2 a_199_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__inv_1 Y A VGND VPWR VNB VPB
X0 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
.ends

.subckt pfet_01v8_w500_l500_nf2 a_n29_0# a_129_0# a_n129_n26# w_n224_n36# a_n187_0#
+ a_29_n26#
X0 a_129_0# a_29_n26# a_n29_0# w_n224_n36# sky130_fd_pr__pfet_01v8 ad=1.45e+11p pd=1.58e+06u as=1.45e+11p ps=1.58e+06u w=500000u l=500000u
X1 a_n29_0# a_n129_n26# a_n187_0# w_n224_n36# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.45e+11p ps=1.58e+06u w=500000u l=500000u
.ends

.subckt sky130_fd_sc_hd__buf_4 VPWR VGND X A VNB VPB
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=8e+11p pd=7.6e+06u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=5.2e+11p ps=5.5e+06u w=650000u l=150000u
X5 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X9 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__dlymetal6s6s_1 VPWR VGND A X VNB VPB
X0 X a_629_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=5.82e+11p ps=5.85e+06u w=650000u l=150000u
X1 a_523_47# a_346_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X2 VGND a_240_47# a_346_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X3 a_240_47# a_63_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X4 VPWR a_240_47# a_346_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=8.445e+11p pd=7.95e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X5 VGND A a_63_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X6 VPWR A a_63_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X7 VPWR a_523_47# a_629_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X8 VGND a_523_47# a_629_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X9 a_523_47# a_346_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X10 a_240_47# a_63_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X11 X a_629_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt adc_noise_decoup_cell1 nmoscap_top nmoscap_bot mimcap_top mimcap_bot pwell
X0 mimcap_top mimcap_bot sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X1 nmoscap_bot nmoscap_top nmoscap_bot pwell sky130_fd_pr__nfet_01v8 ad=2.296e+13p pd=6.84e+07u as=0p ps=0u w=1.64e+07u l=1.6e+07u
.ends

.subckt nfet_01v8_w500_l500_nf2 a_n129_n76# a_n29_n50# a_n187_n50# a_29_n76# a_129_n50#
+ VSUBS
X0 a_129_n50# a_29_n76# a_n29_n50# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45e+11p pd=1.58e+06u as=1.45e+11p ps=1.58e+06u w=500000u l=500000u
X1 a_n29_n50# a_n129_n76# a_n187_n50# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.45e+11p ps=1.58e+06u w=500000u l=500000u
.ends

.subckt adc_vcm_generator clk vcm VDD VSS
Xsky130_fd_sc_hd__inv_1_4 sky130_fd_sc_hd__inv_1_4/Y clk VSS VDD VSS VDD sky130_fd_sc_hd__inv_1
Xpfet_01v8_w500_l500_nf2_0 mimtop2 vcm phi1_n VDD vcm phi1_n pfet_01v8_w500_l500_nf2
Xpfet_01v8_w500_l500_nf2_1 mimtop1 vcm phi1_n VDD vcm phi1_n pfet_01v8_w500_l500_nf2
Xsky130_fd_sc_hd__buf_4_0 VDD VSS phi1_n sky130_fd_sc_hd__inv_1_0/Y VSS VDD sky130_fd_sc_hd__buf_4
Xpfet_01v8_w500_l500_nf2_2 mimbot1 VSS phi1_n VDD VSS phi1_n pfet_01v8_w500_l500_nf2
Xsky130_fd_sc_hd__buf_4_1 VDD VSS phi1 sky130_fd_sc_hd__inv_1_1/Y VSS VDD sky130_fd_sc_hd__buf_4
Xpfet_01v8_w500_l500_nf2_3 mimtop2 mimbot1 phi2_n VDD mimbot1 phi2_n pfet_01v8_w500_l500_nf2
Xsky130_fd_sc_hd__buf_4_2 VDD VSS phi2_n sky130_fd_sc_hd__inv_1_2/Y VSS VDD sky130_fd_sc_hd__buf_4
Xpfet_01v8_w500_l500_nf2_4 VDD mimtop1 phi2_n VDD mimtop1 phi2_n pfet_01v8_w500_l500_nf2
Xsky130_fd_sc_hd__buf_4_3 VDD VSS phi2 sky130_fd_sc_hd__inv_1_3/Y VSS VDD sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__dlymetal6s6s_1_0 VDD VSS sky130_fd_sc_hd__dlymetal6s6s_1_1/X sky130_fd_sc_hd__inv_1_1/A
+ VSS VDD sky130_fd_sc_hd__dlymetal6s6s_1
Xsky130_fd_sc_hd__dlymetal6s6s_1_1 VDD VSS sky130_fd_sc_hd__dlymetal6s6s_1_2/X sky130_fd_sc_hd__dlymetal6s6s_1_1/X
+ VSS VDD sky130_fd_sc_hd__dlymetal6s6s_1
Xsky130_fd_sc_hd__dlymetal6s6s_1_2 VDD VSS sky130_fd_sc_hd__nand2_1_0/Y sky130_fd_sc_hd__dlymetal6s6s_1_2/X
+ VSS VDD sky130_fd_sc_hd__dlymetal6s6s_1
Xsky130_fd_sc_hd__dlymetal6s6s_1_3 VDD VSS sky130_fd_sc_hd__dlymetal6s6s_1_4/X sky130_fd_sc_hd__inv_1_3/A
+ VSS VDD sky130_fd_sc_hd__dlymetal6s6s_1
Xsky130_fd_sc_hd__dlymetal6s6s_1_4 VDD VSS sky130_fd_sc_hd__dlymetal6s6s_1_5/X sky130_fd_sc_hd__dlymetal6s6s_1_4/X
+ VSS VDD sky130_fd_sc_hd__dlymetal6s6s_1
Xsky130_fd_sc_hd__dlymetal6s6s_1_5 VDD VSS sky130_fd_sc_hd__nand2_1_1/Y sky130_fd_sc_hd__dlymetal6s6s_1_5/X
+ VSS VDD sky130_fd_sc_hd__dlymetal6s6s_1
Xadc_noise_decoup_cell1_0[0|0] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_0[1|0] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_0[2|0] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_0[3|0] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_0[4|0] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_0[5|0] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_0[6|0] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_0[7|0] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_0[0|1] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_0[1|1] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_0[2|1] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_0[3|1] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_0[4|1] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_0[5|1] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_0[6|1] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_0[7|1] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_0[0|2] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_0[1|2] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_0[2|2] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_0[3|2] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_0[4|2] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_0[5|2] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_0[6|2] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_0[7|2] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_0[0|3] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_0[1|3] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_0[2|3] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_0[3|3] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_0[4|3] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_0[5|3] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_0[6|3] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_0[7|3] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_0[0|4] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_0[1|4] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_0[2|4] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_0[3|4] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_0[4|4] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_0[5|4] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_0[6|4] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_0[7|4] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[0] VDD VSS VDD VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[1] VDD VSS VDD VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[2] VDD VSS VDD VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_2[0|0] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_2[1|0] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_2[2|0] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_2[3|0] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_2[4|0] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_2[5|0] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_2[6|0] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_2[7|0] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_2[0|1] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_2[1|1] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_2[2|1] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_2[3|1] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_2[4|1] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_2[5|1] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_2[6|1] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_2[7|1] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_2[0|2] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_2[1|2] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_2[2|2] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_2[3|2] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_2[4|2] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_2[5|2] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_2[6|2] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_2[7|2] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_2[0|3] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_2[1|3] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_2[2|3] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_2[3|3] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_2[4|3] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_2[5|3] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_2[6|3] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_2[7|3] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_2[0|4] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_2[1|4] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_2[2|4] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_2[3|4] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_2[4|4] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_2[5|4] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_2[6|4] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_2[7|4] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xnfet_01v8_w500_l500_nf2_0 phi1 mimtop2 vcm phi1 vcm VSS nfet_01v8_w500_l500_nf2
Xnfet_01v8_w500_l500_nf2_1 phi1 mimtop1 vcm phi1 vcm VSS nfet_01v8_w500_l500_nf2
Xsky130_fd_sc_hd__nand2_1_0 sky130_fd_sc_hd__nand2_1_0/Y sky130_fd_sc_hd__inv_1_2/Y
+ clk VSS VDD VSS VDD sky130_fd_sc_hd__nand2_1
Xnfet_01v8_w500_l500_nf2_2 phi1 mimbot1 VSS phi1 VSS VSS nfet_01v8_w500_l500_nf2
Xsky130_fd_sc_hd__nand2_1_1 sky130_fd_sc_hd__nand2_1_1/Y sky130_fd_sc_hd__inv_1_4/Y
+ sky130_fd_sc_hd__inv_1_0/Y VSS VDD VSS VDD sky130_fd_sc_hd__nand2_1
Xnfet_01v8_w500_l500_nf2_3 phi2 mimtop2 mimbot1 phi2 mimbot1 VSS nfet_01v8_w500_l500_nf2
Xnfet_01v8_w500_l500_nf2_4 phi2 VDD mimtop1 phi2 mimtop1 VSS nfet_01v8_w500_l500_nf2
Xsky130_fd_sc_hd__inv_1_1 sky130_fd_sc_hd__inv_1_1/Y sky130_fd_sc_hd__inv_1_1/A VSS
+ VDD VSS VDD sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_0 sky130_fd_sc_hd__inv_1_0/Y sky130_fd_sc_hd__inv_1_1/Y VSS
+ VDD VSS VDD sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_2 sky130_fd_sc_hd__inv_1_2/Y sky130_fd_sc_hd__inv_1_3/Y VSS
+ VDD VSS VDD sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_3 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__inv_1_3/A VSS
+ VDD VSS VDD sky130_fd_sc_hd__inv_1
.ends

.subckt sky130_fd_sc_hd__or2_1 A X B VGND VPWR VNB VPB
X0 VGND A a_68_297# VNB sky130_fd_pr__nfet_01v8 ad=3.097e+11p pd=3.33e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X1 a_68_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 X a_68_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X3 VPWR A a_150_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=2.915e+11p pd=2.67e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X4 X a_68_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=3.4e+11p pd=2.68e+06u as=0p ps=0u w=1e+06u l=150000u
X5 a_150_297# B a_68_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand2_4 Y A B VGND VPWR VNB VPB
X0 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=8.645e+11p pd=9.16e+06u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u
X1 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1.08e+12p pd=1.016e+07u as=1.33e+12p ps=1.266e+07u w=1e+06u l=150000u
X3 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u
X7 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__dfrtp_4 Q RESET_B D CLK VGND VPWR VNB VPB
X0 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X1 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X2 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.998e+11p ps=1.97e+06u w=360000u l=150000u
X3 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X4 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=1.449e+11p ps=1.53e+06u w=420000u l=150000u
X5 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=1.3795e+12p pd=1.312e+07u as=0p ps=0u w=420000u l=150000u
X6 VPWR a_1283_21# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=1.7533e+12p pd=1.756e+07u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X7 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X8 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X9 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VPWR a_1283_21# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X12 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u
X13 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X14 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=2.583e+11p ps=2.37e+06u w=420000u l=150000u
X15 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X16 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X20 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X21 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X24 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 VGND a_1283_21# Q VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 VGND a_1283_21# Q VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X27 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X29 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X30 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X31 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X32 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X33 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a22o_1 A1 A2 X B2 B1 VPWR VGND VNB VPB
X0 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=5.629e+11p pd=5.14e+06u as=5.9e+11p ps=5.18e+06u w=1e+06u l=150000u
X1 a_27_297# B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=3.38e+11p pd=3.64e+06u as=1.495e+11p ps=1.76e+06u w=650000u l=150000u
X2 VGND A2 a_373_47# VNB sky130_fd_pr__nfet_01v8 ad=3.705e+11p pd=3.74e+06u as=2.275e+11p ps=2e+06u w=650000u l=150000u
X3 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X4 a_27_297# B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=5.1285e+11p pd=5.04e+06u as=0p ps=0u w=1e+06u l=150000u
X5 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_373_47# A1 a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X8 a_109_297# B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_109_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand4_1 C B Y D A VPWR VGND VNB VPB
X0 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=8.3e+11p ps=7.66e+06u w=1e+06u l=150000u
X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_193_47# C a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X4 Y A a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=1.95e+11p pd=1.9e+06u as=2.145e+11p ps=1.96e+06u w=650000u l=150000u
X5 a_277_47# B a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_109_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__or4b_1 B D_N A X C VPWR VGND VNB VPB
X0 X a_215_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.75e+11p pd=2.55e+06u as=4.057e+11p ps=4.04e+06u w=1e+06u l=150000u
X1 a_109_53# D_N VGND VNB sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=5.3555e+11p ps=6.08e+06u w=420000u l=150000u
X2 a_215_297# a_109_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=2.415e+11p pd=2.83e+06u as=0p ps=0u w=420000u l=150000u
X3 X a_215_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.7875e+11p pd=1.85e+06u as=0p ps=0u w=650000u l=150000u
X4 a_392_297# C a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=9.03e+10p pd=1.27e+06u as=1.365e+11p ps=1.49e+06u w=420000u l=150000u
X5 a_465_297# B a_392_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=1.281e+11p pd=1.45e+06u as=0p ps=0u w=420000u l=150000u
X6 a_215_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VPWR A a_465_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_297_297# a_109_53# a_215_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X9 a_109_53# D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X10 VGND C a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VGND A a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a211o_1 VGND VPWR X A2 B1 A1 C1 VNB VPB
X0 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=5.45e+11p pd=5.09e+06u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X1 a_80_21# C1 a_472_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=2.65e+11p pd=2.53e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X2 VPWR A2 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.45e+11p ps=5.09e+06u w=1e+06u l=150000u
X3 VGND B1 a_80_21# VNB sky130_fd_pr__nfet_01v8 ad=7.215e+11p pd=4.82e+06u as=3.5425e+11p ps=3.69e+06u w=650000u l=150000u
X4 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=150000u
X5 a_300_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X6 a_217_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_80_21# A1 a_300_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_472_297# B1 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_80_21# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a32o_1 X A3 B2 B1 A1 A2 VGND VPWR VNB VPB
X0 a_93_21# A1 a_346_47# VNB sky130_fd_pr__nfet_01v8 ad=2.86e+11p pd=2.18e+06u as=2.925e+11p ps=2.2e+06u w=650000u l=150000u
X1 a_93_21# B1 a_250_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=9.65e+11p ps=7.93e+06u w=1e+06u l=150000u
X2 a_584_47# B1 a_93_21# VNB sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.72e+06u as=0p ps=0u w=650000u l=150000u
X3 VPWR a_93_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=9.35e+11p pd=5.87e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X4 VGND B2 a_584_47# VNB sky130_fd_pr__nfet_01v8 ad=5.07e+11p pd=4.16e+06u as=0p ps=0u w=650000u l=150000u
X5 a_256_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=1.95e+11p pd=1.9e+06u as=0p ps=0u w=650000u l=150000u
X6 a_250_297# B2 a_93_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND a_93_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.145e+11p ps=1.96e+06u w=650000u l=150000u
X8 a_250_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR A2 a_250_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_250_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_346_47# A2 a_256_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o21ai_1 VGND VPWR A2 A1 B1 Y VNB VPB
X0 Y A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=3.48e+11p pd=2.78e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X1 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=4.42e+11p pd=4.44e+06u as=0p ps=0u w=700000u l=150000u
X2 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=3.445e+11p pd=3.66e+06u as=2.145e+11p ps=1.96e+06u w=650000u l=150000u
X3 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X4 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a31o_2 X B1 A3 A1 A2 VGND VPWR VNB VPB
X0 VPWR A2 a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=8.6e+11p pd=7.72e+06u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X1 a_277_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_79_21# B1 a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=3.2e+11p pd=2.64e+06u as=0p ps=0u w=1e+06u l=150000u
X3 a_277_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X5 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=5.135e+11p pd=5.48e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X6 a_361_47# A2 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X7 a_277_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VGND B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.535e+11p ps=2.08e+06u w=650000u l=150000u
X9 a_79_21# A1 a_361_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__and2b_1 X A_N B VGND VPWR VNB VPB
X0 VPWR B a_207_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=5.986e+11p pd=5e+06u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X1 X a_207_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X2 a_297_47# a_27_413# a_207_413# VNB sky130_fd_pr__nfet_01v8 ad=1.008e+11p pd=1.32e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X3 X a_207_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=3.118e+11p ps=3.34e+06u w=650000u l=150000u
X4 a_207_413# a_27_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VPWR A_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X6 VGND B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_27_413# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__buf_1 VGND VPWR X A VNB VPB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=2.291e+11p pd=2.16e+06u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X1 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=1.508e+11p ps=1.62e+06u w=520000u l=150000u
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X3 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
.ends

.subckt sky130_fd_sc_hd__and4_1 X C A B D VGND VPWR VNB VPB
X0 a_27_47# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.646e+11p pd=2.94e+06u as=8.895e+11p ps=6.3e+06u w=420000u l=150000u
X1 a_197_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=1.596e+11p pd=1.6e+06u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X3 a_303_47# C a_197_47# VNB sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VPWR D a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VGND D a_303_47# VNB sky130_fd_pr__nfet_01v8 ad=3.9255e+11p pd=2.66e+06u as=0p ps=0u w=420000u l=150000u
X7 VPWR B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X9 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkbuf_2 A X VGND VPWR VNB VPB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=5.85e+11p pd=5.17e+06u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X1 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X2 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=2.457e+11p pd=2.85e+06u as=1.113e+11p ps=1.37e+06u w=420000u l=150000u
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X5 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand3_4 Y A B C VGND VPWR VNB VPB
X0 a_27_47# B a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=8.645e+11p pd=9.16e+06u as=8.71e+11p ps=9.18e+06u w=650000u l=150000u
X1 a_27_47# B a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1.62e+12p pd=1.524e+07u as=2.13e+12p ps=2.026e+07u w=1e+06u l=150000u
X3 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 Y A a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u
X5 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 Y A a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_27_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u
X9 a_27_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_445_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_445_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VGND C a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_445_47# B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_445_47# B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VGND C a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nor4_4 A C Y D B VGND VPWR VNB VPB
X0 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=1.35e+12p ps=1.27e+07u w=1e+06u l=150000u
X1 a_807_297# D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=1.33e+12p pd=1.266e+07u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X2 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=1.9175e+12p pd=1.76e+07u as=1.404e+12p ps=1.472e+07u w=650000u l=150000u
X3 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 Y D a_807_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 Y C VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Y D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 Y C VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 Y D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_27_297# B a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.08e+12p ps=1.016e+07u w=1e+06u l=150000u
X12 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_449_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_807_297# C a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 VGND D Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 VGND D Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 a_807_297# C a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_449_297# C a_807_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 a_449_297# C a_807_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 a_27_297# B a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 a_807_297# D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 a_449_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 Y D a_807_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkbuf_4 X A VGND VPWR VNB VPB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=9.1e+11p pd=7.82e+06u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X1 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=3.801e+11p pd=4.33e+06u as=2.352e+11p ps=2.8e+06u w=420000u l=150000u
X2 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=5.6e+11p pd=5.12e+06u as=0p ps=0u w=1e+06u l=150000u
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.113e+11p ps=1.37e+06u w=420000u l=150000u
X6 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__a2bb2o_1 VGND VPWR B1 A1_N A2_N X B2 VNB VPB
X0 a_226_47# A2_N a_226_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=1.113e+11p pd=1.37e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X1 a_489_413# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.226e+11p pd=2.74e+06u as=4.469e+11p ps=4.25e+06u w=420000u l=150000u
X2 a_226_297# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VPWR B2 a_489_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_489_413# a_226_47# a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X5 a_76_199# a_226_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=6.266e+11p ps=5.69e+06u w=420000u l=150000u
X6 VGND B1 a_556_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X7 a_556_47# B2 a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VGND A2_N a_226_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X9 a_226_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__xnor2_2 VGND VPWR Y A B VNB VPB
X0 a_27_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=8.25e+11p pd=7.65e+06u as=1.35e+12p ps=1.27e+07u w=1e+06u l=150000u
X1 a_560_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=5.4925e+11p pd=5.59e+06u as=7.02e+11p ps=7.36e+06u w=650000u l=150000u
X2 VGND B a_560_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y B a_474_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=5.75e+11p pd=5.15e+06u as=8.1e+11p ps=7.62e+06u w=1e+06u l=150000u
X4 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.3625e+11p ps=5.55e+06u w=650000u l=150000u
X5 Y a_27_297# a_560_47# VNB sky130_fd_pr__nfet_01v8 ad=3.38e+11p pd=3.64e+06u as=0p ps=0u w=650000u l=150000u
X6 a_474_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND A a_560_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_27_47# B a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X9 a_27_297# B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_27_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_474_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_560_47# a_27_297# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VPWR A a_474_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 Y a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VPWR a_27_297# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_560_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__dfrtp_2 Q RESET_B D CLK VGND VPWR VNB VPB
X0 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X1 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X2 VGND a_1283_21# Q VNB sky130_fd_pr__nfet_01v8 ad=1.2307e+12p pd=1.144e+07u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X3 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.998e+11p ps=1.97e+06u w=360000u l=150000u
X4 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X5 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=1.449e+11p ps=1.53e+06u w=420000u l=150000u
X6 VPWR a_1283_21# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=1.4795e+12p pd=1.507e+07u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X7 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X10 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X11 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X12 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X13 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=2.583e+11p ps=2.37e+06u w=420000u l=150000u
X14 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X15 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X19 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X20 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X22 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X26 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X27 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X29 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
.ends

.subckt sky130_fd_sc_hd__and3_2 B X A C VPWR VGND VNB VPB
X0 VPWR a_29_311# X VPB sky130_fd_pr__pfet_01v8_hvt ad=6.749e+11p pd=6.59e+06u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1 X a_29_311# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR A a_29_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.5795e+11p ps=2.99e+06u w=420000u l=150000u
X3 VGND a_29_311# X VNB sky130_fd_pr__nfet_01v8 ad=4.3955e+11p pd=4.06e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X4 a_184_53# B a_112_53# VNB sky130_fd_pr__nfet_01v8 ad=1.071e+11p pd=1.35e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X5 VPWR C a_29_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 X a_29_311# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_112_53# A a_29_311# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X8 a_29_311# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 VGND C a_184_53# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand3b_2 Y C A_N B VGND VPWR VNB VPB
X0 a_408_47# B a_218_47# VNB sky130_fd_pr__nfet_01v8 ad=5.135e+11p pd=5.48e+06u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u
X1 a_408_47# a_27_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X2 Y a_27_47# a_408_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=1.4015e+12p pd=1.289e+07u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X4 VGND C a_218_47# VNB sky130_fd_pr__nfet_01v8 ad=4.085e+11p pd=3.91e+06u as=0p ps=0u w=650000u l=150000u
X5 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.1e+11p ps=7.62e+06u w=1e+06u l=150000u
X6 a_218_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_218_47# B a_408_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 Y a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o21ba_1 B1_N A1 X A2 VGND VPWR VNB VPB
X0 a_222_93# B1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=3.76e+11p ps=3.81e+06u w=420000u l=150000u
X1 VPWR A1 a_544_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=9.515e+11p pd=7.99e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X2 VGND a_79_199# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X3 a_222_93# B1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X4 VGND A2 a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.8675e+11p ps=3.79e+06u w=650000u l=150000u
X5 a_448_47# a_222_93# a_79_199# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X6 a_79_199# a_222_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X7 a_544_297# A2 a_79_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_448_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR a_79_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__a21boi_4 Y A1 B1_N A2 VGND VPWR VNB VPB
X0 a_223_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1.96e+12p pd=1.792e+07u as=1.395e+12p ps=1.279e+07u w=1e+06u l=150000u
X1 Y A1 a_658_47# VNB sky130_fd_pr__nfet_01v8 ad=7.28e+11p pd=7.44e+06u as=7.28e+11p ps=7.44e+06u w=650000u l=150000u
X2 VPWR B1_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X3 a_223_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 Y a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.18625e+12p ps=1.015e+07u w=650000u l=150000u
X5 VGND A2 a_658_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_223_297# a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.6e+11p ps=5.12e+06u w=1e+06u l=150000u
X7 Y a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR A2 a_223_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_658_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VPWR A1 a_223_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_223_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_658_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 Y a_27_47# a_223_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_223_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VPWR A2 a_223_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VPWR A1 a_223_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_658_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VGND B1_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.6975e+11p ps=2.13e+06u w=650000u l=150000u
X19 a_223_297# a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 a_658_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 VGND A2 a_658_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 VGND a_27_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 VGND a_27_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 Y A1 a_658_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 Y a_27_47# a_223_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__o21ai_2 B1 Y A2 A1 VGND VPWR VNB VPB
X0 VGND A2 a_29_47# VNB sky130_fd_pr__nfet_01v8 ad=4.355e+11p pd=3.94e+06u as=7.085e+11p ps=7.38e+06u w=650000u l=150000u
X1 Y B1 a_29_47# VNB sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X2 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=8.5e+11p pd=7.7e+06u as=5.6e+11p ps=5.12e+06u w=1e+06u l=150000u
X3 VPWR A1 a_112_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6.3e+11p ps=5.26e+06u w=1e+06u l=150000u
X4 a_29_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y A2 a_112_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND A1 a_29_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_112_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_112_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_29_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_29_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__mux4_1 S0 A1 X S1 A2 A0 A3 VGND VPWR VNB VPB
X0 a_277_47# a_247_21# a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=2.226e+11p pd=2.74e+06u as=2.184e+11p ps=2.72e+06u w=420000u l=150000u
X1 VGND S0 a_247_21# VNB sky130_fd_pr__nfet_01v8 ad=6.142e+11p pd=7.3e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X2 a_834_97# a_247_21# a_750_97# VNB sky130_fd_pr__nfet_01v8 ad=2.1715e+11p pd=2.72e+06u as=2.226e+11p ps=2.74e+06u w=420000u l=150000u
X3 VGND A3 a_668_97# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.171e+11p ps=2.72e+06u w=420000u l=150000u
X4 a_1290_413# S1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=7.039e+11p ps=8e+06u w=420000u l=150000u
X5 a_834_97# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_750_97# S0 a_757_363# VPB sky130_fd_pr__pfet_01v8_hvt ad=3.822e+11p pd=3.5e+06u as=2.171e+11p ps=2.72e+06u w=420000u l=150000u
X7 a_27_47# S0 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=2.184e+11p pd=2.72e+06u as=2.7965e+11p ps=3.21e+06u w=420000u l=150000u
X8 X a_1478_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X9 VPWR A1 a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 VPWR S0 a_247_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.083e+11p ps=1.36e+06u w=420000u l=150000u
X11 X a_1478_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X12 a_193_47# A0 VGND VNB sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X13 a_750_97# a_1290_413# a_1478_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.84175e+11p ps=1.98e+06u w=420000u l=150000u
X14 a_1478_413# S1 a_277_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_1290_413# S1 VGND VNB sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X16 a_277_47# a_247_21# a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 a_750_97# S0 a_668_97# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 a_923_363# a_247_21# a_750_97# VPB sky130_fd_pr__pfet_01v8_hvt ad=1.8025e+11p pd=1.99e+06u as=0p ps=0u w=420000u l=150000u
X19 a_757_363# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 VPWR A3 a_923_363# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 a_277_47# a_1290_413# a_1478_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.0205e+11p ps=2.57e+06u w=420000u l=150000u
X22 a_193_413# A0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.171e+11p pd=2.72e+06u as=0p ps=0u w=420000u l=150000u
X23 a_193_413# S0 a_277_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 a_1478_413# S1 a_750_97# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N X A2_N B2 B1 VPWR VGND VNB VPB
X0 a_206_369# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.58e+11p pd=2.36e+06u as=8.192e+11p ps=6.72e+06u w=420000u l=150000u
X1 a_206_369# A2_N a_205_47# VNB sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.323e+11p ps=1.47e+06u w=420000u l=150000u
X2 VGND B2 a_489_47# VNB sky130_fd_pr__nfet_01v8 ad=3.1065e+11p pd=3.34e+06u as=2.226e+11p ps=2.74e+06u w=420000u l=150000u
X3 a_585_369# B2 a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.344e+11p ps=1.48e+06u w=420000u l=150000u
X4 a_489_47# a_206_369# a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X5 a_489_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VPWR A2_N a_206_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_76_199# a_206_369# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_205_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X10 VPWR B1 a_585_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a21o_2 X B1 A1 A2 VGND VPWR VNB VPB
X0 VPWR a_80_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=8.45e+11p pd=7.69e+06u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X1 X a_80_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND a_80_199# X VNB sky130_fd_pr__nfet_01v8 ad=5.655e+11p pd=5.64e+06u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X3 a_386_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u
X4 X a_80_199# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_80_199# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=3.25e+11p pd=2.3e+06u as=0p ps=0u w=650000u l=150000u
X6 a_386_297# B1 a_80_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X7 a_458_47# A1 a_80_199# VNB sky130_fd_pr__nfet_01v8 ad=2.47e+11p pd=2.06e+06u as=0p ps=0u w=650000u l=150000u
X8 VPWR A1 a_386_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND A2 a_458_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand2b_1 Y A_N B VGND VPWR VNB VPB
X0 VGND A_N a_27_93# VNB sky130_fd_pr__nfet_01v8 ad=2.005e+11p pd=1.97e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X1 Y a_27_93# a_206_47# VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X2 a_206_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR a_27_93# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=5.565e+11p pd=5.2e+06u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X4 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR A_N a_27_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a21oi_2 B1 A2 A1 Y VGND VPWR VNB VPB
X0 VGND A2 a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=6.5975e+11p pd=5.93e+06u as=1.365e+11p ps=1.72e+06u w=650000u l=150000u
X1 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.575e+11p ps=3.7e+06u w=650000u l=150000u
X2 Y A1 a_114_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7875e+11p ps=1.85e+06u w=650000u l=150000u
X3 a_114_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=1.19e+12p pd=1.038e+07u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X5 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.5e+11p ps=5.1e+06u w=1e+06u l=150000u
X6 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_285_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a31oi_1 VGND VPWR Y B1 A2 A1 A3 VNB VPB
X0 Y A1 a_181_47# VNB sky130_fd_pr__nfet_01v8 ad=2.1125e+11p pd=1.95e+06u as=2.3725e+11p ps=2.03e+06u w=650000u l=150000u
X1 a_181_47# A2 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.365e+11p ps=1.72e+06u w=650000u l=150000u
X2 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=3.445e+11p pd=3.66e+06u as=0p ps=0u w=650000u l=150000u
X3 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=5.65e+11p pd=5.13e+06u as=5.95e+11p ps=5.19e+06u w=1e+06u l=150000u
X4 Y B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X5 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_109_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_109_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a21boi_1 Y A1 B1_N A2 VPWR VGND VNB VPB
X0 a_300_297# a_27_413# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=5.45e+11p pd=5.09e+06u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X1 VGND A2 a_384_47# VNB sky130_fd_pr__nfet_01v8 ad=3.76e+11p pd=3.81e+06u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X2 VPWR B1_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=3.913e+11p pd=3.93e+06u as=1.113e+11p ps=1.37e+06u w=420000u l=150000u
X3 Y a_27_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=2.86e+11p pd=2.18e+06u as=0p ps=0u w=650000u l=150000u
X4 VPWR A1 a_300_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_384_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND B1_N a_27_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.113e+11p ps=1.37e+06u w=420000u l=150000u
X7 a_300_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkbuf_8 X A VGND VPWR VNB VPB
X0 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=1.65e+12p pd=1.53e+07u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X1 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.12e+12p ps=1.024e+07u w=1e+06u l=150000u
X2 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=4.704e+11p pd=5.6e+06u as=6.951e+11p ps=8.35e+06u w=420000u l=150000u
X5 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X9 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt adc_array_wafflecap_dummy sample_n colon_n col_n sample vcom row_n ctop VDD
+ VSS
X0 VDD colon_n a_170_252# VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1 a_662_574# row_n VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2 a_170_252# col_n a_662_574# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3 a_566_252# colon_n a_170_252# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4 VSS col_n a_566_252# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5 a_566_252# row_n VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_262_252# sample_n a_170_252# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X7 vcom sample a_262_252# VSS sky130_fd_pr__nfet_01v8 ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X8 a_262_252# sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=2.48e+11p ps=2.22e+06u w=800000u l=150000u
X9 a_170_252# sample a_262_252# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
.ends

.subckt adc_array_wafflecap_drv ctop colon_n col_n vcom row_n sample_i sample_n_i
+ sample_n_o sample_o VDD VSS
X0 VSS sample_i sample_n_o VSS sky130_fd_pr__nfet_01v8 ad=5.208e+11p pd=5.84e+06u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1 sample_n_o sample_i VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VDD sample_i sample_n_o VDD sky130_fd_pr__pfet_01v8 ad=9.92e+11p pd=8.88e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3 sample_n_o sample_i VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4 sample_o sample_n_i VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5 VSS sample_n_i sample_o VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 sample_o sample_n_i VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7 VDD sample_n_i sample_o VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
.ends

.subckt adc_array_wafflecap_1 sample_n colon_n col_n sample vcom row_n en_n ctop VDD
+ VSS
X0 VDD en_n a_170_252# VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1 a_662_574# en_n VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2 a_170_252# en_n a_662_574# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3 a_566_252# en_n a_170_252# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4 VSS en_n a_566_252# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5 a_566_252# en_n VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_262_252# sample_n a_170_252# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X7 vcom sample a_262_252# VSS sky130_fd_pr__nfet_01v8 ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X8 a_262_252# sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=2.48e+11p ps=2.22e+06u w=800000u l=150000u
X9 a_170_252# sample a_262_252# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
.ends

.subckt adc_array_wafflecap_8 sample_n colon_n col_n sample vcom row_n ctop VDD VSS
X0 VDD colon_n a_170_252# VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1 a_662_574# row_n VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2 a_170_252# col_n a_662_574# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3 a_566_252# colon_n a_170_252# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4 VSS col_n a_566_252# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5 a_566_252# row_n VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_262_252# sample_n a_170_252# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X7 vcom sample a_262_252# VSS sky130_fd_pr__nfet_01v8 ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X8 a_262_252# sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=2.48e+11p ps=2.22e+06u w=800000u l=150000u
X9 a_170_252# sample a_262_252# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
.ends

.subckt adc_array_wafflecap_4 sample_n colon_n col_n sample vcom row_n en_n ctop VDD
+ VSS
X0 VDD en_n a_170_252# VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1 a_662_574# en_n VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2 a_170_252# en_n a_662_574# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3 a_566_252# en_n a_170_252# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4 VSS en_n a_566_252# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5 a_566_252# en_n VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_262_252# sample_n a_170_252# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X7 vcom sample a_262_252# VSS sky130_fd_pr__nfet_01v8 ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X8 a_262_252# sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=2.48e+11p ps=2.22e+06u w=800000u l=150000u
X9 a_170_252# sample a_262_252# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
.ends

.subckt adc_array_wafflecap_2 sample_n colon_n col_n sample vcom row_n en_n ctop VDD
+ VSS
X0 VDD en_n a_170_252# VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1 a_662_574# en_n VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2 a_170_252# en_n a_662_574# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3 a_566_252# en_n a_170_252# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4 VSS en_n a_566_252# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5 a_566_252# en_n VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_262_252# sample_n a_170_252# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X7 vcom sample a_262_252# VSS sky130_fd_pr__nfet_01v8 ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X8 a_262_252# sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=2.48e+11p ps=2.22e+06u w=800000u l=150000u
X9 a_170_252# sample a_262_252# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
.ends

.subckt adc_array_wafflecap_gate sample_n colon_n col_n sample vcom row_n analog_in
+ sw sw_n a_169_51# VDD VSS li_854_970#
X0 a_169_51# sw_n analog_in VDD sky130_fd_pr__pfet_01v8 ad=2.7075e+12p pd=2.185e+07u as=1.102e+12p ps=8.76e+06u w=1.9e+06u l=220000u
X1 analog_in sw a_169_51# VSS sky130_fd_pr__nfet_01v8 ad=1.102e+12p pd=8.76e+06u as=2.7645e+12p ps=2.191e+07u w=1.9e+06u l=220000u
X2 analog_in sw_n a_169_51# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.9e+06u l=220000u
X3 a_169_51# sw_n analog_in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.9e+06u l=220000u
X4 a_169_51# sw_n a_169_51# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.9e+06u l=220000u
X5 a_169_51# sw analog_in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.9e+06u l=220000u
X6 a_169_51# sw analog_in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.9e+06u l=220000u
X7 a_169_51# sw a_169_51# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.9e+06u l=220000u
X8 analog_in sw a_169_51# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.9e+06u l=220000u
X9 a_169_51# sw a_169_51# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.9e+06u l=220000u
X10 a_169_51# sw_n a_169_51# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.9e+06u l=220000u
X11 analog_in sw_n a_169_51# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.9e+06u l=220000u
.ends

.subckt adc_array_matrix_12bit vcm sample sample_n row_n[15] row_n[14] row_n[13] row_n[12]
+ row_n[11] row_n[10] row_n[9] row_n[8] row_n[7] row_n[6] row_n[5] row_n[4] row_n[3]
+ row_n[2] row_n[1] row_n[0] rowon_n[15] rowon_n[14] rowon_n[13] rowon_n[12] rowon_n[11]
+ rowon_n[10] rowon_n[9] rowon_n[8] rowon_n[7] rowon_n[6] rowon_n[5] rowon_n[4] rowon_n[3]
+ rowon_n[2] rowon_n[1] rowon_n[0] col_n[31] col_n[30] col_n[29] col_n[28] col_n[27]
+ col_n[26] col_n[25] col_n[24] col_n[23] col_n[22] col_n[21] col_n[20] col_n[19]
+ col_n[18] col_n[17] col_n[16] col_n[15] col_n[14] col_n[13] col_n[12] col_n[11]
+ col_n[10] col_n[9] col_n[8] col_n[7] col_n[6] col_n[5] col_n[4] col_n[3] col_n[2]
+ col_n[1] col_n[0] en_bit_n[2] en_bit_n[1] en_bit_n[0] en_C0_n sw sw_n analog_in
+ ctop VSS VDD
Xadc_array_wafflecap_dummy_5[0] VDD VSS VSS VSS vcm col_n[2] adc_array_wafflecap_dummy_5[0]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_5[1] VDD VSS VSS VSS vcm col_n[3] adc_array_wafflecap_dummy_5[1]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_5[2] VDD VSS VSS VSS vcm col_n[4] adc_array_wafflecap_dummy_5[2]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_5[3] VDD VSS VSS VSS vcm col_n[5] adc_array_wafflecap_dummy_5[3]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_5[4] VDD VSS VSS VSS vcm col_n[6] adc_array_wafflecap_dummy_5[4]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_5[5] VDD VSS VSS VSS vcm col_n[7] adc_array_wafflecap_dummy_5[5]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_5[6] VDD VSS VSS VSS vcm col_n[8] adc_array_wafflecap_dummy_5[6]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_5[7] VDD VSS VSS VSS vcm col_n[9] adc_array_wafflecap_dummy_5[7]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_5[8] VDD VSS VSS VSS vcm col_n[10] adc_array_wafflecap_dummy_5[8]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_5[9] VDD VSS VSS VSS vcm col_n[11] adc_array_wafflecap_dummy_5[9]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_5[10] VDD VSS VSS VSS vcm col_n[12] adc_array_wafflecap_dummy_5[10]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_5[11] VDD VSS VSS VSS vcm col_n[13] adc_array_wafflecap_dummy_5[11]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_5[12] VDD VSS VSS VSS vcm col_n[14] adc_array_wafflecap_dummy_5[12]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_6[0] VDD VSS VSS VSS vcm VDD adc_array_wafflecap_dummy_6[0]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_6[1] VDD VSS VSS VSS vcm col_n[0] adc_array_wafflecap_dummy_6[1]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_drv_0[0] adc_array_wafflecap_drv_0[0]/ctop rowon_n[0] row_n[0]
+ vcm VDD sample sample_n adc_array_wafflecap_8_1[9]/sample_n adc_array_wafflecap_8_1[9]/sample
+ VDD VSS adc_array_wafflecap_drv
Xadc_array_wafflecap_drv_0[1] adc_array_wafflecap_drv_0[1]/ctop rowon_n[1] row_n[1]
+ vcm VDD sample sample_n adc_array_wafflecap_8_0[0|9]/sample_n adc_array_wafflecap_8_0[0|9]/sample
+ VDD VSS adc_array_wafflecap_drv
Xadc_array_wafflecap_drv_0[2] adc_array_wafflecap_drv_0[2]/ctop rowon_n[2] row_n[2]
+ vcm VDD sample sample_n adc_array_wafflecap_8_0[1|9]/sample_n adc_array_wafflecap_8_0[1|9]/sample
+ VDD VSS adc_array_wafflecap_drv
Xadc_array_wafflecap_drv_0[3] adc_array_wafflecap_drv_0[3]/ctop rowon_n[3] row_n[3]
+ vcm VDD sample sample_n adc_array_wafflecap_8_0[2|9]/sample_n adc_array_wafflecap_8_0[2|9]/sample
+ VDD VSS adc_array_wafflecap_drv
Xadc_array_wafflecap_drv_0[4] adc_array_wafflecap_drv_0[4]/ctop rowon_n[4] row_n[4]
+ vcm VDD sample sample_n adc_array_wafflecap_8_0[3|9]/sample_n adc_array_wafflecap_8_0[3|9]/sample
+ VDD VSS adc_array_wafflecap_drv
Xadc_array_wafflecap_drv_0[5] adc_array_wafflecap_drv_0[5]/ctop rowon_n[5] row_n[5]
+ vcm VDD sample sample_n adc_array_wafflecap_8_0[4|9]/sample_n adc_array_wafflecap_8_0[4|9]/sample
+ VDD VSS adc_array_wafflecap_drv
Xadc_array_wafflecap_drv_0[6] adc_array_wafflecap_drv_0[6]/ctop rowon_n[6] row_n[6]
+ vcm VDD sample sample_n adc_array_wafflecap_8_0[5|9]/sample_n adc_array_wafflecap_8_0[5|9]/sample
+ VDD VSS adc_array_wafflecap_drv
Xadc_array_wafflecap_drv_0[7] adc_array_wafflecap_drv_0[7]/ctop rowon_n[7] row_n[7]
+ vcm VDD sample sample_n adc_array_wafflecap_8_0[6|9]/sample_n adc_array_wafflecap_8_0[6|9]/sample
+ VDD VSS adc_array_wafflecap_drv
Xadc_array_wafflecap_drv_0[8] adc_array_wafflecap_drv_0[8]/ctop rowon_n[8] row_n[8]
+ vcm VDD sample sample_n adc_array_wafflecap_8_0[7|9]/sample_n adc_array_wafflecap_8_0[7|9]/sample
+ VDD VSS adc_array_wafflecap_drv
Xadc_array_wafflecap_drv_0[9] adc_array_wafflecap_drv_0[9]/ctop rowon_n[9] row_n[9]
+ vcm VDD sample sample_n adc_array_wafflecap_8_0[8|9]/sample_n adc_array_wafflecap_8_0[8|9]/sample
+ VDD VSS adc_array_wafflecap_drv
Xadc_array_wafflecap_drv_0[10] adc_array_wafflecap_drv_0[10]/ctop rowon_n[10] row_n[10]
+ vcm VDD sample sample_n adc_array_wafflecap_8_0[9|9]/sample_n adc_array_wafflecap_8_0[9|9]/sample
+ VDD VSS adc_array_wafflecap_drv
Xadc_array_wafflecap_drv_0[11] adc_array_wafflecap_drv_0[11]/ctop rowon_n[11] row_n[11]
+ vcm VDD sample sample_n adc_array_wafflecap_8_0[10|9]/sample_n adc_array_wafflecap_8_0[10|9]/sample
+ VDD VSS adc_array_wafflecap_drv
Xadc_array_wafflecap_drv_0[12] adc_array_wafflecap_drv_0[12]/ctop rowon_n[12] row_n[12]
+ vcm VDD sample sample_n adc_array_wafflecap_8_0[11|9]/sample_n adc_array_wafflecap_8_0[11|9]/sample
+ VDD VSS adc_array_wafflecap_drv
Xadc_array_wafflecap_drv_0[13] adc_array_wafflecap_drv_0[13]/ctop rowon_n[13] row_n[13]
+ vcm VDD sample sample_n adc_array_wafflecap_8_0[12|9]/sample_n adc_array_wafflecap_8_0[12|9]/sample
+ VDD VSS adc_array_wafflecap_drv
Xadc_array_wafflecap_drv_0[14] adc_array_wafflecap_drv_0[14]/ctop rowon_n[14] row_n[14]
+ vcm VDD sample sample_n adc_array_wafflecap_8_0[13|9]/sample_n adc_array_wafflecap_8_0[13|9]/sample
+ VDD VSS adc_array_wafflecap_drv
Xadc_array_wafflecap_drv_0[15] adc_array_wafflecap_drv_0[15]/ctop rowon_n[15] row_n[15]
+ vcm VDD sample sample_n adc_array_wafflecap_8_0[14|9]/sample_n adc_array_wafflecap_8_0[14|9]/sample
+ VDD VSS adc_array_wafflecap_drv
Xadc_array_wafflecap_1_0 VDD VSS VSS VSS vcm col_n[1] en_C0_n ctop VDD VSS adc_array_wafflecap_1
Xadc_array_wafflecap_1_1 VDD VSS VSS VSS vcm col_n[17] en_bit_n[0] ctop VDD VSS adc_array_wafflecap_1
Xadc_array_wafflecap_8_0[0|0] adc_array_wafflecap_8_0[0|9]/sample_n rowon_n[1] row_n[1]
+ adc_array_wafflecap_8_0[0|9]/sample vcm col_n[0] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|0] adc_array_wafflecap_8_0[1|9]/sample_n rowon_n[2] row_n[2]
+ adc_array_wafflecap_8_0[1|9]/sample vcm col_n[0] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|0] adc_array_wafflecap_8_0[2|9]/sample_n rowon_n[3] row_n[3]
+ adc_array_wafflecap_8_0[2|9]/sample vcm col_n[0] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|0] adc_array_wafflecap_8_0[3|9]/sample_n rowon_n[4] row_n[4]
+ adc_array_wafflecap_8_0[3|9]/sample vcm col_n[0] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|0] adc_array_wafflecap_8_0[4|9]/sample_n rowon_n[5] row_n[5]
+ adc_array_wafflecap_8_0[4|9]/sample vcm col_n[0] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|0] adc_array_wafflecap_8_0[5|9]/sample_n rowon_n[6] row_n[6]
+ adc_array_wafflecap_8_0[5|9]/sample vcm col_n[0] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|0] adc_array_wafflecap_8_0[6|9]/sample_n rowon_n[7] row_n[7]
+ adc_array_wafflecap_8_0[6|9]/sample vcm col_n[0] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|0] adc_array_wafflecap_8_0[7|9]/sample_n rowon_n[8] row_n[8]
+ adc_array_wafflecap_8_0[7|9]/sample vcm col_n[0] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|0] adc_array_wafflecap_8_0[8|9]/sample_n rowon_n[9] row_n[9]
+ adc_array_wafflecap_8_0[8|9]/sample vcm col_n[0] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|0] adc_array_wafflecap_8_0[9|9]/sample_n rowon_n[10] row_n[10]
+ adc_array_wafflecap_8_0[9|9]/sample vcm col_n[0] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|0] adc_array_wafflecap_8_0[10|9]/sample_n rowon_n[11]
+ row_n[11] adc_array_wafflecap_8_0[10|9]/sample vcm col_n[0] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|0] adc_array_wafflecap_8_0[11|9]/sample_n rowon_n[12]
+ row_n[12] adc_array_wafflecap_8_0[11|9]/sample vcm col_n[0] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|0] adc_array_wafflecap_8_0[12|9]/sample_n rowon_n[13]
+ row_n[13] adc_array_wafflecap_8_0[12|9]/sample vcm col_n[0] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|0] adc_array_wafflecap_8_0[13|9]/sample_n rowon_n[14]
+ row_n[14] adc_array_wafflecap_8_0[13|9]/sample vcm col_n[0] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|0] adc_array_wafflecap_8_0[14|9]/sample_n rowon_n[15]
+ row_n[15] adc_array_wafflecap_8_0[14|9]/sample vcm col_n[0] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|1] adc_array_wafflecap_8_0[0|9]/sample_n rowon_n[1] row_n[1]
+ adc_array_wafflecap_8_0[0|9]/sample vcm col_n[1] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|1] adc_array_wafflecap_8_0[1|9]/sample_n rowon_n[2] row_n[2]
+ adc_array_wafflecap_8_0[1|9]/sample vcm col_n[1] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|1] adc_array_wafflecap_8_0[2|9]/sample_n rowon_n[3] row_n[3]
+ adc_array_wafflecap_8_0[2|9]/sample vcm col_n[1] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|1] adc_array_wafflecap_8_0[3|9]/sample_n rowon_n[4] row_n[4]
+ adc_array_wafflecap_8_0[3|9]/sample vcm col_n[1] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|1] adc_array_wafflecap_8_0[4|9]/sample_n rowon_n[5] row_n[5]
+ adc_array_wafflecap_8_0[4|9]/sample vcm col_n[1] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|1] adc_array_wafflecap_8_0[5|9]/sample_n rowon_n[6] row_n[6]
+ adc_array_wafflecap_8_0[5|9]/sample vcm col_n[1] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|1] adc_array_wafflecap_8_0[6|9]/sample_n rowon_n[7] row_n[7]
+ adc_array_wafflecap_8_0[6|9]/sample vcm col_n[1] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|1] adc_array_wafflecap_8_0[7|9]/sample_n rowon_n[8] row_n[8]
+ adc_array_wafflecap_8_0[7|9]/sample vcm col_n[1] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|1] adc_array_wafflecap_8_0[8|9]/sample_n rowon_n[9] row_n[9]
+ adc_array_wafflecap_8_0[8|9]/sample vcm col_n[1] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|1] adc_array_wafflecap_8_0[9|9]/sample_n rowon_n[10] row_n[10]
+ adc_array_wafflecap_8_0[9|9]/sample vcm col_n[1] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|1] adc_array_wafflecap_8_0[10|9]/sample_n rowon_n[11]
+ row_n[11] adc_array_wafflecap_8_0[10|9]/sample vcm col_n[1] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|1] adc_array_wafflecap_8_0[11|9]/sample_n rowon_n[12]
+ row_n[12] adc_array_wafflecap_8_0[11|9]/sample vcm col_n[1] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|1] adc_array_wafflecap_8_0[12|9]/sample_n rowon_n[13]
+ row_n[13] adc_array_wafflecap_8_0[12|9]/sample vcm col_n[1] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|1] adc_array_wafflecap_8_0[13|9]/sample_n rowon_n[14]
+ row_n[14] adc_array_wafflecap_8_0[13|9]/sample vcm col_n[1] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|1] adc_array_wafflecap_8_0[14|9]/sample_n rowon_n[15]
+ row_n[15] adc_array_wafflecap_8_0[14|9]/sample vcm col_n[1] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|2] adc_array_wafflecap_8_0[0|9]/sample_n rowon_n[1] row_n[1]
+ adc_array_wafflecap_8_0[0|9]/sample vcm col_n[2] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|2] adc_array_wafflecap_8_0[1|9]/sample_n rowon_n[2] row_n[2]
+ adc_array_wafflecap_8_0[1|9]/sample vcm col_n[2] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|2] adc_array_wafflecap_8_0[2|9]/sample_n rowon_n[3] row_n[3]
+ adc_array_wafflecap_8_0[2|9]/sample vcm col_n[2] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|2] adc_array_wafflecap_8_0[3|9]/sample_n rowon_n[4] row_n[4]
+ adc_array_wafflecap_8_0[3|9]/sample vcm col_n[2] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|2] adc_array_wafflecap_8_0[4|9]/sample_n rowon_n[5] row_n[5]
+ adc_array_wafflecap_8_0[4|9]/sample vcm col_n[2] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|2] adc_array_wafflecap_8_0[5|9]/sample_n rowon_n[6] row_n[6]
+ adc_array_wafflecap_8_0[5|9]/sample vcm col_n[2] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|2] adc_array_wafflecap_8_0[6|9]/sample_n rowon_n[7] row_n[7]
+ adc_array_wafflecap_8_0[6|9]/sample vcm col_n[2] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|2] adc_array_wafflecap_8_0[7|9]/sample_n rowon_n[8] row_n[8]
+ adc_array_wafflecap_8_0[7|9]/sample vcm col_n[2] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|2] adc_array_wafflecap_8_0[8|9]/sample_n rowon_n[9] row_n[9]
+ adc_array_wafflecap_8_0[8|9]/sample vcm col_n[2] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|2] adc_array_wafflecap_8_0[9|9]/sample_n rowon_n[10] row_n[10]
+ adc_array_wafflecap_8_0[9|9]/sample vcm col_n[2] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|2] adc_array_wafflecap_8_0[10|9]/sample_n rowon_n[11]
+ row_n[11] adc_array_wafflecap_8_0[10|9]/sample vcm col_n[2] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|2] adc_array_wafflecap_8_0[11|9]/sample_n rowon_n[12]
+ row_n[12] adc_array_wafflecap_8_0[11|9]/sample vcm col_n[2] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|2] adc_array_wafflecap_8_0[12|9]/sample_n rowon_n[13]
+ row_n[13] adc_array_wafflecap_8_0[12|9]/sample vcm col_n[2] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|2] adc_array_wafflecap_8_0[13|9]/sample_n rowon_n[14]
+ row_n[14] adc_array_wafflecap_8_0[13|9]/sample vcm col_n[2] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|2] adc_array_wafflecap_8_0[14|9]/sample_n rowon_n[15]
+ row_n[15] adc_array_wafflecap_8_0[14|9]/sample vcm col_n[2] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|3] adc_array_wafflecap_8_0[0|9]/sample_n rowon_n[1] row_n[1]
+ adc_array_wafflecap_8_0[0|9]/sample vcm col_n[3] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|3] adc_array_wafflecap_8_0[1|9]/sample_n rowon_n[2] row_n[2]
+ adc_array_wafflecap_8_0[1|9]/sample vcm col_n[3] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|3] adc_array_wafflecap_8_0[2|9]/sample_n rowon_n[3] row_n[3]
+ adc_array_wafflecap_8_0[2|9]/sample vcm col_n[3] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|3] adc_array_wafflecap_8_0[3|9]/sample_n rowon_n[4] row_n[4]
+ adc_array_wafflecap_8_0[3|9]/sample vcm col_n[3] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|3] adc_array_wafflecap_8_0[4|9]/sample_n rowon_n[5] row_n[5]
+ adc_array_wafflecap_8_0[4|9]/sample vcm col_n[3] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|3] adc_array_wafflecap_8_0[5|9]/sample_n rowon_n[6] row_n[6]
+ adc_array_wafflecap_8_0[5|9]/sample vcm col_n[3] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|3] adc_array_wafflecap_8_0[6|9]/sample_n rowon_n[7] row_n[7]
+ adc_array_wafflecap_8_0[6|9]/sample vcm col_n[3] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|3] adc_array_wafflecap_8_0[7|9]/sample_n rowon_n[8] row_n[8]
+ adc_array_wafflecap_8_0[7|9]/sample vcm col_n[3] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|3] adc_array_wafflecap_8_0[8|9]/sample_n rowon_n[9] row_n[9]
+ adc_array_wafflecap_8_0[8|9]/sample vcm col_n[3] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|3] adc_array_wafflecap_8_0[9|9]/sample_n rowon_n[10] row_n[10]
+ adc_array_wafflecap_8_0[9|9]/sample vcm col_n[3] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|3] adc_array_wafflecap_8_0[10|9]/sample_n rowon_n[11]
+ row_n[11] adc_array_wafflecap_8_0[10|9]/sample vcm col_n[3] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|3] adc_array_wafflecap_8_0[11|9]/sample_n rowon_n[12]
+ row_n[12] adc_array_wafflecap_8_0[11|9]/sample vcm col_n[3] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|3] adc_array_wafflecap_8_0[12|9]/sample_n rowon_n[13]
+ row_n[13] adc_array_wafflecap_8_0[12|9]/sample vcm col_n[3] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|3] adc_array_wafflecap_8_0[13|9]/sample_n rowon_n[14]
+ row_n[14] adc_array_wafflecap_8_0[13|9]/sample vcm col_n[3] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|3] adc_array_wafflecap_8_0[14|9]/sample_n rowon_n[15]
+ row_n[15] adc_array_wafflecap_8_0[14|9]/sample vcm col_n[3] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|4] adc_array_wafflecap_8_0[0|9]/sample_n rowon_n[1] row_n[1]
+ adc_array_wafflecap_8_0[0|9]/sample vcm col_n[4] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|4] adc_array_wafflecap_8_0[1|9]/sample_n rowon_n[2] row_n[2]
+ adc_array_wafflecap_8_0[1|9]/sample vcm col_n[4] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|4] adc_array_wafflecap_8_0[2|9]/sample_n rowon_n[3] row_n[3]
+ adc_array_wafflecap_8_0[2|9]/sample vcm col_n[4] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|4] adc_array_wafflecap_8_0[3|9]/sample_n rowon_n[4] row_n[4]
+ adc_array_wafflecap_8_0[3|9]/sample vcm col_n[4] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|4] adc_array_wafflecap_8_0[4|9]/sample_n rowon_n[5] row_n[5]
+ adc_array_wafflecap_8_0[4|9]/sample vcm col_n[4] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|4] adc_array_wafflecap_8_0[5|9]/sample_n rowon_n[6] row_n[6]
+ adc_array_wafflecap_8_0[5|9]/sample vcm col_n[4] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|4] adc_array_wafflecap_8_0[6|9]/sample_n rowon_n[7] row_n[7]
+ adc_array_wafflecap_8_0[6|9]/sample vcm col_n[4] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|4] adc_array_wafflecap_8_0[7|9]/sample_n rowon_n[8] row_n[8]
+ adc_array_wafflecap_8_0[7|9]/sample vcm col_n[4] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|4] adc_array_wafflecap_8_0[8|9]/sample_n rowon_n[9] row_n[9]
+ adc_array_wafflecap_8_0[8|9]/sample vcm col_n[4] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|4] adc_array_wafflecap_8_0[9|9]/sample_n rowon_n[10] row_n[10]
+ adc_array_wafflecap_8_0[9|9]/sample vcm col_n[4] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|4] adc_array_wafflecap_8_0[10|9]/sample_n rowon_n[11]
+ row_n[11] adc_array_wafflecap_8_0[10|9]/sample vcm col_n[4] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|4] adc_array_wafflecap_8_0[11|9]/sample_n rowon_n[12]
+ row_n[12] adc_array_wafflecap_8_0[11|9]/sample vcm col_n[4] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|4] adc_array_wafflecap_8_0[12|9]/sample_n rowon_n[13]
+ row_n[13] adc_array_wafflecap_8_0[12|9]/sample vcm col_n[4] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|4] adc_array_wafflecap_8_0[13|9]/sample_n rowon_n[14]
+ row_n[14] adc_array_wafflecap_8_0[13|9]/sample vcm col_n[4] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|4] adc_array_wafflecap_8_0[14|9]/sample_n rowon_n[15]
+ row_n[15] adc_array_wafflecap_8_0[14|9]/sample vcm col_n[4] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|5] adc_array_wafflecap_8_0[0|9]/sample_n rowon_n[1] row_n[1]
+ adc_array_wafflecap_8_0[0|9]/sample vcm col_n[5] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|5] adc_array_wafflecap_8_0[1|9]/sample_n rowon_n[2] row_n[2]
+ adc_array_wafflecap_8_0[1|9]/sample vcm col_n[5] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|5] adc_array_wafflecap_8_0[2|9]/sample_n rowon_n[3] row_n[3]
+ adc_array_wafflecap_8_0[2|9]/sample vcm col_n[5] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|5] adc_array_wafflecap_8_0[3|9]/sample_n rowon_n[4] row_n[4]
+ adc_array_wafflecap_8_0[3|9]/sample vcm col_n[5] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|5] adc_array_wafflecap_8_0[4|9]/sample_n rowon_n[5] row_n[5]
+ adc_array_wafflecap_8_0[4|9]/sample vcm col_n[5] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|5] adc_array_wafflecap_8_0[5|9]/sample_n rowon_n[6] row_n[6]
+ adc_array_wafflecap_8_0[5|9]/sample vcm col_n[5] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|5] adc_array_wafflecap_8_0[6|9]/sample_n rowon_n[7] row_n[7]
+ adc_array_wafflecap_8_0[6|9]/sample vcm col_n[5] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|5] adc_array_wafflecap_8_0[7|9]/sample_n rowon_n[8] row_n[8]
+ adc_array_wafflecap_8_0[7|9]/sample vcm col_n[5] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|5] adc_array_wafflecap_8_0[8|9]/sample_n rowon_n[9] row_n[9]
+ adc_array_wafflecap_8_0[8|9]/sample vcm col_n[5] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|5] adc_array_wafflecap_8_0[9|9]/sample_n rowon_n[10] row_n[10]
+ adc_array_wafflecap_8_0[9|9]/sample vcm col_n[5] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|5] adc_array_wafflecap_8_0[10|9]/sample_n rowon_n[11]
+ row_n[11] adc_array_wafflecap_8_0[10|9]/sample vcm col_n[5] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|5] adc_array_wafflecap_8_0[11|9]/sample_n rowon_n[12]
+ row_n[12] adc_array_wafflecap_8_0[11|9]/sample vcm col_n[5] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|5] adc_array_wafflecap_8_0[12|9]/sample_n rowon_n[13]
+ row_n[13] adc_array_wafflecap_8_0[12|9]/sample vcm col_n[5] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|5] adc_array_wafflecap_8_0[13|9]/sample_n rowon_n[14]
+ row_n[14] adc_array_wafflecap_8_0[13|9]/sample vcm col_n[5] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|5] adc_array_wafflecap_8_0[14|9]/sample_n rowon_n[15]
+ row_n[15] adc_array_wafflecap_8_0[14|9]/sample vcm col_n[5] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|6] adc_array_wafflecap_8_0[0|9]/sample_n rowon_n[1] row_n[1]
+ adc_array_wafflecap_8_0[0|9]/sample vcm col_n[6] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|6] adc_array_wafflecap_8_0[1|9]/sample_n rowon_n[2] row_n[2]
+ adc_array_wafflecap_8_0[1|9]/sample vcm col_n[6] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|6] adc_array_wafflecap_8_0[2|9]/sample_n rowon_n[3] row_n[3]
+ adc_array_wafflecap_8_0[2|9]/sample vcm col_n[6] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|6] adc_array_wafflecap_8_0[3|9]/sample_n rowon_n[4] row_n[4]
+ adc_array_wafflecap_8_0[3|9]/sample vcm col_n[6] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|6] adc_array_wafflecap_8_0[4|9]/sample_n rowon_n[5] row_n[5]
+ adc_array_wafflecap_8_0[4|9]/sample vcm col_n[6] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|6] adc_array_wafflecap_8_0[5|9]/sample_n rowon_n[6] row_n[6]
+ adc_array_wafflecap_8_0[5|9]/sample vcm col_n[6] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|6] adc_array_wafflecap_8_0[6|9]/sample_n rowon_n[7] row_n[7]
+ adc_array_wafflecap_8_0[6|9]/sample vcm col_n[6] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|6] adc_array_wafflecap_8_0[7|9]/sample_n rowon_n[8] row_n[8]
+ adc_array_wafflecap_8_0[7|9]/sample vcm col_n[6] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|6] adc_array_wafflecap_8_0[8|9]/sample_n rowon_n[9] row_n[9]
+ adc_array_wafflecap_8_0[8|9]/sample vcm col_n[6] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|6] adc_array_wafflecap_8_0[9|9]/sample_n rowon_n[10] row_n[10]
+ adc_array_wafflecap_8_0[9|9]/sample vcm col_n[6] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|6] adc_array_wafflecap_8_0[10|9]/sample_n rowon_n[11]
+ row_n[11] adc_array_wafflecap_8_0[10|9]/sample vcm col_n[6] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|6] adc_array_wafflecap_8_0[11|9]/sample_n rowon_n[12]
+ row_n[12] adc_array_wafflecap_8_0[11|9]/sample vcm col_n[6] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|6] adc_array_wafflecap_8_0[12|9]/sample_n rowon_n[13]
+ row_n[13] adc_array_wafflecap_8_0[12|9]/sample vcm col_n[6] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|6] adc_array_wafflecap_8_0[13|9]/sample_n rowon_n[14]
+ row_n[14] adc_array_wafflecap_8_0[13|9]/sample vcm col_n[6] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|6] adc_array_wafflecap_8_0[14|9]/sample_n rowon_n[15]
+ row_n[15] adc_array_wafflecap_8_0[14|9]/sample vcm col_n[6] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|7] adc_array_wafflecap_8_0[0|9]/sample_n rowon_n[1] row_n[1]
+ adc_array_wafflecap_8_0[0|9]/sample vcm col_n[7] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|7] adc_array_wafflecap_8_0[1|9]/sample_n rowon_n[2] row_n[2]
+ adc_array_wafflecap_8_0[1|9]/sample vcm col_n[7] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|7] adc_array_wafflecap_8_0[2|9]/sample_n rowon_n[3] row_n[3]
+ adc_array_wafflecap_8_0[2|9]/sample vcm col_n[7] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|7] adc_array_wafflecap_8_0[3|9]/sample_n rowon_n[4] row_n[4]
+ adc_array_wafflecap_8_0[3|9]/sample vcm col_n[7] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|7] adc_array_wafflecap_8_0[4|9]/sample_n rowon_n[5] row_n[5]
+ adc_array_wafflecap_8_0[4|9]/sample vcm col_n[7] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|7] adc_array_wafflecap_8_0[5|9]/sample_n rowon_n[6] row_n[6]
+ adc_array_wafflecap_8_0[5|9]/sample vcm col_n[7] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|7] adc_array_wafflecap_8_0[6|9]/sample_n rowon_n[7] row_n[7]
+ adc_array_wafflecap_8_0[6|9]/sample vcm col_n[7] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|7] adc_array_wafflecap_8_0[7|9]/sample_n rowon_n[8] row_n[8]
+ adc_array_wafflecap_8_0[7|9]/sample vcm col_n[7] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|7] adc_array_wafflecap_8_0[8|9]/sample_n rowon_n[9] row_n[9]
+ adc_array_wafflecap_8_0[8|9]/sample vcm col_n[7] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|7] adc_array_wafflecap_8_0[9|9]/sample_n rowon_n[10] row_n[10]
+ adc_array_wafflecap_8_0[9|9]/sample vcm col_n[7] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|7] adc_array_wafflecap_8_0[10|9]/sample_n rowon_n[11]
+ row_n[11] adc_array_wafflecap_8_0[10|9]/sample vcm col_n[7] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|7] adc_array_wafflecap_8_0[11|9]/sample_n rowon_n[12]
+ row_n[12] adc_array_wafflecap_8_0[11|9]/sample vcm col_n[7] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|7] adc_array_wafflecap_8_0[12|9]/sample_n rowon_n[13]
+ row_n[13] adc_array_wafflecap_8_0[12|9]/sample vcm col_n[7] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|7] adc_array_wafflecap_8_0[13|9]/sample_n rowon_n[14]
+ row_n[14] adc_array_wafflecap_8_0[13|9]/sample vcm col_n[7] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|7] adc_array_wafflecap_8_0[14|9]/sample_n rowon_n[15]
+ row_n[15] adc_array_wafflecap_8_0[14|9]/sample vcm col_n[7] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|8] adc_array_wafflecap_8_0[0|9]/sample_n rowon_n[1] row_n[1]
+ adc_array_wafflecap_8_0[0|9]/sample vcm col_n[8] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|8] adc_array_wafflecap_8_0[1|9]/sample_n rowon_n[2] row_n[2]
+ adc_array_wafflecap_8_0[1|9]/sample vcm col_n[8] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|8] adc_array_wafflecap_8_0[2|9]/sample_n rowon_n[3] row_n[3]
+ adc_array_wafflecap_8_0[2|9]/sample vcm col_n[8] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|8] adc_array_wafflecap_8_0[3|9]/sample_n rowon_n[4] row_n[4]
+ adc_array_wafflecap_8_0[3|9]/sample vcm col_n[8] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|8] adc_array_wafflecap_8_0[4|9]/sample_n rowon_n[5] row_n[5]
+ adc_array_wafflecap_8_0[4|9]/sample vcm col_n[8] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|8] adc_array_wafflecap_8_0[5|9]/sample_n rowon_n[6] row_n[6]
+ adc_array_wafflecap_8_0[5|9]/sample vcm col_n[8] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|8] adc_array_wafflecap_8_0[6|9]/sample_n rowon_n[7] row_n[7]
+ adc_array_wafflecap_8_0[6|9]/sample vcm col_n[8] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|8] adc_array_wafflecap_8_0[7|9]/sample_n rowon_n[8] row_n[8]
+ adc_array_wafflecap_8_0[7|9]/sample vcm col_n[8] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|8] adc_array_wafflecap_8_0[8|9]/sample_n rowon_n[9] row_n[9]
+ adc_array_wafflecap_8_0[8|9]/sample vcm col_n[8] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|8] adc_array_wafflecap_8_0[9|9]/sample_n rowon_n[10] row_n[10]
+ adc_array_wafflecap_8_0[9|9]/sample vcm col_n[8] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|8] adc_array_wafflecap_8_0[10|9]/sample_n rowon_n[11]
+ row_n[11] adc_array_wafflecap_8_0[10|9]/sample vcm col_n[8] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|8] adc_array_wafflecap_8_0[11|9]/sample_n rowon_n[12]
+ row_n[12] adc_array_wafflecap_8_0[11|9]/sample vcm col_n[8] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|8] adc_array_wafflecap_8_0[12|9]/sample_n rowon_n[13]
+ row_n[13] adc_array_wafflecap_8_0[12|9]/sample vcm col_n[8] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|8] adc_array_wafflecap_8_0[13|9]/sample_n rowon_n[14]
+ row_n[14] adc_array_wafflecap_8_0[13|9]/sample vcm col_n[8] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|8] adc_array_wafflecap_8_0[14|9]/sample_n rowon_n[15]
+ row_n[15] adc_array_wafflecap_8_0[14|9]/sample vcm col_n[8] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|9] adc_array_wafflecap_8_0[0|9]/sample_n rowon_n[1] row_n[1]
+ adc_array_wafflecap_8_0[0|9]/sample vcm col_n[9] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|9] adc_array_wafflecap_8_0[1|9]/sample_n rowon_n[2] row_n[2]
+ adc_array_wafflecap_8_0[1|9]/sample vcm col_n[9] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|9] adc_array_wafflecap_8_0[2|9]/sample_n rowon_n[3] row_n[3]
+ adc_array_wafflecap_8_0[2|9]/sample vcm col_n[9] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|9] adc_array_wafflecap_8_0[3|9]/sample_n rowon_n[4] row_n[4]
+ adc_array_wafflecap_8_0[3|9]/sample vcm col_n[9] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|9] adc_array_wafflecap_8_0[4|9]/sample_n rowon_n[5] row_n[5]
+ adc_array_wafflecap_8_0[4|9]/sample vcm col_n[9] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|9] adc_array_wafflecap_8_0[5|9]/sample_n rowon_n[6] row_n[6]
+ adc_array_wafflecap_8_0[5|9]/sample vcm col_n[9] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|9] adc_array_wafflecap_8_0[6|9]/sample_n rowon_n[7] row_n[7]
+ adc_array_wafflecap_8_0[6|9]/sample vcm col_n[9] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|9] adc_array_wafflecap_8_0[7|9]/sample_n rowon_n[8] row_n[8]
+ adc_array_wafflecap_8_0[7|9]/sample vcm col_n[9] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|9] adc_array_wafflecap_8_0[8|9]/sample_n rowon_n[9] row_n[9]
+ adc_array_wafflecap_8_0[8|9]/sample vcm col_n[9] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|9] adc_array_wafflecap_8_0[9|9]/sample_n rowon_n[10] row_n[10]
+ adc_array_wafflecap_8_0[9|9]/sample vcm col_n[9] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|9] adc_array_wafflecap_8_0[10|9]/sample_n rowon_n[11]
+ row_n[11] adc_array_wafflecap_8_0[10|9]/sample vcm col_n[9] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|9] adc_array_wafflecap_8_0[11|9]/sample_n rowon_n[12]
+ row_n[12] adc_array_wafflecap_8_0[11|9]/sample vcm col_n[9] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|9] adc_array_wafflecap_8_0[12|9]/sample_n rowon_n[13]
+ row_n[13] adc_array_wafflecap_8_0[12|9]/sample vcm col_n[9] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|9] adc_array_wafflecap_8_0[13|9]/sample_n rowon_n[14]
+ row_n[14] adc_array_wafflecap_8_0[13|9]/sample vcm col_n[9] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|9] adc_array_wafflecap_8_0[14|9]/sample_n rowon_n[15]
+ row_n[15] adc_array_wafflecap_8_0[14|9]/sample vcm col_n[9] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|10] adc_array_wafflecap_8_0[0|9]/sample_n rowon_n[1] row_n[1]
+ adc_array_wafflecap_8_0[0|9]/sample vcm col_n[10] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|10] adc_array_wafflecap_8_0[1|9]/sample_n rowon_n[2] row_n[2]
+ adc_array_wafflecap_8_0[1|9]/sample vcm col_n[10] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|10] adc_array_wafflecap_8_0[2|9]/sample_n rowon_n[3] row_n[3]
+ adc_array_wafflecap_8_0[2|9]/sample vcm col_n[10] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|10] adc_array_wafflecap_8_0[3|9]/sample_n rowon_n[4] row_n[4]
+ adc_array_wafflecap_8_0[3|9]/sample vcm col_n[10] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|10] adc_array_wafflecap_8_0[4|9]/sample_n rowon_n[5] row_n[5]
+ adc_array_wafflecap_8_0[4|9]/sample vcm col_n[10] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|10] adc_array_wafflecap_8_0[5|9]/sample_n rowon_n[6] row_n[6]
+ adc_array_wafflecap_8_0[5|9]/sample vcm col_n[10] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|10] adc_array_wafflecap_8_0[6|9]/sample_n rowon_n[7] row_n[7]
+ adc_array_wafflecap_8_0[6|9]/sample vcm col_n[10] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|10] adc_array_wafflecap_8_0[7|9]/sample_n rowon_n[8] row_n[8]
+ adc_array_wafflecap_8_0[7|9]/sample vcm col_n[10] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|10] adc_array_wafflecap_8_0[8|9]/sample_n rowon_n[9] row_n[9]
+ adc_array_wafflecap_8_0[8|9]/sample vcm col_n[10] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|10] adc_array_wafflecap_8_0[9|9]/sample_n rowon_n[10] row_n[10]
+ adc_array_wafflecap_8_0[9|9]/sample vcm col_n[10] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|10] adc_array_wafflecap_8_0[10|9]/sample_n rowon_n[11]
+ row_n[11] adc_array_wafflecap_8_0[10|9]/sample vcm col_n[10] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|10] adc_array_wafflecap_8_0[11|9]/sample_n rowon_n[12]
+ row_n[12] adc_array_wafflecap_8_0[11|9]/sample vcm col_n[10] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|10] adc_array_wafflecap_8_0[12|9]/sample_n rowon_n[13]
+ row_n[13] adc_array_wafflecap_8_0[12|9]/sample vcm col_n[10] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|10] adc_array_wafflecap_8_0[13|9]/sample_n rowon_n[14]
+ row_n[14] adc_array_wafflecap_8_0[13|9]/sample vcm col_n[10] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|10] adc_array_wafflecap_8_0[14|9]/sample_n rowon_n[15]
+ row_n[15] adc_array_wafflecap_8_0[14|9]/sample vcm col_n[10] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|11] adc_array_wafflecap_8_0[0|9]/sample_n rowon_n[1] row_n[1]
+ adc_array_wafflecap_8_0[0|9]/sample vcm col_n[11] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|11] adc_array_wafflecap_8_0[1|9]/sample_n rowon_n[2] row_n[2]
+ adc_array_wafflecap_8_0[1|9]/sample vcm col_n[11] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|11] adc_array_wafflecap_8_0[2|9]/sample_n rowon_n[3] row_n[3]
+ adc_array_wafflecap_8_0[2|9]/sample vcm col_n[11] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|11] adc_array_wafflecap_8_0[3|9]/sample_n rowon_n[4] row_n[4]
+ adc_array_wafflecap_8_0[3|9]/sample vcm col_n[11] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|11] adc_array_wafflecap_8_0[4|9]/sample_n rowon_n[5] row_n[5]
+ adc_array_wafflecap_8_0[4|9]/sample vcm col_n[11] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|11] adc_array_wafflecap_8_0[5|9]/sample_n rowon_n[6] row_n[6]
+ adc_array_wafflecap_8_0[5|9]/sample vcm col_n[11] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|11] adc_array_wafflecap_8_0[6|9]/sample_n rowon_n[7] row_n[7]
+ adc_array_wafflecap_8_0[6|9]/sample vcm col_n[11] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|11] adc_array_wafflecap_8_0[7|9]/sample_n rowon_n[8] row_n[8]
+ adc_array_wafflecap_8_0[7|9]/sample vcm col_n[11] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|11] adc_array_wafflecap_8_0[8|9]/sample_n rowon_n[9] row_n[9]
+ adc_array_wafflecap_8_0[8|9]/sample vcm col_n[11] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|11] adc_array_wafflecap_8_0[9|9]/sample_n rowon_n[10] row_n[10]
+ adc_array_wafflecap_8_0[9|9]/sample vcm col_n[11] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|11] adc_array_wafflecap_8_0[10|9]/sample_n rowon_n[11]
+ row_n[11] adc_array_wafflecap_8_0[10|9]/sample vcm col_n[11] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|11] adc_array_wafflecap_8_0[11|9]/sample_n rowon_n[12]
+ row_n[12] adc_array_wafflecap_8_0[11|9]/sample vcm col_n[11] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|11] adc_array_wafflecap_8_0[12|9]/sample_n rowon_n[13]
+ row_n[13] adc_array_wafflecap_8_0[12|9]/sample vcm col_n[11] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|11] adc_array_wafflecap_8_0[13|9]/sample_n rowon_n[14]
+ row_n[14] adc_array_wafflecap_8_0[13|9]/sample vcm col_n[11] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|11] adc_array_wafflecap_8_0[14|9]/sample_n rowon_n[15]
+ row_n[15] adc_array_wafflecap_8_0[14|9]/sample vcm col_n[11] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|12] adc_array_wafflecap_8_0[0|9]/sample_n rowon_n[1] row_n[1]
+ adc_array_wafflecap_8_0[0|9]/sample vcm col_n[12] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|12] adc_array_wafflecap_8_0[1|9]/sample_n rowon_n[2] row_n[2]
+ adc_array_wafflecap_8_0[1|9]/sample vcm col_n[12] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|12] adc_array_wafflecap_8_0[2|9]/sample_n rowon_n[3] row_n[3]
+ adc_array_wafflecap_8_0[2|9]/sample vcm col_n[12] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|12] adc_array_wafflecap_8_0[3|9]/sample_n rowon_n[4] row_n[4]
+ adc_array_wafflecap_8_0[3|9]/sample vcm col_n[12] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|12] adc_array_wafflecap_8_0[4|9]/sample_n rowon_n[5] row_n[5]
+ adc_array_wafflecap_8_0[4|9]/sample vcm col_n[12] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|12] adc_array_wafflecap_8_0[5|9]/sample_n rowon_n[6] row_n[6]
+ adc_array_wafflecap_8_0[5|9]/sample vcm col_n[12] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|12] adc_array_wafflecap_8_0[6|9]/sample_n rowon_n[7] row_n[7]
+ adc_array_wafflecap_8_0[6|9]/sample vcm col_n[12] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|12] adc_array_wafflecap_8_0[7|9]/sample_n rowon_n[8] row_n[8]
+ adc_array_wafflecap_8_0[7|9]/sample vcm col_n[12] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|12] adc_array_wafflecap_8_0[8|9]/sample_n rowon_n[9] row_n[9]
+ adc_array_wafflecap_8_0[8|9]/sample vcm col_n[12] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|12] adc_array_wafflecap_8_0[9|9]/sample_n rowon_n[10] row_n[10]
+ adc_array_wafflecap_8_0[9|9]/sample vcm col_n[12] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|12] adc_array_wafflecap_8_0[10|9]/sample_n rowon_n[11]
+ row_n[11] adc_array_wafflecap_8_0[10|9]/sample vcm col_n[12] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|12] adc_array_wafflecap_8_0[11|9]/sample_n rowon_n[12]
+ row_n[12] adc_array_wafflecap_8_0[11|9]/sample vcm col_n[12] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|12] adc_array_wafflecap_8_0[12|9]/sample_n rowon_n[13]
+ row_n[13] adc_array_wafflecap_8_0[12|9]/sample vcm col_n[12] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|12] adc_array_wafflecap_8_0[13|9]/sample_n rowon_n[14]
+ row_n[14] adc_array_wafflecap_8_0[13|9]/sample vcm col_n[12] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|12] adc_array_wafflecap_8_0[14|9]/sample_n rowon_n[15]
+ row_n[15] adc_array_wafflecap_8_0[14|9]/sample vcm col_n[12] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|13] adc_array_wafflecap_8_0[0|9]/sample_n rowon_n[1] row_n[1]
+ adc_array_wafflecap_8_0[0|9]/sample vcm col_n[13] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|13] adc_array_wafflecap_8_0[1|9]/sample_n rowon_n[2] row_n[2]
+ adc_array_wafflecap_8_0[1|9]/sample vcm col_n[13] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|13] adc_array_wafflecap_8_0[2|9]/sample_n rowon_n[3] row_n[3]
+ adc_array_wafflecap_8_0[2|9]/sample vcm col_n[13] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|13] adc_array_wafflecap_8_0[3|9]/sample_n rowon_n[4] row_n[4]
+ adc_array_wafflecap_8_0[3|9]/sample vcm col_n[13] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|13] adc_array_wafflecap_8_0[4|9]/sample_n rowon_n[5] row_n[5]
+ adc_array_wafflecap_8_0[4|9]/sample vcm col_n[13] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|13] adc_array_wafflecap_8_0[5|9]/sample_n rowon_n[6] row_n[6]
+ adc_array_wafflecap_8_0[5|9]/sample vcm col_n[13] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|13] adc_array_wafflecap_8_0[6|9]/sample_n rowon_n[7] row_n[7]
+ adc_array_wafflecap_8_0[6|9]/sample vcm col_n[13] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|13] adc_array_wafflecap_8_0[7|9]/sample_n rowon_n[8] row_n[8]
+ adc_array_wafflecap_8_0[7|9]/sample vcm col_n[13] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|13] adc_array_wafflecap_8_0[8|9]/sample_n rowon_n[9] row_n[9]
+ adc_array_wafflecap_8_0[8|9]/sample vcm col_n[13] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|13] adc_array_wafflecap_8_0[9|9]/sample_n rowon_n[10] row_n[10]
+ adc_array_wafflecap_8_0[9|9]/sample vcm col_n[13] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|13] adc_array_wafflecap_8_0[10|9]/sample_n rowon_n[11]
+ row_n[11] adc_array_wafflecap_8_0[10|9]/sample vcm col_n[13] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|13] adc_array_wafflecap_8_0[11|9]/sample_n rowon_n[12]
+ row_n[12] adc_array_wafflecap_8_0[11|9]/sample vcm col_n[13] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|13] adc_array_wafflecap_8_0[12|9]/sample_n rowon_n[13]
+ row_n[13] adc_array_wafflecap_8_0[12|9]/sample vcm col_n[13] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|13] adc_array_wafflecap_8_0[13|9]/sample_n rowon_n[14]
+ row_n[14] adc_array_wafflecap_8_0[13|9]/sample vcm col_n[13] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|13] adc_array_wafflecap_8_0[14|9]/sample_n rowon_n[15]
+ row_n[15] adc_array_wafflecap_8_0[14|9]/sample vcm col_n[13] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|14] adc_array_wafflecap_8_0[0|9]/sample_n rowon_n[1] row_n[1]
+ adc_array_wafflecap_8_0[0|9]/sample vcm col_n[14] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|14] adc_array_wafflecap_8_0[1|9]/sample_n rowon_n[2] row_n[2]
+ adc_array_wafflecap_8_0[1|9]/sample vcm col_n[14] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|14] adc_array_wafflecap_8_0[2|9]/sample_n rowon_n[3] row_n[3]
+ adc_array_wafflecap_8_0[2|9]/sample vcm col_n[14] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|14] adc_array_wafflecap_8_0[3|9]/sample_n rowon_n[4] row_n[4]
+ adc_array_wafflecap_8_0[3|9]/sample vcm col_n[14] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|14] adc_array_wafflecap_8_0[4|9]/sample_n rowon_n[5] row_n[5]
+ adc_array_wafflecap_8_0[4|9]/sample vcm col_n[14] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|14] adc_array_wafflecap_8_0[5|9]/sample_n rowon_n[6] row_n[6]
+ adc_array_wafflecap_8_0[5|9]/sample vcm col_n[14] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|14] adc_array_wafflecap_8_0[6|9]/sample_n rowon_n[7] row_n[7]
+ adc_array_wafflecap_8_0[6|9]/sample vcm col_n[14] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|14] adc_array_wafflecap_8_0[7|9]/sample_n rowon_n[8] row_n[8]
+ adc_array_wafflecap_8_0[7|9]/sample vcm col_n[14] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|14] adc_array_wafflecap_8_0[8|9]/sample_n rowon_n[9] row_n[9]
+ adc_array_wafflecap_8_0[8|9]/sample vcm col_n[14] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|14] adc_array_wafflecap_8_0[9|9]/sample_n rowon_n[10] row_n[10]
+ adc_array_wafflecap_8_0[9|9]/sample vcm col_n[14] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|14] adc_array_wafflecap_8_0[10|9]/sample_n rowon_n[11]
+ row_n[11] adc_array_wafflecap_8_0[10|9]/sample vcm col_n[14] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|14] adc_array_wafflecap_8_0[11|9]/sample_n rowon_n[12]
+ row_n[12] adc_array_wafflecap_8_0[11|9]/sample vcm col_n[14] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|14] adc_array_wafflecap_8_0[12|9]/sample_n rowon_n[13]
+ row_n[13] adc_array_wafflecap_8_0[12|9]/sample vcm col_n[14] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|14] adc_array_wafflecap_8_0[13|9]/sample_n rowon_n[14]
+ row_n[14] adc_array_wafflecap_8_0[13|9]/sample vcm col_n[14] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|14] adc_array_wafflecap_8_0[14|9]/sample_n rowon_n[15]
+ row_n[15] adc_array_wafflecap_8_0[14|9]/sample vcm col_n[14] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|15] adc_array_wafflecap_8_0[0|9]/sample_n rowon_n[1] row_n[1]
+ adc_array_wafflecap_8_0[0|9]/sample vcm col_n[15] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|15] adc_array_wafflecap_8_0[1|9]/sample_n rowon_n[2] row_n[2]
+ adc_array_wafflecap_8_0[1|9]/sample vcm col_n[15] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|15] adc_array_wafflecap_8_0[2|9]/sample_n rowon_n[3] row_n[3]
+ adc_array_wafflecap_8_0[2|9]/sample vcm col_n[15] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|15] adc_array_wafflecap_8_0[3|9]/sample_n rowon_n[4] row_n[4]
+ adc_array_wafflecap_8_0[3|9]/sample vcm col_n[15] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|15] adc_array_wafflecap_8_0[4|9]/sample_n rowon_n[5] row_n[5]
+ adc_array_wafflecap_8_0[4|9]/sample vcm col_n[15] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|15] adc_array_wafflecap_8_0[5|9]/sample_n rowon_n[6] row_n[6]
+ adc_array_wafflecap_8_0[5|9]/sample vcm col_n[15] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|15] adc_array_wafflecap_8_0[6|9]/sample_n rowon_n[7] row_n[7]
+ adc_array_wafflecap_8_0[6|9]/sample vcm col_n[15] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|15] adc_array_wafflecap_8_0[7|9]/sample_n rowon_n[8] row_n[8]
+ adc_array_wafflecap_8_0[7|9]/sample vcm col_n[15] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|15] adc_array_wafflecap_8_0[8|9]/sample_n rowon_n[9] row_n[9]
+ adc_array_wafflecap_8_0[8|9]/sample vcm col_n[15] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|15] adc_array_wafflecap_8_0[9|9]/sample_n rowon_n[10] row_n[10]
+ adc_array_wafflecap_8_0[9|9]/sample vcm col_n[15] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|15] adc_array_wafflecap_8_0[10|9]/sample_n rowon_n[11]
+ row_n[11] adc_array_wafflecap_8_0[10|9]/sample vcm col_n[15] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|15] adc_array_wafflecap_8_0[11|9]/sample_n rowon_n[12]
+ row_n[12] adc_array_wafflecap_8_0[11|9]/sample vcm col_n[15] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|15] adc_array_wafflecap_8_0[12|9]/sample_n rowon_n[13]
+ row_n[13] adc_array_wafflecap_8_0[12|9]/sample vcm col_n[15] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|15] adc_array_wafflecap_8_0[13|9]/sample_n rowon_n[14]
+ row_n[14] adc_array_wafflecap_8_0[13|9]/sample vcm col_n[15] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|15] adc_array_wafflecap_8_0[14|9]/sample_n rowon_n[15]
+ row_n[15] adc_array_wafflecap_8_0[14|9]/sample vcm col_n[15] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|16] adc_array_wafflecap_8_0[0|9]/sample_n rowon_n[1] row_n[1]
+ adc_array_wafflecap_8_0[0|9]/sample vcm col_n[16] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|16] adc_array_wafflecap_8_0[1|9]/sample_n rowon_n[2] row_n[2]
+ adc_array_wafflecap_8_0[1|9]/sample vcm col_n[16] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|16] adc_array_wafflecap_8_0[2|9]/sample_n rowon_n[3] row_n[3]
+ adc_array_wafflecap_8_0[2|9]/sample vcm col_n[16] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|16] adc_array_wafflecap_8_0[3|9]/sample_n rowon_n[4] row_n[4]
+ adc_array_wafflecap_8_0[3|9]/sample vcm col_n[16] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|16] adc_array_wafflecap_8_0[4|9]/sample_n rowon_n[5] row_n[5]
+ adc_array_wafflecap_8_0[4|9]/sample vcm col_n[16] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|16] adc_array_wafflecap_8_0[5|9]/sample_n rowon_n[6] row_n[6]
+ adc_array_wafflecap_8_0[5|9]/sample vcm col_n[16] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|16] adc_array_wafflecap_8_0[6|9]/sample_n rowon_n[7] row_n[7]
+ adc_array_wafflecap_8_0[6|9]/sample vcm col_n[16] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|16] adc_array_wafflecap_8_0[7|9]/sample_n rowon_n[8] row_n[8]
+ adc_array_wafflecap_8_0[7|9]/sample vcm col_n[16] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|16] adc_array_wafflecap_8_0[8|9]/sample_n rowon_n[9] row_n[9]
+ adc_array_wafflecap_8_0[8|9]/sample vcm col_n[16] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|16] adc_array_wafflecap_8_0[9|9]/sample_n rowon_n[10] row_n[10]
+ adc_array_wafflecap_8_0[9|9]/sample vcm col_n[16] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|16] adc_array_wafflecap_8_0[10|9]/sample_n rowon_n[11]
+ row_n[11] adc_array_wafflecap_8_0[10|9]/sample vcm col_n[16] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|16] adc_array_wafflecap_8_0[11|9]/sample_n rowon_n[12]
+ row_n[12] adc_array_wafflecap_8_0[11|9]/sample vcm col_n[16] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|16] adc_array_wafflecap_8_0[12|9]/sample_n rowon_n[13]
+ row_n[13] adc_array_wafflecap_8_0[12|9]/sample vcm col_n[16] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|16] adc_array_wafflecap_8_0[13|9]/sample_n rowon_n[14]
+ row_n[14] adc_array_wafflecap_8_0[13|9]/sample vcm col_n[16] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|16] adc_array_wafflecap_8_0[14|9]/sample_n rowon_n[15]
+ row_n[15] adc_array_wafflecap_8_0[14|9]/sample vcm col_n[16] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|17] adc_array_wafflecap_8_0[0|9]/sample_n rowon_n[1] row_n[1]
+ adc_array_wafflecap_8_0[0|9]/sample vcm col_n[17] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|17] adc_array_wafflecap_8_0[1|9]/sample_n rowon_n[2] row_n[2]
+ adc_array_wafflecap_8_0[1|9]/sample vcm col_n[17] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|17] adc_array_wafflecap_8_0[2|9]/sample_n rowon_n[3] row_n[3]
+ adc_array_wafflecap_8_0[2|9]/sample vcm col_n[17] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|17] adc_array_wafflecap_8_0[3|9]/sample_n rowon_n[4] row_n[4]
+ adc_array_wafflecap_8_0[3|9]/sample vcm col_n[17] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|17] adc_array_wafflecap_8_0[4|9]/sample_n rowon_n[5] row_n[5]
+ adc_array_wafflecap_8_0[4|9]/sample vcm col_n[17] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|17] adc_array_wafflecap_8_0[5|9]/sample_n rowon_n[6] row_n[6]
+ adc_array_wafflecap_8_0[5|9]/sample vcm col_n[17] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|17] adc_array_wafflecap_8_0[6|9]/sample_n rowon_n[7] row_n[7]
+ adc_array_wafflecap_8_0[6|9]/sample vcm col_n[17] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|17] adc_array_wafflecap_8_0[7|9]/sample_n rowon_n[8] row_n[8]
+ adc_array_wafflecap_8_0[7|9]/sample vcm col_n[17] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|17] adc_array_wafflecap_8_0[8|9]/sample_n rowon_n[9] row_n[9]
+ adc_array_wafflecap_8_0[8|9]/sample vcm col_n[17] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|17] adc_array_wafflecap_8_0[9|9]/sample_n rowon_n[10] row_n[10]
+ adc_array_wafflecap_8_0[9|9]/sample vcm col_n[17] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|17] adc_array_wafflecap_8_0[10|9]/sample_n rowon_n[11]
+ row_n[11] adc_array_wafflecap_8_0[10|9]/sample vcm col_n[17] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|17] adc_array_wafflecap_8_0[11|9]/sample_n rowon_n[12]
+ row_n[12] adc_array_wafflecap_8_0[11|9]/sample vcm col_n[17] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|17] adc_array_wafflecap_8_0[12|9]/sample_n rowon_n[13]
+ row_n[13] adc_array_wafflecap_8_0[12|9]/sample vcm col_n[17] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|17] adc_array_wafflecap_8_0[13|9]/sample_n rowon_n[14]
+ row_n[14] adc_array_wafflecap_8_0[13|9]/sample vcm col_n[17] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|17] adc_array_wafflecap_8_0[14|9]/sample_n rowon_n[15]
+ row_n[15] adc_array_wafflecap_8_0[14|9]/sample vcm col_n[17] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|18] adc_array_wafflecap_8_0[0|9]/sample_n rowon_n[1] row_n[1]
+ adc_array_wafflecap_8_0[0|9]/sample vcm col_n[18] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|18] adc_array_wafflecap_8_0[1|9]/sample_n rowon_n[2] row_n[2]
+ adc_array_wafflecap_8_0[1|9]/sample vcm col_n[18] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|18] adc_array_wafflecap_8_0[2|9]/sample_n rowon_n[3] row_n[3]
+ adc_array_wafflecap_8_0[2|9]/sample vcm col_n[18] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|18] adc_array_wafflecap_8_0[3|9]/sample_n rowon_n[4] row_n[4]
+ adc_array_wafflecap_8_0[3|9]/sample vcm col_n[18] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|18] adc_array_wafflecap_8_0[4|9]/sample_n rowon_n[5] row_n[5]
+ adc_array_wafflecap_8_0[4|9]/sample vcm col_n[18] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|18] adc_array_wafflecap_8_0[5|9]/sample_n rowon_n[6] row_n[6]
+ adc_array_wafflecap_8_0[5|9]/sample vcm col_n[18] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|18] adc_array_wafflecap_8_0[6|9]/sample_n rowon_n[7] row_n[7]
+ adc_array_wafflecap_8_0[6|9]/sample vcm col_n[18] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|18] adc_array_wafflecap_8_0[7|9]/sample_n rowon_n[8] row_n[8]
+ adc_array_wafflecap_8_0[7|9]/sample vcm col_n[18] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|18] adc_array_wafflecap_8_0[8|9]/sample_n rowon_n[9] row_n[9]
+ adc_array_wafflecap_8_0[8|9]/sample vcm col_n[18] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|18] adc_array_wafflecap_8_0[9|9]/sample_n rowon_n[10] row_n[10]
+ adc_array_wafflecap_8_0[9|9]/sample vcm col_n[18] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|18] adc_array_wafflecap_8_0[10|9]/sample_n rowon_n[11]
+ row_n[11] adc_array_wafflecap_8_0[10|9]/sample vcm col_n[18] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|18] adc_array_wafflecap_8_0[11|9]/sample_n rowon_n[12]
+ row_n[12] adc_array_wafflecap_8_0[11|9]/sample vcm col_n[18] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|18] adc_array_wafflecap_8_0[12|9]/sample_n rowon_n[13]
+ row_n[13] adc_array_wafflecap_8_0[12|9]/sample vcm col_n[18] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|18] adc_array_wafflecap_8_0[13|9]/sample_n rowon_n[14]
+ row_n[14] adc_array_wafflecap_8_0[13|9]/sample vcm col_n[18] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|18] adc_array_wafflecap_8_0[14|9]/sample_n rowon_n[15]
+ row_n[15] adc_array_wafflecap_8_0[14|9]/sample vcm col_n[18] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|19] adc_array_wafflecap_8_0[0|9]/sample_n rowon_n[1] row_n[1]
+ adc_array_wafflecap_8_0[0|9]/sample vcm col_n[19] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|19] adc_array_wafflecap_8_0[1|9]/sample_n rowon_n[2] row_n[2]
+ adc_array_wafflecap_8_0[1|9]/sample vcm col_n[19] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|19] adc_array_wafflecap_8_0[2|9]/sample_n rowon_n[3] row_n[3]
+ adc_array_wafflecap_8_0[2|9]/sample vcm col_n[19] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|19] adc_array_wafflecap_8_0[3|9]/sample_n rowon_n[4] row_n[4]
+ adc_array_wafflecap_8_0[3|9]/sample vcm col_n[19] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|19] adc_array_wafflecap_8_0[4|9]/sample_n rowon_n[5] row_n[5]
+ adc_array_wafflecap_8_0[4|9]/sample vcm col_n[19] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|19] adc_array_wafflecap_8_0[5|9]/sample_n rowon_n[6] row_n[6]
+ adc_array_wafflecap_8_0[5|9]/sample vcm col_n[19] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|19] adc_array_wafflecap_8_0[6|9]/sample_n rowon_n[7] row_n[7]
+ adc_array_wafflecap_8_0[6|9]/sample vcm col_n[19] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|19] adc_array_wafflecap_8_0[7|9]/sample_n rowon_n[8] row_n[8]
+ adc_array_wafflecap_8_0[7|9]/sample vcm col_n[19] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|19] adc_array_wafflecap_8_0[8|9]/sample_n rowon_n[9] row_n[9]
+ adc_array_wafflecap_8_0[8|9]/sample vcm col_n[19] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|19] adc_array_wafflecap_8_0[9|9]/sample_n rowon_n[10] row_n[10]
+ adc_array_wafflecap_8_0[9|9]/sample vcm col_n[19] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|19] adc_array_wafflecap_8_0[10|9]/sample_n rowon_n[11]
+ row_n[11] adc_array_wafflecap_8_0[10|9]/sample vcm col_n[19] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|19] adc_array_wafflecap_8_0[11|9]/sample_n rowon_n[12]
+ row_n[12] adc_array_wafflecap_8_0[11|9]/sample vcm col_n[19] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|19] adc_array_wafflecap_8_0[12|9]/sample_n rowon_n[13]
+ row_n[13] adc_array_wafflecap_8_0[12|9]/sample vcm col_n[19] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|19] adc_array_wafflecap_8_0[13|9]/sample_n rowon_n[14]
+ row_n[14] adc_array_wafflecap_8_0[13|9]/sample vcm col_n[19] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|19] adc_array_wafflecap_8_0[14|9]/sample_n rowon_n[15]
+ row_n[15] adc_array_wafflecap_8_0[14|9]/sample vcm col_n[19] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|20] adc_array_wafflecap_8_0[0|9]/sample_n rowon_n[1] row_n[1]
+ adc_array_wafflecap_8_0[0|9]/sample vcm col_n[20] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|20] adc_array_wafflecap_8_0[1|9]/sample_n rowon_n[2] row_n[2]
+ adc_array_wafflecap_8_0[1|9]/sample vcm col_n[20] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|20] adc_array_wafflecap_8_0[2|9]/sample_n rowon_n[3] row_n[3]
+ adc_array_wafflecap_8_0[2|9]/sample vcm col_n[20] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|20] adc_array_wafflecap_8_0[3|9]/sample_n rowon_n[4] row_n[4]
+ adc_array_wafflecap_8_0[3|9]/sample vcm col_n[20] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|20] adc_array_wafflecap_8_0[4|9]/sample_n rowon_n[5] row_n[5]
+ adc_array_wafflecap_8_0[4|9]/sample vcm col_n[20] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|20] adc_array_wafflecap_8_0[5|9]/sample_n rowon_n[6] row_n[6]
+ adc_array_wafflecap_8_0[5|9]/sample vcm col_n[20] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|20] adc_array_wafflecap_8_0[6|9]/sample_n rowon_n[7] row_n[7]
+ adc_array_wafflecap_8_0[6|9]/sample vcm col_n[20] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|20] adc_array_wafflecap_8_0[7|9]/sample_n rowon_n[8] row_n[8]
+ adc_array_wafflecap_8_0[7|9]/sample vcm col_n[20] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|20] adc_array_wafflecap_8_0[8|9]/sample_n rowon_n[9] row_n[9]
+ adc_array_wafflecap_8_0[8|9]/sample vcm col_n[20] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|20] adc_array_wafflecap_8_0[9|9]/sample_n rowon_n[10] row_n[10]
+ adc_array_wafflecap_8_0[9|9]/sample vcm col_n[20] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|20] adc_array_wafflecap_8_0[10|9]/sample_n rowon_n[11]
+ row_n[11] adc_array_wafflecap_8_0[10|9]/sample vcm col_n[20] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|20] adc_array_wafflecap_8_0[11|9]/sample_n rowon_n[12]
+ row_n[12] adc_array_wafflecap_8_0[11|9]/sample vcm col_n[20] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|20] adc_array_wafflecap_8_0[12|9]/sample_n rowon_n[13]
+ row_n[13] adc_array_wafflecap_8_0[12|9]/sample vcm col_n[20] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|20] adc_array_wafflecap_8_0[13|9]/sample_n rowon_n[14]
+ row_n[14] adc_array_wafflecap_8_0[13|9]/sample vcm col_n[20] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|20] adc_array_wafflecap_8_0[14|9]/sample_n rowon_n[15]
+ row_n[15] adc_array_wafflecap_8_0[14|9]/sample vcm col_n[20] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|21] adc_array_wafflecap_8_0[0|9]/sample_n rowon_n[1] row_n[1]
+ adc_array_wafflecap_8_0[0|9]/sample vcm col_n[21] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|21] adc_array_wafflecap_8_0[1|9]/sample_n rowon_n[2] row_n[2]
+ adc_array_wafflecap_8_0[1|9]/sample vcm col_n[21] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|21] adc_array_wafflecap_8_0[2|9]/sample_n rowon_n[3] row_n[3]
+ adc_array_wafflecap_8_0[2|9]/sample vcm col_n[21] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|21] adc_array_wafflecap_8_0[3|9]/sample_n rowon_n[4] row_n[4]
+ adc_array_wafflecap_8_0[3|9]/sample vcm col_n[21] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|21] adc_array_wafflecap_8_0[4|9]/sample_n rowon_n[5] row_n[5]
+ adc_array_wafflecap_8_0[4|9]/sample vcm col_n[21] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|21] adc_array_wafflecap_8_0[5|9]/sample_n rowon_n[6] row_n[6]
+ adc_array_wafflecap_8_0[5|9]/sample vcm col_n[21] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|21] adc_array_wafflecap_8_0[6|9]/sample_n rowon_n[7] row_n[7]
+ adc_array_wafflecap_8_0[6|9]/sample vcm col_n[21] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|21] adc_array_wafflecap_8_0[7|9]/sample_n rowon_n[8] row_n[8]
+ adc_array_wafflecap_8_0[7|9]/sample vcm col_n[21] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|21] adc_array_wafflecap_8_0[8|9]/sample_n rowon_n[9] row_n[9]
+ adc_array_wafflecap_8_0[8|9]/sample vcm col_n[21] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|21] adc_array_wafflecap_8_0[9|9]/sample_n rowon_n[10] row_n[10]
+ adc_array_wafflecap_8_0[9|9]/sample vcm col_n[21] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|21] adc_array_wafflecap_8_0[10|9]/sample_n rowon_n[11]
+ row_n[11] adc_array_wafflecap_8_0[10|9]/sample vcm col_n[21] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|21] adc_array_wafflecap_8_0[11|9]/sample_n rowon_n[12]
+ row_n[12] adc_array_wafflecap_8_0[11|9]/sample vcm col_n[21] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|21] adc_array_wafflecap_8_0[12|9]/sample_n rowon_n[13]
+ row_n[13] adc_array_wafflecap_8_0[12|9]/sample vcm col_n[21] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|21] adc_array_wafflecap_8_0[13|9]/sample_n rowon_n[14]
+ row_n[14] adc_array_wafflecap_8_0[13|9]/sample vcm col_n[21] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|21] adc_array_wafflecap_8_0[14|9]/sample_n rowon_n[15]
+ row_n[15] adc_array_wafflecap_8_0[14|9]/sample vcm col_n[21] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|22] adc_array_wafflecap_8_0[0|9]/sample_n rowon_n[1] row_n[1]
+ adc_array_wafflecap_8_0[0|9]/sample vcm col_n[22] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|22] adc_array_wafflecap_8_0[1|9]/sample_n rowon_n[2] row_n[2]
+ adc_array_wafflecap_8_0[1|9]/sample vcm col_n[22] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|22] adc_array_wafflecap_8_0[2|9]/sample_n rowon_n[3] row_n[3]
+ adc_array_wafflecap_8_0[2|9]/sample vcm col_n[22] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|22] adc_array_wafflecap_8_0[3|9]/sample_n rowon_n[4] row_n[4]
+ adc_array_wafflecap_8_0[3|9]/sample vcm col_n[22] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|22] adc_array_wafflecap_8_0[4|9]/sample_n rowon_n[5] row_n[5]
+ adc_array_wafflecap_8_0[4|9]/sample vcm col_n[22] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|22] adc_array_wafflecap_8_0[5|9]/sample_n rowon_n[6] row_n[6]
+ adc_array_wafflecap_8_0[5|9]/sample vcm col_n[22] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|22] adc_array_wafflecap_8_0[6|9]/sample_n rowon_n[7] row_n[7]
+ adc_array_wafflecap_8_0[6|9]/sample vcm col_n[22] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|22] adc_array_wafflecap_8_0[7|9]/sample_n rowon_n[8] row_n[8]
+ adc_array_wafflecap_8_0[7|9]/sample vcm col_n[22] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|22] adc_array_wafflecap_8_0[8|9]/sample_n rowon_n[9] row_n[9]
+ adc_array_wafflecap_8_0[8|9]/sample vcm col_n[22] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|22] adc_array_wafflecap_8_0[9|9]/sample_n rowon_n[10] row_n[10]
+ adc_array_wafflecap_8_0[9|9]/sample vcm col_n[22] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|22] adc_array_wafflecap_8_0[10|9]/sample_n rowon_n[11]
+ row_n[11] adc_array_wafflecap_8_0[10|9]/sample vcm col_n[22] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|22] adc_array_wafflecap_8_0[11|9]/sample_n rowon_n[12]
+ row_n[12] adc_array_wafflecap_8_0[11|9]/sample vcm col_n[22] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|22] adc_array_wafflecap_8_0[12|9]/sample_n rowon_n[13]
+ row_n[13] adc_array_wafflecap_8_0[12|9]/sample vcm col_n[22] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|22] adc_array_wafflecap_8_0[13|9]/sample_n rowon_n[14]
+ row_n[14] adc_array_wafflecap_8_0[13|9]/sample vcm col_n[22] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|22] adc_array_wafflecap_8_0[14|9]/sample_n rowon_n[15]
+ row_n[15] adc_array_wafflecap_8_0[14|9]/sample vcm col_n[22] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|23] adc_array_wafflecap_8_0[0|9]/sample_n rowon_n[1] row_n[1]
+ adc_array_wafflecap_8_0[0|9]/sample vcm col_n[23] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|23] adc_array_wafflecap_8_0[1|9]/sample_n rowon_n[2] row_n[2]
+ adc_array_wafflecap_8_0[1|9]/sample vcm col_n[23] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|23] adc_array_wafflecap_8_0[2|9]/sample_n rowon_n[3] row_n[3]
+ adc_array_wafflecap_8_0[2|9]/sample vcm col_n[23] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|23] adc_array_wafflecap_8_0[3|9]/sample_n rowon_n[4] row_n[4]
+ adc_array_wafflecap_8_0[3|9]/sample vcm col_n[23] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|23] adc_array_wafflecap_8_0[4|9]/sample_n rowon_n[5] row_n[5]
+ adc_array_wafflecap_8_0[4|9]/sample vcm col_n[23] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|23] adc_array_wafflecap_8_0[5|9]/sample_n rowon_n[6] row_n[6]
+ adc_array_wafflecap_8_0[5|9]/sample vcm col_n[23] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|23] adc_array_wafflecap_8_0[6|9]/sample_n rowon_n[7] row_n[7]
+ adc_array_wafflecap_8_0[6|9]/sample vcm col_n[23] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|23] adc_array_wafflecap_8_0[7|9]/sample_n rowon_n[8] row_n[8]
+ adc_array_wafflecap_8_0[7|9]/sample vcm col_n[23] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|23] adc_array_wafflecap_8_0[8|9]/sample_n rowon_n[9] row_n[9]
+ adc_array_wafflecap_8_0[8|9]/sample vcm col_n[23] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|23] adc_array_wafflecap_8_0[9|9]/sample_n rowon_n[10] row_n[10]
+ adc_array_wafflecap_8_0[9|9]/sample vcm col_n[23] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|23] adc_array_wafflecap_8_0[10|9]/sample_n rowon_n[11]
+ row_n[11] adc_array_wafflecap_8_0[10|9]/sample vcm col_n[23] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|23] adc_array_wafflecap_8_0[11|9]/sample_n rowon_n[12]
+ row_n[12] adc_array_wafflecap_8_0[11|9]/sample vcm col_n[23] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|23] adc_array_wafflecap_8_0[12|9]/sample_n rowon_n[13]
+ row_n[13] adc_array_wafflecap_8_0[12|9]/sample vcm col_n[23] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|23] adc_array_wafflecap_8_0[13|9]/sample_n rowon_n[14]
+ row_n[14] adc_array_wafflecap_8_0[13|9]/sample vcm col_n[23] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|23] adc_array_wafflecap_8_0[14|9]/sample_n rowon_n[15]
+ row_n[15] adc_array_wafflecap_8_0[14|9]/sample vcm col_n[23] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|24] adc_array_wafflecap_8_0[0|9]/sample_n rowon_n[1] row_n[1]
+ adc_array_wafflecap_8_0[0|9]/sample vcm col_n[24] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|24] adc_array_wafflecap_8_0[1|9]/sample_n rowon_n[2] row_n[2]
+ adc_array_wafflecap_8_0[1|9]/sample vcm col_n[24] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|24] adc_array_wafflecap_8_0[2|9]/sample_n rowon_n[3] row_n[3]
+ adc_array_wafflecap_8_0[2|9]/sample vcm col_n[24] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|24] adc_array_wafflecap_8_0[3|9]/sample_n rowon_n[4] row_n[4]
+ adc_array_wafflecap_8_0[3|9]/sample vcm col_n[24] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|24] adc_array_wafflecap_8_0[4|9]/sample_n rowon_n[5] row_n[5]
+ adc_array_wafflecap_8_0[4|9]/sample vcm col_n[24] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|24] adc_array_wafflecap_8_0[5|9]/sample_n rowon_n[6] row_n[6]
+ adc_array_wafflecap_8_0[5|9]/sample vcm col_n[24] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|24] adc_array_wafflecap_8_0[6|9]/sample_n rowon_n[7] row_n[7]
+ adc_array_wafflecap_8_0[6|9]/sample vcm col_n[24] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|24] adc_array_wafflecap_8_0[7|9]/sample_n rowon_n[8] row_n[8]
+ adc_array_wafflecap_8_0[7|9]/sample vcm col_n[24] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|24] adc_array_wafflecap_8_0[8|9]/sample_n rowon_n[9] row_n[9]
+ adc_array_wafflecap_8_0[8|9]/sample vcm col_n[24] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|24] adc_array_wafflecap_8_0[9|9]/sample_n rowon_n[10] row_n[10]
+ adc_array_wafflecap_8_0[9|9]/sample vcm col_n[24] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|24] adc_array_wafflecap_8_0[10|9]/sample_n rowon_n[11]
+ row_n[11] adc_array_wafflecap_8_0[10|9]/sample vcm col_n[24] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|24] adc_array_wafflecap_8_0[11|9]/sample_n rowon_n[12]
+ row_n[12] adc_array_wafflecap_8_0[11|9]/sample vcm col_n[24] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|24] adc_array_wafflecap_8_0[12|9]/sample_n rowon_n[13]
+ row_n[13] adc_array_wafflecap_8_0[12|9]/sample vcm col_n[24] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|24] adc_array_wafflecap_8_0[13|9]/sample_n rowon_n[14]
+ row_n[14] adc_array_wafflecap_8_0[13|9]/sample vcm col_n[24] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|24] adc_array_wafflecap_8_0[14|9]/sample_n rowon_n[15]
+ row_n[15] adc_array_wafflecap_8_0[14|9]/sample vcm col_n[24] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|25] adc_array_wafflecap_8_0[0|9]/sample_n rowon_n[1] row_n[1]
+ adc_array_wafflecap_8_0[0|9]/sample vcm col_n[25] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|25] adc_array_wafflecap_8_0[1|9]/sample_n rowon_n[2] row_n[2]
+ adc_array_wafflecap_8_0[1|9]/sample vcm col_n[25] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|25] adc_array_wafflecap_8_0[2|9]/sample_n rowon_n[3] row_n[3]
+ adc_array_wafflecap_8_0[2|9]/sample vcm col_n[25] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|25] adc_array_wafflecap_8_0[3|9]/sample_n rowon_n[4] row_n[4]
+ adc_array_wafflecap_8_0[3|9]/sample vcm col_n[25] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|25] adc_array_wafflecap_8_0[4|9]/sample_n rowon_n[5] row_n[5]
+ adc_array_wafflecap_8_0[4|9]/sample vcm col_n[25] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|25] adc_array_wafflecap_8_0[5|9]/sample_n rowon_n[6] row_n[6]
+ adc_array_wafflecap_8_0[5|9]/sample vcm col_n[25] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|25] adc_array_wafflecap_8_0[6|9]/sample_n rowon_n[7] row_n[7]
+ adc_array_wafflecap_8_0[6|9]/sample vcm col_n[25] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|25] adc_array_wafflecap_8_0[7|9]/sample_n rowon_n[8] row_n[8]
+ adc_array_wafflecap_8_0[7|9]/sample vcm col_n[25] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|25] adc_array_wafflecap_8_0[8|9]/sample_n rowon_n[9] row_n[9]
+ adc_array_wafflecap_8_0[8|9]/sample vcm col_n[25] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|25] adc_array_wafflecap_8_0[9|9]/sample_n rowon_n[10] row_n[10]
+ adc_array_wafflecap_8_0[9|9]/sample vcm col_n[25] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|25] adc_array_wafflecap_8_0[10|9]/sample_n rowon_n[11]
+ row_n[11] adc_array_wafflecap_8_0[10|9]/sample vcm col_n[25] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|25] adc_array_wafflecap_8_0[11|9]/sample_n rowon_n[12]
+ row_n[12] adc_array_wafflecap_8_0[11|9]/sample vcm col_n[25] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|25] adc_array_wafflecap_8_0[12|9]/sample_n rowon_n[13]
+ row_n[13] adc_array_wafflecap_8_0[12|9]/sample vcm col_n[25] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|25] adc_array_wafflecap_8_0[13|9]/sample_n rowon_n[14]
+ row_n[14] adc_array_wafflecap_8_0[13|9]/sample vcm col_n[25] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|25] adc_array_wafflecap_8_0[14|9]/sample_n rowon_n[15]
+ row_n[15] adc_array_wafflecap_8_0[14|9]/sample vcm col_n[25] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|26] adc_array_wafflecap_8_0[0|9]/sample_n rowon_n[1] row_n[1]
+ adc_array_wafflecap_8_0[0|9]/sample vcm col_n[26] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|26] adc_array_wafflecap_8_0[1|9]/sample_n rowon_n[2] row_n[2]
+ adc_array_wafflecap_8_0[1|9]/sample vcm col_n[26] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|26] adc_array_wafflecap_8_0[2|9]/sample_n rowon_n[3] row_n[3]
+ adc_array_wafflecap_8_0[2|9]/sample vcm col_n[26] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|26] adc_array_wafflecap_8_0[3|9]/sample_n rowon_n[4] row_n[4]
+ adc_array_wafflecap_8_0[3|9]/sample vcm col_n[26] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|26] adc_array_wafflecap_8_0[4|9]/sample_n rowon_n[5] row_n[5]
+ adc_array_wafflecap_8_0[4|9]/sample vcm col_n[26] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|26] adc_array_wafflecap_8_0[5|9]/sample_n rowon_n[6] row_n[6]
+ adc_array_wafflecap_8_0[5|9]/sample vcm col_n[26] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|26] adc_array_wafflecap_8_0[6|9]/sample_n rowon_n[7] row_n[7]
+ adc_array_wafflecap_8_0[6|9]/sample vcm col_n[26] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|26] adc_array_wafflecap_8_0[7|9]/sample_n rowon_n[8] row_n[8]
+ adc_array_wafflecap_8_0[7|9]/sample vcm col_n[26] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|26] adc_array_wafflecap_8_0[8|9]/sample_n rowon_n[9] row_n[9]
+ adc_array_wafflecap_8_0[8|9]/sample vcm col_n[26] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|26] adc_array_wafflecap_8_0[9|9]/sample_n rowon_n[10] row_n[10]
+ adc_array_wafflecap_8_0[9|9]/sample vcm col_n[26] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|26] adc_array_wafflecap_8_0[10|9]/sample_n rowon_n[11]
+ row_n[11] adc_array_wafflecap_8_0[10|9]/sample vcm col_n[26] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|26] adc_array_wafflecap_8_0[11|9]/sample_n rowon_n[12]
+ row_n[12] adc_array_wafflecap_8_0[11|9]/sample vcm col_n[26] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|26] adc_array_wafflecap_8_0[12|9]/sample_n rowon_n[13]
+ row_n[13] adc_array_wafflecap_8_0[12|9]/sample vcm col_n[26] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|26] adc_array_wafflecap_8_0[13|9]/sample_n rowon_n[14]
+ row_n[14] adc_array_wafflecap_8_0[13|9]/sample vcm col_n[26] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|26] adc_array_wafflecap_8_0[14|9]/sample_n rowon_n[15]
+ row_n[15] adc_array_wafflecap_8_0[14|9]/sample vcm col_n[26] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|27] adc_array_wafflecap_8_0[0|9]/sample_n rowon_n[1] row_n[1]
+ adc_array_wafflecap_8_0[0|9]/sample vcm col_n[27] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|27] adc_array_wafflecap_8_0[1|9]/sample_n rowon_n[2] row_n[2]
+ adc_array_wafflecap_8_0[1|9]/sample vcm col_n[27] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|27] adc_array_wafflecap_8_0[2|9]/sample_n rowon_n[3] row_n[3]
+ adc_array_wafflecap_8_0[2|9]/sample vcm col_n[27] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|27] adc_array_wafflecap_8_0[3|9]/sample_n rowon_n[4] row_n[4]
+ adc_array_wafflecap_8_0[3|9]/sample vcm col_n[27] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|27] adc_array_wafflecap_8_0[4|9]/sample_n rowon_n[5] row_n[5]
+ adc_array_wafflecap_8_0[4|9]/sample vcm col_n[27] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|27] adc_array_wafflecap_8_0[5|9]/sample_n rowon_n[6] row_n[6]
+ adc_array_wafflecap_8_0[5|9]/sample vcm col_n[27] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|27] adc_array_wafflecap_8_0[6|9]/sample_n rowon_n[7] row_n[7]
+ adc_array_wafflecap_8_0[6|9]/sample vcm col_n[27] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|27] adc_array_wafflecap_8_0[7|9]/sample_n rowon_n[8] row_n[8]
+ adc_array_wafflecap_8_0[7|9]/sample vcm col_n[27] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|27] adc_array_wafflecap_8_0[8|9]/sample_n rowon_n[9] row_n[9]
+ adc_array_wafflecap_8_0[8|9]/sample vcm col_n[27] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|27] adc_array_wafflecap_8_0[9|9]/sample_n rowon_n[10] row_n[10]
+ adc_array_wafflecap_8_0[9|9]/sample vcm col_n[27] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|27] adc_array_wafflecap_8_0[10|9]/sample_n rowon_n[11]
+ row_n[11] adc_array_wafflecap_8_0[10|9]/sample vcm col_n[27] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|27] adc_array_wafflecap_8_0[11|9]/sample_n rowon_n[12]
+ row_n[12] adc_array_wafflecap_8_0[11|9]/sample vcm col_n[27] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|27] adc_array_wafflecap_8_0[12|9]/sample_n rowon_n[13]
+ row_n[13] adc_array_wafflecap_8_0[12|9]/sample vcm col_n[27] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|27] adc_array_wafflecap_8_0[13|9]/sample_n rowon_n[14]
+ row_n[14] adc_array_wafflecap_8_0[13|9]/sample vcm col_n[27] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|27] adc_array_wafflecap_8_0[14|9]/sample_n rowon_n[15]
+ row_n[15] adc_array_wafflecap_8_0[14|9]/sample vcm col_n[27] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|28] adc_array_wafflecap_8_0[0|9]/sample_n rowon_n[1] row_n[1]
+ adc_array_wafflecap_8_0[0|9]/sample vcm col_n[28] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|28] adc_array_wafflecap_8_0[1|9]/sample_n rowon_n[2] row_n[2]
+ adc_array_wafflecap_8_0[1|9]/sample vcm col_n[28] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|28] adc_array_wafflecap_8_0[2|9]/sample_n rowon_n[3] row_n[3]
+ adc_array_wafflecap_8_0[2|9]/sample vcm col_n[28] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|28] adc_array_wafflecap_8_0[3|9]/sample_n rowon_n[4] row_n[4]
+ adc_array_wafflecap_8_0[3|9]/sample vcm col_n[28] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|28] adc_array_wafflecap_8_0[4|9]/sample_n rowon_n[5] row_n[5]
+ adc_array_wafflecap_8_0[4|9]/sample vcm col_n[28] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|28] adc_array_wafflecap_8_0[5|9]/sample_n rowon_n[6] row_n[6]
+ adc_array_wafflecap_8_0[5|9]/sample vcm col_n[28] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|28] adc_array_wafflecap_8_0[6|9]/sample_n rowon_n[7] row_n[7]
+ adc_array_wafflecap_8_0[6|9]/sample vcm col_n[28] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|28] adc_array_wafflecap_8_0[7|9]/sample_n rowon_n[8] row_n[8]
+ adc_array_wafflecap_8_0[7|9]/sample vcm col_n[28] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|28] adc_array_wafflecap_8_0[8|9]/sample_n rowon_n[9] row_n[9]
+ adc_array_wafflecap_8_0[8|9]/sample vcm col_n[28] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|28] adc_array_wafflecap_8_0[9|9]/sample_n rowon_n[10] row_n[10]
+ adc_array_wafflecap_8_0[9|9]/sample vcm col_n[28] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|28] adc_array_wafflecap_8_0[10|9]/sample_n rowon_n[11]
+ row_n[11] adc_array_wafflecap_8_0[10|9]/sample vcm col_n[28] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|28] adc_array_wafflecap_8_0[11|9]/sample_n rowon_n[12]
+ row_n[12] adc_array_wafflecap_8_0[11|9]/sample vcm col_n[28] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|28] adc_array_wafflecap_8_0[12|9]/sample_n rowon_n[13]
+ row_n[13] adc_array_wafflecap_8_0[12|9]/sample vcm col_n[28] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|28] adc_array_wafflecap_8_0[13|9]/sample_n rowon_n[14]
+ row_n[14] adc_array_wafflecap_8_0[13|9]/sample vcm col_n[28] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|28] adc_array_wafflecap_8_0[14|9]/sample_n rowon_n[15]
+ row_n[15] adc_array_wafflecap_8_0[14|9]/sample vcm col_n[28] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|29] adc_array_wafflecap_8_0[0|9]/sample_n rowon_n[1] row_n[1]
+ adc_array_wafflecap_8_0[0|9]/sample vcm col_n[29] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|29] adc_array_wafflecap_8_0[1|9]/sample_n rowon_n[2] row_n[2]
+ adc_array_wafflecap_8_0[1|9]/sample vcm col_n[29] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|29] adc_array_wafflecap_8_0[2|9]/sample_n rowon_n[3] row_n[3]
+ adc_array_wafflecap_8_0[2|9]/sample vcm col_n[29] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|29] adc_array_wafflecap_8_0[3|9]/sample_n rowon_n[4] row_n[4]
+ adc_array_wafflecap_8_0[3|9]/sample vcm col_n[29] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|29] adc_array_wafflecap_8_0[4|9]/sample_n rowon_n[5] row_n[5]
+ adc_array_wafflecap_8_0[4|9]/sample vcm col_n[29] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|29] adc_array_wafflecap_8_0[5|9]/sample_n rowon_n[6] row_n[6]
+ adc_array_wafflecap_8_0[5|9]/sample vcm col_n[29] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|29] adc_array_wafflecap_8_0[6|9]/sample_n rowon_n[7] row_n[7]
+ adc_array_wafflecap_8_0[6|9]/sample vcm col_n[29] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|29] adc_array_wafflecap_8_0[7|9]/sample_n rowon_n[8] row_n[8]
+ adc_array_wafflecap_8_0[7|9]/sample vcm col_n[29] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|29] adc_array_wafflecap_8_0[8|9]/sample_n rowon_n[9] row_n[9]
+ adc_array_wafflecap_8_0[8|9]/sample vcm col_n[29] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|29] adc_array_wafflecap_8_0[9|9]/sample_n rowon_n[10] row_n[10]
+ adc_array_wafflecap_8_0[9|9]/sample vcm col_n[29] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|29] adc_array_wafflecap_8_0[10|9]/sample_n rowon_n[11]
+ row_n[11] adc_array_wafflecap_8_0[10|9]/sample vcm col_n[29] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|29] adc_array_wafflecap_8_0[11|9]/sample_n rowon_n[12]
+ row_n[12] adc_array_wafflecap_8_0[11|9]/sample vcm col_n[29] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|29] adc_array_wafflecap_8_0[12|9]/sample_n rowon_n[13]
+ row_n[13] adc_array_wafflecap_8_0[12|9]/sample vcm col_n[29] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|29] adc_array_wafflecap_8_0[13|9]/sample_n rowon_n[14]
+ row_n[14] adc_array_wafflecap_8_0[13|9]/sample vcm col_n[29] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|29] adc_array_wafflecap_8_0[14|9]/sample_n rowon_n[15]
+ row_n[15] adc_array_wafflecap_8_0[14|9]/sample vcm col_n[29] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|30] adc_array_wafflecap_8_0[0|9]/sample_n rowon_n[1] row_n[1]
+ adc_array_wafflecap_8_0[0|9]/sample vcm col_n[30] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|30] adc_array_wafflecap_8_0[1|9]/sample_n rowon_n[2] row_n[2]
+ adc_array_wafflecap_8_0[1|9]/sample vcm col_n[30] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|30] adc_array_wafflecap_8_0[2|9]/sample_n rowon_n[3] row_n[3]
+ adc_array_wafflecap_8_0[2|9]/sample vcm col_n[30] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|30] adc_array_wafflecap_8_0[3|9]/sample_n rowon_n[4] row_n[4]
+ adc_array_wafflecap_8_0[3|9]/sample vcm col_n[30] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|30] adc_array_wafflecap_8_0[4|9]/sample_n rowon_n[5] row_n[5]
+ adc_array_wafflecap_8_0[4|9]/sample vcm col_n[30] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|30] adc_array_wafflecap_8_0[5|9]/sample_n rowon_n[6] row_n[6]
+ adc_array_wafflecap_8_0[5|9]/sample vcm col_n[30] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|30] adc_array_wafflecap_8_0[6|9]/sample_n rowon_n[7] row_n[7]
+ adc_array_wafflecap_8_0[6|9]/sample vcm col_n[30] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|30] adc_array_wafflecap_8_0[7|9]/sample_n rowon_n[8] row_n[8]
+ adc_array_wafflecap_8_0[7|9]/sample vcm col_n[30] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|30] adc_array_wafflecap_8_0[8|9]/sample_n rowon_n[9] row_n[9]
+ adc_array_wafflecap_8_0[8|9]/sample vcm col_n[30] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|30] adc_array_wafflecap_8_0[9|9]/sample_n rowon_n[10] row_n[10]
+ adc_array_wafflecap_8_0[9|9]/sample vcm col_n[30] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|30] adc_array_wafflecap_8_0[10|9]/sample_n rowon_n[11]
+ row_n[11] adc_array_wafflecap_8_0[10|9]/sample vcm col_n[30] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|30] adc_array_wafflecap_8_0[11|9]/sample_n rowon_n[12]
+ row_n[12] adc_array_wafflecap_8_0[11|9]/sample vcm col_n[30] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|30] adc_array_wafflecap_8_0[12|9]/sample_n rowon_n[13]
+ row_n[13] adc_array_wafflecap_8_0[12|9]/sample vcm col_n[30] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|30] adc_array_wafflecap_8_0[13|9]/sample_n rowon_n[14]
+ row_n[14] adc_array_wafflecap_8_0[13|9]/sample vcm col_n[30] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|30] adc_array_wafflecap_8_0[14|9]/sample_n rowon_n[15]
+ row_n[15] adc_array_wafflecap_8_0[14|9]/sample vcm col_n[30] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|31] adc_array_wafflecap_8_0[0|9]/sample_n rowon_n[1] row_n[1]
+ adc_array_wafflecap_8_0[0|9]/sample vcm col_n[31] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|31] adc_array_wafflecap_8_0[1|9]/sample_n rowon_n[2] row_n[2]
+ adc_array_wafflecap_8_0[1|9]/sample vcm col_n[31] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|31] adc_array_wafflecap_8_0[2|9]/sample_n rowon_n[3] row_n[3]
+ adc_array_wafflecap_8_0[2|9]/sample vcm col_n[31] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|31] adc_array_wafflecap_8_0[3|9]/sample_n rowon_n[4] row_n[4]
+ adc_array_wafflecap_8_0[3|9]/sample vcm col_n[31] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|31] adc_array_wafflecap_8_0[4|9]/sample_n rowon_n[5] row_n[5]
+ adc_array_wafflecap_8_0[4|9]/sample vcm col_n[31] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|31] adc_array_wafflecap_8_0[5|9]/sample_n rowon_n[6] row_n[6]
+ adc_array_wafflecap_8_0[5|9]/sample vcm col_n[31] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|31] adc_array_wafflecap_8_0[6|9]/sample_n rowon_n[7] row_n[7]
+ adc_array_wafflecap_8_0[6|9]/sample vcm col_n[31] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|31] adc_array_wafflecap_8_0[7|9]/sample_n rowon_n[8] row_n[8]
+ adc_array_wafflecap_8_0[7|9]/sample vcm col_n[31] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|31] adc_array_wafflecap_8_0[8|9]/sample_n rowon_n[9] row_n[9]
+ adc_array_wafflecap_8_0[8|9]/sample vcm col_n[31] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|31] adc_array_wafflecap_8_0[9|9]/sample_n rowon_n[10] row_n[10]
+ adc_array_wafflecap_8_0[9|9]/sample vcm col_n[31] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|31] adc_array_wafflecap_8_0[10|9]/sample_n rowon_n[11]
+ row_n[11] adc_array_wafflecap_8_0[10|9]/sample vcm col_n[31] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|31] adc_array_wafflecap_8_0[11|9]/sample_n rowon_n[12]
+ row_n[12] adc_array_wafflecap_8_0[11|9]/sample vcm col_n[31] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|31] adc_array_wafflecap_8_0[12|9]/sample_n rowon_n[13]
+ row_n[13] adc_array_wafflecap_8_0[12|9]/sample vcm col_n[31] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|31] adc_array_wafflecap_8_0[13|9]/sample_n rowon_n[14]
+ row_n[14] adc_array_wafflecap_8_0[13|9]/sample vcm col_n[31] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|31] adc_array_wafflecap_8_0[14|9]/sample_n rowon_n[15]
+ row_n[15] adc_array_wafflecap_8_0[14|9]/sample vcm col_n[31] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[0] adc_array_wafflecap_8_1[9]/sample_n rowon_n[0] row_n[0]
+ adc_array_wafflecap_8_1[9]/sample vcm col_n[1] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[1] adc_array_wafflecap_8_1[9]/sample_n rowon_n[0] row_n[0]
+ adc_array_wafflecap_8_1[9]/sample vcm col_n[2] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[2] adc_array_wafflecap_8_1[9]/sample_n rowon_n[0] row_n[0]
+ adc_array_wafflecap_8_1[9]/sample vcm col_n[3] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[3] adc_array_wafflecap_8_1[9]/sample_n rowon_n[0] row_n[0]
+ adc_array_wafflecap_8_1[9]/sample vcm col_n[4] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[4] adc_array_wafflecap_8_1[9]/sample_n rowon_n[0] row_n[0]
+ adc_array_wafflecap_8_1[9]/sample vcm col_n[5] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[5] adc_array_wafflecap_8_1[9]/sample_n rowon_n[0] row_n[0]
+ adc_array_wafflecap_8_1[9]/sample vcm col_n[6] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[6] adc_array_wafflecap_8_1[9]/sample_n rowon_n[0] row_n[0]
+ adc_array_wafflecap_8_1[9]/sample vcm col_n[7] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[7] adc_array_wafflecap_8_1[9]/sample_n rowon_n[0] row_n[0]
+ adc_array_wafflecap_8_1[9]/sample vcm col_n[8] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[8] adc_array_wafflecap_8_1[9]/sample_n rowon_n[0] row_n[0]
+ adc_array_wafflecap_8_1[9]/sample vcm col_n[9] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[9] adc_array_wafflecap_8_1[9]/sample_n rowon_n[0] row_n[0]
+ adc_array_wafflecap_8_1[9]/sample vcm col_n[10] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[10] adc_array_wafflecap_8_1[9]/sample_n rowon_n[0] row_n[0]
+ adc_array_wafflecap_8_1[9]/sample vcm col_n[11] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[11] adc_array_wafflecap_8_1[9]/sample_n rowon_n[0] row_n[0]
+ adc_array_wafflecap_8_1[9]/sample vcm col_n[12] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[12] adc_array_wafflecap_8_1[9]/sample_n rowon_n[0] row_n[0]
+ adc_array_wafflecap_8_1[9]/sample vcm col_n[13] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[13] adc_array_wafflecap_8_1[9]/sample_n rowon_n[0] row_n[0]
+ adc_array_wafflecap_8_1[9]/sample vcm col_n[14] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[14] adc_array_wafflecap_8_1[9]/sample_n rowon_n[0] row_n[0]
+ adc_array_wafflecap_8_1[9]/sample vcm col_n[15] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[15] adc_array_wafflecap_8_1[9]/sample_n rowon_n[0] row_n[0]
+ adc_array_wafflecap_8_1[9]/sample vcm col_n[16] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[16] adc_array_wafflecap_8_1[9]/sample_n rowon_n[0] row_n[0]
+ adc_array_wafflecap_8_1[9]/sample vcm col_n[17] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[17] adc_array_wafflecap_8_1[9]/sample_n rowon_n[0] row_n[0]
+ adc_array_wafflecap_8_1[9]/sample vcm col_n[18] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[18] adc_array_wafflecap_8_1[9]/sample_n rowon_n[0] row_n[0]
+ adc_array_wafflecap_8_1[9]/sample vcm col_n[19] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[19] adc_array_wafflecap_8_1[9]/sample_n rowon_n[0] row_n[0]
+ adc_array_wafflecap_8_1[9]/sample vcm col_n[20] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[20] adc_array_wafflecap_8_1[9]/sample_n rowon_n[0] row_n[0]
+ adc_array_wafflecap_8_1[9]/sample vcm col_n[21] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[21] adc_array_wafflecap_8_1[9]/sample_n rowon_n[0] row_n[0]
+ adc_array_wafflecap_8_1[9]/sample vcm col_n[22] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[22] adc_array_wafflecap_8_1[9]/sample_n rowon_n[0] row_n[0]
+ adc_array_wafflecap_8_1[9]/sample vcm col_n[23] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[23] adc_array_wafflecap_8_1[9]/sample_n rowon_n[0] row_n[0]
+ adc_array_wafflecap_8_1[9]/sample vcm col_n[24] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[24] adc_array_wafflecap_8_1[9]/sample_n rowon_n[0] row_n[0]
+ adc_array_wafflecap_8_1[9]/sample vcm col_n[25] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[25] adc_array_wafflecap_8_1[9]/sample_n rowon_n[0] row_n[0]
+ adc_array_wafflecap_8_1[9]/sample vcm col_n[26] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[26] adc_array_wafflecap_8_1[9]/sample_n rowon_n[0] row_n[0]
+ adc_array_wafflecap_8_1[9]/sample vcm col_n[27] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[27] adc_array_wafflecap_8_1[9]/sample_n rowon_n[0] row_n[0]
+ adc_array_wafflecap_8_1[9]/sample vcm col_n[28] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[28] adc_array_wafflecap_8_1[9]/sample_n rowon_n[0] row_n[0]
+ adc_array_wafflecap_8_1[9]/sample vcm col_n[29] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[29] adc_array_wafflecap_8_1[9]/sample_n rowon_n[0] row_n[0]
+ adc_array_wafflecap_8_1[9]/sample vcm col_n[30] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[30] adc_array_wafflecap_8_1[9]/sample_n rowon_n[0] row_n[0]
+ adc_array_wafflecap_8_1[9]/sample vcm col_n[31] ctop VDD VSS adc_array_wafflecap_8
Xadc_noise_decoup_cell1_0[0] VDD VSS VDD VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_0[1] VDD VSS VDD VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_0[2] VDD VSS VDD VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_0[3] VDD VSS VDD VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_0[4] VDD VSS VDD VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_0[5] VDD VSS VDD VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[0] VDD VSS VDD VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[1] VDD VSS VDD VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[2] VDD VSS VDD VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[3] VDD VSS VDD VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[4] VDD VSS VDD VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[5] VDD VSS VDD VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[6] VDD VSS VDD VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[7] VDD VSS VDD VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[8] VDD VSS VDD VSS VSS adc_noise_decoup_cell1
Xadc_array_wafflecap_4_0 VDD VSS VSS VSS vcm col_n[16] en_bit_n[2] ctop VDD VSS adc_array_wafflecap_4
Xadc_array_wafflecap_2_0 VDD VSS VSS VSS vcm col_n[15] en_bit_n[1] ctop VDD VSS adc_array_wafflecap_2
Xadc_array_wafflecap_dummy_0[0] adc_array_wafflecap_8_1[9]/sample_n rowon_n[0] row_n[0]
+ adc_array_wafflecap_8_1[9]/sample vcm VDD adc_array_wafflecap_dummy_0[0]/ctop VDD
+ VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_0[1] adc_array_wafflecap_8_0[0|9]/sample_n rowon_n[1] row_n[1]
+ adc_array_wafflecap_8_0[0|9]/sample vcm VDD adc_array_wafflecap_dummy_0[1]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_0[2] adc_array_wafflecap_8_0[1|9]/sample_n rowon_n[2] row_n[2]
+ adc_array_wafflecap_8_0[1|9]/sample vcm VDD adc_array_wafflecap_dummy_0[2]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_0[3] adc_array_wafflecap_8_0[2|9]/sample_n rowon_n[3] row_n[3]
+ adc_array_wafflecap_8_0[2|9]/sample vcm VDD adc_array_wafflecap_dummy_0[3]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_0[4] adc_array_wafflecap_8_0[3|9]/sample_n rowon_n[4] row_n[4]
+ adc_array_wafflecap_8_0[3|9]/sample vcm VDD adc_array_wafflecap_dummy_0[4]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_0[5] adc_array_wafflecap_8_0[4|9]/sample_n rowon_n[5] row_n[5]
+ adc_array_wafflecap_8_0[4|9]/sample vcm VDD adc_array_wafflecap_dummy_0[5]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_0[6] adc_array_wafflecap_8_0[5|9]/sample_n rowon_n[6] row_n[6]
+ adc_array_wafflecap_8_0[5|9]/sample vcm VDD adc_array_wafflecap_dummy_0[6]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_0[7] adc_array_wafflecap_8_0[6|9]/sample_n rowon_n[7] row_n[7]
+ adc_array_wafflecap_8_0[6|9]/sample vcm VDD adc_array_wafflecap_dummy_0[7]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_0[8] adc_array_wafflecap_8_0[7|9]/sample_n rowon_n[8] row_n[8]
+ adc_array_wafflecap_8_0[7|9]/sample vcm VDD adc_array_wafflecap_dummy_0[8]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_0[9] adc_array_wafflecap_8_0[8|9]/sample_n rowon_n[9] row_n[9]
+ adc_array_wafflecap_8_0[8|9]/sample vcm VDD adc_array_wafflecap_dummy_0[9]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_0[10] adc_array_wafflecap_8_0[9|9]/sample_n rowon_n[10]
+ row_n[10] adc_array_wafflecap_8_0[9|9]/sample vcm VDD adc_array_wafflecap_dummy_0[10]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_0[11] adc_array_wafflecap_8_0[10|9]/sample_n rowon_n[11]
+ row_n[11] adc_array_wafflecap_8_0[10|9]/sample vcm VDD adc_array_wafflecap_dummy_0[11]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_0[12] adc_array_wafflecap_8_0[11|9]/sample_n rowon_n[12]
+ row_n[12] adc_array_wafflecap_8_0[11|9]/sample vcm VDD adc_array_wafflecap_dummy_0[12]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_0[13] adc_array_wafflecap_8_0[12|9]/sample_n rowon_n[13]
+ row_n[13] adc_array_wafflecap_8_0[12|9]/sample vcm VDD adc_array_wafflecap_dummy_0[13]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_0[14] adc_array_wafflecap_8_0[13|9]/sample_n rowon_n[14]
+ row_n[14] adc_array_wafflecap_8_0[13|9]/sample vcm VDD adc_array_wafflecap_dummy_0[14]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_0[15] adc_array_wafflecap_8_0[14|9]/sample_n rowon_n[15]
+ row_n[15] adc_array_wafflecap_8_0[14|9]/sample vcm VDD adc_array_wafflecap_dummy_0[15]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_1[0] VDD VDD VDD VSS vcm VDD adc_array_wafflecap_dummy_1[0]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_1[1] VDD VDD VDD VSS vcm col_n[0] adc_array_wafflecap_dummy_1[1]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_1[2] VDD VDD VDD VSS vcm col_n[1] adc_array_wafflecap_dummy_1[2]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_1[3] VDD VDD VDD VSS vcm col_n[2] adc_array_wafflecap_dummy_1[3]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_1[4] VDD VDD VDD VSS vcm col_n[3] adc_array_wafflecap_dummy_1[4]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_1[5] VDD VDD VDD VSS vcm col_n[4] adc_array_wafflecap_dummy_1[5]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_1[6] VDD VDD VDD VSS vcm col_n[5] adc_array_wafflecap_dummy_1[6]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_1[7] VDD VDD VDD VSS vcm col_n[6] adc_array_wafflecap_dummy_1[7]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_1[8] VDD VDD VDD VSS vcm col_n[7] adc_array_wafflecap_dummy_1[8]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_1[9] VDD VDD VDD VSS vcm col_n[8] adc_array_wafflecap_dummy_1[9]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_1[10] VDD VDD VDD VSS vcm col_n[9] adc_array_wafflecap_dummy_1[10]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_1[11] VDD VDD VDD VSS vcm col_n[10] adc_array_wafflecap_dummy_1[11]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_1[12] VDD VDD VDD VSS vcm col_n[11] adc_array_wafflecap_dummy_1[12]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_1[13] VDD VDD VDD VSS vcm col_n[12] adc_array_wafflecap_dummy_1[13]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_1[14] VDD VDD VDD VSS vcm col_n[13] adc_array_wafflecap_dummy_1[14]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_1[15] VDD VDD VDD VSS vcm col_n[14] adc_array_wafflecap_dummy_1[15]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_1[16] VDD VDD VDD VSS vcm col_n[15] adc_array_wafflecap_dummy_1[16]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_1[17] VDD VDD VDD VSS vcm col_n[16] adc_array_wafflecap_dummy_1[17]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_1[18] VDD VDD VDD VSS vcm col_n[17] adc_array_wafflecap_dummy_1[18]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_1[19] VDD VDD VDD VSS vcm col_n[18] adc_array_wafflecap_dummy_1[19]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_1[20] VDD VDD VDD VSS vcm col_n[19] adc_array_wafflecap_dummy_1[20]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_1[21] VDD VDD VDD VSS vcm col_n[20] adc_array_wafflecap_dummy_1[21]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_1[22] VDD VDD VDD VSS vcm col_n[21] adc_array_wafflecap_dummy_1[22]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_1[23] VDD VDD VDD VSS vcm col_n[22] adc_array_wafflecap_dummy_1[23]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_1[24] VDD VDD VDD VSS vcm col_n[23] adc_array_wafflecap_dummy_1[24]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_1[25] VDD VDD VDD VSS vcm col_n[24] adc_array_wafflecap_dummy_1[25]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_1[26] VDD VDD VDD VSS vcm col_n[25] adc_array_wafflecap_dummy_1[26]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_1[27] VDD VDD VDD VSS vcm col_n[26] adc_array_wafflecap_dummy_1[27]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_1[28] VDD VDD VDD VSS vcm col_n[27] adc_array_wafflecap_dummy_1[28]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_1[29] VDD VDD VDD VSS vcm col_n[28] adc_array_wafflecap_dummy_1[29]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_1[30] VDD VDD VDD VSS vcm col_n[29] adc_array_wafflecap_dummy_1[30]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_1[31] VDD VDD VDD VSS vcm col_n[30] adc_array_wafflecap_dummy_1[31]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_1[32] VDD VDD VDD VSS vcm col_n[31] adc_array_wafflecap_dummy_1[32]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_1[33] VDD VDD VDD VSS vcm VDD adc_array_wafflecap_dummy_1[33]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_2 adc_array_wafflecap_8_1[9]/sample_n rowon_n[0] row_n[0]
+ adc_array_wafflecap_8_1[9]/sample vcm col_n[0] adc_array_wafflecap_dummy_2/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_3 VDD VSS VSS VSS vcm VDD adc_array_wafflecap_dummy_3/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_4[0] VDD VSS VSS VSS vcm col_n[18] adc_array_wafflecap_dummy_4[0]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_4[1] VDD VSS VSS VSS vcm col_n[19] adc_array_wafflecap_dummy_4[1]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_4[2] VDD VSS VSS VSS vcm col_n[20] adc_array_wafflecap_dummy_4[2]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_4[3] VDD VSS VSS VSS vcm col_n[21] adc_array_wafflecap_dummy_4[3]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_4[4] VDD VSS VSS VSS vcm col_n[22] adc_array_wafflecap_dummy_4[4]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_4[5] VDD VSS VSS VSS vcm col_n[23] adc_array_wafflecap_dummy_4[5]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_4[6] VDD VSS VSS VSS vcm col_n[24] adc_array_wafflecap_dummy_4[6]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_4[7] VDD VSS VSS VSS vcm col_n[25] adc_array_wafflecap_dummy_4[7]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_4[8] VDD VSS VSS VSS vcm col_n[26] adc_array_wafflecap_dummy_4[8]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_4[9] VDD VSS VSS VSS vcm col_n[27] adc_array_wafflecap_dummy_4[9]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_4[10] VDD VSS VSS VSS vcm col_n[28] adc_array_wafflecap_dummy_4[10]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_4[11] VDD VSS VSS VSS vcm col_n[29] adc_array_wafflecap_dummy_4[11]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_4[12] VDD VSS VSS VSS vcm col_n[30] adc_array_wafflecap_dummy_4[12]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_gate_0 VDD VSS VSS VSS vcm col_n[31] analog_in sw sw_n ctop VDD
+ VSS col_n[31] adc_array_wafflecap_gate
.ends

.subckt sky130_fd_sc_hd__and3b_1 A_N B X C VGND VPWR VNB VPB
X0 a_109_93# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=1.0785e+11p pd=1.36e+06u as=3.5375e+11p ps=3.52e+06u w=420000u l=150000u
X1 X a_209_311# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=5.0705e+11p ps=5.41e+06u w=1e+06u l=150000u
X2 a_109_93# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1.087e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X3 a_296_53# a_109_93# a_209_311# VNB sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=1.07825e+11p ps=1.36e+06u w=420000u l=150000u
X4 VPWR C a_209_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.5725e+11p ps=2.99e+06u w=420000u l=150000u
X5 a_368_53# B a_296_53# VNB sky130_fd_pr__nfet_01v8 ad=1.071e+11p pd=1.35e+06u as=0p ps=0u w=420000u l=150000u
X6 X a_209_311# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X7 a_209_311# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VPWR a_109_93# a_209_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 VGND C a_368_53# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o22ai_1 A2 B1 Y A1 B2 VGND VPWR VNB VPB
X0 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=5.6875e+11p ps=5.65e+06u w=650000u l=150000u
X1 a_27_47# B2 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.8525e+11p ps=1.87e+06u w=650000u l=150000u
X2 VPWR A1 a_307_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=5.3e+11p pd=5.06e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X3 a_307_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.65e+11p ps=2.93e+06u w=1e+06u l=150000u
X4 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.25e+11p ps=2.45e+06u w=1e+06u l=150000u
X6 a_109_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__or2_4 X A B VGND VPWR VNB VPB
X0 a_121_297# B a_35_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X1 VPWR a_35_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=9.05e+11p pd=7.81e+06u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X2 X a_35_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 X a_35_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=7.4425e+11p ps=7.49e+06u w=650000u l=150000u
X4 X a_35_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VPWR a_35_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 X a_35_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND a_35_297# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR A a_121_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND a_35_297# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VGND A a_35_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X11 a_35_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__xor2_4 X B A VGND VPWR VNB VPB
X0 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1.345e+12p pd=1.269e+07u as=1.62e+12p ps=1.524e+07u w=1e+06u l=150000u
X1 a_806_47# B X VNB sky130_fd_pr__nfet_01v8 ad=8.645e+11p pd=9.16e+06u as=7.02e+11p ps=7.36e+06u w=650000u l=150000u
X2 a_806_47# B X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_112_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=7.02e+11p pd=7.36e+06u as=1.75175e+12p ps=1.839e+07u w=650000u l=150000u
X4 a_27_297# B a_112_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X5 a_806_297# a_112_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=1.8668e+12p pd=1.774e+07u as=8.2245e+11p ps=7.66e+06u w=1e+06u l=150000u
X6 VGND a_112_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 X B a_806_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 X a_112_47# a_806_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_112_47# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_806_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VGND A a_806_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 X B a_806_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VGND A a_806_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_806_297# a_112_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND A a_112_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_112_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 VGND A a_112_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 a_806_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VPWR B a_806_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 VGND B a_112_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 VGND B a_112_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 VPWR B a_806_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 a_806_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 a_806_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 a_27_297# B a_112_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 a_112_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X28 VGND a_112_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X29 a_806_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 a_112_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X31 a_112_47# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 VPWR A a_806_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X33 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X34 X a_112_47# a_806_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X35 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X36 a_806_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X37 X a_112_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X38 X a_112_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X39 VPWR A a_806_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__o32a_1 X A3 A1 A2 B1 B2 VPWR VGND VNB VPB
X0 a_77_199# B2 a_227_47# VNB sky130_fd_pr__nfet_01v8 ad=2.665e+11p pd=2.12e+06u as=6.565e+11p ps=5.92e+06u w=650000u l=150000u
X1 a_323_297# A2 a_227_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=3.9e+11p pd=2.78e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X2 a_227_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.6e+11p ps=5.12e+06u w=1e+06u l=150000u
X3 a_227_47# B1 a_77_199# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND a_77_199# X VNB sky130_fd_pr__nfet_01v8 ad=4.29e+11p pd=3.92e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X5 VPWR B1 a_539_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.1e+11p ps=2.82e+06u w=1e+06u l=150000u
X6 a_227_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR a_77_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.35e+11p ps=2.67e+06u w=1e+06u l=150000u
X8 a_77_199# A3 a_323_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=3.9e+11p pd=2.78e+06u as=0p ps=0u w=1e+06u l=150000u
X9 VGND A2 a_227_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_227_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_539_297# B2 a_77_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__buf_6 VPWR VGND X A VNB VPB
X0 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=1.33e+12p pd=1.266e+07u as=8.1e+11p ps=7.62e+06u w=1e+06u l=150000u
X1 a_161_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=8.645e+11p ps=9.16e+06u w=650000u l=150000u
X2 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND A a_161_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.265e+11p ps=5.52e+06u w=650000u l=150000u
X7 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VPWR A a_161_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X14 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_161_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand3_2 A Y B C VGND VPWR VNB VPB
X0 VGND C a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=3.705e+11p pd=3.74e+06u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u
X1 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=1.36e+12p pd=1.272e+07u as=8.1e+11p ps=7.62e+06u w=1e+06u l=150000u
X2 a_277_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=5.135e+11p pd=5.48e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X6 a_27_47# B a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_277_47# B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt adc_inverter out VDD VSS in
X0 out in VDD VDD sky130_fd_pr__pfet_01v8 ad=2.394e+11p pd=2.82e+06u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X1 VDD in out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 out in VSS VSS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
.ends

.subckt adc_nor B Q A VDD VSS
X0 a_312_106# A VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1 VDD B a_120_106# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2 Q B a_312_106# VDD sky130_fd_pr__pfet_01v8 ad=4.96e+11p pd=4.44e+06u as=0p ps=0u w=800000u l=150000u
X3 Q B VSS VSS sky130_fd_pr__nfet_01v8 ad=2.604e+11p pd=2.92e+06u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4 a_120_106# A Q VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5 VSS A Q VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt adc_nor_latch R QN Q S VDD VSS
X0 VSS S QN VSS sky130_fd_pr__nfet_01v8 ad=2.772e+11p pd=3e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1 Q QN VSS VSS sky130_fd_pr__nfet_01v8 ad=2.604e+11p pd=2.92e+06u as=0p ps=0u w=420000u l=150000u
X2 a_624_342# S QN VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=4.96e+11p ps=4.44e+06u w=800000u l=150000u
X3 VDD Q a_624_342# VDD sky130_fd_pr__pfet_01v8 ad=5.28e+11p pd=4.52e+06u as=0p ps=0u w=800000u l=150000u
X4 QN Q a_816_342# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5 a_816_342# S VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6 a_320_342# R VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7 VDD QN a_128_342# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8 Q QN a_320_342# VDD sky130_fd_pr__pfet_01v8 ad=4.96e+11p pd=4.44e+06u as=0p ps=0u w=800000u l=150000u
X9 VSS R Q VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_128_342# R Q VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X11 QN Q VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt adc_noise_decoup_cell2 nmoscap_bot nmoscap_top mimcap_bot mimcap_top pwell
X0 nmoscap_bot nmoscap_top nmoscap_bot pwell sky130_fd_pr__nfet_01v8 ad=2.576e+13p pd=7.64e+07u as=0p ps=0u w=1.84e+07u l=3.9e+06u
X1 mimcap_top mimcap_bot sky130_fd_pr__cap_mim_m3_1 l=5.1e+06u w=1.89e+07u
.ends

.subckt adc_comp_buffer out in VDD VSS
X0 out a_26_n216# VDD VDD sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.66e+06u as=6.4e+11p ps=5.28e+06u w=1e+06u l=150000u
X1 VDD a_26_n216# out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VSS a_26_n216# out VSS sky130_fd_pr__nfet_01v8 ad=3.2e+11p pd=3.28e+06u as=1.65e+11p ps=1.66e+06u w=500000u l=150000u
X3 VSS in a_26_n216# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.55e+11p ps=1.62e+06u w=500000u l=150000u
X4 VDD in a_26_n216# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X5 out a_26_n216# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
.ends

.subckt adc_comp_circuit inp inn outn outp clk nclk VGND VPWR
Xadc_noise_decoup_cell2_0 VGND on VGND VGND VGND adc_noise_decoup_cell2
Xadc_noise_decoup_cell2_1 VGND op VGND VGND VGND adc_noise_decoup_cell2
Xadc_comp_buffer_0 outp bp VPWR VGND adc_comp_buffer
Xadc_comp_buffer_1 outn bn VPWR VGND adc_comp_buffer
X0 bn op a_1306_n446# VPWR sky130_fd_pr__pfet_01v8 ad=1.24e+12p pd=9.24e+06u as=1.32e+12p ps=9.32e+06u w=2e+06u l=150000u
X1 VGND clk a_82_n1170# VGND sky130_fd_pr__nfet_01v8 ad=5.472e+13p pd=1.799e+08u as=4.025e+12p ps=3.144e+07u w=500000u l=150000u
X2 on inp a_82_n1170# VGND sky130_fd_pr__nfet_01v8_lvt ad=1.32e+12p pd=9.32e+06u as=0p ps=0u w=2e+06u l=150000u
X3 VGND clk a_82_n1170# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4 VGND nclk bp VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.6e+11p ps=4.66e+06u w=2e+06u l=150000u
X5 a_82_n1170# clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6 VPWR bp a_1306_n446# VPWR sky130_fd_pr__pfet_01v8 ad=3.985e+12p pd=3.268e+07u as=0p ps=0u w=2e+06u l=150000u
X7 a_82_n1170# inp on VGND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8 a_1820_n446# on bp VPWR sky130_fd_pr__pfet_01v8 ad=1.32e+12p pd=9.32e+06u as=1.24e+12p ps=9.24e+06u w=2e+06u l=150000u
X9 a_82_n1170# clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X10 a_1306_n446# op bn VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11 VGND clk a_82_n1170# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12 a_82_n1170# inn op VGND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.32e+12p ps=9.32e+06u w=2e+06u l=150000u
X13 a_1306_n446# bp VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14 VPWR bn a_1820_n446# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15 op inn a_82_n1170# VGND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X16 VGND clk a_82_n1170# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X17 bn nclk VGND VGND sky130_fd_pr__nfet_01v8 ad=6.6e+11p pd=4.66e+06u as=0p ps=0u w=2e+06u l=150000u
X18 a_82_n1170# inn op VGND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X19 a_82_n1170# clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X20 on inp a_82_n1170# VGND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X21 a_82_n1170# clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X22 VGND bp bn VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X23 bp on a_1820_n446# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X24 bp bn VGND VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X25 op inn a_82_n1170# VGND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X26 a_82_n1170# inp on VGND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X27 op clk VPWR VPWR sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=3.32e+06u as=0p ps=0u w=500000u l=150000u
X28 VPWR clk op VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X29 VPWR clk op VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X30 on clk VPWR VPWR sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=3.32e+06u as=0p ps=0u w=500000u l=150000u
X31 a_1820_n446# bn VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X32 op clk VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X33 on clk VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X34 VPWR clk on VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X35 VPWR clk on VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
.ends

.subckt adc_comp_latch VDD clk inp inn comp_trig latch_qn latch_q VSS
Xadc_inverter_0 adc_inverter_1/in VDD VSS clk adc_inverter
Xadc_inverter_1 adc_inverter_1/out VDD VSS adc_inverter_1/in adc_inverter
Xadc_nor_0 adc_nor_0/B comp_trig adc_nor_0/A VDD VSS adc_nor
Xadc_nor_latch_0 adc_nor_0/A latch_qn latch_q adc_nor_0/B VDD VSS adc_nor_latch
Xadc_comp_circuit_0 inp inn adc_nor_0/A adc_nor_0/B adc_inverter_1/out adc_inverter_1/in
+ VSS VDD adc_comp_circuit
.ends

.subckt sky130_fd_sc_hd__or3_2 A B X C VGND VPWR VNB VPB
X0 VPWR a_30_53# X VPB sky130_fd_pr__pfet_01v8_hvt ad=6.115e+11p pd=5.31e+06u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1 VGND a_30_53# X VNB sky130_fd_pr__nfet_01v8 ad=5.024e+11p pd=5.23e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X2 X a_30_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_112_297# C a_30_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X4 X a_30_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND A a_30_53# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.226e+11p ps=2.74e+06u w=420000u l=150000u
X6 a_30_53# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VGND C a_30_53# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_184_297# B a_112_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X9 VPWR A a_184_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__or3b_2 A B C_N X VPWR VGND VNB VPB
X0 a_388_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=5.88e+11p ps=5.35e+06u w=420000u l=150000u
X1 VPWR C_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X2 VGND a_176_21# X VNB sky130_fd_pr__nfet_01v8 ad=5.1765e+11p pd=5.33e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X3 X a_176_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR a_176_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X5 VGND B a_176_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.226e+11p ps=2.74e+06u w=420000u l=150000u
X6 X a_176_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_176_21# a_27_47# a_472_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X8 a_472_297# B a_388_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_176_21# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_176_21# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VGND C_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o311a_2 X A2 A3 A1 B1 C1 VPWR VGND VNB VPB
X0 X a_91_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=1.245e+12p ps=8.49e+06u w=1e+06u l=150000u
X1 a_91_21# C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=5.35e+11p pd=5.07e+06u as=0p ps=0u w=1e+06u l=150000u
X2 a_360_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=4.6475e+11p pd=4.03e+06u as=8.8725e+11p ps=6.63e+06u w=650000u l=150000u
X3 VPWR B1 a_91_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_360_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=3.5e+11p pd=2.7e+06u as=0p ps=0u w=1e+06u l=150000u
X5 VGND A2 a_360_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_360_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR a_91_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND a_91_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X9 X a_91_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_677_47# B1 a_360_47# VNB sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.72e+06u as=0p ps=0u w=650000u l=150000u
X11 a_460_297# A2 a_360_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=4.2e+11p pd=2.84e+06u as=0p ps=0u w=1e+06u l=150000u
X12 a_91_21# C1 a_677_47# VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X13 a_91_21# A3 a_460_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__or4b_2 C A X B D_N VPWR VGND VNB VPB
X0 a_176_21# C VGND VNB sky130_fd_pr__nfet_01v8 ad=2.52e+11p pd=2.88e+06u as=6.236e+11p ps=6.68e+06u w=420000u l=150000u
X1 VGND D_N a_27_53# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X2 VGND a_176_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X3 X a_176_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR a_176_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=6.753e+11p pd=5.99e+06u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X5 a_555_297# C a_483_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X6 a_176_21# a_27_53# a_555_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X7 X a_176_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_387_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X9 a_483_297# B a_387_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 VGND B a_176_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VGND a_27_53# a_176_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 VPWR D_N a_27_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X13 a_176_21# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o211ai_4 A1 B1 A2 C1 Y VGND VPWR VNB VPB
X0 VPWR A1 a_110_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=2.36e+12p pd=1.872e+07u as=1.12e+12p ps=1.024e+07u w=1e+06u l=150000u
X1 Y A2 a_110_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=1.65e+12p pd=1.53e+07u as=0p ps=0u w=1e+06u l=150000u
X2 a_806_47# B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=3.575e+11p pd=3.7e+06u as=1.3585e+12p ps=1.328e+07u w=650000u l=150000u
X3 a_110_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_110_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=7.345e+11p pd=7.46e+06u as=0p ps=0u w=650000u l=150000u
X6 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_110_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR A1 a_110_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_27_47# B1 a_1314_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.08e+11p ps=1.94e+06u w=650000u l=150000u
X12 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 Y A2 a_110_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 Y C1 a_978_47# VNB sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X20 Y C1 a_806_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 a_27_47# B1 a_806_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 a_110_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 a_806_47# C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X27 a_978_47# B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X28 a_1314_47# C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X29 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a31o_4 B1 A2 A3 A1 X VGND VPWR VNB VPB
X0 VPWR a_277_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=1.9e+12p pd=1.58e+07u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X1 X a_277_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 X a_277_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.39e+12p ps=1.278e+07u w=1e+06u l=150000u
X4 a_27_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_277_47# B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X6 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND a_277_47# X VNB sky130_fd_pr__nfet_01v8 ad=1.2415e+12p pd=1.032e+07u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u
X8 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND a_277_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_193_47# A2 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X12 a_361_47# A1 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u
X13 X a_277_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VGND A3 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.145e+11p ps=1.96e+06u w=650000u l=150000u
X15 X a_277_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_277_47# A1 a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 a_445_47# A2 a_361_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VGND B1 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_27_297# B1 a_277_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VPWR A3 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 VPWR a_277_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_109_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 a_277_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__or2_2 B X A VPWR VGND VNB VPB
X0 a_121_297# B a_39_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X1 X a_39_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=4.917e+11p ps=5.19e+06u w=650000u l=150000u
X2 VPWR a_39_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=5.715e+11p pd=5.23e+06u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X3 X a_39_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND a_39_297# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VPWR A a_121_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VGND A a_39_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X7 a_39_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o211a_2 C1 B1 A2 A1 X VPWR VGND VNB VPB
X0 a_27_47# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1e+12p pd=6e+06u as=9.35e+11p ps=7.87e+06u w=1e+06u l=150000u
X1 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=6.041e+11p pd=5.77e+06u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X2 VPWR C1 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR A1 a_373_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X4 a_182_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=3.4735e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u
X5 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u
X6 a_182_47# B1 a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.365e+11p ps=1.72e+06u w=650000u l=150000u
X7 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_373_297# A2 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_110_47# C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=150000u
X10 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VGND A1 a_182_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nor4_2 C D Y A B VGND VPWR VNB VPB
X0 a_281_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=8.3e+11p ps=7.66e+06u w=1e+06u l=150000u
X1 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=7.02e+11p pd=7.36e+06u as=1.066e+12p ps=1.108e+07u w=650000u l=150000u
X2 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X3 a_475_297# D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=8.1e+11p pd=7.62e+06u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X4 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y D a_475_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND D Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_475_297# C a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_281_297# C a_475_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_27_297# B a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 Y C VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o31a_1 X A2 B1 A1 A3 VGND VPWR VNB VPB
X0 a_103_199# B1 a_253_47# VNB sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=3.9e+11p ps=3.8e+06u w=650000u l=150000u
X1 VPWR a_103_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=7.35e+11p pd=5.47e+06u as=3.6e+11p ps=2.72e+06u w=1e+06u l=150000u
X2 a_337_297# A2 a_253_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=3.3e+11p pd=2.66e+06u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X3 a_103_199# A3 a_337_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=4.25e+11p pd=2.85e+06u as=0p ps=0u w=1e+06u l=150000u
X4 a_253_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR B1 a_103_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND a_103_199# X VNB sky130_fd_pr__nfet_01v8 ad=4.68e+11p pd=4.04e+06u as=2.34e+11p ps=2.02e+06u w=650000u l=150000u
X7 a_253_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_253_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VGND A2 a_253_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__and4b_1 VGND VPWR C A_N X D B VNB VPB
X0 a_297_47# a_27_47# a_193_413# VNB sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X1 a_369_47# B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=1.47e+11p pd=1.54e+06u as=0p ps=0u w=420000u l=150000u
X2 VPWR D a_193_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=6.511e+11p pd=6.09e+06u as=3.297e+11p ps=3.25e+06u w=420000u l=150000u
X3 X a_193_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=3.16e+11p ps=3.36e+06u w=650000u l=150000u
X4 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X5 VGND D a_469_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X6 X a_193_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR B a_193_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_193_413# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_193_413# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_469_47# C a_369_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__dlymetal6s2s_1 VPWR VGND A X VNB VPB
X0 a_558_47# a_381_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=8.445e+11p ps=7.95e+06u w=1e+06u l=150000u
X1 VGND X a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=5.82e+11p pd=5.85e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X2 a_841_47# a_664_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR A a_62_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X4 VGND A a_62_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X5 a_558_47# a_381_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X6 X a_62_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR X a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X8 a_841_47# a_664_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X9 X a_62_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X10 VPWR a_558_47# a_664_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X11 VGND a_558_47# a_664_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 Y C1 VGND VPWR VNB VPB
X0 a_286_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=5.46e+11p pd=5.58e+06u as=5.525e+11p ps=5.6e+06u w=650000u l=150000u
X1 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=1.09e+12p pd=1.018e+07u as=8.4e+11p ps=7.68e+06u w=1e+06u l=150000u
X2 a_286_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y A2 a_487_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.1e+11p ps=7.62e+06u w=1e+06u l=150000u
X4 VGND A1 a_286_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=5.525e+11p ps=5.6e+06u w=650000u l=150000u
X6 VGND A2 a_286_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_487_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_27_47# B1 a_286_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VPWR A1 a_487_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_27_47# C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_487_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_286_47# B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__nor2_4 Y A B VGND VPWR VNB VPB
X0 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=1.36e+12p ps=1.272e+07u w=1e+06u l=150000u
X1 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=7.02e+11p pd=7.36e+06u as=8.775e+11p ps=9.2e+06u w=650000u l=150000u
X2 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X5 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__nor3_4 A C B Y VGND VPWR VNB VPB
X0 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=1.35e+12p ps=1.27e+07u w=1e+06u l=150000u
X1 a_449_297# C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=1.08e+12p pd=1.016e+07u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X2 a_27_297# B a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=1.053e+12p pd=1.104e+07u as=1.2285e+12p ps=1.288e+07u w=650000u l=150000u
X4 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y C a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_449_297# C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 Y C a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_449_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 Y C VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 Y C VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_27_297# B a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 a_449_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__o2111ai_1 D1 C1 A2 A1 B1 Y VGND VPWR VNB VPB
X0 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=9.2e+11p pd=7.84e+06u as=6.85e+11p ps=5.37e+06u w=1e+06u l=150000u
X1 a_235_47# C1 a_163_47# VNB sky130_fd_pr__nfet_01v8 ad=2.535e+11p pd=2.08e+06u as=1.365e+11p ps=1.72e+06u w=650000u l=150000u
X2 a_343_47# B1 a_235_47# VNB sky130_fd_pr__nfet_01v8 ad=4.355e+11p pd=3.94e+06u as=0p ps=0u w=650000u l=150000u
X3 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_454_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=3.9e+11p pd=2.78e+06u as=0p ps=0u w=1e+06u l=150000u
X5 Y D1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR A1 a_454_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_163_47# D1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=150000u
X8 VGND A2 a_343_47# VNB sky130_fd_pr__nfet_01v8 ad=2.535e+11p pd=2.08e+06u as=0p ps=0u w=650000u l=150000u
X9 a_343_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a31oi_4 Y B1 A1 A3 A2 VPWR VGND VNB VPB
X0 a_27_47# A2 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=8.645e+11p pd=9.16e+06u as=7.02e+11p ps=7.36e+06u w=650000u l=150000u
X1 a_27_47# A2 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=1.62e+12p pd=1.524e+07u as=2.99e+12p ps=2.398e+07u w=1e+06u l=150000u
X3 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X5 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_27_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_445_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9.035e+11p ps=9.28e+06u w=650000u l=150000u
X12 VPWR A3 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_445_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=7.02e+11p pd=7.36e+06u as=0p ps=0u w=650000u l=150000u
X16 a_27_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 Y A1 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 Y A1 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 a_445_47# A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 a_445_47# A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X28 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X30 VPWR A3 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__and2_2 VPWR VGND A X B VNB VPB
X0 X a_61_75# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=3.9e+11p pd=2.78e+06u as=8.307e+11p ps=6.94e+06u w=1e+06u l=150000u
X1 VPWR a_61_75# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR B a_61_75# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X3 VGND B a_147_75# VNB sky130_fd_pr__nfet_01v8 ad=4.706e+11p pd=4.14e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X4 X a_61_75# VGND VNB sky130_fd_pr__nfet_01v8 ad=2.535e+11p pd=2.08e+06u as=0p ps=0u w=650000u l=150000u
X5 VGND a_61_75# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_61_75# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_147_75# A a_61_75# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a211oi_4 A2 A1 C1 Y B1 VPWR VGND VNB VPB
X0 Y A1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=1.105e+12p pd=1.12e+07u as=7.02e+11p ps=7.36e+06u w=650000u l=150000u
X1 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=1.2415e+12p pd=1.292e+07u as=0p ps=0u w=650000u l=150000u
X2 VGND A2 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=1.08e+12p pd=1.016e+07u as=1.87e+12p ps=1.774e+07u w=1e+06u l=150000u
X5 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_949_297# B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=3e+11p pd=2.6e+06u as=0p ps=0u w=1e+06u l=150000u
X8 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 Y C1 a_949_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=150000u
X10 a_781_297# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=5.5e+11p pd=5.1e+06u as=0p ps=0u w=1e+06u l=150000u
X11 a_27_297# B1 a_781_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VGND A2 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 Y A1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_781_297# B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_1301_297# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=3.1e+11p pd=2.62e+06u as=0p ps=0u w=1e+06u l=150000u
X16 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 Y C1 a_781_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 a_109_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_109_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_109_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X27 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 a_27_297# B1 a_1301_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X30 a_109_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X31 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nor3_2 C Y A B VGND VPWR VNB VPB
X0 Y C a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=7.9e+11p ps=7.58e+06u w=1e+06u l=150000u
X1 a_281_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.3e+11p ps=7.66e+06u w=1e+06u l=150000u
X2 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=5.265e+11p pd=5.52e+06u as=8.6125e+11p ps=9.15e+06u w=650000u l=150000u
X3 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 Y C VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_281_297# C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_27_297# B a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__or4_4 B C A D X VPWR VGND VNB VPB
X0 VPWR A a_304_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=9.2e+11p pd=7.84e+06u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1 a_304_297# B a_220_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X2 VGND C a_32_297# VNB sky130_fd_pr__nfet_01v8 ad=9.4575e+11p pd=9.41e+06u as=4.225e+11p ps=3.9e+06u w=650000u l=150000u
X3 a_220_297# C a_114_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.8e+11p ps=2.76e+06u w=1e+06u l=150000u
X4 a_32_297# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_32_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR a_32_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X7 X a_32_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND A a_32_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR a_32_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 X a_32_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u
X11 X a_32_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 X a_32_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_114_297# D a_32_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X14 VGND a_32_297# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 VGND a_32_297# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o31ai_1 Y A2 A1 A3 B1 VPWR VGND VNB VPB
X0 Y B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=2.21e+11p pd=1.98e+06u as=5.72e+11p ps=4.36e+06u w=650000u l=150000u
X1 Y A3 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=7.85e+11p pd=3.57e+06u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X2 a_193_297# A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X3 VGND A2 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=3.445e+11p pd=3.66e+06u as=0p ps=0u w=650000u l=150000u
X4 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=5.6e+11p pd=5.12e+06u as=0p ps=0u w=1e+06u l=150000u
X5 a_109_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_109_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a211oi_2 A2 C1 B1 Y A1 VPWR VGND VNB VPB
X0 VGND A2 a_485_47# VNB sky130_fd_pr__nfet_01v8 ad=7.085e+11p pd=7.38e+06u as=5.265e+11p ps=5.52e+06u w=650000u l=150000u
X1 VPWR A1 a_292_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=8.1e+11p pd=7.62e+06u as=8.4e+11p ps=7.68e+06u w=1e+06u l=150000u
X2 a_37_297# B1 a_292_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=8.1e+11p pd=7.62e+06u as=0p ps=0u w=1e+06u l=150000u
X3 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=5.46e+11p pd=5.58e+06u as=0p ps=0u w=650000u l=150000u
X4 a_485_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_292_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR A2 a_292_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_485_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_37_297# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X12 Y A1 a_485_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 Y C1 a_37_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_292_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_292_297# B1 a_37_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__or2b_1 A B_N X VGND VPWR VNB VPB
X0 a_219_297# a_27_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=5.1875e+11p ps=4.32e+06u w=420000u l=150000u
X1 VGND B_N a_27_53# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X2 VPWR A a_301_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=4.057e+11p pd=4.04e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X3 X a_219_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X4 a_301_297# a_27_53# a_219_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X5 X a_219_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X6 a_27_53# B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X7 VGND A a_219_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a221o_1 X B1 A1 B2 A2 VGND VPWR C1 VNB VPB
X0 a_465_47# A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=5.07e+11p ps=5.46e+06u w=650000u l=150000u
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=5.75e+11p ps=5.15e+06u w=1e+06u l=150000u
X2 a_109_297# B1 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=5.3e+11p pd=5.06e+06u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X3 a_193_297# B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=4.1925e+11p ps=3.89e+06u w=650000u l=150000u
X5 a_205_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.72e+06u as=0p ps=0u w=650000u l=150000u
X6 VPWR A2 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_193_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_27_47# B1 a_205_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_109_297# C1 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X10 VGND C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND A2 a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkinv_4 A Y VPWR VGND VNB VPB
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=8.4e+11p pd=7.68e+06u as=1.21e+12p ps=1.042e+07u w=1e+06u l=150000u
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=4.221e+11p pd=4.53e+06u as=2.352e+11p ps=2.8e+06u w=420000u l=150000u
X2 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand3b_1 B C A_N Y VGND VPWR VNB VPB
X0 Y a_53_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=5.5e+11p pd=5.1e+06u as=6.765e+11p ps=5.44e+06u w=1e+06u l=150000u
X1 a_232_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=2.005e+11p ps=1.97e+06u w=650000u l=150000u
X2 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR A_N a_53_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X4 VGND A_N a_53_93# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X5 a_316_47# B a_232_47# VNB sky130_fd_pr__nfet_01v8 ad=2.5025e+11p pd=2.07e+06u as=0p ps=0u w=650000u l=150000u
X6 Y a_53_93# a_316_47# VNB sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X7 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__nor4_1 D C Y A B VGND VPWR VNB VPB
X0 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=4.1275e+11p pd=3.87e+06u as=5.1675e+11p ps=5.49e+06u w=650000u l=150000u
X1 a_191_297# C a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=3.8e+11p pd=2.76e+06u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X2 VPWR A a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X3 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_297_297# B a_191_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_109_297# D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X7 Y D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand3_1 Y A C B VGND VPWR VNB VPB
X0 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=5.9e+11p pd=5.18e+06u as=5.3e+11p ps=5.06e+06u w=1e+06u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_193_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X3 Y A a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X4 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_109_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a2111oi_4 D1 C1 B1 A2 A1 Y VGND VPWR VNB VPB
X0 Y D1 VGND VNB sky130_fd_pr__nfet_01v8 ad=1.4495e+12p pd=1.486e+07u as=1.7615e+12p ps=1.712e+07u w=650000u l=150000u
X1 a_455_297# B1 a_821_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=1.12e+12p pd=1.024e+07u as=2.145e+12p ps=1.829e+07u w=1e+06u l=150000u
X2 a_28_297# D1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=1.365e+12p pd=1.273e+07u as=5.6e+11p ps=5.12e+06u w=1e+06u l=150000u
X3 a_821_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.14e+12p ps=1.028e+07u w=1e+06u l=150000u
X4 a_28_297# C1 a_455_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_455_297# C1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND D1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR A2 a_821_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 Y D1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND D1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 Y D1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_821_297# B1 a_455_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 Y D1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 a_1205_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=9.62e+11p pd=9.46e+06u as=0p ps=0u w=650000u l=150000u
X18 a_28_297# C1 a_455_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 a_1205_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 a_821_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 Y A1 a_1205_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 VPWR A1 a_821_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 Y A1 a_1205_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X27 a_1205_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X28 a_28_297# D1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 VGND A2 a_1205_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X30 a_455_297# B1 a_821_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 a_821_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 a_1205_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X33 VGND A2 a_1205_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X34 VPWR A1 a_821_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X35 a_821_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X36 VPWR A2 a_821_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X37 a_455_297# C1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X38 a_821_297# B1 a_455_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X39 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a2111oi_2 D1 C1 A2 A1 Y B1 VGND VPWR VNB VPB
X0 a_467_297# B1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=1.155e+12p pd=1.031e+07u as=8.65e+11p ps=7.73e+06u w=1e+06u l=150000u
X1 a_287_297# D1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X2 VPWR A2 a_467_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X3 a_923_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=9.1325e+11p ps=8.01e+06u w=650000u l=150000u
X4 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=9.3275e+11p pd=9.37e+06u as=0p ps=0u w=650000u l=150000u
X5 a_28_297# B1 a_467_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_28_297# C1 a_287_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 Y A1 a_923_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VGND A2 a_684_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.575e+11p ps=2.4e+06u w=650000u l=150000u
X10 Y D1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 Y D1 a_115_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X13 a_467_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VGND D1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 VPWR A1 a_467_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_115_297# C1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 a_467_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 a_684_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__or4_2 C A X B D VPWR VGND VNB VPB
X0 a_27_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=2.52e+11p pd=2.88e+06u as=6.246e+11p ps=6.63e+06u w=420000u l=150000u
X1 a_27_297# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_277_297# B a_205_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X3 VPWR A a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=6.015e+11p pd=5.29e+06u as=0p ps=0u w=420000u l=150000u
X4 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X5 a_205_297# C a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X6 VPWR a_27_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X7 VGND a_27_297# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND C a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_109_297# D a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X11 VGND A a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__or2b_2 A B_N X VPWR VGND VNB VPB
X0 VPWR A a_300_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=7.157e+11p pd=6.66e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X1 a_218_297# a_27_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=7.1815e+11p ps=6.23e+06u w=420000u l=150000u
X2 VGND B_N a_27_53# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X3 a_300_297# a_27_53# a_218_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X4 X a_218_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X5 VPWR a_218_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X6 X a_218_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND a_218_297# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_27_53# B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X9 VGND A a_218_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__dfstp_2 Q D VPWR SET_B CLK VGND VNB VPB
X0 VGND a_652_21# a_586_47# VNB sky130_fd_pr__nfet_01v8 ad=1.1373e+12p pd=1.19e+07u as=1.341e+11p ps=1.5e+06u w=420000u l=150000u
X1 a_956_413# a_476_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.5449e+12p ps=1.575e+07u w=420000u l=150000u
X2 a_1136_413# a_193_47# a_1028_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=2.73e+11p ps=2.98e+06u w=420000u l=150000u
X3 VPWR a_476_47# a_652_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X4 a_586_47# a_193_47# a_476_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.44e+11p ps=1.52e+06u w=360000u l=150000u
X5 a_1228_47# a_27_47# a_1028_413# VNB sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=1.47e+11p ps=1.54e+06u w=420000u l=150000u
X6 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X7 a_476_47# a_27_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.87e+11p ps=1.93e+06u w=360000u l=150000u
X8 a_1056_47# a_476_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X9 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.499e+11p pd=2.35e+06u as=0p ps=0u w=840000u l=150000u
X10 a_652_21# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VPWR a_1602_47# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X12 a_562_413# a_27_47# a_476_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=1.89e+11p pd=1.74e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X13 VGND a_1028_413# a_1602_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X14 VGND a_1602_47# Q VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X15 Q a_1602_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 a_1028_413# a_193_47# a_1056_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 a_476_47# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X19 VPWR a_1028_413# a_1602_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X20 VPWR a_652_21# a_562_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 Q a_1602_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 a_1028_413# a_27_47# a_956_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23 VPWR a_1178_261# a_1136_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X25 a_1178_261# a_1028_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.226e+11p pd=2.21e+06u as=0p ps=0u w=840000u l=150000u
X26 a_796_47# SET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X27 a_1300_47# a_1178_261# a_1228_47# VNB sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X28 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X29 a_1178_261# a_1028_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.404e+11p pd=1.6e+06u as=0p ps=0u w=540000u l=150000u
X30 a_652_21# a_476_47# a_796_47# VNB sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X31 VPWR SET_B a_1028_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X32 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X33 VGND SET_B a_1300_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a21oi_4 B1 A2 A1 Y VGND VPWR VNB VPB
X0 a_28_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=1.955e+12p pd=1.791e+07u as=5.6e+11p ps=5.12e+06u w=1e+06u l=150000u
X1 a_462_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=7.28e+11p pd=7.44e+06u as=7.28e+11p ps=7.44e+06u w=650000u l=150000u
X2 Y B1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9.165e+11p ps=9.32e+06u w=650000u l=150000u
X4 a_462_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_28_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.13e+12p ps=1.026e+07u w=1e+06u l=150000u
X6 a_462_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Y B1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y A1 a_462_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_28_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VPWR A2 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VGND A2 a_462_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_28_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VPWR A1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_28_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 VGND A2 a_462_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 VPWR A2 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 a_28_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 Y A1 a_462_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 a_462_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 VPWR A1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__a22o_2 A1 A2 X B2 B1 VPWR VGND VNB VPB
X0 VPWR a_27_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=8.45e+11p pd=7.69e+06u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1 VGND A2 a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=5.4925e+11p pd=5.59e+06u as=2.145e+11p ps=1.96e+06u w=650000u l=150000u
X2 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X3 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_27_297# B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=3.38e+11p pd=3.64e+06u as=1.495e+11p ps=1.76e+06u w=650000u l=150000u
X5 a_27_297# B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=5.2e+11p pd=5.04e+06u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X6 VGND a_27_297# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_381_47# A1 a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_109_297# B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_109_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_mm_sc_hd_dlyPoly5ns VNB VPB out VPWR VGND in
X0 a_851_95# in VGND VNB sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=1.0453e+12p ps=9.52e+06u w=420000u l=3.83e+06u
X1 a_1724_71# a_851_95# VGND VNB sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X2 VPWR out a_1724_71# VNB sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3 VGND out a_1783_329# VPB sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u
X4 a_1783_329# out VGND VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5 a_1724_71# out VPWR VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VGND a_851_95# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X7 a_1783_329# a_851_95# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.72e+11p ps=4.38e+06u w=800000u l=150000u
X8 out a_851_95# a_1783_329# VPB sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X9 a_851_95# in VPWR VPB sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X10 out a_851_95# a_1724_71# VNB sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nor2b_1 B_N Y A VGND VPWR VNB VPB
X0 Y a_74_47# a_265_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X1 VPWR B_N a_74_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=3.146e+11p pd=2.78e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X2 a_265_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=3.695e+11p ps=3.79e+06u w=650000u l=150000u
X4 VGND B_N a_74_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X5 VGND a_74_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt adc_clkgen_with_edgedetect clk_comp_out clk_dig_out dlycontrol1_in[0] dlycontrol1_in[1]
+ dlycontrol1_in[2] dlycontrol1_in[3] dlycontrol1_in[4] dlycontrol2_in[0] dlycontrol2_in[1]
+ dlycontrol2_in[2] dlycontrol2_in[3] dlycontrol2_in[4] dlycontrol3_in[0] dlycontrol3_in[1]
+ dlycontrol3_in[2] dlycontrol3_in[3] dlycontrol3_in[4] dlycontrol4_in[0] dlycontrol4_in[1]
+ dlycontrol4_in[2] dlycontrol4_in[3] dlycontrol4_in[4] dlycontrol4_in[5] ena_in enable_dlycontrol_in
+ ndecision_finish_in nsample_n_in nsample_n_out nsample_p_in nsample_p_out sample_n_in
+ sample_n_out sample_p_in sample_p_out start_conv_in VDD VSS
XFILLER_10_328 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_13_133 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_2.genblk1\[0\].control_invert dlycontrol2_in[0] clkgen.delay_155ns_2.bypass_enable_w\[0\]
+ VDD VSS VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_2_302 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_2.genblk1\[0\].dly_binary.out_mux VSS VDD clkgen.delay_155ns_2.genblk1\[0\].dly_binary.bypass_in
+ clkgen.clk_dig_out clkgen.delay_155ns_2.genblk1\[0\].dly_binary.signal_w\[1\] clkgen.delay_155ns_2.genblk1\[0\].dly_binary.out
+ VSS VDD sky130_fd_sc_hd__mux2_1
Xclkgen.delay_155ns_2.genblk1\[2\].dly_binary.out_mux VSS VDD clkgen.delay_155ns_2.genblk1\[2\].dly_binary.bypass_in
+ clkgen.delay_155ns_2.genblk1\[1\].dly_binary.out clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[4\]
+ clkgen.delay_155ns_2.genblk1\[2\].dly_binary.out VSS VDD sky130_fd_sc_hd__mux2_1
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.out_mux VSS VDD clkgen.delay_155ns_2.genblk1\[4\].dly_binary.bypass_in
+ clkgen.delay_155ns_2.genblk1\[3\].dly_binary.out clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[16\]
+ clkgen.clk_dig_delayed_w VSS VDD sky130_fd_sc_hd__mux2_1
XANTENNA_clkgen.delay_155ns_1.genblk1\[2\].control_invert_A dlycontrol1_in[2] VSS
+ VDD VDD VSS sky130_fd_sc_hd__diode_2
Xedgedetect.or1 edgedetect.start_conv_edge_w clkgen.enable_loop_in edgedetect.ena_in
+ VSS VDD VSS VDD sky130_fd_sc_hd__or2_1
Xclkgen.delay_155ns_3.genblk1\[0\].dly_binary.genblk1\[0\].delay_unit VSS VDD clkgen.delay_155ns_3.genblk1\[0\].dly_binary.signal_w\[1\]
+ VDD VSS clkgen.delay_155ns_3.genblk1\[0\].dly_binary.signal_w\[0\] sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[1\].bypass_enable VDD VSS edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.bypass_in
+ edgedetect.dly_315ns_1.bypass_enable_w\[1\] edgedetect.dly_315ns_1.enable_dlycontrol_w
+ VSS VDD sky130_fd_sc_hd__and2_1
XFILLER_13_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_3_282 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_16_164 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.delay_155ns_2.genblk1\[1\].control_invert_A dlycontrol2_in[1] VSS
+ VDD VDD VSS sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit VSS VDD clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[15\]
+ VDD VSS clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[14\] sky130_mm_sc_hd_dlyPoly5ns
XFILLER_3_57 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.delay_155ns_2.genblk1\[1\].dly_binary.and_bypass_switch_A_N clkgen.delay_155ns_2.genblk1\[1\].dly_binary.bypass_in
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_5_300 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_5_311 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xclkgen.delay_155ns_1.genblk1\[2\].bypass_enable VDD VSS clkgen.delay_155ns_1.genblk1\[2\].dly_binary.bypass_in
+ clkgen.delay_155ns_1.bypass_enable_w\[2\] clkgen.delay_155ns_1.enable_dlycontrol_w
+ VSS VDD sky130_fd_sc_hd__and2_1
Xclkgen.delay_155ns_2.genblk1\[3\].bypass_enable VDD VSS clkgen.delay_155ns_2.genblk1\[3\].dly_binary.bypass_in
+ clkgen.delay_155ns_2.bypass_enable_w\[3\] clkgen.delay_155ns_2.enable_dlycontrol_w
+ VSS VDD sky130_fd_sc_hd__and2_1
XFILLER_2_314 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[4\].bypass_enable VDD VSS clkgen.delay_155ns_3.genblk1\[4\].dly_binary.bypass_in
+ clkgen.delay_155ns_3.bypass_enable_w\[4\] clkgen.delay_155ns_3.enable_dlycontrol_w
+ VSS VDD sky130_fd_sc_hd__and2_1
XANTENNA_clkgen.delay_155ns_3.genblk1\[0\].control_invert_A dlycontrol3_in[0] VSS
+ VDD VDD VSS sky130_fd_sc_hd__diode_2
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[3\].delay_unit VSS VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[4\]
+ VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[3\] sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_clkgen.delay_155ns_3.genblk1\[4\].bypass_enable_A clkgen.delay_155ns_3.enable_dlycontrol_w
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_sampledly04_A nsample_n_in VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_18_32 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_11_276 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_11_243 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_19_321 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit VSS VDD clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[2\]
+ VDD VSS clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[1\] sky130_mm_sc_hd_dlyPoly5ns
XFILLER_4_206 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[1\].control_invert dlycontrol4_in[1] edgedetect.dly_315ns_1.bypass_enable_w\[1\]
+ VDD VSS VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_3_294 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_13_338 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_0_275 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[8\].delay_unit VSS VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[9\]
+ VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[8\] sky130_mm_sc_hd_dlyPoly5ns
XFILLER_9_139 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_8_194 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.delay_155ns_1.genblk1\[4\].dly_binary.and_bypass_switch_A_N clkgen.delay_155ns_1.genblk1\[4\].dly_binary.bypass_in
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit VSS VDD clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[13\]
+ VDD VSS clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[12\] sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit VSS VDD clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[7\]
+ VDD VSS clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[6\] sky130_mm_sc_hd_dlyPoly5ns
XFILLER_14_274 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_0_15 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_3_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xedgedetect.nor1 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.in edgedetect.start_conv_edge_w
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.out VSS VDD VSS VDD sky130_fd_sc_hd__nor2b_1
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[0\].delay_unit VSS VDD clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[1\]
+ VDD VSS clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[0\] sky130_mm_sc_hd_dlyPoly5ns
XFILLER_11_288 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_19_333 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_16_336 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[1\].control_invert dlycontrol3_in[1] clkgen.delay_155ns_3.bypass_enable_w\[1\]
+ VDD VSS VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_13_306 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit VSS VDD edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[4\]
+ VDD VSS edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[3\] sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit VSS VDD clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[6\]
+ VDD VSS clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[5\] sky130_mm_sc_hd_dlyPoly5ns
XFILLER_3_15 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit VSS VDD clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[2\]
+ VDD VSS clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[1\] sky130_mm_sc_hd_dlyPoly5ns
XFILLER_2_124 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[10\].delay_unit VSS VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[11\]
+ VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[10\] sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[10\].delay_unit VSS VDD clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[11\]
+ VDD VSS clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[10\] sky130_mm_sc_hd_dlyPoly5ns
XFILLER_7_216 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit VSS VDD edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[9\]
+ VDD VSS edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[8\] sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_edgedetect.dly_315ns_1.genblk1\[5\].bypass_enable_A edgedetect.dly_315ns_1.enable_dlycontrol_w
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_6_59 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit VSS VDD edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[12\]
+ VDD VSS edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[11\] sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit VSS VDD clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[7\]
+ VDD VSS clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[6\] sky130_mm_sc_hd_dlyPoly5ns
XFILLER_11_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_8_311 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit VSS VDD clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[5\]
+ VDD VSS clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[4\] sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.and_bypass_switch_A_N edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.bypass_in
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[0\].delay_unit VSS VDD clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[1\]
+ VDD VSS clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[0\] sky130_mm_sc_hd_dlyPoly5ns
XFILLER_12_181 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[15\].delay_unit VSS VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[16\]
+ VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[15\] sky130_mm_sc_hd_dlyPoly5ns
XFILLER_5_155 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit VSS VDD clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[16\]
+ VDD VSS clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[15\] sky130_mm_sc_hd_dlyPoly5ns
XFILLER_17_295 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_9_59 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xclkgen.nor1 clkgen.enable_loop_in clkgen.delay_155ns_3.genblk1\[0\].dly_binary.in
+ clkgen.clk_dig_delayed_w VSS VDD VSS VDD sky130_fd_sc_hd__nor2b_1
XANTENNA_sampledly02_A sample_n_in VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit VSS VDD clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[10\]
+ VDD VSS clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[9\] sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit VSS VDD edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[4\]
+ VDD VSS edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[3\] sky130_mm_sc_hd_dlyPoly5ns
XFILLER_10_290 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_1_93 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit VSS VDD clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[6\]
+ VDD VSS clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[5\] sky130_mm_sc_hd_dlyPoly5ns
XFILLER_6_16 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_19_187 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xclkgen.delay_155ns_3.genblk1\[2\].dly_binary.genblk1\[1\].delay_unit VSS VDD clkgen.delay_155ns_3.genblk1\[2\].dly_binary.signal_w\[2\]
+ VDD VSS clkgen.delay_155ns_3.genblk1\[2\].dly_binary.signal_w\[1\] sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_1.genblk1\[2\].control_invert dlycontrol1_in[2] clkgen.delay_155ns_1.bypass_enable_w\[2\]
+ VDD VSS VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_16_124 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[22\].delay_unit VSS VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[23\]
+ VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[22\] sky130_mm_sc_hd_dlyPoly5ns
XFILLER_8_323 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_0_245 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_223 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_3_28 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_8_164 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_18_208 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_12_59 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA_edgedetect.dly_315ns_1.enablebuffer_A enable_dlycontrol_in VSS VDD VDD VSS
+ sky130_fd_sc_hd__diode_2
XFILLER_14_211 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[27\].delay_unit VSS VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[28\]
+ VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[27\] sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_inbuf_3_A ndecision_finish_in VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_11_236 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_1_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xclkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit VSS VDD clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[5\]
+ VDD VSS clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[4\] sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_clkgen.delay_155ns_2.enablebuffer_A enable_dlycontrol_in VSS VDD VDD VSS
+ sky130_fd_sc_hd__diode_2
XANTENNA_clkgen.delay_155ns_1.genblk1\[1\].control_invert_A dlycontrol1_in[1] VSS
+ VDD VDD VSS sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_2.genblk1\[2\].dly_binary.genblk1\[0\].delay_unit VSS VDD clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[1\]
+ VDD VSS clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[0\] sky130_mm_sc_hd_dlyPoly5ns
XFILLER_10_70 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xclkgen.clkdig_inverter clkgen.delay_155ns_1.genblk1\[4\].dly_binary.out clkgen.clk_dig_out
+ VDD VSS VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_3_243 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_3_276 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_12_320 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_8_335 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_15_180 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA_clkgen.delay_155ns_2.genblk1\[0\].control_invert_A dlycontrol2_in[0] VSS
+ VDD VDD VSS sky130_fd_sc_hd__diode_2
XPHY_0 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_7_93 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_12_172 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_8_121 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_12_16 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_2_308 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_17_231 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit VSS VDD edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[4\]
+ VDD VSS edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[3\] sky130_mm_sc_hd_dlyPoly5ns
XFILLER_14_245 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit VSS VDD clkgen.delay_155ns_3.genblk1\[1\].dly_binary.signal_w\[2\]
+ VDD VSS clkgen.delay_155ns_3.genblk1\[1\].dly_binary.signal_w\[1\] sky130_mm_sc_hd_dlyPoly5ns
XFILLER_18_15 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_19_315 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_6_274 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_19_156 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_16_307 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_3_288 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.delay_155ns_1.genblk1\[4\].dly_binary.out_mux_S clkgen.delay_155ns_1.genblk1\[4\].dly_binary.bypass_in
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_12_332 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_0_214 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xedgedetect.dly_315ns_1.genblk1\[0\].dly_binary.out_mux VSS VDD edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.bypass_in
+ edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.in edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.signal_w\[1\]
+ edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.out VSS VDD sky130_fd_sc_hd__mux2_1
XPHY_1 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_7_50 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_edgedetect.dly_315ns_1.genblk1\[0\].bypass_enable_A edgedetect.dly_315ns_1.enable_dlycontrol_w
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xedgedetect.dly_315ns_1.genblk1\[2\].dly_binary.out_mux VSS VDD edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.bypass_in
+ edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.out edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[4\]
+ edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.out VSS VDD sky130_fd_sc_hd__mux2_1
Xedgedetect.dly_315ns_1.genblk1\[0\].dly_binary.and_bypass_switch edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.signal_w\[0\]
+ edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.bypass_in edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.in
+ VSS VDD VSS VDD sky130_fd_sc_hd__and2b_1
XFILLER_5_306 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xinbuf_1 VSS VDD edgedetect.ena_in ena_in VSS VDD sky130_fd_sc_hd__buf_1
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.out_mux VSS VDD edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.bypass_in
+ edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.out edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[16\]
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.out VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_5_125 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsampledly31 VDD VSS sample_p_3 sample_p_4 VSS VDD sky130_fd_sc_hd__dlymetal6s6s_1
XFILLER_4_62 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_2.genblk1\[1\].dly_binary.genblk1\[0\].delay_unit VSS VDD clkgen.delay_155ns_2.genblk1\[1\].dly_binary.signal_w\[1\]
+ VDD VSS clkgen.delay_155ns_2.genblk1\[1\].dly_binary.signal_w\[0\] sky130_mm_sc_hd_dlyPoly5ns
XFILLER_14_202 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_13_93 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_11_227 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_19_327 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_2.genblk1\[3\].control_invert dlycontrol2_in[3] clkgen.delay_155ns_2.bypass_enable_w\[3\]
+ VDD VSS VSS VDD sky130_fd_sc_hd__inv_2
Xedgedetect.dly_315ns_1.genblk1\[2\].bypass_enable VDD VSS edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.bypass_in
+ edgedetect.dly_315ns_1.bypass_enable_w\[2\] edgedetect.dly_315ns_1.enable_dlycontrol_w
+ VSS VDD sky130_fd_sc_hd__and2_1
XFILLER_1_63 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[10\].delay_unit VSS VDD clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[11\]
+ VDD VSS clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[10\] sky130_mm_sc_hd_dlyPoly5ns
XPHY_2 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xclkgen.delay_155ns_1.genblk1\[3\].bypass_enable VDD VSS clkgen.delay_155ns_1.genblk1\[3\].dly_binary.bypass_in
+ clkgen.delay_155ns_1.bypass_enable_w\[3\] clkgen.delay_155ns_1.enable_dlycontrol_w
+ VSS VDD sky130_fd_sc_hd__and2_1
Xclkgen.delay_155ns_2.genblk1\[4\].bypass_enable VDD VSS clkgen.delay_155ns_2.genblk1\[4\].dly_binary.bypass_in
+ clkgen.delay_155ns_2.bypass_enable_w\[4\] clkgen.delay_155ns_2.enable_dlycontrol_w
+ VSS VDD sky130_fd_sc_hd__and2_1
XFILLER_12_163 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xinbuf_2 VSS VDD edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.in start_conv_in VSS
+ VDD sky130_fd_sc_hd__buf_1
XANTENNA_clkgen.delay_155ns_1.genblk1\[2\].dly_binary.out_mux_S clkgen.delay_155ns_1.genblk1\[2\].dly_binary.bypass_in
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit VSS VDD clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[16\]
+ VDD VSS clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[15\] sky130_mm_sc_hd_dlyPoly5ns
XFILLER_17_288 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_17_222 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsampledly21 VDD VSS sample_p_2 sample_p_3 VSS VDD sky130_fd_sc_hd__dlymetal6s6s_1
Xsampledly32 VDD VSS sample_n_3 sample_n_4 VSS VDD sky130_fd_sc_hd__dlymetal6s6s_1
Xclkgen.delay_155ns_1.genblk1\[0\].dly_binary.out_mux VSS VDD clkgen.delay_155ns_1.genblk1\[0\].dly_binary.bypass_in
+ clkgen.delay_155ns_1.genblk1\[0\].dly_binary.in clkgen.delay_155ns_1.genblk1\[0\].dly_binary.signal_w\[1\]
+ clkgen.delay_155ns_1.genblk1\[0\].dly_binary.out VSS VDD sky130_fd_sc_hd__mux2_1
Xclkgen.delay_155ns_1.genblk1\[2\].dly_binary.out_mux VSS VDD clkgen.delay_155ns_1.genblk1\[2\].dly_binary.bypass_in
+ clkgen.delay_155ns_1.genblk1\[1\].dly_binary.out clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[4\]
+ clkgen.delay_155ns_1.genblk1\[2\].dly_binary.out VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_19_306 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.out_mux VSS VDD clkgen.delay_155ns_1.genblk1\[4\].dly_binary.bypass_in
+ clkgen.delay_155ns_1.genblk1\[3\].dly_binary.out clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[16\]
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.out VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_1_31 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[1\].dly_binary.and_bypass_switch edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.signal_w\[0\]
+ edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.bypass_in edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.out
+ VSS VDD VSS VDD sky130_fd_sc_hd__and2b_1
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[4\].delay_unit VSS VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[5\]
+ VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[4\] sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_inbuf_1_A ena_in VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_19_125 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_2_290 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_0_238 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_2.genblk1\[0\].dly_binary.genblk1\[0\].delay_unit VSS VDD clkgen.delay_155ns_2.genblk1\[0\].dly_binary.signal_w\[1\]
+ VDD VSS clkgen.delay_155ns_2.genblk1\[0\].dly_binary.signal_w\[0\] sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[2\].delay_unit VSS VDD clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[3\]
+ VDD VSS clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[2\] sky130_mm_sc_hd_dlyPoly5ns
XPHY_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_7_63 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_16_94 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xinbuf_3 VSS VDD clkgen.delay_155ns_1.genblk1\[0\].dly_binary.in ndecision_finish_in
+ VSS VDD sky130_fd_sc_hd__buf_1
XANTENNA_edgedetect.dly_315ns_1.genblk1\[5\].control_invert_A dlycontrol4_in[5] VSS
+ VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsampledly33 VDD VSS nsample_p_3 nsample_p_4 VSS VDD sky130_fd_sc_hd__dlymetal6s6s_1
Xsampledly11 VDD VSS sample_p_1 sample_p_2 VSS VDD sky130_fd_sc_hd__dlymetal6s6s_1
Xedgedetect.dly_315ns_1.genblk1\[4\].control_invert dlycontrol4_in[4] edgedetect.dly_315ns_1.bypass_enable_w\[4\]
+ VDD VSS VSS VDD sky130_fd_sc_hd__inv_2
Xsampledly22 VDD VSS sample_n_2 sample_n_3 VSS VDD sky130_fd_sc_hd__dlymetal6s6s_1
XANTENNA_clkgen.delay_155ns_1.genblk1\[0\].dly_binary.out_mux_S clkgen.delay_155ns_1.genblk1\[0\].dly_binary.bypass_in
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[9\].delay_unit VSS VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[10\]
+ VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[9\] sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_clkgen.delay_155ns_2.genblk1\[0\].dly_binary.and_bypass_switch_B clkgen.clk_dig_out
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_11_218 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit VSS VDD clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[14\]
+ VDD VSS clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[13\] sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit VSS VDD clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[8\]
+ VDD VSS clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[7\] sky130_mm_sc_hd_dlyPoly5ns
XFILLER_10_284 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_6_211 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA_clkgen.delay_155ns_1.genblk1\[2\].dly_binary.and_bypass_switch_A_N clkgen.delay_155ns_1.genblk1\[2\].dly_binary.bypass_in
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_19_94 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_10_41 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit VSS VDD clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[2\]
+ VDD VSS clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[1\] sky130_mm_sc_hd_dlyPoly5ns
XFILLER_3_236 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[0\].bypass_enable VDD VSS clkgen.delay_155ns_3.genblk1\[0\].dly_binary.bypass_in
+ clkgen.delay_155ns_3.bypass_enable_w\[0\] clkgen.delay_155ns_3.enable_dlycontrol_w
+ VSS VDD sky130_fd_sc_hd__and2_1
XFILLER_12_302 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.delay_155ns_3.genblk1\[2\].bypass_enable_A clkgen.delay_155ns_3.enable_dlycontrol_w
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_8_317 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[1\].dly_binary.out_mux VSS VDD clkgen.delay_155ns_3.genblk1\[1\].dly_binary.bypass_in
+ clkgen.delay_155ns_3.genblk1\[0\].dly_binary.out clkgen.delay_155ns_3.genblk1\[1\].dly_binary.signal_w\[2\]
+ clkgen.delay_155ns_3.genblk1\[1\].dly_binary.out VSS VDD sky130_fd_sc_hd__mux2_1
XPHY_4 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_16_62 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[3\].dly_binary.out_mux VSS VDD clkgen.delay_155ns_3.genblk1\[3\].dly_binary.bypass_in
+ clkgen.delay_155ns_3.genblk1\[2\].dly_binary.out clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[8\]
+ clkgen.delay_155ns_3.genblk1\[3\].dly_binary.out VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_17_279 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsampledly23 VDD VSS nsample_p_2 nsample_p_3 VSS VDD sky130_fd_sc_hd__dlymetal6s6s_1
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit VSS VDD edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[5\]
+ VDD VSS edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[4\] sky130_mm_sc_hd_dlyPoly5ns
Xsampledly01 VDD VSS sample_p_in sample_p_1 VSS VDD sky130_fd_sc_hd__dlymetal6s6s_1
Xclkgen.delay_155ns_3.genblk1\[4\].control_invert dlycontrol3_in[4] clkgen.delay_155ns_3.bypass_enable_w\[4\]
+ VDD VSS VSS VDD sky130_fd_sc_hd__inv_2
Xsampledly34 VDD VSS nsample_n_3 nsample_n_4 VSS VDD sky130_fd_sc_hd__dlymetal6s6s_1
Xsampledly12 VDD VSS sample_n_1 sample_n_2 VSS VDD sky130_fd_sc_hd__dlymetal6s6s_1
XFILLER_4_32 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_4_150 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_13_63 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit VSS VDD clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[7\]
+ VDD VSS clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[6\] sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[2\].dly_binary.and_bypass_switch edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[0\]
+ edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.bypass_in edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.out
+ VSS VDD VSS VDD sky130_fd_sc_hd__and2b_1
XFILLER_13_282 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit VSS VDD clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[3\]
+ VDD VSS clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[2\] sky130_mm_sc_hd_dlyPoly5ns
XFILLER_6_245 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_6_201 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[0\].delay_unit VSS VDD clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[1\]
+ VDD VSS clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[0\] sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_clkgen.delay_155ns_1.genblk1\[0\].control_invert_A dlycontrol1_in[0] VSS
+ VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_18_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_12_314 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[11\].delay_unit VSS VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[12\]
+ VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[11\] sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit VSS VDD clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[12\]
+ VDD VSS clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[11\] sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit VSS VDD edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[10\]
+ VDD VSS edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[9\] sky130_mm_sc_hd_dlyPoly5ns
XPHY_5 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_7_21 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit VSS VDD clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[8\]
+ VDD VSS clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[7\] sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit VSS VDD edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[13\]
+ VDD VSS edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[12\] sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit VSS VDD clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[6\]
+ VDD VSS clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[5\] sky130_mm_sc_hd_dlyPoly5ns
Xsampledly13 VDD VSS nsample_p_1 nsample_p_2 VSS VDD sky130_fd_sc_hd__dlymetal6s6s_1
Xsampledly24 VDD VSS nsample_n_2 nsample_n_3 VSS VDD sky130_fd_sc_hd__dlymetal6s6s_1
Xsampledly02 VDD VSS sample_n_in sample_n_1 VSS VDD sky130_fd_sc_hd__dlymetal6s6s_1
XFILLER_13_31 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit VSS VDD clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[2\]
+ VDD VSS clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[1\] sky130_mm_sc_hd_dlyPoly5ns
XFILLER_13_294 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_9_276 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_9_243 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[16\].delay_unit VSS VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[17\]
+ VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[16\] sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.and_bypass_switch_A_N edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.bypass_in
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_18_331 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_19_63 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_10_87 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_10_32 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_3_227 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_12_326 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[0\].control_invert dlycontrol1_in[0] clkgen.delay_155ns_1.bypass_enable_w\[0\]
+ VDD VSS VSS VDD sky130_fd_sc_hd__inv_2
Xedgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit VSS VDD edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[5\]
+ VDD VSS edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[4\] sky130_mm_sc_hd_dlyPoly5ns
XPHY_6 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_7_11 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit VSS VDD clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[7\]
+ VDD VSS clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[6\] sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_3.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit VSS VDD clkgen.delay_155ns_3.genblk1\[2\].dly_binary.signal_w\[3\]
+ VDD VSS clkgen.delay_155ns_3.genblk1\[2\].dly_binary.signal_w\[2\] sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_edgedetect.dly_315ns_1.genblk1\[3\].bypass_enable_A edgedetect.dly_315ns_1.enable_dlycontrol_w
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[23\].delay_unit VSS VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[24\]
+ VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[23\] sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[3\].dly_binary.and_bypass_switch edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[0\]
+ edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.bypass_in edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.out
+ VSS VDD VSS VDD sky130_fd_sc_hd__and2b_1
XFILLER_1_303 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xsampledly03 VDD VSS nsample_p_in nsample_p_1 VSS VDD sky130_fd_sc_hd__dlymetal6s6s_1
Xsampledly14 VDD VSS nsample_n_1 nsample_n_2 VSS VDD sky130_fd_sc_hd__dlymetal6s6s_1
Xclkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[0\].delay_unit VSS VDD clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[1\]
+ VDD VSS clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[0\] sky130_mm_sc_hd_dlyPoly5ns
XFILLER_4_174 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_8_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_1_155 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.out_mux_S edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.bypass_in
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_2_272 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_18_173 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[28\].delay_unit VSS VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[29\]
+ VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[28\] sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit VSS VDD clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[6\]
+ VDD VSS clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[5\] sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[30\].delay_unit VSS VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[31\]
+ VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[30\] sky130_mm_sc_hd_dlyPoly5ns
XFILLER_12_338 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_7 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA_clkgen.delay_155ns_2.genblk1\[0\].dly_binary.out_mux_S clkgen.delay_155ns_2.genblk1\[0\].dly_binary.bypass_in
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_2.genblk1\[2\].dly_binary.genblk1\[1\].delay_unit VSS VDD clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[2\]
+ VDD VSS clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[1\] sky130_mm_sc_hd_dlyPoly5ns
XFILLER_16_32 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_12_124 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_1_315 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_17_249 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsampledly04 VDD VSS nsample_n_in nsample_n_1 VSS VDD sky130_fd_sc_hd__dlymetal6s6s_1
XFILLER_4_164 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_3_218 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_5_281 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_19_32 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_2_284 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.enablebuffer VDD VSS edgedetect.dly_315ns_1.enable_dlycontrol_w
+ enable_dlycontrol_in VSS VDD sky130_fd_sc_hd__buf_4
XANTENNA_edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.out_mux_S edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.bypass_in
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_1.genblk1\[2\].dly_binary.genblk1\[0\].delay_unit VSS VDD clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[1\]
+ VDD VSS clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[0\] sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.and_bypass_switch edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[0\]
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.bypass_in edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.out
+ VSS VDD VSS VDD sky130_fd_sc_hd__and2b_1
XFILLER_16_3 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_8 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_4_335 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA_edgedetect.dly_315ns_1.genblk1\[4\].control_invert_A dlycontrol4_in[4] VSS
+ VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_1_327 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_4_121 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.enablebuffer VDD VSS clkgen.delay_155ns_1.enable_dlycontrol_w
+ enable_dlycontrol_in VSS VDD sky130_fd_sc_hd__buf_4
Xedgedetect.dly_315ns_1.genblk1\[3\].bypass_enable VDD VSS edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.bypass_in
+ edgedetect.dly_315ns_1.bypass_enable_w\[3\] edgedetect.dly_315ns_1.enable_dlycontrol_w
+ VSS VDD sky130_fd_sc_hd__and2_1
XFILLER_10_245 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_10_212 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_2.genblk1\[1\].control_invert dlycontrol2_in[1] clkgen.delay_155ns_2.bypass_enable_w\[1\]
+ VDD VSS VSS VDD sky130_fd_sc_hd__inv_2
Xclkgen.delay_155ns_2.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit VSS VDD clkgen.delay_155ns_2.genblk1\[1\].dly_binary.signal_w\[2\]
+ VDD VSS clkgen.delay_155ns_2.genblk1\[1\].dly_binary.signal_w\[1\] sky130_mm_sc_hd_dlyPoly5ns
XFILLER_18_164 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[4\].bypass_enable VDD VSS clkgen.delay_155ns_1.genblk1\[4\].dly_binary.bypass_in
+ clkgen.delay_155ns_1.bypass_enable_w\[4\] clkgen.delay_155ns_1.enable_dlycontrol_w
+ VSS VDD sky130_fd_sc_hd__and2_1
XFILLER_2_296 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[0\].dly_binary.and_bypass_switch clkgen.delay_155ns_3.genblk1\[0\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_3.genblk1\[0\].dly_binary.bypass_in clkgen.delay_155ns_3.genblk1\[0\].dly_binary.in
+ VSS VDD VSS VDD sky130_fd_sc_hd__and2b_1
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit VSS VDD clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[12\]
+ VDD VSS clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[11\] sky130_mm_sc_hd_dlyPoly5ns
XPHY_9 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA_edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.out_mux_S edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.bypass_in
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_clkgen.delay_155ns_1.genblk1\[4\].dly_binary.out_mux_A0 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[16\]
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_4_303 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.delay_155ns_1.enablebuffer_A enable_dlycontrol_in VSS VDD VDD VSS
+ sky130_fd_sc_hd__diode_2
XFILLER_19_292 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_1_339 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[0\].delay_unit VSS VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[1\]
+ VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[0\] sky130_mm_sc_hd_dlyPoly5ns
XFILLER_1_125 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_13_276 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_13_243 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_9_214 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_8_280 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xclkgen.delay_155ns_1.genblk1\[1\].dly_binary.genblk1\[0\].delay_unit VSS VDD clkgen.delay_155ns_1.genblk1\[1\].dly_binary.signal_w\[1\]
+ VDD VSS clkgen.delay_155ns_1.genblk1\[1\].dly_binary.signal_w\[0\] sky130_mm_sc_hd_dlyPoly5ns
XFILLER_18_313 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_6_3 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_5_294 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_15_338 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_15_305 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.and_bypass_switch edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[0\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.bypass_in edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.out
+ VSS VDD VSS VDD sky130_fd_sc_hd__and2b_1
XFILLER_12_308 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_11_90 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[5\].delay_unit VSS VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[6\]
+ VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[5\] sky130_mm_sc_hd_dlyPoly5ns
XFILLER_4_315 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xedgedetect.dly_315ns_1.genblk1\[2\].control_invert dlycontrol4_in[2] edgedetect.dly_315ns_1.bypass_enable_w\[2\]
+ VDD VSS VSS VDD sky130_fd_sc_hd__inv_2
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit VSS VDD clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[4\]
+ VDD VSS clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[3\] sky130_mm_sc_hd_dlyPoly5ns
XFILLER_16_274 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_4_16 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_13_288 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_10_203 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_18_325 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_2.genblk1\[0\].bypass_enable VDD VSS clkgen.delay_155ns_2.genblk1\[0\].dly_binary.bypass_in
+ clkgen.delay_155ns_2.bypass_enable_w\[0\] clkgen.delay_155ns_2.enable_dlycontrol_w
+ VSS VDD sky130_fd_sc_hd__and2_1
Xclkgen.delay_155ns_3.genblk1\[1\].dly_binary.and_bypass_switch clkgen.delay_155ns_3.genblk1\[1\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_3.genblk1\[1\].dly_binary.bypass_in clkgen.delay_155ns_3.genblk1\[0\].dly_binary.out
+ VSS VDD VSS VDD sky130_fd_sc_hd__and2b_1
Xclkgen.delay_155ns_3.genblk1\[1\].bypass_enable VDD VSS clkgen.delay_155ns_3.genblk1\[1\].dly_binary.bypass_in
+ clkgen.delay_155ns_3.bypass_enable_w\[1\] clkgen.delay_155ns_3.enable_dlycontrol_w
+ VSS VDD sky130_fd_sc_hd__and2_1
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit VSS VDD clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[9\]
+ VDD VSS clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[8\] sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_clkgen.delay_155ns_3.genblk1\[4\].control_invert_A dlycontrol3_in[4] VSS
+ VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_15_147 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit VSS VDD clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[15\]
+ VDD VSS clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[14\] sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_2.genblk1\[0\].dly_binary.and_bypass_switch clkgen.delay_155ns_2.genblk1\[0\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_2.genblk1\[0\].dly_binary.bypass_in clkgen.clk_dig_out VSS VDD
+ VSS VDD sky130_fd_sc_hd__and2b_1
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[0\].delay_unit VSS VDD edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[1\]
+ VDD VSS edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[0\] sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[2\].delay_unit VSS VDD clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[3\]
+ VDD VSS clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[2\] sky130_mm_sc_hd_dlyPoly5ns
XFILLER_14_3 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_7_187 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_7_154 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[0\].dly_binary.genblk1\[0\].delay_unit VSS VDD clkgen.delay_155ns_1.genblk1\[0\].dly_binary.signal_w\[1\]
+ VDD VSS clkgen.delay_155ns_1.genblk1\[0\].dly_binary.signal_w\[0\] sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_clkgen.delay_155ns_1.genblk1\[0\].dly_binary.and_bypass_switch_A_N clkgen.delay_155ns_1.genblk1\[0\].dly_binary.bypass_in
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_3.genblk1\[2\].control_invert dlycontrol3_in[2] clkgen.delay_155ns_3.bypass_enable_w\[2\]
+ VDD VSS VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_5_93 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_18_337 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit VSS VDD edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[6\]
+ VDD VSS edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[5\] sky130_mm_sc_hd_dlyPoly5ns
XFILLER_10_16 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit VSS VDD clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[8\]
+ VDD VSS clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[7\] sky130_mm_sc_hd_dlyPoly5ns
XFILLER_2_266 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit VSS VDD clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[4\]
+ VDD VSS clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[3\] sky130_mm_sc_hd_dlyPoly5ns
XFILLER_2_94 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_15_137 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_11_321 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit VSS VDD clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[2\]
+ VDD VSS clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[1\] sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[12\].delay_unit VSS VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[13\]
+ VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[12\] sky130_mm_sc_hd_dlyPoly5ns
XFILLER_8_82 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_2.genblk1\[1\].dly_binary.out_mux VSS VDD clkgen.delay_155ns_2.genblk1\[1\].dly_binary.bypass_in
+ clkgen.delay_155ns_2.genblk1\[0\].dly_binary.out clkgen.delay_155ns_2.genblk1\[1\].dly_binary.signal_w\[2\]
+ clkgen.delay_155ns_2.genblk1\[1\].dly_binary.out VSS VDD sky130_fd_sc_hd__mux2_1
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit VSS VDD clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[13\]
+ VDD VSS clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[12\] sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.and_bypass_switch_A_N edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.bypass_in
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_2.genblk1\[3\].dly_binary.out_mux VSS VDD clkgen.delay_155ns_2.genblk1\[3\].dly_binary.bypass_in
+ clkgen.delay_155ns_2.genblk1\[2\].dly_binary.out clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[8\]
+ clkgen.delay_155ns_2.genblk1\[3\].dly_binary.out VSS VDD sky130_fd_sc_hd__mux2_1
XANTENNA_clkgen.delay_155ns_3.genblk1\[0\].bypass_enable_A clkgen.delay_155ns_3.enable_dlycontrol_w
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_3.genblk1\[2\].dly_binary.and_bypass_switch clkgen.delay_155ns_3.genblk1\[2\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_3.genblk1\[2\].dly_binary.bypass_in clkgen.delay_155ns_3.genblk1\[1\].dly_binary.out
+ VSS VDD VSS VDD sky130_fd_sc_hd__and2b_1
XFILLER_0_183 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit VSS VDD edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[14\]
+ VDD VSS edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[13\] sky130_mm_sc_hd_dlyPoly5ns
XFILLER_12_290 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[0\].delay_unit VSS VDD edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[1\]
+ VDD VSS edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[0\] sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_2.genblk1\[1\].dly_binary.and_bypass_switch clkgen.delay_155ns_2.genblk1\[1\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_2.genblk1\[1\].dly_binary.bypass_in clkgen.delay_155ns_2.genblk1\[0\].dly_binary.out
+ VSS VDD VSS VDD sky130_fd_sc_hd__and2b_1
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit VSS VDD clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[7\]
+ VDD VSS clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[6\] sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit VSS VDD clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[3\]
+ VDD VSS clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[2\] sky130_mm_sc_hd_dlyPoly5ns
XFILLER_19_15 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_2_234 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_4_3 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_18_179 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_18_124 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[17\].delay_unit VSS VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[18\]
+ VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[17\] sky130_mm_sc_hd_dlyPoly5ns
XFILLER_2_62 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[0\].dly_binary.and_bypass_switch clkgen.delay_155ns_1.genblk1\[0\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_1.genblk1\[0\].dly_binary.bypass_in clkgen.delay_155ns_1.genblk1\[0\].dly_binary.in
+ VSS VDD VSS VDD sky130_fd_sc_hd__and2b_1
XFILLER_11_333 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_11_300 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_16_16 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_14_193 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit VSS VDD edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[6\]
+ VDD VSS edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[5\] sky130_mm_sc_hd_dlyPoly5ns
XFILLER_0_321 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xclkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit VSS VDD clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[8\]
+ VDD VSS clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[7\] sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_edgedetect.dly_315ns_1.genblk1\[3\].control_invert_A dlycontrol4_in[3] VSS
+ VDD VDD VSS sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_1.genblk1\[3\].control_invert dlycontrol1_in[3] clkgen.delay_155ns_1.bypass_enable_w\[3\]
+ VDD VSS VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_13_214 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit VSS VDD clkgen.delay_155ns_3.genblk1\[2\].dly_binary.signal_w\[4\]
+ VDD VSS clkgen.delay_155ns_3.genblk1\[2\].dly_binary.signal_w\[3\] sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[24\].delay_unit VSS VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[25\]
+ VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[24\] sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit VSS VDD clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[2\]
+ VDD VSS clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[1\] sky130_mm_sc_hd_dlyPoly5ns
XFILLER_5_243 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_7_338 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_7_305 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[29\].delay_unit VSS VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[30\]
+ VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[29\] sky130_mm_sc_hd_dlyPoly5ns
XFILLER_8_40 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_3_341 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xedgedetect.dly_315ns_1.genblk1\[2\].dly_binary.genblk1\[0\].delay_unit VSS VDD edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[1\]
+ VDD VSS edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[0\] sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_3.genblk1\[3\].dly_binary.and_bypass_switch clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_3.genblk1\[3\].dly_binary.bypass_in clkgen.delay_155ns_3.genblk1\[2\].dly_binary.out
+ VSS VDD VSS VDD sky130_fd_sc_hd__and2b_1
Xclkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit VSS VDD clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[7\]
+ VDD VSS clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[6\] sky130_mm_sc_hd_dlyPoly5ns
XFILLER_17_71 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_16_245 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[31\].delay_unit VSS VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[32\]
+ VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[31\] sky130_mm_sc_hd_dlyPoly5ns
XFILLER_0_333 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xclkgen.delay_155ns_2.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit VSS VDD clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[3\]
+ VDD VSS clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[2\] sky130_mm_sc_hd_dlyPoly5ns
XFILLER_12_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xclkgen.delay_155ns_2.genblk1\[2\].dly_binary.and_bypass_switch clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_2.genblk1\[2\].dly_binary.bypass_in clkgen.delay_155ns_2.genblk1\[1\].dly_binary.out
+ VSS VDD VSS VDD sky130_fd_sc_hd__and2b_1
XFILLER_8_274 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_5_63 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_18_307 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[1\].dly_binary.and_bypass_switch clkgen.delay_155ns_1.genblk1\[1\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_1.genblk1\[1\].dly_binary.bypass_in clkgen.delay_155ns_1.genblk1\[0\].dly_binary.out
+ VSS VDD VSS VDD sky130_fd_sc_hd__and2b_1
XFILLER_14_94 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_5_288 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_edgedetect.dly_315ns_1.genblk1\[1\].bypass_enable_A edgedetect.dly_315ns_1.enable_dlycontrol_w
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_14_310 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_2_214 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_2_225 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_17_192 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_1_291 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_sampledly03_A nsample_p_in VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_4_309 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_19_276 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_11_187 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_11_154 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_7_125 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[2\].dly_binary.genblk1\[1\].delay_unit VSS VDD clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[2\]
+ VDD VSS clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[1\] sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[4\].bypass_enable VDD VSS edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.bypass_in
+ edgedetect.dly_315ns_1.bypass_enable_w\[4\] edgedetect.dly_315ns_1.enable_dlycontrol_w
+ VSS VDD sky130_fd_sc_hd__and2_1
XFILLER_12_260 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_5_31 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.delay_155ns_2.genblk1\[4\].control_invert_A dlycontrol2_in[4] VSS
+ VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_18_319 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_14_84 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_2.enablebuffer VDD VSS clkgen.delay_155ns_2.enable_dlycontrol_w
+ enable_dlycontrol_in VSS VDD sky130_fd_sc_hd__buf_4
Xedgedetect.dly_315ns_1.genblk1\[1\].dly_binary.genblk1\[0\].delay_unit VSS VDD edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.signal_w\[1\]
+ VDD VSS edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.signal_w\[0\] sky130_mm_sc_hd_dlyPoly5ns
XFILLER_2_32 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.and_bypass_switch clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.bypass_in clkgen.delay_155ns_3.genblk1\[3\].dly_binary.out
+ VSS VDD VSS VDD sky130_fd_sc_hd__and2b_1
XANTENNA_clkgen.delay_155ns_3.genblk1\[3\].control_invert_A dlycontrol3_in[3] VSS
+ VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.out_mux_A0 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[32\]
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_2_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xclkgen.delay_155ns_2.genblk1\[4\].control_invert dlycontrol2_in[4] clkgen.delay_155ns_2.bypass_enable_w\[4\]
+ VDD VSS VSS VDD sky130_fd_sc_hd__inv_2
Xclkgen.delay_155ns_2.genblk1\[3\].dly_binary.and_bypass_switch clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_2.genblk1\[3\].dly_binary.bypass_in clkgen.delay_155ns_2.genblk1\[2\].dly_binary.out
+ VSS VDD VSS VDD sky130_fd_sc_hd__and2b_1
XFILLER_3_321 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_8_53 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[2\].dly_binary.and_bypass_switch clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_1.genblk1\[2\].dly_binary.bypass_in clkgen.delay_155ns_1.genblk1\[1\].dly_binary.out
+ VSS VDD VSS VDD sky130_fd_sc_hd__and2b_1
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit VSS VDD clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[13\]
+ VDD VSS clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[12\] sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[1\].delay_unit VSS VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[2\]
+ VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[1\] sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_clkgen.delay_155ns_2.genblk1\[0\].dly_binary.and_bypass_switch_A_N clkgen.delay_155ns_2.genblk1\[0\].dly_binary.bypass_in
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_2_205 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit VSS VDD clkgen.delay_155ns_1.genblk1\[1\].dly_binary.signal_w\[2\]
+ VDD VSS clkgen.delay_155ns_1.genblk1\[1\].dly_binary.signal_w\[1\] sky130_mm_sc_hd_dlyPoly5ns
XFILLER_11_315 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.clkdig_inverter_A clkgen.delay_155ns_1.genblk1\[4\].dly_binary.out
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_14_164 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_11_31 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_3_300 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_3_333 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_6_171 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[0\].control_invert dlycontrol4_in[0] edgedetect.dly_315ns_1.bypass_enable_w\[0\]
+ VDD VSS VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_17_85 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_17_30 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[6\].delay_unit VSS VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[7\]
+ VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[6\] sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_1.genblk1\[0\].bypass_enable VDD VSS clkgen.delay_155ns_1.genblk1\[0\].dly_binary.bypass_in
+ clkgen.delay_155ns_1.bypass_enable_w\[0\] clkgen.delay_155ns_1.enable_dlycontrol_w
+ VSS VDD sky130_fd_sc_hd__and2_1
Xedgedetect.dly_315ns_1.genblk1\[0\].dly_binary.genblk1\[0\].delay_unit VSS VDD edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.signal_w\[1\]
+ VDD VSS edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.signal_w\[0\] sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_2.genblk1\[1\].bypass_enable VDD VSS clkgen.delay_155ns_2.genblk1\[1\].dly_binary.bypass_in
+ clkgen.delay_155ns_2.bypass_enable_w\[1\] clkgen.delay_155ns_2.enable_dlycontrol_w
+ VSS VDD sky130_fd_sc_hd__and2_1
XFILLER_12_284 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[2\].bypass_enable VDD VSS clkgen.delay_155ns_3.genblk1\[2\].dly_binary.bypass_in
+ clkgen.delay_155ns_3.bypass_enable_w\[2\] clkgen.delay_155ns_3.enable_dlycontrol_w
+ VSS VDD sky130_fd_sc_hd__and2_1
XFILLER_10_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit VSS VDD clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[5\]
+ VDD VSS clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[4\] sky130_mm_sc_hd_dlyPoly5ns
XFILLER_14_42 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[10\].delay_unit VSS VDD clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[11\]
+ VDD VSS clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[10\] sky130_mm_sc_hd_dlyPoly5ns
XFILLER_5_214 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.delay_155ns_3.genblk1\[3\].bypass_enable_A clkgen.delay_155ns_3.enable_dlycontrol_w
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_4_291 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].control_invert dlycontrol4_in[5] edgedetect.dly_315ns_1.bypass_enable_w\[5\]
+ VDD VSS VSS VDD sky130_fd_sc_hd__inv_2
XPHY_30 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_1_261 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.and_bypass_switch clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.bypass_in clkgen.delay_155ns_2.genblk1\[3\].dly_binary.out
+ VSS VDD VSS VDD sky130_fd_sc_hd__and2b_1
XFILLER_11_327 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.delay_155ns_1.genblk1\[3\].dly_binary.and_bypass_switch_A_N clkgen.delay_155ns_1.genblk1\[3\].dly_binary.bypass_in
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_1.genblk1\[3\].dly_binary.and_bypass_switch clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_1.genblk1\[3\].dly_binary.bypass_in clkgen.delay_155ns_1.genblk1\[2\].dly_binary.out
+ VSS VDD VSS VDD sky130_fd_sc_hd__and2b_1
XANTENNA_sampledly01_A sample_p_in VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit VSS VDD clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[10\]
+ VDD VSS clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[9\] sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit VSS VDD clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[16\]
+ VDD VSS clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[15\] sky130_mm_sc_hd_dlyPoly5ns
XFILLER_0_315 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[0\].control_invert dlycontrol3_in[0] clkgen.delay_155ns_3.bypass_enable_w\[0\]
+ VDD VSS VSS VDD sky130_fd_sc_hd__inv_2
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit VSS VDD edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[2\]
+ VDD VSS edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[1\] sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit VSS VDD clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[4\]
+ VDD VSS clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[3\] sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_edgedetect.dly_315ns_1.genblk1\[2\].control_invert_A dlycontrol4_in[2] VSS
+ VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_12_296 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_12_274 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_8_245 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_8_212 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_14_32 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_17_311 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XPHY_31 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_20 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_1_273 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit VSS VDD edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[7\]
+ VDD VSS edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[6\] sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[1\].dly_binary.out_mux VSS VDD edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.bypass_in
+ edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.out edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.signal_w\[2\]
+ edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.out VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_11_339 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_11_306 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit VSS VDD clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[9\]
+ VDD VSS clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[8\] sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[3\].dly_binary.out_mux VSS VDD edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.bypass_in
+ edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.out edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[8\]
+ edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.out VSS VDD sky130_fd_sc_hd__mux2_1
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.out_mux VSS VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.bypass_in
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.out edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[32\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.out VSS VDD sky130_fd_sc_hd__mux2_1
Xclkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit VSS VDD clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[5\]
+ VDD VSS clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[4\] sky130_mm_sc_hd_dlyPoly5ns
XFILLER_11_125 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_inbuf_2_A start_conv_in VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_6_151 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[2\].delay_unit VSS VDD clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[3\]
+ VDD VSS clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[2\] sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_clkgen.delay_155ns_1.genblk1\[3\].dly_binary.out_mux_A1 clkgen.delay_155ns_1.genblk1\[2\].dly_binary.out
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_3_187 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA_clkgen.delay_155ns_1.genblk1\[3\].dly_binary.out_mux_S clkgen.delay_155ns_1.genblk1\[3\].dly_binary.bypass_in
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[13\].delay_unit VSS VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[14\]
+ VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[13\] sky130_mm_sc_hd_dlyPoly5ns
XFILLER_12_253 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit VSS VDD clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[14\]
+ VDD VSS clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[13\] sky130_mm_sc_hd_dlyPoly5ns
XFILLER_14_55 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_5_249 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XPHY_32 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_21 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.and_bypass_switch clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.bypass_in clkgen.delay_155ns_1.genblk1\[3\].dly_binary.out
+ VSS VDD VSS VDD sky130_fd_sc_hd__and2b_1
XPHY_10 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit VSS VDD edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[15\]
+ VDD VSS edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[14\] sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.and_bypass_switch_A_N edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.bypass_in
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_1_285 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_1_230 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit VSS VDD edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[2\]
+ VDD VSS edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[1\] sky130_mm_sc_hd_dlyPoly5ns
Xoutbuf_1 VDD VSS clk_dig_out clkgen.clk_dig_out VSS VDD sky130_fd_sc_hd__buf_4
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit VSS VDD clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[8\]
+ VDD VSS clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[7\] sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_edgedetect.dly_315ns_1.genblk1\[4\].bypass_enable_A edgedetect.dly_315ns_1.enable_dlycontrol_w
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit VSS VDD clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[4\]
+ VDD VSS clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[3\] sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[18\].delay_unit VSS VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[19\]
+ VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[18\] sky130_mm_sc_hd_dlyPoly5ns
XFILLER_18_292 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA_clkgen.delay_155ns_1.genblk1\[4\].control_invert_A dlycontrol1_in[4] VSS
+ VDD VDD VSS sky130_fd_sc_hd__diode_2
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[20\].delay_unit VSS VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[21\]
+ VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[20\] sky130_mm_sc_hd_dlyPoly5ns
XFILLER_0_306 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[1\].control_invert dlycontrol1_in[1] clkgen.delay_155ns_1.bypass_enable_w\[1\]
+ VDD VSS VSS VDD sky130_fd_sc_hd__inv_2
Xclkgen.delay_155ns_1.genblk1\[1\].dly_binary.out_mux VSS VDD clkgen.delay_155ns_1.genblk1\[1\].dly_binary.bypass_in
+ clkgen.delay_155ns_1.genblk1\[0\].dly_binary.out clkgen.delay_155ns_1.genblk1\[1\].dly_binary.signal_w\[2\]
+ clkgen.delay_155ns_1.genblk1\[1\].dly_binary.out VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_8_203 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_0_125 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xedgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit VSS VDD edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[7\]
+ VDD VSS edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[6\] sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_1.genblk1\[3\].dly_binary.out_mux VSS VDD clkgen.delay_155ns_1.genblk1\[3\].dly_binary.bypass_in
+ clkgen.delay_155ns_1.genblk1\[2\].dly_binary.out clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[8\]
+ clkgen.delay_155ns_1.genblk1\[3\].dly_binary.out VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_17_302 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.delay_155ns_2.genblk1\[3\].control_invert_A dlycontrol2_in[3] VSS
+ VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_clkgen.delay_155ns_1.genblk1\[1\].dly_binary.out_mux_S clkgen.delay_155ns_1.genblk1\[1\].dly_binary.bypass_in
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XPHY_33 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_22 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_17_121 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_1_297 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[25\].delay_unit VSS VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[26\]
+ VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[25\] sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit VSS VDD clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[3\]
+ VDD VSS clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[2\] sky130_mm_sc_hd_dlyPoly5ns
Xoutbuf_2 VDD VSS clk_comp_out clkgen.clk_comp_out VSS VDD sky130_fd_sc_hd__buf_4
XFILLER_14_124 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_9_183 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA_clkgen.delay_155ns_3.genblk1\[2\].control_invert_A dlycontrol3_in[2] VSS
+ VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_3_315 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_19_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_6_164 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_3_178 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[2\].dly_binary.genblk1\[1\].delay_unit VSS VDD edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[2\]
+ VDD VSS edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[1\] sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit VSS VDD clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[8\]
+ VDD VSS clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[7\] sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_2.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit VSS VDD clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[4\]
+ VDD VSS clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[3\] sky130_mm_sc_hd_dlyPoly5ns
XPHY_12 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_17_155 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_34 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_23 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_1_254 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_2_16 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xoutbuf_3 VDD VSS sample_p_out sample_p_4 VSS VDD sky130_fd_sc_hd__buf_4
Xclkgen.delay_155ns_3.genblk1\[0\].dly_binary.out_mux VSS VDD clkgen.delay_155ns_3.genblk1\[0\].dly_binary.bypass_in
+ clkgen.delay_155ns_3.genblk1\[0\].dly_binary.in clkgen.delay_155ns_3.genblk1\[0\].dly_binary.signal_w\[1\]
+ clkgen.delay_155ns_3.genblk1\[0\].dly_binary.out VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_13_180 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xclkgen.delay_155ns_3.genblk1\[2\].dly_binary.out_mux VSS VDD clkgen.delay_155ns_3.genblk1\[2\].dly_binary.bypass_in
+ clkgen.delay_155ns_3.genblk1\[1\].dly_binary.out clkgen.delay_155ns_3.genblk1\[2\].dly_binary.signal_w\[4\]
+ clkgen.delay_155ns_3.genblk1\[2\].dly_binary.out VSS VDD sky130_fd_sc_hd__mux2_1
XANTENNA_outbuf_1_A clkgen.clk_dig_out VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xedgedetect.dly_315ns_1.genblk1\[5\].bypass_enable VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.bypass_in
+ edgedetect.dly_315ns_1.bypass_enable_w\[5\] edgedetect.dly_315ns_1.enable_dlycontrol_w
+ VSS VDD sky130_fd_sc_hd__and2_1
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.out_mux VSS VDD clkgen.delay_155ns_3.genblk1\[4\].dly_binary.bypass_in
+ clkgen.delay_155ns_3.genblk1\[3\].dly_binary.out clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[16\]
+ clkgen.clk_comp_out VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_16_209 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_12_267 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit VSS VDD clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[3\]
+ VDD VSS clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[2\] sky130_mm_sc_hd_dlyPoly5ns
XFILLER_4_274 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_4_285 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_35 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_24 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_13 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_1_244 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xoutbuf_4 VDD VSS sample_n_out sample_n_4 VSS VDD sky130_fd_sc_hd__buf_4
Xclkgen.delay_155ns_3.enablebuffer VDD VSS clkgen.delay_155ns_3.enable_dlycontrol_w
+ enable_dlycontrol_in VSS VDD sky130_fd_sc_hd__buf_4
XFILLER_6_336 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_3_71 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xclkgen.delay_155ns_2.genblk1\[2\].control_invert dlycontrol2_in[2] clkgen.delay_155ns_2.bypass_enable_w\[2\]
+ VDD VSS VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_19_218 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xedgedetect.dly_315ns_1.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit VSS VDD edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.signal_w\[2\]
+ VDD VSS edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.signal_w\[1\] sky130_mm_sc_hd_dlyPoly5ns
XFILLER_8_16 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_3_306 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.delay_155ns_2.genblk1\[4\].dly_binary.out_mux_A0 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[16\]
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_3_147 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_15_276 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_0_94 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_12_246 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_edgedetect.dly_315ns_1.genblk1\[1\].control_invert_A dlycontrol4_in[1] VSS
+ VDD VDD VSS sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit VSS VDD clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[14\]
+ VDD VSS clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[13\] sky130_mm_sc_hd_dlyPoly5ns
XFILLER_4_297 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_36 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_25 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_1_267 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_1_223 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_14 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xedgedetect.dly_315ns_1.genblk1\[0\].bypass_enable VDD VSS edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.bypass_in
+ edgedetect.dly_315ns_1.bypass_enable_w\[0\] edgedetect.dly_315ns_1.enable_dlycontrol_w
+ VSS VDD sky130_fd_sc_hd__and2_1
Xoutbuf_5 VDD VSS nsample_p_out nsample_p_4 VSS VDD sky130_fd_sc_hd__buf_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[2\].delay_unit VSS VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[3\]
+ VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[2\] sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.out_mux_S edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.bypass_in
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_10_322 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_13_171 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_18_274 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_10_174 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[0\].delay_unit VSS VDD clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[1\]
+ VDD VSS clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[0\] sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_1.genblk1\[1\].bypass_enable VDD VSS clkgen.delay_155ns_1.genblk1\[1\].dly_binary.bypass_in
+ clkgen.delay_155ns_1.bypass_enable_w\[1\] clkgen.delay_155ns_1.enable_dlycontrol_w
+ VSS VDD sky130_fd_sc_hd__and2_1
XFILLER_17_59 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xclkgen.delay_155ns_2.genblk1\[2\].bypass_enable VDD VSS clkgen.delay_155ns_2.genblk1\[2\].dly_binary.bypass_in
+ clkgen.delay_155ns_2.bypass_enable_w\[2\] clkgen.delay_155ns_2.enable_dlycontrol_w
+ VSS VDD sky130_fd_sc_hd__and2_1
XFILLER_3_137 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.delay_155ns_2.genblk1\[1\].dly_binary.out_mux_S clkgen.delay_155ns_2.genblk1\[1\].dly_binary.bypass_in
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_3.genblk1\[3\].bypass_enable VDD VSS clkgen.delay_155ns_3.genblk1\[3\].dly_binary.bypass_in
+ clkgen.delay_155ns_3.bypass_enable_w\[3\] clkgen.delay_155ns_3.enable_dlycontrol_w
+ VSS VDD sky130_fd_sc_hd__and2_1
XFILLER_9_93 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[7\].delay_unit VSS VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[8\]
+ VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[7\] sky130_mm_sc_hd_dlyPoly5ns
XFILLER_14_16 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[3\].control_invert dlycontrol4_in[3] edgedetect.dly_315ns_1.bypass_enable_w\[3\]
+ VDD VSS VSS VDD sky130_fd_sc_hd__inv_2
XPHY_37 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_26 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_15 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_17_125 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_17_114 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit VSS VDD clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[6\]
+ VDD VSS clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[5\] sky130_mm_sc_hd_dlyPoly5ns
XFILLER_1_279 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_16_180 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit VSS VDD clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[12\]
+ VDD VSS clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[11\] sky130_mm_sc_hd_dlyPoly5ns
Xoutbuf_6 VDD VSS nsample_n_out nsample_n_4 VSS VDD sky130_fd_sc_hd__buf_4
XFILLER_9_176 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_10_164 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.out_mux_S edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.bypass_in
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_clkgen.delay_155ns_1.genblk1\[3\].control_invert_A dlycontrol1_in[3] VSS
+ VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_3_116 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_0_63 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA_clkgen.delay_155ns_1.genblk1\[1\].dly_binary.and_bypass_switch_A_N clkgen.delay_155ns_1.genblk1\[1\].dly_binary.bypass_in
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_clkgen.delay_155ns_2.genblk1\[0\].dly_binary.out_mux_A1 clkgen.clk_dig_out
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[2\].delay_unit VSS VDD edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[3\]
+ VDD VSS edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[2\] sky130_mm_sc_hd_dlyPoly5ns
XPHY_38 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_27 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit VSS VDD clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[5\]
+ VDD VSS clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[4\] sky130_mm_sc_hd_dlyPoly5ns
XPHY_16 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA_clkgen.delay_155ns_2.genblk1\[2\].control_invert_A dlycontrol2_in[2] VSS
+ VDD VDD VSS sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_3.genblk1\[3\].control_invert dlycontrol3_in[3] clkgen.delay_155ns_3.bypass_enable_w\[3\]
+ VDD VSS VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_15_93 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[0\].delay_unit VSS VDD clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[1\]
+ VDD VSS clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[0\] sky130_mm_sc_hd_dlyPoly5ns
XFILLER_1_214 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.delay_155ns_3.enablebuffer_A enable_dlycontrol_in VSS VDD VDD VSS
+ sky130_fd_sc_hd__diode_2
XANTENNA_clkgen.delay_155ns_3.genblk1\[1\].control_invert_A dlycontrol3_in[1] VSS
+ VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_clkgen.delay_155ns_3.genblk1\[1\].bypass_enable_A clkgen.delay_155ns_3.enable_dlycontrol_w
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_12_94 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_10_121 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_2_320 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit VSS VDD edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[8\]
+ VDD VSS edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[7\] sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit VSS VDD clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[10\]
+ VDD VSS clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[9\] sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.out_mux_S edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.bypass_in
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit VSS VDD clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[6\]
+ VDD VSS clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[5\] sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[10\].delay_unit VSS VDD edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[11\]
+ VDD VSS edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[10\] sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.and_bypass_switch_A_N edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.bypass_in
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_11_282 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.delay_155ns_1.genblk1\[3\].dly_binary.and_bypass_switch_B clkgen.delay_155ns_1.genblk1\[2\].dly_binary.out
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit VSS VDD clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[4\]
+ VDD VSS clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[3\] sky130_mm_sc_hd_dlyPoly5ns
XFILLER_4_245 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_28 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_17 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_39 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_13_300 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_1_237 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[14\].delay_unit VSS VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[15\]
+ VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[14\] sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit VSS VDD clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[15\]
+ VDD VSS clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[14\] sky130_mm_sc_hd_dlyPoly5ns
XFILLER_0_292 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_6_307 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit VSS VDD edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[16\]
+ VDD VSS edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[15\] sky130_mm_sc_hd_dlyPoly5ns
XFILLER_2_332 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xedgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit VSS VDD edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[3\]
+ VDD VSS edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[2\] sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit VSS VDD clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[9\]
+ VDD VSS clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[8\] sky130_mm_sc_hd_dlyPoly5ns
XFILLER_15_214 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_9_30 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.and_bypass_switch_A_N edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.bypass_in
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_0_32 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_2_195 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit VSS VDD clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[5\]
+ VDD VSS clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[4\] sky130_mm_sc_hd_dlyPoly5ns
XFILLER_14_280 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[2\].dly_binary.genblk1\[0\].delay_unit VSS VDD clkgen.delay_155ns_3.genblk1\[2\].dly_binary.signal_w\[1\]
+ VDD VSS clkgen.delay_155ns_3.genblk1\[2\].dly_binary.signal_w\[0\] sky130_mm_sc_hd_dlyPoly5ns
XFILLER_9_63 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_18_94 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[19\].delay_unit VSS VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[20\]
+ VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[19\] sky130_mm_sc_hd_dlyPoly5ns
XFILLER_11_294 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[21\].delay_unit VSS VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[22\]
+ VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[21\] sky130_mm_sc_hd_dlyPoly5ns
XFILLER_15_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_7_276 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_18 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xedgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit VSS VDD edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[8\]
+ VDD VSS edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[7\] sky130_mm_sc_hd_dlyPoly5ns
XFILLER_9_338 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_9_305 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[4\].control_invert dlycontrol1_in[4] clkgen.delay_155ns_1.bypass_enable_w\[4\]
+ VDD VSS VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_13_142 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_9_146 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_3_87 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_6_138 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_6_105 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_18_245 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[26\].delay_unit VSS VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[27\]
+ VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[26\] sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit VSS VDD clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[4\]
+ VDD VSS clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[3\] sky130_mm_sc_hd_dlyPoly5ns
XFILLER_18_62 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_12_218 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA_edgedetect.dly_315ns_1.genblk1\[2\].bypass_enable_A edgedetect.dly_315ns_1.enable_dlycontrol_w
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_edgedetect.dly_315ns_1.genblk1\[0\].control_invert_A dlycontrol4_in[0] VSS
+ VDD VDD VSS sky130_fd_sc_hd__diode_2
XPHY_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xedgedetect.dly_315ns_1.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit VSS VDD edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[3\]
+ VDD VSS edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[2\] sky130_mm_sc_hd_dlyPoly5ns
XFILLER_15_63 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_0_261 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_16_173 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[1\].dly_binary.genblk1\[0\].delay_unit VSS VDD clkgen.delay_155ns_3.genblk1\[1\].dly_binary.signal_w\[1\]
+ VDD VSS clkgen.delay_155ns_3.genblk1\[1\].dly_binary.signal_w\[0\] sky130_mm_sc_hd_dlyPoly5ns
XFILLER_9_125 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_5_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_2_164 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_7_245 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_6_88 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_15_31 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit VSS VDD clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[4\]
+ VDD VSS clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[3\] sky130_mm_sc_hd_dlyPoly5ns
.ends

.subckt sky130_fd_sc_hd__a21bo_2 B1_N A2 X A1 VGND VPWR VNB VPB
X0 VPWR A1 a_485_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=8.93e+11p pd=8.08e+06u as=5.3e+11p ps=5.06e+06u w=1e+06u l=150000u
X1 a_485_297# a_297_93# a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X2 a_297_93# B1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=7.2375e+11p ps=7.48e+06u w=420000u l=150000u
X3 a_581_47# A1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.72e+06u as=2.145e+11p ps=1.96e+06u w=650000u l=150000u
X4 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X5 a_79_21# a_297_93# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND A2 a_581_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X8 a_297_93# B1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X9 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_485_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a2111o_1 VGND VPWR B1 X D1 A1 A2 C1 VNB VPB
X0 VGND A2 a_660_47# VNB sky130_fd_pr__nfet_01v8 ad=9.7175e+11p pd=6.89e+06u as=1.6575e+11p ps=1.81e+06u w=650000u l=150000u
X1 VGND C1 a_85_193# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.72e+11p ps=4.36e+06u w=650000u l=150000u
X2 a_414_297# C1 a_334_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=3.6e+11p pd=2.72e+06u as=2.5e+11p ps=2.5e+06u w=1e+06u l=150000u
X3 VGND a_85_193# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.145e+11p ps=1.96e+06u w=650000u l=150000u
X4 a_334_297# D1 a_85_193# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.85e+11p ps=2.77e+06u w=1e+06u l=150000u
X5 a_516_297# B1 a_414_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=8.5e+11p pd=5.7e+06u as=0p ps=0u w=1e+06u l=150000u
X6 a_516_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.35e+11p ps=5.07e+06u w=1e+06u l=150000u
X7 a_660_47# A1 a_85_193# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_85_193# D1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR A1 a_516_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_85_193# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR a_85_193# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__dfstp_1 D VPWR Q SET_B CLK VGND VNB VPB
X0 VGND a_652_21# a_586_47# VNB sky130_fd_pr__nfet_01v8 ad=9.868e+11p pd=1.019e+07u as=1.341e+11p ps=1.5e+06u w=420000u l=150000u
X1 a_956_413# a_476_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=9.66e+10p pd=1.3e+06u as=1.3171e+12p ps=1.335e+07u w=420000u l=150000u
X2 VPWR a_476_47# a_652_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X3 a_586_47# a_193_47# a_476_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.44e+11p ps=1.52e+06u w=360000u l=150000u
X4 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X5 a_476_47# a_27_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.87e+11p ps=1.93e+06u w=360000u l=150000u
X6 a_1056_47# a_476_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X7 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.499e+11p pd=2.35e+06u as=0p ps=0u w=840000u l=150000u
X8 a_652_21# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_1224_47# a_27_47# a_1032_413# VNB sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X10 a_562_413# a_27_47# a_476_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=1.89e+11p pd=1.74e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X11 VGND a_1032_413# a_1602_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X12 VPWR a_1182_261# a_1140_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X13 Q a_1602_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X14 a_1032_413# a_193_47# a_1056_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_476_47# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 a_1296_47# a_1182_261# a_1224_47# VNB sky130_fd_pr__nfet_01v8 ad=9.66e+10p pd=1.3e+06u as=0p ps=0u w=420000u l=150000u
X17 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X18 VPWR a_652_21# a_562_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 VPWR SET_B a_1032_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.73e+11p ps=2.98e+06u w=420000u l=150000u
X20 a_1032_413# a_27_47# a_956_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 a_1182_261# a_1032_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.184e+11p pd=2.2e+06u as=0p ps=0u w=840000u l=150000u
X22 Q a_1602_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X23 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X24 a_1140_413# a_193_47# a_1032_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 VPWR a_1032_413# a_1602_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X26 a_796_47# SET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X27 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X28 a_1182_261# a_1032_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.404e+11p pd=1.6e+06u as=0p ps=0u w=540000u l=150000u
X29 a_652_21# a_476_47# a_796_47# VNB sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X30 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X31 VGND SET_B a_1296_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a2111oi_1 B1 D1 C1 Y A2 A1 VPWR VGND VNB VPB
X0 a_316_297# C1 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=3.7e+11p pd=2.74e+06u as=3.45e+11p ps=2.69e+06u w=1e+06u l=150000u
X1 Y D1 VGND VNB sky130_fd_pr__nfet_01v8 ad=6.3375e+11p pd=4.55e+06u as=9.1325e+11p ps=6.71e+06u w=650000u l=150000u
X2 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_420_297# B1 a_316_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=8.7e+11p pd=5.74e+06u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR A1 a_420_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=2.75e+11p pd=2.55e+06u as=0p ps=0u w=1e+06u l=150000u
X5 VGND A2 a_568_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X6 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_420_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_217_297# D1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=7.55e+11p ps=3.51e+06u w=1e+06u l=150000u
X9 a_568_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 X VGND VPWR VNB VPB
X0 VGND A4 a_321_47# VNB sky130_fd_pr__nfet_01v8 ad=6.695e+11p pd=5.96e+06u as=6.24e+11p ps=5.82e+06u w=650000u l=150000u
X1 a_321_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_103_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=5.2e+11p pd=3.04e+06u as=5.5e+11p ps=5.1e+06u w=1e+06u l=150000u
X3 VPWR a_103_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.25e+11p ps=2.85e+06u w=1e+06u l=150000u
X4 VGND a_103_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.47e+11p ps=2.06e+06u w=650000u l=150000u
X5 VGND A2 a_321_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_321_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_511_297# A3 a_393_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=3.9e+11p pd=2.78e+06u as=4.4e+11p ps=2.88e+06u w=1e+06u l=150000u
X8 a_619_297# A2 a_511_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=3.9e+11p pd=2.78e+06u as=0p ps=0u w=1e+06u l=150000u
X9 a_321_47# B1 a_103_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X10 a_393_297# A4 a_103_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VPWR A1 a_619_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__dfstp_4 Q D VPWR SET_B CLK VGND VNB VPB
X0 a_1178_261# a_1028_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.184e+11p pd=2.2e+06u as=1.8571e+12p ps=1.843e+07u w=840000u l=150000u
X1 VGND a_652_21# a_586_47# VNB sky130_fd_pr__nfet_01v8 ad=1.3378e+12p pd=1.387e+07u as=1.341e+11p ps=1.5e+06u w=420000u l=150000u
X2 VPWR a_1028_413# a_1598_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X3 a_1178_261# a_1028_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.404e+11p pd=1.6e+06u as=0p ps=0u w=540000u l=150000u
X4 VGND a_1598_47# Q VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.2e+11p ps=5.5e+06u w=650000u l=150000u
X5 a_956_413# a_476_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X6 a_1136_413# a_193_47# a_1028_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=2.73e+11p ps=2.98e+06u w=420000u l=150000u
X7 VPWR a_1598_47# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8e+11p ps=7.6e+06u w=1e+06u l=150000u
X8 VPWR a_476_47# a_652_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X9 a_586_47# a_193_47# a_476_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.44e+11p ps=1.52e+06u w=360000u l=150000u
X10 VGND a_1598_47# Q VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X12 Q a_1598_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_476_47# a_27_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.87e+11p ps=1.93e+06u w=360000u l=150000u
X14 a_1056_47# a_476_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X15 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.499e+11p pd=2.35e+06u as=0p ps=0u w=840000u l=150000u
X16 a_652_21# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 a_1224_47# a_27_47# a_1028_413# VNB sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X18 a_562_413# a_27_47# a_476_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=1.89e+11p pd=1.74e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X19 a_1028_413# a_193_47# a_1056_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 a_476_47# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 Q a_1598_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_1296_47# a_1178_261# a_1224_47# VNB sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X23 VGND a_1028_413# a_1598_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X24 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X25 VPWR a_652_21# a_562_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 VPWR a_1598_47# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 VGND SET_B a_1296_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 Q a_1598_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 a_1028_413# a_27_47# a_956_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X30 VPWR a_1178_261# a_1136_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X31 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X32 Q a_1598_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X33 a_796_47# SET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X34 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X35 Q a_1598_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X36 Q a_1598_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X37 a_652_21# a_476_47# a_796_47# VNB sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X38 VPWR SET_B a_1028_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X39 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nor3b_4 A C_N B Y VGND VPWR VNB VPB
X0 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=1.053e+12p pd=1.104e+07u as=1.56e+12p ps=1.39e+07u w=650000u l=150000u
X1 VPWR A a_197_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=8e+11p pd=7.6e+06u as=1.08e+12p ps=1.016e+07u w=1e+06u l=150000u
X2 Y a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_555_297# a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=1.33e+12p pd=1.266e+07u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X5 a_197_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND a_27_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_197_297# B a_555_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND a_27_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND C_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X12 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 Y a_27_47# a_555_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 Y a_27_47# a_555_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VPWR C_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X16 a_555_297# a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 a_555_297# B a_197_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 a_197_297# B a_555_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 a_555_297# B a_197_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 VPWR A a_197_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 a_197_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 Y a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 Y VGND VPWR VNB VPB
X0 a_27_47# C1 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=8.645e+11p pd=9.16e+06u as=7.02e+11p ps=7.36e+06u w=650000u l=150000u
X1 a_803_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=1.27725e+12p pd=1.303e+07u as=7.02e+11p ps=7.36e+06u w=650000u l=150000u
X2 a_27_47# C1 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VGND A2 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_1163_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=1.08e+12p pd=1.016e+07u as=2.63335e+12p ps=2.328e+07u w=1e+06u l=150000u
X5 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=2.40285e+12p pd=2.282e+07u as=0p ps=0u w=1e+06u l=150000u
X6 VGND A2 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Y D1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 Y A2 a_1163_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_1163_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_445_47# B1 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR D1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_445_47# B1 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 Y D1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VPWR A1 a_1163_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_27_47# D1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u
X16 a_27_47# D1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 VGND A1 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 a_1163_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 a_803_47# B1 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 VPWR A1 a_1163_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 a_803_47# B1 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 Y D1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X27 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 a_445_47# C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X29 a_803_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X30 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 a_1163_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 Y A2 a_1163_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X33 a_445_47# C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X34 a_803_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X35 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X36 a_803_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X37 VPWR D1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X38 Y D1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X39 VGND A1 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt adc_top VDD VSS clk_vcm config_1_in[0] config_1_in[10] config_1_in[11] config_1_in[12]
+ config_1_in[13] config_1_in[14] config_1_in[15] config_1_in[1] config_1_in[2] config_1_in[3]
+ config_1_in[4] config_1_in[5] config_1_in[6] config_1_in[7] config_1_in[8] config_1_in[9]
+ config_2_in[0] config_2_in[10] config_2_in[11] config_2_in[12] config_2_in[13] config_2_in[14]
+ config_2_in[15] config_2_in[1] config_2_in[2] config_2_in[3] config_2_in[4] config_2_in[5]
+ config_2_in[6] config_2_in[7] config_2_in[8] config_2_in[9] conversion_finished_out
+ dummypin[0] dummypin[10] dummypin[11] dummypin[12] dummypin[13] dummypin[14] dummypin[15]
+ dummypin[1] dummypin[2] dummypin[3] dummypin[4] dummypin[5] dummypin[6] dummypin[7]
+ dummypin[8] dummypin[9] inn_analog inp_analog result_out[0] result_out[10] result_out[11]
+ result_out[12] result_out[13] result_out[14] result_out[15] result_out[1] result_out[2]
+ result_out[3] result_out[4] result_out[5] result_out[6] result_out[7] result_out[8]
+ result_out[9] rst_n start_conversion_in
XANTENNA__1725__RESET_B net63 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_50_431 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_139_9 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA_fanout75_A net76 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_26_85 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1445__A1 _0529_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_pmat_col_n[7] core.pdc.col_out_n\[7\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_42_95 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_47_8 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1270_ VSS VDD _0633_ _0631_ core.cnb.average_sum_r\[3\] _0629_ VSS VDD sky130_fd_sc_hd__and3_1
XFILLER_67_81 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_91_375 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_0985_ VDD VSS _0411_ _0365_ core.cnb.data_register_r\[2\] VSS VDD sky130_fd_sc_hd__and2_1
X_1606_ _0234_ _0133_ _0736_ _0221_ VSS VDD VSS VDD sky130_fd_sc_hd__nor3_1
X_1537_ core.pdc.row_out_n\[13\] _0077_ core.ndc.row_out_n\[4\] VSS VDD VSS VDD sky130_fd_sc_hd__nand2_1
X_1468_ _0353_ _0500_ _0463_ _0499_ _0052_ VSS VDD VSS VDD sky130_fd_sc_hd__o211a_1
X_1399_ VSS VDD core.osr.next_result_w\[16\] _0744_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XANTENNA__1747__CLK net81 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_103_57 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_63_28 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_82_375 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_6_129 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_137_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_12_65 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1264__A _0616_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_92_117 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_128_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1322_ VSS VDD _0677_ _0653_ _0651_ _0676_ VSS VDD sky130_fd_sc_hd__and3_1
X_1253_ core.cnb.average_counter_r\[4\] _0621_ VDD VSS VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_83_117 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1184_ _0566_ core.cnb.average_counter_r\[4\] _0568_ _0567_ VSS VDD VSS VDD sky130_fd_sc_hd__a21o_4
XFILLER_80_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_0968_ _0394_ _0393_ core.cnb.data_register_r\[7\] VSS VDD VSS VDD sky130_fd_sc_hd__xnor2_4
XFILLER_119_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_0899_ _0325_ _0318_ core.cnb.data_register_r\[5\] _0322_ _0324_ VSS VDD VSS VDD
+ sky130_fd_sc_hd__a211o_2
XFILLER_58_17 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1531__B core.ndc.row_out_n\[12\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1112__A3 _0468_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_55_386 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_71_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_135_3 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1259__A core.cnb.comparator_in VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_139_53 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_139_97 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_99_35 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1584__B1 core.osr.next_result_w\[5\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_99_57 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1639__A1 core.cnb.result_out\[5\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_0_57 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_62_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_0822_ VSS VDD core.cnb.shift_register_r\[7\] _0248_ core.cnb.shift_register_r\[5\]
+ VSS VDD sky130_fd_sc_hd__xnor2_1
XFILLER_89_90 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1335__C _0634_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_84_404 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1305_ _0661_ _0662_ core.osr.result_r\[5\] VDD VSS VSS VDD sky130_fd_sc_hd__xor2_1
X_1236_ VSS VDD _0609_ _0610_ core.cnb.data_register_r\[10\] VSS VDD sky130_fd_sc_hd__xnor2_1
X_1167_ _0553_ _0552_ _0255_ _0254_ _0554_ VSS VDD VSS VDD sky130_fd_sc_hd__nor4b_1
XANTENNA__1351__B core.cnb.result_out\[8\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1098_ _0513_ _0474_ _0470_ VSS VDD VSS VDD sky130_fd_sc_hd__nand2_2
XFILLER_53_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_100_25 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_60_29 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1079__A _0394_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xadc_top_94 dummypin[9] adc_top_94/HI VDD VSS VSS VDD sky130_fd_sc_hd__conb_1
XFILLER_87_242 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_18_20 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_18_97 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_510 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1688__S _0616_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_44_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XPHY_543 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_532 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_521 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_554 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1557__A0 core.cnb.result_out\[5\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1021__A2 _0427_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1021_ _0426_ _0427_ _0446_ _0441_ _0445_ _0430_ VSS VDD VSS VDD sky130_fd_sc_hd__a311o_1
XFILLER_35_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_98_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_0805_ _0213_ _0232_ _0214_ VSS VDD VSS VDD sky130_fd_sc_hd__nand2b_2
X_1785_ core.osr.result_r\[17\] net71 core.osr.next_result_w\[17\] net59 VSS VDD VSS
+ VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_55_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_1219_ VDD VSS _0596_ _0595_ net53 VSS VDD sky130_fd_sc_hd__and2_1
XFILLER_26_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_111_57 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_52_197 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1537__A core.ndc.row_out_n\[4\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_136_65 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_96_25 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_96_47 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_29_74 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA_input18_A config_2_in[10] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_45_51 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_45_62 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_17_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_90_248 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_340 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_351 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_362 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_373 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_384 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_395 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_77_8 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_1570_ _0101_ _0102_ _0588_ VSS VDD VSS VDD sky130_fd_sc_hd__nor2_1
X_1004_ _0429_ _0428_ _0361_ VSS VDD VSS VDD sky130_fd_sc_hd__nand2_1
XANTENNA__1233__A2 _0579_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__0992__A1 _0364_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1357__A _0709_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1768_ core.osr.result_r\[0\] net65 core.osr.next_result_w\[0\] net55 VSS VDD VSS
+ VDD sky130_fd_sc_hd__dfrtp_1
X_1699_ VSS VDD _0043_ _0201_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_106_35 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_66_39 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_122_56 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_25_120 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_53_484 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1267__A _0616_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xoutput42 VDD VSS result_out[15] net42 VSS VDD sky130_fd_sc_hd__buf_2
XPHY_170 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_181 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_192 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_1622_ _0132_ net48 _0147_ _0134_ VSS VDD VSS VDD sky130_fd_sc_hd__or3b_1
X_1553_ VSS VDD _0089_ core.cnb.next_data_register_w\[3\] core.cnb.result_out\[3\]
+ _0093_ VSS VDD sky130_fd_sc_hd__mux2_1
X_1484_ _0058_ _0598_ core.cnb.data_register_r\[10\] VSS VDD VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_54_204 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_50_421 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1087__A _0466_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_7_8 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_77_27 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_fanout68_A net69 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_85_384 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_53_281 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1696__S _0614_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_9_105 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA_pmat_col_n[6] core.pdc.col_out_n\[6\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_42_63 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_6_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_3_57 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1133__A1 _0353_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_80_3 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_0984_ _0410_ _0409_ _0396_ VSS VDD VSS VDD sky130_fd_sc_hd__xnor2_4
X_1605_ VDD VSS _0132_ _0209_ VSS VDD sky130_fd_sc_hd__buf_2
X_1536_ core.pdc.row_out_n\[12\] core.ndc.row_out_n\[4\] VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_2
X_1467_ _0531_ core.ndc.col_out_n\[23\] _0526_ VSS VDD VSS VDD sky130_fd_sc_hd__nor2_1
XFILLER_86_126 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1398_ VSS VDD _0744_ _0742_ _0635_ _0743_ VSS VDD sky130_fd_sc_hd__and3_1
XFILLER_82_343 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_82_365 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_82_398 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_137_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_128_22 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_12_77 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1545__A core.cnb.shift_register_r\[2\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1363__B2 core.cnb.result_out\[9\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_53_84 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_53_95 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_128_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1321_ _0665_ core.osr.result_r\[7\] core.osr.result_r\[6\] _0676_ _0669_ VDD VSS
+ VSS VDD sky130_fd_sc_hd__a211oi_1
X_1252_ _0620_ core.cnb.next_average_counter_w\[3\] _0616_ VSS VDD VSS VDD sky130_fd_sc_hd__nor2_1
XFILLER_83_129 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1183_ _0567_ core.cnb.average_counter_r\[4\] _0562_ _0566_ VSS VDD VSS VDD sky130_fd_sc_hd__o21a_1
X_0967_ _0393_ _0392_ _0391_ _0388_ _0381_ _0373_ VDD VSS VSS VDD sky130_fd_sc_hd__o2111a_1
XANTENNA__1188__A4 core.cnb.comparator_in VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_119_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_0898_ _0258_ _0324_ _0323_ _0264_ VSS VDD VSS VDD sky130_fd_sc_hd__nor3_1
XFILLER_58_29 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1519_ core.ndc.row_out_n\[10\] core.pdc.row_out_n\[6\] VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_2
XANTENNA__1780__RESET_B net67 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_55_398 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_139_21 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_23_32 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_23_65 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1584__A1 _0110_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_0_69 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_64_72 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_80_60 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_0821_ _0245_ _0244_ _0247_ _0242_ _0246_ VDD VSS VSS VDD sky130_fd_sc_hd__or4_1
XANTENNA__1737__CLK net76 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1304_ _0661_ core.osr.result_r\[4\] _0660_ _0654_ VSS VDD VSS VDD sky130_fd_sc_hd__a21bo_1
X_1235_ _0541_ _0609_ _0554_ _0586_ core.cnb.data_register_r\[9\] _0605_ VSS VDD VSS
+ VDD sky130_fd_sc_hd__o221a_1
X_1166_ _0252_ _0553_ core.cnb.shift_register_r\[12\] _0264_ VDD VSS VSS VDD sky130_fd_sc_hd__or3_1
X_1097_ _0472_ _0512_ _0462_ VSS VDD VSS VDD sky130_fd_sc_hd__nor2_2
XFILLER_100_59 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xadc_top_95 dummypin[10] adc_top_95/HI VDD VSS VSS VDD sky130_fd_sc_hd__conb_1
XANTENNA__1095__A _0466_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_109_57 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_87_221 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_85_16 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_125_89 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XPHY_500 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_544 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_533 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_522 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_511 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_555 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_59_72 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_46_151 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_1020_ _0429_ _0444_ _0425_ _0443_ _0445_ VSS VDD VSS VDD sky130_fd_sc_hd__a31o_1
XFILLER_75_71 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_75_82 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_0804_ _0231_ _0230_ core.osr.sample_count_r\[6\] VSS VDD VSS VDD sky130_fd_sc_hd__nand2_1
XANTENNA__0812__A core.cnb.shift_register_r\[2\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1784_ core.osr.result_r\[16\] net73 core.osr.next_result_w\[16\] net59 VSS VDD VSS
+ VDD sky130_fd_sc_hd__dfrtp_1
XANTENNA__1346__C _0212_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_130_104 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1719__RESET_B net63 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_84_213 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1218_ VSS VDD _0586_ _0394_ core.cnb.data_register_r\[7\] _0595_ VSS VDD sky130_fd_sc_hd__mux2_1
X_1149_ core.cnb.nswitch_out\[1\] core.cnb.pswitch_out\[1\] VDD VSS VSS VDD sky130_fd_sc_hd__inv_2
XANTENNA__1537__B _0077_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_106_112 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_136_77 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1475__B1 _0423_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_83_290 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_330 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_341 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_352 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_363 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_374 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_385 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_61_84 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XPHY_396 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_112_104 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1003_ _0266_ _0404_ _0428_ _0359_ _0415_ VSS VDD VSS VDD sky130_fd_sc_hd__o211ai_1
XANTENNA__1218__A0 core.cnb.data_register_r\[7\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1767_ net42 net70 _0030_ net59 VSS VDD VSS VDD sky130_fd_sc_hd__dfrtp_1
X_1698_ VSS VDD _0614_ _0252_ core.cnb.shift_register_r\[12\] _0201_ VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_122_13 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_122_68 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_15_44 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_31_87 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xoutput43 VDD VSS result_out[1] net43 VSS VDD sky130_fd_sc_hd__buf_2
XANTENNA_input30_A config_2_in[7] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_88_382 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_31_113 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_160 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_193 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_171 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_182 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_82_7 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1621_ core.osr.next_result_w\[8\] _0146_ core.osr.next_result_w\[10\] _0230_ _0124_
+ VSS VDD VSS VDD sky130_fd_sc_hd__o22a_1
X_1552_ VSS VDD _0005_ _0092_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XANTENNA__1193__A core.cnb.shift_register_r\[2\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1483_ _0056_ _0057_ core.cnb.data_register_r\[10\] VSS VDD VSS VDD sky130_fd_sc_hd__nor2_1
XFILLER_50_444 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_50_466 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_89_135 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_117_57 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_89_179 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1678__A0 core.cnb.shift_register_r\[2\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_13_113 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_pmat_col_n[5] core.pdc.col_out_n\[5\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1278__A _0635_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_6_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1770__CLK net55 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_3_69 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_92_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_83_71 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_91_388 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_0983_ VSS VDD _0366_ _0406_ _0405_ _0409_ _0408_ _0359_ VSS VDD sky130_fd_sc_hd__a41o_1
XANTENNA__0820__A core.cnb.shift_register_r\[2\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1604_ core.osr.next_result_w\[2\] _0131_ _0130_ _0115_ _0123_ _0232_ VSS VDD VSS
+ VDD sky130_fd_sc_hd__o221a_1
X_1535_ _0080_ _0079_ net52 core.pdc.row_out_n\[11\] VDD VSS VSS VDD sky130_fd_sc_hd__a21o_1
X_1466_ _0354_ core.ndc.col_out_n\[22\] _0505_ _0525_ VDD VSS VSS VDD sky130_fd_sc_hd__o21bai_1
X_1397_ _0729_ core.osr.result_r\[16\] core.osr.result_r\[12\] _0741_ _0743_ VSS VDD
+ VSS VDD sky130_fd_sc_hd__a31o_1
XFILLER_82_322 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_83_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1793__CLK net76 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_6_109 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1545__B _0568_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_88_38 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1363__A2 core.cnb.result_out\[8\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_fanout80_A net81 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_pmat_col_n[29] core.pdc.col_out_n\[29\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_85_160 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_37_53 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_74_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_53_41 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0905__A core.cnb.data_register_r\[5\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_52_8 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1320_ core.cnb.result_out\[6\] _0674_ core.osr.result_r\[7\] _0675_ core.osr.result_r\[6\]
+ VDD VSS VSS VDD sky130_fd_sc_hd__a211oi_1
XANTENNA__1354__A2 _0635_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_2_871 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1251_ VSS VDD _0561_ _0620_ core.cnb.average_counter_r\[3\] VSS VDD sky130_fd_sc_hd__xnor2_1
X_1182_ _0566_ core.cnb.average_counter_r\[3\] core.cnb.average_counter_r\[2\] _0560_
+ _0564_ _0565_ VSS VDD VSS VDD sky130_fd_sc_hd__o311a_1
XFILLER_65_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_91_174 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_0966_ _0359_ _0370_ _0392_ _0383_ _0325_ _0372_ VSS VDD VSS VDD sky130_fd_sc_hd__a311o_1
X_0897_ core.cnb.data_register_r\[5\] _0323_ VDD VSS VSS VDD sky130_fd_sc_hd__inv_2
X_1518_ _0607_ net52 _0079_ core.pdc.row_out_n\[6\] VSS VDD VSS VDD sky130_fd_sc_hd__o21a_2
XFILLER_87_414 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1449_ _0474_ _0772_ core.ndc.col_out_n\[9\] _0448_ VDD VSS VSS VDD sky130_fd_sc_hd__a21oi_1
XFILLER_114_25 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xvcm clk_vcm vcm/vcm VDD VSS adc_vcm_generator
XFILLER_114_47 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_56_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_130_79 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_136_121 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1033__A1 _0424_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_3_3 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_2_123 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_48_41 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_48_85 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_15 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_46_322 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_47_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_64_40 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_46_377 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_46_399 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_9_57 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_0820_ core.cnb.shift_register_r\[6\] core.cnb.shift_register_r\[2\] _0246_ core.cnb.shift_register_r\[3\]
+ core.cnb.shift_register_r\[16\] VDD VSS VSS VDD sky130_fd_sc_hd__or4_1
X_1303_ _0651_ _0659_ _0658_ _0653_ _0660_ VSS VDD VSS VDD sky130_fd_sc_hd__a31o_1
X_1234_ core.cnb.next_data_register_w\[9\] _0579_ _0608_ _0607_ VSS VDD VSS VDD sky130_fd_sc_hd__o21a_1
XFILLER_49_193 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1165_ core.cnb.data_register_r\[9\] _0552_ VDD VSS VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_38_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_92_461 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1096_ _0511_ _0510_ _0509_ _0448_ core.pdc.col_out_n\[10\] VSS VDD VSS VDD sky130_fd_sc_hd__o211a_1
XFILLER_52_358 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xadc_top_85 dummypin[0] adc_top_85/HI VDD VSS VSS VDD sky130_fd_sc_hd__conb_1
Xadc_top_96 dummypin[11] adc_top_96/HI VDD VSS VSS VDD sky130_fd_sc_hd__conb_1
X_0949_ _0363_ _0375_ _0374_ VSS VDD VSS VDD sky130_fd_sc_hd__or2_1
XFILLER_133_102 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_133_113 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_125_68 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_125_57 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_125_46 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_29_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_18_55 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XPHY_501 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_534 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_523 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_512 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_34_54 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XPHY_556 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_545 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_50_75 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1286__A _0635_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_124_124 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_pmat_sample_n sample_pmatrix_cgen_n VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_46_185 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_91_82 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_0803_ _0230_ core.osr.osr_mode_r\[0\] _0229_ VSS VDD VSS VDD sky130_fd_sc_hd__nand2_2
X_1783_ core.osr.result_r\[15\] net73 core.osr.next_result_w\[15\] net55 VSS VDD VSS
+ VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_115_113 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_115_124 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_130_116 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1217_ VSS VDD core.cnb.next_data_register_w\[6\] _0594_ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_1148_ core.cnb.nswitch_out\[1\] _0538_ _0403_ VSS VDD VSS VDD sky130_fd_sc_hd__xnor2_4
XFILLER_111_26 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1079_ _0394_ _0499_ VDD VSS VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_20_34 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_106_124 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_29_87 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1475__A1 _0450_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1227__B2 core.cnb.data_register_r\[7\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XPHY_320 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_331 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_342 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_353 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_364 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_375 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_386 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_61_63 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_397 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_86_71 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_1002_ _0427_ _0346_ _0350_ VSS VDD VSS VDD sky130_fd_sc_hd__nand2_4
XANTENNA__1466__A1 _0354_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1218__A1 _0394_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1766_ net41 net70 _0029_ net59 VSS VDD VSS VDD sky130_fd_sc_hd__dfrtp_1
X_1697_ VSS VDD _0042_ _0200_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_100_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1457__A1 _0354_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_40_114 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_31_77 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0983__A3 _0366_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xoutput44 VDD VSS result_out[2] net44 VSS VDD sky130_fd_sc_hd__buf_2
XFILLER_48_203 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA_input23_A config_2_in[15] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_56_74 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1448__B2 _0449_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1448__A1 _0466_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XPHY_161 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_150 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_172 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_194 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_183 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_1620_ _0214_ _0145_ _0144_ VSS VDD VSS VDD sky130_fd_sc_hd__or2_1
X_1551_ VSS VDD _0089_ core.cnb.next_data_register_w\[2\] core.cnb.result_out\[2\]
+ _0092_ VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_98_103 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1482_ _0056_ _0541_ _0344_ VSS VDD VSS VDD sky130_fd_sc_hd__nand2_1
XANTENNA__0818__A core.cnb.shift_register_r\[1\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1439__A1 _0354_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1749_ core.cnb.result_out\[9\] net64 _0012_ net79 VSS VDD VSS VDD sky130_fd_sc_hd__dfrtp_4
XFILLER_117_69 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_89_158 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_133_57 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_85_364 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_93_17 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_pmat_col_n[4] core.pdc.col_out_n\[4\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_3_15 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_67_40 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1118__B1 _0514_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_107_80 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_92_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_0982_ _0364_ _0337_ _0408_ core.cnb.data_register_r\[5\] _0407_ VDD VSS VSS VDD
+ sky130_fd_sc_hd__a22o_1
XFILLER_66_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_1603_ VSS VDD _0110_ core.osr.next_result_w\[6\] core.osr.next_result_w\[4\] _0130_
+ VSS VDD sky130_fd_sc_hd__mux2_1
X_1534_ core.pdc.row_out_n\[7\] _0079_ net52 _0080_ VSS VDD VSS VDD sky130_fd_sc_hd__o21a_1
X_1465_ _0474_ _0527_ core.ndc.col_out_n\[21\] _0470_ VDD VSS VSS VDD sky130_fd_sc_hd__a21oi_1
X_1396_ _0729_ core.osr.result_r\[16\] _0742_ _0741_ core.osr.result_r\[12\] VDD VSS
+ VSS VDD sky130_fd_sc_hd__nand4_1
XFILLER_82_356 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_83_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_82_389 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_50_220 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_50_253 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA_fanout73_A net74 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_37_98 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_74_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_2_883 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_1250_ _0618_ _0616_ core.cnb.next_average_counter_w\[2\] _0619_ VDD VSS VSS VDD
+ sky130_fd_sc_hd__a21oi_1
X_1181_ core.cnb.average_counter_r\[3\] core.cnb.sampled_avg_control_r\[1\] core.cnb.sampled_avg_control_r\[2\]
+ _0565_ _0561_ VDD VSS VSS VDD sky130_fd_sc_hd__or4b_1
XFILLER_65_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_91_153 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_94_93 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_91_186 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_0965_ VSS VDD _0391_ _0390_ _0386_ _0389_ _0325_ VSS VDD sky130_fd_sc_hd__a211o_1
X_0896_ _0322_ _0319_ _0321_ _0289_ core.cnb.data_register_r\[4\] _0304_ VSS VDD VSS
+ VDD sky130_fd_sc_hd__a32o_1
X_1517_ VSS VDD _0080_ _0079_ net52 core.ndc.row_out_n\[9\] VSS VDD sky130_fd_sc_hd__o21ai_1
X_1448_ _0772_ _0507_ _0449_ _0503_ _0466_ _0509_ VSS VDD VSS VDD sky130_fd_sc_hd__a32o_1
X_1379_ _0729_ _0728_ _0727_ _0721_ _0722_ VSS VDD VSS VDD sky130_fd_sc_hd__a31o_2
XFILLER_56_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_130_25 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_130_58 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_99_49 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1572__A net12 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_48_97 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_46_356 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_47_879 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_9_14 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_70_871 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_9_69 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_80_73 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_127_100 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_1302_ core.cnb.result_out\[4\] _0659_ VDD VSS VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_49_150 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_1233_ _0552_ _0588_ _0608_ _0579_ VDD VSS VSS VDD sky130_fd_sc_hd__a21oi_1
XANTENNA__1340__A_N core.cnb.result_out\[7\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1164_ _0328_ core.cnb.data_register_r\[8\] _0344_ _0342_ _0551_ VSS VDD VSS VDD
+ sky130_fd_sc_hd__a31o_1
XFILLER_38_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_92_440 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1783__CLK net55 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_52_304 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1095_ _0466_ _0511_ _0475_ VSS VDD VSS VDD sky130_fd_sc_hd__or2_1
XFILLER_52_348 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_0948_ _0374_ _0373_ _0366_ VSS VDD VSS VDD sky130_fd_sc_hd__xnor2_4
Xadc_top_86 dummypin[1] adc_top_86/HI VDD VSS VSS VDD sky130_fd_sc_hd__conb_1
XFILLER_133_125 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xadc_top_97 dummypin[12] adc_top_97/HI VDD VSS VSS VDD sky130_fd_sc_hd__conb_1
X_0879_ _0305_ _0301_ _0304_ _0303_ core.cnb.data_register_r\[6\] _0282_ VSS VDD VSS
+ VDD sky130_fd_sc_hd__a32o_1
XFILLER_87_289 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_29_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_18_45 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_18_78 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XPHY_535 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_524 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_513 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_502 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_557 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_546 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_51_370 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_51_381 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_133_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1567__A net53 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1190__A1 core.cnb.comparator_in VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_46_197 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_0802_ _0229_ _0214_ _0213_ VSS VDD VSS VDD sky130_fd_sc_hd__and2b_1
X_1782_ core.osr.result_r\[14\] net70 core.osr.next_result_w\[14\] net59 VSS VDD VSS
+ VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_130_128 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1216_ VDD VSS _0594_ _0593_ net53 VSS VDD sky130_fd_sc_hd__and2_1
XFILLER_84_259 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1799__RESET_B net63 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1147_ _0538_ _0296_ _0537_ VSS VDD VSS VDD sky130_fd_sc_hd__nand2_2
XFILLER_1_81 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_52_134 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA_nmat_col_n[5] core.ndc.col_out_n\[5\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1078_ _0474_ _0476_ core.pdc.col_out_n\[5\] _0450_ _0498_ VDD VSS VSS VDD sky130_fd_sc_hd__a22o_1
XFILLER_20_79 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_45_76 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_310 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_321 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_332 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_343 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_354 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_365 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_376 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_101_82 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_387 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_398 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_6_15 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_47_440 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1001_ _0426_ _0405_ _0359_ VSS VDD VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_47_462 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1000__A _0364_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1765_ net40 net70 _0028_ net59 VSS VDD VSS VDD sky130_fd_sc_hd__dfrtp_1
X_1696_ VSS VDD _0614_ core.cnb.shift_register_r\[12\] core.cnb.shift_register_r\[11\]
+ _0200_ VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_100_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1670__A _0110_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_122_37 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_53_454 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_40_104 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_15_57 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_31_45 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xoutput45 VDD VSS result_out[3] net45 VSS VDD sky130_fd_sc_hd__buf_2
XFILLER_48_237 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_56_20 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1580__A core.osr.osr_mode_r\[0\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_input16_A config_1_in[9] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_56_64 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_16_123 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0924__A _0347_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XPHY_140 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_151 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_184 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_173 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_162 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_9_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XPHY_195 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_1550_ VSS VDD _0004_ _0091_ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_1481_ VSS VDD _1481_/X _0055_ VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_97_82 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_11_3 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__0818__B core.cnb.is_sampling_w VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1439__A2 _0465_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_54_229 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_50_457 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_1817_ core.osr.data_valid_r net71 core.osr.is_last_sample net57 VSS VDD VSS VDD
+ sky130_fd_sc_hd__dfrtp_1
X_1748_ core.cnb.result_out\[8\] net65 _0011_ net78 VSS VDD VSS VDD sky130_fd_sc_hd__dfrtp_4
XANTENNA__1717__CLK net81 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_117_26 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1679_ VSS VDD _0033_ _0191_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XANTENNA__1127__A1 _0529_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_input8_A config_1_in[1] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_133_69 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_26_34 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_pmat_col_n[3] core.pdc.col_out_n\[3\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_3_27 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1118__A1 _0354_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_67_52 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_88_192 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_83_84 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_83_95 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_0981_ _0364_ _0289_ _0407_ _0318_ _0344_ _0320_ VSS VDD VSS VDD sky130_fd_sc_hd__a311o_1
X_1602_ core.osr.next_result_w\[8\] _0129_ _0124_ VSS VDD VSS VDD sky130_fd_sc_hd__or2_1
X_1533_ core.pdc.row_out_n\[5\] _0079_ net52 _0081_ VSS VDD VSS VDD sky130_fd_sc_hd__o21a_1
X_1464_ VSS VDD _0515_ _0424_ _0511_ core.ndc.col_out_n\[20\] VSS VDD sky130_fd_sc_hd__o21ai_1
X_1395_ VSS VDD _0741_ core.osr.result_r\[14\] core.osr.result_r\[13\] core.osr.result_r\[15\]
+ VSS VDD sky130_fd_sc_hd__and3_1
XFILLER_82_302 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_50_232 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_50_265 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_12_14 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_128_69 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA_nmat_sample_n sample_nmatrix_cgen_n VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_fanout66_A net67 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_85_184 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_53_21 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_38_8 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_49_321 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1180_ core.cnb.average_counter_r\[3\] _0561_ _0564_ _0563_ _0562_ VDD VSS VSS VDD
+ sky130_fd_sc_hd__a22o_1
XFILLER_94_50 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_91_143 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_91_165 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_0964_ _0390_ _0366_ _0331_ _0335_ _0377_ VSS VDD VSS VDD sky130_fd_sc_hd__and4_1
X_0895_ VSS VDD _0321_ core.cnb.data_register_r\[4\] core.cnb.data_register_r\[5\]
+ _0320_ VSS VDD sky130_fd_sc_hd__and3_1
X_1516_ core.pdc.row_out_n\[9\] core.ndc.row_out_n\[7\] VDD VSS VSS VDD sky130_fd_sc_hd__inv_2
X_1447_ _0529_ _0526_ core.ndc.col_out_n\[8\] _0452_ VDD VSS VSS VDD sky130_fd_sc_hd__a21oi_1
XFILLER_87_449 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1378_ VDD VSS _0728_ core.cnb.result_out\[11\] core.osr.result_r\[11\] VSS VDD sky130_fd_sc_hd__and2_1
XANTENNA__1569__B2 core.cnb.result_out\[10\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_139_57 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1572__B net11 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_48_76 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_64_64 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_104_93 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_9_26 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_70_883 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xfanout80 net81 net80 VSS VDD VSS VDD sky130_fd_sc_hd__clkbuf_2
XFILLER_80_85 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_89_50 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_1301_ core.osr.result_r\[4\] _0658_ VDD VSS VSS VDD sky130_fd_sc_hd__inv_2
X_1232_ _0607_ _0606_ _0605_ VSS VDD VSS VDD sky130_fd_sc_hd__xnor2_4
XANTENNA__1702__S _0614_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1163_ _0433_ _0549_ _0344_ _0545_ _0550_ VSS VDD VSS VDD sky130_fd_sc_hd__a31o_1
X_1094_ _0449_ _0510_ _0466_ VSS VDD VSS VDD sky130_fd_sc_hd__or2_1
XFILLER_100_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_0947_ _0373_ _0359_ _0370_ _0372_ VSS VDD VSS VDD sky130_fd_sc_hd__nand3_4
Xadc_top_87 dummypin[2] adc_top_87/HI VDD VSS VSS VDD sky130_fd_sc_hd__conb_1
XFILLER_109_16 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_109_38 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_0878_ _0261_ _0239_ _0304_ _0240_ _0268_ VSS VDD VSS VDD sky130_fd_sc_hd__nor4_4
Xadc_top_98 dummypin[13] adc_top_98/HI VDD VSS VSS VDD sky130_fd_sc_hd__conb_1
XFILLER_125_37 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_87_268 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_55_165 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_525 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_514 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_503 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_558 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_547 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_536 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_34_89 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_34_67 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_126_3 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1567__B _0089_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_50_99 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_75_41 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_75_63 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0927__A _0352_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_46_165 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_0801_ core.osr.osr_mode_r\[0\] _0228_ _0226_ _0222_ _0213_ _0227_ VSS VDD VSS VDD
+ sky130_fd_sc_hd__o221a_1
X_1781_ core.osr.result_r\[13\] net70 core.osr.next_result_w\[13\] net55 VSS VDD VSS
+ VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_115_104 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_41_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_84_205 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_1215_ VSS VDD _0586_ _0410_ core.cnb.data_register_r\[6\] _0593_ VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_84_249 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_1146_ VSS VDD _0295_ _0290_ core.cnb.data_register_r\[1\] _0537_ VSS VDD sky130_fd_sc_hd__o21ai_1
XFILLER_1_93 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA_nmat_col_n[4] core.ndc.col_out_n\[4\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1077_ _0498_ _0497_ _0477_ VSS VDD VSS VDD sky130_fd_sc_hd__nand2_1
XANTENNA__1641__A0 core.osr.next_result_w\[10\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_121_129 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_43_113 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_300 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_311 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_322 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_333 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_344 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_355 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_366 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_377 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_388 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_399 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1773__CLK net56 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1163__A2 _0433_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_86_40 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_1000_ _0365_ _0425_ _0364_ VSS VDD VSS VDD sky130_fd_sc_hd__nor2_1
XFILLER_47_474 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA_pmat_sample sample_pmatrix_cgen VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_cgen_nsample_p_in core.cnb.enable_loop_out VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1764_ net39 net70 _0027_ net59 VSS VDD VSS VDD sky130_fd_sc_hd__dfrtp_1
X_1695_ VSS VDD _0041_ _0199_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_25_113 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_53_400 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_15_14 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_1129_ _0446_ _0432_ _0506_ _0530_ VDD VSS VSS VDD sky130_fd_sc_hd__a21o_1
XFILLER_53_466 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_40_127 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1398__A _0635_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1796__CLK net76 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_31_68 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xoutput35 VDD VSS conversion_finished_out net35 VSS VDD sky130_fd_sc_hd__buf_2
Xoutput46 VDD VSS result_out[4] net46 VSS VDD sky130_fd_sc_hd__buf_2
XFILLER_88_330 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_88_374 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_48_249 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_16_102 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_152 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_141 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_130 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_185 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_163 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_174 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1101__A _0466_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XPHY_196 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__0940__A _0364_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_9_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_68_8 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_1480_ net15 net14 _0055_ net13 net16 VDD VSS VSS VDD sky130_fd_sc_hd__or4_1
XFILLER_98_127 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_95_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1816_ core.osr.osr_mode_r\[2\] net71 _0050_ net57 VSS VDD VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_7_81 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1747_ core.cnb.result_out\[7\] net68 _0010_ net81 VSS VDD VSS VDD sky130_fd_sc_hd__dfrtp_4
X_1678_ VSS VDD _0568_ core.cnb.shift_register_r\[3\] core.cnb.shift_register_r\[2\]
+ _0191_ VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_117_49 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1127__A2 _0506_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_133_15 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_86_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1783__RESET_B net73 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_13_105 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_10_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_3_39 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1118__A2 _0515_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_77_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_123_81 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_83_30 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA_pmat_sw core.cnb.is_sampling_w VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_0980_ _0406_ _0378_ VSS VDD VSS VDD sky130_fd_sc_hd__clkbuf_4
X_1601_ VSS VDD _0018_ _0128_ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_1532_ core.pdc.row_out_n\[4\] core.ndc.row_out_n\[12\] VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_2
X_1463_ VSS VDD core.ndc.col_out_n\[19\] _0051_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_86_119 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_68_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1394_ _0740_ core.osr.next_result_w\[15\] _0736_ VSS VDD VSS VDD sky130_fd_sc_hd__nor2_1
XFILLER_50_244 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_128_59 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_88_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA_pmat_col_n[26] core.pdc.col_out_n\[26\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_59_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_85_130 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_85_152 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_37_89 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA_fanout59_A core.cnb.conv_finished_r VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_53_33 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_91_122 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_91_133 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_0963_ VSS VDD core.cnb.data_register_r\[2\] _0307_ _0313_ _0389_ _0266_ VSS VDD
+ sky130_fd_sc_hd__a2bb2o_1
X_0894_ _0320_ core.cnb.shift_register_r\[9\] core.cnb.shift_register_r\[8\] VSS VDD
+ VSS VDD sky130_fd_sc_hd__and2b_1
X_1515_ core.pdc.row_out_n\[9\] _0556_ _0079_ _0353_ _0607_ VSS VDD VSS VDD sky130_fd_sc_hd__a31o_2
X_1446_ core.ndc.col_out_n\[7\] _0354_ _0506_ _0501_ VSS VDD VSS VDD sky130_fd_sc_hd__o21a_1
X_1377_ core.osr.result_r\[11\] _0727_ core.cnb.result_out\[11\] VSS VDD VSS VDD sky130_fd_sc_hd__or2_1
XFILLER_55_325 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_55_347 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_130_38 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_23_25 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_139_69 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1572__C net10 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_86_461 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_0_29 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_64_21 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_46_369 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_64_54 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_9_38 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_120_60 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xfanout81 VDD VSS net81 core.clk_dig_in VSS VDD sky130_fd_sc_hd__buf_2
Xfanout70 VDD VSS net70 net73 VSS VDD sky130_fd_sc_hd__buf_4
XFILLER_127_113 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_129_91 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1300_ _0657_ core.osr.next_result_w\[4\] VDD VSS VSS VDD sky130_fd_sc_hd__inv_2
X_1231_ VSS VDD _0606_ core.cnb.data_register_r\[9\] _0541_ VSS VDD sky130_fd_sc_hd__xnor2_2
XFILLER_49_174 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_1162_ VSS VDD _0544_ _0548_ _0542_ _0549_ VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_52_317 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1093_ _0427_ _0509_ _0453_ VSS VDD VSS VDD sky130_fd_sc_hd__or2_1
XFILLER_92_453 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_52_328 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_0946_ _0296_ _0371_ _0281_ _0297_ _0372_ VSS VDD VSS VDD sky130_fd_sc_hd__a31o_1
XFILLER_118_102 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xadc_top_99 dummypin[14] adc_top_99/HI VDD VSS VSS VDD sky130_fd_sc_hd__conb_1
X_0877_ _0302_ _0303_ _0252_ _0254_ VSS VDD VSS VDD sky130_fd_sc_hd__nor3_1
Xadc_top_88 dummypin[3] adc_top_88/HI VDD VSS VSS VDD sky130_fd_sc_hd__conb_1
XFILLER_87_225 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_87_236 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_130_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1429_ VDD VSS _0764_ _0762_ core.osr.sample_count_r\[6\] VSS VDD sky130_fd_sc_hd__and2_1
XFILLER_18_14 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1487__A1 _0328_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_83_442 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XPHY_526 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_515 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_504 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_559 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_548 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_537 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_109_113 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_109_124 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_121_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_46_177 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1104__A _0427_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__0943__A core.cnb.data_register_r\[2\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1650__A1 core.cnb.result_out\[7\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_0800_ VDD VSS _0227_ core.osr.sample_count_r\[0\] _0214_ VSS VDD sky130_fd_sc_hd__and2_1
XFILLER_24_90 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_1780_ core.osr.result_r\[12\] net67 core.osr.next_result_w\[12\] net54 VSS VDD VSS
+ VDD sky130_fd_sc_hd__dfrtp_2
XANTENNA__0913__B1 core.cnb.data_register_r\[7\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_112_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_1_50 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1469__A1 _0450_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1214_ VSS VDD core.cnb.next_data_register_w\[5\] _0592_ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_1145_ core.cnb.nswitch_out\[0\] core.cnb.pswitch_out\[0\] VDD VSS VSS VDD sky130_fd_sc_hd__inv_2
XANTENNA_nmat_col_n[3] core.ndc.col_out_n\[3\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_92_272 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1076_ _0491_ _0497_ _0484_ _0496_ VDD VSS VSS VDD sky130_fd_sc_hd__and3_2
X_0929_ _0355_ _0265_ core.cnb.data_register_r\[2\] _0251_ VSS VDD VSS VDD sky130_fd_sc_hd__nand3b_2
XFILLER_103_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_45_45 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_301 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_312 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_323 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_334 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_345 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_356 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_367 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_101_73 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1632__B2 core.osr.next_result_w\[8\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XPHY_378 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_389 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_101_95 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_112_119 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_20_9 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_13_8 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_47_431 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_86_96 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_19_90 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1763_ net38 net66 _0026_ net54 VSS VDD VSS VDD sky130_fd_sc_hd__dfrtp_1
X_1694_ VSS VDD _0614_ core.cnb.shift_register_r\[11\] core.cnb.shift_register_r\[10\]
+ _0199_ VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_89_309 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_103_119 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__0848__A core.cnb.shift_register_r\[2\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1128_ _0352_ _0452_ core.pdc.col_out_n\[24\] _0462_ _0503_ VDD VSS VSS VDD sky130_fd_sc_hd__a22o_1
X_1059_ _0364_ _0480_ _0365_ VSS VDD VSS VDD sky130_fd_sc_hd__or2_1
XANTENNA_nmat_row_n[12] core.ndc.row_out_n\[12\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xoutput36 VDD VSS result_out[0] net36 VSS VDD sky130_fd_sc_hd__buf_2
Xoutput47 VDD VSS result_out[5] net47 VSS VDD sky130_fd_sc_hd__buf_2
XFILLER_88_342 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_56_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_88_397 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1589__A _0110_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_112_50 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_72_21 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_112_72 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_112_94 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_131 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_120 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_142 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_72_65 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_72_76 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_164 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_153 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_175 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1101__B _0468_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XPHY_197 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_186 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_21_91 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_97_51 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_97_95 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_95_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_47_250 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_47_272 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_47_294 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_0 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_50_415 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1815_ core.osr.osr_mode_r\[1\] net71 _0049_ net57 VSS VDD VSS VDD sky130_fd_sc_hd__dfrtp_1
X_1746_ core.cnb.result_out\[6\] net67 _0009_ net79 VSS VDD VSS VDD sky130_fd_sc_hd__dfrtp_4
XFILLER_7_93 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1677_ _0615_ core.cnb.shift_register_r\[1\] _0089_ _0032_ VDD VSS VSS VDD sky130_fd_sc_hd__a21o_1
XFILLER_133_27 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_86_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_85_378 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_26_69 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_13_128 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_pmat_col_n[1] core.pdc.col_out_n\[1\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1599__B1 core.osr.next_result_w\[7\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_10_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_101_3 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_67_87 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_77_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA_input21_A config_2_in[13] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_91_337 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_83_64 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_8_121 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__0801__A2 core.osr.osr_mode_r\[0\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1600_ VSS VDD _0235_ _0127_ _0122_ _0128_ VSS VDD sky130_fd_sc_hd__mux2_1
X_1531_ core.ndc.row_out_n\[12\] core.pdc.row_out_n\[3\] _0074_ VSS VDD VSS VDD sky130_fd_sc_hd__nor2_1
X_1462_ _0516_ _0449_ _0051_ _0512_ VSS VDD VSS VDD sky130_fd_sc_hd__o21ba_1
X_1393_ VSS VDD _0739_ _0740_ core.osr.result_r\[15\] VSS VDD sky130_fd_sc_hd__xnor2_1
XFILLER_68_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__0861__A core.cnb.data_register_r\[0\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_10_109 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1729_ core.cnb.sampled_avg_control_r\[2\] net60 _0002_ net75 VSS VDD VSS VDD sky130_fd_sc_hd__dfrtp_2
XANTENNA_pmat_col_n[25] core.pdc.col_out_n\[25\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_59_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_5_113 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1541__S _0588_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_49_367 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_94_85 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_0962_ _0383_ _0388_ _0384_ _0387_ _0333_ _0385_ VSS VDD VSS VDD sky130_fd_sc_hd__o221a_1
X_0893_ _0259_ _0319_ VDD VSS VSS VDD sky130_fd_sc_hd__inv_2
X_1514_ core.pdc.row_out_n\[10\] core.ndc.row_out_n\[6\] VDD VSS VSS VDD sky130_fd_sc_hd__inv_2
X_1445_ _0529_ _0504_ core.ndc.col_out_n\[6\] _0771_ VDD VSS VSS VDD sky130_fd_sc_hd__a21oi_1
X_1376_ _0726_ core.osr.next_result_w\[11\] VDD VSS VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_114_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_55_304 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_55_359 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_2_116 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_48_34 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_fanout71_A net73 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_46_315 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_86_473 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_46_337 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_46_348 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xfanout71 VDD VSS net71 net73 VSS VDD sky130_fd_sc_hd__buf_4
Xfanout60 net60 net61 VSS VDD VSS VDD sky130_fd_sc_hd__clkbuf_4
XFILLER_80_54 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_13_81 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_50_9 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_43_8 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1230_ _0605_ _0598_ _0551_ _0604_ VSS VDD VSS VDD sky130_fd_sc_hd__a21boi_4
X_1161_ VSS VDD _0548_ core.cnb.data_register_r\[10\] core.cnb.data_register_r\[9\]
+ _0541_ VSS VDD sky130_fd_sc_hd__and3_1
XFILLER_92_410 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_49_186 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1092_ _0508_ core.pdc.col_out_n\[9\] _0507_ _0448_ VSS VDD VSS VDD sky130_fd_sc_hd__o21ai_2
X_0945_ _0307_ _0313_ _0371_ _0251_ _0265_ VSS VDD VSS VDD sky130_fd_sc_hd__o211ai_1
X_0876_ VSS VDD _0255_ _0302_ core.cnb.shift_register_r\[12\] VSS VDD sky130_fd_sc_hd__xnor2_1
Xadc_top_89 dummypin[4] adc_top_89/HI VDD VSS VSS VDD sky130_fd_sc_hd__conb_1
XANTENNA__1708__A0 _0110_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_130_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1428_ _0763_ core.osr.next_sample_count_w\[6\] core.osr.is_last_sample VSS VDD VSS
+ VDD sky130_fd_sc_hd__nor2_1
XFILLER_18_37 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1487__A2 _0342_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1359_ core.cnb.result_out\[8\] core.osr.result_r\[8\] core.osr.result_r\[9\] _0711_
+ VDD VSS VSS VDD sky130_fd_sc_hd__a21o_1
XFILLER_83_454 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XPHY_516 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_505 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_549 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_538 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_527 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1210__A _0364_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_50_57 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_50_68 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_121_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_46_101 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0943__B core.cnb.data_register_r\[1\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_91_53 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_112_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1213_ VDD VSS _0592_ _0591_ net53 VSS VDD sky130_fd_sc_hd__and2_1
XANTENNA__1469__A2 _0506_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1144_ core.cnb.nswitch_out\[0\] _0536_ core.cnb.data_register_r\[0\] VSS VDD VSS
+ VDD sky130_fd_sc_hd__xnor2_4
X_1075_ _0433_ _0493_ _0496_ _0434_ _0494_ _0492_ _0495_ VSS VDD VSS VDD sky130_fd_sc_hd__mux4_1
XANTENNA_pmat_rowon_n[13] core.pdc.row_out_n\[14\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_20_16 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_0928_ VDD VSS _0354_ _0353_ VSS VDD sky130_fd_sc_hd__buf_4
XFILLER_136_16 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_0859_ _0284_ _0285_ _0268_ _0283_ VSS VDD VSS VDD sky130_fd_sc_hd__nor3_1
XFILLER_20_49 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_106_106 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1777__RESET_B net69 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_103_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_28_112 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1205__A _0579_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_45_57 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_302 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_313 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_324 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_61_23 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_335 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_346 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_357 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_368 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_131_3 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XPHY_379 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_6_29 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_86_64 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_47_421 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_47_454 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1320__A1 core.cnb.result_out\[6\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1762_ net37 net70 _0025_ net59 VSS VDD VSS VDD sky130_fd_sc_hd__dfrtp_1
X_1693_ VSS VDD _0040_ _0198_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XANTENNA__1025__A _0449_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1127_ _0529_ _0505_ core.pdc.col_out_n\[23\] _0506_ VDD VSS VSS VDD sky130_fd_sc_hd__a21oi_1
X_1058_ _0345_ _0479_ _0478_ _0406_ VDD VSS VSS VDD sky130_fd_sc_hd__or3_1
XFILLER_31_15 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xoutput37 VDD VSS result_out[10] net37 VSS VDD sky130_fd_sc_hd__buf_2
Xoutput48 VDD VSS result_out[6] net48 VSS VDD sky130_fd_sc_hd__buf_2
XFILLER_88_365 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_48_229 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_16_115 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XPHY_132 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_121 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_110 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_143 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_176 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_165 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_154 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_187 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_198 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_137_81 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XPHY_1 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_94_3 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1814_ core.osr.osr_mode_r\[0\] net70 _0048_ net59 VSS VDD VSS VDD sky130_fd_sc_hd__dfrtp_4
XFILLER_7_50 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_1745_ core.cnb.result_out\[5\] net65 _0008_ net79 VSS VDD VSS VDD sky130_fd_sc_hd__dfrtp_4
X_1676_ _0615_ _0588_ core.cnb.next_conv_finished_w _0031_ VDD VSS VSS VDD sky130_fd_sc_hd__a21o_1
XFILLER_133_39 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_85_324 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_85_346 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_85_357 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_26_15 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_53_276 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_pmat_col_n[0] core.pdc.col_out_n\[0\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_42_14 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA_pmat_analog_in inp_analog VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xpmat_84 net84 pmat_84/HI VDD VSS VSS VDD sky130_fd_sc_hd__conb_1
XFILLER_88_151 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_input14_A config_1_in[7] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__0798__C1 core.osr.osr_mode_r\[0\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1539__S _0588_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_73_8 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1530_ core.ndc.row_out_n\[12\] core.pdc.row_out_n\[1\] _0077_ VSS VDD VSS VDD sky130_fd_sc_hd__nor2_1
X_1461_ VSS VDD _0519_ _0424_ _0514_ core.ndc.col_out_n\[18\] VSS VDD sky130_fd_sc_hd__o21ai_1
X_1392_ _0739_ core.osr.result_r\[14\] core.osr.result_r\[12\] core.osr.result_r\[13\]
+ _0729_ VSS VDD VSS VDD sky130_fd_sc_hd__and4_1
XFILLER_94_121 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_82_316 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_90_382 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1202__A0 core.cnb.nswitch_out\[2\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1728_ core.cnb.sampled_avg_control_r\[1\] net60 _0001_ net75 VSS VDD VSS VDD sky130_fd_sc_hd__dfrtp_2
XANTENNA_pmat_col_n[24] core.pdc.col_out_n\[24\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1659_ core.osr.next_result_w\[11\] _0177_ core.osr.next_result_w\[13\] _0235_ _0219_
+ _0154_ VSS VDD VSS VDD sky130_fd_sc_hd__o221a_1
XANTENNA_input6_A config_1_in[14] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1213__A net53 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_53_57 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_5_125 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_49_357 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_49_379 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_0961_ _0338_ _0387_ _0325_ _0386_ core.cnb.data_register_r\[6\] VDD VSS VSS VDD
+ sky130_fd_sc_hd__o2bb2a_1
X_0892_ _0318_ _0316_ _0317_ _0289_ _0315_ _0282_ VSS VDD VSS VDD sky130_fd_sc_hd__a32o_1
XFILLER_57_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1753__CLK net55 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1513_ core.pdc.row_out_n\[10\] net52 _0607_ _0079_ VSS VDD VSS VDD sky130_fd_sc_hd__a21o_2
XFILLER_87_408 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1444_ _0771_ _0452_ _0497_ VSS VDD VSS VDD sky130_fd_sc_hd__nand2b_1
X_1375_ _0725_ _0726_ core.cnb.result_out\[11\] VDD VSS VSS VDD sky130_fd_sc_hd__xor2_1
XFILLER_82_102 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_82_124 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_48_390 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_82_179 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_128_9 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1208__A core.cnb.is_sampling_w VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_fanout64_A net67 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_64_34 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_104_85 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__0782__A net12 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_80_11 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xfanout72 net73 net72 VSS VDD VSS VDD sky130_fd_sc_hd__clkbuf_2
Xfanout61 net61 net62 VSS VDD VSS VDD sky130_fd_sc_hd__clkbuf_4
XANTENNA__1776__CLK net56 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_13_93 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_129_82 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_89_20 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_49_132 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_89_290 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_49_165 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_1160_ VSS VDD _0547_ _0545_ core.cnb.data_register_r\[8\] _0546_ VSS VDD sky130_fd_sc_hd__and3_1
X_1091_ _0500_ _0353_ _0499_ _0508_ VDD VSS VSS VDD sky130_fd_sc_hd__a21o_1
XFILLER_92_477 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_0944_ _0368_ _0314_ _0355_ _0369_ _0370_ VSS VDD VSS VDD sky130_fd_sc_hd__a31o_1
X_0875_ _0277_ _0301_ _0268_ _0242_ VSS VDD VSS VDD sky130_fd_sc_hd__nor3_1
XANTENNA__1708__A1 net10 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1028__A _0410_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1427_ VSS VDD _0762_ _0763_ core.osr.sample_count_r\[6\] VSS VDD sky130_fd_sc_hd__xnor2_1
XFILLER_83_411 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1358_ core.cnb.result_out\[8\] core.cnb.result_out\[9\] core.osr.result_r\[8\] core.osr.result_r\[9\]
+ _0710_ VSS VDD VSS VDD sky130_fd_sc_hd__a31o_1
XFILLER_83_466 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1289_ VSS VDD _0647_ _0648_ core.osr.result_r\[3\] VSS VDD sky130_fd_sc_hd__xnor2_1
XPHY_517 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_506 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_34_15 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1644__B1 _0236_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XPHY_539 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_528 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1799__CLK net77 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_50_47 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_46_124 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_54_190 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_91_21 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_24_81 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1547__S _0089_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_115_118 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xnmat_82 net82 nmat_82/HI VDD VSS VSS VDD sky130_fd_sc_hd__conb_1
X_1212_ VSS VDD _0586_ _0420_ core.cnb.data_register_r\[5\] _0591_ VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_37_113 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1143_ _0535_ _0270_ _0397_ _0536_ VSS VDD VSS VDD sky130_fd_sc_hd__a21oi_2
XFILLER_92_230 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA_nmat_col_n[1] core.ndc.col_out_n\[1\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_52_105 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1074_ _0347_ _0495_ _0480_ _0444_ VDD VSS VSS VDD sky130_fd_sc_hd__or3_1
XFILLER_52_149 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_nmat_sw core.cnb.is_sampling_w VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1030__B _0374_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_0927_ VDD VSS _0353_ _0352_ VSS VDD sky130_fd_sc_hd__buf_4
X_0858_ _0254_ core.cnb.shift_register_r\[11\] _0284_ core.cnb.shift_register_r\[12\]
+ _0255_ VDD VSS VSS VDD sky130_fd_sc_hd__or4_1
XFILLER_106_118 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_0789_ _0216_ core.osr.osr_mode_r\[0\] VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_2
XFILLER_29_15 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_28_124 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_83_230 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1746__RESET_B net67 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_83_296 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_303 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_314 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_325 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_101_31 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_101_42 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_336 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_347 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_358 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_61_46 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_61_35 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_40_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XPHY_369 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_124_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_120_121 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_19_124 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1131__A _0352_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_31_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1761_ net51 net66 _0024_ net54 VSS VDD VSS VDD sky130_fd_sc_hd__dfrtp_1
X_1692_ VSS VDD _0614_ core.cnb.shift_register_r\[10\] core.cnb.shift_register_r\[9\]
+ _0198_ VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_98_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1306__A _0634_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1126_ _0529_ _0449_ VSS VDD VSS VDD sky130_fd_sc_hd__clkbuf_4
XFILLER_53_425 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_53_436 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_1057_ _0478_ _0365_ _0364_ VSS VDD VSS VDD sky130_fd_sc_hd__nand2_1
XANTENNA_cgen_dlycontrol4_in[5] net7 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_22_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_31_38 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_110_9 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xoutput38 VDD VSS result_out[11] net38 VSS VDD sky130_fd_sc_hd__buf_2
Xoutput49 VDD VSS result_out[7] net49 VSS VDD sky130_fd_sc_hd__buf_2
XFILLER_89_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1216__A net53 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_56_57 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_100 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_112_85 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_133 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_31_108 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_31_119 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_122 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_111 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_144 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_13_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XPHY_155 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_166 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_177 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_188 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_199 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_137_93 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__0949__B _0374_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1126__A _0449_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_47_241 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_2 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_1813_ core.osr.sample_count_r\[8\] net72 core.osr.next_sample_count_w\[8\] net58
+ VSS VDD VSS VDD sky130_fd_sc_hd__dfrtp_2
XANTENNA_nmat_sw_n core.cnb.enable_loop_out VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1744_ core.cnb.result_out\[4\] net65 _0007_ net78 VSS VDD VSS VDD sky130_fd_sc_hd__dfrtp_4
X_1675_ VSS VDD _0187_ _0188_ _0115_ _0030_ _0190_ _0123_ VSS VDD sky130_fd_sc_hd__a41o_1
XFILLER_53_233 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_1109_ _0520_ _0521_ _0466_ VSS VDD VSS VDD sky130_fd_sc_hd__nor2_1
XFILLER_13_119 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_53_299 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_42_37 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_107_63 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_107_74 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_67_34 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_88_163 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_91_317 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_84_380 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_91_328 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_16_93 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xpmat_102 pmat_102/LO net102 VDD VSS VSS VDD sky130_fd_sc_hd__conb_1
XANTENNA__1555__S _0089_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1460_ VSS VDD core.ndc.col_out_n\[17\] core.pdc.col_out_n\[16\] _0463_ _0353_ _0448_
+ VSS VDD sky130_fd_sc_hd__a31oi_1
X_1391_ _0738_ core.osr.next_result_w\[14\] _0736_ VSS VDD VSS VDD sky130_fd_sc_hd__nor2_1
XFILLER_82_328 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_50_214 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_50_258 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_12_29 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_128_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1202__A1 core.cnb.data_register_r\[2\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1727_ core.cnb.sampled_avg_control_r\[0\] net60 _0000_ net75 VSS VDD VSS VDD sky130_fd_sc_hd__dfrtp_2
X_1658_ _0132_ core.cnb.result_out\[9\] _0175_ _0176_ VDD VSS VSS VDD sky130_fd_sc_hd__a21o_1
XFILLER_85_100 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1589_ _0118_ _0657_ _0110_ VSS VDD VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_37_15 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_85_199 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA_pmat_row_n[9] core.pdc.row_out_n\[9\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_53_47 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_139_113 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1441__A1 _0529_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_118_51 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_89_461 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_91_169 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_0960_ _0386_ _0319_ _0304_ VSS VDD VSS VDD sky130_fd_sc_hd__nand2_1
X_0891_ _0317_ core.cnb.shift_register_r\[8\] core.cnb.shift_register_r\[9\] VSS VDD
+ VSS VDD sky130_fd_sc_hd__and2b_1
XANTENNA__1196__A0 core.cnb.nswitch_out\[0\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1512_ _0079_ net52 core.ndc.row_out_n\[5\] _0080_ VDD VSS VSS VDD sky130_fd_sc_hd__a21oi_1
X_1443_ VSS VDD core.ndc.col_out_n\[5\] _0770_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_4_41 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_4_85 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1374_ _0212_ _0725_ _0723_ _0724_ VDD VSS VSS VDD sky130_fd_sc_hd__or3_1
XFILLER_82_169 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1671__A1 _0110_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_133_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_48_47 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_104_20 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA_fanout57_A core.cnb.conv_finished_r VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_104_64 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__0782__B net11 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xfanout62 VDD VSS net62 net74 VSS VDD sky130_fd_sc_hd__buf_2
Xfanout73 VDD VSS net73 net74 VSS VDD sky130_fd_sc_hd__buf_2
XFILLER_80_67 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_124_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_49_199 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1090_ _0507_ _0463_ _0427_ VSS VDD VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_92_467 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_52_309 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1102__B1 _0515_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1653__B2 core.osr.next_result_w\[10\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_0943_ _0290_ core.cnb.data_register_r\[2\] _0369_ core.cnb.data_register_r\[1\]
+ _0295_ VDD VSS VSS VDD sky130_fd_sc_hd__or4_1
X_0874_ _0299_ _0300_ _0264_ VSS VDD VSS VDD sky130_fd_sc_hd__nor2_1
XANTENNA__1309__A core.cnb.result_out\[5\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_115_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1426_ VSS VDD _0762_ core.osr.sample_count_r\[5\] core.osr.sample_count_r\[4\] _0757_
+ VSS VDD sky130_fd_sc_hd__and3_1
X_1357_ _0709_ core.osr.next_result_w\[9\] VDD VSS VSS VDD sky130_fd_sc_hd__inv_2
XANTENNA__1044__A _0410_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_83_423 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_1288_ _0647_ _0640_ _0644_ _0645_ VDD VSS VSS VDD sky130_fd_sc_hd__a21boi_1
XANTENNA__0883__A core.cnb.shift_register_r\[2\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_55_169 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_83_478 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_507 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1644__A1 core.cnb.result_out\[6\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XPHY_529 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_518 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_51_364 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_51_397 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1219__A net53 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_106_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_59_57 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_86_294 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1743__CLK net81 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_91_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_91_33 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_91_88 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1774__D core.osr.next_result_w\[6\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_40_92 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xnmat_83 net83 nmat_83/HI VDD VSS VSS VDD sky130_fd_sc_hd__conb_1
XANTENNA__0968__A core.cnb.data_register_r\[7\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1211_ _0590_ core.cnb.next_data_register_w\[4\] _0588_ VSS VDD VSS VDD sky130_fd_sc_hd__nor2_1
XANTENNA__1323__B1 core.cnb.result_out\[6\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1142_ _0289_ _0286_ _0535_ _0282_ _0285_ VDD VSS VSS VDD sky130_fd_sc_hd__a22o_1
X_1073_ _0345_ _0494_ _0480_ _0444_ VDD VSS VSS VDD sky130_fd_sc_hd__or3_1
X_0926_ _0352_ _0351_ VSS VDD VSS VDD sky130_fd_sc_hd__clkbuf_8
Xpmat pmat/vcm sample_pmatrix_cgen sample_pmatrix_cgen_n core.pdc.row_out_n\[15\]
+ core.pdc.row_out_n\[14\] core.pdc.row_out_n\[13\] core.pdc.row_out_n\[12\] core.pdc.row_out_n\[11\]
+ core.pdc.row_out_n\[10\] core.pdc.row_out_n\[9\] net52 core.pdc.row_out_n\[7\] core.pdc.row_out_n\[6\]
+ core.pdc.row_out_n\[5\] core.pdc.row_out_n\[4\] core.pdc.row_out_n\[3\] core.pdc.row_out_n\[2\]
+ core.pdc.row_out_n\[1\] net84 net103 core.pdc.row_out_n\[15\] core.pdc.row_out_n\[14\]
+ core.pdc.row_out_n\[13\] core.pdc.row_out_n\[12\] core.pdc.row_out_n\[11\] core.pdc.row_out_n\[10\]
+ core.pdc.row_out_n\[9\] core.cnb.nswitch_out\[11\] core.pdc.row_out_n\[7\] core.pdc.row_out_n\[6\]
+ core.pdc.row_out_n\[5\] core.pdc.row_out_n\[4\] core.pdc.row_out_n\[3\] core.pdc.row_out_n\[2\]
+ core.pdc.row_out_n\[1\] core.pdc.col_out_n\[31\] core.pdc.col_out_n\[30\] core.pdc.col_out_n\[29\]
+ core.pdc.col_out_n\[28\] core.pdc.col_out_n\[27\] core.pdc.col_out_n\[26\] core.pdc.col_out_n\[25\]
+ core.pdc.col_out_n\[24\] core.pdc.col_out_n\[23\] core.pdc.col_out_n\[22\] core.pdc.col_out_n\[21\]
+ core.pdc.col_out_n\[20\] core.pdc.col_out_n\[19\] core.pdc.col_out_n\[18\] core.pdc.col_out_n\[17\]
+ core.pdc.col_out_n\[16\] core.pdc.col_out_n\[15\] core.pdc.col_out_n\[14\] core.pdc.col_out_n\[13\]
+ core.pdc.col_out_n\[12\] core.pdc.col_out_n\[11\] core.pdc.col_out_n\[10\] core.pdc.col_out_n\[9\]
+ core.pdc.col_out_n\[8\] core.pdc.col_out_n\[7\] core.pdc.col_out_n\[6\] core.pdc.col_out_n\[5\]
+ core.pdc.col_out_n\[4\] core.pdc.col_out_n\[3\] core.pdc.col_out_n\[2\] core.pdc.col_out_n\[1\]
+ core.pdc.col_out_n\[0\] core.cnb.nswitch_out\[2\] core.cnb.nswitch_out\[1\] core.cnb.nswitch_out\[0\]
+ net102 core.cnb.is_sampling_w core.cnb.enable_loop_out inp_analog ctop_pmatrix_analog
+ VSS VDD adc_array_matrix_12bit
X_0857_ VSS VDD _0252_ _0283_ core.cnb.shift_register_r\[10\] VSS VDD sky130_fd_sc_hd__xnor2_1
XANTENNA__1039__A _0394_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_136_29 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_0788_ VSS VDD _0214_ core.osr.osr_mode_r\[0\] core.osr.sample_count_r\[4\] _0215_
+ VSS VDD sky130_fd_sc_hd__o21ai_1
X_1409_ _0751_ core.osr.next_result_w\[19\] _0736_ VSS VDD VSS VDD sky130_fd_sc_hd__nor2_1
XFILLER_83_242 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_45_15 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1502__A core.ndc.row_out_n\[4\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XPHY_304 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_315 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_61_14 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XPHY_326 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_337 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_348 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_359 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_101_65 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_40_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_126_40 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_34_128 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_34_117 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_35_92 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_31_879 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_1760_ net50 net66 _0023_ net54 VSS VDD VSS VDD sky130_fd_sc_hd__dfrtp_1
X_1691_ VSS VDD _0039_ _0197_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_98_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_111_122 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_1125_ VSS VDD core.pdc.col_out_n\[22\] _0528_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XANTENNA__1322__A _0651_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1056_ _0463_ _0477_ VDD VSS VSS VDD sky130_fd_sc_hd__inv_2
XANTENNA_cgen_dlycontrol4_in[4] net6 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_22_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_0909_ _0335_ _0334_ _0307_ VSS VDD VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_103_9 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xoutput39 VDD VSS result_out[12] net39 VSS VDD sky130_fd_sc_hd__buf_2
XANTENNA__1535__B1 net52 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_89_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_112_42 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_134 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_123 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_112 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_101 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_156 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_145 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_167 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_13_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XPHY_189 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_178 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_97_21 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_97_76 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_47_264 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XPHY_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_46_80 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_50_407 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1812_ core.osr.sample_count_r\[7\] net72 core.osr.next_sample_count_w\[7\] net58
+ VSS VDD VSS VDD sky130_fd_sc_hd__dfrtp_2
X_1743_ core.cnb.result_out\[3\] net68 _0006_ net81 VSS VDD VSS VDD sky130_fd_sc_hd__dfrtp_4
X_1674_ _0115_ _0189_ _0112_ core.osr.next_result_w\[13\] _0190_ VSS VDD VSS VDD sky130_fd_sc_hd__a31o_1
XANTENNA__1517__B1 net52 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_85_315 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1108_ VSS VDD _0520_ _0454_ _0453_ _0455_ VSS VDD sky130_fd_sc_hd__and3_1
XANTENNA__1804__CLK net77 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_53_267 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_53_289 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1039_ _0462_ _0394_ VSS VDD VSS VDD sky130_fd_sc_hd__clkbuf_4
XFILLER_88_131 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_67_57 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_88_175 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_107_86 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_88_197 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_84_370 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xpmat_103 pmat_103/LO net103 VDD VSS VSS VDD sky130_fd_sc_hd__conb_1
XFILLER_59_8 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_1390_ VSS VDD _0737_ _0738_ core.osr.result_r\[14\] VSS VDD sky130_fd_sc_hd__xnor2_1
XFILLER_50_226 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1726_ core.cnb.data_register_r\[11\] net64 core.cnb.next_data_register_w\[11\] net78
+ VSS VDD VSS VDD sky130_fd_sc_hd__dfrtp_1
X_1657_ _0133_ net40 _0175_ _0103_ VSS VDD VSS VDD sky130_fd_sc_hd__and3b_1
X_1588_ VDD VSS _0117_ _0104_ net44 VSS VDD sky130_fd_sc_hd__and2_1
XANTENNA_pmat_row_n[8] net52 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_139_125 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_5_105 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_118_74 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_118_85 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_49_304 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_49_315 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_89_473 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_49_337 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_49_348 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_94_33 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_91_104 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_94_66 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_27_93 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1777__D core.osr.next_result_w\[9\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_43_92 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_0890_ _0237_ _0245_ _0316_ _0242_ _0259_ VSS VDD VSS VDD sky130_fd_sc_hd__o22ai_1
XANTENNA__1196__A1 core.cnb.data_register_r\[0\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1511_ _0080_ _0352_ _0607_ VSS VDD VSS VDD sky130_fd_sc_hd__or2_4
X_1442_ _0471_ _0770_ _0502_ VSS VDD VSS VDD sky130_fd_sc_hd__or2_1
XFILLER_4_53 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_4_97 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1373_ VSS VDD _0724_ _0721_ core.osr.result_r\[11\] _0722_ VSS VDD sky130_fd_sc_hd__and3_1
XFILLER_55_318 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1330__A core.cnb.result_out\[6\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_139_29 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1709_ VSS VDD _0048_ _0206_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_133_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_48_59 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_46_329 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_104_54 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_64_14 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0782__C net10 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_80_24 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xfanout63 net63 net74 VSS VDD VSS VDD sky130_fd_sc_hd__clkbuf_4
Xfanout74 net74 net33 VSS VDD VSS VDD sky130_fd_sc_hd__clkbuf_4
Xfanout52 VDD VSS net52 core.cnb.nswitch_out\[11\] VSS VDD sky130_fd_sc_hd__buf_4
XFILLER_89_99 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_124_879 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_89_281 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1102__A1 _0450_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_0942_ _0295_ _0280_ _0290_ _0368_ _0367_ VDD VSS VSS VDD sky130_fd_sc_hd__or4b_1
X_0873_ core.cnb.shift_register_r\[12\] _0255_ _0252_ _0299_ _0254_ VDD VSS VSS VDD
+ sky130_fd_sc_hd__or4b_1
XFILLER_115_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1425_ core.osr.next_sample_count_w\[5\] _0760_ _0236_ _0761_ VSS VDD VSS VDD sky130_fd_sc_hd__o21a_1
XANTENNA__1325__A core.cnb.result_out\[6\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1356_ _0709_ _0708_ core.cnb.result_out\[9\] VSS VDD VSS VDD sky130_fd_sc_hd__xor2_4
XANTENNA__1044__B _0420_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_55_137 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_1287_ VSS VDD _0646_ core.osr.next_result_w\[2\] _0640_ VSS VDD sky130_fd_sc_hd__xnor2_1
XPHY_508 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1060__A _0347_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_51_310 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_519 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_50_16 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__0907__A1 core.cnb.data_register_r\[5\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_106_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1332__A1 core.cnb.result_out\[6\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_115_97 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_75_57 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_131_41 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_91_45 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1571__A1 core.cnb.result_out\[11\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1145__A core.cnb.nswitch_out\[0\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1210_ _0589_ _0590_ _0364_ VDD VSS VSS VDD sky130_fd_sc_hd__xor2_1
XFILLER_37_104 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1141_ _0423_ core.pdc.col_out_n\[31\] _0450_ VSS VDD VSS VDD sky130_fd_sc_hd__nor2_1
X_1072_ _0345_ _0493_ _0478_ _0444_ VDD VSS VSS VDD sky130_fd_sc_hd__or3_1
XFILLER_52_118 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_0925_ VDD VSS _0351_ _0350_ _0346_ VSS VDD sky130_fd_sc_hd__and2_1
X_0856_ _0240_ _0282_ _0239_ VSS VDD VSS VDD sky130_fd_sc_hd__nor2_2
X_0787_ VDD VSS _0214_ core.osr.osr_mode_r\[2\] VSS VDD sky130_fd_sc_hd__buf_2
X_1408_ VSS VDD _0750_ _0751_ core.osr.result_r\[19\] VSS VDD sky130_fd_sc_hd__xnor2_1
XANTENNA__1055__A _0427_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_28_104 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_1339_ core.osr.result_r\[8\] _0693_ VDD VSS VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_43_118 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1502__B _0074_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XPHY_305 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_316 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_51_151 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_327 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_338 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_349 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1250__B1 _0616_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_10_41 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_105_120 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_126_52 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_10_85 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_126_85 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_47_402 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_47_413 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_47_468 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_89_8 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_1690_ VSS VDD _0616_ core.cnb.shift_register_r\[9\] core.cnb.shift_register_r\[8\]
+ _0197_ VSS VDD sky130_fd_sc_hd__mux2_1
X_1124_ _0526_ _0528_ _0527_ VSS VDD VSS VDD sky130_fd_sc_hd__or2_1
XFILLER_25_129 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_1055_ _0427_ _0476_ _0475_ VSS VDD VSS VDD sky130_fd_sc_hd__or2_1
XFILLER_53_416 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_53_449 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA_cgen_dlycontrol4_in[3] net5 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_0908_ _0334_ _0291_ _0239_ _0294_ _0243_ _0312_ VDD VSS VSS VDD sky130_fd_sc_hd__o32a_1
X_0839_ _0259_ _0258_ _0264_ _0265_ VDD VSS VSS VDD sky130_fd_sc_hd__a21o_1
XFILLER_88_313 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_88_324 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_102_101 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1535__A1 _0079_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XPHY_124 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_113 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_102 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_52_460 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_157 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_135 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1471__B1 _0471_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XPHY_146 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_168 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_179 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_137_51 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_46_70 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_4 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_1811_ core.osr.sample_count_r\[6\] net72 core.osr.next_sample_count_w\[6\] net58
+ VSS VDD VSS VDD sky130_fd_sc_hd__dfrtp_2
X_1742_ core.cnb.result_out\[2\] net68 _0005_ net81 VSS VDD VSS VDD sky130_fd_sc_hd__dfrtp_1
X_1673_ core.cnb.result_out\[11\] _0209_ _0189_ net42 _0236_ VDD VSS VSS VDD sky130_fd_sc_hd__a22o_1
XANTENNA__1517__A1 _0079_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1317__B _0212_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_53_257 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_1107_ _0374_ _0462_ _0468_ _0519_ VSS VDD VSS VDD sky130_fd_sc_hd__o21a_2
X_1038_ VSS VDD core.pdc.col_out_n\[2\] _0461_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XANTENNA__1508__A core.ndc.row_out_n\[4\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_107_21 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_67_69 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1243__A _0614_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1770__RESET_B net67 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_cgen_dlycontrol3_in[4] net22 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_50_238 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_92_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_1725_ core.cnb.data_register_r\[10\] net63 core.cnb.next_data_register_w\[10\] net80
+ VSS VDD VSS VDD sky130_fd_sc_hd__dfrtp_4
XANTENNA_pmat_col_n[21] core.pdc.col_out_n\[21\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1656_ VSS VDD _0027_ _0132_ _0170_ core.cnb.result_out\[8\] _0174_ VSS VDD sky130_fd_sc_hd__a211o_1
X_1587_ VSS VDD _0016_ _0116_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_37_28 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_37_39 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_118_64 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_78_46 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_134_52 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_134_41 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_134_85 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_27_50 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA_input12_A config_1_in[5] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_71_8 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_1510_ VDD VSS _0079_ _0073_ VSS VDD sky130_fd_sc_hd__buf_6
X_1441_ _0529_ _0532_ core.ndc.col_out_n\[4\] _0422_ VDD VSS VSS VDD sky130_fd_sc_hd__a21oi_1
XFILLER_4_65 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1372_ _0721_ core.osr.result_r\[11\] _0723_ _0722_ VDD VSS VSS VDD sky130_fd_sc_hd__a21oi_1
XANTENNA__1353__C1 _0634_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_82_149 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_136_129 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1058__A _0345_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_2_109 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1708_ VSS VDD _0736_ net10 _0110_ _0206_ VSS VDD sky130_fd_sc_hd__mux2_1
XANTENNA__0897__A core.cnb.data_register_r\[5\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1639_ core.cnb.result_out\[5\] _0132_ _0161_ net51 _0236_ VDD VSS VSS VDD sky130_fd_sc_hd__a22o_1
XANTENNA_input4_A config_1_in[12] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_86_477 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_104_99 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_120_10 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xfanout53 net53 core.cnb.enable_loop_out VSS VDD VSS VDD sky130_fd_sc_hd__clkbuf_4
Xfanout64 net64 net67 VSS VDD VSS VDD sky130_fd_sc_hd__clkbuf_4
Xfanout75 VDD VSS net75 net76 VSS VDD sky130_fd_sc_hd__buf_2
XFILLER_13_30 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_129_30 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_89_78 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_49_113 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_89_260 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_92_425 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1102__A2 _0514_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_54_92 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_61_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_0941_ _0275_ _0270_ core.cnb.data_register_r\[2\] _0367_ VDD VSS VSS VDD sky130_fd_sc_hd__a21o_1
X_0872_ _0281_ _0298_ _0296_ _0297_ VSS VDD VSS VDD sky130_fd_sc_hd__nand3_2
XFILLER_70_80 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_118_118 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_1424_ VSS VDD _0761_ _0759_ core.osr.sample_count_r\[4\] _0757_ VSS VDD sky130_fd_sc_hd__and3_1
X_1355_ _0707_ _0708_ _0703_ VSS VDD VSS VDD sky130_fd_sc_hd__nor2_2
XANTENNA__1802__RESET_B net63 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_55_105 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_83_403 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_83_436 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1286_ VSS VDD _0646_ _0644_ _0635_ _0645_ VSS VDD sky130_fd_sc_hd__and3_1
XANTENNA__0883__C core.cnb.shift_register_r\[1\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XPHY_509 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_51_355 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_52_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_50_39 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_109_107 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_109_118 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1516__A core.pdc.row_out_n\[9\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_1_8 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_59_48 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_115_87 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_fanout62_A net74 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_131_53 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_131_64 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_43_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_91_57 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xcomp VDD clk_comp_cgen ctop_pmatrix_analog ctop_nmatrix_analog decision_finish_comp_n
+ comp/latch_qn core.cnb.comparator_in VSS adc_comp_latch
X_1140_ _0354_ core.ndc.col_out_n\[31\] core.pdc.col_out_n\[30\] _0534_ VDD VSS VSS
+ VDD sky130_fd_sc_hd__a21oi_1
X_1071_ _0347_ _0492_ _0478_ _0444_ VDD VSS VSS VDD sky130_fd_sc_hd__or3_1
XFILLER_92_266 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_34_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_0924_ _0347_ _0348_ _0350_ _0349_ VSS VDD VSS VDD sky130_fd_sc_hd__or3_2
X_0855_ core.cnb.data_register_r\[1\] _0276_ _0280_ _0281_ VDD VSS VSS VDD sky130_fd_sc_hd__or3b_2
X_0786_ VDD VSS _0213_ core.osr.osr_mode_r\[1\] VSS VDD sky130_fd_sc_hd__buf_2
XANTENNA__1336__A core.cnb.result_out\[7\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_114_121 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_29_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_1407_ VSS VDD _0750_ _0729_ core.osr.result_r\[18\] _0747_ VSS VDD sky130_fd_sc_hd__and3_1
X_1338_ _0692_ core.cnb.result_out\[8\] VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_2
X_1269_ core.cnb.average_sum_r\[3\] _0631_ _0632_ _0629_ VDD VSS VSS VDD sky130_fd_sc_hd__a21oi_1
XANTENNA__1071__A _0347_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_83_266 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_45_39 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1078__B2 _0450_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_25_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_51_130 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_306 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_51_163 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_317 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_328 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_339 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_51_196 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_10_53 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_10_97 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1724__RESET_B net63 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_126_97 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1680__S _0568_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_19_84 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_16_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_35_83 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__0995__A _0394_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1123_ _0463_ _0524_ _0352_ _0497_ _0527_ VSS VDD VSS VDD sky130_fd_sc_hd__a31o_1
X_1054_ _0475_ _0454_ _0453_ _0455_ VSS VDD VSS VDD sky130_fd_sc_hd__o21a_1
XANTENNA_cgen_dlycontrol4_in[2] net4 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_0907_ _0333_ core.cnb.data_register_r\[4\] _0329_ core.cnb.data_register_r\[5\]
+ _0331_ _0332_ VDD VSS VSS VDD sky130_fd_sc_hd__o311a_2
X_0838_ VDD VSS _0264_ _0263_ VSS VDD sky130_fd_sc_hd__buf_6
XANTENNA__1535__A2 _0080_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_88_336 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_72_15 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_112_66 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_125 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_114 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_103 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_72_37 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XPHY_136 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1471__A1 _0450_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_52_472 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_147 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_158 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_169 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_122_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XPHY_5 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1462__A1 _0449_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1810_ core.osr.sample_count_r\[5\] net71 core.osr.next_sample_count_w\[5\] net57
+ VSS VDD VSS VDD sky130_fd_sc_hd__dfrtp_1
X_1741_ core.cnb.result_out\[1\] net65 _0004_ net78 VSS VDD VSS VDD sky130_fd_sc_hd__dfrtp_2
X_1672_ _0111_ _0188_ core.osr.next_result_w\[19\] VSS VDD VSS VDD sky130_fd_sc_hd__or2_1
XANTENNA__1517__A2 _0080_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_85_306 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1106_ _0518_ core.pdc.col_out_n\[13\] _0517_ VSS VDD VSS VDD sky130_fd_sc_hd__nor2_1
XFILLER_53_247 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1037_ VDD VSS _0461_ _0460_ _0459_ VSS VDD sky130_fd_sc_hd__and2_1
XFILLER_21_122 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1508__B _0077_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_107_11 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_91_309 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_83_47 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1380__B1 _0212_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_82_309 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_50_206 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_90_375 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1199__A0 core.cnb.nswitch_out\[1\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1724_ core.cnb.data_register_r\[9\] net63 core.cnb.next_data_register_w\[9\] net78
+ VSS VDD VSS VDD sky130_fd_sc_hd__dfrtp_4
X_1655_ core.osr.next_result_w\[14\] _0174_ _0172_ _0173_ _0230_ _0214_ VSS VDD VSS
+ VDD sky130_fd_sc_hd__o221a_1
X_1586_ VSS VDD _0115_ _0114_ _0109_ _0116_ VSS VDD sky130_fd_sc_hd__mux2_1
XANTENNA_pmat_row_n[6] core.pdc.row_out_n\[6\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_85_169 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1519__A core.pdc.row_out_n\[6\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_136_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_78_25 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_78_58 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_78_69 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_49_328 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_134_64 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_94_13 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_134_97 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_127_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_64_8 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1440_ _0529_ _0464_ core.ndc.col_out_n\[3\] _0460_ VDD VSS VSS VDD sky130_fd_sc_hd__a21oi_1
XFILLER_4_77 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_1371_ _0713_ core.osr.result_r\[10\] core.cnb.result_out\[10\] _0716_ _0722_ VSS
+ VDD VSS VDD sky130_fd_sc_hd__a31o_1
XFILLER_48_350 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_55_309 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1656__A1 core.cnb.result_out\[8\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_84_90 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_118_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1707_ VSS VDD _0047_ _0205_ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_1638_ core.osr.next_result_w\[7\] _0160_ core.osr.next_result_w\[13\] _0123_ _0124_
+ VSS VDD VSS VDD sky130_fd_sc_hd__o22a_1
XANTENNA__1074__A _0347_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1569_ VSS VDD _0101_ _0610_ _0100_ _0013_ core.cnb.result_out\[10\] VSS VDD sky130_fd_sc_hd__a2bb2o_1
XANTENNA__1344__B1 _0212_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1769__CLK net55 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_46_309 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_54_353 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_54_386 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_54_397 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xfanout65 net67 net65 VSS VDD VSS VDD sky130_fd_sc_hd__clkbuf_2
Xfanout54 VDD VSS net54 net55 VSS VDD sky130_fd_sc_hd__buf_2
Xfanout76 VDD VSS net76 net77 VSS VDD sky130_fd_sc_hd__buf_2
XFILLER_129_75 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_129_64 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_109_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_89_250 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_89_272 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_49_125 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_92_404 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_61_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_0940_ _0366_ _0365_ _0364_ VSS VDD VSS VDD sky130_fd_sc_hd__xor2_4
X_0871_ _0295_ _0276_ _0297_ _0290_ _0280_ VDD VSS VSS VDD sky130_fd_sc_hd__or4b_2
XANTENNA__0998__A _0354_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1423_ core.osr.sample_count_r\[4\] _0759_ _0760_ _0757_ VDD VSS VSS VDD sky130_fd_sc_hd__a21oi_1
XFILLER_48_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_1354_ core.osr.result_r\[9\] _0635_ _0707_ _0705_ _0706_ _0704_ VSS VDD VSS VDD
+ sky130_fd_sc_hd__a311o_1
X_1285_ _0645_ _0643_ core.osr.result_r\[2\] VSS VDD VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_55_128 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0883__D core.cnb.is_sampling_w VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_52_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_50_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1565__A0 core.cnb.result_out\[9\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_119_9 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_115_66 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_75_48 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1532__A core.ndc.row_out_n\[12\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_fanout55_A net56 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_131_76 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_43_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1678__S _0568_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_24_41 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_91_69 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_49_93 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1442__A _0471_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1070_ _0491_ _0490_ _0489_ _0487_ _0486_ _0433_ VDD VSS VSS VDD sky130_fd_sc_hd__o2111a_1
XFILLER_34_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_0923_ _0333_ _0336_ _0306_ _0341_ _0349_ VSS VDD VSS VDD sky130_fd_sc_hd__o211ai_4
X_0854_ _0258_ _0280_ _0278_ _0264_ _0279_ VSS VDD VSS VDD sky130_fd_sc_hd__o22a_1
X_0785_ _0209_ _0210_ _0211_ core.osr.sample_count_r\[0\] _0212_ VSS VDD VSS VDD sky130_fd_sc_hd__a31o_4
X_1406_ _0749_ core.osr.next_result_w\[18\] _0736_ VSS VDD VSS VDD sky130_fd_sc_hd__nor2_1
X_1337_ _0691_ core.osr.next_result_w\[7\] VDD VSS VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_45_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_1268_ core.cnb.average_sum_r\[4\] _0631_ VDD VSS VSS VDD sky130_fd_sc_hd__inv_2
X_1199_ VSS VDD _0579_ core.cnb.data_register_r\[1\] core.cnb.nswitch_out\[1\] _0582_
+ VSS VDD sky130_fd_sc_hd__mux2_1
XPHY_307 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_25_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XPHY_318 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_329 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_101_57 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_51_175 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1235__C1 _0586_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1527__A core.pdc.row_out_n\[2\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_105_100 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_10_65 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_126_76 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1262__A core.cnb.comparator_in VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_19_96 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_16_879 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1437__A _0768_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__0995__B _0410_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1172__A core.cnb.is_sampling_w VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1122_ _0500_ _0526_ _0499_ VSS VDD VSS VDD sky130_fd_sc_hd__nor2_1
X_1053_ VDD VSS _0474_ _0462_ VSS VDD sky130_fd_sc_hd__buf_2
XFILLER_46_470 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_46_481 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA_cgen_dlycontrol4_in[1] net3 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_0906_ _0318_ core.cnb.data_register_r\[4\] _0332_ _0330_ _0329_ VDD VSS VSS VDD
+ sky130_fd_sc_hd__or4_1
X_0837_ _0239_ _0261_ _0263_ _0262_ _0240_ VDD VSS VSS VDD sky130_fd_sc_hd__or4_1
XFILLER_88_348 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_88_359 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_16_109 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_115 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_104 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_148 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_137 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_126 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_159 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_21_64 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__0982__A1 _0364_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_115_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__0982__B2 core.cnb.data_register_r\[5\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_97_57 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_97_68 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_46_61 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_6 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1462__A2 _0512_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_62_60 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1740_ core.cnb.result_out\[0\] net64 _0003_ net78 VSS VDD VSS VDD sky130_fd_sc_hd__dfrtp_2
X_1671_ VSS VDD _0187_ core.osr.next_result_w\[17\] _0186_ _0110_ _0232_ VSS VDD sky130_fd_sc_hd__a211o_1
X_1105_ _0374_ _0474_ _0518_ _0472_ VDD VSS VSS VDD sky130_fd_sc_hd__a21oi_1
X_1036_ _0455_ _0460_ _0422_ VDD VSS VSS VDD sky130_fd_sc_hd__or2_2
XFILLER_21_101 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_88_101 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_12_123 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1686__S _0616_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_32_96 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_5_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_94_104 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_94_115 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1450__A _0529_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XPHY_490 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1199__A1 core.cnb.data_register_r\[1\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1723_ core.cnb.data_register_r\[8\] net63 core.cnb.next_data_register_w\[8\] net80
+ VSS VDD VSS VDD sky130_fd_sc_hd__dfrtp_4
X_1654_ _0173_ core.osr.next_result_w\[16\] _0134_ _0124_ VSS VDD VSS VDD sky130_fd_sc_hd__o21a_1
X_1585_ VDD VSS _0115_ _0235_ VSS VDD sky130_fd_sc_hd__buf_2
XANTENNA__1371__A1 core.cnb.result_out\[10\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1123__A1 _0352_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1659__C1 _0235_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1019_ _0444_ _0331_ _0377_ VSS VDD VSS VDD sky130_fd_sc_hd__nand2_2
XFILLER_118_33 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_136_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_78_37 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1362__B2 core.cnb.result_out\[8\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1362__A1 core.cnb.result_out\[7\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1114__A1 _0353_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_43_40 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_127_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1370_ _0716_ _0713_ core.cnb.result_out\[10\] _0721_ VDD VSS VSS VDD sky130_fd_sc_hd__a21o_1
XFILLER_68_70 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1105__A1 _0374_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_48_384 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_136_109 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1706_ VSS VDD _0614_ _0588_ core.cnb.shift_register_r\[16\] _0205_ VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_118_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1637_ _0159_ _0158_ _0111_ VSS VDD VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_48_18 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_48_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_1568_ _0101_ _0568_ core.cnb.shift_register_r\[2\] VSS VDD VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_86_402 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1499_ VDD VSS _0073_ _0072_ VSS VDD sky130_fd_sc_hd__buf_6
XANTENNA__1090__A _0427_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_54_321 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_54_365 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1789__RESET_B net63 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xfanout55 VDD VSS net55 net56 VSS VDD sky130_fd_sc_hd__buf_2
Xfanout77 core.clk_dig_in net77 VSS VDD VSS VDD sky130_fd_sc_hd__clkbuf_2
XANTENNA__1718__RESET_B net74 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xfanout66 net66 net67 VSS VDD VSS VDD sky130_fd_sc_hd__clkbuf_4
XFILLER_127_109 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_129_98 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_109_879 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_89_69 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_8_3 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_38_95 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1099__B1 _0513_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1638__A2 core.osr.next_result_w\[7\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1271__B1 _0615_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_0870_ core.cnb.data_register_r\[1\] _0290_ _0296_ _0295_ VSS VDD VSS VDD sky130_fd_sc_hd__or3_2
XFILLER_118_109 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0998__B _0423_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1422_ core.osr.sample_count_r\[5\] _0759_ VDD VSS VSS VDD sky130_fd_sc_hd__inv_2
X_1353_ _0706_ _0682_ _0634_ core.osr.result_r\[9\] _0692_ _0693_ VDD VSS VSS VDD
+ sky130_fd_sc_hd__o2111a_1
X_1284_ core.osr.result_r\[2\] _0644_ _0643_ VSS VDD VSS VDD sky130_fd_sc_hd__or2_1
XFILLER_83_449 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_51_324 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_51_346 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_0999_ VDD VSS _0424_ _0353_ VSS VDD sky130_fd_sc_hd__buf_4
XANTENNA__1736__CLK net76 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1085__A _0466_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_59_17 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_59_39 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_115_12 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_86_265 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_131_88 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1694__S _0614_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_49_72 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_1_57 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_0922_ _0327_ _0326_ _0298_ _0267_ _0348_ VDD VSS VSS VDD sky130_fd_sc_hd__o211a_2
XANTENNA__1759__CLK net55 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_0853_ _0239_ _0279_ _0240_ VSS VDD VSS VDD sky130_fd_sc_hd__or2_1
XFILLER_60_3 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_0784_ core.osr.sample_count_r\[6\] core.osr.sample_count_r\[8\] _0211_ core.osr.sample_count_r\[2\]
+ core.osr.sample_count_r\[4\] VSS VDD VSS VDD sky130_fd_sc_hd__nor4_2
X_1405_ _0748_ _0749_ core.osr.result_r\[18\] VDD VSS VSS VDD sky130_fd_sc_hd__xor2_1
X_1336_ VSS VDD _0691_ core.cnb.result_out\[7\] _0690_ VSS VDD sky130_fd_sc_hd__xnor2_2
XFILLER_28_118 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xinput1 VSS VDD net1 config_1_in[0] VSS VDD sky130_fd_sc_hd__clkbuf_1
XANTENNA__1352__B _0634_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1267_ _0630_ core.cnb.next_average_sum_w\[3\] _0616_ VSS VDD VSS VDD sky130_fd_sc_hd__nor2_1
X_1198_ VSS VDD core.cnb.next_data_register_w\[0\] _0581_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XPHY_308 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_319 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_10_77 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_19_118 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_19_107 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1710__A1 net11 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_47_449 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_35_30 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1474__B1 _0465_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1453__A _0512_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__0995__C _0420_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_76_70 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1121_ core.pdc.col_out_n\[21\] _0354_ _0511_ _0525_ VSS VDD VSS VDD sky130_fd_sc_hd__o21a_1
XFILLER_53_408 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1052_ VSS VDD _0471_ _0424_ _0473_ core.pdc.col_out_n\[4\] VSS VDD sky130_fd_sc_hd__o21ai_1
XANTENNA_cgen_dlycontrol4_in[0] net2 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_33_121 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_0905_ core.cnb.data_register_r\[5\] _0330_ _0331_ _0318_ VSS VDD VSS VDD sky130_fd_sc_hd__or3_2
X_0836_ core.cnb.shift_register_r\[9\] _0262_ core.cnb.shift_register_r\[8\] core.cnb.shift_register_r\[16\]
+ VDD VSS VSS VDD sky130_fd_sc_hd__or3_1
XFILLER_102_126 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_56_29 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1319_ _0674_ core.osr.result_r\[4\] _0665_ core.cnb.result_out\[4\] _0664_ VSS VDD
+ VSS VDD sky130_fd_sc_hd__o31a_1
XPHY_116 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_105 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_149 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_138 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_127 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1538__A core.ndc.row_out_n\[4\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1257__B _0615_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_108_3 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1273__A _0634_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_87_360 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_input28_A config_2_in[5] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_46_95 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_7 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1212__S _0586_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_30_102 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1670_ _0740_ _0186_ _0110_ _0736_ VSS VDD VSS VDD sky130_fd_sc_hd__nor3_1
XFILLER_97_113 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_87_80 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_1104_ _0516_ _0517_ _0427_ VSS VDD VSS VDD sky130_fd_sc_hd__nor2_1
X_1035_ _0446_ _0427_ _0432_ _0458_ _0459_ VSS VDD VSS VDD sky130_fd_sc_hd__a31o_1
XFILLER_21_113 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_0819_ core.cnb.shift_register_r\[11\] core.cnb.shift_register_r\[9\] _0245_ core.cnb.shift_register_r\[8\]
+ core.cnb.shift_register_r\[10\] VDD VSS VSS VDD sky130_fd_sc_hd__or4_1
X_1799_ core.cnb.shift_register_r\[11\] net63 _0042_ net77 VSS VDD VSS VDD sky130_fd_sc_hd__dfrtp_2
XFILLER_88_113 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_107_57 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1093__A _0427_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_67_28 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_88_157 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1677__B1 _0089_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_84_396 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_16_65 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_5_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_57_50 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_57_83 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_90_300 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_91_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_90_388 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_480 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_491 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_1722_ core.cnb.data_register_r\[7\] net68 core.cnb.next_data_register_w\[7\] net81
+ VSS VDD VSS VDD sky130_fd_sc_hd__dfrtp_4
X_1653_ _0143_ _0172_ _0171_ core.osr.next_result_w\[12\] core.osr.next_result_w\[10\]
+ VSS VDD VSS VDD sky130_fd_sc_hd__o22a_1
XANTENNA__0810__A _0236_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1584_ _0114_ core.osr.next_result_w\[3\] _0113_ core.osr.next_result_w\[5\] _0110_
+ _0111_ VSS VDD VSS VDD sky130_fd_sc_hd__a32o_1
XFILLER_98_90 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_82_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1018_ VSS VDD _0442_ _0443_ _0345_ VSS VDD sky130_fd_sc_hd__xnor2_1
XFILLER_118_45 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_89_400 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1114__A2 _0519_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_84_182 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_73_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1792__CLK net76 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1105__A2 _0472_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_48_341 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_48_374 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_48_396 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0864__A1 core.cnb.data_register_r\[0\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_64_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_90_185 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_1705_ VSS VDD _0046_ _0204_ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_1636_ VSS VDD _0110_ _0726_ _0709_ _0158_ VSS VDD sky130_fd_sc_hd__mux2_1
X_1567_ _0100_ _0089_ net53 VSS VDD VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_86_414 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_1498_ _0063_ _0071_ _0062_ _0072_ _0064_ VDD VSS VSS VDD sky130_fd_sc_hd__or4b_1
XFILLER_86_425 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_54_300 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_55_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xfanout56 VDD VSS net56 core.cnb.conv_finished_r VSS VDD sky130_fd_sc_hd__buf_2
Xfanout78 VDD VSS net78 net79 VSS VDD sky130_fd_sc_hd__buf_2
Xfanout67 net67 net69 VSS VDD VSS VDD sky130_fd_sc_hd__clkbuf_4
XANTENNA__1032__A1 _0450_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_89_26 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_1_123 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_89_296 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1099__A1 _0424_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_92_417 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA_input10_A config_1_in[3] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_46_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_126_121 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_1421_ _0758_ core.osr.next_sample_count_w\[4\] core.osr.is_last_sample VSS VDD VSS
+ VDD sky130_fd_sc_hd__nor2_1
X_1352_ VSS VDD core.osr.result_r\[8\] core.osr.result_r\[9\] _0705_ core.cnb.result_out\[8\]
+ _0634_ VSS VDD sky130_fd_sc_hd__and4b_1
X_1283_ _0643_ _0642_ _0641_ VSS VDD VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_83_417 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_48_193 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_37_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_51_303 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_91_461 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1069__C _0373_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_0998_ _0423_ core.pdc.col_out_n\[0\] _0354_ VSS VDD VSS VDD sky130_fd_sc_hd__nor2_1
XANTENNA__1014__A1 _0328_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_59_29 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1619_ _0118_ _0144_ _0143_ _0213_ core.osr.next_result_w\[6\] VSS VDD VSS VDD sky130_fd_sc_hd__o22a_1
XANTENNA_input2_A config_1_in[10] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_115_57 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_28_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_54_141 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_54_174 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_91_27 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_24_21 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_138_3 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_123_124 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_123_113 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_1_14 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_49_84 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1215__S _0586_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_37_119 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_19_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_1_69 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_92_258 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_65_83 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_0921_ VSS VDD _0347_ core.cnb.data_register_r\[8\] _0344_ VSS VDD sky130_fd_sc_hd__xnor2_2
X_0852_ _0268_ _0278_ _0241_ _0277_ VDD VSS VSS VDD sky130_fd_sc_hd__or3_1
X_0783_ core.osr.sample_count_r\[1\] core.osr.sample_count_r\[5\] _0210_ core.osr.sample_count_r\[7\]
+ core.osr.sample_count_r\[3\] VSS VDD VSS VDD sky130_fd_sc_hd__nor4_4
XANTENNA_cgen_sample_p_in core.cnb.is_sampling_w VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1404_ _0748_ _0747_ _0729_ VSS VDD VSS VDD sky130_fd_sc_hd__nand2_1
X_1335_ _0682_ _0689_ _0690_ _0634_ VSS VDD VSS VDD sky130_fd_sc_hd__and3b_1
XANTENNA__0867__D_N core.cnb.data_register_r\[0\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xinput2 VDD VSS config_1_in[10] net2 VSS VDD sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_83_203 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_1266_ VSS VDD _0629_ _0630_ core.cnb.average_sum_r\[3\] VSS VDD sky130_fd_sc_hd__xnor2_1
X_1197_ VDD VSS _0581_ _0580_ net53 VSS VDD sky130_fd_sc_hd__and2_1
XFILLER_101_15 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_309 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_126_34 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_86_16 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_86_49 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_35_42 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1474__A1 _0450_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_25_7 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1120_ _0477_ _0499_ _0525_ _0497_ VDD VSS VSS VDD sky130_fd_sc_hd__a21oi_1
X_1051_ _0473_ _0472_ _0466_ VSS VDD VSS VDD sky130_fd_sc_hd__nand2_1
X_0904_ _0258_ _0330_ _0264_ VSS VDD VSS VDD sky130_fd_sc_hd__nor2_1
X_0835_ VDD VSS _0261_ _0260_ VSS VDD sky130_fd_sc_hd__buf_2
XANTENNA__1347__C _0212_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1318_ core.osr.next_result_w\[6\] _0673_ core.cnb.result_out\[6\] VSS VDD VSS VDD
+ sky130_fd_sc_hd__xnor2_4
X_1249_ core.cnb.average_counter_r\[2\] _0619_ _0557_ VSS VDD VSS VDD sky130_fd_sc_hd__or2_1
XFILLER_112_25 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_112_36 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_106 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_24_122 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_72_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XPHY_139 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_128 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_117 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_21_22 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1538__B _0074_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_21_33 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1447__A1 _0529_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XPHY_8 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_7_57 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA_pmat_en_bit_n[2] core.cnb.nswitch_out\[2\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_16_3 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1103_ _0516_ _0420_ _0462_ _0453_ _0455_ VSS VDD VSS VDD sky130_fd_sc_hd__o31a_1
XANTENNA__0808__A _0212_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1034_ VDD VSS _0458_ _0453_ _0394_ VSS VDD sky130_fd_sc_hd__and2_1
X_1798_ core.cnb.shift_register_r\[10\] net62 _0041_ net77 VSS VDD VSS VDD sky130_fd_sc_hd__dfrtp_4
X_0818_ core.cnb.shift_register_r\[1\] _0244_ core.cnb.is_sampling_w VSS VDD VSS VDD
+ sky130_fd_sc_hd__or2_1
XANTENNA__1374__A _0212_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_107_47 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_88_125 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_88_169 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1677__A1 core.cnb.shift_register_r\[1\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_123_57 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_16_11 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_16_77 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_52_261 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_52_283 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_139_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_120_3 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1668__A1 core.cnb.result_out\[10\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_87_191 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_91_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XPHY_470 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_492 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_481 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_1721_ core.cnb.data_register_r\[6\] net64 core.cnb.next_data_register_w\[6\] net79
+ VSS VDD VSS VDD sky130_fd_sc_hd__dfrtp_4
X_1652_ _0213_ _0171_ _0216_ VSS VDD VSS VDD sky130_fd_sc_hd__or2_1
XANTENNA__1194__A core.cnb.comparator_in VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1583_ _0111_ _0113_ _0112_ VSS VDD VSS VDD sky130_fd_sc_hd__nor2_1
XFILLER_85_106 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_85_117 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_85_139 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_82_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1017_ VSS VDD _0306_ _0333_ _0341_ _0442_ VSS VDD sky130_fd_sc_hd__o21ai_1
XANTENNA__1369__A core.cnb.result_out\[10\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_118_57 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_89_412 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_27_32 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_73_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_43_86 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_4_14 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1218__S _0586_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_64_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_90_120 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_83_3 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1704_ VSS VDD _0614_ core.cnb.shift_register_r\[16\] _0254_ _0204_ VSS VDD sky130_fd_sc_hd__mux2_1
X_1635_ _0156_ _0155_ _0157_ _0023_ VDD VSS VSS VDD sky130_fd_sc_hd__a21o_1
X_1566_ VSS VDD _0012_ _0099_ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_1497_ _0071_ _0343_ core.cnb.data_register_r\[10\] _0056_ _0065_ _0070_ VSS VDD
+ VSS VDD sky130_fd_sc_hd__o311a_1
XFILLER_86_437 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_104_37 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_54_345 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_55_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_120_25 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_120_36 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_120_47 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_120_69 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xfanout57 VDD VSS net57 core.cnb.conv_finished_r VSS VDD sky130_fd_sc_hd__buf_2
Xfanout79 VDD VSS net79 net80 VSS VDD sky130_fd_sc_hd__buf_2
Xfanout68 net68 net69 VSS VDD VSS VDD sky130_fd_sc_hd__clkbuf_4
XFILLER_1_113 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1099__A2 _0512_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_46_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_54_52 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_54_85 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_70_40 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1559__A0 core.cnb.result_out\[6\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_62_8 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1420_ VSS VDD _0757_ _0758_ core.osr.sample_count_r\[4\] VSS VDD sky130_fd_sc_hd__xnor2_1
XFILLER_79_82 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1351_ core.cnb.result_out\[8\] _0704_ core.osr.result_r\[8\] VSS VDD VSS VDD sky130_fd_sc_hd__nor2_1
X_1282_ core.cnb.result_out\[1\] core.osr.result_r\[1\] core.osr.result_r\[0\] _0642_
+ core.cnb.result_out\[0\] VSS VDD VSS VDD sky130_fd_sc_hd__o211ai_2
XFILLER_37_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_91_473 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_51_337 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_0997_ _0423_ _0376_ _0422_ VSS VDD VSS VDD sky130_fd_sc_hd__nor2_4
XANTENNA__1014__A2 _0342_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_117_122 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_1618_ _0143_ _0216_ _0213_ VSS VDD VSS VDD sky130_fd_sc_hd__nand2_1
X_1549_ VSS VDD _0089_ core.cnb.next_data_register_w\[1\] core.cnb.result_out\[1\]
+ _0091_ VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_115_36 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_75_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_28_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_91_39 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_50_381 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_40_76 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_40_98 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_1_26 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_19_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_0920_ _0342_ _0328_ _0345_ _0346_ VDD VSS VSS VDD sky130_fd_sc_hd__a21o_1
X_0851_ VSS VDD core.cnb.shift_register_r\[10\] _0277_ core.cnb.shift_register_r\[11\]
+ VSS VDD sky130_fd_sc_hd__xnor2_1
X_0782_ net12 net10 net11 _0209_ VSS VDD VSS VDD sky130_fd_sc_hd__nor3_4
XFILLER_46_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_1403_ _0747_ core.osr.result_r\[17\] core.osr.result_r\[12\] core.osr.result_r\[16\]
+ _0741_ VSS VDD VSS VDD sky130_fd_sc_hd__and4_1
X_1334_ VSS VDD _0689_ _0686_ _0684_ _0688_ VSS VDD sky130_fd_sc_hd__and3_1
X_1265_ VDD VSS _0629_ _0627_ core.cnb.average_sum_r\[2\] VSS VDD sky130_fd_sc_hd__and2_1
XANTENNA__1352__D core.cnb.result_out\[8\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xinput3 VDD VSS config_1_in[11] net3 VSS VDD sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_49_470 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1468__C1 _0353_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1196_ VSS VDD _0579_ core.cnb.data_register_r\[0\] core.cnb.nswitch_out\[0\] _0580_
+ VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_91_281 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_51_123 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_51_145 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_51_189 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_117_9 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA_fanout53_A core.cnb.enable_loop_out VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_55_462 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_82_281 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA_nmat_row_n[4] core.ndc.row_out_n\[4\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1050_ VDD VSS _0472_ _0454_ _0453_ VSS VDD sky130_fd_sc_hd__and2_1
X_0903_ _0304_ _0319_ _0329_ _0320_ _0289_ VDD VSS VSS VDD sky130_fd_sc_hd__a22o_1
X_0834_ core.cnb.shift_register_r\[11\] _0260_ core.cnb.shift_register_r\[10\] VSS
+ VDD VSS VDD sky130_fd_sc_hd__or2_1
XANTENNA__1197__A net53 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1317_ _0671_ _0212_ _0672_ _0673_ VDD VSS VSS VDD sky130_fd_sc_hd__or3b_2
X_1248_ _0618_ _0557_ core.cnb.average_counter_r\[2\] VSS VDD VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_24_101 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1456__A2 _0468_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XPHY_107 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_1179_ _0563_ _0558_ core.cnb.sampled_avg_control_r\[1\] VSS VDD VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_52_443 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_129 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_118 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__0967__A1 _0373_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1570__A _0588_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XPHY_9 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_7_14 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_7_69 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_8_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA_pmat_en_bit_n[1] core.cnb.nswitch_out\[1\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_97_104 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1135__A1 _0529_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1102_ _0514_ _0450_ _0515_ core.pdc.col_out_n\[12\] VDD VSS VSS VDD sky130_fd_sc_hd__a21o_1
XFILLER_53_207 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_1033_ _0457_ core.pdc.col_out_n\[1\] _0448_ _0424_ VSS VDD VSS VDD sky130_fd_sc_hd__o21ai_2
XFILLER_46_281 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_0817_ _0240_ core.cnb.shift_register_r\[16\] _0243_ _0239_ _0242_ VDD VSS VSS VDD
+ sky130_fd_sc_hd__or4_1
X_1797_ core.cnb.shift_register_r\[9\] net62 _0040_ net76 VSS VDD VSS VDD sky130_fd_sc_hd__dfrtp_2
XFILLER_123_25 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1677__A2 _0615_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_123_36 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_84_343 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_84_365 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_52_295 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_32_33 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_139_879 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1117__A1 _0353_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_input33_A rst_n VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_90_313 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_73_51 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_460 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_471 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_493 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_85_7 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XPHY_482 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_1720_ core.cnb.data_register_r\[5\] net64 core.cnb.next_data_register_w\[5\] net79
+ VSS VDD VSS VDD sky130_fd_sc_hd__dfrtp_4
X_1651_ _0134_ net39 _0170_ _0104_ VSS VDD VSS VDD sky130_fd_sc_hd__and3b_1
X_1582_ _0112_ _0213_ _0217_ VSS VDD VSS VDD sky130_fd_sc_hd__and2b_1
XANTENNA_pmat_row_n[2] core.pdc.row_out_n\[2\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1016_ _0440_ _0439_ _0436_ _0433_ _0437_ _0441_ VSS VDD VSS VDD sky130_fd_sc_hd__o2111ai_1
XFILLER_139_109 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1739__CLK net76 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_118_25 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_89_424 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_134_79 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_43_21 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_43_98 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_43_76 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1035__B1 _0427_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_68_40 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_48_332 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_48_365 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XPHY_290 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_1703_ VSS VDD _0045_ _0203_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XANTENNA__1329__A1 _0651_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1634_ core.cnb.result_out\[4\] _0132_ _0157_ net50 _0236_ VDD VSS VSS VDD sky130_fd_sc_hd__a22o_1
X_1565_ VSS VDD _0088_ core.cnb.next_data_register_w\[9\] core.cnb.result_out\[9\]
+ _0099_ VSS VDD sky130_fd_sc_hd__mux2_1
X_1496_ _0070_ _0068_ _0066_ _0067_ _0069_ VSS VDD VSS VDD sky130_fd_sc_hd__and4_1
XFILLER_86_449 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_104_49 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_54_335 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_54_379 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xfanout58 VDD VSS net59 net58 VSS VDD sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout69 VDD VSS net69 net74 VSS VDD sky130_fd_sc_hd__buf_2
XFILLER_129_24 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_13_57 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_38_65 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1256__B1 _0615_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_70_52 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_55_8 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1350_ _0703_ _0702_ _0701_ VSS VDD VSS VDD sky130_fd_sc_hd__nand2_1
X_1281_ _0641_ core.osr.result_r\[1\] core.cnb.result_out\[1\] VSS VDD VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_48_184 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_91_441 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_51_316 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_0996_ VDD VSS _0422_ _0421_ VSS VDD sky130_fd_sc_hd__buf_6
X_1617_ VSS VDD _0020_ _0142_ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_1548_ VSS VDD _0003_ _0090_ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_1479_ VSS VDD net35 _0054_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_115_48 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_54_110 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_54_132 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_54_154 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_82_463 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_40_11 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_6_3 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_49_42 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_1_38 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_92_216 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_92_249 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_65_52 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_65_74 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_81_51 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_0850_ VDD VSS _0276_ _0275_ _0270_ VSS VDD sky130_fd_sc_hd__and2_1
X_1402_ _0745_ _0736_ core.osr.next_result_w\[17\] _0746_ VDD VSS VSS VDD sky130_fd_sc_hd__a21oi_1
X_1333_ VSS VDD _0688_ _0687_ core.osr.result_r\[6\] core.cnb.result_out\[6\] core.osr.result_r\[7\]
+ VSS VDD sky130_fd_sc_hd__a31oi_1
X_1264_ _0628_ core.cnb.next_average_sum_w\[2\] _0616_ VSS VDD VSS VDD sky130_fd_sc_hd__nor2_1
Xinput4 VDD VSS config_1_in[12] net4 VSS VDD sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_83_216 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1195_ _0579_ _0578_ _0239_ _0576_ _0568_ VDD VSS VSS VDD sky130_fd_sc_hd__a31oi_4
XFILLER_91_260 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_51_113 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_0979_ VSS VDD _0405_ _0404_ _0360_ _0355_ _0357_ VSS VDD sky130_fd_sc_hd__a211o_1
XANTENNA__1377__B core.cnb.result_out\[11\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_120_107 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_19_34 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_19_78 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_55_430 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_55_441 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_35_11 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_82_260 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_35_77 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1568__A core.cnb.shift_register_r\[2\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_0902_ _0267_ _0326_ _0298_ _0327_ _0328_ VSS VDD VSS VDD sky130_fd_sc_hd__o211ai_4
X_0833_ core.cnb.shift_register_r\[14\] _0252_ _0259_ core.cnb.shift_register_r\[15\]
+ core.cnb.shift_register_r\[12\] VDD VSS VSS VDD sky130_fd_sc_hd__or4b_2
XANTENNA__1772__CLK net56 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1316_ core.osr.result_r\[6\] _0672_ _0668_ _0670_ VDD VSS VSS VDD sky130_fd_sc_hd__or3_1
X_1247_ _0617_ core.cnb.next_average_counter_w\[1\] _0616_ VSS VDD VSS VDD sky130_fd_sc_hd__nor2_1
X_1178_ core.cnb.sampled_avg_control_r\[1\] core.cnb.sampled_avg_control_r\[2\] _0562_
+ core.cnb.sampled_avg_control_r\[0\] VSS VDD VSS VDD sky130_fd_sc_hd__or3b_1
XPHY_119 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_108 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_52_466 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_52_477 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1388__A _0212_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1613__A0 core.osr.next_result_w\[5\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_21_13 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_21_46 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_21_79 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_137_57 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_47_205 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_55_260 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_15_124 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_15_113 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_55_271 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1298__A _0212_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_7_26 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_8_879 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA_pmat_en_bit_n[0] core.cnb.nswitch_out\[0\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1135__A2 _0465_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1101_ VDD VSS _0466_ _0515_ _0468_ VSS VDD sky130_fd_sc_hd__and2_2
XFILLER_94_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1032_ _0450_ _0456_ _0457_ _0452_ VDD VSS VSS VDD sky130_fd_sc_hd__a21oi_1
XFILLER_46_293 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1700__S _0614_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_0816_ VDD VSS _0242_ _0241_ VSS VDD sky130_fd_sc_hd__buf_2
X_1796_ core.cnb.shift_register_r\[8\] net61 _0039_ net76 VSS VDD VSS VDD sky130_fd_sc_hd__dfrtp_2
XFILLER_84_355 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_85_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_84_388 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_8_109 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_32_56 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_32_89 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_32_78 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_106_3 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_input26_A config_2_in[3] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_76_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XPHY_450 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_461 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_494 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_472 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_483 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_1650_ VSS VDD _0026_ _0132_ _0167_ core.cnb.result_out\[7\] _0169_ VSS VDD sky130_fd_sc_hd__a211o_1
X_1581_ VDD VSS _0111_ _0229_ VSS VDD sky130_fd_sc_hd__buf_2
XFILLER_98_60 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_67_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1015_ _0373_ _0348_ _0440_ _0349_ _0438_ VDD VSS VSS VDD sky130_fd_sc_hd__or4_1
X_1779_ core.osr.result_r\[11\] net67 core.osr.next_result_w\[11\] net54 VSS VDD VSS
+ VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_89_436 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_58_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_84_141 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_84_152 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_138_121 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_4_123 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_68_85 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_49_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XPHY_280 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_291 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_1702_ VSS VDD _0614_ _0254_ _0255_ _0203_ VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_69_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_1633_ core.osr.next_result_w\[6\] _0156_ core.osr.next_result_w\[10\] _0134_ _0123_
+ _0230_ VSS VDD VSS VDD sky130_fd_sc_hd__o221a_1
XANTENNA_cgen_nsample_n_in core.cnb.enable_loop_out VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1564_ VSS VDD _0011_ _0098_ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_1495_ core.cnb.data_register_r\[10\] _0343_ _0069_ _0552_ _0598_ VDD VSS VSS VDD
+ sky130_fd_sc_hd__or4_1
XFILLER_13_14 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xfanout59 VDD VSS net59 core.cnb.conv_finished_r VSS VDD sky130_fd_sc_hd__buf_2
XFILLER_13_36 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_13_69 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_135_113 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_49_108 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_49_119 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_89_266 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_38_22 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA_fanout76_A net77 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_85_461 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_110_60 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_110_71 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_119_91 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_1280_ core.cnb.result_out\[2\] _0640_ VDD VSS VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_48_141 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_95_94 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_0995_ _0394_ _0421_ _0410_ _0420_ VDD VSS VSS VDD sky130_fd_sc_hd__or3_1
X_1616_ _0138_ _0142_ _0141_ VSS VDD VSS VDD sky130_fd_sc_hd__or2_1
XFILLER_5_81 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1547_ VSS VDD _0089_ core.cnb.next_data_register_w\[0\] core.cnb.result_out\[0\]
+ _0090_ VSS VDD sky130_fd_sc_hd__mux2_1
X_1478_ VDD VSS _0054_ core.osr.data_valid_r net57 VSS VDD sky130_fd_sc_hd__and2_1
XFILLER_86_258 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_131_15 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_24_13 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_50_372 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_40_34 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_108_102 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_92_206 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_120_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1401_ core.osr.result_r\[17\] _0746_ _0742_ VSS VDD VSS VDD sky130_fd_sc_hd__or2_1
X_1332_ _0687_ _0669_ _0665_ core.osr.result_r\[7\] core.osr.result_r\[6\] core.cnb.result_out\[6\]
+ VDD VSS VSS VDD sky130_fd_sc_hd__o2111a_1
X_1263_ VSS VDD _0627_ _0628_ core.cnb.average_sum_r\[2\] VSS VDD sky130_fd_sc_hd__xnor2_1
XFILLER_111_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xinput5 VDD VSS config_1_in[13] net5 VSS VDD sky130_fd_sc_hd__dlymetal6s2s_1
X_1194_ VDD VSS _0578_ _0577_ core.cnb.comparator_in VSS VDD sky130_fd_sc_hd__and2_1
XFILLER_91_272 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_51_136 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_51_169 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_0978_ _0296_ _0281_ _0403_ _0401_ _0404_ VSS VDD VSS VDD sky130_fd_sc_hd__o211a_1
XFILLER_10_15 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_126_15 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_102_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_19_57 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1459__A1 _0424_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1613__S core.osr.osr_mode_r\[0\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_27_122 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_42_103 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_82_272 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_42_125 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1568__B _0568_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_nmat_row_n[2] core.ndc.row_out_n\[2\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__0928__A _0353_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_46_464 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_92_95 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_0901_ _0327_ core.cnb.data_register_r\[2\] _0266_ VSS VDD VSS VDD sky130_fd_sc_hd__nand2_2
X_0832_ _0258_ _0256_ _0253_ _0257_ core.cnb.shift_register_r\[12\] VSS VDD VSS VDD
+ sky130_fd_sc_hd__a211o_2
XANTENNA__1386__B1 _0635_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1315_ _0671_ _0668_ core.osr.result_r\[6\] _0670_ VSS VDD VSS VDD sky130_fd_sc_hd__o21a_1
X_1246_ VSS VDD core.cnb.average_counter_r\[0\] _0617_ core.cnb.average_counter_r\[1\]
+ VSS VDD sky130_fd_sc_hd__xnor2_1
X_1177_ VSS VDD _0561_ core.cnb.average_counter_r\[1\] core.cnb.average_counter_r\[2\]
+ core.cnb.average_counter_r\[0\] VSS VDD sky130_fd_sc_hd__and3_1
XPHY_109 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1613__A1 core.osr.next_result_w\[7\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_137_69 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1129__B1 _0506_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_87_342 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_47_217 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_46_33 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_46_44 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_62_21 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_62_54 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_7_38 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1368__B1 _0635_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1100_ _0514_ _0466_ _0454_ _0376_ _0463_ VSS VDD VSS VDD sky130_fd_sc_hd__a31o_2
XFILLER_94_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1031_ _0456_ _0454_ _0394_ _0453_ _0455_ VSS VDD VSS VDD sky130_fd_sc_hd__and4_1
Xinput30 VSS VDD net30 config_2_in[7] VSS VDD sky130_fd_sc_hd__clkbuf_1
X_1795_ core.cnb.shift_register_r\[7\] net61 _0038_ net75 VSS VDD VSS VDD sky130_fd_sc_hd__dfrtp_4
X_0815_ core.cnb.shift_register_r\[15\] core.cnb.shift_register_r\[13\] _0241_ core.cnb.shift_register_r\[12\]
+ core.cnb.shift_register_r\[14\] VDD VSS VSS VDD sky130_fd_sc_hd__or4_1
XFILLER_84_334 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_85_879 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_1229_ _0428_ _0442_ _0361_ _0603_ _0604_ VSS VDD VSS VDD sky130_fd_sc_hd__a31o_1
XFILLER_52_253 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_52_242 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_57_43 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_76_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA_input19_A config_2_in[11] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_90_326 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_90_359 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_440 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_451 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_462 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_495 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_473 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_484 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_22_90 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1580_ _0110_ core.osr.osr_mode_r\[0\] VSS VDD VSS VDD sky130_fd_sc_hd__clkbuf_4
XANTENNA__1513__B1 net52 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_67_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1014_ VSS VDD _0439_ _0342_ _0434_ _0328_ _0438_ VSS VDD sky130_fd_sc_hd__a211o_1
X_1778_ core.osr.result_r\[10\] net69 core.osr.next_result_w\[10\] net56 VSS VDD VSS
+ VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_134_15 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_58_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_84_131 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_27_57 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_43_34 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_68_53 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_49_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_84_85 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_90_145 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_90_156 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_17_90 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_270 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_281 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_292 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_1701_ VSS VDD _0044_ _0202_ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_1632_ _0124_ _0155_ _0154_ core.osr.next_result_w\[12\] core.osr.next_result_w\[8\]
+ VSS VDD VSS VDD sky130_fd_sc_hd__o22a_1
XANTENNA__1706__S _0614_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1563_ VSS VDD _0088_ core.cnb.next_data_register_w\[8\] core.cnb.result_out\[8\]
+ _0098_ VSS VDD sky130_fd_sc_hd__mux2_1
X_1494_ _0059_ core.cnb.data_register_r\[8\] _0068_ core.cnb.data_register_r\[9\]
+ _0330_ VDD VSS VSS VDD sky130_fd_sc_hd__or4_1
XFILLER_120_17 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_13_48 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_129_48 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_135_125 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_1_105 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA_fanout69_A net74 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_85_473 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_54_44 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_54_66 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_54_99 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1776__RESET_B net69 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1192__A1 core.cnb.comparator_in VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_0994_ _0413_ _0406_ _0419_ _0420_ _0418_ VDD VSS VSS VDD sky130_fd_sc_hd__a211oi_4
XFILLER_117_103 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1615_ _0124_ _0141_ _0139_ _0140_ core.osr.next_result_w\[9\] _0232_ VSS VDD VSS
+ VDD sky130_fd_sc_hd__o221a_1
XANTENNA_cgen_enable_dlycontrol_in net23 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1546_ _0089_ _0088_ VSS VDD VSS VDD sky130_fd_sc_hd__clkbuf_4
XFILLER_5_93 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1477_ VSS VDD core.cnb.next_conv_finished_w _0053_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_39_120 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_54_123 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_82_421 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_54_167 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_24_69 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1200__A net53 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_49_66 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_49_99 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_120_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_105_61 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_105_72 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_65_43 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_85_281 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_105_94 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1400_ _0745_ _0742_ core.osr.result_r\[17\] VSS VDD VSS VDD sky130_fd_sc_hd__nand2_1
X_1331_ VSS VDD _0686_ _0653_ _0667_ _0651_ _0685_ VSS VDD sky130_fd_sc_hd__a211o_1
X_1262_ VSS VDD _0627_ core.cnb.average_sum_r\[1\] core.cnb.comparator_in core.cnb.average_sum_r\[0\]
+ VSS VDD sky130_fd_sc_hd__and3_1
XFILLER_49_440 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_111_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xinput6 VSS VDD net6 config_1_in[14] VSS VDD sky130_fd_sc_hd__clkbuf_1
X_1193_ _0308_ _0577_ core.cnb.shift_register_r\[2\] core.cnb.shift_register_r\[3\]
+ VSS VDD VSS VDD sky130_fd_sc_hd__nor3_1
XFILLER_91_251 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_51_104 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0843__B core.cnb.shift_register_r\[1\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_0977_ _0403_ _0276_ _0282_ _0402_ VSS VDD VSS VDD sky130_fd_sc_hd__a21o_2
X_1529_ VSS VDD core.ndc.row_out_n\[15\] _0084_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_102_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_19_69 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_55_421 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1459__A2 _0520_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_35_24 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_42_115 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_82_295 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_35_68 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_51_45 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_51_67 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_51_78 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_51_89 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA_nmat_row_n[1] core.ndc.row_out_n\[1\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_111_109 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_90 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_0900_ _0325_ _0326_ _0306_ _0314_ VSS VDD VSS VDD sky130_fd_sc_hd__nor3_2
X_0831_ _0257_ _0254_ _0252_ _0255_ VSS VDD VSS VDD sky130_fd_sc_hd__o21a_1
X_1314_ VDD VSS _0670_ _0669_ _0665_ VSS VDD sky130_fd_sc_hd__and2_1
X_1245_ _0616_ _0613_ VSS VDD VSS VDD sky130_fd_sc_hd__clkbuf_4
XFILLER_49_281 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1176_ core.cnb.average_counter_r\[0\] _0560_ _0559_ core.cnb.average_counter_r\[1\]
+ core.cnb.sampled_avg_control_r\[1\] VSS VDD VSS VDD sky130_fd_sc_hd__o22a_1
XFILLER_112_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_137_15 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_47_229 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_46_89 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_102_40 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_102_95 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_30_129 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_11_81 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_97_118 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_97_129 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_1030_ VDD VSS _0455_ _0374_ _0363_ VSS VDD sky130_fd_sc_hd__and2_1
XFILLER_21_107 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_0814_ core.cnb.is_sampling_w core.cnb.shift_register_r\[7\] core.cnb.shift_register_r\[1\]
+ core.cnb.shift_register_r\[6\] _0240_ VDD VSS VSS VDD sky130_fd_sc_hd__or4_4
Xinput31 VSS VDD net31 config_2_in[8] VSS VDD sky130_fd_sc_hd__clkbuf_1
Xinput20 VSS VDD net20 config_2_in[12] VSS VDD sky130_fd_sc_hd__clkbuf_1
X_1794_ core.cnb.shift_register_r\[6\] net61 _0037_ net77 VSS VDD VSS VDD sky130_fd_sc_hd__dfrtp_4
X_1228_ _0408_ _0603_ _0602_ VSS VDD VSS VDD sky130_fd_sc_hd__nor2_1
XFILLER_52_210 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_16_37 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_52_221 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1159_ _0342_ _0328_ _0344_ _0546_ VDD VSS VSS VDD sky130_fd_sc_hd__a21o_1
XFILLER_52_276 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_57_66 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_57_77 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_90_338 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_113_61 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_73_76 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_430 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_441 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_452 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_463 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_474 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_485 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_496 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_1013_ _0438_ _0366_ _0345_ VSS VDD VSS VDD sky130_fd_sc_hd__nand2_1
X_1777_ core.osr.result_r\[9\] net69 core.osr.next_result_w\[9\] net56 VSS VDD VSS
+ VDD sky130_fd_sc_hd__dfrtp_4
XFILLER_89_449 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_84_165 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_84_176 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1203__A net53 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_4_29 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA_input31_A config_2_in[8] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_48_357 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_17_80 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XPHY_260 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_271 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_282 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_293 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_1700_ VSS VDD _0614_ _0255_ _0252_ _0202_ VSS VDD sky130_fd_sc_hd__mux2_1
X_1631_ _0154_ _0111_ _0216_ VSS VDD VSS VDD sky130_fd_sc_hd__nand2_1
X_1562_ VSS VDD _0010_ _0097_ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_1493_ _0264_ _0552_ _0067_ core.cnb.data_register_r\[10\] _0540_ VDD VSS VSS VDD
+ sky130_fd_sc_hd__or4_1
XFILLER_86_408 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_120_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_129_16 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1752__CLK net55 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1489__B1 _0433_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_70_66 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_79_42 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_135_81 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_48_121 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_95_63 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_0993_ VSS VDD _0419_ _0406_ _0364_ _0417_ VSS VDD sky130_fd_sc_hd__and3_1
XANTENNA_pmat_row_n[14] core.pdc.row_out_n\[14\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1775__CLK net56 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_132_118 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1614_ _0140_ _0219_ _0134_ core.osr.next_result_w\[3\] VSS VDD VSS VDD sky130_fd_sc_hd__o21a_1
X_1545_ VDD VSS _0088_ _0568_ core.cnb.shift_register_r\[2\] VSS VDD sky130_fd_sc_hd__and2_1
XANTENNA__1018__A _0345_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1476_ VDD VSS _0053_ _0614_ core.cnb.shift_register_r\[1\] VSS VDD sky130_fd_sc_hd__and2_1
XFILLER_115_29 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_82_477 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_40_25 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_40_69 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_40_58 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_40_47 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_49_34 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_45_124 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_45_113 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_121_50 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1634__B1 _0236_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1798__CLK net77 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_53_8 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1330_ _0685_ core.osr.result_r\[7\] core.cnb.result_out\[6\] VSS VDD VSS VDD sky130_fd_sc_hd__nand2_1
X_1261_ _0626_ core.cnb.next_average_sum_w\[1\] _0616_ VSS VDD VSS VDD sky130_fd_sc_hd__nor2_1
XFILLER_49_430 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xinput7 VSS VDD net7 config_1_in[15] VSS VDD sky130_fd_sc_hd__clkbuf_1
X_1192_ _0576_ _0575_ _0572_ _0570_ _0569_ core.cnb.comparator_in VDD VSS VSS VDD
+ sky130_fd_sc_hd__o2111a_1
XFILLER_49_463 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_36_124 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0843__C core.cnb.is_sampling_w VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1625__A0 _0691_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_0976_ _0402_ _0268_ _0261_ _0258_ _0278_ VDD VSS VSS VDD sky130_fd_sc_hd__o31ai_1
X_1528_ _0077_ _0084_ core.ndc.row_out_n\[12\] VSS VDD VSS VDD sky130_fd_sc_hd__or2_1
XFILLER_19_26 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1459_ _0424_ _0474_ core.ndc.col_out_n\[16\] _0520_ VDD VSS VSS VDD sky130_fd_sc_hd__a21oi_1
XFILLER_27_113 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_55_477 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_82_241 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1211__A _0588_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_50_182 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_46_444 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_91 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_80 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_30_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_0830_ VSS VDD _0255_ _0256_ _0254_ VSS VDD sky130_fd_sc_hd__xnor2_1
X_1313_ core.cnb.result_out\[4\] core.osr.result_r\[4\] _0669_ core.osr.result_r\[5\]
+ core.cnb.result_out\[5\] VDD VSS VSS VDD sky130_fd_sc_hd__a22o_1
XFILLER_97_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1244_ core.cnb.next_average_counter_w\[0\] _0615_ core.cnb.average_counter_r\[0\]
+ VSS VDD VSS VDD sky130_fd_sc_hd__nand2_1
X_1175_ _0559_ _0558_ _0557_ VSS VDD VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_24_116 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_52_425 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1031__A _0394_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__0870__A core.cnb.data_register_r\[1\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_21_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_137_27 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_0959_ core.cnb.data_register_r\[6\] _0385_ VDD VSS VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_88_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_101_121 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_87_366 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_87_377 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_62_45 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_12_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_11_93 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_87_42 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_79_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__0955__A _0366_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_0813_ VDD VSS _0239_ _0238_ VSS VDD sky130_fd_sc_hd__buf_6
Xinput10 VDD VSS net10 config_1_in[3] VSS VDD sky130_fd_sc_hd__buf_2
Xinput21 VSS VDD net21 config_2_in[13] VSS VDD sky130_fd_sc_hd__clkbuf_1
X_1793_ core.cnb.shift_register_r\[5\] net62 _0036_ net76 VSS VDD VSS VDD sky130_fd_sc_hd__dfrtp_4
Xinput32 VSS VDD net32 config_2_in[9] VSS VDD sky130_fd_sc_hd__clkbuf_1
XANTENNA__1359__A2 core.cnb.result_out\[8\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1026__A _0394_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_84_303 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1227_ VSS VDD _0601_ _0385_ _0599_ _0602_ core.cnb.data_register_r\[7\] VSS VDD
+ sky130_fd_sc_hd__a2bb2o_1
X_1158_ _0545_ _0542_ _0544_ VSS VDD VSS VDD sky130_fd_sc_hd__and2b_1
XFILLER_52_233 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1089_ VSS VDD _0505_ _0424_ _0506_ core.pdc.col_out_n\[8\] VSS VDD sky130_fd_sc_hd__o21ai_1
XANTENNA__1047__A1 _0354_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_87_185 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_113_95 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_73_66 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_420 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_431 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_442 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_453 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_486 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_464 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_475 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_497 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_22_81 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_98_74 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_98_85 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1513__A2 _0079_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1012_ _0349_ _0435_ _0348_ _0437_ _0434_ VDD VSS VSS VDD sky130_fd_sc_hd__or4b_1
X_1776_ core.osr.result_r\[8\] net69 core.osr.next_result_w\[8\] net56 VSS VDD VSS
+ VDD sky130_fd_sc_hd__dfrtp_2
XFILLER_27_26 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_43_14 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1440__A1 _0529_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__0951__B1 core.cnb.data_register_r\[5\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_68_22 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_68_33 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_48_325 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_input24_A config_2_in[1] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_90_114 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_261 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_250 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_129_113 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XPHY_272 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_283 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_294 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_1630_ _0150_ _0153_ _0115_ _0151_ _0022_ VSS VDD VSS VDD sky130_fd_sc_hd__a31o_1
X_1561_ VSS VDD _0089_ core.cnb.next_data_register_w\[7\] core.cnb.result_out\[7\]
+ _0097_ VSS VDD sky130_fd_sc_hd__mux2_1
X_1492_ core.cnb.data_register_r\[9\] _0066_ _0059_ _0541_ VDD VSS VSS VDD sky130_fd_sc_hd__or3_1
XFILLER_47_380 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_135_105 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_1759_ net49 net66 _0022_ net55 VSS VDD VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_132_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_38_36 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_54_35 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_54_79 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_110_41 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_110_85 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_123_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_135_93 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_48_166 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_48_177 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_0992_ _0417_ _0406_ _0413_ _0418_ _0364_ VDD VSS VSS VDD sky130_fd_sc_hd__a211oi_2
X_1613_ VSS VDD core.osr.osr_mode_r\[0\] core.osr.next_result_w\[7\] core.osr.next_result_w\[5\]
+ _0139_ VSS VDD sky130_fd_sc_hd__mux2_1
X_1544_ VSS VDD _0002_ _0087_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_114_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1475_ _0533_ _0450_ _0423_ core.ndc.col_out_n\[30\] VDD VSS VSS VDD sky130_fd_sc_hd__a21o_1
XFILLER_86_239 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1034__A _0394_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_82_445 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_108_127 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1209__A _0579_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_105_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_49_57 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_65_67 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1634__A1 core.cnb.result_out\[4\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_14_60 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1553__S _0089_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1260_ _0625_ _0626_ core.cnb.average_sum_r\[1\] VDD VSS VSS VDD sky130_fd_sc_hd__xor2_1
X_1191_ _0574_ core.cnb.sampled_avg_control_r\[1\] _0575_ VSS VDD VSS VDD sky130_fd_sc_hd__or2b_1
Xinput8 VSS VDD net8 config_1_in[1] VSS VDD sky130_fd_sc_hd__clkbuf_1
XANTENNA__1742__CLK net81 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1625__A1 _0709_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_0975_ _0401_ _0397_ _0289_ _0399_ _0287_ VSS VDD _0400_ VSS VDD sky130_fd_sc_hd__a221o_1
XFILLER_10_29 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1029__A _0420_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1527_ core.pdc.row_out_n\[2\] core.ndc.row_out_n\[14\] VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_4
XANTENNA__1561__A0 core.cnb.result_out\[7\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1458_ _0529_ _0474_ core.ndc.col_out_n\[15\] _0520_ VDD VSS VSS VDD sky130_fd_sc_hd__a21oi_1
XFILLER_82_220 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1313__B1 core.cnb.result_out\[5\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1389_ VSS VDD _0737_ core.osr.result_r\[13\] core.osr.result_r\[12\] _0729_ VSS
+ VDD sky130_fd_sc_hd__and3_1
XFILLER_82_253 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_51_25 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_76_22 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_76_33 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_116_95 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_46_412 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_46_456 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_25_81 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_92 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_81 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_70 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_30_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1312_ _0651_ _0667_ _0668_ _0653_ VDD VSS VSS VDD sky130_fd_sc_hd__a21oi_1
XFILLER_97_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_2_41 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1243_ _0614_ _0615_ VDD VSS VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_2_85 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1015__C _0373_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1174_ _0558_ core.cnb.sampled_avg_control_r\[2\] core.cnb.sampled_avg_control_r\[0\]
+ VSS VDD VSS VDD sky130_fd_sc_hd__and2b_1
XFILLER_52_437 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_21_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_0958_ _0325_ _0338_ _0384_ _0379_ VDD VSS VSS VDD sky130_fd_sc_hd__a21oi_1
XFILLER_137_39 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_0889_ core.cnb.shift_register_r\[16\] _0315_ VDD VSS VSS VDD sky130_fd_sc_hd__inv_2
XANTENNA__1534__B1 net52 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1206__B _0579_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_88_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_46_25 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_87_389 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_15_106 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1222__A _0588_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_102_64 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_62_79 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_134_3 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_12_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_127_50 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1116__B _0394_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_79_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_46_253 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_36_91 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_0812_ core.cnb.shift_register_r\[4\] core.cnb.shift_register_r\[2\] _0238_ core.cnb.shift_register_r\[3\]
+ core.cnb.shift_register_r\[5\] VDD VSS VSS VDD sky130_fd_sc_hd__or4_1
Xinput11 net11 config_1_in[4] VSS VDD VSS VDD sky130_fd_sc_hd__clkbuf_4
Xinput22 VSS VDD net22 config_2_in[14] VSS VDD sky130_fd_sc_hd__clkbuf_1
Xinput33 VSS VDD net33 rst_n VSS VDD sky130_fd_sc_hd__clkbuf_1
X_1792_ core.cnb.shift_register_r\[4\] net60 _0035_ net76 VSS VDD VSS VDD sky130_fd_sc_hd__dfrtp_4
XANTENNA__1307__A core.cnb.result_out\[5\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1026__B _0410_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1226_ VSS VDD _0600_ _0385_ _0382_ _0601_ VSS VDD sky130_fd_sc_hd__o21ai_1
XFILLER_16_17 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_1157_ VSS VDD _0543_ _0544_ core.cnb.data_register_r\[11\] VSS VDD sky130_fd_sc_hd__xnor2_1
XFILLER_12_109 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_52_267 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1088_ _0506_ _0462_ _0463_ VSS VDD VSS VDD sky130_fd_sc_hd__nand2_2
XFILLER_52_289 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1047__A2 _0465_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_32_49 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_57_35 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_57_57 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_87_175 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_87_197 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_113_52 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_73_45 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_410 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1803__CLK net77 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XPHY_421 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_432 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_443 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_454 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_465 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_476 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_498 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_487 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_7_113 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_98_42 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_21_7 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1561__S _0089_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1011_ _0436_ _0435_ _0434_ VSS VDD VSS VDD sky130_fd_sc_hd__nand2_1
XANTENNA__0788__A1 core.osr.osr_mode_r\[0\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1775_ core.osr.result_r\[7\] net68 core.osr.next_result_w\[7\] net56 VSS VDD VSS
+ VDD sky130_fd_sc_hd__dfrtp_4
Xnmat nmat/vcm sample_nmatrix_cgen sample_nmatrix_cgen_n core.ndc.row_out_n\[15\]
+ core.ndc.row_out_n\[14\] core.ndc.row_out_n\[13\] core.ndc.row_out_n\[12\] core.ndc.row_out_n\[11\]
+ core.ndc.row_out_n\[10\] core.ndc.row_out_n\[9\] core.cnb.pswitch_out\[11\] core.ndc.row_out_n\[7\]
+ core.ndc.row_out_n\[6\] core.ndc.row_out_n\[5\] core.ndc.row_out_n\[4\] core.ndc.row_out_n\[3\]
+ core.ndc.row_out_n\[2\] core.ndc.row_out_n\[1\] net83 net101 core.ndc.row_out_n\[15\]
+ core.ndc.row_out_n\[14\] core.ndc.row_out_n\[13\] core.ndc.row_out_n\[12\] core.ndc.row_out_n\[11\]
+ core.ndc.row_out_n\[10\] core.ndc.row_out_n\[9\] core.cnb.pswitch_out\[11\] core.ndc.row_out_n\[7\]
+ core.ndc.row_out_n\[6\] core.ndc.row_out_n\[5\] core.ndc.row_out_n\[4\] core.ndc.row_out_n\[3\]
+ core.ndc.row_out_n\[2\] core.ndc.row_out_n\[1\] core.ndc.col_out_n\[31\] core.ndc.col_out_n\[30\]
+ core.ndc.col_out_n\[29\] core.ndc.col_out_n\[28\] core.ndc.col_out_n\[27\] core.ndc.col_out_n\[26\]
+ core.ndc.col_out_n\[25\] core.ndc.col_out_n\[24\] core.ndc.col_out_n\[23\] core.ndc.col_out_n\[22\]
+ core.ndc.col_out_n\[21\] core.ndc.col_out_n\[20\] core.ndc.col_out_n\[19\] core.ndc.col_out_n\[18\]
+ core.ndc.col_out_n\[17\] core.ndc.col_out_n\[16\] core.ndc.col_out_n\[15\] core.ndc.col_out_n\[14\]
+ core.ndc.col_out_n\[13\] core.ndc.col_out_n\[12\] core.ndc.col_out_n\[11\] core.ndc.col_out_n\[10\]
+ core.ndc.col_out_n\[9\] core.ndc.col_out_n\[8\] core.ndc.col_out_n\[7\] core.ndc.col_out_n\[6\]
+ core.ndc.col_out_n\[5\] core.ndc.col_out_n\[4\] core.ndc.col_out_n\[3\] core.ndc.col_out_n\[2\]
+ core.ndc.col_out_n\[1\] core.ndc.col_out_n\[0\] core.cnb.pswitch_out\[2\] core.cnb.pswitch_out\[1\]
+ core.cnb.pswitch_out\[0\] net82 core.cnb.is_sampling_w core.cnb.enable_loop_out
+ inn_analog ctop_nmatrix_analog VSS VDD adc_array_matrix_12bit
XFILLER_134_29 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_27_38 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1209_ _0579_ _0417_ _0589_ _0413_ VSS VDD VSS VDD sky130_fd_sc_hd__or3b_1
XFILLER_84_189 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1440__A2 _0460_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_108_96 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_1_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_124_62 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA_input17_A config_2_in[0] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XPHY_240 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_251 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_129_125 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XPHY_273 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_262 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_284 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_295 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_76_8 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_1560_ VSS VDD _0009_ _0096_ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_1491_ core.cnb.data_register_r\[8\] _0065_ _0059_ _0344_ VDD VSS VSS VDD sky130_fd_sc_hd__or3_1
X_1758_ net48 net70 _0021_ net54 VSS VDD VSS VDD sky130_fd_sc_hd__dfrtp_1
X_1689_ VSS VDD _0038_ _0196_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_132_879 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA_input9_A config_1_in[2] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_38_59 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1110__A1 _0449_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_70_46 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_123_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_0991_ _0359_ _0417_ _0414_ _0416_ _0365_ _0415_ VSS VDD VSS VDD sky130_fd_sc_hd__o221a_1
X_1612_ _0132_ core.cnb.result_out\[1\] _0137_ _0138_ VDD VSS VSS VDD sky130_fd_sc_hd__a21o_1
X_1543_ VSS VDD _0588_ net9 core.cnb.sampled_avg_control_r\[2\] _0087_ VSS VDD sky130_fd_sc_hd__mux2_1
X_1474_ core.ndc.col_out_n\[29\] _0450_ _0465_ _0534_ VSS VDD VSS VDD sky130_fd_sc_hd__o21a_1
XFILLER_114_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_82_457 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_50_332 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_50_365 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_50_387 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_50_398 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1196__S _0579_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_123_109 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1159__A1 _0328_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_105_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_105_31 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA_fanout67_A net69 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_85_240 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1331__A1 _0651_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_45_104 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_53_181 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_81_45 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_14_72 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_114_109 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_46_9 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_39_80 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1190_ VSS VDD core.cnb.sampled_avg_control_r\[2\] core.cnb.comparator_in _0573_
+ _0574_ VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_49_454 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_49_476 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__0974__A core.cnb.data_register_r\[0\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xinput9 VSS VDD net9 config_1_in[2] VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_91_221 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_91_232 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_0974_ VSS VDD _0400_ _0282_ core.cnb.data_register_r\[0\] _0285_ VSS VDD sky130_fd_sc_hd__and3_1
X_1526_ VDD VSS core.pdc.row_out_n\[2\] _0083_ VSS VDD sky130_fd_sc_hd__buf_6
X_1457_ _0775_ _0354_ _0518_ core.ndc.col_out_n\[14\] VDD VSS VSS VDD sky130_fd_sc_hd__a21o_1
XANTENNA__1313__A1 core.cnb.result_out\[4\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1388_ _0736_ _0212_ VSS VDD VSS VDD sky130_fd_sc_hd__clkbuf_4
XFILLER_55_468 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_50_173 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_51_37 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_116_85 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_76_78 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_18_126 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_46_435 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_33_107 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_33_129 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_82 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_71 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_60 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_93 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1775__D core.osr.next_result_w\[7\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1311_ _0665_ _0666_ _0664_ _0667_ VSS VDD VSS VDD sky130_fd_sc_hd__nand3b_1
X_1242_ _0614_ _0613_ VSS VDD VSS VDD sky130_fd_sc_hd__clkbuf_4
XFILLER_2_53 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1173_ _0557_ core.cnb.average_counter_r\[0\] core.cnb.average_counter_r\[1\] VSS
+ VDD VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_2_97 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_52_416 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_52_449 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_0957_ core.cnb.data_register_r\[6\] _0383_ _0382_ VSS VDD VSS VDD sky130_fd_sc_hd__or2_1
X_0888_ _0313_ _0314_ _0307_ VSS VDD VSS VDD sky130_fd_sc_hd__nor2_1
XANTENNA__1534__A1 _0079_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1509_ VSS VDD core.ndc.row_out_n\[3\] _0078_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_87_324 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_51_471 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1470__B1 core.pdc.col_out_n\[24\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_11_51 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0789__A core.osr.osr_mode_r\[0\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_86_390 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1559__S _0089_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1461__B1 _0514_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_0811_ core.cnb.shift_register_r\[10\] core.cnb.shift_register_r\[9\] _0237_ core.cnb.shift_register_r\[8\]
+ core.cnb.shift_register_r\[11\] VDD VSS VSS VDD sky130_fd_sc_hd__or4b_2
X_1791_ core.cnb.shift_register_r\[3\] net62 _0034_ net75 VSS VDD VSS VDD sky130_fd_sc_hd__dfrtp_4
Xinput12 VDD VSS net12 config_1_in[5] VSS VDD sky130_fd_sc_hd__buf_2
Xinput34 VSS VDD net34 start_conversion_in VSS VDD sky130_fd_sc_hd__clkbuf_1
Xinput23 VSS VDD net23 config_2_in[15] VSS VDD sky130_fd_sc_hd__clkbuf_1
X_1225_ _0242_ _0268_ _0600_ _0279_ _0277_ VDD VSS VSS VDD sky130_fd_sc_hd__or4_1
XFILLER_84_349 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1156_ _0242_ _0315_ _0543_ _0279_ _0245_ VDD VSS VSS VDD sky130_fd_sc_hd__or4_1
X_1087_ _0503_ _0505_ _0466_ VSS VDD VSS VDD sky130_fd_sc_hd__nor2_1
XFILLER_20_110 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_32_39 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_113_9 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_73_35 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_83_393 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_113_75 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XPHY_400 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_411 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_422 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_433 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_444 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_455 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_466 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_477 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_499 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_488 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1779__RESET_B net67 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_98_54 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1010_ VDD VSS _0435_ _0366_ _0347_ VSS VDD sky130_fd_sc_hd__and2_1
XFILLER_8_41 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1778__CLK net56 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_8_85 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1774_ core.osr.result_r\[6\] net68 core.osr.next_result_w\[6\] net56 VSS VDD VSS
+ VDD sky130_fd_sc_hd__dfrtp_4
XANTENNA__1318__A core.cnb.result_out\[6\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1037__B _0460_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1208_ VDD VSS _0588_ core.cnb.is_sampling_w VSS VDD sky130_fd_sc_hd__buf_4
X_1139_ _0456_ core.ndc.col_out_n\[31\] _0352_ VSS VDD VSS VDD sky130_fd_sc_hd__nor2_1
XANTENNA__1673__B1 _0236_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1199__S _0579_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1425__B1 _0236_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1801__RESET_B net63 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_1_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_124_85 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_84_67 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1410__B _0236_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XPHY_241 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_252 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_230 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_274 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_263 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_285 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_296 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1195__A2 _0568_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1138__A _0374_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1490_ _0064_ _0059_ core.cnb.data_register_r\[9\] _0433_ _0344_ core.cnb.data_register_r\[8\]
+ VDD VSS VSS VDD sky130_fd_sc_hd__o2111a_1
XFILLER_47_393 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1757_ net47 net70 _0020_ net54 VSS VDD VSS VDD sky130_fd_sc_hd__dfrtp_1
X_1688_ VSS VDD _0616_ core.cnb.shift_register_r\[8\] core.cnb.shift_register_r\[7\]
+ _0196_ VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_89_216 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_38_49 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_85_433 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1511__A _0352_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_53_374 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1110__A2 _0519_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_53_385 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_110_98 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_126_129 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_119_63 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_119_85 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_135_51 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_60_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1778__D core.osr.next_result_w\[10\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_0990_ _0281_ _0296_ _0416_ _0371_ _0365_ _0297_ VSS VDD VSS VDD sky130_fd_sc_hd__a311o_1
XANTENNA__1723__RESET_B net63 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1611_ _0133_ net47 _0137_ _0103_ VSS VDD VSS VDD sky130_fd_sc_hd__and3b_1
XFILLER_5_31 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1542_ VSS VDD _0001_ _0086_ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_1473_ _0424_ _0464_ core.ndc.col_out_n\[28\] _0460_ VDD VSS VSS VDD sky130_fd_sc_hd__a21oi_1
XFILLER_82_414 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_24_29 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_51_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1809_ core.osr.sample_count_r\[4\] net72 core.osr.next_sample_count_w\[4\] net57
+ VSS VDD VSS VDD sky130_fd_sc_hd__dfrtp_4
XANTENNA__1159__A2 _0342_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1506__A core.pdc.row_out_n\[14\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_49_48 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_85_252 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_85_263 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_105_87 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_81_24 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_42_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_30_61 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_49_400 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_91_244 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1086__A1 _0450_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_91_266 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_33_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_0973_ _0398_ _0242_ _0399_ _0261_ _0268_ VSS VDD VSS VDD sky130_fd_sc_hd__nor4_1
X_1525_ VSS VDD _0083_ _0607_ _0556_ _0079_ VSS VDD sky130_fd_sc_hd__and3_1
X_1456_ VSS VDD _0468_ _0376_ _0474_ _0775_ VSS VDD sky130_fd_sc_hd__o21ai_1
X_1387_ _0735_ core.osr.next_result_w\[13\] VSS VDD VSS VDD sky130_fd_sc_hd__clkbuf_2
XANTENNA__1061__A _0347_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_82_266 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_24_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_76_57 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_132_85 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1068__A1 _0328_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XPHY_83 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_72 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_15_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XPHY_61 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_50 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_92_89 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_94 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_41_82 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_41_71 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_nmat_rowon_n[3] core.ndc.row_out_n\[4\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1310_ core.osr.result_r\[4\] _0666_ core.cnb.result_out\[4\] VDD VSS VSS VDD sky130_fd_sc_hd__xor2_1
XANTENNA__0985__A core.cnb.data_register_r\[2\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1241_ _0577_ _0613_ _0568_ VSS VDD VSS VDD sky130_fd_sc_hd__or2_1
XFILLER_2_65 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1172_ core.cnb.is_sampling_w core.cnb.enable_loop_out VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_4
XFILLER_24_108 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_0956_ _0382_ _0303_ _0304_ VSS VDD VSS VDD sky130_fd_sc_hd__nand2_1
X_0887_ _0313_ _0310_ _0308_ _0291_ _0243_ _0312_ VDD VSS VSS VDD sky130_fd_sc_hd__o32a_1
XANTENNA__1534__A2 _0080_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1508_ VDD VSS _0078_ _0077_ core.ndc.row_out_n\[4\] VSS VDD sky130_fd_sc_hd__and2_1
XFILLER_87_314 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0895__A core.cnb.data_register_r\[5\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1439_ _0354_ _0465_ core.ndc.col_out_n\[2\] _0448_ _0769_ VDD VSS VSS VDD sky130_fd_sc_hd__a22o_1
XFILLER_55_233 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_55_244 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_102_77 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1470__A1 _0424_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__0972__C_N core.cnb.data_register_r\[0\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_127_63 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_2_3 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1461__A1 _0424_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_0810_ core.osr.is_last_sample _0236_ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_2
X_1790_ core.cnb.shift_register_r\[2\] net62 _0033_ net77 VSS VDD VSS VDD sky130_fd_sc_hd__dfrtp_4
Xinput13 VSS VDD net13 config_1_in[6] VSS VDD sky130_fd_sc_hd__clkbuf_1
Xinput24 VSS VDD net24 config_2_in[1] VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_35_3 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1224_ _0553_ _0255_ _0599_ _0254_ VSS VDD VSS VDD sky130_fd_sc_hd__or3b_1
X_1155_ VSS VDD _0541_ core.cnb.data_register_r\[9\] core.cnb.data_register_r\[10\]
+ _0542_ VSS VDD sky130_fd_sc_hd__o21ai_1
XFILLER_92_350 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1086_ core.pdc.col_out_n\[7\] _0450_ _0452_ _0504_ VSS VDD VSS VDD sky130_fd_sc_hd__o21a_1
XFILLER_20_122 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1452__A1 _0449_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_0939_ VDD VSS _0365_ _0329_ VSS VDD sky130_fd_sc_hd__buf_6
XANTENNA__0963__B1 core.cnb.data_register_r\[2\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1063__S0 _0373_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_57_26 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_87_144 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_87_133 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1514__A core.pdc.row_out_n\[10\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_113_21 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_83_361 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_401 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_412 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_423 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_434 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_445 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_456 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_467 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_489 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_478 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_98_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_8_53 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_8_97 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1773_ core.osr.result_r\[5\] net68 core.osr.next_result_w\[5\] net56 VSS VDD VSS
+ VDD sky130_fd_sc_hd__dfrtp_1
XANTENNA__1370__B1 core.cnb.result_out\[10\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1207_ net53 _0587_ _0586_ core.cnb.data_register_r\[3\] core.cnb.next_data_register_w\[3\]
+ VSS VDD VSS VDD sky130_fd_sc_hd__o211a_1
X_1138_ _0422_ _0534_ _0374_ VSS VDD VSS VDD sky130_fd_sc_hd__nor2_1
XANTENNA__1673__A1 core.cnb.result_out\[11\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1069_ _0373_ _0348_ _0490_ _0349_ _0488_ VDD VSS VSS VDD sky130_fd_sc_hd__or4_1
XANTENNA__1722__CLK net81 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_135_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_108_76 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_48_317 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_17_51 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_220 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_231 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_242 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_253 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_264 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_275 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_286 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_297 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_126_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__0993__A _0364_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_54_309 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1756_ net46 net66 _0019_ net54 VSS VDD VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_117_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1687_ VSS VDD _0037_ _0195_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XANTENNA__1591__B1 core.osr.next_result_w\[6\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_85_445 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_53_320 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_110_77 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1239__A net53 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_108_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_48_103 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1768__CLK net55 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_input22_A config_2_in[14] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_95_78 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_28_72 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_44_93 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_60_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_81_8 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA_pmat_row_n[10] core.pdc.row_out_n\[10\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1149__A core.cnb.nswitch_out\[1\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_60_70 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1610_ _0131_ _0129_ _0136_ _0019_ VDD VSS VSS VDD sky130_fd_sc_hd__a21o_1
X_1541_ VSS VDD _0588_ net8 core.cnb.sampled_avg_control_r\[1\] _0086_ VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_5_43 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1472_ _0424_ _0532_ core.ndc.col_out_n\[27\] _0422_ VDD VSS VSS VDD sky130_fd_sc_hd__a21oi_1
XFILLER_86_209 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_39_103 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_82_437 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_51_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1808_ core.osr.sample_count_r\[3\] net71 core.osr.next_sample_count_w\[3\] net57
+ VSS VDD VSS VDD sky130_fd_sc_hd__dfrtp_1
XANTENNA__1059__A _0364_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1739_ core.cnb.average_sum_r\[4\] net60 core.cnb.next_average_sum_w\[4\] net76 VSS
+ VDD VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_131_100 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_85_220 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_85_297 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1619__B2 core.osr.next_result_w\[6\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1241__B _0568_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_42_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_121_98 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_14_41 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1555__A0 core.cnb.result_out\[4\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_33_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_0972_ _0244_ core.cnb.data_register_r\[0\] _0398_ core.cnb.shift_register_r\[4\]
+ VSS VDD VSS VDD sky130_fd_sc_hd__or3b_1
X_1524_ VSS VDD core.ndc.row_out_n\[13\] _0082_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_113_122 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_1455_ VSS VDD _0519_ _0449_ _0514_ core.ndc.col_out_n\[13\] VSS VDD sky130_fd_sc_hd__o21ai_1
X_1386_ _0735_ _0733_ _0635_ _0734_ VSS VDD VSS VDD sky130_fd_sc_hd__o21a_1
XFILLER_82_201 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_35_18 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_82_289 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_24_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_136_9 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_116_10 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_pmat_col_n[18] core.pdc.col_out_n\[18\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_116_54 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_fanout72_A net73 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1252__A _0616_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_132_64 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_40 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1068__A2 _0342_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_92_57 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_92_79 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_73 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_62 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_15_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XPHY_51 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_95 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_84 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_41_61 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_41_94 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_1240_ VSS VDD core.cnb.next_data_register_w\[11\] _0612_ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_1171_ core.cnb.pswitch_out\[11\] net52 VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_2
XFILLER_2_77 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_49_297 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_0955_ _0381_ _0366_ _0380_ _0378_ VSS VDD VSS VDD sky130_fd_sc_hd__nand3_1
X_0886_ _0312_ _0311_ _0237_ _0286_ VDD VSS VSS VDD sky130_fd_sc_hd__a21boi_1
XANTENNA__1337__A _0691_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1507_ _0077_ _0352_ _0607_ VSS VDD VSS VDD sky130_fd_sc_hd__nand2_4
X_1438_ _0452_ _0769_ _0353_ VSS VDD VSS VDD sky130_fd_sc_hd__nor2_1
XANTENNA__1072__A _0345_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1369_ core.osr.next_result_w\[10\] _0720_ core.cnb.result_out\[10\] VSS VDD VSS
+ VDD sky130_fd_sc_hd__xnor2_4
XFILLER_102_89 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1207__C1 net53 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1247__A _0616_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__0981__A1 _0364_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_127_75 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_99_9 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1461__A2 _0519_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_52_60 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xinput14 VSS VDD net14 config_1_in[7] VSS VDD sky130_fd_sc_hd__clkbuf_1
Xinput25 VSS VDD net25 config_2_in[2] VSS VDD sky130_fd_sc_hd__clkbuf_1
X_1223_ _0264_ _0598_ _0258_ VSS VDD VSS VDD sky130_fd_sc_hd__or2_1
X_1154_ _0540_ _0541_ _0264_ VSS VDD VSS VDD sky130_fd_sc_hd__nor2_2
XFILLER_52_204 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1085_ VDD VSS _0504_ _0503_ _0466_ VSS VDD sky130_fd_sc_hd__and2_1
XFILLER_92_373 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1452__A2 _0515_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_0938_ VDD VSS _0364_ core.cnb.data_register_r\[4\] VSS VDD sky130_fd_sc_hd__buf_4
X_0869_ _0294_ core.cnb.shift_register_r\[4\] _0293_ _0291_ _0274_ _0295_ VSS VDD
+ VSS VDD sky130_fd_sc_hd__a2111oi_4
XANTENNA__1063__S1 _0433_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1140__A1 _0354_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_83_373 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_113_88 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1530__A _0077_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XPHY_402 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_413 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_424 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_435 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_446 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_457 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_468 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_7_105 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XPHY_479 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_138_41 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_22_85 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_138_85 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_4_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_98_67 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_47_93 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_8_65 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1772_ core.osr.result_r\[4\] net68 core.osr.next_result_w\[4\] net56 VSS VDD VSS
+ VDD sky130_fd_sc_hd__dfrtp_4
XFILLER_84_115 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_1206_ _0363_ _0587_ _0579_ VSS VDD VSS VDD sky130_fd_sc_hd__or2_1
X_1137_ core.pdc.col_out_n\[29\] _0354_ _0533_ _0460_ VSS VDD VSS VDD sky130_fd_sc_hd__a21bo_1
XFILLER_92_181 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1068_ VSS VDD _0489_ _0342_ _0434_ _0328_ _0488_ VSS VDD sky130_fd_sc_hd__a211o_1
XFILLER_135_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_108_22 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_108_33 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_68_59 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_88_421 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1244__B _0615_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1361__A1 core.cnb.result_out\[6\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1113__A1 _0352_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_90_107 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_90_129 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1629__A1_N _0235_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XPHY_210 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_232 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_221 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_243 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_265 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_276 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_254 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_287 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_298 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_126_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1435__A _0450_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1755_ net45 net66 _0018_ net54 VSS VDD VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_117_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1686_ VSS VDD _0616_ core.cnb.shift_register_r\[7\] core.cnb.shift_register_r\[6\]
+ _0195_ VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_89_207 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_85_402 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_126_109 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_108_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_119_76 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_88_262 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_95_57 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_48_148 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_88_295 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_input15_A config_1_in[8] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_91_449 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_44_72 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1540_ VSS VDD _0000_ _0085_ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_1471_ _0530_ _0450_ _0471_ core.ndc.col_out_n\[26\] VDD VSS VSS VDD sky130_fd_sc_hd__a21o_1
XFILLER_10_3 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_82_405 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_82_427 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_82_449 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1089__B1 _0506_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_50_346 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_50_357 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_1807_ core.osr.sample_count_r\[2\] net71 core.osr.next_sample_count_w\[2\] net57
+ VSS VDD VSS VDD sky130_fd_sc_hd__dfrtp_2
XFILLER_40_19 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1738_ core.cnb.average_sum_r\[3\] net61 core.cnb.next_average_sum_w\[3\] net76 VSS
+ VDD VSS VDD sky130_fd_sc_hd__dfrtp_1
X_1669_ VSS VDD _0183_ _0182_ _0185_ _0029_ VSS VDD sky130_fd_sc_hd__o21ai_1
XANTENNA_input7_A config_1_in[15] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_45_118 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_65_16 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_85_287 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_121_66 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_121_77 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_121_88 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1684__S _0616_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1735__CLK net76 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_39_50 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_49_424 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_91_202 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_91_213 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_0971_ core.cnb.shift_register_r\[5\] core.cnb.shift_register_r\[3\] _0291_ _0274_
+ _0397_ _0292_ VSS VDD VSS VDD sky130_fd_sc_hd__a2111oi_2
XANTENNA__0999__A _0353_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_58_3 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1523_ _0074_ _0082_ core.ndc.row_out_n\[12\] VSS VDD VSS VDD sky130_fd_sc_hd__or2_1
XFILLER_113_101 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_1454_ VSS VDD core.ndc.col_out_n\[12\] _0774_ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_1385_ VSS VDD _0734_ _0732_ core.osr.result_r\[12\] _0729_ VSS VDD sky130_fd_sc_hd__and3_1
XFILLER_55_449 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_82_246 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_129_9 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_4_8 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_104_123 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_116_22 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA_fanout65_A net67 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_132_21 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_46_449 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_132_76 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_30 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_92_69 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_74 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_63 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_41 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_52 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_96 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_85 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA_nmat_rowon_n[1] core.ndc.row_out_n\[2\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1443__A _0770_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1170_ VSS VDD core.cnb.nswitch_out\[11\] _0556_ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_0954_ _0379_ core.cnb.data_register_r\[6\] _0338_ _0380_ VDD VSS VSS VDD sky130_fd_sc_hd__a21o_1
X_0885_ core.cnb.shift_register_r\[10\] _0311_ core.cnb.shift_register_r\[11\] VSS
+ VDD VSS VDD sky130_fd_sc_hd__nor2_1
X_1506_ core.pdc.row_out_n\[14\] core.ndc.row_out_n\[2\] VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_4
XFILLER_87_305 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1437_ VSS VDD core.ndc.col_out_n\[1\] _0768_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_87_349 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_1368_ _0635_ _0720_ _0719_ _0718_ VSS VDD VSS VDD sky130_fd_sc_hd__o21ai_2
X_1299_ VSS VDD _0657_ core.cnb.result_out\[4\] _0656_ VSS VDD sky130_fd_sc_hd__xnor2_2
XANTENNA__1455__B1 _0514_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_62_39 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_51_441 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1528__A _0077_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_86_360 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_86_371 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1446__B1 _0506_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1202__S _0579_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_52_94 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xinput15 VSS VDD net15 config_1_in[8] VSS VDD sky130_fd_sc_hd__clkbuf_1
Xinput26 VSS VDD net26 config_2_in[3] VSS VDD sky130_fd_sc_hd__clkbuf_1
XANTENNA__1438__A _0353_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_96_102 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1222_ _0597_ core.cnb.next_data_register_w\[8\] _0588_ VSS VDD VSS VDD sky130_fd_sc_hd__nor2_1
XFILLER_84_319 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_1153_ core.cnb.shift_register_r\[12\] _0254_ _0252_ _0540_ _0255_ VDD VSS VSS VDD
+ sky130_fd_sc_hd__or4b_1
X_1084_ _0503_ _0376_ _0453_ _0454_ VSS VDD VSS VDD sky130_fd_sc_hd__o21a_1
XFILLER_92_385 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_52_249 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_93_90 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_0937_ VSS VDD _0362_ _0363_ _0358_ VSS VDD sky130_fd_sc_hd__xnor2_1
X_0868_ _0244_ _0261_ _0294_ _0268_ _0241_ VDD VSS VSS VDD sky130_fd_sc_hd__or4_2
X_0799_ core.osr.sample_count_r\[0\] _0226_ _0214_ VSS VDD VSS VDD sky130_fd_sc_hd__nor2_1
XFILLER_87_113 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_87_157 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1530__B core.ndc.row_out_n\[12\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XPHY_403 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_414 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_425 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_11_113 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_436 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_447 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_458 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_469 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1258__A core.cnb.comparator_in VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_138_53 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_22_97 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_138_97 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1692__S _0614_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_4_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_47_72 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_90_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_8_77 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_1771_ core.osr.result_r\[3\] net68 core.osr.next_result_w\[3\] net56 VSS VDD VSS
+ VDD sky130_fd_sc_hd__dfrtp_2
XFILLER_40_3 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1205_ _0579_ _0586_ VDD VSS VSS VDD sky130_fd_sc_hd__inv_2
X_1136_ _0533_ _0464_ _0374_ VSS VDD VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_81_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1067_ _0488_ _0435_ _0406_ VSS VDD VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_138_129 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_4_109 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_111_9 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_108_12 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_68_16 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_88_433 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_88_477 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_124_99 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_17_31 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_83_160 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_200 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_72_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XPHY_233 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_211 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_222 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_244 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_277 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_255 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_266 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_288 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_299 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_63_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1597__S core.osr.osr_mode_r\[0\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1754_ net44 net66 _0017_ net54 VSS VDD VSS VDD sky130_fd_sc_hd__dfrtp_1
X_1685_ VSS VDD _0036_ _0194_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_54_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1119_ VSS VDD _0512_ _0449_ _0513_ core.pdc.col_out_n\[20\] VSS VDD sky130_fd_sc_hd__o21ai_1
XFILLER_134_121 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1536__A core.ndc.row_out_n\[4\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_79_48 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_91_417 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_28_85 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_45_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_44_51 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_60_61 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_5_12 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1470_ _0424_ core.pdc.col_out_n\[24\] core.ndc.col_out_n\[25\] _0448_ VDD VSS VSS
+ VDD sky130_fd_sc_hd__a21oi_1
XFILLER_85_91 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1089__A1 _0424_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_36_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1806_ core.osr.sample_count_r\[1\] net71 core.osr.next_sample_count_w\[1\] net57
+ VSS VDD VSS VDD sky130_fd_sc_hd__dfrtp_2
X_1737_ core.cnb.average_sum_r\[2\] net61 core.cnb.next_average_sum_w\[2\] net76 VSS
+ VDD VSS VDD sky130_fd_sc_hd__dfrtp_1
XANTENNA__1356__A core.cnb.result_out\[9\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_131_113 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1668_ core.cnb.result_out\[10\] _0184_ _0185_ _0132_ VDD VSS VSS VDD sky130_fd_sc_hd__a21oi_1
X_1599_ core.osr.next_result_w\[1\] _0127_ core.osr.next_result_w\[7\] _0126_ _0123_
+ _0124_ VSS VDD VSS VDD sky130_fd_sc_hd__o221a_1
XFILLER_85_233 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_85_277 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_105_79 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_27_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_81_38 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_107_121 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_122_124 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_18_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_0970_ VSS VDD _0396_ _0385_ _0395_ VSS VDD sky130_fd_sc_hd__xnor2_2
X_1522_ core.ndc.row_out_n\[12\] _0556_ _0073_ VSS VDD VSS VDD sky130_fd_sc_hd__nand2_4
X_1453_ _0512_ _0774_ _0517_ VSS VDD VSS VDD sky130_fd_sc_hd__or2_1
X_1384_ core.osr.result_r\[12\] _0732_ _0733_ _0729_ VDD VSS VSS VDD sky130_fd_sc_hd__a21oi_1
XFILLER_27_108 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_50_111 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1234__A1 _0579_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_pmat_col_n[16] core.pdc.col_out_n\[16\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_116_78 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_46_406 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_25_20 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_20 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_31 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_64 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_42 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_53 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1473__A1 _0424_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XPHY_97 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_86 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_75 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA_nmat_rowon_n[0] core.ndc.row_out_n\[1\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_49_211 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_49_288 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_52_409 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_32_122 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1464__A1 _0424_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_0953_ _0300_ _0379_ _0337_ VSS VDD VSS VDD sky130_fd_sc_hd__nor2_1
X_0884_ _0309_ _0261_ _0310_ _0268_ _0242_ VDD VSS VSS VDD sky130_fd_sc_hd__or4_1
XANTENNA__0803__A core.osr.osr_mode_r\[0\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1075__S0 _0433_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1505_ VDD VSS core.pdc.row_out_n\[14\] _0076_ VSS VDD sky130_fd_sc_hd__buf_6
XFILLER_101_105 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_1436_ _0423_ _0459_ _0768_ VDD VSS VSS VDD sky130_fd_sc_hd__or2b_2
XFILLER_101_127 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1367_ VSS VDD _0719_ _0713_ _0717_ _0716_ VSS VDD sky130_fd_sc_hd__and3_1
XFILLER_46_19 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_55_225 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_1298_ _0655_ _0656_ _0212_ VSS VDD VSS VDD sky130_fd_sc_hd__nor2_1
XFILLER_102_25 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1455__A1 _0449_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_102_47 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_102_58 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_62_29 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_51_464 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1528__B core.ndc.row_out_n\[12\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_127_44 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_87_26 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1446__A1 _0354_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_36_85 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xinput16 VSS VDD net16 config_1_in[9] VSS VDD sky130_fd_sc_hd__clkbuf_1
Xinput27 VSS VDD net27 config_2_in[4] VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_96_125 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_1221_ VSS VDD _0586_ _0427_ _0343_ _0597_ VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_84_309 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1134__B1 _0471_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1152_ core.cnb.nswitch_out\[2\] core.cnb.pswitch_out\[2\] VDD VSS VSS VDD sky130_fd_sc_hd__inv_2
X_1083_ _0502_ core.pdc.col_out_n\[6\] _0501_ VSS VDD VSS VDD sky130_fd_sc_hd__nor2_1
XFILLER_92_397 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_20_103 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_0936_ VDD VSS _0362_ _0361_ _0359_ VSS VDD sky130_fd_sc_hd__and2_1
X_0867_ core.cnb.shift_register_r\[5\] core.cnb.data_register_r\[0\] core.cnb.shift_register_r\[3\]
+ _0293_ _0292_ VDD VSS VSS VDD sky130_fd_sc_hd__or4b_1
X_0798_ _0224_ core.osr.osr_mode_r\[0\] _0213_ _0225_ _0223_ VDD VSS VSS VDD sky130_fd_sc_hd__a211oi_2
XFILLER_87_125 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_1419_ VDD VSS _0757_ _0755_ core.osr.sample_count_r\[3\] VSS VDD sky130_fd_sc_hd__and2_1
XFILLER_87_169 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1676__A1 _0588_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XPHY_404 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_415 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_426 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_437 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_448 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_459 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_138_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_138_65 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_98_25 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_3 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_93_117 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_86_191 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_90_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1770_ core.osr.result_r\[2\] net67 core.osr.next_result_w\[2\] net55 VSS VDD VSS
+ VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_129_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_33_3 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_88_80 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_cgen_sample_n_in core.cnb.is_sampling_w VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1204_ VSS VDD core.cnb.next_data_register_w\[2\] _0585_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XANTENNA__1658__A1 core.cnb.result_out\[9\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1135_ _0529_ _0469_ core.pdc.col_out_n\[28\] _0465_ VDD VSS VSS VDD sky130_fd_sc_hd__a21oi_1
X_1066_ _0434_ _0348_ _0487_ _0349_ _0485_ VDD VSS VSS VDD sky130_fd_sc_hd__or4_1
XFILLER_81_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA_pmat_rowon_n[9] core.pdc.row_out_n\[10\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_0919_ _0345_ _0344_ _0343_ VSS VDD VSS VDD sky130_fd_sc_hd__xnor2_4
XFILLER_104_9 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1094__A _0449_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1525__C _0079_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_88_445 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_48_309 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_84_16 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_84_38 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1113__A3 _0468_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XPHY_201 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_72_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XPHY_212 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_234 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_223 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_245 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_256 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_267 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_33_64 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XPHY_278 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_289 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__0901__A core.cnb.data_register_r\[2\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_12_8 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_63_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1753_ net43 net66 _0016_ net55 VSS VDD VSS VDD sky130_fd_sc_hd__dfrtp_1
X_1684_ VSS VDD _0616_ core.cnb.shift_register_r\[6\] core.cnb.shift_register_r\[5\]
+ _0194_ VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_99_90 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_53_312 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_54_879 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_1118_ core.pdc.col_out_n\[19\] _0354_ _0514_ _0515_ VSS VDD VSS VDD sky130_fd_sc_hd__o21a_1
XFILLER_53_367 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1049_ _0470_ _0471_ _0462_ VSS VDD VSS VDD sky130_fd_sc_hd__nor2_2
XFILLER_110_25 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_70_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_0_113 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_88_253 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_48_128 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_28_42 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_28_97 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_91_429 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1698__S _0614_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_45_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_44_85 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_5_57 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_36_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_50_304 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_50_315 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA_pmat_sw_n core.cnb.enable_loop_out VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1805_ core.osr.sample_count_r\[0\] core.osr.next_sample_count_w\[0\] VDD net71 net57
+ VSS VSS VDD sky130_fd_sc_hd__dfstp_2
X_1736_ core.cnb.average_sum_r\[1\] net61 core.cnb.next_average_sum_w\[1\] net76 VSS
+ VDD VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_49_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_1667_ _0134_ net41 _0184_ _0104_ VSS VDD VSS VDD sky130_fd_sc_hd__and3b_1
XFILLER_131_125 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_1598_ _0232_ _0126_ _0125_ VSS VDD VSS VDD sky130_fd_sc_hd__or2_1
XFILLER_105_25 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_27_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_53_131 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_53_120 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_81_17 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_121_57 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_49_415 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1712__A0 net12 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_input20_A config_2_in[12] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_18_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_55_40 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1781__CLK net55 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_55_73 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_55_95 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1221__S _0586_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_72_7 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_1521_ VSS VDD _0081_ _0079_ net52 core.ndc.row_out_n\[11\] VSS VDD sky130_fd_sc_hd__o21ai_1
X_1452_ VSS VDD _0515_ _0449_ _0511_ core.ndc.col_out_n\[11\] VSS VDD sky130_fd_sc_hd__o21ai_1
X_1383_ core.osr.result_r\[13\] _0732_ VDD VSS VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_50_167 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1719_ core.cnb.data_register_r\[4\] net63 core.cnb.next_data_register_w\[4\] net80
+ VSS VDD VSS VDD sky130_fd_sc_hd__dfrtp_1
XANTENNA_pmat_col_n[15] core.pdc.col_out_n\[15\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__0929__A_N core.cnb.data_register_r\[2\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_132_34 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_46_429 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_10 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_21 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_54_462 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_65 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_54 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_32 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_43 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1473__A2 _0460_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_25_87 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_98 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_87 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_76 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_110_117 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1464__A2 _0515_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_0952_ VDD VSS _0378_ _0377_ _0331_ VSS VDD sky130_fd_sc_hd__and2_1
X_0883_ core.cnb.shift_register_r\[1\] core.cnb.shift_register_r\[2\] _0309_ core.cnb.shift_register_r\[3\]
+ core.cnb.is_sampling_w VDD VSS VSS VDD sky130_fd_sc_hd__or4_1
X_1504_ _0556_ _0076_ _0607_ _0073_ VDD VSS VSS VDD sky130_fd_sc_hd__or3_1
XFILLER_99_123 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1435_ _0456_ core.ndc.col_out_n\[0\] _0450_ VSS VDD VSS VDD sky130_fd_sc_hd__nor2_1
X_1366_ _0713_ _0717_ _0718_ _0716_ VDD VSS VSS VDD sky130_fd_sc_hd__a21oi_1
X_1297_ VSS VDD _0654_ _0655_ core.osr.result_r\[4\] VSS VDD sky130_fd_sc_hd__xnor2_1
XANTENNA__1455__A2 _0519_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_51_432 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_51_454 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1207__A2 _0586_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_fanout70_A net73 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_36_42 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_14_123 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xinput17 VSS VDD net17 config_2_in[0] VSS VDD sky130_fd_sc_hd__clkbuf_1
Xinput28 VSS VDD net28 config_2_in[5] VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_7_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_42_8 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1220_ VSS VDD core.cnb.next_data_register_w\[7\] _0596_ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_1151_ core.cnb.nswitch_out\[2\] _0539_ _0356_ VSS VDD VSS VDD sky130_fd_sc_hd__xnor2_4
XANTENNA__1134__A1 _0529_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1082_ _0458_ _0427_ _0502_ _0497_ VDD VSS VSS VDD sky130_fd_sc_hd__a21oi_1
XFILLER_93_70 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0814__A core.cnb.shift_register_r\[1\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_0935_ _0360_ _0361_ VDD VSS VSS VDD sky130_fd_sc_hd__inv_2
X_0866_ _0292_ core.cnb.shift_register_r\[7\] core.cnb.shift_register_r\[2\] core.cnb.shift_register_r\[6\]
+ VSS VDD VSS VDD sky130_fd_sc_hd__o21a_1
X_0797_ _0214_ core.osr.sample_count_r\[0\] _0224_ core.osr.sample_count_r\[8\] VSS
+ VDD VSS VDD sky130_fd_sc_hd__or3b_1
X_1418_ _0756_ core.osr.next_sample_count_w\[3\] core.osr.is_last_sample VSS VDD VSS
+ VDD sky130_fd_sc_hd__nor2_1
XANTENNA__1676__A2 _0615_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1349_ _0694_ _0635_ _0692_ _0693_ core.osr.result_r\[9\] _0702_ VSS VDD VSS VDD
+ sky130_fd_sc_hd__o2111ai_1
XFILLER_83_343 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_405 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_416 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_51_251 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_427 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_438 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_449 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_22_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_138_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_22_66 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_138_77 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1274__B _0635_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1290__A _0212_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_97_9 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_129_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1107__A1 _0374_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1203_ VDD VSS _0585_ _0584_ net53 VSS VDD sky130_fd_sc_hd__and2_1
XANTENNA__0866__B1 core.cnb.shift_register_r\[2\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1134_ _0529_ _0471_ core.pdc.col_out_n\[27\] _0473_ VDD VSS VSS VDD sky130_fd_sc_hd__a21oi_1
X_1065_ _0373_ _0486_ _0485_ VSS VDD VSS VDD sky130_fd_sc_hd__or2_1
XFILLER_138_109 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA_pmat_rowon_n[8] core.pdc.row_out_n\[9\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_0918_ VDD VSS _0344_ _0330_ VSS VDD sky130_fd_sc_hd__buf_6
X_0849_ _0275_ _0274_ _0273_ _0272_ _0271_ core.cnb.shift_register_r\[7\] VDD VSS
+ VSS VDD sky130_fd_sc_hd__o2111a_1
XANTENNA__1375__A core.cnb.result_out\[11\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_108_69 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1094__B _0466_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_88_457 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1649__A2 core.osr.next_result_w\[9\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XPHY_224 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_213 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_202 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_33_32 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_257 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_268 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_235 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_246 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_33_76 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_279 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1738__CLK net76 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_47_387 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_74_50 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_114_90 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1752_ net36 net66 _0015_ net55 VSS VDD VSS VDD sky130_fd_sc_hd__dfrtp_1
X_1683_ VSS VDD _0035_ _0193_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_85_427 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_85_449 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1117_ _0353_ _0463_ core.pdc.col_out_n\[18\] _0516_ _0524_ _0448_ VSS VDD VSS VDD
+ sky130_fd_sc_hd__a311o_1
XFILLER_53_357 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1048_ _0454_ _0376_ _0453_ _0470_ VDD VSS VSS VDD sky130_fd_sc_hd__a21o_1
XFILLER_79_28 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1319__A1 core.cnb.result_out\[4\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_0_125 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_88_221 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_95_16 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_95_49 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_28_65 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_100_70 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_125_101 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_5_69 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1804_ core.cnb.shift_register_r\[16\] net62 _0047_ net77 VSS VDD VSS VDD sky130_fd_sc_hd__dfrtp_2
X_1735_ core.cnb.average_sum_r\[0\] net61 core.cnb.next_average_sum_w\[0\] net76 VSS
+ VDD VSS VDD sky130_fd_sc_hd__dfrtp_1
X_1666_ VSS VDD core.osr.next_result_w\[12\] _0123_ _0115_ _0183_ VSS VDD sky130_fd_sc_hd__o21ai_1
X_1597_ VSS VDD core.osr.osr_mode_r\[0\] core.osr.next_result_w\[5\] core.osr.next_result_w\[3\]
+ _0125_ VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_105_48 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_53_143 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_81_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_14_89 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_30_55 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_input13_A config_1_in[6] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_91_238 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_55_63 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_65_7 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_1520_ VDD VSS _0352_ _0081_ _0607_ VSS VDD sky130_fd_sc_hd__and2_2
X_1451_ _0773_ _0513_ _0507_ _0448_ core.ndc.col_out_n\[10\] VSS VDD VSS VDD sky130_fd_sc_hd__o211a_1
X_1382_ VDD VSS _0731_ core.osr.next_result_w\[12\] VSS VDD sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_55_408 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_50_157 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_1718_ core.cnb.data_register_r\[3\] net74 core.cnb.next_data_register_w\[3\] net81
+ VSS VDD VSS VDD sky130_fd_sc_hd__dfrtp_1
X_1649_ core.osr.next_result_w\[9\] _0169_ core.osr.next_result_w\[15\] _0168_ _0123_
+ _0124_ VSS VDD VSS VDD sky130_fd_sc_hd__o221a_1
XANTENNA_input5_A config_1_in[13] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_54_430 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_22 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_25_44 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XPHY_55 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_33 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_44 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_88 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_77 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_66 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_25_99 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XPHY_99 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_2_15 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_49_268 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_66_51 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_66_62 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_0951_ VSS VDD _0318_ _0330_ core.cnb.data_register_r\[5\] _0377_ VSS VDD sky130_fd_sc_hd__o21ai_1
XANTENNA__1621__B1 core.osr.next_result_w\[10\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_0882_ core.cnb.shift_register_r\[4\] _0308_ core.cnb.shift_register_r\[5\] VSS VDD
+ VSS VDD sky130_fd_sc_hd__or2_1
XFILLER_56_3 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1503_ VSS VDD core.ndc.row_out_n\[1\] _0075_ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_1434_ _0767_ core.osr.next_sample_count_w\[8\] core.osr.is_last_sample VSS VDD VSS
+ VDD sky130_fd_sc_hd__nor2_1
X_1365_ core.osr.result_r\[10\] _0717_ VDD VSS VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_55_205 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_1296_ _0654_ _0653_ _0651_ VSS VDD VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_23_113 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_51_422 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_23_124 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_51_477 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1097__B _0472_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_11_57 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_127_57 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1771__CLK net56 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_fanout63_A net74 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_46_249 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_86_396 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_36_76 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_36_65 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_36_98 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_52_20 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xinput18 VSS VDD net18 config_2_in[10] VSS VDD sky130_fd_sc_hd__clkbuf_1
Xinput29 VSS VDD net29 config_2_in[6] VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_7_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_96_116 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_28_7 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1150_ _0539_ _0327_ _0355_ VSS VDD VSS VDD sky130_fd_sc_hd__nand2_2
XFILLER_77_83 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1081_ VDD VSS _0501_ _0500_ _0499_ VSS VDD sky130_fd_sc_hd__and2_1
XFILLER_92_344 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_93_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__0814__B core.cnb.is_sampling_w VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_20_116 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1794__CLK net77 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_0934_ _0334_ _0360_ _0307_ VSS VDD VSS VDD sky130_fd_sc_hd__nor2_1
X_0865_ _0291_ core.cnb.shift_register_r\[6\] core.cnb.shift_register_r\[7\] VSS VDD
+ VSS VDD sky130_fd_sc_hd__xnor2_4
XANTENNA__1070__A1 _0433_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_0796_ core.osr.sample_count_r\[0\] core.osr.osr_mode_r\[2\] _0223_ _0222_ VSS VDD
+ VSS VDD sky130_fd_sc_hd__or3b_1
X_1417_ VSS VDD _0755_ _0756_ core.osr.sample_count_r\[3\] VSS VDD sky130_fd_sc_hd__xnor2_1
XFILLER_87_138 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1348_ VSS VDD _0701_ _0700_ _0682_ _0699_ _0694_ VSS VDD sky130_fd_sc_hd__a211o_1
XFILLER_84_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1279_ VSS VDD _0639_ core.osr.next_result_w\[1\] core.cnb.result_out\[1\] VSS VDD
+ sky130_fd_sc_hd__xnor2_1
XFILLER_83_388 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_51_230 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_406 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_417 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_11_105 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_51_241 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1600__S _0235_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XPHY_428 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_439 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1349__C1 _0635_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1364__A2 core.cnb.result_out\[9\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_93_108 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_47_86 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_75_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_103_70 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1052__A1 _0424_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1107__A2 _0468_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1202_ VSS VDD _0579_ core.cnb.data_register_r\[2\] core.cnb.nswitch_out\[2\] _0584_
+ VSS VDD sky130_fd_sc_hd__mux2_1
XANTENNA__0809__B _0235_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1133_ VSS VDD core.pdc.col_out_n\[26\] _0448_ _0531_ _0353_ _0532_ VSS VDD sky130_fd_sc_hd__a211o_1
XFILLER_66_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_92_141 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_1064_ _0444_ _0485_ _0438_ VSS VDD VSS VDD sky130_fd_sc_hd__or2_1
X_0917_ _0343_ core.cnb.data_register_r\[8\] VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_2
X_0848_ core.cnb.shift_register_r\[2\] _0274_ VDD VSS VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_108_48 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_108_59 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_88_403 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_88_469 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_84_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_57_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XPHY_225 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_203 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_214 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_33_11 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_236 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_247 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_258 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_269 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_3_123 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_47_344 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_48_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1476__A core.cnb.shift_register_r\[1\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1751_ core.cnb.result_out\[11\] net64 _0014_ net79 VSS VDD VSS VDD sky130_fd_sc_hd__dfrtp_4
X_1682_ VSS VDD _0568_ core.cnb.shift_register_r\[5\] core.cnb.shift_register_r\[4\]
+ _0193_ VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_85_417 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_39_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1116_ VDD VSS _0524_ _0394_ _0351_ VSS VDD sky130_fd_sc_hd__and2_1
XFILLER_0_81 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_1047_ _0354_ _0469_ core.pdc.col_out_n\[3\] _0465_ VDD VSS VSS VDD sky130_fd_sc_hd__a21oi_1
XFILLER_110_49 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1016__A1 _0433_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_88_233 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_135_57 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_28_33 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_60_42 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1296__A _0651_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_100_93 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_125_113 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_69_40 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_50_339 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1803_ core.cnb.shift_register_r\[15\] net63 _0046_ net77 VSS VDD VSS VDD sky130_fd_sc_hd__dfrtp_1
X_1734_ core.cnb.average_counter_r\[4\] net60 core.cnb.next_average_counter_w\[4\]
+ net75 VSS VDD VSS VDD sky130_fd_sc_hd__dfrtp_1
XANTENNA_pmat_col_n[30] core.pdc.col_out_n\[30\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1665_ _0182_ _0736_ _0111_ _0749_ _0181_ _0123_ VSS VDD VSS VDD sky130_fd_sc_hd__o311a_1
X_1596_ VDD VSS _0124_ _0105_ VSS VDD sky130_fd_sc_hd__buf_2
XFILLER_85_214 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_85_225 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_53_155 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_121_37 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_107_113 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_30_89 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_30_67 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_49_406 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_39_87 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__0920__B1 _0345_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_111_81 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_1450_ _0773_ _0474_ _0529_ VSS VDD VSS VDD sky130_fd_sc_hd__nand2_1
X_1381_ _0731_ core.osr.result_r\[12\] _0730_ _0729_ VSS VDD VSS VDD sky130_fd_sc_hd__o21a_1
XFILLER_96_71 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_96_93 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_110_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_50_125 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_90_294 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1717_ core.cnb.data_register_r\[2\] net68 core.cnb.next_data_register_w\[2\] net81
+ VSS VDD VSS VDD sky130_fd_sc_hd__dfrtp_4
XANTENNA_nmat_rowon_n[11] core.ndc.row_out_n\[12\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_pmat_col_n[13] core.pdc.col_out_n\[13\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1648_ core.osr.next_result_w\[13\] _0168_ _0154_ _0134_ _0230_ core.osr.next_result_w\[11\]
+ VSS VDD VSS VDD sky130_fd_sc_hd__o221a_1
X_1579_ VDD VSS _0109_ _0104_ net43 VSS VDD sky130_fd_sc_hd__and2_1
XFILLER_101_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1603__S _0110_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1458__A1 _0529_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_26_122 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_12 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_54_442 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_92_29 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_56 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_23 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_34 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_45 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_89 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_78 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_67 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1146__B1 core.cnb.data_register_r\[1\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_49_225 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_0950_ _0376_ _0375_ VSS VDD VSS VDD sky130_fd_sc_hd__clkbuf_4
X_0881_ core.cnb.data_register_r\[3\] _0307_ VDD VSS VSS VDD sky130_fd_sc_hd__inv_2
X_1502_ VDD VSS _0075_ _0074_ core.ndc.row_out_n\[4\] VSS VDD sky130_fd_sc_hd__and2_1
XFILLER_99_103 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1433_ _0766_ _0767_ core.osr.sample_count_r\[8\] VDD VSS VSS VDD sky130_fd_sc_hd__xor2_1
XFILLER_49_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_1364_ core.cnb.result_out\[9\] _0716_ _0680_ _0715_ core.osr.result_r\[9\] _0712_
+ VSS VDD VSS VDD sky130_fd_sc_hd__o221a_1
X_1295_ _0652_ core.osr.result_r\[3\] core.cnb.result_out\[3\] _0653_ VSS VDD VSS
+ VDD sky130_fd_sc_hd__a21oi_4
XFILLER_55_217 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1378__B core.cnb.result_out\[11\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_11_69 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_46_217 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_36_33 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA_fanout56_A core.cnb.conv_finished_r VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_54_294 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_52_76 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1603__A1 core.osr.next_result_w\[6\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xinput19 VSS VDD net19 config_2_in[11] VSS VDD sky130_fd_sc_hd__clkbuf_1
XANTENNA__1119__B1 _0513_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_77_62 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1080_ _0454_ _0463_ _0500_ _0455_ VDD VSS VSS VDD sky130_fd_sc_hd__a21oi_1
XFILLER_92_356 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_93_879 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_0933_ VDD VSS _0359_ _0335_ VSS VDD sky130_fd_sc_hd__buf_2
X_0864_ _0290_ _0285_ _0289_ _0287_ core.cnb.data_register_r\[0\] _0282_ VSS VDD VSS
+ VDD sky130_fd_sc_hd__a32o_1
X_0795_ core.osr.sample_count_r\[8\] _0222_ VDD VSS VSS VDD sky130_fd_sc_hd__inv_2
XANTENNA__1358__B1 core.cnb.result_out\[9\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1416_ VSS VDD _0755_ core.osr.sample_count_r\[1\] core.osr.sample_count_r\[0\] core.osr.sample_count_r\[2\]
+ VSS VDD sky130_fd_sc_hd__and3_1
XFILLER_3_81 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1347_ _0693_ _0700_ core.osr.result_r\[9\] _0212_ VDD VSS VSS VDD sky130_fd_sc_hd__or3_1
XFILLER_84_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1278_ _0639_ _0638_ _0635_ VSS VDD VSS VDD sky130_fd_sc_hd__nand2_1
XPHY_407 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_418 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_429 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_11_128 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_51_275 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_98_17 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1521__B1 net52 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_47_32 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_47_65 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_75_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_63_42 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1299__A core.cnb.result_out\[4\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_8_15 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__0931__A core.cnb.data_register_r\[2\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1052__A2 _0471_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_6_121 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1238__S _0586_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1201_ VSS VDD core.cnb.next_data_register_w\[1\] _0583_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XANTENNA__1512__B1 net52 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1132_ _0532_ _0454_ _0458_ _0455_ VSS VDD VSS VDD sky130_fd_sc_hd__o21a_1
XFILLER_66_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_92_131 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1063_ _0373_ _0481_ _0484_ _0433_ _0482_ _0479_ _0483_ VSS VDD VSS VDD sky130_fd_sc_hd__mux4_1
XFILLER_92_175 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0841__A core.cnb.data_register_r\[2\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_0916_ _0341_ _0336_ _0306_ _0333_ _0342_ VDD VSS VSS VDD sky130_fd_sc_hd__o211a_2
X_0847_ core.cnb.shift_register_r\[6\] _0273_ VDD VSS VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_124_37 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_124_15 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_124_48 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_57_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_83_142 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_83_153 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_17_57 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XPHY_204 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_215 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_237 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_248 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_226 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_259 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_33_89 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_116_3 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_3_113 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_48_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_88_7 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1750_ core.cnb.result_out\[10\] net64 _0013_ net79 VSS VDD VSS VDD sky130_fd_sc_hd__dfrtp_4
XANTENNA__1476__B _0614_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1681_ VSS VDD _0034_ _0192_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_99_71 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_nmat_analog_in inn_analog VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_39_879 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_1115_ VSS VDD core.pdc.col_out_n\[17\] _0523_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_53_337 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_53_348 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1046_ _0468_ _0469_ _0466_ VSS VDD VSS VDD sky130_fd_sc_hd__nor2_1
XFILLER_119_15 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_119_122 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_119_37 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_135_69 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_95_29 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_48_109 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_84_473 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_44_66 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_60_21 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_60_76 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_125_125 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_90_421 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1802_ core.cnb.shift_register_r\[14\] net63 _0045_ net80 VSS VDD VSS VDD sky130_fd_sc_hd__dfrtp_1
X_1733_ core.cnb.average_counter_r\[3\] net60 core.cnb.next_average_counter_w\[3\]
+ net75 VSS VDD VSS VDD sky130_fd_sc_hd__dfrtp_2
XFILLER_116_103 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1664_ _0738_ _0216_ _0180_ _0181_ VDD VSS VSS VDD sky130_fd_sc_hd__a21o_1
X_1595_ VDD VSS _0123_ _0219_ VSS VDD sky130_fd_sc_hd__buf_2
X_1029_ _0420_ _0454_ VSS VDD VSS VDD sky130_fd_sc_hd__clkbuf_2
XFILLER_122_106 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_39_44 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0920__A1 _0328_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_71_20 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_71_53 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_1380_ core.osr.result_r\[12\] _0212_ _0730_ _0729_ VDD VSS VSS VDD sky130_fd_sc_hd__a21oi_1
XFILLER_82_207 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_110_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_82_229 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_50_137 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1010__A _0347_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1716_ core.cnb.data_register_r\[1\] net67 core.cnb.next_data_register_w\[1\] net79
+ VSS VDD VSS VDD sky130_fd_sc_hd__dfrtp_2
X_1647_ _0134_ net38 _0167_ _0104_ VSS VDD VSS VDD sky130_fd_sc_hd__and3b_1
XFILLER_104_117 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_116_16 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1578_ VSS VDD _0015_ _0108_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_101_879 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1458__A2 _0520_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_54_421 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_13 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_41_104 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_24 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_35 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_46 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_25_57 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XPHY_79 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_68 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_57 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_41_34 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_89_384 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1590__A _0110_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_49_259 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_17_123 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_122_81 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1082__B1 _0427_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1621__A2 core.osr.next_result_w\[8\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_0880_ core.cnb.data_register_r\[6\] _0300_ _0306_ core.cnb.data_register_r\[7\]
+ _0305_ VDD VSS VSS VDD sky130_fd_sc_hd__a22o_2
XANTENNA__1718__CLK net81 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1501_ _0074_ _0352_ _0607_ VSS VDD VSS VDD sky130_fd_sc_hd__nor2_4
X_1432_ _0766_ _0764_ core.osr.sample_count_r\[7\] VSS VDD VSS VDD sky130_fd_sc_hd__nand2_1
XANTENNA__1137__A1 _0354_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1704__S _0614_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1363_ _0715_ core.osr.result_r\[9\] core.osr.result_r\[8\] core.cnb.result_out\[9\]
+ core.cnb.result_out\[8\] VSS VDD _0714_ VSS VDD sky130_fd_sc_hd__a221o_1
X_1294_ core.osr.result_r\[2\] core.cnb.result_out\[2\] core.osr.result_r\[3\] core.cnb.result_out\[3\]
+ _0652_ VSS VDD VSS VDD sky130_fd_sc_hd__o211a_1
XFILLER_48_270 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1005__A _0364_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_102_29 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_11_15 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_127_26 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1128__A1 _0352_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_86_365 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1585__A _0235_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1119__A1 _0449_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_77_74 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_93_40 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_92_379 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_0932_ _0355_ _0357_ _0358_ _0356_ VDD VSS VSS VDD sky130_fd_sc_hd__a21oi_1
X_0863_ _0288_ _0240_ _0289_ _0242_ _0239_ VSS VDD VSS VDD sky130_fd_sc_hd__nor4_4
X_0794_ VSS VDD core.osr.sample_count_r\[2\] _0220_ _0218_ _0221_ VSS VDD sky130_fd_sc_hd__mux2_1
X_1415_ _0754_ core.osr.next_sample_count_w\[2\] core.osr.is_last_sample VSS VDD VSS
+ VDD sky130_fd_sc_hd__nor2_1
X_1346_ _0692_ _0699_ core.osr.result_r\[9\] _0212_ VDD VSS VSS VDD sky130_fd_sc_hd__or3_1
XFILLER_3_93 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_83_302 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_113_28 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1277_ VSS VDD _0637_ _0638_ core.osr.result_r\[1\] VSS VDD sky130_fd_sc_hd__xnor2_1
XPHY_408 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_419 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_132_9 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_22_25 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1597__A1 core.osr.next_result_w\[5\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_98_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1521__A1 _0079_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_103_83 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_63_65 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_63_76 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_88_51 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1200_ VDD VSS _0583_ _0582_ net53 VSS VDD sky130_fd_sc_hd__and2_1
XANTENNA__1512__A1 _0079_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1131_ VDD VSS _0531_ _0452_ _0352_ VSS VDD sky130_fd_sc_hd__and2_1
X_1062_ _0345_ _0483_ _0480_ _0406_ VDD VSS VSS VDD sky130_fd_sc_hd__or3_1
XFILLER_92_187 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_pmat_rowon_n[5] core.pdc.row_out_n\[6\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_0915_ _0340_ _0341_ _0300_ VSS VDD VSS VDD sky130_fd_sc_hd__or2_1
X_0846_ VSS VDD core.cnb.shift_register_r\[5\] core.cnb.shift_register_r\[3\] core.cnb.shift_register_r\[7\]
+ _0272_ VSS VDD sky130_fd_sc_hd__o21ai_1
XFILLER_17_14 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1329_ VSS VDD _0684_ _0653_ _0667_ _0651_ _0683_ VSS VDD sky130_fd_sc_hd__a211o_1
XFILLER_17_69 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_83_176 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_216 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_205 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_249 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_227 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_238 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_33_46 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_109_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xcgen clk_comp_cgen core.clk_dig_in net17 net24 net25 net26 net27 net28 net29 net30
+ net31 net32 net18 net19 net20 net21 net22 net2 net3 net4 net5 net6 net7 net53 net23
+ decision_finish_comp_n core.cnb.enable_loop_out sample_nmatrix_cgen_n core.cnb.enable_loop_out
+ sample_pmatrix_cgen_n core.cnb.is_sampling_w sample_nmatrix_cgen core.cnb.is_sampling_w
+ sample_pmatrix_cgen net34 VDD VSS adc_clkgen_with_edgedetect
XFILLER_47_313 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA_input29_A config_2_in[6] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_47_368 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_95_9 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1680_ VSS VDD _0568_ core.cnb.shift_register_r\[4\] core.cnb.shift_register_r\[3\]
+ _0192_ VSS VDD sky130_fd_sc_hd__mux2_1
XANTENNA__1712__S _0635_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1114_ _0521_ _0353_ _0523_ _0519_ VSS VDD VSS VDD sky130_fd_sc_hd__o21ba_1
XANTENNA__1013__A _0345_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1045_ VDD VSS _0468_ _0467_ VSS VDD sky130_fd_sc_hd__buf_2
XFILLER_110_29 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_9_81 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_0829_ VDD VSS _0255_ core.cnb.shift_register_r\[14\] VSS VDD sky130_fd_sc_hd__buf_2
XFILLER_135_15 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_88_268 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_84_441 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_44_45 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1007__A3 _0427_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_69_64 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_47_121 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_47_176 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_90_400 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_90_433 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_90_477 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_1801_ core.cnb.shift_register_r\[13\] net63 _0044_ net80 VSS VDD VSS VDD sky130_fd_sc_hd__dfrtp_1
X_1732_ core.cnb.average_counter_r\[2\] net60 core.cnb.next_average_counter_w\[2\]
+ net75 VSS VDD VSS VDD sky130_fd_sc_hd__dfrtp_1
X_1663_ _0635_ _0111_ _0743_ _0216_ _0742_ _0180_ VSS VDD VSS VDD sky130_fd_sc_hd__o2111ai_1
XANTENNA__1706__A1 _0588_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1594_ VDD VSS _0122_ _0104_ net45 VSS VDD sky130_fd_sc_hd__and2_1
XFILLER_53_113 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1028_ VDD VSS _0453_ _0410_ VSS VDD sky130_fd_sc_hd__buf_2
XFILLER_14_48 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1774__CLK net56 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_122_118 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_39_34 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_29_121 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0920__A2 _0342_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_84_293 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_111_72 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1633__B1 core.osr.next_result_w\[10\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1164__A2 _0328_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_48_463 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_35_124 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_90_241 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1797__CLK net76 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_50_149 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_91_3 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1010__B _0366_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1715_ core.cnb.data_register_r\[0\] net64 core.cnb.next_data_register_w\[0\] net78
+ VSS VDD VSS VDD sky130_fd_sc_hd__dfrtp_4
XFILLER_104_107 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_1646_ VSS VDD _0163_ _0164_ _0115_ _0025_ _0166_ _0123_ VSS VDD sky130_fd_sc_hd__a41o_1
X_1577_ VDD VSS _0108_ _0107_ _0104_ VSS VDD sky130_fd_sc_hd__and2_1
XFILLER_25_14 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_14 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_25 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_36 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_47 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_54_477 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_25_69 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_69 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_58 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1091__A1 _0353_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_49_205 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_2_29 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_49_238 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_106_61 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_106_72 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_49_249 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_66_21 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA_input11_A config_1_in[4] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_82_42 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_82_64 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1500_ core.ndc.row_out_n\[4\] _0556_ _0073_ VSS VDD VSS VDD sky130_fd_sc_hd__nor2_4
X_1431_ _0765_ core.osr.next_sample_count_w\[7\] core.osr.is_last_sample VSS VDD VSS
+ VDD sky130_fd_sc_hd__nor2_1
XANTENNA__1137__A2 _0460_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1362_ core.osr.result_r\[7\] _0714_ core.osr.result_r\[8\] core.cnb.result_out\[7\]
+ core.cnb.result_out\[8\] VSS VDD VSS VDD sky130_fd_sc_hd__o22a_1
X_1293_ _0650_ _0642_ _0651_ _0641_ VSS VDD VSS VDD sky130_fd_sc_hd__a21bo_2
XFILLER_96_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_20_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_11_27 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1629_ VSS VDD core.cnb.result_out\[3\] _0235_ _0152_ _0153_ _0132_ VSS VDD sky130_fd_sc_hd__a2bb2o_1
XANTENNA_input3_A config_1_in[11] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_86_300 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_86_344 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_86_333 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_87_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_46_208 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_11_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA_cgen_ena_in net53 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1119__A2 _0512_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_77_53 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_78_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_92_314 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_0931_ VDD VSS _0357_ _0266_ core.cnb.data_register_r\[2\] VSS VDD sky130_fd_sc_hd__and2_1
X_0862_ core.cnb.shift_register_r\[11\] _0288_ core.cnb.shift_register_r\[10\] core.cnb.shift_register_r\[16\]
+ VDD VSS VSS VDD sky130_fd_sc_hd__or3_1
X_0793_ core.osr.sample_count_r\[4\] _0220_ _0219_ VSS VDD VSS VDD sky130_fd_sc_hd__or2_1
XFILLER_54_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1358__A2 core.cnb.result_out\[8\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1414_ _0753_ _0754_ core.osr.sample_count_r\[2\] VDD VSS VSS VDD sky130_fd_sc_hd__xor2_1
XFILLER_69_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1345_ core.osr.next_result_w\[8\] _0698_ _0692_ VSS VDD VSS VDD sky130_fd_sc_hd__xnor2_4
X_1276_ _0637_ core.cnb.result_out\[0\] core.osr.result_r\[0\] VSS VDD VSS VDD sky130_fd_sc_hd__nand2_1
XANTENNA__0855__A core.cnb.data_register_r\[1\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XPHY_409 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_11_119 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_51_266 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_51_288 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_138_15 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_125_9 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_22_37 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_22_59 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1625__S _0110_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1521__A2 _0081_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_86_152 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_86_163 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_63_88 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1512__A2 _0080_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1130_ _0501_ _0530_ _0529_ core.pdc.col_out_n\[25\] VSS VDD VSS VDD sky130_fd_sc_hd__a21oi_2
X_1061_ _0347_ _0482_ _0478_ _0406_ VDD VSS VSS VDD sky130_fd_sc_hd__or3_1
Xnmat_101 nmat_101/LO net101 VDD VSS VSS VDD sky130_fd_sc_hd__conb_1
X_0914_ _0340_ _0337_ _0339_ core.cnb.data_register_r\[6\] _0338_ VSS VDD VSS VDD
+ sky130_fd_sc_hd__o31a_1
X_0845_ core.cnb.shift_register_r\[5\] _0271_ core.cnb.shift_register_r\[3\] VDD VSS
+ VSS VDD sky130_fd_sc_hd__xor2_1
XANTENNA__1784__RESET_B net73 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_88_417 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_1328_ _0683_ core.osr.result_r\[7\] core.osr.result_r\[6\] VSS VDD VSS VDD sky130_fd_sc_hd__nand2_1
X_1259_ _0625_ core.cnb.average_sum_r\[0\] core.cnb.comparator_in VSS VDD VSS VDD
+ sky130_fd_sc_hd__nand2_1
XFILLER_17_26 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_206 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_33_25 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_228 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_217 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_239 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_137_113 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_87_461 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_47_358 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_74_21 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1663__D1 _0635_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_128_102 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_99_84 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0941__B1 core.cnb.data_register_r\[2\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_85_409 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1113_ core.pdc.col_out_n\[16\] _0376_ _0462_ _0352_ _0468_ VSS VDD VSS VDD sky130_fd_sc_hd__o31a_1
XFILLER_53_328 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1044_ _0410_ _0467_ _0420_ VSS VDD VSS VDD sky130_fd_sc_hd__or2_1
XANTENNA__1013__B _0366_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_9_93 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_119_28 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_0828_ VDD VSS _0254_ core.cnb.shift_register_r\[15\] VSS VDD sky130_fd_sc_hd__buf_2
XFILLER_135_27 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_131_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_28_25 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1488__A1 _0433_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_84_453 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_52_372 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_121_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_69_21 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_122_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_47_144 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_85_64 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_47_188 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_47_199 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_90_445 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1100__B1 _0466_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1800_ core.cnb.shift_register_r\[12\] net63 _0043_ net80 VSS VDD VSS VDD sky130_fd_sc_hd__dfrtp_4
X_1731_ core.cnb.average_counter_r\[1\] net60 core.cnb.next_average_counter_w\[1\]
+ net75 VSS VDD VSS VDD sky130_fd_sc_hd__dfrtp_1
X_1662_ VSS VDD _0028_ _0179_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_116_127 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1593_ VSS VDD _0017_ _0121_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_113_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1024__A _0427_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_121_29 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_53_169 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1027_ _0451_ _0452_ VSS VDD VSS VDD sky130_fd_sc_hd__clkbuf_2
XFILLER_107_127 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_104_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_39_57 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_39_68 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_71_88 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1109__A _0466_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1543__S _0588_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__0948__A _0366_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1164__A3 _0342_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_96_41 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_96_85 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_48_431 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_48_442 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_48_453 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_90_253 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_1714_ core.cnb.conv_finished_r net64 core.cnb.next_conv_finished_w net78 VSS VDD
+ VSS VDD sky130_fd_sc_hd__dfrtp_1
XANTENNA_pmat_col_n[10] core.pdc.col_out_n\[10\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1645_ _0115_ _0165_ _0112_ core.osr.next_result_w\[8\] _0166_ VSS VDD VSS VDD sky130_fd_sc_hd__a31o_1
X_1576_ VSS VDD _0235_ _0106_ net36 _0107_ VSS VDD sky130_fd_sc_hd__mux2_1
XPHY_15 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_26 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_37 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_59 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_48 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1615__A1 core.osr.next_result_w\[9\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_41_25 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_66_33 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_122_94 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_99_117 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1430_ VSS VDD _0764_ _0765_ core.osr.sample_count_r\[7\] VSS VDD sky130_fd_sc_hd__xnor2_1
X_1361_ VSS VDD _0668_ _0713_ _0712_ core.cnb.result_out\[6\] core.osr.result_r\[6\]
+ _0670_ VSS VDD sky130_fd_sc_hd__a2111o_1
X_1292_ core.osr.result_r\[2\] _0650_ core.cnb.result_out\[3\] core.cnb.result_out\[2\]
+ core.osr.result_r\[3\] VSS VDD VSS VDD sky130_fd_sc_hd__o22a_1
XFILLER_96_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1302__A core.cnb.result_out\[4\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_20_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_11_39 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1628_ _0152_ _0104_ net49 VSS VDD VSS VDD sky130_fd_sc_hd__nand2_1
X_1559_ VSS VDD _0089_ core.cnb.next_data_register_w\[6\] core.cnb.result_out\[6\]
+ _0096_ VSS VDD sky130_fd_sc_hd__mux2_1
XANTENNA__1533__B1 net52 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_87_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_54_286 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_54_264 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_50_481 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_11_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_77_21 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_96_109 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_117_94 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_78_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_92_326 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_92_337 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_0930_ _0296_ _0356_ _0281_ _0297_ VDD VSS VSS VDD sky130_fd_sc_hd__and3_2
X_0861_ VDD VSS _0287_ _0286_ core.cnb.data_register_r\[0\] VSS VDD sky130_fd_sc_hd__and2_1
X_0792_ core.osr.osr_mode_r\[1\] _0216_ _0219_ core.osr.osr_mode_r\[2\] VSS VDD VSS
+ VDD sky130_fd_sc_hd__or3_2
X_1413_ _0753_ core.osr.sample_count_r\[1\] core.osr.sample_count_r\[0\] VSS VDD VSS
+ VDD sky130_fd_sc_hd__nand2_1
XFILLER_3_51 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_69_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1344_ _0212_ _0697_ _0696_ _0698_ VSS VDD VSS VDD sky130_fd_sc_hd__a21oi_2
X_1275_ VSS VDD _0636_ core.osr.next_result_w\[0\] core.cnb.result_out\[0\] VSS VDD
+ sky130_fd_sc_hd__xnor2_1
XFILLER_83_337 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_22_49 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_86_197 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1641__S _0110_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_fanout54_A net55 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_103_30 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_103_96 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_8_29 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1551__S _0089_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_92_123 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1060_ _0347_ _0481_ _0480_ _0406_ VDD VSS VSS VDD sky130_fd_sc_hd__or3_1
X_0913_ _0304_ core.cnb.data_register_r\[7\] core.cnb.data_register_r\[6\] _0319_
+ _0339_ VSS VDD VSS VDD sky130_fd_sc_hd__a31o_1
X_0844_ _0242_ _0269_ _0270_ _0261_ _0268_ VSS VDD VSS VDD sky130_fd_sc_hd__nor4_2
XFILLER_124_29 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_83_123 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1327_ _0679_ _0675_ _0682_ _0677_ _0681_ VDD VSS VSS VDD sky130_fd_sc_hd__or4b_2
X_1258_ VSS VDD _0624_ core.cnb.next_average_sum_w\[0\] core.cnb.comparator_in VSS
+ VDD sky130_fd_sc_hd__xnor2_1
X_1189_ VSS VDD core.cnb.sampled_avg_control_r\[0\] core.cnb.average_sum_r\[3\] core.cnb.average_sum_r\[2\]
+ _0573_ VSS VDD sky130_fd_sc_hd__mux2_1
XPHY_207 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_229 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_218 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_137_125 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_3_105 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1636__S _0110_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_58_56 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_0_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_47_304 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_87_473 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_74_11 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_74_33 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_74_44 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_130_50 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_90_43 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_90_54 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_90_76 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_139_81 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_99_41 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_1112_ core.pdc.col_out_n\[15\] _0376_ _0474_ _0449_ _0468_ VSS VDD VSS VDD sky130_fd_sc_hd__o31a_1
XFILLER_0_41 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1043_ VDD VSS _0466_ _0462_ VSS VDD sky130_fd_sc_hd__buf_2
XFILLER_0_85 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1310__A core.cnb.result_out\[4\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_9_50 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_0827_ _0252_ _0253_ VDD VSS VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_88_215 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_135_39 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_131_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_84_410 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_28_59 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_84_465 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_52_340 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_5_19 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_109_51 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_122_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA_input34_A start_conversion_in VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_87_281 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_47_156 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_90_457 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_93_8 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_1730_ core.cnb.next_average_counter_w\[0\] VDD core.cnb.average_counter_r\[0\] net60
+ net75 VSS VSS VDD sky130_fd_sc_hd__dfstp_1
X_1661_ _0176_ _0179_ _0178_ VSS VDD VSS VDD sky130_fd_sc_hd__or2_1
X_1592_ VSS VDD _0115_ _0120_ _0117_ _0121_ VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_113_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_53_104 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1026_ _0394_ _0451_ _0410_ VSS VDD VSS VDD sky130_fd_sc_hd__or2_1
XFILLER_104_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_84_240 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_44_104 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_55_57 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_52_170 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1633__A2 core.osr.next_result_w\[6\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1109__B _0520_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_113_109 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__0948__B _0373_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1125__A _0528_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_35_104 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_90_221 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_90_232 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XPHY_390 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_1713_ VSS VDD _0050_ _0208_ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_1644_ core.cnb.result_out\[6\] _0209_ _0165_ net37 _0236_ VDD VSS VSS VDD sky130_fd_sc_hd__a22o_1
X_1575_ _0105_ _0106_ _0657_ VSS VDD VSS VDD sky130_fd_sc_hd__nor2_1
XANTENNA__1312__A1 _0651_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XPHY_16 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_27 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_38 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_54_468 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_49 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_1009_ _0370_ _0434_ _0359_ _0372_ VDD VSS VSS VDD sky130_fd_sc_hd__and3_2
XFILLER_49_218 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_106_41 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_106_96 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_17_104 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_122_51 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_82_33 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_82_77 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA_vcm_clk clk_vcm VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1360_ core.cnb.result_out\[7\] core.osr.result_r\[7\] _0712_ _0711_ _0710_ VDD VSS
+ VSS VDD sky130_fd_sc_hd__a22o_1
X_1291_ VSS VDD core.osr.next_result_w\[3\] core.cnb.result_out\[3\] _0649_ VSS VDD
+ sky130_fd_sc_hd__xnor2_2
XANTENNA__1778__RESET_B net69 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_23_118 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_23_107 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_51_416 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_51_449 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_1627_ core.osr.next_result_w\[5\] _0151_ core.osr.next_result_w\[11\] _0123_ _0124_
+ VSS VDD VSS VDD sky130_fd_sc_hd__o22a_1
X_1558_ VSS VDD _0008_ _0095_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XANTENNA__1533__A1 _0079_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1489_ _0433_ _0059_ core.cnb.data_register_r\[9\] _0063_ _0344_ core.cnb.data_register_r\[8\]
+ VDD VSS VSS VDD sky130_fd_sc_hd__a2111oi_1
XFILLER_100_123 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_86_379 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_36_59 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_36_48 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_14_129 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_52_14 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_52_69 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_77_44 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_26_81 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1800__RESET_B net63 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1460__B1 core.pdc.col_out_n\[16\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1549__S _0089_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_0860_ core.cnb.shift_register_r\[8\] _0286_ core.cnb.shift_register_r\[9\] VDD VSS
+ VSS VDD sky130_fd_sc_hd__xor2_1
X_0791_ _0213_ _0218_ _0215_ core.osr.sample_count_r\[4\] _0217_ VDD VSS VSS VDD sky130_fd_sc_hd__o2bb2a_1
XANTENNA__1212__A0 core.cnb.data_register_r\[5\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1412_ _0752_ core.osr.next_sample_count_w\[1\] core.osr.is_last_sample VSS VDD VSS
+ VDD sky130_fd_sc_hd__nor2_1
XANTENNA__1515__A1 _0353_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1343_ _0697_ _0695_ _0693_ VSS VDD VSS VDD sky130_fd_sc_hd__nand2_1
X_1274_ _0636_ _0635_ core.osr.result_r\[0\] VSS VDD VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_83_349 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_51_213 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_51_202 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_91_382 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_51_257 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1451__B1 _0513_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_0989_ VSS VDD _0415_ _0368_ _0355_ _0369_ VSS VDD sky130_fd_sc_hd__and3_1
XFILLER_86_132 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_47_14 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_63_57 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_128_94 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_3_876 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_26_9 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_0912_ _0278_ _0338_ _0279_ VSS VDD VSS VDD sky130_fd_sc_hd__nor2_1
X_0843_ core.cnb.shift_register_r\[4\] _0269_ core.cnb.shift_register_r\[1\] core.cnb.is_sampling_w
+ VDD VSS VSS VDD sky130_fd_sc_hd__or3_1
XANTENNA__1308__A core.cnb.result_out\[5\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1326_ core.osr.result_r\[7\] _0681_ _0680_ VSS VDD VSS VDD sky130_fd_sc_hd__or2_1
X_1257_ _0624_ _0615_ core.cnb.average_sum_r\[0\] VSS VDD VSS VDD sky130_fd_sc_hd__nand2_1
X_1188_ core.cnb.sampled_avg_control_r\[1\] core.cnb.sampled_avg_control_r\[0\] core.cnb.sampled_avg_control_r\[2\]
+ core.cnb.comparator_in _0571_ _0572_ VSS VDD VSS VDD sky130_fd_sc_hd__o41a_1
XPHY_208 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_219 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1777__CLK net56 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_0_879 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_47_327 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_114_41 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_114_85 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1773__D core.osr.next_result_w\[5\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1111_ VSS VDD core.pdc.col_out_n\[14\] _0522_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_0_53 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_1042_ _0465_ _0376_ _0464_ VSS VDD VSS VDD sky130_fd_sc_hd__nand2_2
XFILLER_0_97 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_119_104 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_134_129 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_0826_ VDD VSS _0252_ core.cnb.shift_register_r\[13\] VSS VDD sky130_fd_sc_hd__buf_2
XFILLER_0_109 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_88_205 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1038__A _0461_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_88_227 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_28_49 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_1309_ core.osr.result_r\[5\] _0665_ core.cnb.result_out\[5\] VDD VSS VSS VDD sky130_fd_sc_hd__or2_2
XFILLER_84_477 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1501__A _0352_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_52_385 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_60_36 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_69_12 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xadc_top_90 dummypin[5] adc_top_90/HI VDD VSS VSS VDD sky130_fd_sc_hd__conb_1
XFILLER_107_3 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_69_34 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_109_96 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_69_78 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_47_135 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_input27_A config_2_in[4] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1636__A0 _0709_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_90_469 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XPHY_550 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_86_8 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1557__S _0089_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1660_ core.osr.next_result_w\[15\] _0178_ core.osr.next_result_w\[17\] _0177_ _0230_
+ _0124_ VSS VDD VSS VDD sky130_fd_sc_hd__o221a_1
XFILLER_50_91 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_1591_ _0120_ _0119_ _0113_ core.osr.next_result_w\[6\] _0111_ _0118_ VSS VDD VSS
+ VDD sky130_fd_sc_hd__a32o_1
XFILLER_85_208 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1025_ _0450_ _0449_ VSS VDD VSS VDD sky130_fd_sc_hd__clkbuf_4
XFILLER_14_29 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_50_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_0809_ _0236_ _0209_ _0235_ VSS VDD VSS VDD sky130_fd_sc_hd__nor2_4
X_1789_ core.cnb.shift_register_r\[1\] net63 _0032_ net78 VSS VDD VSS VDD sky130_fd_sc_hd__dfrtp_2
XFILLER_29_102 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_29_113 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_44_127 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_111_20 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_41_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_71_57 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_20_61 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_48_411 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_96_65 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_48_477 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1141__A _0450_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_50_119 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_90_288 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_32_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XPHY_380 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_391 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_1712_ VSS VDD _0635_ _0214_ net12 _0208_ VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_6_41 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1643_ _0111_ _0164_ core.osr.next_result_w\[14\] VSS VDD VSS VDD sky130_fd_sc_hd__or2_1
XFILLER_6_85 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1574_ _0105_ _0232_ _0219_ VSS VDD VSS VDD sky130_fd_sc_hd__nand2_1
XANTENNA__0899__A1 core.cnb.data_register_r\[5\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_99_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_112_110 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_54_436 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_17 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_28 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1051__A _0466_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_41_119 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_39 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_1008_ _0433_ _0348_ _0349_ VSS VDD VSS VDD sky130_fd_sc_hd__nor2_4
XFILLER_23_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_41_49 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_89_366 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_106_53 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1303__A2 _0651_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_122_85 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_14_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_82_89 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_15_94 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_31_93 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1136__A _0374_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1290_ _0212_ _0649_ _0648_ VSS VDD VSS VDD sky130_fd_sc_hd__or2_1
XFILLER_48_296 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1626_ _0150_ _0149_ _0111_ VSS VDD VSS VDD sky130_fd_sc_hd__nand2_1
X_1557_ VSS VDD _0089_ core.cnb.next_data_register_w\[5\] core.cnb.result_out\[5\]
+ _0095_ VSS VDD sky130_fd_sc_hd__mux2_1
XANTENNA__1046__A _0466_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1533__A2 _0081_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1488_ _0062_ _0433_ _0061_ _0057_ VSS VDD VSS VDD sky130_fd_sc_hd__a21bo_1
XFILLER_54_222 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_54_277 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_52_37 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_52_48 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_50_472 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1221__A1 _0427_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_133_95 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_93_77 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1460__A1 _0353_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1776__D core.osr.next_result_w\[8\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_0790_ _0214_ _0217_ _0216_ VSS VDD VSS VDD sky130_fd_sc_hd__nor2_1
XANTENNA__1212__A1 _0420_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1411_ VSS VDD core.osr.sample_count_r\[1\] _0752_ core.osr.sample_count_r\[0\] VSS
+ VDD sky130_fd_sc_hd__xnor2_1
XANTENNA_nmat_en_bit_n[2] core.cnb.pswitch_out\[2\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1342_ _0693_ _0696_ _0695_ VSS VDD VSS VDD sky130_fd_sc_hd__or2_1
X_1273_ VDD VSS _0635_ _0634_ VSS VDD sky130_fd_sc_hd__buf_4
XFILLER_83_328 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_22_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_138_29 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_0988_ _0365_ _0414_ _0360_ VSS VDD VSS VDD sky130_fd_sc_hd__or2_1
X_1609_ _0132_ core.cnb.result_out\[0\] _0135_ _0136_ VDD VSS VSS VDD sky130_fd_sc_hd__a21o_1
XANTENNA_input1_A config_1_in[0] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_47_26 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_47_48 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_103_21 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_137_3 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_50_291 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_3_888 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_92_169 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_pmat_rowon_n[1] core.pdc.row_out_n\[2\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_0911_ _0259_ _0337_ _0264_ VSS VDD VSS VDD sky130_fd_sc_hd__nor2_1
X_0842_ _0268_ _0262_ VSS VDD VSS VDD sky130_fd_sc_hd__clkbuf_4
XFILLER_88_409 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_1325_ core.cnb.result_out\[6\] _0680_ core.osr.result_r\[6\] VSS VDD VSS VDD sky130_fd_sc_hd__or2_1
XANTENNA__1324__A _0651_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1256_ core.cnb.next_average_counter_w\[4\] _0622_ _0615_ _0623_ VSS VDD VSS VDD
+ sky130_fd_sc_hd__o21a_1
X_1187_ core.cnb.sampled_avg_control_r\[0\] core.cnb.sampled_avg_control_r\[2\] core.cnb.sampled_avg_control_r\[1\]
+ _0571_ core.cnb.average_sum_r\[4\] VDD VSS VSS VDD sky130_fd_sc_hd__or4b_1
XFILLER_83_169 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_91_180 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_209 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_33_17 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_137_105 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_134_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_58_47 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_58_36 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_87_420 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_114_53 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_114_64 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_114_97 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_130_85 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_90_67 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_128_127 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_125_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_24_7 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1144__A core.cnb.data_register_r\[0\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1110_ _0521_ _0449_ _0522_ _0519_ VSS VDD VSS VDD sky130_fd_sc_hd__o21ba_1
X_1041_ VSS VDD _0464_ _0463_ _0462_ _0454_ VSS VDD sky130_fd_sc_hd__and3_1
X_0825_ _0243_ _0251_ _0247_ _0237_ _0250_ VSS VDD VSS VDD sky130_fd_sc_hd__o22a_1
XFILLER_116_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_88_239 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1308_ VDD VSS _0664_ core.osr.result_r\[5\] core.cnb.result_out\[5\] VSS VDD sky130_fd_sc_hd__and2_1
X_1239_ VDD VSS _0612_ _0611_ net53 VSS VDD sky130_fd_sc_hd__and2_1
XFILLER_52_397 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_60_15 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_60_48 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_100_99 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xadc_top_91 dummypin[6] adc_top_91/HI VDD VSS VSS VDD sky130_fd_sc_hd__conb_1
XFILLER_107_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_47_169 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_551 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_540 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1139__A _0352_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1590_ _0110_ _0119_ core.osr.next_result_w\[2\] VSS VDD VSS VDD sky130_fd_sc_hd__or2_1
X_1024_ _0449_ _0427_ VSS VDD VSS VDD sky130_fd_sc_hd__clkbuf_4
XANTENNA__1602__A core.osr.next_result_w\[8\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_50_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_30_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_0808_ _0212_ _0234_ _0221_ _0235_ VSS VDD VSS VDD sky130_fd_sc_hd__nor3_4
X_1788_ core.cnb.is_sampling_w _0031_ VDD net64 net78 VSS VSS VDD sky130_fd_sc_hd__dfstp_4
XANTENNA__1563__A0 core.cnb.result_out\[8\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_55_15 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_84_253 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_44_117 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_55_48 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_111_32 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_71_47 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_41_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_71_69 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_121_122 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0964__C _0366_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1141__B _0423_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_32_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XPHY_370 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_381 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_392 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_1711_ VSS VDD _0049_ _0207_ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_1642_ _0232_ _0163_ _0162_ VSS VDD VSS VDD sky130_fd_sc_hd__or2_1
XFILLER_6_53 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_6_97 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1573_ VDD VSS _0104_ _0103_ VSS VDD sky130_fd_sc_hd__buf_2
XFILLER_99_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XPHY_18 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_54_448 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1007_ _0425_ _0426_ _0432_ _0406_ _0431_ _0427_ VSS VDD VSS VDD sky130_fd_sc_hd__a311o_1
XANTENNA__1051__B _0472_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_23_879 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_9_8 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1507__A _0352_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_66_69 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_17_117 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_82_13 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_122_75 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_82_57 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_14_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_15_51 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_99_109 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xoutput50 VDD VSS result_out[8] net50 VSS VDD sky130_fd_sc_hd__buf_2
XANTENNA__1152__A core.cnb.nswitch_out\[2\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_48_264 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_51_407 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1716__RESET_B net67 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1518__B1 net52 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1625_ VSS VDD _0110_ _0709_ _0691_ _0149_ VSS VDD sky130_fd_sc_hd__mux2_1
X_1556_ VSS VDD _0007_ _0094_ VSS VDD sky130_fd_sc_hd__clkbuf_1
XANTENNA__1046__B _0468_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1487_ _0328_ _0342_ _0061_ _0060_ _0058_ VDD VSS VSS VDD sky130_fd_sc_hd__a22o_1
XFILLER_86_315 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1062__A _0345_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1237__A _0588_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_89_142 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_77_57 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_77_68 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_9_113 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA_pmat_col_n[9] core.pdc.col_out_n\[9\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_61_8 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1410_ core.osr.next_sample_count_w\[0\] _0236_ core.osr.sample_count_r\[0\] VSS
+ VDD VSS VDD sky130_fd_sc_hd__nand2_1
XANTENNA__1515__A3 _0079_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_nmat_en_bit_n[1] core.cnb.pswitch_out\[1\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1341_ _0694_ _0695_ _0682_ VSS VDD VSS VDD sky130_fd_sc_hd__nor2_1
X_1272_ _0634_ _0209_ core.osr.sample_count_r\[0\] _0211_ _0210_ VDD VSS VSS VDD sky130_fd_sc_hd__a31oi_4
XFILLER_83_318 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_0987_ _0356_ _0412_ _0359_ _0411_ _0413_ VSS VDD VSS VDD sky130_fd_sc_hd__a31o_1
XANTENNA__1057__A _0364_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1608_ _0134_ net46 _0135_ _0104_ VSS VDD VSS VDD sky130_fd_sc_hd__and3b_1
X_1539_ VSS VDD _0588_ net1 core.cnb.sampled_avg_control_r\[0\] _0085_ VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_47_38 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1520__A _0352_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_10_123 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_12_41 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_12_85 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_88_45 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_88_89 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1130__A1 _0529_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_0910_ _0306_ _0336_ _0335_ _0325_ VDD VSS VSS VDD sky130_fd_sc_hd__or3_1
XFILLER_53_70 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_0841_ _0266_ _0267_ core.cnb.data_register_r\[2\] VSS VDD VSS VDD sky130_fd_sc_hd__nor2_1
XANTENNA__1576__S _0235_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_45_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_1324_ VSS VDD _0679_ _0653_ _0651_ _0678_ VSS VDD sky130_fd_sc_hd__and3_1
XFILLER_83_104 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1255_ VSS VDD _0623_ core.cnb.average_counter_r\[3\] _0621_ _0561_ VSS VDD sky130_fd_sc_hd__and3_1
X_1186_ core.cnb.sampled_avg_control_r\[2\] core.cnb.sampled_avg_control_r\[0\] core.cnb.sampled_avg_control_r\[1\]
+ _0570_ core.cnb.average_sum_r\[1\] VDD VSS VSS VDD sky130_fd_sc_hd__or4b_1
XANTENNA__1121__A1 _0354_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_91_192 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_134_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_87_432 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1360__A1 core.cnb.result_out\[7\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_114_76 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1112__A1 _0449_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_82_192 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_130_97 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_90_35 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_23_73 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_99_22 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_125_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_48_70 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1040_ _0463_ _0453_ VSS VDD VSS VDD sky130_fd_sc_hd__clkbuf_4
X_0824_ VSS VDD core.cnb.shift_register_r\[4\] _0249_ _0248_ _0250_ VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_134_109 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_116_879 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_28_18 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_84_435 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1307_ core.osr.next_result_w\[5\] _0663_ core.cnb.result_out\[5\] VSS VDD VSS VDD
+ sky130_fd_sc_hd__xnor2_4
X_1238_ VSS VDD _0586_ _0556_ core.cnb.data_register_r\[11\] _0611_ VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_44_39 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1169_ _0547_ _0555_ _0550_ _0556_ VSS VDD VSS VDD sky130_fd_sc_hd__nor3b_4
XFILLER_125_109 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_109_32 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xadc_top_92 dummypin[7] adc_top_92/HI VDD VSS VSS VDD sky130_fd_sc_hd__conb_1
XFILLER_109_65 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_107_879 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_109_87 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_47_104 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_85_24 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1333__A1 core.cnb.result_out\[6\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_85_57 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_87_295 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_552 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_541 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_530 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_1023_ VDD VSS _0448_ _0447_ VSS VDD sky130_fd_sc_hd__buf_6
XANTENNA__1627__A2 core.osr.next_result_w\[5\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1787_ core.osr.result_r\[19\] net72 core.osr.next_result_w\[19\] net58 VSS VDD VSS
+ VDD sky130_fd_sc_hd__dfrtp_1
X_0807_ _0225_ _0228_ _0210_ _0231_ _0233_ _0234_ VSS VDD VSS VDD sky130_fd_sc_hd__o2111ai_4
XFILLER_39_28 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1065__A _0373_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_84_265 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_84_276 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_84_287 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_111_44 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_71_26 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_136_41 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_136_85 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_20_96 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_48_402 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_29_61 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_input32_A config_2_in[9] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_90_279 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1490__B1 _0433_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XPHY_360 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_61_70 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XPHY_371 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_382 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_393 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_1710_ VSS VDD _0736_ net11 _0213_ _0207_ VSS VDD sky130_fd_sc_hd__mux2_1
X_1641_ VSS VDD _0110_ core.osr.next_result_w\[12\] core.osr.next_result_w\[10\] _0162_
+ VSS VDD sky130_fd_sc_hd__mux2_1
XFILLER_6_65 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1572_ net12 _0103_ net11 net10 VDD VSS VSS VDD sky130_fd_sc_hd__or3_1
XFILLER_54_405 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_1006_ _0431_ _0350_ _0429_ _0346_ _0430_ VSS VDD VSS VDD sky130_fd_sc_hd__and4_1
XANTENNA__1233__B1 _0588_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_89_346 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_89_357 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_66_15 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1523__A _0074_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_122_21 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_122_43 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xoutput40 VDD VSS result_out[13] net40 VSS VDD sky130_fd_sc_hd__buf_2
Xoutput51 VDD VSS result_out[9] net51 VSS VDD sky130_fd_sc_hd__buf_2
XFILLER_88_390 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_190 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_1624_ _0145_ _0148_ _0115_ _0146_ _0021_ VSS VDD VSS VDD sky130_fd_sc_hd__a31o_1
X_1555_ VSS VDD _0089_ core.cnb.next_data_register_w\[4\] core.cnb.result_out\[4\]
+ _0094_ VSS VDD sky130_fd_sc_hd__mux2_1
X_1486_ core.cnb.data_register_r\[8\] _0060_ _0059_ _0541_ VDD VSS VSS VDD sky130_fd_sc_hd__or3_1
XFILLER_86_327 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_54_235 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_54_246 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_22_121 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_117_32 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_77_36 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_117_87 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_85_371 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_85_393 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_93_46 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_93_57 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_26_40 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_26_95 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_pmat_col_n[8] core.pdc.col_out_n\[8\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_42_72 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1340_ VSS VDD _0686_ core.cnb.result_out\[7\] _0694_ _0688_ _0684_ VSS VDD sky130_fd_sc_hd__and4b_1
XANTENNA_nmat_en_bit_n[0] core.cnb.pswitch_out\[0\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_95_113 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_1271_ core.cnb.next_average_sum_w\[4\] _0632_ _0615_ _0633_ VSS VDD VSS VDD sky130_fd_sc_hd__o21a_1
XFILLER_95_124 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_83_308 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_91_363 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_0986_ _0412_ _0411_ _0365_ _0314_ _0266_ _0359_ VSS VDD VSS VDD sky130_fd_sc_hd__a32o_1
XANTENNA__1338__A core.cnb.result_out\[8\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xadc_top_100 dummypin[15] adc_top_100/HI VDD VSS VSS VDD sky130_fd_sc_hd__conb_1
X_1607_ VDD VSS _0134_ _0133_ VSS VDD sky130_fd_sc_hd__buf_2
XFILLER_86_102 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
X_1538_ core.pdc.row_out_n\[15\] _0074_ core.ndc.row_out_n\[4\] VSS VDD VSS VDD sky130_fd_sc_hd__nand2_1
XANTENNA__1073__A _0345_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1469_ _0506_ _0450_ _0052_ core.ndc.col_out_n\[24\] VDD VSS VSS VDD sky130_fd_sc_hd__a21o_1
XFILLER_12_53 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_12_97 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_88_13 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1682__S _0568_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_5_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_88_68 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_88_57 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_92_149 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_37_72 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_37_61 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_0840_ _0266_ _0251_ _0265_ VSS VDD VSS VDD sky130_fd_sc_hd__nand2_2
X_1323_ _0665_ core.osr.result_r\[7\] core.cnb.result_out\[6\] _0678_ _0669_ VDD VSS
+ VSS VDD sky130_fd_sc_hd__a211oi_1
X_1254_ core.cnb.average_counter_r\[3\] _0621_ _0622_ _0561_ VDD VSS VSS VDD sky130_fd_sc_hd__a21oi_1
XFILLER_49_393 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1185_ _0569_ core.cnb.sampled_avg_control_r\[2\] core.cnb.sampled_avg_control_r\[0\]
+ VSS VDD VSS VDD sky130_fd_sc_hd__nand2_1
XANTENNA__0880__B2 core.cnb.data_register_r\[7\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_80_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_0969_ _0300_ _0395_ _0338_ VSS VDD VSS VDD sky130_fd_sc_hd__nor2_1
XFILLER_87_400 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_87_444 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1531__A _0074_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_55_374 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_82_160 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_71_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_90_25 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_139_41 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_23_96 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_139_85 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_99_78 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_17_8 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1103__A2 _0420_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1639__B1 _0236_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_62_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_0823_ core.cnb.shift_register_r\[5\] _0249_ core.cnb.shift_register_r\[7\] VSS VDD
+ VSS VDD sky130_fd_sc_hd__or2_1
XFILLER_80_80 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1306_ _0663_ _0662_ _0634_ VSS VDD VSS VDD sky130_fd_sc_hd__nand2_1
XFILLER_84_425 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1237_ _0610_ core.cnb.next_data_register_w\[10\] _0588_ VSS VDD VSS VDD sky130_fd_sc_hd__nor2_1
X_1168_ VSS VDD _0555_ _0546_ _0544_ _0551_ _0554_ VSS VDD sky130_fd_sc_hd__a211o_1
XFILLER_44_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_53_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1645__A3 core.osr.next_result_w\[8\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1099_ VSS VDD _0512_ _0424_ _0513_ core.pdc.col_out_n\[11\] VSS VDD sky130_fd_sc_hd__o21ai_1
XANTENNA__1790__CLK net77 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xadc_top_93 dummypin[8] adc_top_93/HI VDD VSS VSS VDD sky130_fd_sc_hd__conb_1
XFILLER_109_44 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_109_77 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_87_230 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1261__A _0616_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_18_85 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_90_406 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_44_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XPHY_553 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_542 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_531 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_520 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_34_73 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1436__A _0423_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1171__A net52 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1022_ VDD VSS _0447_ _0446_ _0432_ VSS VDD sky130_fd_sc_hd__and2_1
XFILLER_35_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
X_1786_ core.osr.result_r\[18\] net71 core.osr.next_result_w\[18\] net58 VSS VDD VSS
+ VDD sky130_fd_sc_hd__dfrtp_1
X_0806_ VSS VDD _0233_ core.osr.sample_count_r\[4\] core.osr.sample_count_r\[6\] _0216_
+ _0232_ VSS VDD sky130_fd_sc_hd__a211o_1
XFILLER_26_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_52_141 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_136_53 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_96_35 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_136_97 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XANTENNA__1690__S _0616_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_96_57 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_29_40 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_input25_A config_2_in[2] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_48_469 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_17_867 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_45_94 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1803__RESET_B net63 VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XPHY_350 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_361 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_84_8 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_372 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_383 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_394 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
X_1640_ _0159_ _0161_ _0134_ _0160_ _0024_ VSS VDD VSS VDD sky130_fd_sc_hd__a31o_1
X_1571_ core.cnb.result_out\[11\] _0101_ _0014_ _0611_ _0102_ VDD VSS VSS VDD sky130_fd_sc_hd__a22o_1
XFILLER_6_77 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
X_1005_ VDD VSS _0430_ _0365_ _0364_ VSS VDD sky130_fd_sc_hd__and2_1
XFILLER_41_19 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
X_1769_ core.osr.result_r\[1\] net66 core.osr.next_result_w\[1\] net55 VSS VDD VSS
+ VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_89_325 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_106_12 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_106_23 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_106_78 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1523__B core.ndc.row_out_n\[12\] VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_82_48 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1472__A1 _0424_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_53_472 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_15_86 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_31_30 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xoutput41 VDD VSS result_out[14] net41 VSS VDD sky130_fd_sc_hd__buf_2
XPHY_180 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_191 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1215__A1 _0410_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA__1518__A2 _0079_ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
X_1623_ VSS VDD _0104_ _0640_ _0147_ _0148_ VSS VDD sky130_fd_sc_hd__o21ai_1
X_1554_ VSS VDD _0006_ _0093_ VSS VDD sky130_fd_sc_hd__clkbuf_1
X_1485_ core.cnb.data_register_r\[10\] _0059_ VDD VSS VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_100_105 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_100_116 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
.ends

