* NGSPICE file created from adc_clkgen_with_edgedetect.ext - technology: sky130A

.subckt sky130_fd_sc_hd__inv_2 A Y VPWR VGND VNB VPB
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=5.2e+11p ps=5.04e+06u w=1e+06u l=150000u
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=3.38e+11p pd=3.64e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
C0 VPWR Y 0.19fF
C1 Y VGND 0.14fF
C2 VGND VNB 0.27fF
C3 VPWR VNB 0.27fF
C4 A VNB 0.28fF
C5 VPB VNB 0.34fF
.ends

.subckt sky130_fd_sc_hd__decap_3 VPWR VGND VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=4.524e+11p pd=4.52e+06u as=0p ps=0u w=870000u l=590000u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=2.86e+11p pd=3.24e+06u as=0p ps=0u w=550000u l=590000u
C0 VGND VPWR 0.33fF
C1 VPWR VNB 0.47fF
C2 VGND VNB 0.44fF
C3 VPB VNB 0.34fF
.ends

.subckt sky130_fd_sc_hd__decap_4 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=4.524e+11p pd=4.52e+06u as=0p ps=0u w=870000u l=1.05e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=2.86e+11p pd=3.24e+06u as=0p ps=0u w=550000u l=1.05e+06u
C0 VGND VPWR 0.52fF
C1 VPWR VNB 0.61fF
C2 VGND VNB 0.56fF
C3 VPB VNB 0.43fF
.ends

.subckt sky130_fd_sc_hd__mux2_1 VGND VPWR S A1 A0 X VNB VPB a_505_21#
X0 VPWR a_505_21# a_535_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=4.553e+11p pd=4.29e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X1 a_505_21# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X2 a_218_374# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X3 VGND a_505_21# a_439_47# VNB sky130_fd_pr__nfet_01v8 ad=5.155e+11p pd=4.31e+06u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4 a_76_199# A0 a_218_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X5 a_505_21# S VGND VNB sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X6 a_439_47# A0 a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X7 a_535_374# A1 a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_76_199# A1 a_218_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X9 a_218_47# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
C0 A1 a_76_199# 0.17fF
C1 VGND a_76_199# 0.11fF
C2 A0 A1 0.24fF
C3 a_76_199# S 0.28fF
C4 X VPWR 0.11fF
C5 a_505_21# S 0.14fF
C6 VPWR S 0.29fF
C7 VGND VNB 0.50fF
C8 A1 VNB 0.11fF
C9 A0 VNB 0.12fF
C10 S VNB 0.29fF
C11 VPWR VNB 0.45fF
C12 VPB VNB 0.87fF
C13 a_505_21# VNB 0.21fF
C14 a_76_199# VNB 0.15fF
.ends

.subckt sky130_fd_sc_hd__decap_6 VPWR VGND VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=4.524e+11p pd=4.52e+06u as=0p ps=0u w=870000u l=1.97e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=2.86e+11p pd=3.24e+06u as=0p ps=0u w=550000u l=1.97e+06u
C0 VPWR VGND 0.89fF
C1 VPWR VPB 0.10fF
C2 VPWR VNB 0.85fF
C3 VGND VNB 0.77fF
C4 VPB VNB 0.60fF
.ends

.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VPWR VPB VNB
D0 VNB DIODE sky130_fd_pr__diode_pw2nd_05v5 pj=2.64e+06 area=4.347e+11
C0 VGND VNB 0.15fF
C1 VPWR VNB 0.14fF
C2 DIODE VNB 0.19fF
C3 VPB VNB 0.25fF
.ends

.subckt sky130_fd_sc_hd__or2_1 A X B VGND VPWR VNB VPB
X0 VGND A a_68_297# VNB sky130_fd_pr__nfet_01v8 ad=3.097e+11p pd=3.33e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X1 a_68_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 X a_68_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X3 VPWR A a_150_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=2.915e+11p pd=2.67e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X4 X a_68_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=3.4e+11p pd=2.68e+06u as=0p ps=0u w=1e+06u l=150000u
X5 a_150_297# B a_68_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
C0 A a_68_297# 0.15fF
C1 VGND VNB 0.32fF
C2 X VNB 0.11fF
C3 B VNB 0.19fF
C4 VPWR VNB 0.29fF
C5 VPB VNB 0.52fF
C6 a_68_297# VNB 0.18fF
.ends

.subckt sky130_mm_sc_hd_dlyPoly5ns VPWR VGND in out VNB VPB mid a_1632_71# a_1691_329#
X0 a_1691_329# out VGND VPB sky130_fd_pr__pfet_01v8_hvt ad=7.52e+11p pd=6.68e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1 a_1691_329# mid VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.72e+11p ps=4.38e+06u w=800000u l=150000u
X2 out mid a_1691_329# VPB sky130_fd_pr__pfet_01v8_hvt ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X3 VGND out a_1691_329# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4 VGND mid VGND VNB sky130_fd_pr__nfet_01v8 ad=1.0453e+12p pd=9.52e+06u as=0p ps=0u w=1.375e+06u l=2.045e+06u
X5 a_1632_71# mid VGND VNB sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X6 VPWR out a_1632_71# VNB sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X7 a_1632_71# out VPWR VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 out mid a_1632_71# VNB sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X9 mid in VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=1.42e+06u
X10 mid in VGND VNB sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=3.69e+06u
C0 mid VGND 2.09fF
C1 VGND VPWR 0.40fF
C2 mid VPB 0.19fF
C3 VPB VPWR 0.28fF
C4 a_1691_329# VPWR 0.52fF
C5 in VGND 0.14fF
C6 out VPWR 0.17fF
C7 VPB in 0.15fF
C8 mid VPWR 0.70fF
C9 VPB VGND 0.12fF
C10 a_1691_329# VGND 0.31fF
C11 mid in 0.16fF
C12 a_1632_71# VGND 0.48fF
C13 VGND VNB 1.42fF
C14 VPWR VNB 1.15fF
C15 in VNB 1.04fF
C16 out VNB 0.34fF
C17 VPB VNB 1.93fF
C18 mid VNB 1.08fF
.ends

.subckt sky130_fd_sc_hd__and2_1 VPWR VGND X B A VNB VPB
X0 VPWR B a_59_75# VPB sky130_fd_pr__pfet_01v8_hvt ad=4.507e+11p pd=4.18e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X1 X a_59_75# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=4.75e+11p pd=2.95e+06u as=0p ps=0u w=1e+06u l=150000u
X2 VGND B a_145_75# VNB sky130_fd_pr__nfet_01v8 ad=2.236e+11p pd=2.08e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X3 a_59_75# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 X a_59_75# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X5 a_145_75# A a_59_75# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
C0 a_59_75# VPWR 0.13fF
C1 B a_59_75# 0.13fF
C2 VGND VNB 0.31fF
C3 X VNB 0.11fF
C4 B VNB 0.12fF
C5 A VNB 0.19fF
C6 VPWR VNB 0.30fF
C7 VPB VNB 0.52fF
C8 a_59_75# VNB 0.20fF
.ends

.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=4.524e+11p pd=4.52e+06u as=0p ps=0u w=870000u l=4.73e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=2.86e+11p pd=3.24e+06u as=0p ps=0u w=550000u l=4.73e+06u
C0 VPWR VPB 0.21fF
C1 VPB VGND 0.20fF
C2 VPWR VGND 1.27fF
C3 VPWR VNB 1.62fF
C4 VGND VNB 1.45fF
C5 VPB VNB 1.14fF
.ends

.subckt sky130_fd_sc_hd__nor2b_1 B_N Y A VGND VPWR VNB VPB
X0 Y a_74_47# a_265_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X1 VPWR B_N a_74_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=3.146e+11p pd=2.78e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X2 a_265_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=3.695e+11p ps=3.79e+06u w=650000u l=150000u
X4 VGND B_N a_74_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X5 VGND a_74_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
C0 VGND Y 0.17fF
C1 A a_74_47# 0.14fF
C2 VGND VNB 0.33fF
C3 B_N VNB 0.23fF
C4 VPWR VNB 0.30fF
C5 VPB VNB 0.52fF
C6 a_74_47# VNB 0.18fF
.ends

.subckt sky130_fd_sc_hd__decap_8 VPWR VGND VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=4.524e+11p pd=4.52e+06u as=0p ps=0u w=870000u l=2.89e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=2.86e+11p pd=3.24e+06u as=0p ps=0u w=550000u l=2.89e+06u
C0 VPB VPWR 0.13fF
C1 VPB VGND 0.12fF
C2 VPWR VGND 1.26fF
C3 VPWR VNB 1.11fF
C4 VGND VNB 1.00fF
C5 VPB VNB 0.78fF
.ends

.subckt sky130_fd_sc_hd__and2b_1 X A_N B VGND VPWR VNB VPB
X0 VPWR B a_207_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=5.986e+11p pd=5e+06u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X1 X a_207_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X2 a_297_47# a_27_413# a_207_413# VNB sky130_fd_pr__nfet_01v8 ad=1.008e+11p pd=1.32e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X3 X a_207_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=3.118e+11p ps=3.34e+06u w=650000u l=150000u
X4 a_207_413# a_27_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VPWR A_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X6 VGND B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_27_413# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
C0 a_207_413# B 0.14fF
C1 A_N a_27_413# 0.13fF
C2 a_207_413# a_27_413# 0.14fF
C3 VGND VNB 0.37fF
C4 VPWR VNB 0.32fF
C5 B VNB 0.13fF
C6 A_N VNB 0.21fF
C7 VPB VNB 0.60fF
C8 a_207_413# VNB 0.15fF
C9 a_27_413# VNB 0.17fF
.ends

.subckt sky130_fd_sc_hd__buf_1 VGND VPWR X A VNB VPB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=2.291e+11p pd=2.16e+06u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X1 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=1.508e+11p ps=1.62e+06u w=520000u l=150000u
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X3 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
C0 a_27_47# VPWR 0.11fF
C1 a_27_47# A 0.13fF
C2 VGND VNB 0.21fF
C3 VPWR VNB 0.19fF
C4 A VNB 0.17fF
C5 VPB VNB 0.34fF
C6 a_27_47# VNB 0.22fF
.ends

.subckt sky130_fd_sc_hd__dlymetal6s6s_1 VPWR VGND A X VNB VPB a_523_47#
X0 X a_629_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=5.82e+11p ps=5.85e+06u w=650000u l=150000u
X1 a_523_47# a_346_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X2 VGND a_240_47# a_346_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X3 a_240_47# a_63_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X4 VPWR a_240_47# a_346_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=8.445e+11p pd=7.95e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X5 VGND A a_63_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X6 VPWR A a_63_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X7 VPWR a_523_47# a_629_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X8 VGND a_523_47# a_629_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X9 a_523_47# a_346_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X10 a_240_47# a_63_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X11 X a_629_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
C0 VPWR a_629_47# 0.11fF
C1 a_63_47# VPWR 0.11fF
C2 a_346_47# a_240_47# 0.25fF
C3 a_346_47# a_523_47# 0.14fF
C4 VGND VPWR 0.11fF
C5 VGND a_629_47# 0.10fF
C6 VGND a_63_47# 0.11fF
C7 X a_629_47# 0.11fF
C8 A a_63_47# 0.20fF
C9 a_523_47# a_629_47# 0.25fF
C10 a_63_47# a_240_47# 0.14fF
C11 VGND VNB 0.54fF
C12 X VNB 0.10fF
C13 VPWR VNB 0.48fF
C14 A VNB 0.23fF
C15 VPB VNB 0.96fF
C16 a_629_47# VNB 0.14fF
C17 a_523_47# VNB 0.18fF
C18 a_240_47# VNB 0.18fF
C19 a_63_47# VNB 0.16fF
.ends

.subckt sky130_fd_sc_hd__buf_4 VPWR VGND X A VNB VPB a_27_47#
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=8e+11p pd=7.6e+06u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=5.2e+11p ps=5.5e+06u w=650000u l=150000u
X5 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X9 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
C0 a_27_47# VPWR 0.14fF
C1 X VGND 0.18fF
C2 X VPWR 0.26fF
C3 a_27_47# A 0.14fF
C4 a_27_47# VGND 0.11fF
C5 a_27_47# X 0.11fF
C6 VGND VNB 0.38fF
C7 VPWR VNB 0.35fF
C8 A VNB 0.14fF
C9 VPB VNB 0.60fF
C10 a_27_47# VNB 0.45fF
.ends

.subckt adc_clkgen_with_edgedetect VDD VSS clk_comp_out clk_dig_out dlycontrol1_in[0]
+ dlycontrol1_in[1] dlycontrol1_in[2] dlycontrol1_in[3] dlycontrol1_in[4] dlycontrol2_in[0]
+ dlycontrol2_in[1] dlycontrol2_in[2] dlycontrol2_in[3] dlycontrol2_in[4] dlycontrol3_in[0]
+ dlycontrol3_in[1] dlycontrol3_in[2] dlycontrol3_in[3] dlycontrol3_in[4] dlycontrol4_in[0]
+ dlycontrol4_in[1] dlycontrol4_in[2] dlycontrol4_in[3] dlycontrol4_in[4] dlycontrol4_in[5]
+ ena_in enable_dlycontrol_in ndecision_finish_in nsample_n_in nsample_n_out nsample_p_in
+ nsample_p_out sample_n_in sample_n_out sample_p_in sample_p_out start_conv_in
Xclkgen.delay_155ns_2.genblk1\[0\].control_invert dlycontrol2_in[0] clkgen.delay_155ns_2.bypass_enable_w\[0\]
+ VDD VSS VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_18_214 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_10_125 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_2.genblk1\[0\].dly_binary.out_mux VSS VDD clkgen.delay_155ns_2.genblk1\[0\].dly_binary.bypass_in
+ clkgen.clk_dig_out clkgen.delay_155ns_2.genblk1\[0\].dly_binary.signal_w\[1\] clkgen.delay_155ns_2.genblk1\[0\].dly_binary.out
+ VSS VDD clkgen.delay_155ns_2.genblk1\[0\].dly_binary.out_mux/a_505_21# sky130_fd_sc_hd__mux2_1
XFILLER_17_291 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_2.genblk1\[2\].dly_binary.out_mux VSS VDD clkgen.delay_155ns_2.genblk1\[2\].dly_binary.bypass_in
+ clkgen.delay_155ns_2.genblk1\[1\].dly_binary.out clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[4\]
+ clkgen.delay_155ns_2.genblk1\[2\].dly_binary.out VSS VDD clkgen.delay_155ns_2.genblk1\[2\].dly_binary.out_mux/a_505_21#
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_272 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.out_mux VSS VDD clkgen.delay_155ns_2.genblk1\[4\].dly_binary.bypass_in
+ clkgen.delay_155ns_2.genblk1\[3\].dly_binary.out clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[16\]
+ clkgen.clk_dig_delayed_w VSS VDD clkgen.delay_155ns_2.genblk1\[4\].dly_binary.out_mux/a_505_21#
+ sky130_fd_sc_hd__mux2_1
XANTENNA_clkgen.delay_155ns_1.genblk1\[2\].control_invert_A dlycontrol1_in[2] VSS
+ VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_2_143 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xedgedetect.or1 edgedetect.start_conv_edge_w clkgen.enable_loop_in edgedetect.ena_in
+ VSS VDD VSS VDD sky130_fd_sc_hd__or2_1
XFILLER_11_275 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_11_242 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_16_334 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xclkgen.delay_155ns_3.genblk1\[0\].dly_binary.genblk1\[0\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[0\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_3.genblk1\[0\].dly_binary.signal_w\[1\] VSS VDD clkgen.delay_155ns_3.genblk1\[0\].dly_binary.genblk1\[0\].delay_unit/mid
+ clkgen.delay_155ns_3.genblk1\[0\].dly_binary.genblk1\[0\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_3.genblk1\[0\].dly_binary.genblk1\[0\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XFILLER_4_205 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[1\].bypass_enable VDD VSS edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.bypass_in
+ edgedetect.dly_315ns_1.bypass_enable_w\[1\] edgedetect.dly_315ns_1.enable_dlycontrol_w
+ VSS VDD sky130_fd_sc_hd__and2_1
XFILLER_13_3 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_6_56 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_1_208 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_0_241 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA_clkgen.delay_155ns_2.genblk1\[1\].control_invert_A dlycontrol2_in[1] VSS
+ VDD VDD VSS sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[14\]
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[15\] VSS VDD clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit/mid
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XFILLER_13_156 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.delay_155ns_2.genblk1\[1\].dly_binary.and_bypass_switch_A_N clkgen.delay_155ns_2.genblk1\[1\].dly_binary.bypass_in
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_5_311 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xclkgen.delay_155ns_1.genblk1\[2\].bypass_enable VDD VSS clkgen.delay_155ns_1.genblk1\[2\].dly_binary.bypass_in
+ clkgen.delay_155ns_1.bypass_enable_w\[2\] clkgen.delay_155ns_1.enable_dlycontrol_w
+ VSS VDD sky130_fd_sc_hd__and2_1
Xclkgen.delay_155ns_2.genblk1\[3\].bypass_enable VDD VSS clkgen.delay_155ns_2.genblk1\[3\].dly_binary.bypass_in
+ clkgen.delay_155ns_2.bypass_enable_w\[3\] clkgen.delay_155ns_2.enable_dlycontrol_w
+ VSS VDD sky130_fd_sc_hd__and2_1
Xclkgen.delay_155ns_3.genblk1\[4\].bypass_enable VDD VSS clkgen.delay_155ns_3.genblk1\[4\].dly_binary.bypass_in
+ clkgen.delay_155ns_3.bypass_enable_w\[4\] clkgen.delay_155ns_3.enable_dlycontrol_w
+ VSS VDD sky130_fd_sc_hd__and2_1
XANTENNA_clkgen.delay_155ns_3.genblk1\[0\].control_invert_A dlycontrol3_in[0] VSS
+ VDD VDD VSS sky130_fd_sc_hd__diode_2
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[3\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[3\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[4\] VSS VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[3\].delay_unit/mid
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[3\].delay_unit/a_1632_71#
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[3\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XFILLER_0_58 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_sampledly04_A nsample_n_in VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_18_32 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_11_287 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_19_321 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[1\]
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[2\] VSS VDD clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit/mid
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[1\].control_invert dlycontrol4_in[1] edgedetect.dly_315ns_1.bypass_enable_w\[1\]
+ VDD VSS VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_13_305 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_10_319 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[8\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[8\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[9\] VSS VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[8\].delay_unit/mid
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[8\].delay_unit/a_1632_71#
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[8\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XFILLER_5_323 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_2_304 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[12\]
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[13\] VSS VDD clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit/mid
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[6\]
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[7\] VSS VDD clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit/mid
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XFILLER_5_153 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_3_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xedgedetect.nor1 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.in edgedetect.start_conv_edge_w
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.out VSS VDD VSS VDD sky130_fd_sc_hd__nor2b_1
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[0\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[1\] VSS VDD clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[0\].delay_unit/mid
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[0\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[0\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XFILLER_11_299 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_19_333 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xclkgen.delay_155ns_3.genblk1\[1\].control_invert dlycontrol3_in[1] clkgen.delay_155ns_3.bypass_enable_w\[1\]
+ VDD VSS VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_0_276 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[3\]
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[4\] VSS VDD edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit/mid
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit/a_1632_71#
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XFILLER_13_125 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[5\]
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[6\] VSS VDD clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit/mid
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XFILLER_8_173 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_5_335 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_2_316 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xclkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[1\]
+ clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[2\] VSS VDD clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit/mid
+ clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[10\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[10\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[11\] VSS VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[10\].delay_unit/mid
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[10\].delay_unit/a_1632_71#
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[10\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XFILLER_7_216 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[10\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[10\]
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[11\] VSS VDD clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[10\].delay_unit/mid
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[10\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[10\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[8\]
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[9\] VSS VDD edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit/mid
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit/a_1632_71#
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XFILLER_3_241 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[11\]
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[12\] VSS VDD edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit/mid
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit/a_1632_71#
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XFILLER_15_57 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[6\]
+ clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[7\] VSS VDD clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit/mid
+ clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XFILLER_0_222 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_11_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[4\]
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[5\] VSS VDD clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit/mid
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.and_bypass_switch_A_N edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.bypass_in
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[0\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[1\] VSS VDD clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[0\].delay_unit/mid
+ clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[0\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[0\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XFILLER_18_207 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[15\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[15\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[16\] VSS VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[15\].delay_unit/mid
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[15\].delay_unit/a_1632_71#
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[15\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XFILLER_12_58 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[15\]
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[16\] VSS VDD clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit/mid
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XFILLER_2_328 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_17_284 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.nor1 clkgen.enable_loop_in clkgen.delay_155ns_3.genblk1\[0\].dly_binary.in
+ clkgen.clk_dig_delayed_w VSS VDD VSS VDD sky130_fd_sc_hd__nor2b_1
XFILLER_11_235 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_sampledly02_A sample_n_in VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[9\]
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[10\] VSS VDD clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit/mid
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[3\]
+ edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[4\] VSS VDD edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit/mid
+ edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit/a_1632_71#
+ edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XFILLER_10_290 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_6_272 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xclkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[5\]
+ clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[6\] VSS VDD clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit/mid
+ clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XFILLER_19_187 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_3_275 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[2\].dly_binary.genblk1\[1\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[2\].dly_binary.signal_w\[1\]
+ clkgen.delay_155ns_3.genblk1\[2\].dly_binary.signal_w\[2\] VSS VDD clkgen.delay_155ns_3.genblk1\[2\].dly_binary.genblk1\[1\].delay_unit/mid
+ clkgen.delay_155ns_3.genblk1\[2\].dly_binary.genblk1\[1\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_3.genblk1\[2\].dly_binary.genblk1\[1\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XFILLER_0_212 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[2\].control_invert dlycontrol1_in[2] clkgen.delay_155ns_1.bypass_enable_w\[2\]
+ VDD VSS VSS VDD sky130_fd_sc_hd__inv_2
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[22\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[22\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[23\] VSS VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[22\].delay_unit/mid
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[22\].delay_unit/a_1632_71#
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[22\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XFILLER_12_171 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_8_164 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_8_120 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA_edgedetect.dly_315ns_1.enablebuffer_A enable_dlycontrol_in VSS VDD VDD VSS
+ sky130_fd_sc_hd__diode_2
XFILLER_5_112 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_14_244 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_14_211 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_2_115 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[27\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[27\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[28\] VSS VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[27\].delay_unit/mid
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[27\].delay_unit/a_1632_71#
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[27\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[4\]
+ clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[5\] VSS VDD clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit/mid
+ clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XFILLER_1_3 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.delay_155ns_1.genblk1\[1\].control_invert_A dlycontrol1_in[1] VSS
+ VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_clkgen.delay_155ns_2.enablebuffer_A enable_dlycontrol_in VSS VDD VDD VSS
+ sky130_fd_sc_hd__diode_2
XANTENNA_inbuf_3_A ndecision_finish_in VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_1_94 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_16_306 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_2.genblk1\[2\].dly_binary.genblk1\[0\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[1\] VSS VDD clkgen.delay_155ns_2.genblk1\[2\].dly_binary.genblk1\[0\].delay_unit/mid
+ clkgen.delay_155ns_2.genblk1\[2\].dly_binary.genblk1\[0\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_2.genblk1\[2\].dly_binary.genblk1\[0\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XFILLER_19_90 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xclkgen.clkdig_inverter clkgen.delay_155ns_1.genblk1\[4\].dly_binary.out clkgen.clk_dig_out
+ VDD VSS VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_15_15 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_16_125 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.delay_155ns_2.genblk1\[0\].control_invert_A dlycontrol2_in[0] VSS
+ VDD VDD VSS sky130_fd_sc_hd__diode_2
XPHY_0 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_7_93 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_3_18 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_12_16 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_17_297 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[3\]
+ edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[4\] VSS VDD edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit/mid
+ edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit/a_1632_71#
+ edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XFILLER_5_146 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_4_94 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xclkgen.delay_155ns_3.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[1\].dly_binary.signal_w\[1\]
+ clkgen.delay_155ns_3.genblk1\[1\].dly_binary.signal_w\[2\] VSS VDD clkgen.delay_155ns_3.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit/mid
+ clkgen.delay_155ns_3.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_3.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XFILLER_19_315 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_3_222 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_15_181 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[0\].dly_binary.out_mux VSS VDD edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.bypass_in
+ edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.in edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.signal_w\[1\]
+ edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.out VSS VDD edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.out_mux/a_505_21#
+ sky130_fd_sc_hd__mux2_1
XPHY_1 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xedgedetect.dly_315ns_1.genblk1\[2\].dly_binary.out_mux VSS VDD edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.bypass_in
+ edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.out edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[4\]
+ edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.out VSS VDD edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.out_mux/a_505_21#
+ sky130_fd_sc_hd__mux2_1
Xedgedetect.dly_315ns_1.genblk1\[0\].dly_binary.and_bypass_switch edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.signal_w\[0\]
+ edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.bypass_in edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.in
+ VSS VDD VSS VDD sky130_fd_sc_hd__and2b_1
Xinbuf_1 VSS VDD edgedetect.ena_in ena_in VSS VDD sky130_fd_sc_hd__buf_1
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.out_mux VSS VDD edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.bypass_in
+ edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.out edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[16\]
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.out VSS VDD edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.out_mux/a_505_21#
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_136 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsampledly31 VDD VSS sample_p_3 sample_p_4 VSS VDD sampledly31/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1
Xclkgen.delay_155ns_2.genblk1\[1\].dly_binary.genblk1\[0\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[1\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_2.genblk1\[1\].dly_binary.signal_w\[1\] VSS VDD clkgen.delay_155ns_2.genblk1\[1\].dly_binary.genblk1\[0\].delay_unit/mid
+ clkgen.delay_155ns_2.genblk1\[1\].dly_binary.genblk1\[0\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_2.genblk1\[1\].dly_binary.genblk1\[0\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XFILLER_2_106 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_1_194 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[2\].bypass_enable VDD VSS edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.bypass_in
+ edgedetect.dly_315ns_1.bypass_enable_w\[2\] edgedetect.dly_315ns_1.enable_dlycontrol_w
+ VSS VDD sky130_fd_sc_hd__and2_1
Xclkgen.delay_155ns_2.genblk1\[3\].control_invert dlycontrol2_in[3] clkgen.delay_155ns_2.bypass_enable_w\[3\]
+ VDD VSS VSS VDD sky130_fd_sc_hd__inv_2
XANTENNA_clkgen.delay_155ns_3.genblk1\[4\].dly_binary.out_mux_A0 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[16\]
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_1_63 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[10\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[10\]
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[11\] VSS VDD clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[10\].delay_unit/mid
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[10\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[10\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_clkgen.delay_155ns_2.genblk1\[4\].dly_binary.and_bypass_switch_A_N clkgen.delay_155ns_2.genblk1\[4\].dly_binary.bypass_in
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_10_94 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_15_171 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_2 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xclkgen.delay_155ns_1.genblk1\[3\].bypass_enable VDD VSS clkgen.delay_155ns_1.genblk1\[3\].dly_binary.bypass_in
+ clkgen.delay_155ns_1.bypass_enable_w\[3\] clkgen.delay_155ns_1.enable_dlycontrol_w
+ VSS VDD sky130_fd_sc_hd__and2_1
Xclkgen.delay_155ns_2.genblk1\[4\].bypass_enable VDD VSS clkgen.delay_155ns_2.genblk1\[4\].dly_binary.bypass_in
+ clkgen.delay_155ns_2.bypass_enable_w\[4\] clkgen.delay_155ns_2.enable_dlycontrol_w
+ VSS VDD sky130_fd_sc_hd__and2_1
Xinbuf_2 VSS VDD edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.in start_conv_in VSS
+ VDD sky130_fd_sc_hd__buf_1
XFILLER_5_307 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[15\]
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[16\] VSS VDD clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit/mid
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
Xsampledly21 VDD VSS sample_p_2 sample_p_3 VSS VDD sampledly21/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1
Xsampledly32 VDD VSS sample_n_3 sample_n_4 VSS VDD sampledly32/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1
XFILLER_4_63 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[0\].dly_binary.out_mux VSS VDD clkgen.delay_155ns_1.genblk1\[0\].dly_binary.bypass_in
+ clkgen.delay_155ns_1.genblk1\[0\].dly_binary.in clkgen.delay_155ns_1.genblk1\[0\].dly_binary.signal_w\[1\]
+ clkgen.delay_155ns_1.genblk1\[0\].dly_binary.out VSS VDD clkgen.delay_155ns_1.genblk1\[0\].dly_binary.out_mux/a_505_21#
+ sky130_fd_sc_hd__mux2_1
XFILLER_13_94 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_9_19 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_11_228 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[2\].dly_binary.out_mux VSS VDD clkgen.delay_155ns_1.genblk1\[2\].dly_binary.bypass_in
+ clkgen.delay_155ns_1.genblk1\[1\].dly_binary.out clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[4\]
+ clkgen.delay_155ns_1.genblk1\[2\].dly_binary.out VSS VDD clkgen.delay_155ns_1.genblk1\[2\].dly_binary.out_mux/a_505_21#
+ sky130_fd_sc_hd__mux2_1
XFILLER_19_306 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_6_210 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.out_mux VSS VDD clkgen.delay_155ns_1.genblk1\[4\].dly_binary.bypass_in
+ clkgen.delay_155ns_1.genblk1\[3\].dly_binary.out clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[16\]
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.out VSS VDD clkgen.delay_155ns_1.genblk1\[4\].dly_binary.out_mux/a_505_21#
+ sky130_fd_sc_hd__mux2_1
Xedgedetect.dly_315ns_1.genblk1\[1\].dly_binary.and_bypass_switch edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.signal_w\[0\]
+ edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.bypass_in edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.out
+ VSS VDD VSS VDD sky130_fd_sc_hd__and2b_1
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[4\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[4\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[5\] VSS VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[4\].delay_unit/mid
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[4\].delay_unit/a_1632_71#
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[4\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_inbuf_1_A ena_in VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_3_235 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_19_125 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_15_29 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[2\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[2\]
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[3\] VSS VDD clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[2\].delay_unit/mid
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[2\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[2\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_2.genblk1\[0\].dly_binary.genblk1\[0\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[0\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_2.genblk1\[0\].dly_binary.signal_w\[1\] VSS VDD clkgen.delay_155ns_2.genblk1\[0\].dly_binary.genblk1\[0\].delay_unit/mid
+ clkgen.delay_155ns_2.genblk1\[0\].dly_binary.genblk1\[0\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_2.genblk1\[0\].dly_binary.genblk1\[0\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XPHY_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_7_63 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_16_94 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xinbuf_3 VSS VDD clkgen.delay_155ns_1.genblk1\[0\].dly_binary.in ndecision_finish_in
+ VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_12_164 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_4_330 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA_edgedetect.dly_315ns_1.genblk1\[5\].control_invert_A dlycontrol4_in[5] VSS
+ VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsampledly33 VDD VSS nsample_p_3 nsample_p_4 VSS VDD sampledly33/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1
Xedgedetect.dly_315ns_1.genblk1\[4\].control_invert dlycontrol4_in[4] edgedetect.dly_315ns_1.bypass_enable_w\[4\]
+ VDD VSS VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_17_256 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_17_223 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xsampledly11 VDD VSS sample_p_1 sample_p_2 VSS VDD sampledly11/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1
XFILLER_1_311 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xsampledly22 VDD VSS sample_n_2 sample_n_3 VSS VDD sampledly22/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[9\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[9\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[10\] VSS VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[9\].delay_unit/mid
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[9\].delay_unit/a_1632_71#
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[9\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_clkgen.delay_155ns_2.genblk1\[0\].dly_binary.and_bypass_switch_B clkgen.clk_dig_out
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_13_281 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[13\]
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[14\] VSS VDD clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit/mid
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[7\]
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[8\] VSS VDD clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit/mid
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XFILLER_10_284 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_6_244 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_1_32 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_19_94 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[1\]
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[2\] VSS VDD clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit/mid
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_3.genblk1\[0\].bypass_enable VDD VSS clkgen.delay_155ns_3.genblk1\[0\].dly_binary.bypass_in
+ clkgen.delay_155ns_3.bypass_enable_w\[0\] clkgen.delay_155ns_3.enable_dlycontrol_w
+ VSS VDD sky130_fd_sc_hd__and2_1
XFILLER_0_206 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_2_280 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_12_302 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[1\].dly_binary.out_mux VSS VDD clkgen.delay_155ns_3.genblk1\[1\].dly_binary.bypass_in
+ clkgen.delay_155ns_3.genblk1\[0\].dly_binary.out clkgen.delay_155ns_3.genblk1\[1\].dly_binary.signal_w\[2\]
+ clkgen.delay_155ns_3.genblk1\[1\].dly_binary.out VSS VDD clkgen.delay_155ns_3.genblk1\[1\].dly_binary.out_mux/a_505_21#
+ sky130_fd_sc_hd__mux2_1
XPHY_4 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_12_143 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[3\].dly_binary.out_mux VSS VDD clkgen.delay_155ns_3.genblk1\[3\].dly_binary.bypass_in
+ clkgen.delay_155ns_3.genblk1\[2\].dly_binary.out clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[8\]
+ clkgen.delay_155ns_3.genblk1\[3\].dly_binary.out VSS VDD clkgen.delay_155ns_3.genblk1\[3\].dly_binary.out_mux/a_505_21#
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_301 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_1_323 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xsampledly23 VDD VSS nsample_p_2 nsample_p_3 VSS VDD sampledly23/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[4\]
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[5\] VSS VDD edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit/mid
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit/a_1632_71#
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
Xsampledly01 VDD VSS sample_p_in sample_p_1 VSS VDD sampledly01/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1
Xsampledly34 VDD VSS nsample_n_3 nsample_n_4 VSS VDD sampledly34/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1
XFILLER_4_32 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xsampledly12 VDD VSS sample_n_1 sample_n_2 VSS VDD sampledly12/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1
Xclkgen.delay_155ns_3.genblk1\[4\].control_invert dlycontrol3_in[4] clkgen.delay_155ns_3.bypass_enable_w\[4\]
+ VDD VSS VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_13_63 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[6\]
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[7\] VSS VDD clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit/mid
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[2\].dly_binary.and_bypass_switch edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[0\]
+ edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.bypass_in edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.out
+ VSS VDD VSS VDD sky130_fd_sc_hd__and2b_1
XFILLER_13_293 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_9_275 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_9_220 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_1_175 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.delay_155ns_2.genblk1\[4\].dly_binary.out_mux_S clkgen.delay_155ns_2.genblk1\[4\].dly_binary.bypass_in
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_11_219 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[2\]
+ clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[3\] VSS VDD clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit/mid
+ clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XFILLER_6_201 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.delay_155ns_1.genblk1\[0\].control_invert_A dlycontrol1_in[0] VSS
+ VDD VDD VSS sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[0\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[1\] VSS VDD clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[0\].delay_unit/mid
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[0\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[0\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XFILLER_3_215 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_2_270 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_2_292 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[11\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[11\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[12\] VSS VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[11\].delay_unit/mid
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[11\].delay_unit/a_1632_71#
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[11\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XFILLER_8_307 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[11\]
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[12\] VSS VDD clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit/mid
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[9\]
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[10\] VSS VDD edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit/mid
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit/a_1632_71#
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XPHY_5 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_7_32 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_16_63 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_12_199 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[7\]
+ clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[8\] VSS VDD clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit/mid
+ clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[12\]
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[13\] VSS VDD edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit/mid
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit/a_1632_71#
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XFILLER_1_335 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[5\]
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[6\] VSS VDD clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit/mid
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
Xsampledly13 VDD VSS nsample_p_1 nsample_p_2 VSS VDD sampledly13/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1
Xsampledly24 VDD VSS nsample_n_2 nsample_n_3 VSS VDD sampledly24/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1
Xsampledly02 VDD VSS sample_n_in sample_n_1 VSS VDD sampledly02/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1
Xclkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[1\]
+ clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[2\] VSS VDD clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit/mid
+ clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XFILLER_9_243 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_1_143 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[16\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[16\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[17\] VSS VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[16\].delay_unit/mid
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[16\].delay_unit/a_1632_71#
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[16\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.and_bypass_switch_A_N edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.bypass_in
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_19_63 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_10_87 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xclkgen.delay_155ns_1.genblk1\[0\].control_invert dlycontrol1_in[0] clkgen.delay_155ns_1.bypass_enable_w\[0\]
+ VDD VSS VSS VDD sky130_fd_sc_hd__inv_2
Xedgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[4\]
+ edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[5\] VSS VDD edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit/mid
+ edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit/a_1632_71#
+ edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XPHY_6 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xclkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[6\]
+ clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[7\] VSS VDD clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit/mid
+ clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_3.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[2\].dly_binary.signal_w\[2\]
+ clkgen.delay_155ns_3.genblk1\[2\].dly_binary.signal_w\[3\] VSS VDD clkgen.delay_155ns_3.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit/mid
+ clkgen.delay_155ns_3.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_3.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[3\].dly_binary.and_bypass_switch edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[0\]
+ edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.bypass_in edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.out
+ VSS VDD VSS VDD sky130_fd_sc_hd__and2b_1
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[23\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[23\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[24\] VSS VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[23\].delay_unit/mid
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[23\].delay_unit/a_1632_71#
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[23\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
Xsampledly03 VDD VSS nsample_p_in nsample_p_1 VSS VDD sampledly03/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1
Xsampledly14 VDD VSS nsample_n_1 nsample_n_2 VSS VDD sampledly14/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1
Xclkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[0\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[1\] VSS VDD clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[0\].delay_unit/mid
+ clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[0\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[0\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XFILLER_4_196 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_13_32 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_8_3 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_1_133 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_10_210 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_18_310 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.out_mux_S edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.bypass_in
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_10_77 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[28\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[28\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[29\] VSS VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[28\].delay_unit/mid
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[28\].delay_unit/a_1632_71#
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[28\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[5\]
+ clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[6\] VSS VDD clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit/mid
+ clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XFILLER_15_143 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[30\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[30\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[31\] VSS VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[30\].delay_unit/mid
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[30\].delay_unit/a_1632_71#
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[30\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XFILLER_12_338 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA_clkgen.delay_155ns_2.genblk1\[0\].dly_binary.out_mux_S clkgen.delay_155ns_2.genblk1\[0\].dly_binary.bypass_in
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XPHY_7 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xclkgen.delay_155ns_2.genblk1\[2\].dly_binary.genblk1\[1\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[1\]
+ clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[2\] VSS VDD clkgen.delay_155ns_2.genblk1\[2\].dly_binary.genblk1\[1\].delay_unit/mid
+ clkgen.delay_155ns_2.genblk1\[2\].dly_binary.genblk1\[1\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_2.genblk1\[2\].dly_binary.genblk1\[1\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XFILLER_16_32 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_12_102 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsampledly04 VDD VSS nsample_n_in nsample_n_1 VSS VDD sampledly04/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1
XFILLER_4_164 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_10_244 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_18_322 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_3_229 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_5_281 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_19_32 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_2_240 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_18_174 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_18_152 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xedgedetect.dly_315ns_1.enablebuffer VDD VSS edgedetect.dly_315ns_1.enable_dlycontrol_w
+ enable_dlycontrol_in VSS VDD edgedetect.dly_315ns_1.enablebuffer/a_27_47# sky130_fd_sc_hd__buf_4
XANTENNA_edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.out_mux_S edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.bypass_in
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_1.genblk1\[2\].dly_binary.genblk1\[0\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[1\] VSS VDD clkgen.delay_155ns_1.genblk1\[2\].dly_binary.genblk1\[0\].delay_unit/mid
+ clkgen.delay_155ns_1.genblk1\[2\].dly_binary.genblk1\[0\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_1.genblk1\[2\].dly_binary.genblk1\[0\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.and_bypass_switch edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[0\]
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.bypass_in edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.out
+ VSS VDD VSS VDD sky130_fd_sc_hd__and2b_1
XFILLER_16_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_15_133 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_8 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_11_191 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_edgedetect.dly_315ns_1.genblk1\[4\].control_invert_A dlycontrol4_in[4] VSS
+ VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_17_239 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_16_272 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xclkgen.delay_155ns_1.enablebuffer VDD VSS clkgen.delay_155ns_1.enable_dlycontrol_w
+ enable_dlycontrol_in VSS VDD clkgen.delay_155ns_1.enablebuffer/a_27_47# sky130_fd_sc_hd__buf_4
Xedgedetect.dly_315ns_1.genblk1\[3\].bypass_enable VDD VSS edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.bypass_in
+ edgedetect.dly_315ns_1.bypass_enable_w\[3\] edgedetect.dly_315ns_1.enable_dlycontrol_w
+ VSS VDD sky130_fd_sc_hd__and2_1
XFILLER_13_275 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_10_201 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_2.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[1\].dly_binary.signal_w\[1\]
+ clkgen.delay_155ns_2.genblk1\[1\].dly_binary.signal_w\[2\] VSS VDD clkgen.delay_155ns_2.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit/mid
+ clkgen.delay_155ns_2.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_2.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_2.genblk1\[1\].control_invert dlycontrol2_in[1] clkgen.delay_155ns_2.bypass_enable_w\[1\]
+ VDD VSS VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_5_293 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_15_337 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_18_164 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[4\].bypass_enable VDD VSS clkgen.delay_155ns_1.genblk1\[4\].dly_binary.bypass_in
+ clkgen.delay_155ns_1.bypass_enable_w\[4\] clkgen.delay_155ns_1.enable_dlycontrol_w
+ VSS VDD sky130_fd_sc_hd__and2_1
XFILLER_2_252 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[0\].dly_binary.and_bypass_switch clkgen.delay_155ns_3.genblk1\[0\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_3.genblk1\[0\].dly_binary.bypass_in clkgen.delay_155ns_3.genblk1\[0\].dly_binary.in
+ VSS VDD VSS VDD sky130_fd_sc_hd__and2b_1
XPHY_9 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[11\]
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[12\] VSS VDD clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit/mid
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.out_mux_S edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.bypass_in
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_12_115 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.delay_155ns_1.enablebuffer_A enable_dlycontrol_in VSS VDD VDD VSS
+ sky130_fd_sc_hd__diode_2
XANTENNA_clkgen.delay_155ns_1.genblk1\[4\].dly_binary.out_mux_A0 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[16\]
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_19_292 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[0\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[0\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[1\] VSS VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[0\].delay_unit/mid
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[0\].delay_unit/a_1632_71#
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[0\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XFILLER_13_287 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_9_236 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_8_280 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xclkgen.delay_155ns_1.genblk1\[1\].dly_binary.genblk1\[0\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[1\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_1.genblk1\[1\].dly_binary.signal_w\[1\] VSS VDD clkgen.delay_155ns_1.genblk1\[1\].dly_binary.genblk1\[0\].delay_unit/mid
+ clkgen.delay_155ns_1.genblk1\[1\].dly_binary.genblk1\[0\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_1.genblk1\[1\].dly_binary.genblk1\[0\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.and_bypass_switch edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[0\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.bypass_in edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.out
+ VSS VDD VSS VDD sky130_fd_sc_hd__and2b_1
XFILLER_10_36 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_2_264 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_12_308 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[5\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[5\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[6\] VSS VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[5\].delay_unit/mid
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[5\].delay_unit/a_1632_71#
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[5\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[2\].control_invert dlycontrol4_in[2] edgedetect.dly_315ns_1.bypass_enable_w\[2\]
+ VDD VSS VSS VDD sky130_fd_sc_hd__inv_2
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[3\]
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[4\] VSS VDD clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit/mid
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XFILLER_4_16 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_13_299 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_0_192 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_2.genblk1\[0\].bypass_enable VDD VSS clkgen.delay_155ns_2.genblk1\[0\].dly_binary.bypass_in
+ clkgen.delay_155ns_2.bypass_enable_w\[0\] clkgen.delay_155ns_2.enable_dlycontrol_w
+ VSS VDD sky130_fd_sc_hd__and2_1
Xclkgen.delay_155ns_3.genblk1\[1\].bypass_enable VDD VSS clkgen.delay_155ns_3.genblk1\[1\].dly_binary.bypass_in
+ clkgen.delay_155ns_3.bypass_enable_w\[1\] clkgen.delay_155ns_3.enable_dlycontrol_w
+ VSS VDD sky130_fd_sc_hd__and2_1
Xclkgen.delay_155ns_3.genblk1\[1\].dly_binary.and_bypass_switch clkgen.delay_155ns_3.genblk1\[1\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_3.genblk1\[1\].dly_binary.bypass_in clkgen.delay_155ns_3.genblk1\[0\].dly_binary.out
+ VSS VDD VSS VDD sky130_fd_sc_hd__and2b_1
XFILLER_2_276 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[8\]
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[9\] VSS VDD clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit/mid
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_clkgen.delay_155ns_3.genblk1\[4\].control_invert_A dlycontrol3_in[4] VSS
+ VDD VDD VSS sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[14\]
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[15\] VSS VDD clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit/mid
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_2.genblk1\[0\].dly_binary.and_bypass_switch clkgen.delay_155ns_2.genblk1\[0\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_2.genblk1\[0\].dly_binary.bypass_in clkgen.clk_dig_out VSS VDD
+ VSS VDD sky130_fd_sc_hd__and2b_1
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[0\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[0\]
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[1\] VSS VDD edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[0\].delay_unit/mid
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[0\].delay_unit/a_1632_71#
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[0\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[2\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[2\]
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[3\] VSS VDD clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[2\].delay_unit/mid
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[2\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[2\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XFILLER_4_338 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_11_183 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_7_187 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[0\].dly_binary.genblk1\[0\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[0\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_1.genblk1\[0\].dly_binary.signal_w\[1\] VSS VDD clkgen.delay_155ns_1.genblk1\[0\].dly_binary.genblk1\[0\].delay_unit/mid
+ clkgen.delay_155ns_1.genblk1\[0\].dly_binary.genblk1\[0\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_1.genblk1\[0\].dly_binary.genblk1\[0\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XFILLER_19_261 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[2\].control_invert dlycontrol3_in[2] clkgen.delay_155ns_3.bypass_enable_w\[2\]
+ VDD VSS VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_13_245 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_182 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_18_304 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[5\]
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[6\] VSS VDD edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit/mid
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit/a_1632_71#
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XFILLER_5_241 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_10_49 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_10_16 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[7\]
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[8\] VSS VDD clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit/mid
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XFILLER_2_222 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[3\]
+ clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[4\] VSS VDD clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit/mid
+ clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XFILLER_7_303 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[1\]
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[2\] VSS VDD clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit/mid
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XFILLER_16_15 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_4_306 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_7_155 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[12\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[12\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[13\] VSS VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[12\].delay_unit/mid
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[12\].delay_unit/a_1632_71#
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[12\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_2.genblk1\[1\].dly_binary.out_mux VSS VDD clkgen.delay_155ns_2.genblk1\[1\].dly_binary.bypass_in
+ clkgen.delay_155ns_2.genblk1\[0\].dly_binary.out clkgen.delay_155ns_2.genblk1\[1\].dly_binary.signal_w\[2\]
+ clkgen.delay_155ns_2.genblk1\[1\].dly_binary.out VSS VDD clkgen.delay_155ns_2.genblk1\[1\].dly_binary.out_mux/a_505_21#
+ sky130_fd_sc_hd__mux2_1
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[12\]
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[13\] VSS VDD clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit/mid
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XFILLER_4_125 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.and_bypass_switch_A_N edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.bypass_in
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_16_210 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xclkgen.delay_155ns_2.genblk1\[3\].dly_binary.out_mux VSS VDD clkgen.delay_155ns_2.genblk1\[3\].dly_binary.bypass_in
+ clkgen.delay_155ns_2.genblk1\[2\].dly_binary.out clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[8\]
+ clkgen.delay_155ns_2.genblk1\[3\].dly_binary.out VSS VDD clkgen.delay_155ns_2.genblk1\[3\].dly_binary.out_mux/a_505_21#
+ sky130_fd_sc_hd__mux2_1
Xclkgen.delay_155ns_3.genblk1\[2\].dly_binary.and_bypass_switch clkgen.delay_155ns_3.genblk1\[2\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_3.genblk1\[2\].dly_binary.bypass_in clkgen.delay_155ns_3.genblk1\[1\].dly_binary.out
+ VSS VDD VSS VDD sky130_fd_sc_hd__and2b_1
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[13\]
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[14\] VSS VDD edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit/mid
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit/a_1632_71#
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XFILLER_12_290 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_8_272 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_18_316 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[0\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[0\]
+ edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[1\] VSS VDD edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[0\].delay_unit/mid
+ edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[0\].delay_unit/a_1632_71#
+ edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[0\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[6\]
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[7\] VSS VDD clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit/mid
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_2.genblk1\[1\].dly_binary.and_bypass_switch clkgen.delay_155ns_2.genblk1\[1\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_2.genblk1\[1\].dly_binary.bypass_in clkgen.delay_155ns_2.genblk1\[0\].dly_binary.out
+ VSS VDD VSS VDD sky130_fd_sc_hd__and2b_1
Xclkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[2\]
+ clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[3\] VSS VDD clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit/mid
+ clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XFILLER_5_275 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_2_234 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_4_3 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_18_124 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[17\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[17\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[18\] VSS VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[17\].delay_unit/mid
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[17\].delay_unit/a_1632_71#
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[17\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_1.genblk1\[0\].dly_binary.and_bypass_switch clkgen.delay_155ns_1.genblk1\[0\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_1.genblk1\[0\].dly_binary.bypass_in clkgen.delay_155ns_1.genblk1\[0\].dly_binary.in
+ VSS VDD VSS VDD sky130_fd_sc_hd__and2b_1
XFILLER_11_311 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_7_337 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_14_182 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_4_318 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xedgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[5\]
+ edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[6\] VSS VDD edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit/mid
+ edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit/a_1632_71#
+ edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XFILLER_16_244 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[7\]
+ clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[8\] VSS VDD clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit/mid
+ clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_edgedetect.dly_315ns_1.genblk1\[3\].control_invert_A dlycontrol4_in[3] VSS
+ VDD VDD VSS sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_1.genblk1\[3\].control_invert dlycontrol1_in[3] clkgen.delay_155ns_1.bypass_enable_w\[3\]
+ VDD VSS VSS VDD sky130_fd_sc_hd__inv_2
XANTENNA_edgedetect.nor1_A edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.out VSS
+ VDD VDD VSS sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_3.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[2\].dly_binary.signal_w\[3\]
+ clkgen.delay_155ns_3.genblk1\[2\].dly_binary.signal_w\[4\] VSS VDD clkgen.delay_155ns_3.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit/mid
+ clkgen.delay_155ns_3.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_3.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XFILLER_9_229 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_0_173 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[24\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[24\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[25\] VSS VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[24\].delay_unit/mid
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[24\].delay_unit/a_1632_71#
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[24\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XFILLER_5_84 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_18_328 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xclkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[1\]
+ clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[2\] VSS VDD clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit/mid
+ clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XFILLER_5_287 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_2_202 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_2_246 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_19_275 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[29\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[29\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[30\] VSS VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[29\].delay_unit/mid
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[29\].delay_unit/a_1632_71#
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[29\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[2\].dly_binary.genblk1\[0\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[0\]
+ edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[1\] VSS VDD edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.genblk1\[0\].delay_unit/mid
+ edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.genblk1\[0\].delay_unit/a_1632_71#
+ edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.genblk1\[0\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_3.genblk1\[3\].dly_binary.and_bypass_switch clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_3.genblk1\[3\].dly_binary.bypass_in clkgen.delay_155ns_3.genblk1\[2\].dly_binary.out
+ VSS VDD VSS VDD sky130_fd_sc_hd__and2b_1
Xclkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[6\]
+ clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[7\] VSS VDD clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit/mid
+ clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XFILLER_17_71 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[31\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[31\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[32\] VSS VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[31\].delay_unit/mid
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[31\].delay_unit/a_1632_71#
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[31\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XFILLER_0_311 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xclkgen.delay_155ns_2.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[2\]
+ clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[3\] VSS VDD clkgen.delay_155ns_2.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit/mid
+ clkgen.delay_155ns_2.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_2.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XFILLER_12_3 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_2.genblk1\[2\].dly_binary.and_bypass_switch clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_2.genblk1\[2\].dly_binary.bypass_in clkgen.delay_155ns_2.genblk1\[1\].dly_binary.out
+ VSS VDD VSS VDD sky130_fd_sc_hd__and2b_1
Xclkgen.delay_155ns_1.genblk1\[1\].dly_binary.and_bypass_switch clkgen.delay_155ns_1.genblk1\[1\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_1.genblk1\[1\].dly_binary.bypass_in clkgen.delay_155ns_1.genblk1\[0\].dly_binary.out
+ VSS VDD VSS VDD sky130_fd_sc_hd__and2b_1
XFILLER_5_299 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_2_258 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_sampledly03_A nsample_p_in VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_7_125 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xclkgen.delay_155ns_1.genblk1\[2\].dly_binary.genblk1\[1\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[1\]
+ clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[2\] VSS VDD clkgen.delay_155ns_1.genblk1\[2\].dly_binary.genblk1\[1\].delay_unit/mid
+ clkgen.delay_155ns_1.genblk1\[2\].dly_binary.genblk1\[1\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_1.genblk1\[2\].dly_binary.genblk1\[1\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[4\].bypass_enable VDD VSS edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.bypass_in
+ edgedetect.dly_315ns_1.bypass_enable_w\[4\] edgedetect.dly_315ns_1.enable_dlycontrol_w
+ VSS VDD sky130_fd_sc_hd__and2_1
XFILLER_0_323 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_0_164 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_5_75 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.delay_155ns_2.genblk1\[4\].control_invert_A dlycontrol2_in[4] VSS
+ VDD VDD VSS sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_2.enablebuffer VDD VSS clkgen.delay_155ns_2.enable_dlycontrol_w
+ enable_dlycontrol_in VSS VDD clkgen.delay_155ns_2.enablebuffer/a_27_47# sky130_fd_sc_hd__buf_4
Xedgedetect.dly_315ns_1.genblk1\[1\].dly_binary.genblk1\[0\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.signal_w\[0\]
+ edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.signal_w\[1\] VSS VDD edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.genblk1\[0\].delay_unit/mid
+ edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.genblk1\[0\].delay_unit/a_1632_71#
+ edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.genblk1\[0\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.and_bypass_switch clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.bypass_in clkgen.delay_155ns_3.genblk1\[3\].dly_binary.out
+ VSS VDD VSS VDD sky130_fd_sc_hd__and2b_1
XANTENNA_edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.out_mux_A0 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[32\]
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_clkgen.delay_155ns_3.genblk1\[3\].control_invert_A dlycontrol3_in[3] VSS
+ VDD VDD VSS sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_2.genblk1\[4\].control_invert dlycontrol2_in[4] clkgen.delay_155ns_2.bypass_enable_w\[4\]
+ VDD VSS VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_11_155 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_2.genblk1\[3\].dly_binary.and_bypass_switch clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_2.genblk1\[3\].dly_binary.bypass_in clkgen.delay_155ns_2.genblk1\[2\].dly_binary.out
+ VSS VDD VSS VDD sky130_fd_sc_hd__and2b_1
XFILLER_8_86 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_0_335 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xclkgen.delay_155ns_1.genblk1\[2\].dly_binary.and_bypass_switch clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_1.genblk1\[2\].dly_binary.bypass_in clkgen.delay_155ns_1.genblk1\[1\].dly_binary.out
+ VSS VDD VSS VDD sky130_fd_sc_hd__and2b_1
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[12\]
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[13\] VSS VDD clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit/mid
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XFILLER_3_151 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_13_217 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_12_261 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_8_210 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_0_143 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_0_121 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_5_32 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_14_63 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_5_213 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[1\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[1\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[2\] VSS VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[1\].delay_unit/mid
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[1\].delay_unit/a_1632_71#
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[1\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_clkgen.delay_155ns_2.genblk1\[0\].dly_binary.and_bypass_switch_A_N clkgen.delay_155ns_2.genblk1\[0\].dly_binary.bypass_in
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_17_194 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_14_334 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_1_271 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[1\].dly_binary.signal_w\[1\]
+ clkgen.delay_155ns_1.genblk1\[1\].dly_binary.signal_w\[2\] VSS VDD clkgen.delay_155ns_1.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit/mid
+ clkgen.delay_155ns_1.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_1.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XFILLER_3_311 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xedgedetect.dly_315ns_1.genblk1\[0\].control_invert dlycontrol4_in[0] edgedetect.dly_315ns_1.bypass_enable_w\[0\]
+ VDD VSS VSS VDD sky130_fd_sc_hd__inv_2
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[6\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[6\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[7\] VSS VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[6\].delay_unit/mid
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[6\].delay_unit/a_1632_71#
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[6\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_1.genblk1\[0\].bypass_enable VDD VSS clkgen.delay_155ns_1.genblk1\[0\].dly_binary.bypass_in
+ clkgen.delay_155ns_1.bypass_enable_w\[0\] clkgen.delay_155ns_1.enable_dlycontrol_w
+ VSS VDD sky130_fd_sc_hd__and2_1
Xedgedetect.dly_315ns_1.genblk1\[0\].dly_binary.genblk1\[0\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.signal_w\[0\]
+ edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.signal_w\[1\] VSS VDD edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.genblk1\[0\].delay_unit/mid
+ edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.genblk1\[0\].delay_unit/a_1632_71#
+ edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.genblk1\[0\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_2.genblk1\[1\].bypass_enable VDD VSS clkgen.delay_155ns_2.genblk1\[1\].dly_binary.bypass_in
+ clkgen.delay_155ns_2.bypass_enable_w\[1\] clkgen.delay_155ns_2.enable_dlycontrol_w
+ VSS VDD sky130_fd_sc_hd__and2_1
XFILLER_0_199 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_0_133 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_12_284 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_12_273 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xclkgen.delay_155ns_3.genblk1\[2\].bypass_enable VDD VSS clkgen.delay_155ns_3.genblk1\[2\].dly_binary.bypass_in
+ clkgen.delay_155ns_3.bypass_enable_w\[2\] clkgen.delay_155ns_3.enable_dlycontrol_w
+ VSS VDD sky130_fd_sc_hd__and2_1
XFILLER_10_3 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_8_244 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[4\]
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[5\] VSS VDD clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit/mid
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[10\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[10\]
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[11\] VSS VDD clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[10\].delay_unit/mid
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[10\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[10\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[5\].control_invert dlycontrol4_in[5] edgedetect.dly_315ns_1.bypass_enable_w\[5\]
+ VDD VSS VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_2_228 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_30 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_17_151 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.and_bypass_switch clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.bypass_in clkgen.delay_155ns_2.genblk1\[3\].dly_binary.out
+ VSS VDD VSS VDD sky130_fd_sc_hd__and2b_1
XFILLER_11_305 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_11_32 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.delay_155ns_1.genblk1\[3\].dly_binary.and_bypass_switch_A_N clkgen.delay_155ns_1.genblk1\[3\].dly_binary.bypass_in
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_1.genblk1\[3\].dly_binary.and_bypass_switch clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_1.genblk1\[3\].dly_binary.bypass_in clkgen.delay_155ns_1.genblk1\[2\].dly_binary.out
+ VSS VDD VSS VDD sky130_fd_sc_hd__and2b_1
XANTENNA_sampledly01_A sample_p_in VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[9\]
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[10\] VSS VDD clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit/mid
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XFILLER_3_323 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[15\]
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[16\] VSS VDD clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit/mid
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[1\]
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[2\] VSS VDD edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit/mid
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit/a_1632_71#
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XFILLER_17_86 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[0\].control_invert dlycontrol3_in[0] clkgen.delay_155ns_3.bypass_enable_w\[0\]
+ VDD VSS VSS VDD sky130_fd_sc_hd__inv_2
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[3\]
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[4\] VSS VDD clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit/mid
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XFILLER_12_296 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_edgedetect.dly_315ns_1.genblk1\[2\].control_invert_A dlycontrol4_in[2] VSS
+ VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_8_201 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_14_32 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XPHY_31 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_20 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[6\]
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[7\] VSS VDD edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit/mid
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit/a_1632_71#
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[1\].dly_binary.out_mux VSS VDD edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.bypass_in
+ edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.out edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.signal_w\[2\]
+ edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.out VSS VDD edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.out_mux/a_505_21#
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_144 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[8\]
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[9\] VSS VDD clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit/mid
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[3\].dly_binary.out_mux VSS VDD edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.bypass_in
+ edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.out edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[8\]
+ edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.out VSS VDD edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.out_mux/a_505_21#
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_192 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_9_181 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_inbuf_2_A start_conv_in VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.out_mux VSS VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.bypass_in
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.out edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[32\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.out VSS VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.out_mux/a_505_21#
+ sky130_fd_sc_hd__mux2_1
Xclkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[4\]
+ clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[5\] VSS VDD clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit/mid
+ clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XFILLER_11_125 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_3_335 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_6_173 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_17_32 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[2\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[2\]
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[3\] VSS VDD clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[2\].delay_unit/mid
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[2\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[2\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XFILLER_3_187 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_0_90 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA_clkgen.delay_155ns_1.genblk1\[3\].dly_binary.out_mux_S clkgen.delay_155ns_1.genblk1\[3\].dly_binary.bypass_in
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[13\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[13\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[14\] VSS VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[13\].delay_unit/mid
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[13\].delay_unit/a_1632_71#
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[13\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[13\]
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[14\] VSS VDD clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit/mid
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XPHY_32 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_21 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.and_bypass_switch clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.bypass_in clkgen.delay_155ns_1.genblk1\[3\].dly_binary.out
+ VSS VDD VSS VDD sky130_fd_sc_hd__and2b_1
XPHY_10 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[14\]
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[15\] VSS VDD edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit/mid
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit/a_1632_71#
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.and_bypass_switch_A_N edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.bypass_in
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_2_58 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xedgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[1\]
+ edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[2\] VSS VDD edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit/mid
+ edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit/a_1632_71#
+ edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XFILLER_11_89 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xoutbuf_1 VDD VSS clk_dig_out clkgen.clk_dig_out VSS VDD outbuf_1/a_27_47# sky130_fd_sc_hd__buf_4
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[7\]
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[8\] VSS VDD clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit/mid
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XFILLER_14_134 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[3\]
+ clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[4\] VSS VDD clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit/mid
+ clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[18\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[18\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[19\] VSS VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[18\].delay_unit/mid
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[18\].delay_unit/a_1632_71#
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[18\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XFILLER_3_303 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_18_292 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.delay_155ns_1.genblk1\[4\].control_invert_A dlycontrol1_in[4] VSS
+ VDD VDD VSS sky130_fd_sc_hd__diode_2
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[20\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[20\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[21\] VSS VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[20\].delay_unit/mid
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[20\].delay_unit/a_1632_71#
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[20\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XFILLER_15_240 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[1\].control_invert dlycontrol1_in[1] clkgen.delay_155ns_1.bypass_enable_w\[1\]
+ VDD VSS VSS VDD sky130_fd_sc_hd__inv_2
Xclkgen.delay_155ns_1.genblk1\[1\].dly_binary.out_mux VSS VDD clkgen.delay_155ns_1.genblk1\[1\].dly_binary.bypass_in
+ clkgen.delay_155ns_1.genblk1\[0\].dly_binary.out clkgen.delay_155ns_1.genblk1\[1\].dly_binary.signal_w\[2\]
+ clkgen.delay_155ns_1.genblk1\[1\].dly_binary.out VSS VDD clkgen.delay_155ns_1.genblk1\[1\].dly_binary.out_mux/a_505_21#
+ sky130_fd_sc_hd__mux2_1
Xedgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[6\]
+ edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[7\] VSS VDD edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit/mid
+ edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit/a_1632_71#
+ edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_1.genblk1\[3\].dly_binary.out_mux VSS VDD clkgen.delay_155ns_1.genblk1\[3\].dly_binary.bypass_in
+ clkgen.delay_155ns_1.genblk1\[2\].dly_binary.out clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[8\]
+ clkgen.delay_155ns_1.genblk1\[3\].dly_binary.out VSS VDD clkgen.delay_155ns_1.genblk1\[3\].dly_binary.out_mux/a_505_21#
+ sky130_fd_sc_hd__mux2_1
XANTENNA_clkgen.delay_155ns_2.genblk1\[3\].control_invert_A dlycontrol2_in[3] VSS
+ VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.and_bypass_switch_B edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.out
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_4_272 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XPHY_33 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_22 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_2_209 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_17_121 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_1_253 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[25\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[25\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[26\] VSS VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[25\].delay_unit/mid
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[25\].delay_unit/a_1632_71#
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[25\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[2\]
+ clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[3\] VSS VDD clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit/mid
+ clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
Xoutbuf_2 VDD VSS clk_comp_out clkgen.clk_comp_out VSS VDD outbuf_2/a_27_47# sky130_fd_sc_hd__buf_4
XFILLER_6_334 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA_clkgen.delay_155ns_3.genblk1\[2\].control_invert_A dlycontrol3_in[2] VSS
+ VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_8_58 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_6_164 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_0_307 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_12_255 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[2\].dly_binary.genblk1\[1\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[1\]
+ edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[2\] VSS VDD edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.genblk1\[1\].delay_unit/mid
+ edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.genblk1\[1\].delay_unit/a_1632_71#
+ edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.genblk1\[1\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[7\]
+ clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[8\] VSS VDD clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit/mid
+ clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XFILLER_17_303 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xclkgen.delay_155ns_2.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[3\]
+ clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[4\] VSS VDD clkgen.delay_155ns_2.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit/mid
+ clkgen.delay_155ns_2.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_2.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XPHY_12 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_34 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_14_306 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_23 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_1_221 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_1_265 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xoutbuf_3 VDD VSS sample_p_out sample_p_4 VSS VDD outbuf_3/a_27_47# sky130_fd_sc_hd__buf_4
Xclkgen.delay_155ns_3.genblk1\[0\].dly_binary.out_mux VSS VDD clkgen.delay_155ns_3.genblk1\[0\].dly_binary.bypass_in
+ clkgen.delay_155ns_3.genblk1\[0\].dly_binary.in clkgen.delay_155ns_3.genblk1\[0\].dly_binary.signal_w\[1\]
+ clkgen.delay_155ns_3.genblk1\[0\].dly_binary.out VSS VDD clkgen.delay_155ns_3.genblk1\[0\].dly_binary.out_mux/a_505_21#
+ sky130_fd_sc_hd__mux2_1
Xclkgen.delay_155ns_3.genblk1\[2\].dly_binary.out_mux VSS VDD clkgen.delay_155ns_3.genblk1\[2\].dly_binary.bypass_in
+ clkgen.delay_155ns_3.genblk1\[1\].dly_binary.out clkgen.delay_155ns_3.genblk1\[2\].dly_binary.signal_w\[4\]
+ clkgen.delay_155ns_3.genblk1\[2\].dly_binary.out VSS VDD clkgen.delay_155ns_3.genblk1\[2\].dly_binary.out_mux/a_505_21#
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_151 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA_outbuf_1_A clkgen.clk_dig_out VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xedgedetect.dly_315ns_1.genblk1\[5\].bypass_enable VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.bypass_in
+ edgedetect.dly_315ns_1.bypass_enable_w\[5\] edgedetect.dly_315ns_1.enable_dlycontrol_w
+ VSS VDD sky130_fd_sc_hd__and2_1
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.out_mux VSS VDD clkgen.delay_155ns_3.genblk1\[4\].dly_binary.bypass_in
+ clkgen.delay_155ns_3.genblk1\[3\].dly_binary.out clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[16\]
+ clkgen.clk_comp_out VSS VDD clkgen.delay_155ns_3.genblk1\[4\].dly_binary.out_mux/a_505_21#
+ sky130_fd_sc_hd__mux2_1
XFILLER_18_272 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_15_275 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_15_231 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_12_267 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[2\]
+ clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[3\] VSS VDD clkgen.delay_155ns_1.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit/mid
+ clkgen.delay_155ns_1.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_1.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XFILLER_17_337 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XPHY_35 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_24 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_9_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_13 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_1_233 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_1_277 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xoutbuf_4 VDD VSS sample_n_out sample_n_4 VSS VDD outbuf_4/a_27_47# sky130_fd_sc_hd__buf_4
Xclkgen.delay_155ns_3.enablebuffer VDD VSS clkgen.delay_155ns_3.enable_dlycontrol_w
+ enable_dlycontrol_in VSS VDD clkgen.delay_155ns_3.enablebuffer/a_27_47# sky130_fd_sc_hd__buf_4
Xclkgen.delay_155ns_2.genblk1\[2\].control_invert dlycontrol2_in[2] clkgen.delay_155ns_2.bypass_enable_w\[2\]
+ VDD VSS VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_19_218 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.signal_w\[1\]
+ edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.signal_w\[2\] VSS VDD edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit/mid
+ edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit/a_1632_71#
+ edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XFILLER_10_173 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_8_16 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.delay_155ns_2.genblk1\[4\].dly_binary.out_mux_A0 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[16\]
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_0_94 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA_edgedetect.dly_315ns_1.genblk1\[1\].control_invert_A dlycontrol4_in[1] VSS
+ VDD VDD VSS sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[13\]
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[14\] VSS VDD clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit/mid
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XPHY_36 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_25 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_1_245 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_1_201 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_14 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xedgedetect.dly_315ns_1.genblk1\[0\].bypass_enable VDD VSS edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.bypass_in
+ edgedetect.dly_315ns_1.bypass_enable_w\[0\] edgedetect.dly_315ns_1.enable_dlycontrol_w
+ VSS VDD sky130_fd_sc_hd__and2_1
XFILLER_1_289 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xoutbuf_5 VDD VSS nsample_p_out nsample_p_4 VSS VDD outbuf_5/a_27_47# sky130_fd_sc_hd__buf_4
XANTENNA_edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.out_mux_S edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.bypass_in
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[2\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[2\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[3\] VSS VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[2\].delay_unit/mid
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[2\].delay_unit/a_1632_71#
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[2\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XFILLER_11_119 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_3_94 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_18_285 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[1\].bypass_enable VDD VSS clkgen.delay_155ns_1.genblk1\[1\].dly_binary.bypass_in
+ clkgen.delay_155ns_1.bypass_enable_w\[1\] clkgen.delay_155ns_1.enable_dlycontrol_w
+ VSS VDD sky130_fd_sc_hd__and2_1
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[0\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[1\] VSS VDD clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[0\].delay_unit/mid
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[0\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[0\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_2.genblk1\[2\].bypass_enable VDD VSS clkgen.delay_155ns_2.genblk1\[2\].dly_binary.bypass_in
+ clkgen.delay_155ns_2.bypass_enable_w\[2\] clkgen.delay_155ns_2.enable_dlycontrol_w
+ VSS VDD sky130_fd_sc_hd__and2_1
XANTENNA_clkgen.delay_155ns_2.genblk1\[1\].dly_binary.out_mux_S clkgen.delay_155ns_2.genblk1\[1\].dly_binary.bypass_in
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_15_222 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_17_3 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[3\].bypass_enable VDD VSS clkgen.delay_155ns_3.genblk1\[3\].dly_binary.bypass_in
+ clkgen.delay_155ns_3.bypass_enable_w\[3\] clkgen.delay_155ns_3.enable_dlycontrol_w
+ VSS VDD sky130_fd_sc_hd__and2_1
XFILLER_0_107 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_12_225 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[7\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[7\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[8\] VSS VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[7\].delay_unit/mid
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[7\].delay_unit/a_1632_71#
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[7\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[3\].control_invert dlycontrol4_in[3] edgedetect.dly_315ns_1.bypass_enable_w\[3\]
+ VDD VSS VSS VDD sky130_fd_sc_hd__inv_2
XPHY_37 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_26 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_15 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_6_94 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_17_114 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[5\]
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[6\] VSS VDD clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit/mid
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[11\]
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[12\] VSS VDD clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit/mid
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
Xoutbuf_6 VDD VSS nsample_n_out nsample_n_4 VSS VDD outbuf_6/a_27_47# sky130_fd_sc_hd__buf_4
XFILLER_14_106 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_10_164 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.out_mux_S edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.bypass_in
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.out_mux_A0 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[16\]
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XANTENNA_clkgen.delay_155ns_1.genblk1\[3\].control_invert_A dlycontrol1_in[3] VSS
+ VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_9_94 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_0_63 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_5_19 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_11_281 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.delay_155ns_2.genblk1\[0\].dly_binary.out_mux_A1 clkgen.clk_dig_out
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[2\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[2\]
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[3\] VSS VDD edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[2\].delay_unit/mid
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[2\].delay_unit/a_1632_71#
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[2\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XFILLER_4_244 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_38 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_27 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA_clkgen.delay_155ns_2.genblk1\[2\].control_invert_A dlycontrol2_in[2] VSS
+ VDD VDD VSS sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[4\]
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[5\] VSS VDD clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit/mid
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XPHY_16 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_6_84 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[0\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[1\] VSS VDD clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[0\].delay_unit/mid
+ clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[0\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[0\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XFILLER_9_303 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xclkgen.delay_155ns_3.genblk1\[3\].control_invert dlycontrol3_in[3] clkgen.delay_155ns_3.bypass_enable_w\[3\]
+ VDD VSS VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_0_280 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_6_306 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.delay_155ns_3.enablebuffer_A enable_dlycontrol_in VSS VDD VDD VSS
+ sky130_fd_sc_hd__diode_2
XFILLER_7_3 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_3_63 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA_clkgen.delay_155ns_3.genblk1\[1\].control_invert_A dlycontrol3_in[1] VSS
+ VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_6_125 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_18_298 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[7\]
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[8\] VSS VDD edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit/mid
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit/a_1632_71#
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XFILLER_15_213 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.out_mux_A1 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.out
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[9\]
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[10\] VSS VDD clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit/mid
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.out_mux_S edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.bypass_in
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[5\]
+ clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[6\] VSS VDD clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit/mid
+ clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[10\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[10\]
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[11\] VSS VDD edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[10\].delay_unit/mid
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[10\].delay_unit/a_1632_71#
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[10\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.and_bypass_switch_A_N edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.bypass_in
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_11_293 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_7_275 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[3\]
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[4\] VSS VDD clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit/mid
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XPHY_28 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_17 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_39 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_13_311 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_1_215 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_1_259 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_16_182 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[14\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[14\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[15\] VSS VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[14\].delay_unit/mid
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[14\].delay_unit/a_1632_71#
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[14\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XFILLER_15_94 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_9_337 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[14\]
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[15\] VSS VDD clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit/mid
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XFILLER_11_19 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_10_325 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[15\]
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[16\] VSS VDD edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit/mid
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit/a_1632_71#
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XFILLER_18_244 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[2\]
+ edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[3\] VSS VDD edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit/mid
+ edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit/a_1632_71#
+ edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[8\]
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[9\] VSS VDD clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit/mid
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.and_bypass_switch_A_N edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.bypass_in
+ VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit VDD VSS clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[4\]
+ clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[5\] VSS VDD clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit/mid
+ clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_3.genblk1\[2\].dly_binary.genblk1\[0\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[2\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_3.genblk1\[2\].dly_binary.signal_w\[1\] VSS VDD clkgen.delay_155ns_3.genblk1\[2\].dly_binary.genblk1\[0\].delay_unit/mid
+ clkgen.delay_155ns_3.genblk1\[2\].dly_binary.genblk1\[0\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_3.genblk1\[2\].dly_binary.genblk1\[0\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XFILLER_9_63 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_18_94 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[19\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[19\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[20\] VSS VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[19\].delay_unit/mid
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[19\].delay_unit/a_1632_71#
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[19\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[21\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[21\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[22\] VSS VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[21\].delay_unit/mid
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[21\].delay_unit/a_1632_71#
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[21\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XFILLER_15_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_18 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_1_227 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[7\]
+ edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[8\] VSS VDD edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit/mid
+ edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit/a_1632_71#
+ edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XFILLER_0_293 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xclkgen.delay_155ns_1.genblk1\[4\].control_invert dlycontrol1_in[4] clkgen.delay_155ns_1.bypass_enable_w\[4\]
+ VDD VSS VSS VDD sky130_fd_sc_hd__inv_2
XFILLER_10_337 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_3_32 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[26\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[26\]
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[27\] VSS VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[26\].delay_unit/mid
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[26\].delay_unit/a_1632_71#
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[26\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[3\]
+ clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[4\] VSS VDD clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit/mid
+ clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XFILLER_5_182 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_2_174 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_7_244 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_4_214 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA_edgedetect.dly_315ns_1.genblk1\[0\].control_invert_A dlycontrol4_in[0] VSS
+ VDD VDD VSS sky130_fd_sc_hd__diode_2
XFILLER_6_43 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_9_9 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_1_239 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_15_63 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xedgedetect.dly_315ns_1.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit VDD VSS edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[2\]
+ edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[3\] VSS VDD edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit/mid
+ edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit/a_1632_71#
+ edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XFILLER_0_261 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_13_187 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xclkgen.delay_155ns_3.genblk1\[1\].dly_binary.genblk1\[0\].delay_unit VDD VSS clkgen.delay_155ns_3.genblk1\[1\].dly_binary.signal_w\[0\]
+ clkgen.delay_155ns_3.genblk1\[1\].dly_binary.signal_w\[1\] VSS VDD clkgen.delay_155ns_3.genblk1\[1\].dly_binary.genblk1\[0\].delay_unit/mid
+ clkgen.delay_155ns_3.genblk1\[1\].dly_binary.genblk1\[0\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_3.genblk1\[1\].dly_binary.genblk1\[0\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
XFILLER_5_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_2_164 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_9_32 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_18_63 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_12_208 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_19_182 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit VDD VSS clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[3\]
+ clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[4\] VSS VDD clkgen.delay_155ns_1.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit/mid
+ clkgen.delay_155ns_1.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit/a_1632_71#
+ clkgen.delay_155ns_1.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit/a_1691_329#
+ sky130_mm_sc_hd_dlyPoly5ns
C0 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[9\] sample_p_in 0.12fF
C1 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[11\].delay_unit/a_1691_329# VDD 0.11fF
C2 dlycontrol3_in[4] dlycontrol3_in[3] 0.66fF
C3 VDD clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[9\] 0.74fF
C4 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[16\] clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[14\] 0.13fF
C5 VDD clkgen.delay_155ns_3.bypass_enable_w\[3\] 0.86fF
C6 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit/mid VDD 0.17fF
C7 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[16\] edgedetect.dly_315ns_1.bypass_enable_w\[0\] 0.32fF
C8 clkgen.delay_155ns_2.genblk1\[0\].dly_binary.bypass_in VDD 3.00fF
C9 edgedetect.dly_315ns_1.enable_dlycontrol_w edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.bypass_in 0.48fF
C10 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[10\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[13\] 0.11fF
C11 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[16\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[0\].delay_unit/mid 0.16fF
C12 nsample_p_1 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.bypass_in 0.37fF
C13 edgedetect.dly_315ns_1.bypass_enable_w\[4\] edgedetect.dly_315ns_1.bypass_enable_w\[5\] 0.28fF
C14 clkgen.delay_155ns_3.genblk1\[2\].dly_binary.signal_w\[3\] clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[0\].delay_unit/mid 0.12fF
C15 clkgen.delay_155ns_1.genblk1\[1\].dly_binary.bypass_in clk_dig_out 0.15fF
C16 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[3\] clkgen.delay_155ns_3.genblk1\[4\].dly_binary.bypass_in 0.18fF
C17 clkgen.delay_155ns_3.genblk1\[1\].dly_binary.signal_w\[1\] clkgen.delay_155ns_3.genblk1\[2\].dly_binary.bypass_in 0.18fF
C18 dlycontrol1_in[4] clkgen.clk_comp_out 0.51fF
C19 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[0\] clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit/mid 0.10fF
C20 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.out clkgen.delay_155ns_1.genblk1\[0\].dly_binary.out 0.22fF
C21 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit/a_1632_71# clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[3\] 0.13fF
C22 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.bypass_in clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[8\] 0.11fF
C23 VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[19\].delay_unit/mid 0.50fF
C24 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.bypass_in dlycontrol2_in[4] 2.08fF
C25 clkgen.delay_155ns_2.genblk1\[1\].dly_binary.signal_w\[0\] clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[3\] 0.12fF
C26 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit/a_1632_71# clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[4\] 0.13fF
C27 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[5\] VDD 0.91fF
C28 clkgen.enable_loop_in clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[0\] 0.11fF
C29 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit/mid edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[2\] 0.22fF
C30 dlycontrol2_in[0] clkgen.delay_155ns_1.genblk1\[1\].dly_binary.out 0.75fF
C31 VDD clkgen.delay_155ns_1.bypass_enable_w\[1\] 0.66fF
C32 clkgen.delay_155ns_2.genblk1\[1\].dly_binary.signal_w\[0\] clkgen.delay_155ns_3.genblk1\[3\].dly_binary.out 0.10fF
C33 clkgen.delay_155ns_2.genblk1\[0\].dly_binary.bypass_in dlycontrol1_in[3] 0.13fF
C34 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.out sample_p_in 1.53fF
C35 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.bypass_in clkgen.delay_155ns_1.enable_dlycontrol_w 0.63fF
C36 dlycontrol3_in[2] start_conv_in 0.21fF
C37 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.bypass_in clkgen.delay_155ns_2.genblk1\[1\].dly_binary.signal_w\[0\] 2.10fF
C38 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.bypass_in dlycontrol2_in[3] 2.49fF
C39 edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.bypass_in dlycontrol4_in[2] 0.10fF
C40 clkgen.clk_dig_out clkgen.delay_155ns_2.genblk1\[0\].dly_binary.signal_w\[0\] 2.37fF
C41 sample_p_in edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.bypass_in 3.16fF
C42 clkgen.delay_155ns_3.genblk1\[2\].dly_binary.signal_w\[0\] dlycontrol3_in[3] 0.11fF
C43 sample_p_in edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.bypass_in 0.63fF
C44 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.bypass_in dlycontrol4_in[4] 0.19fF
C45 ena_in clkgen.delay_155ns_1.genblk1\[1\].dly_binary.bypass_in 0.14fF
C46 clkgen.delay_155ns_2.genblk1\[1\].dly_binary.signal_w\[1\] clkgen.delay_155ns_2.genblk1\[1\].dly_binary.bypass_in 0.30fF
C47 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit/mid clkgen.delay_155ns_2.genblk1\[4\].dly_binary.bypass_in 0.10fF
C48 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit/mid VDD 0.45fF
C49 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[10\] dlycontrol1_in[4] 0.33fF
C50 clkgen.delay_155ns_3.genblk1\[0\].dly_binary.bypass_in clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[4\] 0.30fF
C51 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[0\].delay_unit/mid VDD 0.26fF
C52 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[9\] dlycontrol3_in[1] 0.30fF
C53 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[16\] edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit/mid 0.11fF
C54 clkgen.clk_dig_out clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[2\] 0.20fF
C55 dlycontrol1_in[2] ena_in 4.36fF
C56 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[8\] enable_dlycontrol_in 4.48fF
C57 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit/mid edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[2\] 0.13fF
C58 edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.bypass_in edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[18\] 0.11fF
C59 dlycontrol4_in[4] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.out 0.45fF
C60 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.out clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[1\] 0.26fF
C61 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.out clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[16\] 0.44fF
C62 clkgen.delay_155ns_2.bypass_enable_w\[1\] clkgen.delay_155ns_2.enable_dlycontrol_w 0.16fF
C63 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit/mid clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[6\] 0.13fF
C64 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[4\] dlycontrol3_in[1] 0.33fF
C65 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.bypass_in clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[16\] 0.11fF
C66 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.bypass_in dlycontrol3_in[0] 0.13fF
C67 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[8\] VDD 1.34fF
C68 dlycontrol3_in[2] enable_dlycontrol_in 0.14fF
C69 clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[4\] sample_n_1 0.12fF
C70 sample_n_2 start_conv_in 0.15fF
C71 VDD dlycontrol2_in[4] 3.36fF
C72 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.bypass_in clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[16\] 1.24fF
C73 VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[26\] 0.96fF
C74 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.bypass_in dlycontrol3_in[2] 0.31fF
C75 dlycontrol4_in[2] edgedetect.dly_315ns_1.bypass_enable_w\[4\] 0.15fF
C76 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.bypass_in edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[0\] 0.20fF
C77 edgedetect.dly_315ns_1.bypass_enable_w\[3\] VDD 0.53fF
C78 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[1\] clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[8\] 0.23fF
C79 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.bypass_in VDD 2.36fF
C80 VDD clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit/a_1691_329# 0.10fF
C81 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit/mid VDD 0.34fF
C82 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[13\] clkgen.delay_155ns_3.enable_dlycontrol_w 0.12fF
C83 clkgen.delay_155ns_1.genblk1\[0\].dly_binary.in clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[8\] 1.44fF
C84 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[12\] VDD 0.96fF
C85 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit/mid clkgen.delay_155ns_2.enable_dlycontrol_w 0.14fF
C86 VDD dlycontrol2_in[3] 2.69fF
C87 VDD clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[6\] 0.95fF
C88 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.out clkgen.delay_155ns_3.genblk1\[4\].dly_binary.bypass_in 0.11fF
C89 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[31\].delay_unit/mid sample_p_in 0.12fF
C90 ena_in dlycontrol1_in[0] 0.13fF
C91 start_conv_in clkgen.delay_155ns_3.genblk1\[2\].dly_binary.signal_w\[4\] 0.21fF
C92 VDD clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[7\] 0.68fF
C93 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[16\] edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.signal_w\[0\] 0.10fF
C94 dlycontrol4_in[4] VDD 1.18fF
C95 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[29\].delay_unit/mid edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[18\].delay_unit/mid 0.12fF
C96 sample_n_in clk_dig_out 0.80fF
C97 clkgen.delay_155ns_2.genblk1\[0\].dly_binary.signal_w\[0\] clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[8\] 2.36fF
C98 dlycontrol3_in[4] edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.signal_w\[0\] 0.11fF
C99 edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.signal_w\[1\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.out 0.24fF
C100 VDD edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.genblk1\[0\].delay_unit/mid 0.29fF
C101 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.bypass_in clk_dig_out 0.62fF
C102 clkgen.delay_155ns_1.genblk1\[1\].dly_binary.bypass_in dlycontrol1_in[4] 0.21fF
C103 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[6\] clkgen.delay_155ns_1.genblk1\[2\].dly_binary.bypass_in 0.19fF
C104 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.bypass_in edgedetect.dly_315ns_1.bypass_enable_w\[4\] 0.21fF
C105 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.out clkgen.delay_155ns_3.genblk1\[1\].dly_binary.bypass_in 0.12fF
C106 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.bypass_in enable_dlycontrol_in 0.52fF
C107 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[0\] clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[7\] 0.42fF
C108 edgedetect.start_conv_edge_w clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[5\] 0.22fF
C109 clkgen.delay_155ns_2.genblk1\[1\].dly_binary.bypass_in clk_dig_out 1.30fF
C110 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit/a_1632_71# edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[6\] 0.13fF
C111 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.bypass_in edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.out 2.52fF
C112 dlycontrol1_in[2] dlycontrol1_in[4] 0.55fF
C113 clkgen.delay_155ns_3.genblk1\[1\].dly_binary.bypass_in clkgen.delay_155ns_3.bypass_enable_w\[0\] 1.24fF
C114 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[28\].delay_unit/mid VDD 0.40fF
C115 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.out clkgen.delay_155ns_3.genblk1\[2\].dly_binary.signal_w\[3\] 0.68fF
C116 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[0\] clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[16\] 0.83fF
C117 VDD clkgen.delay_155ns_1.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit/mid 0.24fF
C118 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit/mid edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[4\] 0.11fF
C119 edgedetect.dly_315ns_1.bypass_enable_w\[3\] edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.bypass_in 0.16fF
C120 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[4\] clkgen.delay_155ns_2.genblk1\[0\].dly_binary.signal_w\[0\] 0.12fF
C121 VDD clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit/mid 0.44fF
C122 edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.bypass_in VDD 6.52fF
C123 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.bypass_in clkgen.clk_comp_out 0.14fF
C124 sample_p_in edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.out 0.19fF
C125 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[2\] clkgen.delay_155ns_3.genblk1\[2\].dly_binary.bypass_in 0.29fF
C126 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.bypass_in clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[0\] 0.51fF
C127 edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.bypass_in edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[1\] 0.31fF
C128 nsample_p_in edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[14\] 0.24fF
C129 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.bypass_in clkgen.delay_155ns_2.genblk1\[1\].dly_binary.bypass_in 3.11fF
C130 VDD clkgen.delay_155ns_3.genblk1\[2\].dly_binary.bypass_in 3.44fF
C131 clkgen.delay_155ns_1.genblk1\[2\].dly_binary.bypass_in clkgen.delay_155ns_1.genblk1\[2\].dly_binary.out 1.42fF
C132 clkgen.delay_155ns_2.enable_dlycontrol_w clkgen.delay_155ns_2.bypass_enable_w\[2\] 0.96fF
C133 edgedetect.dly_315ns_1.bypass_enable_w\[2\] clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[6\] 0.23fF
C134 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[25\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[24\] 0.16fF
C135 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[22\].delay_unit/mid edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[23\] 0.12fF
C136 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.genblk1\[0\].delay_unit/mid VDD 0.37fF
C137 clkgen.delay_155ns_3.genblk1\[1\].dly_binary.signal_w\[0\] VDD 0.60fF
C138 clkgen.delay_155ns_2.genblk1\[0\].dly_binary.bypass_in clkgen.delay_155ns_1.genblk1\[1\].dly_binary.bypass_in 0.11fF
C139 ena_in sample_n_in 0.74fF
C140 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[27\].delay_unit/mid edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[24\] 0.14fF
C141 ndecision_finish_in clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit/mid 0.14fF
C142 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit/a_1632_71# clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[16\] 0.13fF
C143 dlycontrol4_in[4] edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.bypass_in 0.32fF
C144 clkgen.delay_155ns_1.genblk1\[0\].dly_binary.bypass_in dlycontrol1_in[4] 2.67fF
C145 dlycontrol2_in[1] dlycontrol2_in[2] 1.27fF
C146 ena_in clkgen.delay_155ns_1.genblk1\[3\].dly_binary.bypass_in 2.83fF
C147 VDD edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.signal_w\[1\] 1.56fF
C148 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.out clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[0\] 1.06fF
C149 dlycontrol4_in[4] edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[1\] 0.12fF
C150 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.genblk1\[1\].delay_unit/mid clkgen.delay_155ns_3.genblk1\[1\].dly_binary.bypass_in 0.11fF
C151 clkgen.delay_155ns_2.genblk1\[1\].dly_binary.genblk1\[0\].delay_unit/mid clkgen.delay_155ns_1.genblk1\[4\].dly_binary.out 0.14fF
C152 VDD clkgen.delay_155ns_3.genblk1\[2\].dly_binary.genblk1\[0\].delay_unit/mid 0.26fF
C153 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[22\].delay_unit/a_1691_329# VDD 0.13fF
C154 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.bypass_in edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.signal_w\[0\] 0.97fF
C155 ena_in clkgen.delay_155ns_2.genblk1\[1\].dly_binary.bypass_in 1.49fF
C156 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[8\].delay_unit/mid clkgen.delay_155ns_3.enable_dlycontrol_w 0.16fF
C157 edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[1\] edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[2\] 0.14fF
C158 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[11\].delay_unit/mid edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[29\] 0.14fF
C159 clkgen.delay_155ns_2.genblk1\[0\].dly_binary.signal_w\[0\] clkgen.delay_155ns_1.genblk1\[4\].dly_binary.bypass_in 0.34fF
C160 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[1\] clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[4\] 0.10fF
C161 sample_n_in clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[3\] 0.18fF
C162 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[7\] VDD 0.96fF
C163 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[0\] clkgen.delay_155ns_2.genblk1\[4\].dly_binary.bypass_in 2.35fF
C164 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[5\] clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[3\] 0.14fF
C165 clkgen.clk_dig_delayed_w clkgen.delay_155ns_1.genblk1\[1\].dly_binary.signal_w\[1\] 0.60fF
C166 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[16\].delay_unit/mid nsample_p_in 0.11fF
C167 VDD edgedetect.dly_315ns_1.bypass_enable_w\[4\] 1.88fF
C168 dlycontrol4_in[2] dlycontrol3_in[3] 2.29fF
C169 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit/mid VDD 0.46fF
C170 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[8\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[7\].delay_unit/mid 0.24fF
C171 VDD clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[2\] 0.41fF
C172 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[13\].delay_unit/mid edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[14\].delay_unit/mid 0.14fF
C173 dlycontrol1_in[4] clkgen.delay_155ns_3.enable_dlycontrol_w 0.11fF
C174 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit/mid clkgen.delay_155ns_1.genblk1\[0\].dly_binary.out 0.13fF
C175 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit/mid clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[16\] 0.11fF
C176 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.out VDD 1.93fF
C177 VDD edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[2\] 0.75fF
C178 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[16\] clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit/mid 0.11fF
C179 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[16\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[19\].delay_unit/mid 0.13fF
C180 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit/mid dlycontrol3_in[4] 0.11fF
C181 dlycontrol2_in[0] clkgen.delay_155ns_1.genblk1\[2\].dly_binary.genblk1\[0\].delay_unit/mid 0.18fF
C182 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[3\] VDD 0.81fF
C183 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[4\] ena_in 0.78fF
C184 nsample_p_1 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[15\] 0.17fF
C185 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[1\].delay_unit/mid edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.out 0.20fF
C186 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[10\].delay_unit/mid VDD 0.23fF
C187 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit/mid dlycontrol2_in[2] 0.29fF
C188 clkgen.delay_155ns_2.genblk1\[0\].dly_binary.bypass_in dlycontrol1_in[0] 0.17fF
C189 clkgen.delay_155ns_1.genblk1\[0\].dly_binary.out sample_n_out 0.38fF
C190 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[4\] VDD 0.60fF
C191 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.bypass_in dlycontrol3_in[3] 2.52fF
C192 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[8\] start_conv_in 0.25fF
C193 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.out clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[5\] 0.14fF
C194 clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[0\] dlycontrol1_in[4] 0.19fF
C195 clkgen.clk_dig_out clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[16\] 1.94fF
C196 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[0\] clkgen.delay_155ns_2.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit/mid 0.13fF
C197 dlycontrol4_in[4] edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[7\] 0.77fF
C198 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[20\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[19\].delay_unit/a_1632_71# 0.13fF
C199 clkgen.delay_155ns_1.genblk1\[0\].dly_binary.signal_w\[0\] clkgen.delay_155ns_3.genblk1\[4\].dly_binary.bypass_in 0.49fF
C200 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[16\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[16\].delay_unit/mid 0.13fF
C201 clkgen.delay_155ns_2.enable_dlycontrol_w clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[5\] 0.28fF
C202 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[1\] clkgen.delay_155ns_3.genblk1\[2\].dly_binary.bypass_in 0.71fF
C203 VDD clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[8\] 0.57fF
C204 VDD clkgen.delay_155ns_3.genblk1\[3\].dly_binary.bypass_in 2.00fF
C205 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.out clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[0\] 0.15fF
C206 clkgen.delay_155ns_3.genblk1\[0\].dly_binary.in VDD 3.42fF
C207 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[5\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[6\] 0.21fF
C208 clkgen.clk_dig_out VDD 6.19fF
C209 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.bypass_in dlycontrol1_in[4] 3.17fF
C210 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.out dlycontrol3_in[3] 0.14fF
C211 VDD clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit/mid 0.24fF
C212 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[12\].delay_unit/mid edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[13\] 0.10fF
C213 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[2\] VDD 0.73fF
C214 clkgen.delay_155ns_2.genblk1\[1\].dly_binary.bypass_in dlycontrol1_in[4] 0.10fF
C215 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.out edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.bypass_in 0.16fF
C216 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[5\] edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[0\] 0.36fF
C217 clkgen.delay_155ns_3.genblk1\[0\].dly_binary.in clkgen.delay_155ns_1.genblk1\[0\].dly_binary.genblk1\[0\].delay_unit/mid 0.17fF
C218 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[3\] enable_dlycontrol_in 0.13fF
C219 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[0\].delay_unit/mid edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.out 0.13fF
C220 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit/mid clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit/mid 0.14fF
C221 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[27\].delay_unit/a_1632_71# edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[28\] 0.13fF
C222 ndecision_finish_in VDD 5.57fF
C223 clkgen.clk_dig_out clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[0\] 0.38fF
C224 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit/mid clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[6\] 0.16fF
C225 VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[1\].delay_unit/mid 0.38fF
C226 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[16\] dlycontrol2_in[4] 2.69fF
C227 start_conv_in clkgen.delay_155ns_1.genblk1\[2\].dly_binary.out 0.16fF
C228 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[22\].delay_unit/mid edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[25\].delay_unit/mid 0.14fF
C229 clkgen.delay_155ns_3.genblk1\[0\].dly_binary.signal_w\[0\] dlycontrol3_in[1] 3.03fF
C230 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[4\].delay_unit/mid edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[4\] 0.16fF
C231 edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[4\] dlycontrol3_in[4] 0.12fF
C232 clkgen.delay_155ns_3.genblk1\[0\].dly_binary.signal_w\[0\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[6\].delay_unit/mid 0.13fF
C233 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[16\] edgedetect.dly_315ns_1.bypass_enable_w\[3\] 0.13fF
C234 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit/mid clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[8\] 0.11fF
C235 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.in edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[5\] 0.19fF
C236 clkgen.delay_155ns_2.bypass_enable_w\[1\] clkgen.delay_155ns_2.bypass_enable_w\[2\] 0.49fF
C237 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[8\] enable_dlycontrol_in 3.21fF
C238 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[6\] enable_dlycontrol_in 0.12fF
C239 clkgen.delay_155ns_1.genblk1\[2\].dly_binary.bypass_in enable_dlycontrol_in 2.08fF
C240 edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[4\] start_conv_in 0.18fF
C241 clkgen.clk_dig_delayed_w sample_n_1 0.17fF
C242 clkgen.delay_155ns_2.genblk1\[0\].dly_binary.signal_w\[0\] sample_n_4 0.28fF
C243 clkgen.delay_155ns_2.genblk1\[0\].dly_binary.bypass_in sample_n_in 0.16fF
C244 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[0\] dlycontrol4_in[0] 0.29fF
C245 VDD edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[2\] 0.47fF
C246 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[7\] VDD 0.73fF
C247 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit/mid edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[5\].delay_unit/mid 0.13fF
C248 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit/mid dlycontrol1_in[1] 0.14fF
C249 clkgen.delay_155ns_2.genblk1\[0\].dly_binary.bypass_in clkgen.delay_155ns_1.genblk1\[3\].dly_binary.bypass_in 1.91fF
C250 nsample_p_in start_conv_in 0.54fF
C251 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[8\] clkgen.delay_155ns_2.genblk1\[1\].dly_binary.signal_w\[0\] 0.33fF
C252 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[16\] dlycontrol2_in[3] 7.25fF
C253 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.bypass_in clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[8\] 0.16fF
C254 clkgen.delay_155ns_1.enable_dlycontrol_w dlycontrol3_in[4] 0.36fF
C255 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[0\].delay_unit/mid edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[1\] 0.12fF
C256 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[28\] sample_p_in 0.17fF
C257 VDD dlycontrol3_in[3] 2.83fF
C258 clkgen.delay_155ns_2.genblk1\[0\].dly_binary.bypass_in clkgen.delay_155ns_2.genblk1\[1\].dly_binary.bypass_in 0.23fF
C259 edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.signal_w\[1\] edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.signal_w\[2\] 0.14fF
C260 sample_p_in edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[32\] 3.54fF
C261 dlycontrol1_in[4] dlycontrol1_in[1] 0.34fF
C262 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit/mid VDD 0.37fF
C263 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[16\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[19\] 0.10fF
C264 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit/mid clkgen.clk_comp_out 0.15fF
C265 VDD clkgen.delay_155ns_1.genblk1\[3\].dly_binary.out_mux/a_505_21# 0.12fF
C266 VDD clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[14\] 0.72fF
C267 clkgen.delay_155ns_1.genblk1\[0\].dly_binary.signal_w\[0\] clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[0\] 0.41fF
C268 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit/mid dlycontrol2_in[3] 0.17fF
C269 dlycontrol2_in[4] dlycontrol3_in[0] 3.39fF
C270 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit/a_1691_329# VDD 0.11fF
C271 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[0\].delay_unit/mid VDD 0.42fF
C272 VDD clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[9\] 0.60fF
C273 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[13\] edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.bypass_in 0.14fF
C274 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.bypass_in edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit/mid 0.15fF
C275 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.out clkgen.delay_155ns_3.bypass_enable_w\[0\] 0.26fF
C276 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.out edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.bypass_in 0.40fF
C277 VDD clkgen.delay_155ns_2.enablebuffer/a_27_47# 0.27fF
C278 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[0\] edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[1\] 0.37fF
C279 VDD clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[8\] 1.33fF
C280 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.bypass_in clkgen.delay_155ns_1.bypass_enable_w\[1\] 0.26fF
C281 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.out edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.signal_w\[2\] 1.79fF
C282 dlycontrol3_in[0] dlycontrol2_in[3] 0.50fF
C283 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.bypass_in clkgen.delay_155ns_1.genblk1\[3\].dly_binary.out 0.18fF
C284 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[12\] ndecision_finish_in 0.28fF
C285 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[1\] clkgen.delay_155ns_3.genblk1\[0\].dly_binary.in 0.26fF
C286 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[7\] VDD 0.77fF
C287 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[16\] dlycontrol3_in[4] 0.80fF
C288 sample_p_in dlycontrol4_in[3] 0.32fF
C289 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[4\] sample_p_out 0.50fF
C290 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit/mid edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[5\] 0.12fF
C291 dlycontrol3_in[2] VDD 3.24fF
C292 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[16\] start_conv_in 0.69fF
C293 clkgen.delay_155ns_1.genblk1\[0\].dly_binary.in clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[0\] 0.23fF
C294 VDD clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit/mid 0.38fF
C295 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.bypass_in clkgen.delay_155ns_3.enable_dlycontrol_w 0.12fF
C296 edgedetect.dly_315ns_1.bypass_enable_w\[2\] edgedetect.dly_315ns_1.enable_dlycontrol_w 0.14fF
C297 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[4\] edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[0\].delay_unit/mid 0.11fF
C298 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit/mid edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[0\] 0.16fF
C299 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.bypass_in clkgen.delay_155ns_3.genblk1\[2\].dly_binary.signal_w\[1\] 0.23fF
C300 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[8\] edgedetect.dly_315ns_1.bypass_enable_w\[5\] 1.74fF
C301 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[4\] VDD 0.46fF
C302 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.bypass_in dlycontrol2_in[1] 1.40fF
C303 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[16\] clkgen.delay_155ns_3.genblk1\[2\].dly_binary.bypass_in 0.11fF
C304 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.signal_w\[0\] dlycontrol3_in[1] 0.18fF
C305 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[6\].delay_unit/mid edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.signal_w\[0\] 0.12fF
C306 clkgen.clk_dig_delayed_w clkgen.delay_155ns_1.genblk1\[0\].dly_binary.in 0.12fF
C307 clkgen.delay_155ns_2.bypass_enable_w\[4\] clkgen.delay_155ns_2.genblk1\[4\].dly_binary.bypass_in 0.11fF
C308 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[23\] dlycontrol4_in[4] 0.45fF
C309 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit/a_1632_71# clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[5\] 0.13fF
C310 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[12\] clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[16\] 1.06fF
C311 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.out clkgen.delay_155ns_3.genblk1\[3\].dly_binary.out 0.29fF
C312 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit/mid clkgen.delay_155ns_1.genblk1\[0\].dly_binary.out 0.10fF
C313 VDD clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[6\] 0.60fF
C314 dlycontrol2_in[0] clkgen.delay_155ns_1.genblk1\[4\].dly_binary.out 0.37fF
C315 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[13\] VDD 0.87fF
C316 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[32\] dlycontrol3_in[1] 1.99fF
C317 clkgen.delay_155ns_3.genblk1\[0\].dly_binary.bypass_in clkgen.delay_155ns_3.genblk1\[0\].dly_binary.signal_w\[1\] 0.34fF
C318 clkgen.delay_155ns_1.genblk1\[0\].dly_binary.bypass_in clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit/mid 0.11fF
C319 clkgen.delay_155ns_3.genblk1\[1\].dly_binary.bypass_in clkgen.delay_155ns_3.genblk1\[0\].dly_binary.bypass_in 0.50fF
C320 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.out dlycontrol2_in[1] 1.94fF
C321 VDD edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit/mid 0.29fF
C322 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[23\].delay_unit/mid VDD 0.42fF
C323 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.out clkgen.delay_155ns_2.genblk1\[3\].dly_binary.bypass_in 0.57fF
C324 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.in dlycontrol4_in[4] 0.21fF
C325 dlycontrol1_in[1] clkgen.delay_155ns_1.bypass_enable_w\[1\] 0.19fF
C326 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[0\] edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.out 3.11fF
C327 sample_n_2 VDD 0.70fF
C328 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[17\].delay_unit/mid edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[19\] 0.22fF
C329 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[16\] edgedetect.dly_315ns_1.bypass_enable_w\[4\] 1.33fF
C330 dlycontrol3_in[4] clkgen.delay_155ns_1.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit/mid 0.11fF
C331 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.out VDD 1.61fF
C332 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.bypass_in clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[0\] 1.77fF
C333 dlycontrol3_in[0] clkgen.delay_155ns_3.genblk1\[2\].dly_binary.bypass_in 2.26fF
C334 edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.bypass_in edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[0\] 0.24fF
C335 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.bypass_in VDD 1.19fF
C336 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[22\].delay_unit/mid edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.bypass_in 0.18fF
C337 VDD nsample_p_out 0.14fF
C338 edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.bypass_in edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.out 1.48fF
C339 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.bypass_in clkgen.delay_155ns_1.genblk1\[3\].dly_binary.bypass_in 0.80fF
C340 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.bypass_in clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[16\] 0.58fF
C341 start_conv_in enable_dlycontrol_in 1.13fF
C342 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[6\] VDD 0.79fF
C343 edgedetect.dly_315ns_1.enable_dlycontrol_w edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.bypass_in 0.35fF
C344 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit/mid VDD 0.24fF
C345 sample_n_2 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[0\] 0.21fF
C346 VDD clkgen.delay_155ns_3.genblk1\[2\].dly_binary.out_mux/a_505_21# 0.12fF
C347 edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.bypass_in clkgen.delay_155ns_3.enable_dlycontrol_w 0.88fF
C348 clkgen.delay_155ns_2.genblk1\[1\].dly_binary.out clkgen.delay_155ns_2.genblk1\[0\].dly_binary.signal_w\[0\] 0.11fF
C349 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.bypass_in dlycontrol3_in[4] 0.11fF
C350 edgedetect.dly_315ns_1.enable_dlycontrol_w edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.bypass_in 0.82fF
C351 dlycontrol3_in[0] clkgen.delay_155ns_3.genblk1\[2\].dly_binary.genblk1\[0\].delay_unit/mid 0.10fF
C352 clkgen.delay_155ns_1.genblk1\[1\].dly_binary.signal_w\[2\] dlycontrol1_in[4] 0.12fF
C353 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[16\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[17\].delay_unit/mid 0.13fF
C354 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.bypass_in start_conv_in 0.24fF
C355 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit/a_1632_71# clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[10\] 0.13fF
C356 clkgen.delay_155ns_2.genblk1\[1\].dly_binary.bypass_in dlycontrol2_in[3] 0.11fF
C357 VDD clkgen.delay_155ns_3.genblk1\[2\].dly_binary.signal_w\[4\] 1.03fF
C358 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.out edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[1\] 0.71fF
C359 clkgen.delay_155ns_1.genblk1\[0\].dly_binary.in clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[16\] 1.00fF
C360 clkgen.clk_dig_delayed_w clkgen.delay_155ns_1.genblk1\[1\].dly_binary.signal_w\[0\] 0.17fF
C361 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.bypass_in dlycontrol1_in[3] 0.48fF
C362 clkgen.clk_dig_out clkgen.delay_155ns_1.genblk1\[1\].dly_binary.bypass_in 0.32fF
C363 clkgen.delay_155ns_2.genblk1\[0\].dly_binary.bypass_in clkgen.delay_155ns_1.genblk1\[0\].dly_binary.out 1.07fF
C364 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[31\] VDD 0.99fF
C365 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[11\] VDD 0.82fF
C366 dlycontrol2_in[0] clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit/mid 0.10fF
C367 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[13\] clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit/mid 0.16fF
C368 clkgen.delay_155ns_3.genblk1\[2\].dly_binary.signal_w\[3\] clkgen.delay_155ns_3.bypass_enable_w\[0\] 0.93fF
C369 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[1\] sample_p_in 0.15fF
C370 VDD edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.signal_w\[0\] 1.78fF
C371 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.bypass_in edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[30\] 0.16fF
C372 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.out edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[11\] 0.22fF
C373 clkgen.delay_155ns_3.genblk1\[1\].dly_binary.out clkgen.delay_155ns_3.genblk1\[2\].dly_binary.signal_w\[0\] 0.15fF
C374 dlycontrol4_in[1] edgedetect.dly_315ns_1.enable_dlycontrol_w 0.12fF
C375 edgedetect.dly_315ns_1.bypass_enable_w\[1\] VDD 0.39fF
C376 dlycontrol4_in[1] nsample_p_1 0.21fF
C377 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[8\] dlycontrol4_in[2] 0.11fF
C378 ena_in clkgen.delay_155ns_2.genblk1\[0\].dly_binary.out 0.57fF
C379 dlycontrol2_in[0] dlycontrol1_in[4] 0.60fF
C380 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.out clkgen.delay_155ns_2.genblk1\[0\].dly_binary.out 0.47fF
C381 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[6\] VDD 0.72fF
C382 clkgen.delay_155ns_2.bypass_enable_w\[4\] edgedetect.dly_315ns_1.enable_dlycontrol_w 0.15fF
C383 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[0\] edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[0\] 1.59fF
C384 edgedetect.start_conv_edge_w clkgen.delay_155ns_3.genblk1\[0\].dly_binary.bypass_in 0.10fF
C385 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[16\] edgedetect.dly_315ns_1.bypass_enable_w\[5\] 0.17fF
C386 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[13\].delay_unit/mid edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.bypass_in 0.14fF
C387 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit/a_1691_329# VDD 0.16fF
C388 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.bypass_in enable_dlycontrol_in 0.61fF
C389 clkgen.delay_155ns_3.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit/a_1632_71# clkgen.delay_155ns_3.genblk1\[2\].dly_binary.signal_w\[3\] 0.13fF
C390 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit/mid clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[12\] 0.12fF
C391 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[20\].delay_unit/mid edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[21\] 0.16fF
C392 VDD clkgen.delay_155ns_1.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit/mid 0.32fF
C393 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.bypass_in clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit/mid 0.14fF
C394 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[2\] VDD 0.68fF
C395 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[1\] VDD 0.54fF
C396 clkgen.delay_155ns_1.genblk1\[0\].dly_binary.bypass_in clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[8\] 0.31fF
C397 start_conv_in clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[2\] 0.11fF
C398 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.bypass_in dlycontrol2_in[2] 5.29fF
C399 clkgen.delay_155ns_3.genblk1\[0\].dly_binary.in clkgen.delay_155ns_1.genblk1\[0\].dly_binary.bypass_in 0.13fF
C400 clkgen.delay_155ns_1.genblk1\[1\].dly_binary.out clkgen.delay_155ns_1.genblk1\[1\].dly_binary.signal_w\[0\] 0.98fF
C401 clkgen.delay_155ns_3.genblk1\[1\].dly_binary.bypass_in clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit/mid 0.12fF
C402 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.bypass_in dlycontrol1_in[4] 0.12fF
C403 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[20\] edgedetect.dly_315ns_1.bypass_enable_w\[5\] 0.22fF
C404 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[10\].delay_unit/mid VDD 0.51fF
C405 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[0\] clkgen.delay_155ns_2.genblk1\[4\].dly_binary.bypass_in 0.42fF
C406 dlycontrol2_in[0] clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[9\] 0.24fF
C407 VDD edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[11\] 0.51fF
C408 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[5\] edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.bypass_in 0.15fF
C409 edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[4\] dlycontrol4_in[2] 2.12fF
C410 clkgen.clk_dig_out dlycontrol1_in[0] 2.55fF
C411 dlycontrol2_in[0] clkgen.delay_155ns_2.genblk1\[0\].dly_binary.bypass_in 0.27fF
C412 sample_n_4 VDD 0.16fF
C413 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[7\] VDD 0.69fF
C414 edgedetect.dly_315ns_1.bypass_enable_w\[2\] dlycontrol2_in[4] 0.14fF
C415 clkgen.delay_155ns_1.genblk1\[0\].dly_binary.signal_w\[0\] clkgen.delay_155ns_2.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit/mid 0.13fF
C416 clkgen.clk_dig_out clkgen.delay_155ns_3.enable_dlycontrol_w 0.16fF
C417 clkgen.delay_155ns_2.genblk1\[0\].dly_binary.signal_w\[0\] enable_dlycontrol_in 0.38fF
C418 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[1\] clkgen.delay_155ns_3.genblk1\[2\].dly_binary.signal_w\[4\] 0.38fF
C419 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[1\] dlycontrol1_in[3] 0.35fF
C420 sample_p_2 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[3\] 0.69fF
C421 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.genblk1\[1\].delay_unit/mid clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[2\] 0.11fF
C422 nsample_n_2 VDD 0.32fF
C423 dlycontrol1_in[2] clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[8\] 0.11fF
C424 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[1\] VDD 0.48fF
C425 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit/mid VDD 0.36fF
C426 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[8\] dlycontrol2_in[2] 0.59fF
C427 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[12\] VDD 0.54fF
C428 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit/mid VDD 0.24fF
C429 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.bypass_in edgedetect.dly_315ns_1.bypass_enable_w\[5\] 0.36fF
C430 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[3\] VDD 0.74fF
C431 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.out clkgen.delay_155ns_1.genblk1\[2\].dly_binary.out 0.22fF
C432 clkgen.delay_155ns_1.genblk1\[1\].dly_binary.genblk1\[0\].delay_unit/mid VDD 0.48fF
C433 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit/mid VDD 0.35fF
C434 VDD clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[3\] 0.47fF
C435 VDD edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[14\] 0.67fF
C436 dlycontrol3_in[0] dlycontrol3_in[3] 0.16fF
C437 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.bypass_in clkgen.delay_155ns_1.genblk1\[0\].dly_binary.out 0.16fF
C438 clkgen.delay_155ns_3.genblk1\[1\].dly_binary.signal_w\[1\] clkgen.delay_155ns_3.genblk1\[1\].dly_binary.out 0.12fF
C439 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[2\] edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[3\] 0.12fF
C440 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[4\].delay_unit/a_1632_71# edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[5\] 0.14fF
C441 clkgen.delay_155ns_1.bypass_enable_w\[3\] clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[9\] 0.22fF
C442 clkgen.delay_155ns_2.genblk1\[1\].dly_binary.signal_w\[0\] clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[0\] 0.33fF
C443 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[10\].delay_unit/mid clkgen.clk_comp_out 0.16fF
C444 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.bypass_in edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[11\] 0.19fF
C445 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[7\] clkgen.delay_155ns_3.enable_dlycontrol_w 0.14fF
C446 clkgen.delay_155ns_2.genblk1\[0\].dly_binary.bypass_in clkgen.delay_155ns_1.bypass_enable_w\[3\] 0.12fF
C447 clkgen.delay_155ns_3.genblk1\[0\].dly_binary.in clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[0\] 0.91fF
C448 clkgen.clk_dig_out sample_n_in 0.31fF
C449 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[0\].delay_unit/mid clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[1\] 0.15fF
C450 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[0\] dlycontrol1_in[4] 0.41fF
C451 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[8\] VDD 2.99fF
C452 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[6\] VDD 0.64fF
C453 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.out edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[0\] 0.18fF
C454 VDD clkgen.delay_155ns_1.genblk1\[2\].dly_binary.bypass_in 2.23fF
C455 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[6\] clkgen.delay_155ns_1.genblk1\[1\].dly_binary.bypass_in 0.62fF
C456 clkgen.delay_155ns_3.genblk1\[0\].dly_binary.in clkgen.delay_155ns_1.genblk1\[3\].dly_binary.bypass_in 0.11fF
C457 dlycontrol4_in[2] dlycontrol3_in[4] 0.71fF
C458 clkgen.clk_dig_out clkgen.delay_155ns_1.genblk1\[3\].dly_binary.bypass_in 1.53fF
C459 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.bypass_in clkgen.delay_155ns_1.genblk1\[1\].dly_binary.signal_w\[2\] 0.83fF
C460 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[0\] edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.genblk1\[0\].delay_unit/mid 0.11fF
C461 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.bypass_in clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[0\].delay_unit/mid 0.18fF
C462 clkgen.clk_dig_out clkgen.delay_155ns_2.genblk1\[1\].dly_binary.bypass_in 1.49fF
C463 clkgen.delay_155ns_2.genblk1\[0\].dly_binary.bypass_in clkgen.delay_155ns_2.genblk1\[0\].dly_binary.out 0.67fF
C464 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit/mid clkgen.delay_155ns_3.enable_dlycontrol_w 0.11fF
C465 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[24\].delay_unit/mid VDD 0.39fF
C466 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[29\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[12\] 0.62fF
C467 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[16\].delay_unit/mid VDD 0.51fF
C468 dlycontrol1_in[0] clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[8\] 0.49fF
C469 dlycontrol3_in[1] clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[10\] 0.14fF
C470 VDD clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[13\] 0.72fF
C471 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[12\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.bypass_in 0.56fF
C472 VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[3\] 0.88fF
C473 VDD edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit/mid 0.29fF
C474 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit/mid clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit/mid 0.13fF
C475 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[30\].delay_unit/mid sample_p_in 0.12fF
C476 start_conv_in clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit/mid 0.16fF
C477 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[0\] dlycontrol4_in[5] 0.12fF
C478 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[0\] dlycontrol4_in[3] 4.45fF
C479 edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.out_mux/a_505_21# VDD 0.12fF
C480 clkgen.delay_155ns_3.genblk1\[1\].dly_binary.signal_w\[2\] dlycontrol2_in[4] 1.19fF
C481 clkgen.delay_155ns_2.bypass_enable_w\[3\] clkgen.delay_155ns_2.enable_dlycontrol_w 0.19fF
C482 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[4\] clkgen.delay_155ns_3.genblk1\[2\].dly_binary.bypass_in 0.16fF
C483 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.bypass_in edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[14\] 0.38fF
C484 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.out clkgen.delay_155ns_2.genblk1\[4\].dly_binary.bypass_in 0.15fF
C485 VDD clkgen.delay_155ns_1.genblk1\[2\].dly_binary.out 1.34fF
C486 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.bypass_in clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[16\] 0.15fF
C487 dlycontrol1_in[3] clkgen.delay_155ns_1.genblk1\[2\].dly_binary.bypass_in 0.54fF
C488 clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[1\] clkgen.delay_155ns_1.genblk1\[2\].dly_binary.bypass_in 0.71fF
C489 dlycontrol4_in[4] dlycontrol4_in[0] 6.62fF
C490 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[7\] clkgen.delay_155ns_1.genblk1\[3\].dly_binary.bypass_in 0.18fF
C491 VDD clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit/mid 0.27fF
C492 edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[4\] VDD 1.68fF
C493 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.bypass_in start_conv_in 0.23fF
C494 clkgen.delay_155ns_1.genblk1\[0\].dly_binary.in clkgen.delay_155ns_1.genblk1\[0\].dly_binary.signal_w\[0\] 1.08fF
C495 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[16\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.out 0.12fF
C496 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[7\] clkgen.delay_155ns_2.genblk1\[1\].dly_binary.bypass_in 0.21fF
C497 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.out edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.bypass_in 0.18fF
C498 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit/mid edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.out 0.16fF
C499 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[8\] clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[16\] 0.18fF
C500 VDD nsample_p_in 1.76fF
C501 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[28\].delay_unit/mid edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.bypass_in 0.12fF
C502 clkgen.delay_155ns_1.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit/mid clkgen.delay_155ns_1.genblk1\[1\].dly_binary.signal_w\[2\] 0.10fF
C503 VDD outbuf_2/a_27_47# 0.27fF
C504 dlycontrol3_in[4] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.out 1.09fF
C505 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[5\].delay_unit/mid VDD 0.36fF
C506 clkgen.delay_155ns_2.genblk1\[1\].dly_binary.out VDD 3.18fF
C507 clkgen.clk_dig_out dlycontrol1_in[1] 1.26fF
C508 clkgen.delay_155ns_1.enable_dlycontrol_w VDD 1.30fF
C509 edgedetect.start_conv_edge_w edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[6\] 0.11fF
C510 edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.bypass_in edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.bypass_in 0.13fF
C511 ndecision_finish_in edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[25\].delay_unit/mid 0.12fF
C512 edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.bypass_in edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.bypass_in 4.10fF
C513 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[10\].delay_unit/mid enable_dlycontrol_in 0.12fF
C514 dlycontrol4_in[1] dlycontrol4_in[4] 0.11fF
C515 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit/mid VDD 0.39fF
C516 sample_n_in clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[8\] 0.17fF
C517 VDD clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit/mid 0.40fF
C518 clkgen.delay_155ns_2.genblk1\[1\].dly_binary.signal_w\[0\] clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[16\] 0.57fF
C519 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[2\] clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[6\] 0.23fF
C520 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[23\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[23\].delay_unit/mid 0.14fF
C521 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.bypass_in clkgen.delay_155ns_3.genblk1\[4\].dly_binary.bypass_in 0.77fF
C522 VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[19\] 0.67fF
C523 clkgen.delay_155ns_1.enable_dlycontrol_w clkgen.delay_155ns_1.bypass_enable_w\[4\] 0.19fF
C524 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.bypass_in clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[8\] 0.30fF
C525 clkgen.delay_155ns_3.genblk1\[0\].dly_binary.bypass_in clkgen.delay_155ns_3.genblk1\[2\].dly_binary.out 0.20fF
C526 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.bypass_in dlycontrol1_in[0] 0.39fF
C527 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[12\] VDD 0.94fF
C528 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.out_mux/a_505_21# VDD 0.12fF
C529 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.bypass_in clkgen.delay_155ns_3.bypass_enable_w\[4\] 0.78fF
C530 clkgen.delay_155ns_3.genblk1\[1\].dly_binary.signal_w\[0\] edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.bypass_in 0.18fF
C531 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[23\].delay_unit/a_1691_329# VDD 0.16fF
C532 VDD clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit/mid 0.39fF
C533 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.out clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[8\] 2.44fF
C534 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.out clkgen.delay_155ns_3.enable_dlycontrol_w 1.18fF
C535 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.bypass_in enable_dlycontrol_in 0.32fF
C536 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit/mid edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit/mid 0.11fF
C537 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.bypass_in clkgen.delay_155ns_3.enable_dlycontrol_w 0.96fF
C538 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.out enable_dlycontrol_in 0.11fF
C539 dlycontrol3_in[0] clkgen.delay_155ns_3.genblk1\[2\].dly_binary.signal_w\[4\] 0.10fF
C540 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[14\] clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[16\] 0.11fF
C541 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[16\] dlycontrol3_in[4] 0.14fF
C542 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.out clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[1\] 0.21fF
C543 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[16\] VDD 6.30fF
C544 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit/mid VDD 0.35fF
C545 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.bypass_in clkgen.delay_155ns_2.genblk1\[3\].dly_binary.bypass_in 0.17fF
C546 ndecision_finish_in edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[26\].delay_unit/mid 0.11fF
C547 nsample_p_in edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.bypass_in 0.94fF
C548 dlycontrol3_in[4] VDD 5.54fF
C549 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[5\] VDD 0.63fF
C550 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.out clkgen.delay_155ns_2.genblk1\[1\].dly_binary.signal_w\[0\] 1.02fF
C551 VDD start_conv_in 6.19fF
C552 edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.signal_w\[0\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[6\] 0.12fF
C553 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.bypass_in edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.out 0.37fF
C554 dlycontrol4_in[2] edgedetect.dly_315ns_1.bypass_enable_w\[5\] 1.84fF
C555 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.out clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[0\] 0.18fF
C556 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.out dlycontrol4_in[0] 0.16fF
C557 VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[20\] 0.77fF
C558 sample_n_2 clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[0\] 0.75fF
C559 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.out clkgen.delay_155ns_2.genblk1\[3\].dly_binary.bypass_in 1.07fF
C560 clkgen.delay_155ns_3.genblk1\[2\].dly_binary.genblk1\[0\].delay_unit/mid clkgen.delay_155ns_3.genblk1\[2\].dly_binary.signal_w\[1\] 0.12fF
C561 clkgen.clk_dig_out clkgen.delay_155ns_1.genblk1\[0\].dly_binary.out 0.14fF
C562 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[30\] VDD 0.61fF
C563 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[0\] clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit/mid 0.10fF
C564 dlycontrol4_in[4] edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.out 1.65fF
C565 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.bypass_in sample_n_in 0.68fF
C566 clkgen.delay_155ns_3.genblk1\[1\].dly_binary.out VDD 0.79fF
C567 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit/mid start_conv_in 0.19fF
C568 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.out edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[10\] 0.20fF
C569 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[1\] edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[2\].delay_unit/mid 0.12fF
C570 VDD clkgen.delay_155ns_1.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit/mid 0.41fF
C571 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.out edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[8\] 4.69fF
C572 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit/a_1632_71# clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[2\] 0.13fF
C573 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[16\] edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.bypass_in 0.55fF
C574 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.bypass_in edgedetect.dly_315ns_1.bypass_enable_w\[5\] 0.29fF
C575 VDD enable_dlycontrol_in 6.13fF
C576 clkgen.delay_155ns_2.bypass_enable_w\[4\] edgedetect.dly_315ns_1.bypass_enable_w\[4\] 0.39fF
C577 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit/mid VDD 0.28fF
C578 clkgen.delay_155ns_3.genblk1\[0\].dly_binary.in clkgen.delay_155ns_1.genblk1\[1\].dly_binary.signal_w\[2\] 0.15fF
C579 edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[4\] edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[0\].delay_unit/mid 0.10fF
C580 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[1\] VDD 0.57fF
C581 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.out ndecision_finish_in 0.50fF
C582 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit/mid clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[8\] 0.18fF
C583 dlycontrol3_in[4] clkgen.clk_comp_out 2.39fF
C584 VDD nsample_n_out 0.37fF
C585 clkgen.delay_155ns_3.genblk1\[2\].dly_binary.signal_w\[0\] VDD 0.92fF
C586 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.bypass_in clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit/mid 0.16fF
C587 VDD clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit/mid 0.37fF
C588 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.bypass_in VDD 3.75fF
C589 edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.bypass_in edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.out 0.11fF
C590 clkgen.delay_155ns_2.enable_dlycontrol_w clk_dig_out 0.54fF
C591 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[0\] enable_dlycontrol_in 0.11fF
C592 clkgen.delay_155ns_1.genblk1\[1\].dly_binary.bypass_in clkgen.delay_155ns_1.genblk1\[2\].dly_binary.bypass_in 0.12fF
C593 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit/mid clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit/mid 0.16fF
C594 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[17\].delay_unit/mid VDD 0.31fF
C595 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[0\] VDD 0.68fF
C596 dlycontrol4_in[1] edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[4\] 0.11fF
C597 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[26\].delay_unit/a_1632_71# edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[27\] 0.13fF
C598 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[8\] clkgen.delay_155ns_3.genblk1\[2\].dly_binary.signal_w\[4\] 0.25fF
C599 ndecision_finish_in edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.bypass_in 0.64fF
C600 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[8\] dlycontrol2_in[2] 4.13fF
C601 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[4\] clkgen.delay_155ns_1.genblk1\[4\].dly_binary.bypass_in 0.11fF
C602 clkgen.delay_155ns_3.genblk1\[0\].dly_binary.in clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[1\] 0.15fF
C603 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[16\] clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[8\] 0.13fF
C604 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit/mid edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[4\] 0.20fF
C605 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[3\].delay_unit/mid edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[4\] 0.11fF
C606 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[10\].delay_unit/a_1691_329# VDD 0.13fF
C607 dlycontrol1_in[3] enable_dlycontrol_in 0.12fF
C608 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit/mid dlycontrol2_in[3] 0.15fF
C609 VDD edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[10\] 1.59fF
C610 sample_n_1 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit/mid 0.11fF
C611 dlycontrol2_in[0] clkgen.delay_155ns_3.genblk1\[0\].dly_binary.in 0.61fF
C612 dlycontrol2_in[0] clkgen.clk_dig_out 1.23fF
C613 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.bypass_in clkgen.delay_155ns_2.enable_dlycontrol_w 0.15fF
C614 VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[21\].delay_unit/mid 0.30fF
C615 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[5\] clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit/mid 0.15fF
C616 sample_p_3 sample_p_4 0.37fF
C617 dlycontrol4_in[4] edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[0\] 4.06fF
C618 edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.genblk1\[1\].delay_unit/mid edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[2\] 0.20fF
C619 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit/mid clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[4\] 0.26fF
C620 clkgen.delay_155ns_2.genblk1\[0\].dly_binary.signal_w\[0\] VDD 1.10fF
C621 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.bypass_in dlycontrol3_in[3] 0.13fF
C622 VDD outbuf_3/a_27_47# 0.18fF
C623 dlycontrol1_in[2] clkgen.delay_155ns_1.genblk1\[2\].dly_binary.out 2.34fF
C624 VDD edgedetect.dly_315ns_1.bypass_enable_w\[5\] 1.46fF
C625 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[1\] clkgen.delay_155ns_3.genblk1\[1\].dly_binary.out 0.63fF
C626 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.out clkgen.delay_155ns_2.enable_dlycontrol_w 0.40fF
C627 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[3\] clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[0\] 0.29fF
C628 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[16\] edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.signal_w\[2\] 0.58fF
C629 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[13\] VDD 0.87fF
C630 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[2\] clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[2\].delay_unit/mid 0.17fF
C631 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit/a_1691_329# VDD 0.10fF
C632 VDD clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[2\] 0.61fF
C633 dlycontrol2_in[2] clkgen.delay_155ns_2.bypass_enable_w\[2\] 0.20fF
C634 VDD edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit/mid 0.23fF
C635 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[2\].delay_unit/mid VDD 0.27fF
C636 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit/mid VDD 0.45fF
C637 clkgen.delay_155ns_1.genblk1\[0\].dly_binary.signal_w\[0\] clkgen.delay_155ns_2.genblk1\[1\].dly_binary.signal_w\[0\] 0.17fF
C638 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.bypass_in clkgen.delay_155ns_3.bypass_enable_w\[3\] 0.69fF
C639 clkgen.delay_155ns_2.bypass_enable_w\[3\] clkgen.delay_155ns_2.bypass_enable_w\[2\] 0.77fF
C640 VDD clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[0\].delay_unit/mid 0.22fF
C641 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.bypass_in dlycontrol4_in[2] 0.97fF
C642 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.out clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[4\] 0.19fF
C643 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[8\] clkgen.delay_155ns_3.enable_dlycontrol_w 0.17fF
C644 clkgen.delay_155ns_2.genblk1\[0\].dly_binary.signal_w\[0\] dlycontrol1_in[3] 0.34fF
C645 dlycontrol3_in[3] clkgen.delay_155ns_3.genblk1\[2\].dly_binary.signal_w\[1\] 0.14fF
C646 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[2\] clkgen.delay_155ns_1.genblk1\[2\].dly_binary.bypass_in 0.50fF
C647 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[4\] edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.out 0.26fF
C648 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.bypass_in edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[21\].delay_unit/mid 0.11fF
C649 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[7\] VDD 0.62fF
C650 clkgen.delay_155ns_3.genblk1\[1\].dly_binary.signal_w\[1\] VDD 0.66fF
C651 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[10\] start_conv_in 0.12fF
C652 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[11\] ndecision_finish_in 0.22fF
C653 clkgen.delay_155ns_1.bypass_enable_w\[2\] clkgen.delay_155ns_1.enable_dlycontrol_w 0.50fF
C654 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[4\] clkgen.delay_155ns_1.genblk1\[1\].dly_binary.signal_w\[2\] 0.71fF
C655 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[3\] clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[0\] 0.48fF
C656 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.bypass_in clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[10\].delay_unit/mid 0.10fF
C657 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[5\] clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[0\] 0.20fF
C658 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit/a_1632_71# edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[13\] 0.13fF
C659 clkgen.clk_dig_out clkgen.delay_155ns_2.genblk1\[0\].dly_binary.out 0.30fF
C660 clkgen.delay_155ns_3.genblk1\[0\].dly_binary.bypass_in clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[4\] 0.16fF
C661 sample_n_in clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[3\] 0.28fF
C662 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit/mid clkgen.delay_155ns_3.genblk1\[0\].dly_binary.bypass_in 0.15fF
C663 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[16\].delay_unit/a_1691_329# VDD 0.12fF
C664 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit/mid clkgen.delay_155ns_3.enable_dlycontrol_w 0.13fF
C665 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[1\] clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[0\].delay_unit/mid 0.11fF
C666 clkgen.delay_155ns_1.genblk1\[1\].dly_binary.genblk1\[0\].delay_unit/mid clkgen.delay_155ns_1.genblk1\[3\].dly_binary.bypass_in 0.12fF
C667 dlycontrol2_in[4] clkgen.delay_155ns_3.bypass_enable_w\[0\] 1.59fF
C668 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.bypass_in clkgen.delay_155ns_1.genblk1\[0\].dly_binary.out 3.91fF
C669 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit/mid VDD 0.20fF
C670 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.out edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.signal_w\[1\] 0.22fF
C671 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.bypass_in clkgen.delay_155ns_3.genblk1\[0\].dly_binary.bypass_in 1.73fF
C672 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit/mid clkgen.delay_155ns_2.genblk1\[1\].dly_binary.bypass_in 0.12fF
C673 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[5\] start_conv_in 0.15fF
C674 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[10\].delay_unit/mid edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[13\] 0.22fF
C675 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[13\] edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[14\] 0.11fF
C676 VDD edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[8\] 0.61fF
C677 clkgen.delay_155ns_2.genblk1\[1\].dly_binary.out clkgen.delay_155ns_1.genblk1\[0\].dly_binary.bypass_in 0.96fF
C678 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[3\] clkgen.delay_155ns_3.genblk1\[2\].dly_binary.bypass_in 0.15fF
C679 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[5\].delay_unit/mid edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[6\] 0.19fF
C680 clkgen.delay_155ns_1.genblk1\[1\].dly_binary.bypass_in start_conv_in 0.23fF
C681 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[16\] clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[16\] 0.16fF
C682 clkgen.enable_loop_in clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[4\] 0.25fF
C683 clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[0\] clkgen.delay_155ns_1.genblk1\[2\].dly_binary.bypass_in 0.45fF
C684 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.bypass_in clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit/mid 0.16fF
C685 sample_n_in clkgen.delay_155ns_1.genblk1\[2\].dly_binary.bypass_in 0.16fF
C686 clkgen.delay_155ns_2.enable_dlycontrol_w dlycontrol1_in[4] 1.01fF
C687 dlycontrol4_in[2] edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[1\] 0.96fF
C688 clkgen.delay_155ns_3.genblk1\[0\].dly_binary.in clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[0\] 0.71fF
C689 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[23\].delay_unit/mid edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.bypass_in 0.13fF
C690 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[4\] clkgen.delay_155ns_3.genblk1\[2\].dly_binary.signal_w\[4\] 0.11fF
C691 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[6\] clkgen.delay_155ns_1.genblk1\[3\].dly_binary.bypass_in 0.22fF
C692 edgedetect.dly_315ns_1.bypass_enable_w\[1\] edgedetect.dly_315ns_1.bypass_enable_w\[2\] 0.11fF
C693 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.out edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.bypass_in 1.25fF
C694 clkgen.delay_155ns_1.genblk1\[2\].dly_binary.bypass_in clkgen.delay_155ns_1.genblk1\[3\].dly_binary.bypass_in 0.40fF
C695 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.out edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.bypass_in 0.22fF
C696 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.in edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[4\] 0.23fF
C697 clkgen.delay_155ns_2.genblk1\[1\].dly_binary.bypass_in clkgen.delay_155ns_1.genblk1\[2\].dly_binary.bypass_in 0.34fF
C698 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.out clkgen.delay_155ns_3.genblk1\[0\].dly_binary.bypass_in 1.98fF
C699 edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.genblk1\[0\].delay_unit/mid edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.genblk1\[0\].delay_unit/mid 0.10fF
C700 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[2\].delay_unit/a_1632_71# clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[3\] 0.14fF
C701 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[16\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[14\].delay_unit/mid 0.13fF
C702 dlycontrol4_in[2] VDD 3.49fF
C703 edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.bypass_in edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[28\] 0.11fF
C704 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[5\].delay_unit/a_1691_329# VDD 0.11fF
C705 dlycontrol2_in[2] clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[11\] 0.23fF
C706 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.in edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[5\].delay_unit/mid 0.17fF
C707 dlycontrol4_in[4] dlycontrol4_in[5] 9.57fF
C708 dlycontrol4_in[4] dlycontrol4_in[3] 0.71fF
C709 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit/mid VDD 0.50fF
C710 clkgen.delay_155ns_3.genblk1\[0\].dly_binary.signal_w\[0\] clkgen.delay_155ns_3.genblk1\[3\].dly_binary.bypass_in 0.34fF
C711 clkgen.delay_155ns_2.bypass_enable_w\[3\] clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[5\] 0.29fF
C712 clkgen.delay_155ns_3.genblk1\[0\].dly_binary.in clkgen.delay_155ns_3.genblk1\[0\].dly_binary.signal_w\[0\] 0.16fF
C713 VDD clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit/mid 0.43fF
C714 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.out clkgen.delay_155ns_3.genblk1\[1\].dly_binary.signal_w\[2\] 0.34fF
C715 ndecision_finish_in clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit/mid 0.15fF
C716 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit/mid edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[6\] 0.10fF
C717 VDD clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[10\].delay_unit/mid 0.26fF
C718 VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[18\] 0.62fF
C719 clkgen.delay_155ns_1.genblk1\[1\].dly_binary.bypass_in enable_dlycontrol_in 0.16fF
C720 dlycontrol3_in[4] clkgen.delay_155ns_1.genblk1\[0\].dly_binary.bypass_in 1.68fF
C721 clkgen.delay_155ns_1.genblk1\[0\].dly_binary.bypass_in start_conv_in 0.59fF
C722 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[16\] edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[0\] 1.01fF
C723 edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.bypass_in clkgen.delay_155ns_3.bypass_enable_w\[0\] 0.23fF
C724 sample_p_in clkgen.delay_155ns_3.genblk1\[1\].dly_binary.genblk1\[0\].delay_unit/mid 0.11fF
C725 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[16\] edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.out 1.62fF
C726 clkgen.delay_155ns_2.genblk1\[0\].dly_binary.out clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[8\] 0.36fF
C727 clkgen.delay_155ns_2.genblk1\[1\].dly_binary.bypass_in clkgen.delay_155ns_1.genblk1\[2\].dly_binary.out 0.69fF
C728 dlycontrol4_in[1] nsample_p_out 0.30fF
C729 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.out clkgen.delay_155ns_2.bypass_enable_w\[1\] 0.31fF
C730 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[16\] clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[15\] 0.31fF
C731 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[16\] enable_dlycontrol_in 0.12fF
C732 clkgen.delay_155ns_3.genblk1\[1\].dly_binary.bypass_in clkgen.delay_155ns_3.genblk1\[0\].dly_binary.out 0.15fF
C733 dlycontrol3_in[4] edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.out 0.21fF
C734 edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[1\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.out 0.15fF
C735 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.out clkgen.clk_dig_delayed_w 0.26fF
C736 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.bypass_in VDD 6.70fF
C737 edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[0\] start_conv_in 0.17fF
C738 clkgen.delay_155ns_3.bypass_enable_w\[0\] clkgen.delay_155ns_3.genblk1\[2\].dly_binary.bypass_in 1.28fF
C739 edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.out start_conv_in 0.19fF
C740 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit/mid edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.out 0.14fF
C741 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.out VDD 0.61fF
C742 edgedetect.dly_315ns_1.bypass_enable_w\[1\] edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.bypass_in 0.34fF
C743 clkgen.delay_155ns_1.genblk1\[2\].dly_binary.bypass_in dlycontrol1_in[1] 0.12fF
C744 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.bypass_in edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[16\] 0.11fF
C745 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[0\] clkgen.delay_155ns_1.genblk1\[1\].dly_binary.bypass_in 0.10fF
C746 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[28\] edgedetect.dly_315ns_1.bypass_enable_w\[4\] 0.22fF
C747 clkgen.delay_155ns_3.genblk1\[1\].dly_binary.signal_w\[0\] clkgen.delay_155ns_3.bypass_enable_w\[0\] 0.94fF
C748 clkgen.delay_155ns_3.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit/mid start_conv_in 0.14fF
C749 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.in clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[16\] 0.43fF
C750 clkgen.delay_155ns_3.genblk1\[1\].dly_binary.out dlycontrol3_in[0] 0.15fF
C751 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit/mid clkgen.delay_155ns_3.genblk1\[1\].dly_binary.bypass_in 0.32fF
C752 start_conv_in clkgen.delay_155ns_3.enable_dlycontrol_w 0.12fF
C753 VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.out 3.92fF
C754 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.in dlycontrol3_in[4] 3.63fF
C755 clkgen.delay_155ns_2.bypass_enable_w\[0\] VDD 0.19fF
C756 clkgen.delay_155ns_3.genblk1\[0\].dly_binary.signal_w\[0\] dlycontrol3_in[3] 0.18fF
C757 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.bypass_in clkgen.delay_155ns_2.genblk1\[1\].dly_binary.signal_w\[0\] 1.28fF
C758 dlycontrol3_in[0] enable_dlycontrol_in 1.49fF
C759 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit/mid clkgen.delay_155ns_2.genblk1\[4\].dly_binary.bypass_in 0.11fF
C760 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.out edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.genblk1\[0\].delay_unit/mid 0.10fF
C761 VDD clkgen.delay_155ns_1.bypass_enable_w\[0\] 0.45fF
C762 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit/mid VDD 0.36fF
C763 clkgen.delay_155ns_2.genblk1\[0\].dly_binary.out clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[6\] 0.82fF
C764 VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[7\] 0.68fF
C765 dlycontrol1_in[1] clkgen.delay_155ns_1.genblk1\[2\].dly_binary.out 1.22fF
C766 dlycontrol1_in[0] enable_dlycontrol_in 0.79fF
C767 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[0\].delay_unit/a_1632_71# clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[1\] 0.13fF
C768 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit/mid edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[4\] 0.16fF
C769 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[4\] clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[0\] 0.47fF
C770 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit/mid clkgen.delay_155ns_3.bypass_enable_w\[3\] 0.11fF
C771 VDD edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[1\] 0.87fF
C772 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[25\].delay_unit/a_1632_71# edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[26\] 0.13fF
C773 VDD clkgen.delay_155ns_1.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit/a_1691_329# 0.12fF
C774 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.bypass_in edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.bypass_in 0.34fF
C775 clkgen.delay_155ns_1.genblk1\[1\].dly_binary.genblk1\[0\].delay_unit/mid clkgen.delay_155ns_1.genblk1\[0\].dly_binary.out 0.10fF
C776 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit/mid VDD 0.30fF
C777 dlycontrol3_in[4] clkgen.delay_155ns_1.genblk1\[3\].dly_binary.bypass_in 0.43fF
C778 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[2\] VDD 0.57fF
C779 VDD edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit/mid 0.24fF
C780 enable_dlycontrol_in clkgen.delay_155ns_3.enable_dlycontrol_w 1.75fF
C781 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[16\] clkgen.delay_155ns_2.genblk1\[1\].dly_binary.bypass_in 1.12fF
C782 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.out clkgen.delay_155ns_2.genblk1\[1\].dly_binary.signal_w\[0\] 0.25fF
C783 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[16\] VDD 6.50fF
C784 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[1\] edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.out 0.34fF
C785 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.bypass_in start_conv_in 0.89fF
C786 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[24\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[27\] 0.17fF
C787 edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit/a_1632_71# edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[3\] 0.14fF
C788 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[32\] clkgen.delay_155ns_3.genblk1\[3\].dly_binary.bypass_in 1.16fF
C789 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.bypass_in clkgen.delay_155ns_3.enable_dlycontrol_w 1.69fF
C790 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[16\] edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit/mid 0.10fF
C791 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.bypass_in edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.out 1.40fF
C792 clkgen.delay_155ns_2.genblk1\[1\].dly_binary.bypass_in start_conv_in 2.08fF
C793 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[10\].delay_unit/mid edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[13\].delay_unit/mid 0.11fF
C794 dlycontrol1_in[3] clkgen.delay_155ns_1.bypass_enable_w\[0\] 0.17fF
C795 VDD clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit/a_1691_329# 0.16fF
C796 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[16\] clkgen.delay_155ns_1.bypass_enable_w\[4\] 0.17fF
C797 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[4\] clkgen.delay_155ns_1.genblk1\[0\].dly_binary.signal_w\[1\] 0.48fF
C798 clkgen.delay_155ns_1.genblk1\[0\].dly_binary.genblk1\[0\].delay_unit/mid VDD 0.26fF
C799 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[4\] edgedetect.start_conv_edge_w 0.11fF
C800 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[0\] VDD 1.49fF
C801 clkgen.delay_155ns_1.bypass_enable_w\[4\] VDD 0.83fF
C802 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.out clkgen.delay_155ns_2.bypass_enable_w\[2\] 0.56fF
C803 VDD clkgen.delay_155ns_2.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit/mid 0.36fF
C804 clkgen.delay_155ns_3.genblk1\[0\].dly_binary.genblk1\[0\].delay_unit/mid VDD 0.40fF
C805 sample_n_in enable_dlycontrol_in 0.57fF
C806 clkgen.delay_155ns_2.genblk1\[0\].dly_binary.signal_w\[0\] dlycontrol1_in[0] 0.10fF
C807 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.signal_w\[0\] dlycontrol3_in[3] 1.41fF
C808 dlycontrol1_in[3] VDD 2.33fF
C809 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[13\] dlycontrol3_in[0] 0.11fF
C810 clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[1\] VDD 0.89fF
C811 clkgen.delay_155ns_2.bypass_enable_w\[4\] clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[7\] 0.14fF
C812 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[8\] dlycontrol1_in[4] 0.32fF
C813 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.bypass_in enable_dlycontrol_in 1.11fF
C814 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[0\].delay_unit/mid clkgen.delay_155ns_3.genblk1\[1\].dly_binary.bypass_in 0.15fF
C815 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[15\].delay_unit/mid VDD 0.47fF
C816 ndecision_finish_in clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit/mid 0.11fF
C817 clkgen.delay_155ns_1.genblk1\[0\].dly_binary.signal_w\[0\] clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[0\] 0.31fF
C818 clkgen.delay_155ns_2.genblk1\[1\].dly_binary.bypass_in enable_dlycontrol_in 0.57fF
C819 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[16\] clkgen.clk_comp_out 0.33fF
C820 edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[4\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[4\] 0.11fF
C821 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit/a_1632_71# clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[16\] 0.14fF
C822 clkgen.delay_155ns_1.bypass_enable_w\[4\] dlycontrol1_in[3] 0.83fF
C823 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit/a_1632_71# edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[5\] 0.14fF
C824 VDD edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.bypass_in 4.06fF
C825 dlycontrol2_in[3] clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[4\] 0.10fF
C826 edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.signal_w\[1\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[1\] 0.12fF
C827 VDD clkgen.clk_comp_out 4.67fF
C828 clkgen.delay_155ns_1.genblk1\[0\].dly_binary.signal_w\[0\] clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[3\] 0.66fF
C829 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[1\] VDD 0.64fF
C830 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[6\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[7\].delay_unit/mid 0.13fF
C831 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.bypass_in edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[8\] 0.18fF
C832 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[0\].delay_unit/mid edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.out 0.14fF
C833 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[12\] VDD 0.76fF
C834 VDD clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit/mid 0.55fF
C835 edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.bypass_in edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[0\] 1.23fF
C836 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.out edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[7\] 0.25fF
C837 clkgen.delay_155ns_3.bypass_enable_w\[0\] dlycontrol3_in[3] 1.30fF
C838 dlycontrol3_in[2] edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.signal_w\[0\] 0.12fF
C839 dlycontrol2_in[0] clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[6\] 0.13fF
C840 dlycontrol4_in[5] edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[2\] 0.11fF
C841 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.out edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.signal_w\[2\] 0.12fF
C842 clkgen.delay_155ns_2.genblk1\[1\].dly_binary.out clkgen.delay_155ns_1.genblk1\[0\].dly_binary.out 0.13fF
C843 dlycontrol2_in[0] clkgen.delay_155ns_1.genblk1\[2\].dly_binary.bypass_in 0.22fF
C844 edgedetect.ena_in clkgen.delay_155ns_2.genblk1\[0\].dly_binary.bypass_in 0.30fF
C845 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.bypass_in clkgen.delay_155ns_3.genblk1\[3\].dly_binary.bypass_in 0.32fF
C846 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[5\] VDD 0.61fF
C847 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[1\] VDD 0.72fF
C848 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[16\] dlycontrol4_in[2] 1.07fF
C849 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[28\] dlycontrol3_in[2] 0.38fF
C850 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.out clkgen.delay_155ns_2.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit/mid 0.12fF
C851 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[29\] nsample_p_in 0.15fF
C852 edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[4\] edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.bypass_in 1.51fF
C853 sample_p_1 VDD 0.25fF
C854 dlycontrol3_in[2] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[32\] 8.19fF
C855 nsample_p_in edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.bypass_in 0.38fF
C856 dlycontrol1_in[1] enable_dlycontrol_in 0.16fF
C857 VDD outbuf_4/a_27_47# 0.14fF
C858 clkgen.clk_dig_delayed_w clkgen.delay_155ns_2.genblk1\[1\].dly_binary.signal_w\[1\] 0.37fF
C859 dlycontrol2_in[4] clkgen.delay_155ns_3.genblk1\[0\].dly_binary.bypass_in 0.11fF
C860 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[0\] edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.signal_w\[0\] 0.17fF
C861 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[15\].delay_unit/mid edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.bypass_in 0.15fF
C862 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[9\] start_conv_in 0.14fF
C863 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[4\] clkgen.delay_155ns_1.genblk1\[1\].dly_binary.signal_w\[1\] 0.63fF
C864 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[2\] clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[0\] 0.18fF
C865 edgedetect.dly_315ns_1.bypass_enable_w\[2\] start_conv_in 0.28fF
C866 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[10\] VDD 0.77fF
C867 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[8\] edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit/mid 0.17fF
C868 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[4\] start_conv_in 0.12fF
C869 dlycontrol2_in[0] clkgen.delay_155ns_1.genblk1\[2\].dly_binary.out 3.22fF
C870 clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[4\] clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit/mid 0.12fF
C871 sample_p_in dlycontrol3_in[1] 0.21fF
C872 edgedetect.ena_in clkgen.delay_155ns_1.bypass_enable_w\[1\] 1.24fF
C873 VDD clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit/mid 0.48fF
C874 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[0\].delay_unit/mid VDD 0.43fF
C875 dlycontrol2_in[3] clkgen.delay_155ns_3.genblk1\[0\].dly_binary.bypass_in 0.11fF
C876 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[7\] clkgen.delay_155ns_2.enable_dlycontrol_w 0.31fF
C877 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.out edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.signal_w\[0\] 1.69fF
C878 clkgen.delay_155ns_2.genblk1\[1\].dly_binary.bypass_in clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[2\] 0.38fF
C879 ndecision_finish_in clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[12\] 0.57fF
C880 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.bypass_in edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[16\] 1.70fF
C881 VDD edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[7\] 0.49fF
C882 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.bypass_in clkgen.delay_155ns_3.genblk1\[1\].dly_binary.bypass_in 0.36fF
C883 VDD outbuf_1/a_27_47# 0.19fF
C884 VDD edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.signal_w\[2\] 0.69fF
C885 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit/mid dlycontrol3_in[0] 0.20fF
C886 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.bypass_in dlycontrol3_in[3] 0.12fF
C887 VDD clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit/mid 0.32fF
C888 dlycontrol4_in[2] edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.out 2.48fF
C889 clkgen.delay_155ns_2.genblk1\[0\].dly_binary.bypass_in clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[4\] 0.16fF
C890 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.out_mux/a_505_21# VDD 0.12fF
C891 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[0\].delay_unit/mid clk_dig_out 0.14fF
C892 clkgen.delay_155ns_1.enable_dlycontrol_w dlycontrol2_in[1] 0.22fF
C893 clkgen.enable_loop_in clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[16\] 0.29fF
C894 clkgen.delay_155ns_2.genblk1\[1\].dly_binary.out_mux/a_505_21# VDD 0.12fF
C895 clkgen.delay_155ns_2.genblk1\[0\].dly_binary.out clkgen.delay_155ns_1.genblk1\[2\].dly_binary.bypass_in 0.22fF
C896 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[3\].delay_unit/mid VDD 0.35fF
C897 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[10\] VDD 0.81fF
C898 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[16\] edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.bypass_in 2.09fF
C899 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[29\] start_conv_in 0.54fF
C900 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[15\] clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[14\] 0.27fF
C901 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.out clkgen.delay_155ns_3.genblk1\[1\].dly_binary.bypass_in 2.12fF
C902 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[16\] dlycontrol4_in[0] 0.26fF
C903 clkgen.delay_155ns_1.genblk1\[1\].dly_binary.signal_w\[2\] start_conv_in 0.10fF
C904 start_conv_in edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.bypass_in 1.41fF
C905 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.bypass_in dlycontrol3_in[0] 3.12fF
C906 dlycontrol3_in[4] dlycontrol4_in[0] 0.44fF
C907 clkgen.delay_155ns_2.bypass_enable_w\[0\] clkgen.delay_155ns_1.bypass_enable_w\[2\] 0.21fF
C908 start_conv_in edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.bypass_in 2.90fF
C909 clkgen.delay_155ns_2.genblk1\[1\].dly_binary.signal_w\[2\] VDD 0.36fF
C910 clkgen.delay_155ns_3.genblk1\[0\].dly_binary.in clkgen.delay_155ns_1.genblk1\[0\].dly_binary.in 0.11fF
C911 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[11\] clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[7\] 0.10fF
C912 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[5\] VDD 0.90fF
C913 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.out_mux/a_505_21# VDD 0.14fF
C914 clkgen.delay_155ns_3.genblk1\[0\].dly_binary.bypass_in clkgen.delay_155ns_3.genblk1\[2\].dly_binary.bypass_in 0.62fF
C915 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.out dlycontrol1_in[0] 0.16fF
C916 VDD clkgen.delay_155ns_1.genblk1\[1\].dly_binary.bypass_in 3.56fF
C917 nsample_p_out dlycontrol4_in[3] 0.35fF
C918 edgedetect.start_conv_edge_w clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[4\] 0.12fF
C919 clkgen.delay_155ns_1.genblk1\[0\].dly_binary.in ndecision_finish_in 0.71fF
C920 dlycontrol2_in[0] dlycontrol3_in[4] 0.68fF
C921 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.bypass_in clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[8\] 0.99fF
C922 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.bypass_in clkgen.delay_155ns_3.enable_dlycontrol_w 0.93fF
C923 clkgen.delay_155ns_3.genblk1\[1\].dly_binary.out edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.bypass_in 0.22fF
C924 dlycontrol1_in[2] VDD 2.63fF
C925 dlycontrol4_in[1] dlycontrol3_in[4] 0.21fF
C926 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[17\].delay_unit/a_1632_71# edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[18\] 0.14fF
C927 clkgen.delay_155ns_1.enable_dlycontrol_w clkgen.delay_155ns_1.bypass_enable_w\[3\] 1.02fF
C928 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[16\] VDD 3.99fF
C929 clkgen.delay_155ns_3.bypass_enable_w\[0\] clkgen.delay_155ns_3.genblk1\[2\].dly_binary.signal_w\[4\] 1.96fF
C930 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[0\].delay_unit/mid edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[1\] 0.10fF
C931 edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[4\] edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.out 0.17fF
C932 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[0\] clkgen.delay_155ns_1.genblk1\[0\].dly_binary.out 3.32fF
C933 sample_p_2 sample_p_3 0.31fF
C934 clkgen.delay_155ns_1.bypass_enable_w\[2\] VDD 0.29fF
C935 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit/mid VDD 0.37fF
C936 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.bypass_in edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[29\] 0.13fF
C937 dlycontrol1_in[0] clkgen.delay_155ns_1.bypass_enable_w\[0\] 0.19fF
C938 VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[14\].delay_unit/mid 0.27fF
C939 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.in edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.out 0.31fF
C940 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.bypass_in edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.bypass_in 5.15fF
C941 dlycontrol1_in[3] clkgen.delay_155ns_1.genblk1\[1\].dly_binary.bypass_in 2.83fF
C942 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.bypass_in edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.bypass_in 0.82fF
C943 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit/mid clkgen.delay_155ns_2.genblk1\[4\].dly_binary.bypass_in 0.12fF
C944 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[7\] clkgen.delay_155ns_2.enable_dlycontrol_w 0.45fF
C945 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit/mid dlycontrol2_in[4] 0.14fF
C946 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[31\].delay_unit/mid start_conv_in 0.14fF
C947 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.out edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[10\] 0.49fF
C948 dlycontrol1_in[2] dlycontrol1_in[3] 0.64fF
C949 edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[1\] edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.out 0.75fF
C950 VDD dlycontrol3_in[0] 4.79fF
C951 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[11\] clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[16\] 0.49fF
C952 VDD clkgen.delay_155ns_1.genblk1\[0\].dly_binary.bypass_in 1.82fF
C953 clkgen.delay_155ns_3.genblk1\[0\].dly_binary.in clkgen.delay_155ns_1.genblk1\[1\].dly_binary.signal_w\[0\] 0.44fF
C954 VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[6\] 1.23fF
C955 clkgen.delay_155ns_2.genblk1\[0\].dly_binary.signal_w\[0\] clkgen.delay_155ns_1.genblk1\[0\].dly_binary.out 0.38fF
C956 edgedetect.start_conv_edge_w edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[7\].delay_unit/mid 0.11fF
C957 dlycontrol2_in[0] enable_dlycontrol_in 0.20fF
C958 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[12\] clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit/a_1632_71# 0.13fF
C959 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[6\] clkgen.delay_155ns_2.genblk1\[3\].dly_binary.bypass_in 0.14fF
C960 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.in edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[7\] 0.50fF
C961 dlycontrol1_in[0] VDD 3.50fF
C962 nsample_n_3 VDD 0.38fF
C963 clkgen.delay_155ns_2.genblk1\[1\].dly_binary.out clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[0\] 0.46fF
C964 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[7\] clkgen.delay_155ns_2.bypass_enable_w\[1\] 0.19fF
C965 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[8\] edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit/a_1632_71# 0.13fF
C966 VDD edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[0\] 1.10fF
C967 VDD edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.out 1.71fF
C968 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[23\] VDD 1.17fF
C969 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[15\] VDD 0.57fF
C970 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.bypass_in clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit/mid 0.16fF
C971 edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.bypass_in edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[21\].delay_unit/mid 0.10fF
C972 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.out clkgen.delay_155ns_2.genblk1\[1\].dly_binary.bypass_in 0.92fF
C973 dlycontrol2_in[3] clkgen.delay_155ns_2.bypass_enable_w\[2\] 0.12fF
C974 clkgen.delay_155ns_3.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit/mid VDD 0.24fF
C975 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[16\] edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.out 0.76fF
C976 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[2\] VDD 0.54fF
C977 VDD clkgen.delay_155ns_3.enable_dlycontrol_w 2.36fF
C978 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit/mid clkgen.delay_155ns_1.genblk1\[2\].dly_binary.bypass_in 0.12fF
C979 dlycontrol1_in[0] clkgen.delay_155ns_1.bypass_enable_w\[4\] 0.16fF
C980 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[8\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.out 0.49fF
C981 clkgen.delay_155ns_3.genblk1\[0\].dly_binary.bypass_in clkgen.delay_155ns_3.genblk1\[3\].dly_binary.bypass_in 0.25fF
C982 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit/mid clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[0\] 0.14fF
C983 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.in VDD 3.02fF
C984 sample_p_in edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit/mid 0.12fF
C985 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.bypass_in clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[16\] 0.13fF
C986 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[3\].delay_unit/mid edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[7\] 0.13fF
C987 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit/mid clkgen.delay_155ns_1.genblk1\[3\].dly_binary.bypass_in 0.13fF
C988 nsample_n_in enable_dlycontrol_in 0.36fF
C989 dlycontrol1_in[0] dlycontrol1_in[3] 2.07fF
C990 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[0\].delay_unit/mid clkgen.delay_155ns_2.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit/mid 0.12fF
C991 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[15\] clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit/a_1632_71# 0.14fF
C992 VDD edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[15\] 0.51fF
C993 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.genblk1\[0\].delay_unit/mid clkgen.delay_155ns_2.genblk1\[1\].dly_binary.signal_w\[0\] 0.33fF
C994 edgedetect.start_conv_edge_w edgedetect.dly_315ns_1.enable_dlycontrol_w 0.18fF
C995 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[7\] edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[8\] 0.26fF
C996 sample_n_3 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit/mid 0.11fF
C997 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[0\] start_conv_in 0.13fF
C998 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit/mid enable_dlycontrol_in 0.14fF
C999 clkgen.clk_dig_out clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit/mid 0.11fF
C1000 clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[0\] VDD 1.49fF
C1001 sample_n_in VDD 4.98fF
C1002 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.out clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[16\] 1.58fF
C1003 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit/mid clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[4\] 0.32fF
C1004 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[8\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[32\] 1.85fF
C1005 VDD clkgen.delay_155ns_1.genblk1\[3\].dly_binary.bypass_in 4.43fF
C1006 clkgen.delay_155ns_2.genblk1\[1\].dly_binary.genblk1\[0\].delay_unit/mid VDD 0.36fF
C1007 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.out edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[0\] 0.24fF
C1008 VDD clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[0\].delay_unit/mid 0.41fF
C1009 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[13\] VDD 0.81fF
C1010 clkgen.delay_155ns_2.genblk1\[1\].dly_binary.bypass_in VDD 6.80fF
C1011 VDD edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[8\] 2.04fF
C1012 sample_n_in clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[0\] 0.20fF
C1013 VDD clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit/mid 0.51fF
C1014 edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.signal_w\[0\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[1\] 0.21fF
C1015 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[1\] sample_n_1 0.15fF
C1016 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[10\].delay_unit/a_1632_71# clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[11\] 0.13fF
C1017 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[0\] clkgen.delay_155ns_1.genblk1\[3\].dly_binary.bypass_in 0.33fF
C1018 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.in edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.bypass_in 1.53fF
C1019 clkgen.delay_155ns_1.bypass_enable_w\[4\] clkgen.delay_155ns_1.genblk1\[3\].dly_binary.bypass_in 0.15fF
C1020 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit/a_1632_71# clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[6\] 0.14fF
C1021 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit/mid VDD 0.53fF
C1022 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[0\] clkgen.delay_155ns_2.genblk1\[1\].dly_binary.bypass_in 0.25fF
C1023 clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[1\] clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[0\] 0.12fF
C1024 sample_n_in dlycontrol1_in[3] 0.54fF
C1025 nsample_p_in edgedetect.dly_315ns_1.bypass_enable_w\[0\] 0.15fF
C1026 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[0\].delay_unit/mid clkgen.delay_155ns_3.genblk1\[1\].dly_binary.bypass_in 0.20fF
C1027 inbuf_2/a_27_47# VDD 0.10fF
C1028 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[7\] clkgen.delay_155ns_2.bypass_enable_w\[2\] 0.10fF
C1029 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit/a_1632_71# clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[7\] 0.13fF
C1030 dlycontrol1_in[3] clkgen.delay_155ns_1.genblk1\[3\].dly_binary.bypass_in 0.54fF
C1031 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[4\] VDD 0.49fF
C1032 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[0\] VDD 1.17fF
C1033 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[28\] nsample_p_in 0.28fF
C1034 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[16\] dlycontrol1_in[1] 0.29fF
C1035 clkgen.delay_155ns_1.genblk1\[1\].dly_binary.out dlycontrol1_in[4] 0.12fF
C1036 VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[25\].delay_unit/mid 0.28fF
C1037 sample_n_in clkgen.clk_comp_out 0.24fF
C1038 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit/mid edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[10\] 0.10fF
C1039 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[0\] edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.signal_w\[0\] 3.33fF
C1040 ndecision_finish_in clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[8\] 0.96fF
C1041 VDD dlycontrol1_in[1] 4.00fF
C1042 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.bypass_in clkgen.delay_155ns_2.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit/mid 0.13fF
C1043 clkgen.delay_155ns_3.genblk1\[1\].dly_binary.bypass_in dlycontrol2_in[4] 0.24fF
C1044 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[9\].delay_unit/mid dlycontrol3_in[1] 0.21fF
C1045 clkgen.delay_155ns_3.genblk1\[0\].dly_binary.in clkgen.delay_155ns_2.genblk1\[1\].dly_binary.signal_w\[0\] 0.25fF
C1046 dlycontrol4_in[2] edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.bypass_in 0.13fF
C1047 dlycontrol1_in[4] clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[16\] 2.76fF
C1048 dlycontrol1_in[2] clkgen.delay_155ns_1.genblk1\[1\].dly_binary.bypass_in 0.28fF
C1049 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.bypass_in edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[8\] 0.68fF
C1050 clkgen.delay_155ns_2.genblk1\[1\].dly_binary.bypass_in clkgen.clk_comp_out 0.95fF
C1051 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[8\] clkgen.delay_155ns_3.genblk1\[3\].dly_binary.out 0.30fF
C1052 edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.out edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.signal_w\[2\] 1.06fF
C1053 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[1\] VDD 0.58fF
C1054 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[4\] dlycontrol1_in[3] 0.43fF
C1055 ndecision_finish_in clkgen.delay_155ns_2.genblk1\[1\].dly_binary.signal_w\[0\] 0.74fF
C1056 clkgen.delay_155ns_3.genblk1\[1\].dly_binary.bypass_in dlycontrol2_in[3] 3.92fF
C1057 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.bypass_in dlycontrol3_in[1] 0.20fF
C1058 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.bypass_in edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.out 3.87fF
C1059 clkgen.delay_155ns_3.enable_dlycontrol_w clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit/mid 0.12fF
C1060 VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[26\].delay_unit/mid 0.28fF
C1061 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.signal_w\[1\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.out 0.46fF
C1062 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit/mid clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[8\] 0.16fF
C1063 dlycontrol4_in[1] dlycontrol4_in[2] 0.71fF
C1064 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[16\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[28\] 0.18fF
C1065 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.bypass_in edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.bypass_in 0.16fF
C1066 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.out edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.out 5.02fF
C1067 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.bypass_in dlycontrol2_in[2] 1.23fF
C1068 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.out dlycontrol1_in[4] 0.77fF
C1069 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[12\].delay_unit/mid VDD 0.33fF
C1070 clkgen.delay_155ns_1.genblk1\[1\].dly_binary.bypass_in clkgen.delay_155ns_1.genblk1\[0\].dly_binary.bypass_in 0.49fF
C1071 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[9\] VDD 0.61fF
C1072 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[28\] start_conv_in 0.10fF
C1073 edgedetect.dly_315ns_1.bypass_enable_w\[2\] VDD 0.54fF
C1074 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[0\] edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[10\] 0.14fF
C1075 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.out edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.bypass_in 0.20fF
C1076 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[1\].delay_unit/a_1632_71# edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[2\] 0.14fF
C1077 start_conv_in edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[32\] 0.15fF
C1078 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.bypass_in edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[1\] 0.16fF
C1079 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[4\] VDD 0.68fF
C1080 dlycontrol1_in[0] clkgen.delay_155ns_1.genblk1\[1\].dly_binary.bypass_in 2.60fF
C1081 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[16\] dlycontrol3_in[0] 6.20fF
C1082 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[16\] edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.genblk1\[0\].delay_unit/mid 0.12fF
C1083 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.out dlycontrol3_in[4] 0.49fF
C1084 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.out edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[7\] 0.13fF
C1085 dlycontrol3_in[4] edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.genblk1\[0\].delay_unit/mid 0.16fF
C1086 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[0\] clkgen.delay_155ns_3.genblk1\[2\].dly_binary.out 0.43fF
C1087 dlycontrol4_in[5] edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[2\].delay_unit/mid 0.12fF
C1088 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[1\] clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[0\] 0.29fF
C1089 dlycontrol1_in[2] dlycontrol1_in[0] 0.81fF
C1090 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[4\] VDD 1.05fF
C1091 clkgen.delay_155ns_1.bypass_enable_w\[2\] clkgen.delay_155ns_1.genblk1\[0\].dly_binary.bypass_in 0.44fF
C1092 clkgen.delay_155ns_1.genblk1\[1\].dly_binary.bypass_in clkgen.delay_155ns_3.enable_dlycontrol_w 1.32fF
C1093 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[2\] clkgen.delay_155ns_1.genblk1\[1\].dly_binary.bypass_in 0.12fF
C1094 sample_p_4 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[3\] 0.12fF
C1095 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[28\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[30\] 0.24fF
C1096 sample_p_2 edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.bypass_in 1.31fF
C1097 clkgen.delay_155ns_3.bypass_enable_w\[0\] start_conv_in 0.12fF
C1098 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.in edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[5\] 0.17fF
C1099 VDD clkgen.delay_155ns_1.genblk1\[0\].dly_binary.out 0.98fF
C1100 clkgen.delay_155ns_3.genblk1\[1\].dly_binary.bypass_in clkgen.delay_155ns_3.genblk1\[2\].dly_binary.bypass_in 0.69fF
C1101 edgedetect.start_conv_edge_w clkgen.delay_155ns_2.genblk1\[2\].dly_binary.bypass_in 0.13fF
C1102 clkgen.delay_155ns_3.genblk1\[1\].dly_binary.signal_w\[0\] clkgen.delay_155ns_3.genblk1\[0\].dly_binary.signal_w\[1\] 0.16fF
C1103 clkgen.delay_155ns_2.genblk1\[1\].dly_binary.out clkgen.delay_155ns_2.genblk1\[3\].dly_binary.bypass_in 0.34fF
C1104 dlycontrol3_in[4] dlycontrol4_in[3] 0.32fF
C1105 VDD edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.signal_w\[1\] 0.39fF
C1106 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.bypass_in clkgen.delay_155ns_2.bypass_enable_w\[4\] 0.28fF
C1107 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.bypass_in clkgen.clk_dig_delayed_w 0.21fF
C1108 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.bypass_in edgedetect.dly_315ns_1.bypass_enable_w\[0\] 0.10fF
C1109 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.out VDD 5.28fF
C1110 dlycontrol4_in[1] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.out 3.67fF
C1111 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.bypass_in edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.signal_w\[0\] 0.21fF
C1112 VDD clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[2\].delay_unit/mid 0.19fF
C1113 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.out clkgen.delay_155ns_3.genblk1\[1\].dly_binary.out 0.21fF
C1114 edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[4\] sample_p_4 1.10fF
C1115 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[29\] VDD 1.03fF
C1116 VDD clkgen.delay_155ns_1.genblk1\[1\].dly_binary.signal_w\[2\] 0.89fF
C1117 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit/a_1691_329# VDD 0.13fF
C1118 VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.bypass_in 4.52fF
C1119 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.bypass_in edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[28\] 0.19fF
C1120 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit/mid clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[13\] 0.21fF
C1121 VDD edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.bypass_in 5.94fF
C1122 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[10\].delay_unit/mid clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit/mid 0.11fF
C1123 VDD clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[5\] 0.58fF
C1124 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.bypass_in edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[32\] 0.18fF
C1125 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[24\].delay_unit/mid edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[25\] 0.30fF
C1126 dlycontrol1_in[3] clkgen.delay_155ns_1.genblk1\[0\].dly_binary.out 0.14fF
C1127 VDD dlycontrol4_in[0] 1.88fF
C1128 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[29\].delay_unit/mid start_conv_in 0.11fF
C1129 clkgen.delay_155ns_3.genblk1\[2\].dly_binary.signal_w\[2\] clkgen.delay_155ns_3.genblk1\[2\].dly_binary.out 0.25fF
C1130 clkgen.delay_155ns_3.genblk1\[1\].dly_binary.out_mux/a_505_21# VDD 0.11fF
C1131 clkgen.delay_155ns_2.enable_dlycontrol_w clkgen.delay_155ns_1.genblk1\[2\].dly_binary.bypass_in 0.22fF
C1132 clkgen.delay_155ns_1.genblk1\[1\].dly_binary.bypass_in clkgen.delay_155ns_1.genblk1\[3\].dly_binary.bypass_in 0.84fF
C1133 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit/mid edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.out 0.16fF
C1134 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.out edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.bypass_in 0.44fF
C1135 edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[0\] edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.out 0.28fF
C1136 dlycontrol1_in[2] sample_n_in 0.80fF
C1137 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit/a_1632_71# clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[7\] 0.13fF
C1138 clkgen.delay_155ns_2.genblk1\[1\].dly_binary.bypass_in clkgen.delay_155ns_1.genblk1\[1\].dly_binary.bypass_in 0.13fF
C1139 dlycontrol2_in[0] clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[16\] 2.80fF
C1140 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[1\] VDD 1.64fF
C1141 dlycontrol1_in[2] clkgen.delay_155ns_1.genblk1\[3\].dly_binary.bypass_in 0.26fF
C1142 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit/mid dlycontrol4_in[1] 0.11fF
C1143 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[5\] clkgen.delay_155ns_2.genblk1\[3\].dly_binary.bypass_in 0.12fF
C1144 clkgen.delay_155ns_3.genblk1\[1\].dly_binary.signal_w\[2\] VDD 1.21fF
C1145 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.in edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[6\] 0.61fF
C1146 dlycontrol2_in[0] VDD 2.93fF
C1147 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[30\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[29\].delay_unit/mid 0.14fF
C1148 clkgen.delay_155ns_3.genblk1\[2\].dly_binary.genblk1\[1\].delay_unit/mid dlycontrol3_in[3] 0.12fF
C1149 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.bypass_in clkgen.delay_155ns_1.genblk1\[1\].dly_binary.out 4.51fF
C1150 dlycontrol1_in[2] clkgen.delay_155ns_2.genblk1\[1\].dly_binary.bypass_in 0.38fF
C1151 VDD clkgen.delay_155ns_3.genblk1\[2\].dly_binary.signal_w\[1\] 0.49fF
C1152 dlycontrol4_in[1] VDD 6.14fF
C1153 clkgen.delay_155ns_1.genblk1\[2\].dly_binary.genblk1\[1\].delay_unit/a_1632_71# clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[2\] 0.13fF
C1154 dlycontrol2_in[1] VDD 2.47fF
C1155 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.out edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.bypass_in 1.58fF
C1156 sample_n_1 start_conv_in 0.36fF
C1157 VDD edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit/mid 0.24fF
C1158 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.out clkgen.delay_155ns_2.genblk1\[0\].dly_binary.out 3.80fF
C1159 clkgen.delay_155ns_3.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit/a_1691_329# VDD 0.10fF
C1160 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit/mid VDD 0.29fF
C1161 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[8\] VDD 0.67fF
C1162 clkgen.delay_155ns_2.enable_dlycontrol_w clkgen.delay_155ns_1.genblk1\[2\].dly_binary.out 0.51fF
C1163 clkgen.delay_155ns_2.bypass_enable_w\[4\] VDD 0.75fF
C1164 clkgen.delay_155ns_3.bypass_enable_w\[1\] VDD 0.22fF
C1165 dlycontrol2_in[0] clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[0\] 0.17fF
C1166 clkgen.delay_155ns_2.genblk1\[0\].dly_binary.signal_w\[0\] clkgen.delay_155ns_1.genblk1\[1\].dly_binary.signal_w\[1\] 0.27fF
C1167 dlycontrol2_in[0] clkgen.delay_155ns_1.bypass_enable_w\[4\] 0.10fF
C1168 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[28\] edgedetect.dly_315ns_1.bypass_enable_w\[5\] 0.15fF
C1169 edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.out edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.out 0.49fF
C1170 clkgen.delay_155ns_3.genblk1\[0\].dly_binary.in clkgen.delay_155ns_3.genblk1\[0\].dly_binary.signal_w\[1\] 0.17fF
C1171 clkgen.delay_155ns_1.bypass_enable_w\[3\] clkgen.delay_155ns_1.bypass_enable_w\[0\] 0.16fF
C1172 dlycontrol2_in[1] clkgen.delay_155ns_1.bypass_enable_w\[4\] 1.20fF
C1173 clkgen.delay_155ns_3.genblk1\[0\].dly_binary.in clkgen.delay_155ns_3.genblk1\[1\].dly_binary.bypass_in 0.11fF
C1174 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[32\] edgedetect.dly_315ns_1.bypass_enable_w\[5\] 0.14fF
C1175 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[16\] clkgen.delay_155ns_3.genblk1\[4\].dly_binary.bypass_in 0.13fF
C1176 dlycontrol4_in[0] edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.bypass_in 3.56fF
C1177 VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[31\].delay_unit/mid 0.43fF
C1178 clkgen.delay_155ns_1.genblk1\[2\].dly_binary.genblk1\[0\].delay_unit/mid clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit/mid 0.14fF
C1179 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.bypass_in edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[29\].delay_unit/mid 0.15fF
C1180 dlycontrol2_in[0] dlycontrol1_in[3] 0.34fF
C1181 clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[4\] sample_n_2 0.15fF
C1182 VDD clkgen.delay_155ns_3.genblk1\[4\].dly_binary.bypass_in 1.51fF
C1183 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[15\] VDD 1.32fF
C1184 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit/mid VDD 0.36fF
C1185 sample_n_in dlycontrol1_in[0] 1.01fF
C1186 nsample_n_in VDD 1.51fF
C1187 dlycontrol2_in[1] dlycontrol1_in[3] 0.10fF
C1188 clkgen.delay_155ns_1.enable_dlycontrol_w clkgen.delay_155ns_2.enable_dlycontrol_w 0.11fF
C1189 clkgen.delay_155ns_3.bypass_enable_w\[4\] VDD 0.39fF
C1190 dlycontrol1_in[0] clkgen.delay_155ns_1.genblk1\[3\].dly_binary.bypass_in 0.36fF
C1191 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[7\] clkgen.delay_155ns_2.bypass_enable_w\[1\] 0.25fF
C1192 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[6\] edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[8\] 0.34fF
C1193 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[11\] VDD 0.85fF
C1194 dlycontrol1_in[2] dlycontrol1_in[1] 3.45fF
C1195 VDD clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit/mid 0.38fF
C1196 clkgen.delay_155ns_1.bypass_enable_w\[3\] VDD 0.46fF
C1197 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.out clkgen.delay_155ns_2.genblk1\[2\].dly_binary.bypass_in 0.18fF
C1198 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit/mid edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[6\] 0.14fF
C1199 VDD edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.genblk1\[1\].delay_unit/mid 0.12fF
C1200 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit/a_1632_71# clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[5\] 0.13fF
C1201 edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.out edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[8\] 0.16fF
C1202 VDD clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit/mid 0.23fF
C1203 dlycontrol4_in[1] edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.bypass_in 2.23fF
C1204 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[8\] clkgen.delay_155ns_3.genblk1\[0\].dly_binary.bypass_in 0.21fF
C1205 clkgen.delay_155ns_2.genblk1\[1\].dly_binary.bypass_in clkgen.delay_155ns_3.enable_dlycontrol_w 0.10fF
C1206 clkgen.delay_155ns_2.genblk1\[0\].dly_binary.out VDD 1.23fF
C1207 clkgen.clk_dig_out clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[0\].delay_unit/mid 0.12fF
C1208 clkgen.enable_loop_in clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit/mid 0.10fF
C1209 VDD edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.out 2.18fF
C1210 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[16\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[0\] 0.15fF
C1211 VDD clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit/a_1691_329# 0.13fF
C1212 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit/mid VDD 0.68fF
C1213 clkgen.delay_155ns_2.genblk1\[1\].dly_binary.signal_w\[0\] clkgen.delay_155ns_1.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit/mid 0.12fF
C1214 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit/mid VDD 0.12fF
C1215 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[4\] dlycontrol1_in[0] 0.23fF
C1216 start_conv_in edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[7\] 0.38fF
C1217 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[0\] start_conv_in 0.50fF
C1218 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[0\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.out 0.71fF
C1219 clkgen.delay_155ns_3.bypass_enable_w\[2\] start_conv_in 0.24fF
C1220 sample_n_in clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[0\] 1.30fF
C1221 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[16\] clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit/mid 0.16fF
C1222 VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[2\] 0.63fF
C1223 edgedetect.start_conv_edge_w clkgen.delay_155ns_3.genblk1\[0\].dly_binary.in 0.34fF
C1224 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit/mid clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[12\] 0.17fF
C1225 clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[0\] clkgen.delay_155ns_1.genblk1\[3\].dly_binary.bypass_in 0.78fF
C1226 dlycontrol1_in[0] dlycontrol1_in[1] 0.87fF
C1227 sample_n_in clkgen.delay_155ns_1.genblk1\[3\].dly_binary.bypass_in 1.43fF
C1228 VDD clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit/mid 0.41fF
C1229 VDD clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[0\] 2.27fF
C1230 clkgen.delay_155ns_3.genblk1\[0\].dly_binary.signal_w\[0\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[7\] 0.17fF
C1231 clkgen.delay_155ns_2.genblk1\[0\].dly_binary.out dlycontrol1_in[3] 0.17fF
C1232 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit/mid clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[9\] 0.11fF
C1233 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.out clkgen.delay_155ns_2.genblk1\[4\].dly_binary.bypass_in 4.10fF
C1234 sample_n_in clkgen.delay_155ns_2.genblk1\[1\].dly_binary.bypass_in 2.74fF
C1235 clkgen.delay_155ns_1.genblk1\[0\].dly_binary.genblk1\[0\].delay_unit/mid clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[0\] 0.11fF
C1236 edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.bypass_in sample_p_in 0.10fF
C1237 clkgen.delay_155ns_1.genblk1\[0\].dly_binary.out_mux/a_505_21# VDD 0.11fF
C1238 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[2\].delay_unit/mid clkgen.delay_155ns_3.genblk1\[3\].dly_binary.out 0.11fF
C1239 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit/mid clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[0\].delay_unit/mid 0.12fF
C1240 clkgen.delay_155ns_2.genblk1\[1\].dly_binary.bypass_in clkgen.delay_155ns_1.genblk1\[3\].dly_binary.bypass_in 0.73fF
C1241 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit/mid dlycontrol2_in[3] 0.14fF
C1242 clkgen.delay_155ns_1.genblk1\[1\].dly_binary.bypass_in clkgen.delay_155ns_1.genblk1\[0\].dly_binary.out 0.11fF
C1243 VDD clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit/mid 0.26fF
C1244 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[3\].delay_unit/mid edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.bypass_in 0.15fF
C1245 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit/mid clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[16\] 0.12fF
C1246 dlycontrol4_in[2] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[32\] 0.95fF
C1247 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit/a_1632_71# clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[2\] 0.14fF
C1248 clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[4\] clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[1\] 0.27fF
C1249 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit/mid edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[12\] 0.21fF
C1250 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.bypass_in edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.out 0.14fF
C1251 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.out dlycontrol4_in[2] 0.10fF
C1252 clkgen.delay_155ns_3.genblk1\[0\].dly_binary.signal_w\[0\] VDD 2.02fF
C1253 clkgen.delay_155ns_1.genblk1\[0\].dly_binary.signal_w\[1\] VDD 0.35fF
C1254 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[8\] dlycontrol2_in[2] 0.17fF
C1255 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[0\] VDD 1.40fF
C1256 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[0\] VDD 0.89fF
C1257 dlycontrol2_in[3] dlycontrol3_in[1] 1.79fF
C1258 edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.signal_w\[1\] sample_p_in 0.19fF
C1259 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit/mid VDD 0.31fF
C1260 clkgen.delay_155ns_1.genblk1\[1\].dly_binary.bypass_in clkgen.delay_155ns_1.genblk1\[1\].dly_binary.signal_w\[2\] 1.34fF
C1261 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.bypass_in dlycontrol2_in[2] 0.14fF
C1262 VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[26\].delay_unit/a_1691_329# 0.13fF
C1263 enable_dlycontrol_in clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[10\] 0.17fF
C1264 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.signal_w\[0\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.out 0.34fF
C1265 dlycontrol4_in[2] dlycontrol4_in[3] 0.76fF
C1266 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit/mid clkgen.delay_155ns_3.genblk1\[0\].dly_binary.bypass_in 0.18fF
C1267 clkgen.delay_155ns_3.genblk1\[0\].dly_binary.in clkgen.delay_155ns_1.genblk1\[1\].dly_binary.out 0.86fF
C1268 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.bypass_in edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[32\] 0.51fF
C1269 sample_n_in dlycontrol1_in[1] 4.94fF
C1270 dlycontrol2_in[3] dlycontrol2_in[2] 0.62fF
C1271 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[12\].delay_unit/mid clkgen.delay_155ns_3.enable_dlycontrol_w 0.17fF
C1272 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.out clkgen.delay_155ns_3.genblk1\[0\].dly_binary.signal_w\[1\] 0.15fF
C1273 clkgen.delay_155ns_3.genblk1\[2\].dly_binary.genblk1\[1\].delay_unit/a_1632_71# clkgen.delay_155ns_3.genblk1\[2\].dly_binary.signal_w\[2\] 0.14fF
C1274 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.bypass_in dlycontrol1_in[1] 0.18fF
C1275 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.out sample_p_in 0.12fF
C1276 VDD clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[5\] 0.72fF
C1277 nsample_n_4 VDD 0.36fF
C1278 dlycontrol2_in[1] clkgen.delay_155ns_2.genblk1\[1\].dly_binary.signal_w\[2\] 0.97fF
C1279 clkgen.delay_155ns_3.genblk1\[0\].dly_binary.in clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[16\] 0.25fF
C1280 VDD clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit/mid 0.46fF
C1281 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[3\] VDD 0.70fF
C1282 VDD clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit/mid 0.19fF
C1283 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.out dlycontrol3_in[0] 1.62fF
C1284 sample_n_3 clk_dig_out 0.22fF
C1285 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.genblk1\[0\].delay_unit/mid clkgen.delay_155ns_2.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit/mid 0.14fF
C1286 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.out edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.out 0.15fF
C1287 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[4\] clkgen.delay_155ns_2.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit/a_1632_71# 0.17fF
C1288 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit/a_1632_71# edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[2\] 0.14fF
C1289 ndecision_finish_in clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[16\] 2.58fF
C1290 dlycontrol2_in[0] dlycontrol1_in[2] 1.24fF
C1291 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.bypass_in dlycontrol4_in[5] 0.19fF
C1292 clkgen.delay_155ns_3.genblk1\[2\].dly_binary.out clkgen.delay_155ns_3.genblk1\[2\].dly_binary.bypass_in 0.10fF
C1293 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[0\] edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.bypass_in 0.44fF
C1294 clkgen.delay_155ns_3.genblk1\[2\].dly_binary.bypass_in dlycontrol3_in[1] 0.18fF
C1295 VDD outbuf_5/a_27_47# 0.16fF
C1296 clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[4\] clkgen.delay_155ns_1.genblk1\[2\].dly_binary.bypass_in 0.70fF
C1297 nsample_p_4 VDD 0.17fF
C1298 VDD edgedetect.dly_315ns_1.bypass_enable_w\[0\] 0.34fF
C1299 clkgen.delay_155ns_2.genblk1\[1\].dly_binary.out clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[8\] 1.41fF
C1300 VDD edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.signal_w\[0\] 2.31fF
C1301 clkgen.delay_155ns_3.genblk1\[1\].dly_binary.out clkgen.delay_155ns_3.genblk1\[0\].dly_binary.bypass_in 0.16fF
C1302 sample_p_2 clkgen.delay_155ns_3.genblk1\[2\].dly_binary.signal_w\[4\] 0.12fF
C1303 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[30\].delay_unit/mid edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[30\] 0.25fF
C1304 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.out dlycontrol1_in[4] 0.75fF
C1305 dlycontrol4_in[5] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.out 0.12fF
C1306 VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.out_mux/a_505_21# 0.13fF
C1307 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.out clkgen.delay_155ns_3.genblk1\[3\].dly_binary.bypass_in 0.29fF
C1308 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.out dlycontrol4_in[3] 4.42fF
C1309 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[4\] clkgen.clk_dig_delayed_w 0.23fF
C1310 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.out clkgen.delay_155ns_3.genblk1\[0\].dly_binary.in 2.05fF
C1311 clkgen.delay_155ns_2.bypass_enable_w\[1\] dlycontrol3_in[4] 0.15fF
C1312 sample_p_in clkgen.delay_155ns_3.genblk1\[3\].dly_binary.bypass_in 1.14fF
C1313 edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[0\] edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.bypass_in 0.56fF
C1314 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[13\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[13\].delay_unit/mid 0.31fF
C1315 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[23\] edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.bypass_in 0.31fF
C1316 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.in edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.out 0.23fF
C1317 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[28\] VDD 3.29fF
C1318 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[1\] clkgen.delay_155ns_1.genblk1\[0\].dly_binary.bypass_in 0.24fF
C1319 edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.bypass_in edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[1\] 0.44fF
C1320 dlycontrol2_in[4] clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[6\] 0.23fF
C1321 VDD clkgen.delay_155ns_1.genblk1\[1\].dly_binary.signal_w\[1\] 1.06fF
C1322 clkgen.delay_155ns_3.genblk1\[1\].dly_binary.signal_w\[2\] dlycontrol3_in[0] 0.28fF
C1323 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit/mid clkgen.delay_155ns_2.enable_dlycontrol_w 0.14fF
C1324 clkgen.delay_155ns_2.genblk1\[0\].dly_binary.bypass_in clkgen.delay_155ns_2.genblk1\[4\].dly_binary.bypass_in 0.14fF
C1325 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.genblk1\[0\].delay_unit/mid dlycontrol2_in[2] 0.10fF
C1326 VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[32\] 3.95fF
C1327 clkgen.delay_155ns_2.genblk1\[1\].dly_binary.out clkgen.delay_155ns_2.genblk1\[1\].dly_binary.signal_w\[0\] 0.65fF
C1328 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit/a_1632_71# clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[14\] 0.13fF
C1329 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit/mid clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[16\] 0.11fF
C1330 dlycontrol4_in[2] sample_p_4 1.21fF
C1331 VDD clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[4\] 0.62fF
C1332 edgedetect.start_conv_edge_w edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit/mid 0.11fF
C1333 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.in edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.bypass_in 0.13fF
C1334 clkgen.delay_155ns_2.genblk1\[1\].dly_binary.signal_w\[2\] clkgen.delay_155ns_2.genblk1\[0\].dly_binary.out 0.37fF
C1335 clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[4\] clkgen.delay_155ns_1.genblk1\[2\].dly_binary.out 2.26fF
C1336 dlycontrol2_in[1] clkgen.delay_155ns_1.genblk1\[0\].dly_binary.bypass_in 0.16fF
C1337 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.bypass_in clkgen.delay_155ns_3.genblk1\[0\].dly_binary.bypass_in 0.49fF
C1338 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.in edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.bypass_in 1.86fF
C1339 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.out VDD 1.60fF
C1340 VDD edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.genblk1\[0\].delay_unit/mid 0.33fF
C1341 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.bypass_in edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[30\].delay_unit/mid 0.12fF
C1342 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.in dlycontrol4_in[0] 0.34fF
C1343 clkgen.clk_dig_delayed_w sample_n_2 0.39fF
C1344 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[25\].delay_unit/mid edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[26\].delay_unit/mid 0.12fF
C1345 VDD clkgen.delay_155ns_3.bypass_enable_w\[0\] 1.46fF
C1346 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit/mid clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[12\] 0.11fF
C1347 clkgen.delay_155ns_2.genblk1\[1\].dly_binary.bypass_in clkgen.delay_155ns_1.genblk1\[0\].dly_binary.out 0.11fF
C1348 clkgen.delay_155ns_2.genblk1\[0\].dly_binary.out clkgen.delay_155ns_1.genblk1\[1\].dly_binary.bypass_in 0.16fF
C1349 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[11\].delay_unit/mid edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[28\].delay_unit/mid 0.13fF
C1350 sample_n_in clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[2\].delay_unit/mid 0.21fF
C1351 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit/mid edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.bypass_in 0.22fF
C1352 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit/mid VDD 0.41fF
C1353 nsample_p_4 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.bypass_in 0.28fF
C1354 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit/mid clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[3\] 0.11fF
C1355 clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[1\] clkgen.delay_155ns_1.genblk1\[1\].dly_binary.signal_w\[1\] 0.12fF
C1356 VDD dlycontrol4_in[5] 2.06fF
C1357 nsample_p_1 edgedetect.dly_315ns_1.enable_dlycontrol_w 0.20fF
C1358 VDD dlycontrol4_in[3] 1.19fF
C1359 VDD clkgen.delay_155ns_1.genblk1\[2\].dly_binary.genblk1\[1\].delay_unit/mid 0.29fF
C1360 clkgen.delay_155ns_3.genblk1\[0\].dly_binary.in clkgen.delay_155ns_2.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit/mid 0.18fF
C1361 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.bypass_in clkgen.delay_155ns_1.genblk1\[0\].dly_binary.bypass_in 0.17fF
C1362 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.out edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[8\] 0.24fF
C1363 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[20\].delay_unit/mid edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[21\].delay_unit/mid 0.11fF
C1364 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[8\] clkgen.delay_155ns_3.enable_dlycontrol_w 0.11fF
C1365 sample_p_in dlycontrol3_in[3] 0.14fF
C1366 clkgen.delay_155ns_3.bypass_enable_w\[1\] clkgen.delay_155ns_3.enable_dlycontrol_w 0.25fF
C1367 dlycontrol4_in[1] edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.in 0.11fF
C1368 clkgen.delay_155ns_3.genblk1\[2\].dly_binary.out clkgen.delay_155ns_3.genblk1\[3\].dly_binary.bypass_in 0.43fF
C1369 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[2\].delay_unit/mid VDD 0.47fF
C1370 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.bypass_in edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[32\] 0.32fF
C1371 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[8\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.bypass_in 4.47fF
C1372 dlycontrol4_in[1] edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[15\] 0.25fF
C1373 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[2\] clkgen.delay_155ns_3.genblk1\[3\].dly_binary.out 0.10fF
C1374 VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[29\].delay_unit/mid 0.23fF
C1375 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[13\] dlycontrol4_in[0] 0.17fF
C1376 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.genblk1\[1\].delay_unit/mid VDD 0.33fF
C1377 VDD clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[3\] 0.62fF
C1378 VDD clkgen.delay_155ns_2.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit/mid 0.28fF
C1379 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[0\].delay_unit/mid clkgen.delay_155ns_2.genblk1\[4\].dly_binary.bypass_in 0.16fF
C1380 VDD clkgen.delay_155ns_3.genblk1\[3\].dly_binary.out 0.87fF
C1381 dlycontrol2_in[0] sample_n_in 0.10fF
C1382 clkgen.delay_155ns_1.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit/a_1632_71# clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[3\] 0.13fF
C1383 edgedetect.ena_in enable_dlycontrol_in 1.61fF
C1384 dlycontrol2_in[0] clkgen.delay_155ns_1.genblk1\[3\].dly_binary.bypass_in 0.16fF
C1385 dlycontrol2_in[0] clkgen.delay_155ns_2.genblk1\[1\].dly_binary.genblk1\[0\].delay_unit/mid 0.11fF
C1386 dlycontrol3_in[2] sample_p_in 1.60fF
C1387 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[11\] VDD 0.74fF
C1388 clkgen.enable_loop_in clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[2\] 0.59fF
C1389 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.bypass_in VDD 2.58fF
C1390 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[10\] VDD 0.55fF
C1391 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[3\] clkgen.delay_155ns_1.genblk1\[0\].dly_binary.signal_w\[0\] 0.25fF
C1392 sample_n_2 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[16\] 0.24fF
C1393 dlycontrol1_in[0] clkgen.delay_155ns_2.genblk1\[0\].dly_binary.out 0.25fF
C1394 dlycontrol2_in[0] clkgen.delay_155ns_2.genblk1\[1\].dly_binary.bypass_in 0.13fF
C1395 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.out clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[4\] 0.38fF
C1396 dlycontrol4_in[5] edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.bypass_in 0.13fF
C1397 sample_n_1 VDD 0.88fF
C1398 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.bypass_in dlycontrol4_in[3] 0.39fF
C1399 dlycontrol2_in[1] clkgen.delay_155ns_2.genblk1\[1\].dly_binary.bypass_in 1.24fF
C1400 sampledly04/a_523_47# VDD 0.11fF
C1401 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit/mid VDD 0.54fF
C1402 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[7\] clk_dig_out 0.48fF
C1403 ndecision_finish_in dlycontrol2_in[2] 0.19fF
C1404 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit/mid clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[2\] 0.21fF
C1405 VDD clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[12\] 0.97fF
C1406 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[0\] clkgen.delay_155ns_1.genblk1\[0\].dly_binary.bypass_in 1.05fF
C1407 clkgen.delay_155ns_3.genblk1\[2\].dly_binary.out dlycontrol3_in[3] 0.65fF
C1408 VDD edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit/mid 0.29fF
C1409 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.bypass_in clkgen.delay_155ns_2.enable_dlycontrol_w 0.10fF
C1410 VDD sample_p_4 0.88fF
C1411 dlycontrol3_in[3] dlycontrol3_in[1] 1.01fF
C1412 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.bypass_in dlycontrol2_in[3] 0.17fF
C1413 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[4\] VDD 0.70fF
C1414 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[8\] VDD 0.86fF
C1415 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit/mid enable_dlycontrol_in 0.17fF
C1416 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[0\] dlycontrol2_in[1] 4.02fF
C1417 VDD edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit/mid 0.20fF
C1418 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit/mid VDD 0.33fF
C1419 VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[1\] 0.55fF
C1420 sample_p_2 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[3\] 0.40fF
C1421 clkgen.enable_loop_in clkgen.delay_155ns_3.genblk1\[0\].dly_binary.in 0.13fF
C1422 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit/a_1632_71# clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[13\] 0.13fF
C1423 ndecision_finish_in clkgen.delay_155ns_1.genblk1\[0\].dly_binary.signal_w\[0\] 0.19fF
C1424 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit/mid clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[14\] 0.12fF
C1425 dlycontrol2_in[0] dlycontrol1_in[1] 1.54fF
C1426 clkgen.delay_155ns_2.bypass_enable_w\[0\] clkgen.delay_155ns_2.enable_dlycontrol_w 0.10fF
C1427 clkgen.delay_155ns_3.genblk1\[0\].dly_binary.signal_w\[0\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[6\] 0.19fF
C1428 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.out dlycontrol2_in[3] 0.44fF
C1429 VDD clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit/mid 0.36fF
C1430 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[12\].delay_unit/mid edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.bypass_in 0.10fF
C1431 clkgen.delay_155ns_2.genblk1\[1\].dly_binary.genblk1\[0\].delay_unit/mid clkgen.delay_155ns_2.genblk1\[0\].dly_binary.out 0.13fF
C1432 dlycontrol3_in[2] dlycontrol3_in[1] 6.19fF
C1433 VDD clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit/a_1691_329# 0.10fF
C1434 edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[4\] sample_p_2 0.58fF
C1435 clkgen.delay_155ns_3.genblk1\[2\].dly_binary.bypass_in clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[4\] 0.13fF
C1436 clkgen.clk_dig_delayed_w clkgen.delay_155ns_1.genblk1\[1\].dly_binary.genblk1\[0\].delay_unit/mid 0.10fF
C1437 clkgen.delay_155ns_2.genblk1\[1\].dly_binary.bypass_in clkgen.delay_155ns_2.genblk1\[0\].dly_binary.out 0.18fF
C1438 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[2\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[3\] 0.51fF
C1439 edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.bypass_in clkgen.delay_155ns_2.genblk1\[4\].dly_binary.bypass_in 0.16fF
C1440 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[16\] clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[11\] 0.23fF
C1441 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[25\] VDD 1.42fF
C1442 clkgen.delay_155ns_3.genblk1\[0\].dly_binary.signal_w\[0\] clkgen.delay_155ns_3.enable_dlycontrol_w 0.23fF
C1443 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[27\].delay_unit/mid VDD 0.45fF
C1444 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[17\] VDD 0.70fF
C1445 clkgen.delay_155ns_1.genblk1\[0\].dly_binary.in VDD 2.01fF
C1446 VDD edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[7\] 0.59fF
C1447 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[0\] VDD 1.48fF
C1448 VDD clkgen.delay_155ns_3.bypass_enable_w\[2\] 0.18fF
C1449 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.in clkgen.delay_155ns_3.genblk1\[0\].dly_binary.signal_w\[0\] 0.12fF
C1450 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[0\].delay_unit/mid clkgen.delay_155ns_3.genblk1\[0\].dly_binary.in 0.12fF
C1451 edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.signal_w\[0\] sample_p_in 0.37fF
C1452 edgedetect.start_conv_edge_w clkgen.delay_155ns_1.genblk1\[2\].dly_binary.bypass_in 0.56fF
C1453 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit/mid clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[2\] 0.30fF
C1454 clkgen.delay_155ns_1.genblk1\[0\].dly_binary.out clkgen.delay_155ns_1.genblk1\[1\].dly_binary.signal_w\[2\] 0.53fF
C1455 nsample_p_2 VDD 0.20fF
C1456 VDD clkgen.delay_155ns_2.enable_dlycontrol_w 2.35fF
C1457 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit/mid clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[15\] 0.14fF
C1458 edgedetect.dly_315ns_1.enable_dlycontrol_w dlycontrol2_in[4] 2.20fF
C1459 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit/a_1632_71# edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[4\] 0.13fF
C1460 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[1\] edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit/mid 0.25fF
C1461 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.signal_w\[1\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.bypass_in 0.27fF
C1462 clkgen.delay_155ns_2.genblk1\[1\].dly_binary.signal_w\[0\] clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[0\].delay_unit/mid 0.10fF
C1463 clkgen.delay_155ns_2.genblk1\[0\].dly_binary.signal_w\[0\] clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[4\] 0.40fF
C1464 VDD clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[10\] 0.61fF
C1465 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[16\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[32\] 0.14fF
C1466 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[5\] clkgen.delay_155ns_3.bypass_enable_w\[0\] 0.13fF
C1467 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit/a_1632_71# clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[8\] 0.13fF
C1468 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.bypass_in edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[20\].delay_unit/mid 0.14fF
C1469 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.bypass_in clkgen.delay_155ns_3.genblk1\[0\].dly_binary.bypass_in 0.10fF
C1470 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.out edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.bypass_in 0.12fF
C1471 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.bypass_in dlycontrol1_in[4] 0.49fF
C1472 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[12\] edgedetect.dly_315ns_1.enable_dlycontrol_w 0.12fF
C1473 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.out dlycontrol4_in[0] 0.32fF
C1474 VDD clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[4\] 0.97fF
C1475 edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit/mid VDD 0.26fF
C1476 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[29\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.bypass_in 0.19fF
C1477 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit/mid edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[3\] 0.17fF
C1478 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[1\] clkgen.delay_155ns_1.genblk1\[0\].dly_binary.out 0.39fF
C1479 clkgen.clk_comp_out clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit/mid 0.12fF
C1480 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.bypass_in edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.bypass_in 1.07fF
C1481 dlycontrol2_in[0] clkgen.delay_155ns_1.genblk1\[0\].dly_binary.out 0.11fF
C1482 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.bypass_in edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[2\] 0.15fF
C1483 sample_p_2 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[16\] 2.21fF
C1484 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit/mid VDD 0.41fF
C1485 clkgen.delay_155ns_3.genblk1\[1\].dly_binary.bypass_in start_conv_in 0.16fF
C1486 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[4\] clkgen.delay_155ns_1.genblk1\[0\].dly_binary.signal_w\[0\] 0.65fF
C1487 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.out clkgen.delay_155ns_3.genblk1\[1\].dly_binary.signal_w\[2\] 0.14fF
C1488 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[17\].delay_unit/mid edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[18\].delay_unit/mid 0.14fF
C1489 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[5\] dlycontrol3_in[4] 0.35fF
C1490 clkgen.delay_155ns_1.genblk1\[1\].dly_binary.signal_w\[1\] clkgen.delay_155ns_1.genblk1\[0\].dly_binary.bypass_in 0.24fF
C1491 dlycontrol3_in[0] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[32\] 1.79fF
C1492 dlycontrol4_in[1] edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.out 3.78fF
C1493 VDD clkgen.delay_155ns_1.genblk1\[1\].dly_binary.signal_w\[0\] 1.65fF
C1494 clkgen.clk_dig_out clk_dig_out 1.84fF
C1495 nsample_p_2 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.bypass_in 0.31fF
C1496 clkgen.delay_155ns_1.genblk1\[1\].dly_binary.out clkgen.delay_155ns_1.genblk1\[2\].dly_binary.bypass_in 1.37fF
C1497 clkgen.delay_155ns_1.genblk1\[0\].dly_binary.bypass_in clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[4\] 0.12fF
C1498 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[10\].delay_unit/mid clkgen.delay_155ns_2.genblk1\[4\].dly_binary.bypass_in 0.14fF
C1499 clkgen.enable_loop_in clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[4\] 0.10fF
C1500 clkgen.delay_155ns_2.enable_dlycontrol_w clkgen.clk_comp_out 1.59fF
C1501 VDD edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[3\] 0.44fF
C1502 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[4\] clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[2\] 0.31fF
C1503 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[16\] edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[2\] 0.12fF
C1504 clkgen.delay_155ns_3.genblk1\[1\].dly_binary.out clkgen.delay_155ns_3.genblk1\[0\].dly_binary.signal_w\[1\] 0.23fF
C1505 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit/mid VDD 0.41fF
C1506 clkgen.delay_155ns_3.genblk1\[0\].dly_binary.in clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[4\] 0.23fF
C1507 clkgen.delay_155ns_2.genblk1\[1\].dly_binary.out clkgen.clk_dig_delayed_w 0.45fF
C1508 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[10\].delay_unit/a_1632_71# edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[11\] 0.13fF
C1509 dlycontrol3_in[0] clkgen.delay_155ns_3.bypass_enable_w\[0\] 0.40fF
C1510 edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.bypass_in edgedetect.dly_315ns_1.enable_dlycontrol_w 0.27fF
C1511 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[0\] clkgen.delay_155ns_1.genblk1\[1\].dly_binary.signal_w\[0\] 0.52fF
C1512 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[2\] clkgen.delay_155ns_1.genblk1\[1\].dly_binary.signal_w\[1\] 0.52fF
C1513 dlycontrol2_in[1] clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[5\] 0.14fF
C1514 clkgen.delay_155ns_2.genblk1\[1\].dly_binary.bypass_in clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[5\] 0.15fF
C1515 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit/mid VDD 0.40fF
C1516 dlycontrol4_in[1] dlycontrol4_in[0] 4.05fF
C1517 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[0\] clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[0\] 0.19fF
C1518 clkgen.delay_155ns_3.genblk1\[0\].dly_binary.in clkgen.delay_155ns_2.genblk1\[4\].dly_binary.bypass_in 0.37fF
C1519 clkgen.clk_dig_out clkgen.delay_155ns_2.genblk1\[4\].dly_binary.bypass_in 0.13fF
C1520 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.bypass_in clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit/mid 0.12fF
C1521 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.bypass_in edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[10\].delay_unit/mid 0.16fF
C1522 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[4\] clkgen.delay_155ns_3.enable_dlycontrol_w 0.11fF
C1523 VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[20\].delay_unit/mid 0.36fF
C1524 VDD clkgen.delay_155ns_3.genblk1\[0\].dly_binary.bypass_in 2.61fF
C1525 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit/mid clkgen.delay_155ns_3.genblk1\[1\].dly_binary.bypass_in 0.12fF
C1526 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit/mid edgedetect.dly_315ns_1.bypass_enable_w\[2\] 0.12fF
C1527 edgedetect.dly_315ns_1.bypass_enable_w\[3\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[19\].delay_unit/mid 0.19fF
C1528 edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit/mid dlycontrol3_in[3] 0.14fF
C1529 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[30\].delay_unit/mid VDD 0.23fF
C1530 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[5\] clkgen.delay_155ns_1.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit/mid 0.21fF
C1531 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[10\].delay_unit/mid VDD 0.26fF
C1532 clkgen.delay_155ns_2.bypass_enable_w\[1\] clkgen.delay_155ns_1.bypass_enable_w\[0\] 0.70fF
C1533 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit/mid clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit/mid 0.11fF
C1534 clkgen.enable_loop_in sample_n_2 0.19fF
C1535 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[7\] clk_dig_out 0.51fF
C1536 sample_n_2 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[2\] 0.16fF
C1537 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[16\].delay_unit/a_1632_71# edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[17\] 0.14fF
C1538 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[31\].delay_unit/mid edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.bypass_in 0.20fF
C1539 ndecision_finish_in clkgen.delay_155ns_2.genblk1\[4\].dly_binary.bypass_in 0.20fF
C1540 edgedetect.ena_in clkgen.delay_155ns_1.genblk1\[3\].dly_binary.out 0.27fF
C1541 edgedetect.start_conv_edge_w clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[16\] 0.65fF
C1542 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.out edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.in 0.35fF
C1543 VDD edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.out_mux/a_505_21# 0.11fF
C1544 dlycontrol2_in[0] dlycontrol2_in[1] 0.68fF
C1545 dlycontrol1_in[2] sample_n_1 0.44fF
C1546 edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.signal_w\[0\] edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[1\] 0.13fF
C1547 clkgen.clk_dig_out ena_in 0.30fF
C1548 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[2\].delay_unit/mid clkgen.delay_155ns_1.genblk1\[0\].dly_binary.bypass_in 0.17fF
C1549 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[5\] sample_p_4 0.15fF
C1550 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit/a_1632_71# edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[7\] 0.13fF
C1551 clkgen.delay_155ns_2.genblk1\[0\].dly_binary.out clkgen.delay_155ns_1.genblk1\[0\].dly_binary.out 0.64fF
C1552 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[0\] clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[5\] 0.38fF
C1553 clkgen.clk_dig_out clkgen.delay_155ns_1.genblk1\[4\].dly_binary.out 0.28fF
C1554 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[8\] sample_p_in 0.14fF
C1555 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[13\] edgedetect.dly_315ns_1.bypass_enable_w\[0\] 0.17fF
C1556 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit/mid dlycontrol4_in[1] 0.10fF
C1557 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[4\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[5\] 0.15fF
C1558 clkgen.delay_155ns_1.genblk1\[0\].dly_binary.bypass_in clkgen.delay_155ns_2.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit/mid 0.19fF
C1559 clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[0\] clkgen.delay_155ns_1.genblk1\[1\].dly_binary.signal_w\[1\] 0.26fF
C1560 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.signal_w\[0\] edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[8\] 0.25fF
C1561 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.signal_w\[1\] edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.out 0.28fF
C1562 clkgen.delay_155ns_3.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit/mid start_conv_in 0.14fF
C1563 clkgen.delay_155ns_2.bypass_enable_w\[1\] VDD 2.26fF
C1564 VDD outbuf_6/a_27_47# 0.13fF
C1565 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.in dlycontrol4_in[5] 0.13fF
C1566 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit/mid edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.out 0.14fF
C1567 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[0\] clkgen.delay_155ns_3.genblk1\[3\].dly_binary.bypass_in 0.89fF
C1568 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit/mid dlycontrol3_in[4] 0.31fF
C1569 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[2\] VDD 0.67fF
C1570 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.out edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit/mid 0.16fF
C1571 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.bypass_in dlycontrol3_in[3] 0.11fF
C1572 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[0\].delay_unit/mid VDD 0.41fF
C1573 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[20\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[21\] 0.10fF
C1574 edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.out edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.bypass_in 1.51fF
C1575 dlycontrol4_in[0] edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.out 0.30fF
C1576 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.out_mux/a_505_21# VDD 0.11fF
C1577 VDD edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[10\].delay_unit/mid 0.30fF
C1578 sample_n_1 dlycontrol1_in[0] 0.26fF
C1579 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[12\] clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[16\] 0.50fF
C1580 nsample_n_1 VDD 0.25fF
C1581 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit/mid edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[14\] 0.18fF
C1582 dlycontrol2_in[1] clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit/mid 0.12fF
C1583 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit/mid clkgen.delay_155ns_2.genblk1\[1\].dly_binary.signal_w\[0\] 0.12fF
C1584 clkgen.delay_155ns_2.bypass_enable_w\[1\] dlycontrol1_in[3] 0.62fF
C1585 edgedetect.start_conv_edge_w enable_dlycontrol_in 0.20fF
C1586 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit/mid VDD 0.42fF
C1587 edgedetect.ena_in VDD 1.02fF
C1588 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[8\] VDD 2.27fF
C1589 clkgen.delay_155ns_1.genblk1\[1\].dly_binary.out dlycontrol3_in[4] 0.74fF
C1590 nsample_p_in sample_p_in 0.72fF
C1591 dlycontrol2_in[0] clkgen.delay_155ns_2.genblk1\[0\].dly_binary.out 0.12fF
C1592 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[23\].delay_unit/a_1632_71# edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[24\] 0.13fF
C1593 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.out clkgen.delay_155ns_2.genblk1\[1\].dly_binary.out 3.32fF
C1594 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[1\] clkgen.delay_155ns_3.genblk1\[0\].dly_binary.bypass_in 0.18fF
C1595 VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[22\] 0.67fF
C1596 dlycontrol2_in[4] dlycontrol2_in[3] 0.58fF
C1597 clkgen.enable_loop_in clkgen.delay_155ns_1.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit/mid 0.20fF
C1598 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit/mid clkgen.delay_155ns_1.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit/mid 0.10fF
C1599 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[2\] clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit/mid 0.21fF
C1600 dlycontrol4_in[1] edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.out 0.45fF
C1601 clkgen.delay_155ns_3.bypass_enable_w\[4\] clkgen.delay_155ns_3.genblk1\[4\].dly_binary.bypass_in 0.31fF
C1602 edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[0\] sample_p_4 0.26fF
C1603 edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.out sample_p_4 0.41fF
C1604 clkgen.delay_155ns_3.genblk1\[0\].dly_binary.in dlycontrol1_in[4] 0.14fF
C1605 dlycontrol3_in[4] clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[16\] 0.43fF
C1606 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit/mid dlycontrol2_in[2] 0.10fF
C1607 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit/mid VDD 0.36fF
C1608 clkgen.clk_dig_out dlycontrol1_in[4] 0.10fF
C1609 clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[0\] clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[3\] 0.16fF
C1610 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[10\].delay_unit/a_1632_71# edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[11\] 0.13fF
C1611 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[8\] dlycontrol3_in[1] 0.18fF
C1612 ena_in clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[8\] 0.12fF
C1613 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit/mid VDD 0.23fF
C1614 start_conv_in clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[16\] 0.97fF
C1615 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit/mid VDD 0.22fF
C1616 clkgen.delay_155ns_2.genblk1\[1\].dly_binary.signal_w\[0\] VDD 2.15fF
C1617 inbuf_3/a_27_47# VDD 0.10fF
C1618 dlycontrol3_in[4] edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit/mid 0.18fF
C1619 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.out edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[0\] 0.22fF
C1620 VDD clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit/mid 0.22fF
C1621 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit/mid VDD 0.36fF
C1622 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[1\] clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[0\] 0.59fF
C1623 ndecision_finish_in dlycontrol1_in[4] 0.22fF
C1624 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit/a_1632_71# clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[7\] 0.13fF
C1625 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[8\] dlycontrol1_in[3] 0.11fF
C1626 clkgen.delay_155ns_1.genblk1\[2\].dly_binary.out_mux/a_505_21# VDD 0.13fF
C1627 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[0\] clkgen.delay_155ns_2.genblk1\[1\].dly_binary.signal_w\[0\] 0.31fF
C1628 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.out clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit/mid 0.14fF
C1629 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[0\] clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit/mid 0.11fF
C1630 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[0\].delay_unit/mid clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[2\] 0.17fF
C1631 clkgen.clk_dig_out sample_n_3 0.45fF
C1632 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit/mid clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[15\] 0.14fF
C1633 sample_n_1 clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[0\] 0.37fF
C1634 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[21\].delay_unit/mid edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[21\] 0.23fF
C1635 VDD edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[3\] 0.98fF
C1636 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit/mid VDD 0.32fF
C1637 sample_n_in sample_n_1 0.30fF
C1638 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[0\] dlycontrol4_in[0] 0.44fF
C1639 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[16\] clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[4\] 0.73fF
C1640 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[14\] VDD 0.64fF
C1641 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[3\] VDD 0.59fF
C1642 clkgen.delay_155ns_3.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit/mid VDD 0.51fF
C1643 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.bypass_in clkgen.delay_155ns_2.genblk1\[1\].dly_binary.bypass_in 0.17fF
C1644 VDD clkgen.delay_155ns_2.bypass_enable_w\[2\] 1.31fF
C1645 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[10\] clkgen.delay_155ns_2.genblk1\[1\].dly_binary.bypass_in 0.25fF
C1646 clkgen.delay_155ns_1.genblk1\[0\].dly_binary.in clkgen.delay_155ns_1.genblk1\[0\].dly_binary.bypass_in 0.28fF
C1647 clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[4\] VDD 2.09fF
C1648 VDD clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[1\] 0.67fF
C1649 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[8\] clkgen.delay_155ns_3.genblk1\[2\].dly_binary.signal_w\[3\] 0.35fF
C1650 dlycontrol3_in[4] sample_p_in 0.31fF
C1651 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.out edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[4\].delay_unit/mid 0.11fF
C1652 edgedetect.dly_315ns_1.enable_dlycontrol_w dlycontrol3_in[3] 1.33fF
C1653 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[7\] edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[6\] 0.10fF
C1654 clkgen.delay_155ns_2.genblk1\[0\].dly_binary.bypass_in clkgen.clk_dig_out 1.75fF
C1655 VDD clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit/mid 0.27fF
C1656 sample_p_in start_conv_in 0.32fF
C1657 dlycontrol2_in[4] clkgen.delay_155ns_3.genblk1\[2\].dly_binary.bypass_in 2.31fF
C1658 clkgen.delay_155ns_3.genblk1\[0\].dly_binary.signal_w\[0\] clkgen.delay_155ns_3.genblk1\[2\].dly_binary.signal_w\[1\] 0.15fF
C1659 VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[2\].delay_unit/mid 0.18fF
C1660 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.bypass_in clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit/mid 0.14fF
C1661 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[0\] edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[0\] 2.48fF
C1662 edgedetect.dly_315ns_1.enablebuffer/a_27_47# VDD 0.18fF
C1663 clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[4\] clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[0\] 2.64fF
C1664 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[0\] clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[0\].delay_unit/mid 0.32fF
C1665 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit/mid dlycontrol1_in[4] 0.13fF
C1666 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit/mid clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[16\] 0.10fF
C1667 clkgen.delay_155ns_2.genblk1\[1\].dly_binary.bypass_in clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[12\] 0.10fF
C1668 dlycontrol4_in[1] edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[0\] 0.37fF
C1669 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[24\] VDD 1.64fF
C1670 clkgen.delay_155ns_3.bypass_enable_w\[4\] clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[0\] 0.38fF
C1671 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[16\] VDD 0.77fF
C1672 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[2\].delay_unit/a_1632_71# edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[3\] 0.13fF
C1673 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit/mid clkgen.clk_comp_out 0.16fF
C1674 VDD edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[6\] 0.76fF
C1675 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[6\] VDD 0.74fF
C1676 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit/a_1632_71# clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[3\] 0.14fF
C1677 clkgen.delay_155ns_2.enable_dlycontrol_w clkgen.delay_155ns_3.enable_dlycontrol_w 0.17fF
C1678 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit/mid clkgen.delay_155ns_1.genblk1\[3\].dly_binary.bypass_in 0.17fF
C1679 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[4\].delay_unit/mid clkgen.delay_155ns_3.genblk1\[2\].dly_binary.signal_w\[4\] 0.15fF
C1680 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit/a_1632_71# clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[3\] 0.13fF
C1681 clkgen.delay_155ns_1.genblk1\[0\].dly_binary.signal_w\[1\] clkgen.delay_155ns_1.genblk1\[0\].dly_binary.genblk1\[0\].delay_unit/a_1632_71# 0.13fF
C1682 sample_n_2 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[3\] 0.26fF
C1683 edgedetect.dly_315ns_1.bypass_enable_w\[4\] dlycontrol2_in[4] 1.83fF
C1684 edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[4\] edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[1\] 1.19fF
C1685 clkgen.delay_155ns_2.genblk1\[1\].dly_binary.out dlycontrol2_in[2] 2.30fF
C1686 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.bypass_in clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[7\] 0.28fF
C1687 sample_n_in clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit/mid 0.12fF
C1688 clkgen.delay_155ns_3.genblk1\[2\].dly_binary.genblk1\[1\].delay_unit/mid VDD 0.21fF
C1689 edgedetect.dly_315ns_1.bypass_enable_w\[3\] edgedetect.dly_315ns_1.bypass_enable_w\[4\] 0.41fF
C1690 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.signal_w\[0\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.bypass_in 2.77fF
C1691 sample_p_in enable_dlycontrol_in 1.27fF
C1692 VDD clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[9\] 0.58fF
C1693 sample_n_1 dlycontrol1_in[1] 0.64fF
C1694 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[16\] clkgen.delay_155ns_3.genblk1\[0\].dly_binary.bypass_in 2.19fF
C1695 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[7\] clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[6\] 0.16fF
C1696 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.bypass_in sample_p_in 0.14fF
C1697 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[28\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.bypass_in 0.12fF
C1698 clkgen.delay_155ns_1.genblk1\[1\].dly_binary.signal_w\[2\] clkgen.delay_155ns_1.genblk1\[1\].dly_binary.signal_w\[1\] 0.11fF
C1699 VDD clk_comp_out 1.31fF
C1700 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[16\] clkgen.delay_155ns_3.genblk1\[0\].dly_binary.out 0.14fF
C1701 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.bypass_in edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[32\] 0.11fF
C1702 VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[18\].delay_unit/mid 0.22fF
C1703 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.out clkgen.delay_155ns_3.bypass_enable_w\[0\] 0.45fF
C1704 start_conv_in dlycontrol3_in[1] 0.69fF
C1705 VDD clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[5\] 0.77fF
C1706 VDD clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[11\] 0.79fF
C1707 dlycontrol4_in[4] edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[2\] 0.63fF
C1708 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.out edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.bypass_in 0.84fF
C1709 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.out dlycontrol4_in[5] 1.24fF
C1710 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.out dlycontrol4_in[3] 0.64fF
C1711 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[0\] edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.out 0.19fF
C1712 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.out edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.genblk1\[0\].delay_unit/mid 0.10fF
C1713 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit/mid edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.out 0.14fF
C1714 clkgen.delay_155ns_2.genblk1\[1\].dly_binary.bypass_in clkgen.delay_155ns_2.enable_dlycontrol_w 0.19fF
C1715 sample_p_out edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[8\] 0.31fF
C1716 clkgen.delay_155ns_3.genblk1\[1\].dly_binary.out clkgen.delay_155ns_3.genblk1\[2\].dly_binary.out 1.13fF
C1717 clkgen.delay_155ns_1.genblk1\[2\].dly_binary.genblk1\[1\].delay_unit/mid clkgen.delay_155ns_1.genblk1\[1\].dly_binary.signal_w\[2\] 0.21fF
C1718 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.bypass_in clkgen.delay_155ns_3.genblk1\[0\].dly_binary.in 0.15fF
C1719 ndecision_finish_in clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[8\] 0.92fF
C1720 clkgen.delay_155ns_2.genblk1\[1\].dly_binary.bypass_in clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[10\] 0.21fF
C1721 edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.bypass_in edgedetect.dly_315ns_1.bypass_enable_w\[4\] 0.61fF
C1722 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit/mid clkgen.delay_155ns_3.enable_dlycontrol_w 0.17fF
C1723 dlycontrol4_in[4] edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[4\] 0.73fF
C1724 dlycontrol4_in[0] dlycontrol4_in[5] 0.37fF
C1725 ndecision_finish_in edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[26\] 0.18fF
C1726 clkgen.delay_155ns_2.genblk1\[1\].dly_binary.out clkgen.delay_155ns_2.genblk1\[1\].dly_binary.signal_w\[1\] 0.27fF
C1727 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[25\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[25\].delay_unit/mid 0.23fF
C1728 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.out edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.bypass_in 3.34fF
C1729 clkgen.delay_155ns_3.genblk1\[1\].dly_binary.signal_w\[2\] clkgen.delay_155ns_3.bypass_enable_w\[0\] 1.18fF
C1730 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[2\] clkgen.delay_155ns_3.genblk1\[1\].dly_binary.bypass_in 0.15fF
C1731 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.out dlycontrol4_in[1] 0.47fF
C1732 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.bypass_in ndecision_finish_in 0.82fF
C1733 enable_dlycontrol_in dlycontrol3_in[1] 1.61fF
C1734 VDD clkgen.delay_155ns_3.genblk1\[0\].dly_binary.signal_w\[1\] 0.35fF
C1735 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[2\].delay_unit/a_1632_71# edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[3\] 0.13fF
C1736 clkgen.delay_155ns_3.genblk1\[1\].dly_binary.bypass_in VDD 3.58fF
C1737 clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[0\] clkgen.delay_155ns_1.genblk1\[1\].dly_binary.signal_w\[0\] 0.59fF
C1738 sample_n_in clkgen.delay_155ns_1.genblk1\[1\].dly_binary.signal_w\[0\] 1.02fF
C1739 edgedetect.ena_in dlycontrol1_in[2] 0.19fF
C1740 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.in clkgen.delay_155ns_3.genblk1\[0\].dly_binary.bypass_in 0.23fF
C1741 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[6\] clk_dig_out 0.31fF
C1742 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.bypass_in dlycontrol3_in[1] 0.33fF
C1743 clkgen.delay_155ns_1.genblk1\[2\].dly_binary.bypass_in clk_dig_out 0.19fF
C1744 sample_p_2 VDD 0.82fF
C1745 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.bypass_in clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit/mid 0.15fF
C1746 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit/mid dlycontrol2_in[1] 0.15fF
C1747 clkgen.delay_155ns_1.genblk1\[1\].dly_binary.signal_w\[0\] clkgen.delay_155ns_1.genblk1\[3\].dly_binary.bypass_in 0.50fF
C1748 edgedetect.dly_315ns_1.bypass_enable_w\[1\] edgedetect.dly_315ns_1.enable_dlycontrol_w 0.67fF
C1749 dlycontrol4_in[1] dlycontrol4_in[5] 4.28fF
C1750 dlycontrol4_in[1] dlycontrol4_in[3] 0.21fF
C1751 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.out edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.signal_w\[1\] 0.92fF
C1752 enable_dlycontrol_in dlycontrol2_in[2] 0.13fF
C1753 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[5\] VDD 0.50fF
C1754 VDD edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit/mid 0.13fF
C1755 edgedetect.ena_in clkgen.delay_155ns_1.bypass_enable_w\[2\] 0.24fF
C1756 clkgen.delay_155ns_2.genblk1\[0\].dly_binary.bypass_in clkgen.delay_155ns_1.genblk1\[4\].dly_binary.bypass_in 0.58fF
C1757 dlycontrol2_in[4] dlycontrol3_in[3] 1.15fF
C1758 clkgen.enable_loop_in start_conv_in 0.37fF
C1759 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[25\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[26\].delay_unit/mid 0.18fF
C1760 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[2\] start_conv_in 0.12fF
C1761 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[11\].delay_unit/mid start_conv_in 0.14fF
C1762 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[6\] edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[7\] 0.22fF
C1763 clkgen.delay_155ns_2.genblk1\[0\].dly_binary.signal_w\[1\] VDD 0.27fF
C1764 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit/mid dlycontrol3_in[3] 0.19fF
C1765 ena_in clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[3\] 0.14fF
C1766 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[9\] VDD 0.44fF
C1767 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit/mid clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit/mid 0.11fF
C1768 VDD edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[2\] 0.58fF
C1769 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.out_mux/a_505_21# VDD 0.10fF
C1770 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit/a_1632_71# clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[2\] 0.14fF
C1771 VDD clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit/mid 0.27fF
C1772 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[0\].delay_unit/mid VDD 0.24fF
C1773 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[8\] clkgen.delay_155ns_1.genblk1\[0\].dly_binary.bypass_in 0.51fF
C1774 clkgen.delay_155ns_3.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit/a_1632_71# clkgen.delay_155ns_3.genblk1\[2\].dly_binary.signal_w\[4\] 0.13fF
C1775 clkgen.delay_155ns_3.genblk1\[0\].dly_binary.in clkgen.delay_155ns_3.genblk1\[2\].dly_binary.bypass_in 0.24fF
C1776 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[13\].delay_unit/a_1632_71# edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[14\] 0.15fF
C1777 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[8\] clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[7\] 0.40fF
C1778 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.bypass_in clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[13\] 0.14fF
C1779 start_conv_in clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[6\] 0.22fF
C1780 edgedetect.ena_in dlycontrol1_in[0] 1.07fF
C1781 clkgen.delay_155ns_3.genblk1\[0\].dly_binary.in clkgen.delay_155ns_2.genblk1\[2\].dly_binary.genblk1\[0\].delay_unit/mid 0.13fF
C1782 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[16\] clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit/mid 0.14fF
C1783 ena_in clkgen.delay_155ns_1.genblk1\[2\].dly_binary.bypass_in 3.09fF
C1784 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.genblk1\[0\].delay_unit/mid dlycontrol3_in[3] 0.20fF
C1785 VDD clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[0\] 0.64fF
C1786 dlycontrol2_in[1] clkgen.delay_155ns_2.genblk1\[3\].dly_binary.bypass_in 2.94fF
C1787 dlycontrol2_in[0] sample_n_1 0.52fF
C1788 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.in edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[10\].delay_unit/mid 0.11fF
C1789 clkgen.delay_155ns_1.genblk1\[1\].dly_binary.signal_w\[0\] dlycontrol1_in[1] 1.04fF
C1790 VDD clkgen.delay_155ns_3.genblk1\[1\].dly_binary.genblk1\[0\].delay_unit/mid 0.42fF
C1791 edgedetect.start_conv_edge_w VDD 2.36fF
C1792 VDD clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[3\] 0.55fF
C1793 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[1\] edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.bypass_in 0.30fF
C1794 clkgen.delay_155ns_2.bypass_enable_w\[1\] clkgen.delay_155ns_1.genblk1\[3\].dly_binary.bypass_in 0.15fF
C1795 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.bypass_in clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit/mid 0.18fF
C1796 clkgen.delay_155ns_3.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit/mid VDD 0.44fF
C1797 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.bypass_in clkgen.delay_155ns_3.genblk1\[3\].dly_binary.out 0.38fF
C1798 clkgen.delay_155ns_2.genblk1\[1\].dly_binary.bypass_in clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit/mid 0.23fF
C1799 clkgen.clk_dig_delayed_w VDD 0.66fF
C1800 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[8\] clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[0\] 0.45fF
C1801 dlycontrol4_in[2] sample_p_in 2.46fF
C1802 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[0\] clkgen.delay_155ns_3.genblk1\[0\].dly_binary.bypass_in 1.81fF
C1803 clkgen.delay_155ns_3.genblk1\[0\].dly_binary.in clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[2\] 0.45fF
C1804 VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[21\] 0.78fF
C1805 dlycontrol4_in[5] edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.out 3.79fF
C1806 edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.out dlycontrol4_in[3] 0.58fF
C1807 clkgen.delay_155ns_3.genblk1\[0\].dly_binary.signal_w\[0\] edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.signal_w\[0\] 2.99fF
C1808 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit/mid clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[15\] 0.15fF
C1809 edgedetect.start_conv_edge_w clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[0\] 0.22fF
C1810 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[14\] dlycontrol3_in[0] 0.12fF
C1811 clkgen.delay_155ns_3.genblk1\[1\].dly_binary.signal_w\[1\] clkgen.delay_155ns_3.genblk1\[2\].dly_binary.out 0.11fF
C1812 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit/mid VDD 0.27fF
C1813 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit/mid VDD 0.43fF
C1814 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit/mid dlycontrol2_in[2] 0.13fF
C1815 clkgen.delay_155ns_3.genblk1\[2\].dly_binary.bypass_in dlycontrol3_in[3] 0.14fF
C1816 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.out edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit/mid 0.11fF
C1817 nsample_p_1 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[14\] 0.12fF
C1818 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit/mid clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[0\].delay_unit/mid 0.11fF
C1819 clkgen.delay_155ns_1.genblk1\[0\].dly_binary.in clkgen.delay_155ns_1.genblk1\[1\].dly_binary.signal_w\[2\] 0.52fF
C1820 clkgen.delay_155ns_1.genblk1\[0\].dly_binary.signal_w\[1\] clkgen.delay_155ns_1.genblk1\[1\].dly_binary.signal_w\[1\] 0.45fF
C1821 VDD sample_p_out 0.30fF
C1822 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[16\] clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[15\] 0.15fF
C1823 edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.out edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[3\] 0.73fF
C1824 edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit/mid edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[4\] 0.19fF
C1825 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.bypass_in edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[7\] 0.31fF
C1826 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit/mid clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit/mid 0.11fF
C1827 VDD clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[15\] 1.53fF
C1828 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[0\] edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.bypass_in 1.36fF
C1829 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.bypass_in clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[12\] 0.14fF
C1830 dlycontrol3_in[3] clkgen.delay_155ns_3.genblk1\[2\].dly_binary.genblk1\[0\].delay_unit/mid 0.20fF
C1831 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.bypass_in sample_p_in 0.50fF
C1832 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[21\].delay_unit/a_1632_71# edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[22\] 0.14fF
C1833 start_conv_in clk_dig_out 2.59fF
C1834 sample_p_3 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[3\] 0.18fF
C1835 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.out edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[0\] 0.12fF
C1836 clkgen.delay_155ns_3.genblk1\[0\].dly_binary.signal_w\[0\] clkgen.delay_155ns_3.bypass_enable_w\[0\] 0.46fF
C1837 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[9\].delay_unit/mid start_conv_in 0.13fF
C1838 clkgen.delay_155ns_1.genblk1\[1\].dly_binary.out VDD 1.60fF
C1839 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit/mid clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[0\] 0.17fF
C1840 clkgen.delay_155ns_3.genblk1\[0\].dly_binary.in clkgen.delay_155ns_3.genblk1\[3\].dly_binary.bypass_in 0.15fF
C1841 clkgen.clk_dig_out clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[8\] 0.13fF
C1842 clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[0\] clkgen.delay_155ns_2.genblk1\[1\].dly_binary.signal_w\[0\] 0.19fF
C1843 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[16\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[18\].delay_unit/mid 0.13fF
C1844 sample_p_2 edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.signal_w\[2\] 0.13fF
C1845 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[16\] clkgen.delay_155ns_2.genblk1\[4\].dly_binary.bypass_in 0.14fF
C1846 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[16\] clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[16\] 0.31fF
C1847 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[8\].delay_unit/mid edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit/mid 0.10fF
C1848 sample_n_out enable_dlycontrol_in 0.45fF
C1849 clkgen.delay_155ns_3.genblk1\[1\].dly_binary.bypass_in clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit/mid 0.12fF
C1850 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.bypass_in edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[21\] 0.11fF
C1851 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.genblk1\[1\].delay_unit/mid clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[0\] 0.13fF
C1852 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit/mid edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[7\] 0.19fF
C1853 clkgen.delay_155ns_2.genblk1\[1\].dly_binary.signal_w\[0\] clkgen.delay_155ns_1.genblk1\[3\].dly_binary.bypass_in 0.10fF
C1854 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[12\] edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit/mid 0.33fF
C1855 VDD clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[16\] 4.64fF
C1856 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[0\] dlycontrol4_in[5] 5.25fF
C1857 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.bypass_in start_conv_in 0.23fF
C1858 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[0\] dlycontrol4_in[3] 0.67fF
C1859 clkgen.delay_155ns_3.genblk1\[0\].dly_binary.in ndecision_finish_in 1.89fF
C1860 clkgen.delay_155ns_2.genblk1\[1\].dly_binary.bypass_in clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit/mid 0.16fF
C1861 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[10\].delay_unit/mid edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[12\].delay_unit/mid 0.10fF
C1862 clkgen.clk_dig_out ndecision_finish_in 0.53fF
C1863 dlycontrol4_in[2] dlycontrol3_in[1] 0.12fF
C1864 VDD edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit/mid 0.26fF
C1865 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit/mid clkgen.clk_comp_out 0.13fF
C1866 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[8\] clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit/a_1632_71# 0.13fF
C1867 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[6\] clkgen.delay_155ns_3.enable_dlycontrol_w 0.12fF
C1868 clkgen.delay_155ns_1.genblk1\[0\].dly_binary.genblk1\[0\].delay_unit/mid clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[16\] 0.10fF
C1869 dlycontrol2_in[3] clkgen.delay_155ns_3.genblk1\[2\].dly_binary.signal_w\[4\] 1.29fF
C1870 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.out clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[16\] 0.16fF
C1871 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit/mid clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[2\] 0.13fF
C1872 clk_dig_out enable_dlycontrol_in 0.71fF
C1873 clkgen.delay_155ns_1.genblk1\[1\].dly_binary.out dlycontrol1_in[3] 0.20fF
C1874 clkgen.delay_155ns_1.genblk1\[1\].dly_binary.out clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[1\] 0.77fF
C1875 clkgen.delay_155ns_2.bypass_enable_w\[4\] clkgen.delay_155ns_2.enable_dlycontrol_w 0.22fF
C1876 clkgen.delay_155ns_1.genblk1\[1\].dly_binary.signal_w\[0\] clkgen.delay_155ns_1.genblk1\[1\].dly_binary.signal_w\[2\] 0.16fF
C1877 ena_in start_conv_in 0.52fF
C1878 nsample_p_in edgedetect.dly_315ns_1.enable_dlycontrol_w 0.29fF
C1879 clkgen.delay_155ns_1.genblk1\[0\].dly_binary.in clkgen.delay_155ns_3.genblk1\[4\].dly_binary.bypass_in 0.47fF
C1880 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[10\] clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit/mid 0.15fF
C1881 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[10\].delay_unit/mid clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[9\] 0.11fF
C1882 clkgen.delay_155ns_2.genblk1\[0\].dly_binary.bypass_in clkgen.delay_155ns_1.genblk1\[2\].dly_binary.bypass_in 0.11fF
C1883 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.bypass_in clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[6\] 0.18fF
C1884 clkgen.delay_155ns_2.genblk1\[1\].dly_binary.bypass_in clkgen.delay_155ns_2.bypass_enable_w\[2\] 0.13fF
C1885 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit/mid clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[15\] 0.11fF
C1886 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.out VDD 1.57fF
C1887 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.bypass_in clkgen.delay_155ns_3.genblk1\[2\].dly_binary.out 1.71fF
C1888 VDD sample_p_in 5.66fF
C1889 clkgen.delay_155ns_1.genblk1\[1\].dly_binary.out clkgen.clk_comp_out 0.83fF
C1890 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.bypass_in dlycontrol3_in[1] 0.12fF
C1891 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.bypass_in enable_dlycontrol_in 1.40fF
C1892 clkgen.clk_dig_out clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[14\] 0.16fF
C1893 clkgen.delay_155ns_2.genblk1\[0\].dly_binary.signal_w\[0\] sample_n_out 0.43fF
C1894 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.bypass_in edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[13\] 0.34fF
C1895 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[2\].delay_unit/a_1632_71# clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[3\] 0.14fF
C1896 clkgen.clk_comp_out clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[16\] 0.88fF
C1897 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.bypass_in clkgen.delay_155ns_2.genblk1\[4\].dly_binary.bypass_in 0.25fF
C1898 dlycontrol2_in[0] clkgen.delay_155ns_1.genblk1\[1\].dly_binary.signal_w\[0\] 0.53fF
C1899 edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.bypass_in edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[20\].delay_unit/mid 0.11fF
C1900 edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.bypass_in clkgen.delay_155ns_3.genblk1\[0\].dly_binary.bypass_in 0.23fF
C1901 clkgen.clk_dig_out clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[8\] 0.32fF
C1902 nsample_p_4 dlycontrol4_in[3] 0.49fF
C1903 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[16\] clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit/mid 0.13fF
C1904 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[8\] edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[6\] 0.18fF
C1905 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[0\].delay_unit/a_1632_71# clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[1\] 0.13fF
C1906 ena_in enable_dlycontrol_in 0.48fF
C1907 edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.genblk1\[0\].delay_unit/mid edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.out 0.12fF
C1908 clkgen.delay_155ns_3.genblk1\[0\].dly_binary.genblk1\[0\].delay_unit/mid sample_p_in 0.23fF
C1909 clkgen.delay_155ns_3.genblk1\[2\].dly_binary.bypass_in clkgen.delay_155ns_3.genblk1\[2\].dly_binary.signal_w\[4\] 0.18fF
C1910 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[10\].delay_unit/mid dlycontrol2_in[3] 0.17fF
C1911 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[0\].delay_unit/mid clkgen.delay_155ns_1.genblk1\[0\].dly_binary.out 0.13fF
C1912 edgedetect.dly_315ns_1.bypass_enable_w\[1\] edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.bypass_in 0.76fF
C1913 clkgen.delay_155ns_3.genblk1\[1\].dly_binary.bypass_in dlycontrol3_in[0] 0.44fF
C1914 clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[4\] dlycontrol1_in[1] 1.92fF
C1915 clkgen.delay_155ns_3.genblk1\[1\].dly_binary.signal_w\[2\] clkgen.delay_155ns_3.genblk1\[0\].dly_binary.bypass_in 0.73fF
C1916 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit/mid VDD 0.39fF
C1917 clkgen.delay_155ns_2.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit/mid VDD 0.36fF
C1918 edgedetect.dly_315ns_1.enable_dlycontrol_w start_conv_in 0.15fF
C1919 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[7\] clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[6\] 0.12fF
C1920 dlycontrol3_in[4] dlycontrol1_in[4] 0.54fF
C1921 sample_p_in edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.bypass_in 0.11fF
C1922 clkgen.delay_155ns_1.genblk1\[0\].dly_binary.in clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[0\] 0.73fF
C1923 dlycontrol2_in[1] clkgen.delay_155ns_3.genblk1\[0\].dly_binary.bypass_in 0.28fF
C1924 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.out dlycontrol4_in[3] 0.12fF
C1925 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[5\] clkgen.delay_155ns_3.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit/mid 0.15fF
C1926 sample_p_2 edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[0\] 0.14fF
C1927 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit/mid VDD 0.34fF
C1928 sample_p_2 edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.out 0.14fF
C1929 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.out edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[10\].delay_unit/mid 0.10fF
C1930 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.bypass_in clkgen.delay_155ns_1.genblk1\[1\].dly_binary.genblk1\[0\].delay_unit/mid 0.13fF
C1931 VDD clkgen.delay_155ns_3.genblk1\[2\].dly_binary.out 1.41fF
C1932 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[4\] ndecision_finish_in 0.13fF
C1933 edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.genblk1\[0\].delay_unit/mid edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[1\] 0.19fF
C1934 clkgen.delay_155ns_2.enable_dlycontrol_w clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit/mid 0.10fF
C1935 clkgen.clk_dig_out clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[6\] 0.11fF
C1936 VDD dlycontrol3_in[1] 3.74fF
C1937 VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[15\] 0.75fF
C1938 VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[6\].delay_unit/mid 0.71fF
C1939 clkgen.delay_155ns_3.genblk1\[0\].dly_binary.out VDD 0.94fF
C1940 edgedetect.start_conv_edge_w dlycontrol1_in[2] 1.66fF
C1941 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[5\].delay_unit/mid edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[5\] 0.11fF
C1942 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[13\] clkgen.delay_155ns_2.genblk1\[4\].dly_binary.bypass_in 0.14fF
C1943 clkgen.delay_155ns_2.genblk1\[0\].dly_binary.genblk1\[0\].delay_unit/mid VDD 0.30fF
C1944 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit/mid dlycontrol2_in[3] 0.16fF
C1945 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit/mid clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[2\] 0.17fF
C1946 dlycontrol4_in[5] dlycontrol4_in[3] 0.28fF
C1947 VDD edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.genblk1\[0\].delay_unit/mid 0.37fF
C1948 clkgen.delay_155ns_1.enable_dlycontrol_w clkgen.delay_155ns_1.bypass_enable_w\[1\] 0.10fF
C1949 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.out edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.signal_w\[0\] 4.08fF
C1950 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[4\] VDD 0.69fF
C1951 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit/mid VDD 0.39fF
C1952 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[5\] sample_p_out 0.49fF
C1953 ndecision_finish_in clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[13\] 0.29fF
C1954 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit/mid VDD 0.19fF
C1955 edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[1\] edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[1\] 0.21fF
C1956 VDD dlycontrol2_in[2] 4.17fF
C1957 dlycontrol3_in[2] dlycontrol3_in[3] 1.21fF
C1958 edgedetect.dly_315ns_1.enable_dlycontrol_w enable_dlycontrol_in 0.13fF
C1959 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[0\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[0\] 0.10fF
C1960 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit/a_1632_71# edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[6\] 0.13fF
C1961 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[5\] clkgen.delay_155ns_3.bypass_enable_w\[3\] 0.16fF
C1962 clkgen.delay_155ns_2.bypass_enable_w\[3\] VDD 0.28fF
C1963 sample_n_1 clkgen.delay_155ns_1.genblk1\[1\].dly_binary.signal_w\[1\] 0.17fF
C1964 clkgen.delay_155ns_2.bypass_enable_w\[4\] clkgen.delay_155ns_2.bypass_enable_w\[1\] 0.41fF
C1965 clkgen.delay_155ns_3.genblk1\[0\].dly_binary.genblk1\[0\].delay_unit/mid dlycontrol3_in[1] 0.15fF
C1966 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[4\] clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[0\] 0.14fF
C1967 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[0\] clkgen.delay_155ns_1.genblk1\[0\].dly_binary.bypass_in 0.11fF
C1968 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.bypass_in edgedetect.dly_315ns_1.enable_dlycontrol_w 0.52fF
C1969 VDD edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[1\] 0.93fF
C1970 edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.bypass_in edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[22\] 0.16fF
C1971 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.out clkgen.delay_155ns_2.genblk1\[3\].dly_binary.bypass_in 0.37fF
C1972 clkgen.delay_155ns_3.genblk1\[2\].dly_binary.signal_w\[3\] VDD 0.87fF
C1973 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[0\].delay_unit/mid VDD 0.26fF
C1974 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[15\].delay_unit/mid edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[15\] 0.16fF
C1975 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[3\] clkgen.delay_155ns_1.genblk1\[0\].dly_binary.bypass_in 0.17fF
C1976 ndecision_finish_in clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit/mid 0.12fF
C1977 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[16\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[19\].delay_unit/mid 0.14fF
C1978 VDD edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit/mid 0.27fF
C1979 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[8\] clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit/mid 0.11fF
C1980 clkgen.delay_155ns_2.genblk1\[1\].dly_binary.signal_w\[2\] clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[16\] 1.37fF
C1981 clkgen.clk_dig_delayed_w clkgen.delay_155ns_1.genblk1\[0\].dly_binary.bypass_in 0.16fF
C1982 sample_p_in edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.signal_w\[2\] 0.10fF
C1983 clkgen.delay_155ns_1.genblk1\[0\].dly_binary.out clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit/mid 0.12fF
C1984 dlycontrol2_in[0] clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[8\] 0.17fF
C1985 clkgen.delay_155ns_1.genblk1\[0\].dly_binary.signal_w\[0\] VDD 0.87fF
C1986 dlycontrol1_in[2] clkgen.delay_155ns_1.genblk1\[1\].dly_binary.out 0.10fF
C1987 sample_p_2 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[8\] 0.46fF
C1988 clkgen.delay_155ns_1.genblk1\[2\].dly_binary.genblk1\[0\].delay_unit/mid VDD 0.35fF
C1989 clkgen.delay_155ns_2.enable_dlycontrol_w clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit/mid 0.17fF
C1990 clkgen.delay_155ns_1.genblk1\[1\].dly_binary.bypass_in clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[16\] 0.16fF
C1991 edgedetect.start_conv_edge_w clkgen.delay_155ns_3.enable_dlycontrol_w 0.12fF
C1992 clkgen.enable_loop_in VDD 0.90fF
C1993 VDD clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[2\] 0.89fF
C1994 clkgen.delay_155ns_2.genblk1\[0\].dly_binary.bypass_in enable_dlycontrol_in 2.20fF
C1995 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[11\].delay_unit/mid VDD 0.45fF
C1996 dlycontrol2_in[0] clkgen.delay_155ns_2.genblk1\[1\].dly_binary.signal_w\[0\] 0.13fF
C1997 edgedetect.start_conv_edge_w edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.in 1.30fF
C1998 nsample_n_in nsample_n_1 0.59fF
C1999 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[0\] clkgen.delay_155ns_3.genblk1\[1\].dly_binary.bypass_in 0.12fF
C2000 edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.signal_w\[0\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[1\].delay_unit/mid 0.13fF
C2001 edgedetect.dly_315ns_1.enable_dlycontrol_w edgedetect.dly_315ns_1.bypass_enable_w\[5\] 0.26fF
C2002 edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.out sample_p_out 0.12fF
C2003 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit/mid clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit/mid 0.11fF
C2004 clkgen.delay_155ns_3.genblk1\[0\].dly_binary.in clkgen.delay_155ns_1.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit/mid 0.12fF
C2005 clkgen.delay_155ns_2.genblk1\[1\].dly_binary.signal_w\[1\] VDD 0.74fF
C2006 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.out edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[6\] 0.37fF
C2007 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit/mid clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[9\] 0.12fF
C2008 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit/a_1691_329# VDD 0.10fF
C2009 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[0\].delay_unit/mid edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.bypass_in 0.14fF
C2010 edgedetect.dly_315ns_1.bypass_enable_w\[3\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[19\] 0.23fF
C2011 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[0\].delay_unit/mid edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[1\] 0.17fF
C2012 clkgen.delay_155ns_1.genblk1\[2\].dly_binary.genblk1\[0\].delay_unit/mid clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[1\] 0.13fF
C2013 clkgen.delay_155ns_2.genblk1\[0\].dly_binary.bypass_in clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[0\] 4.18fF
C2014 VDD clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[6\] 1.00fF
C2015 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.bypass_in edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit/mid 0.15fF
C2016 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.out edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit/mid 0.21fF
C2017 clkgen.delay_155ns_1.genblk1\[0\].dly_binary.in clkgen.delay_155ns_1.genblk1\[1\].dly_binary.signal_w\[1\] 0.15fF
C2018 nsample_p_3 VDD 0.19fF
C2019 edgedetect.ena_in clkgen.delay_155ns_1.bypass_enable_w\[3\] 0.16fF
C2020 enable_dlycontrol_in clkgen.delay_155ns_1.bypass_enable_w\[1\] 0.86fF
C2021 edgedetect.start_conv_edge_w clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[0\] 1.27fF
C2022 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[0\] edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.out 0.14fF
C2023 edgedetect.start_conv_edge_w sample_n_in 0.16fF
C2024 dlycontrol2_in[0] clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[4\] 1.06fF
C2025 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit/mid VDD 0.37fF
C2026 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[0\].delay_unit/mid VDD 0.41fF
C2027 VDD clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[14\] 0.83fF
C2028 clkgen.delay_155ns_1.genblk1\[0\].dly_binary.bypass_in clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[16\] 1.93fF
C2029 clkgen.clk_dig_delayed_w clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[0\] 0.26fF
C2030 edgedetect.start_conv_edge_w clkgen.delay_155ns_1.genblk1\[3\].dly_binary.bypass_in 0.49fF
C2031 clkgen.clk_dig_out sample_n_4 0.28fF
C2032 clkgen.delay_155ns_2.genblk1\[0\].dly_binary.signal_w\[0\] sample_n_3 0.17fF
C2033 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit/a_1632_71# edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[15\] 0.13fF
C2034 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[1\] clkgen.delay_155ns_3.genblk1\[1\].dly_binary.bypass_in 0.60fF
C2035 edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[4\] edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.bypass_in 0.80fF
C2036 clkgen.delay_155ns_2.bypass_enable_w\[4\] clkgen.delay_155ns_2.bypass_enable_w\[2\] 0.28fF
C2037 edgedetect.ena_in clkgen.delay_155ns_2.genblk1\[0\].dly_binary.out 1.14fF
C2038 edgedetect.start_conv_edge_w clkgen.delay_155ns_2.genblk1\[1\].dly_binary.bypass_in 0.41fF
C2039 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[10\].delay_unit/a_1632_71# clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[11\] 0.13fF
C2040 VDD clkgen.delay_155ns_1.genblk1\[1\].dly_binary.out_mux/a_505_21# 0.11fF
C2041 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit/mid clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[16\] 0.11fF
C2042 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.bypass_in dlycontrol3_in[4] 0.18fF
C2043 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[11\] clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[12\] 0.22fF
C2044 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.bypass_in clkgen.delay_155ns_2.genblk1\[4\].dly_binary.bypass_in 0.54fF
C2045 edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.bypass_in nsample_p_in 0.11fF
C2046 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.bypass_in start_conv_in 0.87fF
C2047 clkgen.delay_155ns_2.genblk1\[0\].dly_binary.bypass_in clkgen.delay_155ns_2.genblk1\[0\].dly_binary.signal_w\[0\] 0.36fF
C2048 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit/mid VDD 0.42fF
C2049 clkgen.delay_155ns_2.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit/mid clkgen.delay_155ns_2.genblk1\[1\].dly_binary.signal_w\[2\] 0.10fF
C2050 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[0\] edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[1\] 0.13fF
C2051 clkgen.delay_155ns_3.genblk1\[1\].dly_binary.out dlycontrol2_in[4] 1.16fF
C2052 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[0\].delay_unit/mid edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[1\] 0.12fF
C2053 edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.bypass_in edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[18\].delay_unit/mid 0.10fF
C2054 VDD edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit/mid 0.39fF
C2055 clkgen.delay_155ns_2.genblk1\[1\].dly_binary.out clkgen.delay_155ns_2.genblk1\[2\].dly_binary.genblk1\[0\].delay_unit/mid 0.14fF
C2056 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.bypass_in clkgen.delay_155ns_1.genblk1\[4\].dly_binary.out 0.81fF
C2057 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.in edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit/mid 0.15fF
C2058 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[8\] clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[0\] 0.10fF
C2059 nsample_p_3 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.bypass_in 0.44fF
C2060 ena_in clkgen.delay_155ns_1.genblk1\[3\].dly_binary.out 1.47fF
C2061 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[0\] VDD 0.74fF
C2062 clkgen.delay_155ns_1.genblk1\[1\].dly_binary.out clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[0\] 0.13fF
C2063 VDD clk_dig_out 2.26fF
C2064 sample_p_in edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.out 0.23fF
C2065 clkgen.delay_155ns_1.genblk1\[1\].dly_binary.out clkgen.delay_155ns_1.genblk1\[3\].dly_binary.bypass_in 0.50fF
C2066 clkgen.delay_155ns_1.genblk1\[0\].dly_binary.in clkgen.delay_155ns_3.genblk1\[3\].dly_binary.out 0.60fF
C2067 VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[27\] 1.08fF
C2068 clkgen.clk_dig_out clkgen.delay_155ns_1.genblk1\[2\].dly_binary.bypass_in 1.15fF
C2069 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[9\].delay_unit/mid VDD 0.38fF
C2070 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[28\].delay_unit/mid start_conv_in 0.12fF
C2071 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[16\] edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.bypass_in 0.53fF
C2072 dlycontrol4_in[2] edgedetect.dly_315ns_1.enable_dlycontrol_w 0.84fF
C2073 clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[0\] clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[16\] 1.05fF
C2074 VDD clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[4\] 0.73fF
C2075 clkgen.delay_155ns_2.bypass_enable_w\[0\] clkgen.delay_155ns_1.genblk1\[4\].dly_binary.out 0.12fF
C2076 VDD clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit/mid 0.31fF
C2077 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.out clkgen.delay_155ns_3.genblk1\[2\].dly_binary.signal_w\[4\] 0.52fF
C2078 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[0\] clk_dig_out 3.78fF
C2079 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[16\] clkgen.delay_155ns_2.genblk1\[4\].dly_binary.bypass_in 1.54fF
C2080 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.bypass_in clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[16\] 0.13fF
C2081 edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.bypass_in start_conv_in 0.10fF
C2082 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.out clkgen.delay_155ns_3.genblk1\[1\].dly_binary.bypass_in 0.10fF
C2083 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[13\] VDD 0.77fF
C2084 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit/mid clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[13\] 0.14fF
C2085 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[0\].delay_unit/mid clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[1\] 0.13fF
C2086 clkgen.delay_155ns_2.genblk1\[1\].dly_binary.bypass_in clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[16\] 1.67fF
C2087 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.bypass_in VDD 6.64fF
C2088 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[4\].delay_unit/mid VDD 0.28fF
C2089 start_conv_in clkgen.delay_155ns_3.genblk1\[2\].dly_binary.bypass_in 0.16fF
C2090 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[4\] dlycontrol1_in[2] 0.19fF
C2091 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[16\] dlycontrol2_in[2] 1.55fF
C2092 dlycontrol3_in[4] edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.signal_w\[1\] 0.23fF
C2093 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit/a_1632_71# clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[16\] 0.14fF
C2094 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[14\].delay_unit/mid edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[15\] 0.14fF
C2095 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[7\] clkgen.delay_155ns_1.genblk1\[2\].dly_binary.bypass_in 0.11fF
C2096 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[0\] edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.bypass_in 0.14fF
C2097 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.bypass_in edgedetect.dly_315ns_1.enable_dlycontrol_w 0.62fF
C2098 ena_in VDD 2.47fF
C2099 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[16\] edgedetect.dly_315ns_1.bypass_enable_w\[4\] 0.62fF
C2100 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.out VDD 2.87fF
C2101 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit/mid clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[9\] 0.13fF
C2102 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit/mid dlycontrol2_in[2] 0.15fF
C2103 dlycontrol3_in[0] dlycontrol3_in[1] 1.17fF
C2104 clkgen.delay_155ns_3.genblk1\[0\].dly_binary.out dlycontrol3_in[0] 0.45fF
C2105 clkgen.delay_155ns_3.genblk1\[1\].dly_binary.out clkgen.delay_155ns_3.genblk1\[2\].dly_binary.bypass_in 0.89fF
C2106 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.out clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[16\] 0.69fF
C2107 VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[7\].delay_unit/mid 0.37fF
C2108 clkgen.delay_155ns_3.genblk1\[1\].dly_binary.signal_w\[2\] clkgen.delay_155ns_3.genblk1\[0\].dly_binary.signal_w\[1\] 0.21fF
C2109 VDD clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[3\] 0.72fF
C2110 VDD clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[0\] 0.57fF
C2111 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[0\] clkgen.delay_155ns_3.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit/mid 0.11fF
C2112 dlycontrol3_in[0] dlycontrol2_in[2] 0.84fF
C2113 dlycontrol2_in[1] clkgen.delay_155ns_3.genblk1\[1\].dly_binary.bypass_in 0.14fF
C2114 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.bypass_in edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.bypass_in 4.54fF
C2115 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit/mid clkgen.delay_155ns_3.genblk1\[2\].dly_binary.bypass_in 0.11fF
C2116 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit/a_1691_329# VDD 0.12fF
C2117 clkgen.delay_155ns_2.genblk1\[1\].dly_binary.out ndecision_finish_in 1.40fF
C2118 dlycontrol1_in[2] clkgen.delay_155ns_1.genblk1\[2\].dly_binary.genblk1\[0\].delay_unit/mid 0.19fF
C2119 clkgen.delay_155ns_2.genblk1\[1\].dly_binary.signal_w\[1\] clkgen.delay_155ns_2.genblk1\[1\].dly_binary.signal_w\[2\] 1.05fF
C2120 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[8\] clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[10\] 0.15fF
C2121 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[5\] dlycontrol2_in[0] 0.13fF
C2122 ena_in dlycontrol1_in[3] 0.26fF
C2123 VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[14\] 0.57fF
C2124 clkgen.clk_dig_delayed_w clkgen.delay_155ns_1.genblk1\[0\].dly_binary.out 0.51fF
C2125 clkgen.delay_155ns_3.genblk1\[2\].dly_binary.signal_w\[0\] clkgen.delay_155ns_3.genblk1\[2\].dly_binary.bypass_in 0.17fF
C2126 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.out clkgen.delay_155ns_3.genblk1\[1\].dly_binary.genblk1\[0\].delay_unit/mid 0.16fF
C2127 dlycontrol4_in[1] edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit/mid 0.15fF
C2128 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[27\].delay_unit/mid edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[25\] 0.19fF
C2129 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.in dlycontrol3_in[1] 0.12fF
C2130 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[8\] dlycontrol3_in[2] 2.31fF
C2131 sample_p_3 VDD 1.16fF
C2132 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[7\] dlycontrol2_in[4] 0.14fF
C2133 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[22\].delay_unit/mid VDD 0.29fF
C2134 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.bypass_in edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.signal_w\[1\] 0.22fF
C2135 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit/a_1632_71# edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[8\] 0.13fF
C2136 clkgen.delay_155ns_2.genblk1\[0\].dly_binary.bypass_in clkgen.delay_155ns_1.genblk1\[3\].dly_binary.out 4.87fF
C2137 clkgen.clk_dig_out clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[16\] 0.54fF
C2138 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[8\].delay_unit/mid VDD 0.27fF
C2139 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit/mid VDD 0.38fF
C2140 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit/a_1632_71# edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[9\] 0.14fF
C2141 clkgen.delay_155ns_3.genblk1\[0\].dly_binary.in dlycontrol3_in[4] 0.52fF
C2142 clkgen.clk_dig_delayed_w clkgen.delay_155ns_1.genblk1\[1\].dly_binary.signal_w\[2\] 0.71fF
C2143 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[2\] edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit/mid 0.21fF
C2144 clkgen.clk_dig_out dlycontrol3_in[4] 0.17fF
C2145 clkgen.delay_155ns_1.genblk1\[0\].dly_binary.signal_w\[0\] clkgen.delay_155ns_1.genblk1\[0\].dly_binary.bypass_in 0.10fF
C2146 VDD edgedetect.dly_315ns_1.enable_dlycontrol_w 2.04fF
C2147 clkgen.delay_155ns_3.genblk1\[0\].dly_binary.genblk1\[0\].delay_unit/a_1632_71# clkgen.delay_155ns_3.genblk1\[0\].dly_binary.signal_w\[1\] 0.13fF
C2148 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[8\] clkgen.delay_155ns_1.genblk1\[2\].dly_binary.out 0.47fF
C2149 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[16\] dlycontrol1_in[4] 2.55fF
C2150 nsample_p_1 VDD 0.36fF
C2151 start_conv_in clkgen.delay_155ns_3.genblk1\[3\].dly_binary.bypass_in 0.62fF
C2152 clkgen.delay_155ns_3.genblk1\[2\].dly_binary.genblk1\[1\].delay_unit/mid clkgen.delay_155ns_3.genblk1\[0\].dly_binary.signal_w\[0\] 0.11fF
C2153 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.out clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[8\] 0.10fF
C2154 VDD edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[3\] 0.61fF
C2155 VDD dlycontrol1_in[4] 3.26fF
C2156 clkgen.delay_155ns_3.genblk1\[2\].dly_binary.signal_w\[2\] VDD 0.74fF
C2157 clkgen.delay_155ns_2.bypass_enable_w\[0\] clkgen.delay_155ns_2.genblk1\[0\].dly_binary.bypass_in 0.33fF
C2158 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit/mid clkgen.delay_155ns_3.genblk1\[0\].dly_binary.bypass_in 0.12fF
C2159 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[6\] clkgen.delay_155ns_1.genblk1\[2\].dly_binary.bypass_in 0.13fF
C2160 edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.bypass_in edgedetect.dly_315ns_1.bypass_enable_w\[5\] 0.18fF
C2161 VDD clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit/mid 0.25fF
C2162 clkgen.clk_dig_delayed_w clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[1\] 0.24fF
C2163 clkgen.delay_155ns_1.bypass_enable_w\[4\] dlycontrol1_in[4] 0.24fF
C2164 clkgen.delay_155ns_3.genblk1\[0\].dly_binary.in clkgen.delay_155ns_3.genblk1\[1\].dly_binary.out 0.25fF
C2165 clkgen.delay_155ns_1.genblk1\[1\].dly_binary.bypass_in sample_n_out 0.11fF
C2166 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[5\] VDD 0.67fF
C2167 sample_n_3 VDD 0.35fF
C2168 edgedetect.start_conv_edge_w edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[8\] 0.14fF
C2169 dlycontrol4_in[2] dlycontrol2_in[4] 1.29fF
C2170 dlycontrol1_in[3] dlycontrol1_in[4] 0.73fF
C2171 clkgen.delay_155ns_2.genblk1\[1\].dly_binary.bypass_in dlycontrol2_in[2] 1.07fF
C2172 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[2\].delay_unit/mid clkgen.delay_155ns_3.genblk1\[2\].dly_binary.bypass_in 0.15fF
C2173 clkgen.delay_155ns_2.genblk1\[0\].dly_binary.bypass_in clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[16\] 0.19fF
C2174 VDD edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[13\].delay_unit/mid 0.22fF
C2175 clkgen.clk_dig_out enable_dlycontrol_in 0.72fF
C2176 clkgen.delay_155ns_1.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit/mid VSS 1.27fF
C2177 clkgen.delay_155ns_3.genblk1\[1\].dly_binary.genblk1\[0\].delay_unit/mid VSS 1.31fF
C2178 edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[2\] VSS 2.04fF
C2179 edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[3\] VSS 1.24fF
C2180 edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit/mid VSS 1.31fF
C2181 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit/mid VSS 1.20fF
C2182 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[26\] VSS 1.09fF
C2183 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[27\] VSS 1.46fF
C2184 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[26\].delay_unit/mid VSS 1.27fF
C2185 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit/mid VSS 1.25fF
C2186 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[21\] VSS 1.43fF
C2187 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[22\] VSS 1.18fF
C2188 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[21\].delay_unit/mid VSS 1.28fF
C2189 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[19\].delay_unit/mid VSS 1.27fF
C2190 clkgen.delay_155ns_3.genblk1\[2\].dly_binary.signal_w\[1\] VSS 1.08fF
C2191 clkgen.delay_155ns_3.genblk1\[2\].dly_binary.genblk1\[0\].delay_unit/mid VSS 1.33fF
C2192 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[4\] VSS 1.13fF
C2193 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[5\] VSS 1.16fF
C2194 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit/mid VSS 1.23fF
C2195 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[8\] VSS 1.05fF
C2196 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[9\] VSS 1.17fF
C2197 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit/mid VSS 1.50fF
C2198 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[3\] VSS 1.25fF
C2199 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit/mid VSS 1.33fF
C2200 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[15\] VSS 1.14fF
C2201 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit/mid VSS 1.24fF
C2202 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[14\] VSS 1.02fF
C2203 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[15\] VSS 2.42fF
C2204 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit/mid VSS 1.29fF
C2205 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[14\] VSS 1.36fF
C2206 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[15\] VSS 1.09fF
C2207 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[14\].delay_unit/mid VSS 1.42fF
C2208 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit/mid VSS 1.40fF
C2209 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[10\] VSS 1.14fF
C2210 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[11\] VSS 1.23fF
C2211 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[10\].delay_unit/mid VSS 1.24fF
C2212 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[6\] VSS 1.12fF
C2213 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit/mid VSS 1.28fF
C2214 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[9\] VSS 1.06fF
C2215 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[10\] VSS 1.05fF
C2216 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit/mid VSS 1.30fF
C2217 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[7\] VSS 2.04fF
C2218 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[8\] VSS 1.43fF
C2219 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit/mid VSS 1.26fF
C2220 dlycontrol3_in[1] VSS 2.84fF
C2221 dlycontrol3_in[3] VSS 1.87fF
C2222 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[0\].delay_unit/mid VSS 1.23fF
C2223 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[4\] VSS 1.25fF
C2224 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit/mid VSS 1.32fF
C2225 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[3\] VSS 1.50fF
C2226 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[2\].delay_unit/mid VSS 1.19fF
C2227 nsample_n_out VSS 0.61fF
C2228 outbuf_6/a_27_47# VSS 0.62fF
C2229 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[11\] VSS 1.26fF
C2230 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit/mid VSS 1.53fF
C2231 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[6\] VSS 1.28fF
C2232 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit/mid VSS 1.41fF
C2233 dlycontrol4_in[3] VSS 2.98fF
C2234 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[7\].delay_unit/mid VSS 1.15fF
C2235 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.bypass_in VSS 0.90fF
C2236 clkgen.delay_155ns_3.bypass_enable_w\[3\] VSS 0.30fF
C2237 clkgen.delay_155ns_3.genblk1\[3\].bypass_enable/a_59_75# VSS 0.24fF $ **FLOATING
C2238 clkgen.delay_155ns_2.bypass_enable_w\[2\] VSS 0.44fF
C2239 clkgen.delay_155ns_2.genblk1\[2\].bypass_enable/a_59_75# VSS 0.26fF $ **FLOATING
C2240 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[1\] VSS 1.24fF
C2241 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[0\].delay_unit/mid VSS 1.25fF
C2242 clkgen.delay_155ns_1.bypass_enable_w\[1\] VSS 3.25fF
C2243 clkgen.delay_155ns_1.genblk1\[1\].bypass_enable/a_59_75# VSS 0.23fF $ **FLOATING
C2244 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[3\] VSS 1.18fF
C2245 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[2\].delay_unit/mid VSS 1.32fF
C2246 nsample_p_out VSS 0.36fF
C2247 outbuf_5/a_27_47# VSS 0.53fF
C2248 edgedetect.dly_315ns_1.bypass_enable_w\[0\] VSS 0.69fF
C2249 edgedetect.dly_315ns_1.genblk1\[0\].bypass_enable/a_59_75# VSS 0.24fF $ **FLOATING
C2250 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[13\] VSS 1.33fF
C2251 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[14\] VSS 1.62fF
C2252 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit/mid VSS 1.27fF
C2253 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[16\] VSS 3.68fF
C2254 edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.signal_w\[2\] VSS 0.51fF
C2255 edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit/mid VSS 1.25fF
C2256 dlycontrol2_in[2] VSS 3.49fF
C2257 clkgen.delay_155ns_3.enable_dlycontrol_w VSS 1.40fF
C2258 enable_dlycontrol_in VSS 4.96fF
C2259 clkgen.delay_155ns_3.enablebuffer/a_27_47# VSS 0.50fF
C2260 sample_n_out VSS 0.18fF
C2261 outbuf_4/a_27_47# VSS 0.52fF
C2262 clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[3\] VSS 1.30fF
C2263 clkgen.delay_155ns_1.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit/mid VSS 1.24fF
C2264 clkgen.clk_comp_out VSS 1.06fF
C2265 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.out_mux/a_505_21# VSS 0.25fF
C2266 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.out_mux/a_76_199# VSS 0.17fF $ **FLOATING
C2267 edgedetect.dly_315ns_1.bypass_enable_w\[5\] VSS 1.33fF
C2268 edgedetect.dly_315ns_1.genblk1\[5\].bypass_enable/a_59_75# VSS 0.23fF $ **FLOATING
C2269 clkgen.delay_155ns_3.genblk1\[2\].dly_binary.signal_w\[4\] VSS 2.55fF
C2270 clkgen.delay_155ns_3.genblk1\[2\].dly_binary.bypass_in VSS 2.04fF
C2271 clkgen.delay_155ns_3.genblk1\[2\].dly_binary.out VSS 0.81fF
C2272 clkgen.delay_155ns_3.genblk1\[2\].dly_binary.out_mux/a_505_21# VSS 0.25fF
C2273 clkgen.delay_155ns_3.genblk1\[2\].dly_binary.out_mux/a_76_199# VSS 0.18fF $ **FLOATING
C2274 clkgen.delay_155ns_3.genblk1\[0\].dly_binary.signal_w\[1\] VSS 0.50fF
C2275 clkgen.delay_155ns_3.genblk1\[0\].dly_binary.bypass_in VSS 1.26fF
C2276 clkgen.delay_155ns_3.genblk1\[0\].dly_binary.out_mux/a_505_21# VSS 0.23fF
C2277 clkgen.delay_155ns_3.genblk1\[0\].dly_binary.out_mux/a_76_199# VSS 0.18fF $ **FLOATING
C2278 sample_p_out VSS 0.30fF
C2279 sample_p_4 VSS 0.72fF
C2280 outbuf_3/a_27_47# VSS 0.51fF
C2281 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit/mid VSS 1.22fF
C2282 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit/mid VSS 1.32fF
C2283 edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.genblk1\[1\].delay_unit/mid VSS 1.21fF
C2284 clk_comp_out VSS 0.46fF
C2285 outbuf_2/a_27_47# VSS 0.61fF
C2286 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[2\] VSS 1.42fF
C2287 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[3\] VSS 1.45fF
C2288 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit/mid VSS 1.18fF
C2289 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[25\].delay_unit/mid VSS 1.20fF
C2290 dlycontrol2_in[3] VSS 2.84fF
C2291 clkgen.delay_155ns_1.genblk1\[2\].dly_binary.out VSS 1.86fF
C2292 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[8\] VSS 1.30fF
C2293 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.out_mux/a_505_21# VSS 0.25fF
C2294 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.out_mux/a_76_199# VSS 0.17fF $ **FLOATING
C2295 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[6\] VSS 1.30fF
C2296 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[7\] VSS 1.22fF
C2297 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit/mid VSS 1.32fF
C2298 clkgen.delay_155ns_1.genblk1\[1\].dly_binary.out_mux/a_505_21# VSS 0.24fF
C2299 clkgen.delay_155ns_1.genblk1\[1\].dly_binary.out_mux/a_76_199# VSS 0.17fF $ **FLOATING
C2300 dlycontrol1_in[1] VSS 2.64fF
C2301 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[20\] VSS 1.42fF
C2302 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[20\].delay_unit/mid VSS 1.45fF
C2303 dlycontrol1_in[4] VSS 1.94fF
C2304 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[18\] VSS 1.29fF
C2305 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[19\] VSS 1.00fF
C2306 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[18\].delay_unit/mid VSS 1.27fF
C2307 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit/mid VSS 1.30fF
C2308 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit/a_1691_329# VSS 0.11fF
C2309 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit/mid VSS 1.27fF
C2310 clk_dig_out VSS 1.71fF
C2311 outbuf_1/a_27_47# VSS 0.54fF
C2312 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[1\] VSS 1.20fF
C2313 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[2\] VSS 1.12fF
C2314 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit/a_1691_329# VSS 0.10fF
C2315 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit/mid VSS 1.31fF
C2316 edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.bypass_in VSS 4.54fF
C2317 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[14\] VSS 2.14fF
C2318 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit/mid VSS 1.19fF
C2319 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.and_bypass_switch/a_207_413# VSS 0.18fF $ **FLOATING
C2320 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.and_bypass_switch/a_27_413# VSS 0.18fF $ **FLOATING
C2321 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit/mid VSS 1.27fF
C2322 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[13\].delay_unit/a_1691_329# VSS 0.11fF
C2323 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[13\].delay_unit/mid VSS 1.26fF
C2324 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[3\] VSS 1.41fF
C2325 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[2\].delay_unit/mid VSS 1.27fF
C2326 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[5\] VSS 0.93fF
C2327 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit/mid VSS 1.33fF
C2328 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[32\] VSS 6.07fF
C2329 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.bypass_in VSS 2.51fF
C2330 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.out VSS 4.86fF
C2331 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.out_mux/a_505_21# VSS 0.25fF
C2332 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.out_mux/a_76_199# VSS 0.18fF $ **FLOATING
C2333 start_conv_in VSS 7.11fF
C2334 edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.out VSS 2.49fF
C2335 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[8\] VSS 2.15fF
C2336 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.bypass_in VSS 4.38fF
C2337 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.out_mux/a_505_21# VSS 0.24fF
C2338 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.out_mux/a_76_199# VSS 0.20fF $ **FLOATING
C2339 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit/mid VSS 1.24fF
C2340 edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.out VSS 1.64fF
C2341 edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.out_mux/a_505_21# VSS 0.25fF
C2342 edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.out_mux/a_76_199# VSS 0.17fF $ **FLOATING
C2343 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit/mid VSS 1.25fF
C2344 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit/mid VSS 1.27fF
C2345 clkgen.delay_155ns_3.bypass_enable_w\[0\] VSS 1.24fF
C2346 dlycontrol3_in[0] VSS 3.86fF
C2347 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[2\] VSS 1.31fF
C2348 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit/mid VSS 1.16fF
C2349 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit/mid VSS 1.37fF
C2350 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[9\] VSS 1.03fF
C2351 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit/mid VSS 1.30fF
C2352 sample_p_in VSS 5.14fF
C2353 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.bypass_in VSS 3.30fF
C2354 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.and_bypass_switch/a_207_413# VSS 0.16fF $ **FLOATING
C2355 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.and_bypass_switch/a_27_413# VSS 0.19fF $ **FLOATING
C2356 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.and_bypass_switch/a_207_413# VSS 0.17fF $ **FLOATING
C2357 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.and_bypass_switch/a_27_413# VSS 0.19fF $ **FLOATING
C2358 dlycontrol4_in[5] VSS 1.33fF
C2359 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[10\].delay_unit/mid VSS 1.25fF
C2360 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[4\] VSS 1.07fF
C2361 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[5\] VSS 1.14fF
C2362 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit/mid VSS 1.43fF
C2363 clkgen.delay_155ns_3.bypass_enable_w\[2\] VSS 0.43fF
C2364 clkgen.delay_155ns_3.genblk1\[2\].bypass_enable/a_59_75# VSS 0.26fF $ **FLOATING
C2365 clkgen.delay_155ns_2.genblk1\[1\].bypass_enable/a_59_75# VSS 0.25fF $ **FLOATING
C2366 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.signal_w\[0\] VSS 1.27fF
C2367 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.signal_w\[1\] VSS 0.42fF
C2368 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.genblk1\[0\].delay_unit/mid VSS 1.28fF
C2369 clkgen.delay_155ns_1.genblk1\[0\].dly_binary.bypass_in VSS 1.87fF
C2370 clkgen.delay_155ns_1.bypass_enable_w\[0\] VSS 0.14fF
C2371 clkgen.delay_155ns_1.genblk1\[0\].bypass_enable/a_59_75# VSS 0.28fF $ **FLOATING
C2372 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[6\] VSS 1.03fF
C2373 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[7\] VSS 1.02fF
C2374 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[6\].delay_unit/mid VSS 1.32fF
C2375 dlycontrol4_in[0] VSS 9.33fF
C2376 clkgen.delay_155ns_1.genblk1\[1\].dly_binary.signal_w\[1\] VSS 1.10fF
C2377 clkgen.delay_155ns_1.genblk1\[1\].dly_binary.signal_w\[2\] VSS 0.59fF
C2378 clkgen.delay_155ns_1.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit/mid VSS 1.28fF
C2379 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[1\] VSS 1.10fF
C2380 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[2\] VSS 1.08fF
C2381 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[1\].delay_unit/mid VSS 1.27fF
C2382 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[12\] VSS 1.01fF
C2383 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit/mid VSS 1.30fF
C2384 clkgen.delay_155ns_1.genblk1\[2\].dly_binary.bypass_in VSS 2.91fF
C2385 clkgen.delay_155ns_1.genblk1\[2\].dly_binary.and_bypass_switch/a_207_413# VSS 0.16fF $ **FLOATING
C2386 clkgen.delay_155ns_1.genblk1\[2\].dly_binary.and_bypass_switch/a_27_413# VSS 0.19fF $ **FLOATING
C2387 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.and_bypass_switch/a_207_413# VSS 0.16fF $ **FLOATING
C2388 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.and_bypass_switch/a_27_413# VSS 0.18fF $ **FLOATING
C2389 dlycontrol2_in[4] VSS 1.83fF
C2390 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[0\] VSS 1.28fF
C2391 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.out VSS 0.68fF
C2392 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.bypass_in VSS 1.24fF
C2393 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.and_bypass_switch/a_207_413# VSS 0.17fF $ **FLOATING
C2394 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.and_bypass_switch/a_27_413# VSS 0.18fF $ **FLOATING
C2395 edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.signal_w\[0\] VSS 1.25fF
C2396 edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.signal_w\[1\] VSS 1.11fF
C2397 edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.genblk1\[0\].delay_unit/mid VSS 1.27fF
C2398 clkgen.delay_155ns_2.enable_dlycontrol_w VSS 1.43fF
C2399 clkgen.delay_155ns_2.enablebuffer/a_27_47# VSS 0.53fF
C2400 edgedetect.dly_315ns_1.bypass_enable_w\[4\] VSS 0.96fF
C2401 edgedetect.dly_315ns_1.enable_dlycontrol_w VSS 1.11fF
C2402 edgedetect.dly_315ns_1.genblk1\[4\].bypass_enable/a_59_75# VSS 0.25fF $ **FLOATING
C2403 clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[2\] VSS 1.16fF
C2404 clkgen.delay_155ns_1.genblk1\[2\].dly_binary.genblk1\[1\].delay_unit/mid VSS 1.38fF
C2405 nsample_p_in VSS 1.55fF
C2406 clkgen.delay_155ns_1.genblk1\[1\].dly_binary.signal_w\[0\] VSS 1.69fF
C2407 clkgen.delay_155ns_1.genblk1\[0\].dly_binary.out VSS 1.67fF
C2408 clkgen.delay_155ns_1.genblk1\[1\].dly_binary.bypass_in VSS 1.16fF
C2409 clkgen.delay_155ns_1.genblk1\[1\].dly_binary.and_bypass_switch/a_207_413# VSS 0.16fF $ **FLOATING
C2410 clkgen.delay_155ns_1.genblk1\[1\].dly_binary.and_bypass_switch/a_27_413# VSS 0.19fF $ **FLOATING
C2411 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[0\] VSS 1.34fF
C2412 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.and_bypass_switch/a_207_413# VSS 0.16fF $ **FLOATING
C2413 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.and_bypass_switch/a_27_413# VSS 0.18fF $ **FLOATING
C2414 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[2\] VSS 1.06fF
C2415 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[3\] VSS 1.47fF
C2416 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit/mid VSS 1.43fF
C2417 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[31\].delay_unit/mid VSS 1.40fF
C2418 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[6\] VSS 2.09fF
C2419 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[7\] VSS 1.23fF
C2420 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit/mid VSS 1.32fF
C2421 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[0\] VSS 0.88fF
C2422 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.and_bypass_switch/a_207_413# VSS 0.18fF $ **FLOATING
C2423 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.and_bypass_switch/a_27_413# VSS 0.21fF $ **FLOATING
C2424 edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[0\] VSS 1.44fF
C2425 edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[1\] VSS 1.21fF
C2426 edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.genblk1\[0\].delay_unit/mid VSS 1.31fF
C2427 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[29\].delay_unit/mid VSS 1.31fF
C2428 VDD VSS 665.58fF
C2429 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[1\] VSS 1.38fF
C2430 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit/mid VSS 1.20fF
C2431 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[24\] VSS 1.35fF
C2432 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[25\] VSS 1.24fF
C2433 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[24\].delay_unit/mid VSS 1.28fF
C2434 clkgen.delay_155ns_3.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit/mid VSS 1.23fF
C2435 clkgen.delay_155ns_1.bypass_enable_w\[3\] VSS 0.72fF
C2436 dlycontrol1_in[3] VSS 4.43fF
C2437 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit/a_1691_329# VSS 0.10fF
C2438 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit/mid VSS 1.36fF
C2439 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[5\] VSS 1.91fF
C2440 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit/mid VSS 1.26fF
C2441 clkgen.delay_155ns_1.genblk1\[0\].dly_binary.and_bypass_switch/a_207_413# VSS 0.17fF $ **FLOATING
C2442 clkgen.delay_155ns_1.genblk1\[0\].dly_binary.and_bypass_switch/a_27_413# VSS 0.20fF $ **FLOATING
C2443 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[17\].delay_unit/mid VSS 1.33fF
C2444 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[3\] VSS 1.18fF
C2445 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit/mid VSS 1.35fF
C2446 clkgen.delay_155ns_2.genblk1\[1\].dly_binary.signal_w\[0\] VSS 2.12fF
C2447 clkgen.delay_155ns_2.genblk1\[0\].dly_binary.out VSS 3.22fF
C2448 clkgen.delay_155ns_2.genblk1\[1\].dly_binary.bypass_in VSS 3.31fF
C2449 clkgen.delay_155ns_2.genblk1\[1\].dly_binary.and_bypass_switch/a_207_413# VSS 0.16fF $ **FLOATING
C2450 clkgen.delay_155ns_2.genblk1\[1\].dly_binary.and_bypass_switch/a_27_413# VSS 0.19fF $ **FLOATING
C2451 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[6\] VSS 1.04fF
C2452 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[7\] VSS 1.09fF
C2453 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit/mid VSS 1.24fF
C2454 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[0\] VSS 1.52fF
C2455 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[0\].delay_unit/mid VSS 1.29fF
C2456 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit/mid VSS 1.22fF
C2457 clkgen.delay_155ns_3.genblk1\[2\].dly_binary.signal_w\[0\] VSS 0.79fF
C2458 clkgen.delay_155ns_3.genblk1\[2\].dly_binary.and_bypass_switch/a_207_413# VSS 0.17fF $ **FLOATING
C2459 clkgen.delay_155ns_3.genblk1\[2\].dly_binary.and_bypass_switch/a_27_413# VSS 0.20fF $ **FLOATING
C2460 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[8\] VSS 1.05fF
C2461 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.bypass_in VSS 2.42fF
C2462 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.out_mux/a_505_21# VSS 0.24fF
C2463 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.out_mux/a_76_199# VSS 0.16fF $ **FLOATING
C2464 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[12\] VSS 2.13fF
C2465 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[13\] VSS 1.28fF
C2466 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit/mid VSS 1.35fF
C2467 clkgen.delay_155ns_2.genblk1\[1\].dly_binary.signal_w\[2\] VSS 0.57fF
C2468 clkgen.delay_155ns_2.genblk1\[1\].dly_binary.out_mux/a_505_21# VSS 0.25fF
C2469 clkgen.delay_155ns_2.genblk1\[1\].dly_binary.out_mux/a_76_199# VSS 0.17fF $ **FLOATING
C2470 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[12\] VSS 1.22fF
C2471 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[13\] VSS 1.32fF
C2472 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[12\].delay_unit/a_1691_329# VSS 0.11fF
C2473 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[12\].delay_unit/mid VSS 1.34fF
C2474 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[2\] VSS 1.36fF
C2475 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit/mid VSS 1.26fF
C2476 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[3\] VSS 0.99fF
C2477 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[4\] VSS 0.97fF
C2478 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit/mid VSS 1.47fF
C2479 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[8\] VSS 1.29fF
C2480 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit/mid VSS 1.33fF
C2481 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[6\] VSS 1.62fF
C2482 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit/mid VSS 1.24fF
C2483 dlycontrol3_in[2] VSS 2.05fF
C2484 clkgen.delay_155ns_1.genblk1\[0\].dly_binary.signal_w\[0\] VSS 1.72fF
C2485 clkgen.delay_155ns_1.genblk1\[0\].dly_binary.genblk1\[0\].delay_unit/mid VSS 1.27fF
C2486 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[3\] VSS 1.14fF
C2487 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[2\].delay_unit/mid VSS 1.19fF
C2488 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[0\] VSS 1.13fF
C2489 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[1\] VSS 1.36fF
C2490 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[0\].delay_unit/mid VSS 1.29fF
C2491 clkgen.delay_155ns_2.genblk1\[0\].dly_binary.signal_w\[0\] VSS 4.06fF
C2492 clkgen.clk_dig_out VSS 3.15fF
C2493 clkgen.delay_155ns_2.genblk1\[0\].dly_binary.bypass_in VSS 4.89fF
C2494 clkgen.delay_155ns_2.genblk1\[0\].dly_binary.and_bypass_switch/a_207_413# VSS 0.16fF $ **FLOATING
C2495 clkgen.delay_155ns_2.genblk1\[0\].dly_binary.and_bypass_switch/a_27_413# VSS 0.18fF $ **FLOATING
C2496 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[14\] VSS 1.00fF
C2497 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[15\] VSS 1.42fF
C2498 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit/mid VSS 1.28fF
C2499 dlycontrol3_in[4] VSS 2.81fF
C2500 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit/a_1691_329# VSS 0.10fF
C2501 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit/mid VSS 1.31fF
C2502 clkgen.delay_155ns_3.genblk1\[1\].dly_binary.signal_w\[0\] VSS 1.87fF
C2503 clkgen.delay_155ns_3.genblk1\[0\].dly_binary.out VSS 0.28fF
C2504 clkgen.delay_155ns_3.genblk1\[1\].dly_binary.bypass_in VSS 1.64fF
C2505 clkgen.delay_155ns_3.genblk1\[1\].dly_binary.and_bypass_switch/a_207_413# VSS 0.19fF $ **FLOATING
C2506 clkgen.delay_155ns_3.genblk1\[1\].dly_binary.and_bypass_switch/a_27_413# VSS 0.18fF $ **FLOATING
C2507 clkgen.delay_155ns_3.bypass_enable_w\[1\] VSS 0.26fF
C2508 clkgen.delay_155ns_3.genblk1\[1\].bypass_enable/a_59_75# VSS 0.24fF $ **FLOATING
C2509 clkgen.delay_155ns_2.genblk1\[0\].bypass_enable/a_59_75# VSS 0.26fF $ **FLOATING
C2510 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit/mid VSS 1.36fF
C2511 edgedetect.dly_315ns_1.bypass_enable_w\[2\] VSS 0.32fF
C2512 dlycontrol4_in[2] VSS 1.71fF
C2513 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[5\].delay_unit/mid VSS 1.27fF
C2514 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.and_bypass_switch/a_207_413# VSS 0.18fF $ **FLOATING
C2515 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.and_bypass_switch/a_27_413# VSS 0.20fF $ **FLOATING
C2516 clkgen.delay_155ns_1.genblk1\[1\].dly_binary.genblk1\[0\].delay_unit/mid VSS 1.19fF
C2517 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[0\] VSS 1.39fF
C2518 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[0\].delay_unit/mid VSS 1.25fF
C2519 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit/mid VSS 1.26fF
C2520 clkgen.delay_155ns_3.genblk1\[0\].dly_binary.signal_w\[0\] VSS 1.96fF
C2521 clkgen.delay_155ns_3.genblk1\[0\].dly_binary.and_bypass_switch/a_207_413# VSS 0.16fF $ **FLOATING
C2522 clkgen.delay_155ns_3.genblk1\[0\].dly_binary.and_bypass_switch/a_27_413# VSS 0.18fF $ **FLOATING
C2523 clkgen.delay_155ns_1.bypass_enable_w\[4\] VSS 0.81fF
C2524 clkgen.delay_155ns_1.genblk1\[4\].bypass_enable/a_59_75# VSS 0.24fF $ **FLOATING
C2525 clkgen.delay_155ns_2.bypass_enable_w\[1\] VSS 0.38fF
C2526 dlycontrol2_in[1] VSS 3.88fF
C2527 clkgen.delay_155ns_2.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit/mid VSS 1.21fF
C2528 edgedetect.dly_315ns_1.bypass_enable_w\[3\] VSS 1.14fF
C2529 edgedetect.dly_315ns_1.genblk1\[3\].bypass_enable/a_59_75# VSS 0.23fF $ **FLOATING
C2530 clkgen.delay_155ns_1.enable_dlycontrol_w VSS 1.46fF
C2531 clkgen.delay_155ns_1.enablebuffer/a_27_47# VSS 0.50fF
C2532 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.and_bypass_switch/a_207_413# VSS 0.17fF $ **FLOATING
C2533 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.and_bypass_switch/a_27_413# VSS 0.20fF $ **FLOATING
C2534 clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[0\] VSS 1.61fF
C2535 clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[1\] VSS 1.05fF
C2536 clkgen.delay_155ns_1.genblk1\[2\].dly_binary.genblk1\[0\].delay_unit/mid VSS 1.26fF
C2537 edgedetect.dly_315ns_1.enablebuffer/a_27_47# VSS 0.50fF
C2538 nsample_n_1 VSS 0.53fF
C2539 nsample_n_in VSS 1.10fF
C2540 sampledly04/a_629_47# VSS 0.16fF $ **FLOATING
C2541 sampledly04/a_523_47# VSS 0.19fF
C2542 sampledly04/a_346_47# VSS 0.11fF $ **FLOATING
C2543 sampledly04/a_240_47# VSS 0.22fF $ **FLOATING
C2544 sampledly04/a_63_47# VSS 0.19fF $ **FLOATING
C2545 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.genblk1\[1\].delay_unit/mid VSS 1.28fF
C2546 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[30\] VSS 1.20fF
C2547 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[31\] VSS 1.42fF
C2548 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[30\].delay_unit/mid VSS 1.23fF
C2549 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit/mid VSS 1.25fF
C2550 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[28\] VSS 2.03fF
C2551 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[29\] VSS 1.02fF
C2552 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[28\].delay_unit/mid VSS 1.28fF
C2553 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[0\] VSS 2.60fF
C2554 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[0\].delay_unit/mid VSS 1.27fF
C2555 nsample_n_2 VSS 0.41fF
C2556 sampledly14/a_629_47# VSS 0.16fF $ **FLOATING
C2557 sampledly14/a_523_47# VSS 0.19fF
C2558 sampledly14/a_346_47# VSS 0.11fF $ **FLOATING
C2559 sampledly14/a_240_47# VSS 0.22fF $ **FLOATING
C2560 sampledly14/a_63_47# VSS 0.18fF $ **FLOATING
C2561 nsample_p_1 VSS 0.68fF
C2562 sampledly03/a_629_47# VSS 0.16fF $ **FLOATING
C2563 sampledly03/a_523_47# VSS 0.20fF
C2564 sampledly03/a_346_47# VSS 0.11fF $ **FLOATING
C2565 sampledly03/a_240_47# VSS 0.20fF $ **FLOATING
C2566 sampledly03/a_63_47# VSS 0.22fF $ **FLOATING
C2567 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[23\].delay_unit/mid VSS 1.27fF
C2568 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.and_bypass_switch/a_207_413# VSS 0.16fF $ **FLOATING
C2569 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.and_bypass_switch/a_27_413# VSS 0.19fF $ **FLOATING
C2570 clkgen.delay_155ns_3.genblk1\[2\].dly_binary.signal_w\[2\] VSS 1.30fF
C2571 clkgen.delay_155ns_3.genblk1\[2\].dly_binary.signal_w\[3\] VSS 1.32fF
C2572 clkgen.delay_155ns_3.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit/mid VSS 1.33fF
C2573 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[6\] VSS 1.03fF
C2574 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[7\] VSS 1.41fF
C2575 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit/mid VSS 1.51fF
C2576 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit/mid VSS 1.25fF
C2577 dlycontrol1_in[0] VSS 3.57fF
C2578 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[16\] VSS 1.00fF
C2579 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[17\] VSS 1.08fF
C2580 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[16\].delay_unit/mid VSS 1.24fF
C2581 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[2\] VSS 1.23fF
C2582 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit/mid VSS 1.27fF
C2583 sample_n_1 VSS 0.23fF
C2584 sample_n_in VSS 4.62fF
C2585 sampledly02/a_629_47# VSS 0.15fF $ **FLOATING
C2586 sampledly02/a_523_47# VSS 0.19fF
C2587 sampledly02/a_346_47# VSS 0.10fF $ **FLOATING
C2588 sampledly02/a_240_47# VSS 0.19fF $ **FLOATING
C2589 sampledly02/a_63_47# VSS 0.21fF $ **FLOATING
C2590 nsample_n_3 VSS 0.48fF
C2591 sampledly24/a_629_47# VSS 0.16fF $ **FLOATING
C2592 sampledly24/a_523_47# VSS 0.22fF
C2593 sampledly24/a_346_47# VSS 0.11fF $ **FLOATING
C2594 sampledly24/a_240_47# VSS 0.19fF $ **FLOATING
C2595 sampledly24/a_63_47# VSS 0.19fF $ **FLOATING
C2596 nsample_p_2 VSS 0.31fF
C2597 sampledly13/a_629_47# VSS 0.16fF $ **FLOATING
C2598 sampledly13/a_523_47# VSS 0.19fF
C2599 sampledly13/a_346_47# VSS 0.10fF $ **FLOATING
C2600 sampledly13/a_240_47# VSS 0.19fF $ **FLOATING
C2601 sampledly13/a_63_47# VSS 0.17fF $ **FLOATING
C2602 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit/mid VSS 1.25fF
C2603 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[13\] VSS 1.19fF
C2604 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit/mid VSS 1.22fF
C2605 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[7\] VSS 1.02fF
C2606 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[8\] VSS 2.53fF
C2607 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit/mid VSS 1.27fF
C2608 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit/mid VSS 1.26fF
C2609 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit/a_1691_329# VSS 0.10fF
C2610 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit/mid VSS 1.51fF
C2611 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[11\].delay_unit/mid VSS 1.31fF
C2612 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[0\] VSS 1.42fF
C2613 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[1\] VSS 0.91fF
C2614 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[0\].delay_unit/mid VSS 1.27fF
C2615 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit/mid VSS 1.28fF
C2616 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.bypass_in VSS 5.00fF
C2617 edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.and_bypass_switch/a_207_413# VSS 0.17fF $ **FLOATING
C2618 edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.and_bypass_switch/a_27_413# VSS 0.20fF $ **FLOATING
C2619 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[7\] VSS 1.04fF
C2620 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit/mid VSS 1.33fF
C2621 clkgen.delay_155ns_3.bypass_enable_w\[4\] VSS 0.20fF
C2622 sampledly12/a_629_47# VSS 0.16fF $ **FLOATING
C2623 sampledly12/a_523_47# VSS 0.19fF
C2624 sampledly12/a_346_47# VSS 0.10fF $ **FLOATING
C2625 sampledly12/a_240_47# VSS 0.19fF $ **FLOATING
C2626 sampledly12/a_63_47# VSS 0.19fF $ **FLOATING
C2627 nsample_n_4 VSS 0.47fF
C2628 sampledly34/a_629_47# VSS 0.20fF $ **FLOATING
C2629 sampledly34/a_523_47# VSS 0.24fF
C2630 sampledly34/a_346_47# VSS 0.18fF $ **FLOATING
C2631 sampledly34/a_240_47# VSS 0.29fF $ **FLOATING
C2632 sampledly34/a_63_47# VSS 0.27fF $ **FLOATING
C2633 sample_p_1 VSS 0.30fF
C2634 sampledly01/a_629_47# VSS 0.16fF $ **FLOATING
C2635 sampledly01/a_523_47# VSS 0.20fF
C2636 sampledly01/a_346_47# VSS 0.11fF $ **FLOATING
C2637 sampledly01/a_240_47# VSS 0.20fF $ **FLOATING
C2638 sampledly01/a_63_47# VSS 0.21fF $ **FLOATING
C2639 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[4\] VSS 2.06fF
C2640 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[5\] VSS 1.23fF
C2641 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit/mid VSS 1.26fF
C2642 nsample_p_3 VSS 0.41fF
C2643 sampledly23/a_629_47# VSS 0.18fF $ **FLOATING
C2644 sampledly23/a_523_47# VSS 0.20fF
C2645 sampledly23/a_346_47# VSS 0.11fF $ **FLOATING
C2646 sampledly23/a_240_47# VSS 0.20fF $ **FLOATING
C2647 sampledly23/a_63_47# VSS 0.21fF $ **FLOATING
C2648 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.out_mux/a_505_21# VSS 0.26fF
C2649 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.out_mux/a_76_199# VSS 0.18fF $ **FLOATING
C2650 clkgen.delay_155ns_3.genblk1\[1\].dly_binary.signal_w\[2\] VSS 0.38fF
C2651 clkgen.delay_155ns_3.genblk1\[1\].dly_binary.out VSS 0.33fF
C2652 clkgen.delay_155ns_3.genblk1\[1\].dly_binary.out_mux/a_505_21# VSS 0.24fF
C2653 clkgen.delay_155ns_3.genblk1\[1\].dly_binary.out_mux/a_76_199# VSS 0.17fF $ **FLOATING
C2654 clkgen.delay_155ns_3.genblk1\[0\].bypass_enable/a_59_75# VSS 0.22fF $ **FLOATING
C2655 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[2\] VSS 1.32fF
C2656 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit/mid VSS 1.30fF
C2657 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[7\] VSS 0.95fF
C2658 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[8\] VSS 1.15fF
C2659 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit/mid VSS 1.31fF
C2660 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit/mid VSS 1.35fF
C2661 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[9\] VSS 1.00fF
C2662 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[10\] VSS 1.40fF
C2663 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[9\].delay_unit/mid VSS 1.36fF
C2664 sample_n_2 VSS 0.60fF
C2665 sampledly22/a_629_47# VSS 0.16fF $ **FLOATING
C2666 sampledly22/a_523_47# VSS 0.20fF
C2667 sampledly22/a_346_47# VSS 0.11fF $ **FLOATING
C2668 sampledly22/a_240_47# VSS 0.20fF $ **FLOATING
C2669 sampledly22/a_63_47# VSS 0.21fF $ **FLOATING
C2670 sampledly11/a_629_47# VSS 0.15fF $ **FLOATING
C2671 sampledly11/a_523_47# VSS 0.19fF
C2672 sampledly11/a_346_47# VSS 0.11fF $ **FLOATING
C2673 sampledly11/a_240_47# VSS 0.20fF $ **FLOATING
C2674 sampledly11/a_63_47# VSS 0.22fF $ **FLOATING
C2675 dlycontrol4_in[4] VSS 3.31fF
C2676 nsample_p_4 VSS 0.23fF
C2677 sampledly33/a_629_47# VSS 0.16fF $ **FLOATING
C2678 sampledly33/a_523_47# VSS 0.23fF
C2679 sampledly33/a_346_47# VSS 0.18fF $ **FLOATING
C2680 sampledly33/a_240_47# VSS 0.26fF $ **FLOATING
C2681 sampledly33/a_63_47# VSS 0.19fF $ **FLOATING
C2682 ndecision_finish_in VSS 3.63fF
C2683 inbuf_3/a_27_47# VSS 0.27fF $ **FLOATING
C2684 clkgen.delay_155ns_2.genblk1\[0\].dly_binary.genblk1\[0\].delay_unit/mid VSS 1.21fF
C2685 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[2\] VSS 0.94fF
C2686 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[3\] VSS 2.09fF
C2687 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[2\].delay_unit/mid VSS 1.25fF
C2688 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[4\] VSS 1.37fF
C2689 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[5\] VSS 1.30fF
C2690 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[4\].delay_unit/mid VSS 1.24fF
C2691 edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.bypass_in VSS 3.49fF
C2692 edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.and_bypass_switch/a_207_413# VSS 0.17fF $ **FLOATING
C2693 edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.and_bypass_switch/a_27_413# VSS 0.20fF $ **FLOATING
C2694 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.out VSS 1.50fF
C2695 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[16\] VSS 4.47fF
C2696 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.bypass_in VSS 2.08fF
C2697 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.out VSS 1.79fF
C2698 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.out_mux/a_505_21# VSS 0.25fF
C2699 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.out_mux/a_76_199# VSS 0.18fF $ **FLOATING
C2700 clkgen.delay_155ns_1.genblk1\[1\].dly_binary.out VSS 0.61fF
C2701 clkgen.delay_155ns_1.genblk1\[2\].dly_binary.signal_w\[4\] VSS 0.73fF
C2702 clkgen.delay_155ns_1.genblk1\[2\].dly_binary.out_mux/a_505_21# VSS 0.25fF
C2703 clkgen.delay_155ns_1.genblk1\[2\].dly_binary.out_mux/a_76_199# VSS 0.16fF $ **FLOATING
C2704 clkgen.delay_155ns_1.genblk1\[0\].dly_binary.in VSS 1.26fF
C2705 clkgen.delay_155ns_1.genblk1\[0\].dly_binary.signal_w\[1\] VSS 0.49fF
C2706 clkgen.delay_155ns_1.genblk1\[0\].dly_binary.out_mux/a_505_21# VSS 0.29fF
C2707 clkgen.delay_155ns_1.genblk1\[0\].dly_binary.out_mux/a_76_199# VSS 0.17fF $ **FLOATING
C2708 sample_n_4 VSS 0.24fF
C2709 sample_n_3 VSS 0.35fF
C2710 sampledly32/a_629_47# VSS 0.16fF $ **FLOATING
C2711 sampledly32/a_523_47# VSS 0.20fF
C2712 sampledly32/a_346_47# VSS 0.11fF $ **FLOATING
C2713 sampledly32/a_240_47# VSS 0.20fF $ **FLOATING
C2714 sampledly32/a_63_47# VSS 0.22fF $ **FLOATING
C2715 sample_p_3 VSS 0.42fF
C2716 sample_p_2 VSS 1.20fF
C2717 sampledly21/a_629_47# VSS 0.17fF $ **FLOATING
C2718 sampledly21/a_523_47# VSS 0.21fF
C2719 sampledly21/a_346_47# VSS 0.11fF $ **FLOATING
C2720 sampledly21/a_240_47# VSS 0.20fF $ **FLOATING
C2721 sampledly21/a_63_47# VSS 0.22fF $ **FLOATING
C2722 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[15\] VSS 1.33fF
C2723 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit/mid VSS 1.64fF
C2724 inbuf_2/a_27_47# VSS 0.28fF $ **FLOATING
C2725 clkgen.delay_155ns_2.bypass_enable_w\[4\] VSS 0.39fF
C2726 clkgen.delay_155ns_2.genblk1\[4\].bypass_enable/a_59_75# VSS 0.26fF $ **FLOATING
C2727 clkgen.delay_155ns_1.genblk1\[3\].bypass_enable/a_59_75# VSS 0.26fF $ **FLOATING
C2728 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[11\] VSS 1.14fF
C2729 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[10\].delay_unit/mid VSS 1.25fF
C2730 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[16\] VSS 2.79fF
C2731 edgedetect.dly_315ns_1.genblk1\[2\].bypass_enable/a_59_75# VSS 0.24fF $ **FLOATING
C2732 clkgen.delay_155ns_2.genblk1\[1\].dly_binary.signal_w\[1\] VSS 1.17fF
C2733 clkgen.delay_155ns_2.genblk1\[1\].dly_binary.genblk1\[0\].delay_unit/mid VSS 1.26fF
C2734 sampledly31/a_629_47# VSS 0.17fF $ **FLOATING
C2735 sampledly31/a_523_47# VSS 0.21fF
C2736 sampledly31/a_346_47# VSS 0.12fF $ **FLOATING
C2737 sampledly31/a_240_47# VSS 0.21fF $ **FLOATING
C2738 sampledly31/a_63_47# VSS 0.20fF $ **FLOATING
C2739 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.out VSS 2.81fF
C2740 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[16\] VSS 2.59fF
C2741 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.bypass_in VSS 2.96fF
C2742 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.out VSS 3.22fF
C2743 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.out_mux/a_505_21# VSS 0.25fF
C2744 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.out_mux/a_76_199# VSS 0.17fF $ **FLOATING
C2745 ena_in VSS 3.72fF
C2746 inbuf_1/a_27_47# VSS 0.29fF $ **FLOATING
C2747 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.and_bypass_switch/a_207_413# VSS 0.17fF $ **FLOATING
C2748 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.and_bypass_switch/a_27_413# VSS 0.19fF $ **FLOATING
C2749 edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.signal_w\[4\] VSS 1.83fF
C2750 edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.out_mux/a_505_21# VSS 0.24fF
C2751 edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.out_mux/a_76_199# VSS 0.17fF $ **FLOATING
C2752 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.in VSS 2.41fF
C2753 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.bypass_in VSS 3.53fF
C2754 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.out VSS 0.53fF
C2755 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.out_mux/a_505_21# VSS 0.23fF
C2756 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.out_mux/a_76_199# VSS 0.17fF $ **FLOATING
C2757 clkgen.delay_155ns_3.genblk1\[1\].dly_binary.signal_w\[1\] VSS 0.90fF
C2758 clkgen.delay_155ns_3.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit/mid VSS 1.23fF
C2759 edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit/mid VSS 1.37fF
C2760 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[1\] VSS 1.20fF
C2761 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.genblk1\[0\].delay_unit/mid VSS 1.23fF
C2762 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[4\] VSS 2.01fF
C2763 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.signal_w\[5\] VSS 1.48fF
C2764 clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit/mid VSS 1.27fF
C2765 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[27\].delay_unit/mid VSS 1.28fF
C2766 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[23\] VSS 1.68fF
C2767 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[22\].delay_unit/mid VSS 1.29fF
C2768 dlycontrol1_in[2] VSS 2.28fF
C2769 clkgen.delay_155ns_3.genblk1\[2\].dly_binary.genblk1\[1\].delay_unit/mid VSS 1.33fF
C2770 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit/a_1691_329# VSS 0.10fF
C2771 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit/mid VSS 1.30fF
C2772 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.signal_w\[4\] VSS 1.17fF
C2773 edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit/mid VSS 1.30fF
C2774 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[10\] VSS 1.48fF
C2775 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit/mid VSS 1.37fF
C2776 clkgen.delay_155ns_3.genblk1\[0\].dly_binary.in VSS 1.91fF
C2777 clkgen.clk_dig_delayed_w VSS 0.51fF
C2778 clkgen.nor1/a_74_47# VSS 0.22fF $ **FLOATING
C2779 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit/mid VSS 1.21fF
C2780 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[15\].delay_unit/mid VSS 1.32fF
C2781 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[0\] VSS 1.54fF
C2782 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.signal_w\[1\] VSS 1.61fF
C2783 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[0\].delay_unit/mid VSS 1.21fF
C2784 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[4\] VSS 0.93fF
C2785 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.signal_w\[5\] VSS 1.25fF
C2786 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit/mid VSS 1.21fF
C2787 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit/mid VSS 1.27fF
C2788 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[12\] VSS 1.59fF
C2789 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit/mid VSS 1.48fF
C2790 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.signal_w\[9\] VSS 1.49fF
C2791 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit/mid VSS 1.20fF
C2792 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[10\] VSS 1.09fF
C2793 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.signal_w\[11\] VSS 1.32fF
C2794 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[10\].delay_unit/mid VSS 1.28fF
C2795 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[11\] VSS 1.33fF
C2796 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[10\].delay_unit/mid VSS 1.31fF
C2797 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[1\] VSS 1.00fF
C2798 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.signal_w\[2\] VSS 1.16fF
C2799 clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit/mid VSS 1.18fF
C2800 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[5\] VSS 1.01fF
C2801 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[6\] VSS 1.05fF
C2802 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit/a_1691_329# VSS 0.10fF
C2803 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit/mid VSS 1.49fF
C2804 edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit/mid VSS 1.23fF
C2805 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[0\] VSS 1.05fF
C2806 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[1\] VSS 1.40fF
C2807 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[0\].delay_unit/mid VSS 1.26fF
C2808 edgedetect.nor1/a_74_47# VSS 0.27fF $ **FLOATING
C2809 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit/mid VSS 1.29fF
C2810 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[12\] VSS 1.19fF
C2811 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.signal_w\[13\] VSS 1.34fF
C2812 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit/a_1691_329# VSS 0.14fF
C2813 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit/mid VSS 1.41fF
C2814 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.signal_w\[8\] VSS 1.10fF
C2815 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[8\].delay_unit/a_1691_329# VSS 0.11fF
C2816 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[8\].delay_unit/mid VSS 1.34fF
C2817 dlycontrol4_in[1] VSS 4.77fF
C2818 clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit/mid VSS 1.28fF
C2819 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[3\].delay_unit/mid VSS 1.39fF
C2820 clkgen.delay_155ns_3.genblk1\[4\].bypass_enable/a_59_75# VSS 0.24fF $ **FLOATING
C2821 clkgen.delay_155ns_2.bypass_enable_w\[3\] VSS 1.40fF
C2822 clkgen.delay_155ns_2.genblk1\[3\].bypass_enable/a_59_75# VSS 0.25fF $ **FLOATING
C2823 clkgen.delay_155ns_1.bypass_enable_w\[2\] VSS 0.81fF
C2824 clkgen.delay_155ns_1.genblk1\[2\].bypass_enable/a_59_75# VSS 0.23fF $ **FLOATING
C2825 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit/a_1691_329# VSS 0.14fF
C2826 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit/mid VSS 1.51fF
C2827 edgedetect.dly_315ns_1.bypass_enable_w\[1\] VSS 0.20fF
C2828 edgedetect.dly_315ns_1.genblk1\[1\].bypass_enable/a_59_75# VSS 0.25fF $ **FLOATING
C2829 clkgen.delay_155ns_3.genblk1\[0\].dly_binary.genblk1\[0\].delay_unit/mid VSS 1.28fF
C2830 clkgen.enable_loop_in VSS 0.65fF
C2831 edgedetect.start_conv_edge_w VSS 1.32fF
C2832 edgedetect.ena_in VSS 3.12fF
C2833 edgedetect.or1/a_68_297# VSS 0.22fF $ **FLOATING
C2834 clkgen.delay_155ns_2.genblk1\[3\].dly_binary.out VSS 0.67fF
C2835 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.out_mux/a_505_21# VSS 0.25fF
C2836 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.out_mux/a_76_199# VSS 0.16fF $ **FLOATING
C2837 clkgen.delay_155ns_2.genblk1\[1\].dly_binary.out VSS 0.73fF
C2838 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.signal_w\[4\] VSS 2.74fF
C2839 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.bypass_in VSS 1.32fF
C2840 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.out VSS 1.34fF
C2841 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.out_mux/a_505_21# VSS 0.25fF
C2842 clkgen.delay_155ns_2.genblk1\[2\].dly_binary.out_mux/a_76_199# VSS 0.17fF $ **FLOATING
C2843 clkgen.delay_155ns_2.genblk1\[0\].dly_binary.signal_w\[1\] VSS 0.74fF
C2844 clkgen.delay_155ns_2.genblk1\[0\].dly_binary.out_mux/a_505_21# VSS 0.24fF
C2845 clkgen.delay_155ns_2.genblk1\[0\].dly_binary.out_mux/a_76_199# VSS 0.20fF $ **FLOATING
C2846 clkgen.delay_155ns_2.bypass_enable_w\[0\] VSS 0.43fF
C2847 dlycontrol2_in[0] VSS 2.24fF
.ends

