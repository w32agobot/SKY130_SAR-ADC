* SPICE3 file created from adc_array_fingercap_8(8).ext - technology: sky130A

C0 cbot ctop 5.96fF
