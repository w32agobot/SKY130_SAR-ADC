* SPICE3 file created from sky130_mm_sc_hd_dlyPoly6ns.ext - technology: sky130A

.subckt sky130_mm_sc_hd_dlyPoly6ns_postlayout VPWR in out VGND VNB VPB
X0 cap_top in VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.0453e+12p ps=9.52e+06u w=420000u l=3.83e+06u
X1 a_1724_71# cap_top VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VPWR out a_1724_71# VNB sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3 VGND out a_1783_329# VPB sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4 a_1783_329# out VGND VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5 a_1724_71# out VPWR VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VGND cap_top VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X7 a_1783_329# cap_top VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.72e+11p ps=4.38e+06u w=800000u l=150000u
X8 out cap_top a_1783_329# VPB sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X9 cap_top in VPWR VPB sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=800000u l=3.83e+06u
X10 out cap_top a_1724_71# VNB sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
C0 VGND VPWR 0.34fF
C1 VGND in 0.38fF
C2 cap_top VPB 0.17fF
C3 a_1783_329# a_1724_71# 0.00fF
C4 VGND out 0.11fF
C5 VPWR a_1724_71# 0.07fF
C6 a_1724_71# in 0.00fF
C7 VGND VPB 0.15fF
C8 a_1724_71# out 0.13fF
C9 VGND cap_top 2.50fF
C10 a_1783_329# VPWR 0.98fF
C11 a_1783_329# in 0.00fF
C12 VPB a_1724_71# 0.00fF
C13 a_1783_329# out 0.06fF
C14 cap_top a_1724_71# 0.13fF
C15 VPWR in 0.22fF
C16 VPWR out 0.29fF
C17 a_1783_329# VPB 0.02fF
C18 out in 0.00fF
C19 a_1783_329# cap_top 0.03fF
C20 VGND a_1724_71# 0.77fF
C21 VPWR VPB 0.28fF
C22 VPB in 0.23fF
C23 cap_top VPWR 0.52fF
C24 VPB out 0.05fF
C25 cap_top in 0.19fF
C26 a_1783_329# VGND 0.46fF
C27 cap_top out 0.05fF
C28 VPWR VNB 1.20fF
C29 in VNB 1.50fF
C30 out VNB 0.34fF
C31 VPB VNB 2.04fF
C32 a_1724_71# VNB 0.04fF **FLOATING
C33 a_1783_329# VNB 0.07fF **FLOATING
C34 cap_top VNB 0.90fF **FLOATING
.ends
