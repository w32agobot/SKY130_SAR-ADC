* NGSPICE file created from sky130_mm_sc_hd_dlyxns.ext - technology: sky130A

.subckt sky130_mm_sc_hd_dlyxns in out VPWR VGND VNB VPB
X0 a_1184_80# out VPWR VNB sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1 VPWR out a_1184_80# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 cap_top in VGND VNB sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=1.0337e+12p ps=9.44e+06u w=420000u l=350000u
X3 VGND out a_1162_296# VPB sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u
X4 a_1162_296# out VGND VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5 a_1162_296# cap_top VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.72e+11p ps=4.38e+06u w=800000u l=150000u
X6 out cap_top a_1162_296# VPB sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X7 cap_top in VPWR VPB sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=350000u
X8 out cap_top a_1184_80# VNB sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X9 VGND cap_top VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.355e+06u l=2.25e+06u
X10 a_1184_80# cap_top VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
C0 m1_394_79# out 0.00fF
C1 VGND VPB 0.08fF
C2 a_1184_80# cap_top 0.01fF
C3 m1_394_79# in 0.00fF
C4 VGND a_1162_296# 0.16fF
C5 a_1184_80# VPWR 0.10fF
C6 cap_top VPWR 0.68fF
C7 a_1184_80# out 0.35fF
C8 VPB m1_394_79# 0.00fF
C9 cap_top out 0.09fF
C10 a_1184_80# in 0.00fF
C11 cap_top in 0.03fF
C12 VPWR out 0.14fF
C13 VPWR in 0.02fF
C14 a_1184_80# VPB 0.00fF
C15 in out 0.00fF
C16 cap_top VPB 0.14fF
C17 a_1184_80# a_1162_296# 0.02fF
C18 VGND m1_394_79# 1.04fF
C19 a_1162_296# cap_top 0.04fF
C20 VPWR VPB 0.25fF
C21 VPB out 0.07fF
C22 a_1162_296# VPWR 1.11fF
C23 VPB in 0.05fF
C24 a_1162_296# out 0.41fF
C25 a_1184_80# VGND 1.06fF
C26 a_1162_296# in 0.00fF
C27 VGND cap_top 0.88fF
C28 VGND VPWR 0.25fF
C29 VGND out 0.15fF
C30 a_1162_296# VPB 0.03fF
C31 a_1184_80# m1_394_79# 0.02fF
C32 VGND in 0.02fF
C33 cap_top m1_394_79# 1.16fF
C34 VPWR m1_394_79# 0.00fF
.ends

