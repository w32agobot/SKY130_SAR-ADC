magic
tech sky130A
magscale 1 2
timestamp 1681461446
<< nwell >>
rect 180 224 3820 3776
<< pwell >>
rect 0 3776 4000 4000
rect 0 224 180 3776
rect 3820 224 4000 3776
rect 0 0 4000 224
<< varactor >>
rect 360 400 3640 3600
<< psubdiff >>
rect 890 3900 1350 3920
rect 890 3850 920 3900
rect 1320 3850 1350 3900
rect 890 3830 1350 3850
rect 2650 3900 3110 3920
rect 2650 3850 2680 3900
rect 3080 3850 3110 3900
rect 2650 3830 3110 3850
rect 80 3080 154 3110
rect 80 2680 100 3080
rect 150 2680 154 3080
rect 80 2650 154 2680
rect 80 1320 154 1350
rect 80 920 100 1320
rect 150 920 154 1320
rect 80 890 154 920
rect 3846 3080 3920 3110
rect 3846 2680 3850 3080
rect 3900 2680 3920 3080
rect 3846 2650 3920 2680
rect 3846 1320 3920 1350
rect 3846 920 3850 1320
rect 3900 920 3920 1320
rect 3846 890 3920 920
rect 890 150 1350 170
rect 890 100 920 150
rect 1320 100 1350 150
rect 890 80 1350 100
rect 2650 150 3110 170
rect 2650 100 2680 150
rect 3080 100 3110 150
rect 2650 80 3110 100
<< nsubdiff >>
rect 360 3720 3640 3740
rect 360 3653 420 3720
rect 3570 3653 3640 3720
rect 360 3600 3640 3653
rect 360 347 3640 400
rect 360 280 420 347
rect 3570 280 3640 347
rect 360 260 3640 280
<< psubdiffcont >>
rect 920 3850 1320 3900
rect 2680 3850 3080 3900
rect 100 2680 150 3080
rect 100 920 150 1320
rect 3850 2680 3900 3080
rect 3850 920 3900 1320
rect 920 100 1320 150
rect 2680 100 3080 150
<< nsubdiffcont >>
rect 420 3653 3570 3720
rect 420 280 3570 347
<< poly >>
rect 320 3150 360 3600
rect 210 2960 360 3150
rect 210 1050 240 2960
rect 313 1050 360 2960
rect 210 840 360 1050
rect 320 400 360 840
rect 3640 3150 3680 3600
rect 3640 2960 3790 3150
rect 3640 1050 3687 2960
rect 3760 1050 3790 2960
rect 3640 840 3790 1050
rect 3640 400 3680 840
<< polycont >>
rect 240 1050 313 2960
rect 3687 1050 3760 2960
<< locali >>
rect 890 3920 1350 4000
rect 2650 3920 3110 4000
rect 80 3900 3920 3920
rect 80 3850 920 3900
rect 1320 3850 2680 3900
rect 3080 3850 3920 3900
rect 80 3840 3920 3850
rect 80 3110 160 3840
rect 890 3830 1350 3840
rect 2650 3830 3110 3840
rect 360 3620 420 3720
rect 540 3620 580 3653
rect 700 3620 740 3653
rect 860 3620 900 3653
rect 1020 3620 1060 3653
rect 1180 3620 2820 3653
rect 2940 3620 2980 3653
rect 3100 3620 3140 3653
rect 3260 3620 3300 3653
rect 3420 3620 3460 3653
rect 3570 3620 3640 3720
rect 360 3600 3640 3620
rect 240 3520 1040 3560
rect 240 3400 320 3520
rect 1080 3480 1150 3600
rect 360 3440 1150 3480
rect 240 3360 1040 3400
rect 240 3240 320 3360
rect 1080 3320 1150 3440
rect 360 3280 1150 3320
rect 240 3200 1040 3240
rect 0 3080 170 3110
rect 0 2680 100 3080
rect 150 2680 170 3080
rect 0 2650 170 2680
rect 240 3080 320 3200
rect 1080 3160 1150 3280
rect 360 3120 1150 3160
rect 240 3040 1040 3080
rect 240 2960 320 3040
rect 1080 3000 1150 3120
rect 360 2960 1150 3000
rect 80 1350 160 2650
rect 0 1320 170 1350
rect 0 920 100 1320
rect 150 920 170 1320
rect 0 890 170 920
rect 313 2920 320 2960
rect 313 2880 1040 2920
rect 313 2760 320 2880
rect 1080 2840 1150 2960
rect 360 2800 1150 2840
rect 313 2720 1040 2760
rect 313 2600 320 2720
rect 1080 2680 1150 2800
rect 360 2640 1150 2680
rect 313 2560 1040 2600
rect 313 2440 320 2560
rect 1080 2520 1150 2640
rect 360 2480 1150 2520
rect 313 2400 1040 2440
rect 313 2280 320 2400
rect 1080 2360 1150 2480
rect 360 2320 1150 2360
rect 313 2240 1040 2280
rect 313 2120 320 2240
rect 1080 2200 1150 2320
rect 360 2160 1150 2200
rect 313 2080 1040 2120
rect 1080 2080 1150 2160
rect 313 2040 320 2080
rect 1190 2040 1230 3560
rect 1270 2080 1310 3600
rect 1350 2040 1390 3560
rect 1430 2080 1470 3600
rect 1510 2040 1550 3560
rect 1590 2080 1630 3600
rect 1670 2040 1710 3560
rect 1750 2080 1790 3600
rect 1830 2040 1870 3560
rect 313 1960 1870 2040
rect 313 1920 320 1960
rect 313 1880 1040 1920
rect 313 1760 320 1880
rect 1080 1840 1150 1920
rect 360 1800 1150 1840
rect 313 1720 1040 1760
rect 313 1600 320 1720
rect 1080 1680 1150 1800
rect 360 1640 1150 1680
rect 313 1560 1040 1600
rect 313 1440 320 1560
rect 1080 1520 1150 1640
rect 360 1480 1150 1520
rect 313 1400 1040 1440
rect 313 1280 320 1400
rect 1080 1360 1150 1480
rect 360 1320 1150 1360
rect 313 1240 1040 1280
rect 313 1120 320 1240
rect 1080 1200 1150 1320
rect 360 1160 1150 1200
rect 313 1080 1040 1120
rect 313 1050 320 1080
rect 240 960 320 1050
rect 1080 1040 1150 1160
rect 360 1000 1150 1040
rect 240 920 1040 960
rect 80 160 160 890
rect 240 800 320 920
rect 1080 880 1150 1000
rect 360 840 1150 880
rect 240 760 1040 800
rect 240 640 320 760
rect 1080 720 1150 840
rect 360 680 1150 720
rect 240 600 1040 640
rect 240 480 320 600
rect 1080 560 1150 680
rect 360 520 1150 560
rect 240 440 1040 480
rect 1080 400 1150 520
rect 1190 440 1230 1960
rect 1270 400 1310 1920
rect 1350 440 1390 1960
rect 1430 400 1470 1920
rect 1510 440 1550 1960
rect 1590 400 1630 1920
rect 1670 440 1710 1960
rect 1750 400 1790 1920
rect 1830 440 1870 1960
rect 1910 400 2090 3600
rect 2130 2040 2170 3560
rect 2210 2080 2250 3600
rect 2290 2040 2330 3560
rect 2370 2080 2410 3600
rect 2450 2040 2490 3560
rect 2530 2080 2570 3600
rect 2610 2040 2650 3560
rect 2690 2080 2730 3600
rect 2770 2040 2810 3560
rect 2850 3480 2920 3600
rect 2960 3520 3760 3560
rect 2850 3440 3640 3480
rect 2850 3320 2920 3440
rect 3680 3400 3760 3520
rect 2960 3360 3760 3400
rect 2850 3280 3640 3320
rect 2850 3160 2920 3280
rect 3680 3240 3760 3360
rect 2960 3200 3760 3240
rect 2850 3120 3640 3160
rect 2850 3000 2920 3120
rect 3680 3080 3760 3200
rect 3840 3110 3920 3840
rect 2960 3040 3760 3080
rect 2850 2960 3640 3000
rect 3680 2960 3760 3040
rect 2850 2840 2920 2960
rect 3680 2920 3687 2960
rect 2960 2880 3687 2920
rect 2850 2800 3640 2840
rect 2850 2680 2920 2800
rect 3680 2760 3687 2880
rect 2960 2720 3687 2760
rect 2850 2640 3640 2680
rect 2850 2520 2920 2640
rect 3680 2600 3687 2720
rect 2960 2560 3687 2600
rect 2850 2480 3640 2520
rect 2850 2360 2920 2480
rect 3680 2440 3687 2560
rect 2960 2400 3687 2440
rect 2850 2320 3640 2360
rect 2850 2200 2920 2320
rect 3680 2280 3687 2400
rect 2960 2240 3687 2280
rect 2850 2160 3640 2200
rect 2850 2080 2920 2160
rect 3680 2120 3687 2240
rect 2960 2080 3687 2120
rect 3680 2040 3687 2080
rect 2130 1960 3687 2040
rect 2130 440 2170 1960
rect 2210 400 2250 1920
rect 2290 440 2330 1960
rect 2370 400 2410 1920
rect 2450 440 2490 1960
rect 2530 400 2570 1920
rect 2610 440 2650 1960
rect 2690 400 2730 1920
rect 2770 440 2810 1960
rect 3680 1920 3687 1960
rect 2850 1840 2920 1920
rect 2960 1880 3687 1920
rect 2850 1800 3640 1840
rect 2850 1680 2920 1800
rect 3680 1760 3687 1880
rect 2960 1720 3687 1760
rect 2850 1640 3640 1680
rect 2850 1520 2920 1640
rect 3680 1600 3687 1720
rect 2960 1560 3687 1600
rect 2850 1480 3640 1520
rect 2850 1360 2920 1480
rect 3680 1440 3687 1560
rect 2960 1400 3687 1440
rect 2850 1320 3640 1360
rect 2850 1200 2920 1320
rect 3680 1280 3687 1400
rect 2960 1240 3687 1280
rect 2850 1160 3640 1200
rect 2850 1040 2920 1160
rect 3680 1120 3687 1240
rect 2960 1080 3687 1120
rect 3680 1050 3687 1080
rect 3830 3080 4000 3110
rect 3830 2680 3850 3080
rect 3900 2680 4000 3080
rect 3830 2650 4000 2680
rect 3840 1350 3920 2650
rect 2850 1000 3640 1040
rect 2850 880 2920 1000
rect 3680 960 3760 1050
rect 2960 920 3760 960
rect 2850 840 3640 880
rect 2850 720 2920 840
rect 3680 800 3760 920
rect 3830 1320 4000 1350
rect 3830 920 3850 1320
rect 3900 920 4000 1320
rect 3830 890 4000 920
rect 2960 760 3760 800
rect 2850 680 3640 720
rect 2850 560 2920 680
rect 3680 640 3760 760
rect 2960 600 3760 640
rect 2850 520 3640 560
rect 2850 400 2920 520
rect 3680 480 3760 600
rect 2960 440 3760 480
rect 360 380 3640 400
rect 360 280 420 380
rect 540 347 580 380
rect 700 347 740 380
rect 860 347 900 380
rect 1020 347 1060 380
rect 1180 347 2820 380
rect 2940 347 2980 380
rect 3100 347 3140 380
rect 3260 347 3300 380
rect 3420 347 3460 380
rect 3570 280 3640 380
rect 890 160 1350 170
rect 2650 160 3110 170
rect 3840 160 3920 890
rect 80 150 3920 160
rect 80 100 920 150
rect 1320 100 2680 150
rect 3080 100 3920 150
rect 80 80 3920 100
rect 890 0 1350 80
rect 2650 0 3110 80
<< viali >>
rect 420 3653 540 3720
rect 580 3653 700 3720
rect 740 3653 860 3720
rect 900 3653 1020 3720
rect 1060 3653 1180 3720
rect 2820 3653 2940 3720
rect 2980 3653 3100 3720
rect 3140 3653 3260 3720
rect 3300 3653 3420 3720
rect 3460 3653 3570 3720
rect 420 3620 540 3653
rect 580 3620 700 3653
rect 740 3620 860 3653
rect 900 3620 1020 3653
rect 1060 3620 1180 3653
rect 2820 3620 2940 3653
rect 2980 3620 3100 3653
rect 3140 3620 3260 3653
rect 3300 3620 3420 3653
rect 3460 3620 3570 3653
rect 250 1060 310 2950
rect 3690 1060 3750 2950
rect 420 347 540 380
rect 580 347 700 380
rect 740 347 860 380
rect 900 347 1020 380
rect 1060 347 1180 380
rect 2820 347 2940 380
rect 2980 347 3100 380
rect 3140 347 3260 380
rect 3300 347 3420 380
rect 3460 347 3570 380
rect 420 280 540 347
rect 580 280 700 347
rect 740 280 860 347
rect 900 280 1020 347
rect 1060 280 1180 347
rect 2820 280 2940 347
rect 2980 280 3100 347
rect 3140 280 3260 347
rect 3300 280 3420 347
rect 3460 280 3570 347
<< metal1 >>
rect 0 3980 880 4000
rect 0 3780 20 3980
rect 220 3780 340 3980
rect 540 3780 660 3980
rect 860 3970 880 3980
rect 1360 3980 2640 4000
rect 860 3790 1200 3970
rect 860 3780 880 3790
rect 0 3760 880 3780
rect 0 3660 240 3760
rect 910 3730 1200 3790
rect 1360 3780 1380 3980
rect 1580 3780 1610 3980
rect 1810 3780 1840 3980
rect 2160 3780 2190 3980
rect 2390 3780 2420 3980
rect 2620 3780 2640 3980
rect 3120 3980 4000 4000
rect 3120 3960 3140 3980
rect 1360 3760 2640 3780
rect 2800 3780 3140 3960
rect 3340 3780 3460 3980
rect 3660 3780 3780 3980
rect 3980 3780 4000 3980
rect 0 3460 20 3660
rect 220 3460 240 3660
rect 0 3340 240 3460
rect 0 3140 20 3340
rect 220 3140 240 3340
rect 0 3120 240 3140
rect 360 3720 1200 3730
rect 360 3620 420 3720
rect 540 3620 580 3720
rect 700 3620 740 3720
rect 860 3620 900 3720
rect 1020 3620 1060 3720
rect 1180 3690 1200 3720
rect 1180 3660 1870 3690
rect 1180 3620 1200 3660
rect 1900 3630 2100 3760
rect 2800 3730 3090 3780
rect 3120 3760 4000 3780
rect 2800 3720 3640 3730
rect 2800 3690 2820 3720
rect 2140 3660 2820 3690
rect 360 3600 1200 3620
rect 1230 3600 2770 3630
rect 2800 3620 2820 3660
rect 2940 3620 2980 3720
rect 3100 3620 3140 3720
rect 3260 3620 3300 3720
rect 3420 3620 3460 3720
rect 3570 3620 3640 3720
rect 2800 3600 3640 3620
rect 360 3030 390 3600
rect 240 2950 390 3000
rect 240 2640 250 2950
rect 0 2620 250 2640
rect 0 2480 20 2620
rect 160 2480 250 2620
rect 0 2450 250 2480
rect 0 2310 20 2450
rect 160 2310 250 2450
rect 0 2280 250 2310
rect 0 2140 20 2280
rect 160 2140 250 2280
rect 0 2090 250 2140
rect 0 1910 30 2090
rect 160 1910 250 2090
rect 0 1860 250 1910
rect 0 1720 20 1860
rect 160 1720 250 1860
rect 0 1690 250 1720
rect 0 1550 20 1690
rect 160 1550 250 1690
rect 0 1520 250 1550
rect 0 1380 20 1520
rect 160 1380 250 1520
rect 0 1360 250 1380
rect 240 1060 250 1360
rect 310 2060 390 2950
rect 420 2060 450 3570
rect 480 2090 510 3600
rect 540 2060 570 3570
rect 600 2090 630 3600
rect 660 2060 690 3570
rect 720 2090 750 3600
rect 780 2060 810 3570
rect 840 2090 870 3600
rect 900 2060 930 3570
rect 960 2090 990 3600
rect 1080 3570 1200 3600
rect 1020 2060 1050 3570
rect 1080 3540 1870 3570
rect 1080 3450 1200 3540
rect 1900 3510 2100 3600
rect 2800 3570 2920 3600
rect 2130 3540 2920 3570
rect 1230 3480 2770 3510
rect 1080 3420 1870 3450
rect 1080 3330 1200 3420
rect 1900 3390 2100 3480
rect 2800 3450 2920 3540
rect 2130 3420 2920 3450
rect 1230 3360 2770 3390
rect 1080 3300 1870 3330
rect 1080 3210 1200 3300
rect 1900 3270 2100 3360
rect 2800 3330 2920 3420
rect 2130 3300 2920 3330
rect 1230 3240 2770 3270
rect 1080 3180 1870 3210
rect 1080 3090 1200 3180
rect 1900 3150 2100 3240
rect 2800 3210 2920 3300
rect 2130 3180 2920 3210
rect 1230 3120 2770 3150
rect 1080 3060 1870 3090
rect 1080 2970 1200 3060
rect 1900 3030 2100 3120
rect 2800 3090 2920 3180
rect 2130 3060 2920 3090
rect 1230 3000 2770 3030
rect 1080 2940 1870 2970
rect 1080 2850 1200 2940
rect 1900 2910 2100 3000
rect 2800 2970 2920 3060
rect 2130 2940 2920 2970
rect 1230 2880 2770 2910
rect 1080 2820 1870 2850
rect 1080 2730 1200 2820
rect 1900 2790 2100 2880
rect 2800 2850 2920 2940
rect 2130 2820 2920 2850
rect 1230 2760 2770 2790
rect 1080 2700 1870 2730
rect 1080 2610 1200 2700
rect 1900 2670 2100 2760
rect 2800 2730 2920 2820
rect 2130 2700 2920 2730
rect 1230 2640 2770 2670
rect 1080 2580 1870 2610
rect 1080 2490 1200 2580
rect 1900 2550 2100 2640
rect 2800 2610 2920 2700
rect 2130 2580 2920 2610
rect 1230 2520 2770 2550
rect 1080 2460 1870 2490
rect 1080 2370 1200 2460
rect 1900 2430 2100 2520
rect 2800 2490 2920 2580
rect 2130 2460 2920 2490
rect 1230 2400 2770 2430
rect 1080 2340 1870 2370
rect 1080 2250 1200 2340
rect 1900 2310 2100 2400
rect 2800 2370 2920 2460
rect 2130 2340 2920 2370
rect 1230 2280 2770 2310
rect 1080 2220 1870 2250
rect 1080 2130 1200 2220
rect 1900 2190 2100 2280
rect 2800 2250 2920 2340
rect 2130 2220 2920 2250
rect 1230 2160 2770 2190
rect 1080 2090 1870 2130
rect 1900 2060 2100 2160
rect 2800 2130 2920 2220
rect 2130 2090 2920 2130
rect 2950 2060 2980 3570
rect 3010 2090 3040 3600
rect 3070 2060 3100 3570
rect 3130 2090 3160 3600
rect 3190 2060 3220 3570
rect 3250 2090 3280 3600
rect 3310 2060 3340 3570
rect 3370 2090 3400 3600
rect 3430 2060 3460 3570
rect 3490 2090 3520 3600
rect 3550 2060 3580 3570
rect 3610 3030 3640 3600
rect 3760 3660 4000 3760
rect 3760 3460 3780 3660
rect 3980 3460 4000 3660
rect 3760 3340 4000 3460
rect 3760 3140 3780 3340
rect 3980 3140 4000 3340
rect 3760 3120 4000 3140
rect 3610 2950 3760 3000
rect 3610 2060 3690 2950
rect 310 1940 3690 2060
rect 310 1060 390 1940
rect 240 1010 390 1060
rect 0 860 240 880
rect 0 660 20 860
rect 220 660 240 860
rect 0 540 240 660
rect 0 340 20 540
rect 220 340 240 540
rect 0 240 240 340
rect 360 400 390 980
rect 420 430 450 1940
rect 480 400 510 1910
rect 540 430 570 1940
rect 600 400 630 1910
rect 660 430 690 1940
rect 720 400 750 1910
rect 780 430 810 1940
rect 840 400 870 1910
rect 900 430 930 1940
rect 960 400 990 1910
rect 1020 430 1050 1940
rect 1080 1870 1870 1910
rect 1080 1780 1200 1870
rect 1900 1840 2100 1940
rect 2130 1870 2920 1910
rect 1230 1810 2770 1840
rect 1080 1750 1870 1780
rect 1080 1660 1200 1750
rect 1900 1720 2100 1810
rect 2800 1780 2920 1870
rect 2130 1750 2920 1780
rect 1230 1690 2770 1720
rect 1080 1630 1870 1660
rect 1080 1540 1200 1630
rect 1900 1600 2100 1690
rect 2800 1660 2920 1750
rect 2130 1630 2920 1660
rect 1230 1570 2770 1600
rect 1080 1510 1870 1540
rect 1080 1420 1200 1510
rect 1900 1480 2100 1570
rect 2800 1540 2920 1630
rect 2130 1510 2920 1540
rect 1230 1450 2770 1480
rect 1080 1390 1870 1420
rect 1080 1300 1200 1390
rect 1900 1360 2100 1450
rect 2800 1420 2920 1510
rect 2130 1390 2920 1420
rect 1230 1330 2770 1360
rect 1080 1270 1870 1300
rect 1080 1180 1200 1270
rect 1900 1240 2100 1330
rect 2800 1300 2920 1390
rect 2130 1270 2920 1300
rect 1230 1210 2770 1240
rect 1080 1150 1870 1180
rect 1080 1060 1200 1150
rect 1900 1120 2100 1210
rect 2800 1180 2920 1270
rect 2130 1150 2920 1180
rect 1230 1090 2770 1120
rect 1080 1030 1870 1060
rect 1080 940 1200 1030
rect 1900 1000 2100 1090
rect 2800 1060 2920 1150
rect 2130 1030 2920 1060
rect 1230 970 2770 1000
rect 1080 910 1870 940
rect 1080 820 1200 910
rect 1900 880 2100 970
rect 2800 940 2920 1030
rect 2130 910 2920 940
rect 1230 850 2770 880
rect 1080 790 1870 820
rect 1080 700 1200 790
rect 1900 760 2100 850
rect 2800 820 2920 910
rect 2130 790 2920 820
rect 1230 730 2770 760
rect 1080 670 1870 700
rect 1080 580 1200 670
rect 1900 640 2100 730
rect 2800 700 2920 790
rect 2130 670 2920 700
rect 1230 610 2770 640
rect 1080 550 1870 580
rect 1080 460 1200 550
rect 1900 520 2100 610
rect 2800 580 2920 670
rect 2130 550 2920 580
rect 1230 490 2770 520
rect 1080 430 1870 460
rect 1080 400 1200 430
rect 1900 400 2100 490
rect 2800 460 2920 550
rect 2130 430 2920 460
rect 2950 430 2980 1940
rect 2800 400 2920 430
rect 3010 400 3040 1910
rect 3070 430 3100 1940
rect 3130 400 3160 1910
rect 3190 430 3220 1940
rect 3250 400 3280 1910
rect 3310 430 3340 1940
rect 3370 400 3400 1910
rect 3430 430 3460 1940
rect 3490 400 3520 1910
rect 3550 430 3580 1940
rect 3610 1060 3690 1940
rect 3750 2640 3760 2950
rect 3750 2620 4000 2640
rect 3750 2480 3840 2620
rect 3980 2480 4000 2620
rect 3750 2450 4000 2480
rect 3750 2310 3840 2450
rect 3980 2310 4000 2450
rect 3750 2280 4000 2310
rect 3750 2140 3840 2280
rect 3980 2140 4000 2280
rect 3750 2090 4000 2140
rect 3750 1910 3840 2090
rect 3970 1910 4000 2090
rect 3750 1860 4000 1910
rect 3750 1720 3840 1860
rect 3980 1720 4000 1860
rect 3750 1690 4000 1720
rect 3750 1550 3840 1690
rect 3980 1550 4000 1690
rect 3750 1520 4000 1550
rect 3750 1380 3840 1520
rect 3980 1380 4000 1520
rect 3750 1360 4000 1380
rect 3750 1060 3760 1360
rect 3610 1010 3760 1060
rect 3610 400 3640 980
rect 360 380 1200 400
rect 360 280 420 380
rect 540 280 580 380
rect 700 280 740 380
rect 860 280 900 380
rect 1020 280 1060 380
rect 1180 340 1200 380
rect 1230 370 2770 400
rect 2800 380 3640 400
rect 1180 310 1870 340
rect 1180 280 1200 310
rect 360 270 1200 280
rect 0 220 880 240
rect 0 20 20 220
rect 220 20 340 220
rect 540 20 660 220
rect 860 210 880 220
rect 910 210 1200 270
rect 1900 240 2100 370
rect 2800 340 2820 380
rect 2130 310 2820 340
rect 2800 280 2820 310
rect 2940 280 2980 380
rect 3100 280 3140 380
rect 3260 280 3300 380
rect 3420 280 3460 380
rect 3570 280 3640 380
rect 2800 270 3640 280
rect 3760 860 4000 880
rect 3760 660 3780 860
rect 3980 660 4000 860
rect 3760 540 4000 660
rect 3760 340 3780 540
rect 3980 340 4000 540
rect 860 30 1200 210
rect 1360 220 2640 240
rect 860 20 880 30
rect 0 0 880 20
rect 1360 20 1380 220
rect 1580 20 1600 220
rect 1800 20 1830 220
rect 2150 20 2190 220
rect 2390 20 2420 220
rect 2620 20 2640 220
rect 2800 210 3090 270
rect 3760 240 4000 340
rect 3120 220 4000 240
rect 3120 210 3140 220
rect 2800 30 3140 210
rect 1360 0 2640 20
rect 3120 20 3140 30
rect 3340 20 3460 220
rect 3660 20 3780 220
rect 3980 20 4000 220
rect 3120 0 4000 20
<< via1 >>
rect 20 3780 220 3980
rect 340 3780 540 3980
rect 660 3780 860 3980
rect 1380 3780 1580 3980
rect 1610 3780 1810 3980
rect 1840 3780 2160 3980
rect 2190 3780 2390 3980
rect 2420 3780 2620 3980
rect 3140 3780 3340 3980
rect 3460 3780 3660 3980
rect 3780 3780 3980 3980
rect 20 3460 220 3660
rect 20 3140 220 3340
rect 20 2480 160 2620
rect 20 2310 160 2450
rect 20 2140 160 2280
rect 20 1720 160 1860
rect 20 1550 160 1690
rect 20 1380 160 1520
rect 3780 3460 3980 3660
rect 3780 3140 3980 3340
rect 20 660 220 860
rect 20 340 220 540
rect 3840 2480 3980 2620
rect 3840 2310 3980 2450
rect 3840 2140 3980 2280
rect 3840 1720 3980 1860
rect 3840 1550 3980 1690
rect 3840 1380 3980 1520
rect 20 20 220 220
rect 340 20 540 220
rect 660 20 860 220
rect 3780 660 3980 860
rect 3780 340 3980 540
rect 1380 20 1580 220
rect 1600 20 1800 220
rect 1830 20 2150 220
rect 2190 20 2390 220
rect 2420 20 2620 220
rect 3140 20 3340 220
rect 3460 20 3660 220
rect 3780 20 3980 220
<< metal2 >>
rect 0 3980 880 4000
rect 0 3780 20 3980
rect 220 3780 340 3980
rect 540 3780 660 3980
rect 860 3780 880 3980
rect 1360 3980 2640 4000
rect 1360 3820 1380 3980
rect 0 3760 880 3780
rect 980 3780 1380 3820
rect 1580 3780 1610 3980
rect 1810 3780 1840 3980
rect 2160 3780 2190 3980
rect 2390 3780 2420 3980
rect 2620 3820 2640 3980
rect 3120 3980 4000 4000
rect 2620 3780 3020 3820
rect 0 3660 242 3760
rect 980 3720 3020 3780
rect 3120 3780 3140 3980
rect 3340 3780 3460 3980
rect 3660 3780 3780 3980
rect 3980 3780 4000 3980
rect 3120 3760 4000 3780
rect 0 3460 20 3660
rect 220 3570 242 3660
rect 360 3710 3640 3720
rect 360 3600 1120 3710
rect 220 3540 1030 3570
rect 220 3460 320 3540
rect 1060 3510 1120 3600
rect 350 3480 1120 3510
rect 0 3450 320 3460
rect 0 3420 1030 3450
rect 0 3340 320 3420
rect 1060 3390 1120 3480
rect 350 3360 1120 3390
rect 0 3140 20 3340
rect 220 3330 320 3340
rect 220 3300 1030 3330
rect 220 3210 320 3300
rect 1060 3270 1120 3360
rect 350 3240 1120 3270
rect 220 3180 1030 3210
rect 220 3140 320 3180
rect 1060 3150 1120 3240
rect 0 3120 320 3140
rect 350 3120 1120 3150
rect 240 3090 320 3120
rect 240 3060 1030 3090
rect 240 2970 320 3060
rect 1060 3030 1120 3120
rect 350 3000 1120 3030
rect 240 2940 1030 2970
rect 240 2850 320 2940
rect 1060 2910 1120 3000
rect 350 2880 1120 2910
rect 240 2820 1030 2850
rect 240 2730 320 2820
rect 1060 2790 1120 2880
rect 350 2760 1120 2790
rect 240 2700 1030 2730
rect 0 2620 180 2640
rect 0 2480 20 2620
rect 160 2480 180 2620
rect 0 2450 180 2480
rect 0 2310 20 2450
rect 160 2310 180 2450
rect 0 2280 180 2310
rect 0 2140 20 2280
rect 160 2140 180 2280
rect 0 1860 180 2140
rect 0 1720 20 1860
rect 160 1720 180 1860
rect 0 1690 180 1720
rect 0 1550 20 1690
rect 160 1550 180 1690
rect 0 1520 180 1550
rect 0 1380 20 1520
rect 160 1380 180 1520
rect 0 1360 180 1380
rect 240 2610 320 2700
rect 1060 2670 1120 2760
rect 350 2640 1120 2670
rect 240 2580 1030 2610
rect 240 2490 320 2580
rect 1060 2550 1120 2640
rect 350 2520 1120 2550
rect 240 2460 1030 2490
rect 240 2370 320 2460
rect 1060 2430 1120 2520
rect 350 2400 1120 2430
rect 240 2340 1030 2370
rect 240 2250 320 2340
rect 1060 2310 1120 2400
rect 350 2280 1120 2310
rect 240 2220 1030 2250
rect 240 2130 320 2220
rect 1060 2190 1120 2280
rect 350 2160 1120 2190
rect 240 2100 1030 2130
rect 240 2040 320 2100
rect 1060 2070 1120 2160
rect 1150 2040 1180 3680
rect 1210 2070 1240 3710
rect 1270 2040 1300 3680
rect 1330 2070 1360 3710
rect 1390 2040 1420 3680
rect 1450 2070 1480 3710
rect 1510 2040 1540 3680
rect 1570 2070 1600 3710
rect 1630 2040 1660 3680
rect 1690 2070 1720 3710
rect 1750 2040 1780 3680
rect 1810 2070 1840 3710
rect 1870 2040 1900 3680
rect 240 1960 1900 2040
rect 240 1900 320 1960
rect 240 1870 1030 1900
rect 240 1780 320 1870
rect 1060 1840 1120 1930
rect 350 1810 1120 1840
rect 240 1750 1030 1780
rect 240 1660 320 1750
rect 1060 1720 1120 1810
rect 350 1690 1120 1720
rect 240 1630 1030 1660
rect 240 1540 320 1630
rect 1060 1600 1120 1690
rect 350 1570 1120 1600
rect 240 1510 1030 1540
rect 240 1420 320 1510
rect 1060 1480 1120 1570
rect 350 1450 1120 1480
rect 240 1390 1030 1420
rect 240 1300 320 1390
rect 1060 1360 1120 1450
rect 350 1330 1120 1360
rect 240 1270 1030 1300
rect 240 1180 320 1270
rect 1060 1240 1120 1330
rect 350 1210 1120 1240
rect 240 1150 1030 1180
rect 240 1060 320 1150
rect 1060 1120 1120 1210
rect 350 1090 1120 1120
rect 240 1030 1030 1060
rect 240 940 320 1030
rect 1060 1000 1120 1090
rect 350 970 1120 1000
rect 240 910 1030 940
rect 240 880 320 910
rect 1060 880 1120 970
rect 0 860 320 880
rect 0 660 20 860
rect 220 820 320 860
rect 350 850 1120 880
rect 220 790 1030 820
rect 220 700 320 790
rect 1060 760 1120 850
rect 350 730 1120 760
rect 220 670 1030 700
rect 220 660 320 670
rect 0 580 320 660
rect 1060 640 1120 730
rect 350 610 1120 640
rect 0 550 1030 580
rect 0 540 320 550
rect 0 340 20 540
rect 220 460 320 540
rect 1060 520 1120 610
rect 350 490 1120 520
rect 220 430 1030 460
rect 220 340 240 430
rect 1060 400 1120 490
rect 0 240 240 340
rect 360 290 1120 400
rect 1150 320 1180 1960
rect 1210 290 1240 1930
rect 1270 320 1300 1960
rect 1330 290 1360 1930
rect 1390 320 1420 1960
rect 1450 290 1480 1930
rect 1510 320 1540 1960
rect 1570 290 1600 1930
rect 1630 320 1660 1960
rect 1690 290 1720 1930
rect 1750 320 1780 1960
rect 1810 290 1840 1930
rect 1870 320 1900 1960
rect 1930 290 2070 3710
rect 2100 2040 2130 3680
rect 2160 2070 2190 3710
rect 2220 2040 2250 3680
rect 2280 2070 2310 3710
rect 2340 2040 2370 3680
rect 2400 2070 2430 3710
rect 2460 2040 2490 3680
rect 2520 2070 2550 3710
rect 2580 2040 2610 3680
rect 2640 2070 2670 3710
rect 2700 2040 2730 3680
rect 2760 2070 2790 3710
rect 2820 2040 2850 3680
rect 2880 3600 3640 3710
rect 3760 3660 4000 3760
rect 2880 3510 2940 3600
rect 3760 3570 3780 3660
rect 2970 3540 3780 3570
rect 2880 3480 3650 3510
rect 2880 3390 2940 3480
rect 3680 3460 3780 3540
rect 3980 3460 4000 3660
rect 3680 3450 4000 3460
rect 2970 3420 4000 3450
rect 2880 3360 3650 3390
rect 2880 3270 2940 3360
rect 3680 3340 4000 3420
rect 3680 3330 3780 3340
rect 2970 3300 3780 3330
rect 2880 3240 3650 3270
rect 2880 3150 2940 3240
rect 3680 3210 3780 3300
rect 2970 3180 3780 3210
rect 2880 3120 3650 3150
rect 3680 3140 3780 3180
rect 3980 3140 4000 3340
rect 3680 3120 4000 3140
rect 2880 3030 2940 3120
rect 3680 3090 3760 3120
rect 2970 3060 3760 3090
rect 2880 3000 3650 3030
rect 2880 2910 2940 3000
rect 3680 2970 3760 3060
rect 2970 2940 3760 2970
rect 2880 2880 3650 2910
rect 2880 2790 2940 2880
rect 3680 2850 3760 2940
rect 2970 2820 3760 2850
rect 2880 2760 3650 2790
rect 2880 2670 2940 2760
rect 3680 2730 3760 2820
rect 2970 2700 3760 2730
rect 2880 2640 3650 2670
rect 2880 2550 2940 2640
rect 3680 2610 3760 2700
rect 2970 2580 3760 2610
rect 2880 2520 3650 2550
rect 2880 2430 2940 2520
rect 3680 2490 3760 2580
rect 2970 2460 3760 2490
rect 2880 2400 3650 2430
rect 2880 2310 2940 2400
rect 3680 2370 3760 2460
rect 2970 2340 3760 2370
rect 2880 2280 3650 2310
rect 2880 2190 2940 2280
rect 3680 2250 3760 2340
rect 2970 2220 3760 2250
rect 2880 2160 3650 2190
rect 2880 2070 2940 2160
rect 3680 2130 3760 2220
rect 2970 2100 3760 2130
rect 3680 2040 3760 2100
rect 2100 1960 3760 2040
rect 2100 320 2130 1960
rect 2160 290 2190 1930
rect 2220 320 2250 1960
rect 2280 290 2310 1930
rect 2340 320 2370 1960
rect 2400 290 2430 1930
rect 2460 320 2490 1960
rect 2520 290 2550 1930
rect 2580 320 2610 1960
rect 2640 290 2670 1930
rect 2700 320 2730 1960
rect 2760 290 2790 1930
rect 2820 320 2850 1960
rect 2880 1840 2940 1930
rect 3680 1900 3760 1960
rect 2970 1870 3760 1900
rect 2880 1810 3650 1840
rect 2880 1720 2940 1810
rect 3680 1780 3760 1870
rect 2970 1750 3760 1780
rect 2880 1690 3650 1720
rect 2880 1600 2940 1690
rect 3680 1660 3760 1750
rect 2970 1630 3760 1660
rect 2880 1570 3650 1600
rect 2880 1480 2940 1570
rect 3680 1540 3760 1630
rect 2970 1510 3760 1540
rect 2880 1450 3650 1480
rect 2880 1360 2940 1450
rect 3680 1420 3760 1510
rect 2970 1390 3760 1420
rect 2880 1330 3650 1360
rect 2880 1240 2940 1330
rect 3680 1300 3760 1390
rect 3820 2620 4000 2640
rect 3820 2480 3840 2620
rect 3980 2480 4000 2620
rect 3820 2450 4000 2480
rect 3820 2310 3840 2450
rect 3980 2310 4000 2450
rect 3820 2280 4000 2310
rect 3820 2140 3840 2280
rect 3980 2140 4000 2280
rect 3820 1860 4000 2140
rect 3820 1720 3840 1860
rect 3980 1720 4000 1860
rect 3820 1690 4000 1720
rect 3820 1550 3840 1690
rect 3980 1550 4000 1690
rect 3820 1520 4000 1550
rect 3820 1380 3840 1520
rect 3980 1380 4000 1520
rect 3820 1360 4000 1380
rect 2970 1270 3760 1300
rect 2880 1210 3650 1240
rect 2880 1120 2940 1210
rect 3680 1180 3760 1270
rect 2970 1150 3760 1180
rect 2880 1090 3650 1120
rect 2880 1000 2940 1090
rect 3680 1060 3760 1150
rect 2970 1030 3760 1060
rect 2880 970 3650 1000
rect 2880 880 2940 970
rect 3680 940 3760 1030
rect 2970 910 3760 940
rect 3680 880 3760 910
rect 2880 850 3650 880
rect 3680 860 4000 880
rect 2880 760 2940 850
rect 3680 820 3780 860
rect 2970 790 3780 820
rect 2880 730 3650 760
rect 2880 640 2940 730
rect 3680 700 3780 790
rect 2970 670 3780 700
rect 3680 660 3780 670
rect 3980 660 4000 860
rect 2880 610 3650 640
rect 2880 520 2940 610
rect 3680 580 4000 660
rect 2970 550 4000 580
rect 3680 540 4000 550
rect 2880 490 3650 520
rect 2880 400 2940 490
rect 3680 460 3780 540
rect 2970 430 3780 460
rect 2880 290 3640 400
rect 360 280 3640 290
rect 3760 340 3780 430
rect 3980 340 4000 540
rect 0 220 880 240
rect 0 20 20 220
rect 220 20 340 220
rect 540 20 660 220
rect 860 20 880 220
rect 980 220 3020 280
rect 3760 240 4000 340
rect 980 180 1380 220
rect 0 0 880 20
rect 1360 20 1380 180
rect 1580 20 1600 220
rect 1800 20 1830 220
rect 2150 20 2190 220
rect 2390 20 2420 220
rect 2620 180 3020 220
rect 3120 220 4000 240
rect 2620 20 2640 180
rect 1360 0 2640 20
rect 3120 20 3140 220
rect 3340 20 3460 220
rect 3660 20 3780 220
rect 3980 20 4000 220
rect 3120 0 4000 20
<< metal3 >>
rect 0 3980 880 4000
rect 0 3810 20 3980
rect 190 3810 210 3980
rect 380 3810 500 3980
rect 670 3810 690 3980
rect 860 3810 880 3980
rect 1360 3980 2640 4000
rect 1360 3850 1380 3980
rect 1510 3850 1540 3980
rect 1670 3850 1700 3980
rect 1830 3850 2170 3980
rect 2300 3850 2330 3980
rect 2460 3850 2490 3980
rect 2620 3850 2640 3980
rect 1360 3830 2640 3850
rect 3120 3980 4000 4000
rect 0 3790 880 3810
rect 0 3620 20 3790
rect 190 3750 880 3790
rect 3120 3810 3140 3980
rect 3310 3810 3330 3980
rect 3500 3810 3620 3980
rect 3790 3810 3810 3980
rect 3980 3810 4000 3980
rect 3120 3790 4000 3810
rect 3120 3750 3810 3790
rect 190 3620 3810 3750
rect 3980 3620 4000 3790
rect 0 3500 4000 3620
rect 0 3330 20 3500
rect 190 3330 3810 3500
rect 3980 3330 4000 3500
rect 0 3310 4000 3330
rect 0 3140 20 3310
rect 190 3140 3810 3310
rect 3980 3140 4000 3310
rect 0 3120 4000 3140
rect 0 2620 170 2640
rect 0 2490 20 2620
rect 150 2490 170 2620
rect 0 2460 170 2490
rect 0 2330 20 2460
rect 150 2330 170 2460
rect 0 2300 170 2330
rect 0 2170 20 2300
rect 150 2170 170 2300
rect 0 1830 170 2170
rect 0 1700 20 1830
rect 150 1700 170 1830
rect 0 1670 170 1700
rect 0 1540 20 1670
rect 150 1540 170 1670
rect 0 1510 170 1540
rect 0 1380 20 1510
rect 150 1380 170 1510
rect 0 1360 170 1380
rect 250 880 3750 3120
rect 3830 2620 4000 2640
rect 3830 2490 3850 2620
rect 3980 2490 4000 2620
rect 3830 2460 4000 2490
rect 3830 2330 3850 2460
rect 3980 2330 4000 2460
rect 3830 2300 4000 2330
rect 3830 2170 3850 2300
rect 3980 2170 4000 2300
rect 3830 1830 4000 2170
rect 3830 1700 3850 1830
rect 3980 1700 4000 1830
rect 3830 1670 4000 1700
rect 3830 1540 3850 1670
rect 3980 1540 4000 1670
rect 3830 1510 4000 1540
rect 3830 1380 3850 1510
rect 3980 1380 4000 1510
rect 3830 1360 4000 1380
rect 0 860 4000 880
rect 0 690 20 860
rect 190 690 3810 860
rect 3980 690 4000 860
rect 0 670 4000 690
rect 0 500 20 670
rect 190 500 3810 670
rect 3980 500 4000 670
rect 0 380 4000 500
rect 0 210 20 380
rect 190 250 3810 380
rect 190 210 880 250
rect 0 190 880 210
rect 0 20 20 190
rect 190 20 210 190
rect 380 20 500 190
rect 670 20 690 190
rect 860 20 880 190
rect 3120 210 3810 250
rect 3980 210 4000 380
rect 3120 190 4000 210
rect 0 0 880 20
rect 1360 150 2640 170
rect 1360 20 1380 150
rect 1510 20 1540 150
rect 1670 20 1700 150
rect 1830 20 2170 150
rect 2300 20 2330 150
rect 2460 20 2490 150
rect 2620 20 2640 150
rect 1360 0 2640 20
rect 3120 20 3140 190
rect 3310 20 3330 190
rect 3500 20 3620 190
rect 3790 20 3810 190
rect 3980 20 4000 190
rect 3120 0 4000 20
<< via3 >>
rect 20 3810 190 3980
rect 210 3810 380 3980
rect 500 3810 670 3980
rect 690 3810 860 3980
rect 1380 3850 1510 3980
rect 1540 3850 1670 3980
rect 1700 3850 1830 3980
rect 2170 3850 2300 3980
rect 2330 3850 2460 3980
rect 2490 3850 2620 3980
rect 20 3620 190 3790
rect 3140 3810 3310 3980
rect 3330 3810 3500 3980
rect 3620 3810 3790 3980
rect 3810 3810 3980 3980
rect 3810 3620 3980 3790
rect 20 3330 190 3500
rect 3810 3330 3980 3500
rect 20 3140 190 3310
rect 3810 3140 3980 3310
rect 20 2490 150 2620
rect 20 2330 150 2460
rect 20 2170 150 2300
rect 20 1700 150 1830
rect 20 1540 150 1670
rect 20 1380 150 1510
rect 3850 2490 3980 2620
rect 3850 2330 3980 2460
rect 3850 2170 3980 2300
rect 3850 1700 3980 1830
rect 3850 1540 3980 1670
rect 3850 1380 3980 1510
rect 20 690 190 860
rect 3810 690 3980 860
rect 20 500 190 670
rect 3810 500 3980 670
rect 20 210 190 380
rect 20 20 190 190
rect 210 20 380 190
rect 500 20 670 190
rect 690 20 860 190
rect 3810 210 3980 380
rect 1380 20 1510 150
rect 1540 20 1670 150
rect 1700 20 1830 150
rect 2170 20 2300 150
rect 2330 20 2460 150
rect 2490 20 2620 150
rect 3140 20 3310 190
rect 3330 20 3500 190
rect 3620 20 3790 190
rect 3810 20 3980 190
<< mimcap >>
rect 280 3690 3720 3720
rect 280 310 310 3690
rect 3690 310 3720 3690
rect 280 280 3720 310
<< mimcapcontact >>
rect 310 310 3690 3690
<< metal4 >>
rect 0 3980 880 4000
rect 0 3810 20 3980
rect 190 3810 210 3980
rect 380 3810 500 3980
rect 670 3810 690 3980
rect 860 3810 880 3980
rect 0 3790 880 3810
rect 1360 3980 2640 4000
rect 1360 3850 1380 3980
rect 1510 3850 1540 3980
rect 1670 3850 1700 3980
rect 1830 3850 2170 3980
rect 2300 3850 2330 3980
rect 2460 3850 2490 3980
rect 2620 3850 2640 3980
rect 0 3620 20 3790
rect 190 3620 210 3790
rect 1360 3710 2640 3850
rect 3120 3980 4000 4000
rect 3120 3810 3140 3980
rect 3310 3810 3330 3980
rect 3500 3810 3620 3980
rect 3790 3810 3810 3980
rect 3980 3810 4000 3980
rect 3120 3790 4000 3810
rect 0 3500 210 3620
rect 0 3330 20 3500
rect 190 3330 210 3500
rect 0 3310 210 3330
rect 0 3140 20 3310
rect 190 3140 210 3310
rect 0 3120 210 3140
rect 290 3690 3710 3710
rect 290 2640 310 3690
rect 0 2620 310 2640
rect 0 2490 20 2620
rect 150 2490 310 2620
rect 0 2460 310 2490
rect 0 2330 20 2460
rect 150 2330 310 2460
rect 0 2300 310 2330
rect 0 2170 20 2300
rect 150 2170 310 2300
rect 0 1830 310 2170
rect 0 1700 20 1830
rect 150 1700 310 1830
rect 0 1670 310 1700
rect 0 1540 20 1670
rect 150 1540 310 1670
rect 0 1510 310 1540
rect 0 1380 20 1510
rect 150 1380 310 1510
rect 0 1360 310 1380
rect 0 860 210 880
rect 0 690 20 860
rect 190 690 210 860
rect 0 670 210 690
rect 0 500 20 670
rect 190 500 210 670
rect 0 380 210 500
rect 0 210 20 380
rect 190 210 210 380
rect 290 310 310 1360
rect 3690 2640 3710 3690
rect 3790 3620 3810 3790
rect 3980 3620 4000 3790
rect 3790 3500 4000 3620
rect 3790 3330 3810 3500
rect 3980 3330 4000 3500
rect 3790 3310 4000 3330
rect 3790 3140 3810 3310
rect 3980 3140 4000 3310
rect 3790 3120 4000 3140
rect 3690 2620 4000 2640
rect 3690 2490 3850 2620
rect 3980 2490 4000 2620
rect 3690 2460 4000 2490
rect 3690 2330 3850 2460
rect 3980 2330 4000 2460
rect 3690 2300 4000 2330
rect 3690 2170 3850 2300
rect 3980 2170 4000 2300
rect 3690 1830 4000 2170
rect 3690 1700 3850 1830
rect 3980 1700 4000 1830
rect 3690 1670 4000 1700
rect 3690 1540 3850 1670
rect 3980 1540 4000 1670
rect 3690 1510 4000 1540
rect 3690 1380 3850 1510
rect 3980 1380 4000 1510
rect 3690 1360 4000 1380
rect 3690 310 3710 1360
rect 290 290 3710 310
rect 3790 860 4000 880
rect 3790 690 3810 860
rect 3980 690 4000 860
rect 3790 670 4000 690
rect 3790 500 3810 670
rect 3980 500 4000 670
rect 3790 380 4000 500
rect 0 190 880 210
rect 0 20 20 190
rect 190 20 210 190
rect 380 20 500 190
rect 670 20 690 190
rect 860 20 880 190
rect 0 0 880 20
rect 1360 150 2640 290
rect 3790 210 3810 380
rect 3980 210 4000 380
rect 1360 20 1380 150
rect 1510 20 1540 150
rect 1670 20 1700 150
rect 1830 20 2170 150
rect 2300 20 2330 150
rect 2460 20 2490 150
rect 2620 20 2640 150
rect 1360 0 2640 20
rect 3120 190 4000 210
rect 3120 20 3140 190
rect 3310 20 3330 190
rect 3500 20 3620 190
rect 3790 20 3810 190
rect 3980 20 4000 190
rect 3120 0 4000 20
<< labels >>
flabel metal1 s 1360 0 2640 180 5 FreeSans 320 0 0 0 nmoscap_top
port 1 s
flabel metal1 s 1360 3820 2640 4000 1 FreeSans 320 0 0 0 nmoscap_top
port 1 n
flabel metal1 s 3974 1360 4000 2640 3 FreeSans 320 90 0 0 nmoscap_top
port 1 e
flabel metal1 s 0 1360 26 2640 7 FreeSans 320 90 0 0 nmoscap_top
port 1 w
flabel metal1 s 0 3120 240 4000 7 FreeSans 320 90 0 0 nmoscap_bot
port 2 w
flabel metal1 s 0 0 240 880 7 FreeSans 320 90 0 0 nmoscap_bot
port 2 w
flabel metal1 s 3760 0 4000 880 3 FreeSans 320 90 0 0 nmoscap_bot
port 2 e
flabel metal1 s 3760 3120 4000 4000 3 FreeSans 320 90 0 0 nmoscap_bot
port 2 e
flabel metal1 s 3120 3760 4000 4000 1 FreeSans 320 0 0 0 nmoscap_bot
port 2 n
flabel metal1 s 0 3760 880 4000 1 FreeSans 320 0 0 0 nmoscap_bot
port 2 n
flabel metal1 s 0 0 880 240 5 FreeSans 320 0 0 0 nmoscap_bot
port 2 s
flabel metal1 s 3120 0 4000 240 5 FreeSans 320 0 0 0 nmoscap_bot
port 2 s
flabel locali s 890 0 1350 80 5 FreeSans 320 0 0 0 pwell
port 3 s
flabel locali s 2650 0 3110 80 5 FreeSans 320 0 0 0 pwell
port 3 s
flabel locali s 2650 3920 3110 4000 1 FreeSans 320 0 0 0 pwell
port 3 n
flabel locali s 890 3920 1350 4000 1 FreeSans 320 0 0 0 pwell
port 3 n
flabel locali s 3920 2650 4000 3110 3 FreeSans 320 90 0 0 pwell
port 3 e
flabel locali s 3920 890 4000 1350 3 FreeSans 320 90 0 0 pwell
port 3 e
flabel locali s 0 890 80 1350 7 FreeSans 320 90 0 0 pwell
port 3 w
flabel locali s 0 2650 80 3110 7 FreeSans 320 90 0 0 pwell
port 3 w
flabel metal4 1360 3830 2640 4000 1 FreeSans 320 0 0 0 mimcap_top
port 4 n
flabel metal4 1360 0 2640 170 5 FreeSans 320 0 0 0 mimcap_top
port 4 s
flabel metal4 3830 1360 4000 2640 3 FreeSans 320 90 0 0 mimcap_top
port 4 e
flabel metal4 0 1360 170 2640 7 FreeSans 320 90 0 0 mimcap_top
port 4 w
flabel metal4 3120 0 4000 210 5 FreeSans 320 0 0 0 mimcap_bot
port 5 s
flabel metal4 0 0 880 210 5 FreeSans 320 0 0 0 mimcap_bot
port 5 s
flabel metal4 0 3790 880 4000 1 FreeSans 320 0 0 0 mimcap_bot
port 5 n
flabel metal4 3120 3790 4000 4000 1 FreeSans 320 0 0 0 mimcap_bot
port 5 n
flabel metal4 3790 3120 4000 4000 3 FreeSans 320 90 0 0 mimcap_bot
port 5 e
flabel metal4 3790 0 4000 880 3 FreeSans 320 90 0 0 mimcap_bot
port 5 e
flabel metal4 0 0 210 880 7 FreeSans 320 90 0 0 mimcap_bot
port 5 w
flabel metal4 0 3120 210 4000 7 FreeSans 320 90 0 0 mimcap_bot
port 5 w
<< properties >>
string FIXED_BBOX 0 0 4000 4000
<< end >>
