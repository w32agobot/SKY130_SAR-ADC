magic
tech sky130A
magscale 1 2
timestamp 1663935273
<< nwell >>
rect 3477 34899 3539 34909
rect 3477 34819 3541 34899
rect 1557 34596 1583 34597
rect 1557 34594 2167 34596
rect 1557 34264 2169 34594
rect 3477 34584 3539 34819
rect 2063 33176 2257 33421
<< psubdiff >>
rect 944 35679 5768 35727
rect 944 35519 1306 35679
rect 1466 35519 1706 35679
rect 1866 35519 2106 35679
rect 2266 35519 2506 35679
rect 2666 35519 2906 35679
rect 3066 35519 3306 35679
rect 3466 35519 3706 35679
rect 3866 35519 4106 35679
rect 4266 35519 4506 35679
rect 4666 35519 4906 35679
rect 5066 35519 5306 35679
rect 5462 35519 5768 35679
rect 944 35496 5768 35519
rect 944 35336 1008 35496
rect 1168 35476 5547 35496
rect 1168 35336 1237 35476
rect 944 35096 1237 35336
rect 944 34936 1008 35096
rect 1168 34936 1237 35096
rect 5479 35336 5547 35476
rect 5707 35476 5768 35496
rect 5707 35336 5767 35476
rect 5479 35096 5767 35336
rect 944 34696 1237 34936
rect 5479 34936 5547 35096
rect 5707 34936 5767 35096
rect 944 34536 1008 34696
rect 1168 34536 1237 34696
rect 944 34296 1237 34536
rect 944 34136 1008 34296
rect 1168 34136 1237 34296
rect 944 33896 1237 34136
rect 944 33736 1008 33896
rect 1168 33736 1237 33896
rect 944 33496 1237 33736
rect 944 33336 1008 33496
rect 1168 33336 1237 33496
rect 944 33096 1237 33336
rect 5479 34696 5767 34936
rect 5479 34536 5547 34696
rect 5707 34536 5767 34696
rect 5479 34296 5767 34536
rect 5479 34136 5547 34296
rect 5707 34136 5767 34296
rect 5479 33896 5767 34136
rect 5479 33736 5547 33896
rect 5707 33736 5767 33896
rect 5479 33496 5767 33736
rect 5479 33336 5547 33496
rect 5707 33336 5767 33496
rect 944 32936 1008 33096
rect 1168 32936 1237 33096
rect 5479 33096 5767 33336
rect 944 32650 1237 32936
rect 5479 32936 5547 33096
rect 5707 32936 5767 33096
rect 5479 32732 5767 32936
rect 5479 32650 5768 32732
rect 944 32649 3138 32650
rect 3285 32649 5768 32650
rect 944 32614 5768 32649
rect 944 32454 1008 32614
rect 1168 32454 1408 32614
rect 1568 32454 1808 32614
rect 1968 32454 2208 32614
rect 2368 32454 2608 32614
rect 2768 32454 3008 32614
rect 3168 32454 3408 32614
rect 3568 32454 3808 32614
rect 3968 32454 4208 32614
rect 4368 32454 4608 32614
rect 4768 32454 5008 32614
rect 5168 32454 5547 32614
rect 5707 32454 5768 32614
rect 944 32449 5768 32454
rect 944 32411 5767 32449
<< psubdiffcont >>
rect 1306 35519 1466 35679
rect 1706 35519 1866 35679
rect 2106 35519 2266 35679
rect 2506 35519 2666 35679
rect 2906 35519 3066 35679
rect 3306 35519 3466 35679
rect 3706 35519 3866 35679
rect 4106 35519 4266 35679
rect 4506 35519 4666 35679
rect 4906 35519 5066 35679
rect 5306 35519 5462 35679
rect 1008 35336 1168 35496
rect 1008 34936 1168 35096
rect 5547 35336 5707 35496
rect 5547 34936 5707 35096
rect 1008 34536 1168 34696
rect 1008 34136 1168 34296
rect 1008 33736 1168 33896
rect 1008 33336 1168 33496
rect 5547 34536 5707 34696
rect 5547 34136 5707 34296
rect 5547 33736 5707 33896
rect 5547 33336 5707 33496
rect 1008 32936 1168 33096
rect 5547 32936 5707 33096
rect 1008 32454 1168 32614
rect 1408 32454 1568 32614
rect 1808 32454 1968 32614
rect 2208 32454 2368 32614
rect 2608 32454 2768 32614
rect 3008 32454 3168 32614
rect 3408 32454 3568 32614
rect 3808 32454 3968 32614
rect 4208 32454 4368 32614
rect 4608 32454 4768 32614
rect 5008 32454 5168 32614
rect 5547 32454 5707 32614
<< poly >>
rect 3485 34981 3551 34994
rect 3485 34966 3501 34981
rect 2639 34964 3501 34966
rect 1752 34947 3501 34964
rect 3535 34947 3551 34981
rect 1752 34934 3551 34947
rect 1652 34870 3565 34892
rect 1652 34862 3521 34870
rect 3511 34836 3521 34862
rect 3555 34836 3565 34870
rect 3511 34820 3565 34836
rect 3544 33172 3612 33182
rect 3544 33144 3562 33172
rect 2244 33138 3562 33144
rect 3596 33138 3612 33172
rect 2244 33114 3612 33138
rect 2244 33040 3569 33070
rect 3500 33038 3569 33040
rect 3500 33003 3516 33038
rect 3553 33003 3569 33038
rect 3500 32992 3569 33003
<< polycont >>
rect 3501 34947 3535 34981
rect 3521 34836 3555 34870
rect 3562 33138 3596 33172
rect 3516 33003 3553 33038
<< locali >>
rect 463 63060 946 63109
rect 463 62984 504 63060
rect 576 62984 626 63060
rect 698 62984 752 63060
rect 824 62984 946 63060
rect 463 62913 946 62984
rect 463 62837 504 62913
rect 576 62837 626 62913
rect 698 62837 752 62913
rect 824 62837 946 62913
rect 463 62776 946 62837
rect 463 62700 504 62776
rect 576 62700 626 62776
rect 698 62700 752 62776
rect 824 62700 946 62776
rect 463 62650 946 62700
rect 463 61300 946 61349
rect 463 61224 504 61300
rect 576 61224 626 61300
rect 698 61224 752 61300
rect 824 61224 946 61300
rect 463 61153 946 61224
rect 463 61077 504 61153
rect 576 61077 626 61153
rect 698 61077 752 61153
rect 824 61077 946 61153
rect 463 61016 946 61077
rect 463 60940 504 61016
rect 576 60940 626 61016
rect 698 60940 752 61016
rect 824 60940 946 61016
rect 463 60890 946 60940
rect 463 59060 946 59109
rect 463 58984 504 59060
rect 576 58984 626 59060
rect 698 58984 752 59060
rect 824 58984 946 59060
rect 463 58913 946 58984
rect 463 58837 504 58913
rect 576 58837 626 58913
rect 698 58837 752 58913
rect 824 58837 946 58913
rect 463 58776 946 58837
rect 463 58700 504 58776
rect 576 58700 626 58776
rect 698 58700 752 58776
rect 824 58700 946 58776
rect 463 58650 946 58700
rect 463 57301 946 57350
rect 463 57225 504 57301
rect 576 57225 626 57301
rect 698 57225 752 57301
rect 824 57225 946 57301
rect 463 57154 946 57225
rect 463 57078 504 57154
rect 576 57078 626 57154
rect 698 57078 752 57154
rect 824 57078 946 57154
rect 463 57017 946 57078
rect 463 56941 504 57017
rect 576 56941 626 57017
rect 698 56941 752 57017
rect 824 56941 946 57017
rect 463 56891 946 56941
rect 464 55068 947 55109
rect 463 55060 947 55068
rect 463 54984 504 55060
rect 576 54984 626 55060
rect 698 54984 752 55060
rect 824 54984 947 55060
rect 463 54913 947 54984
rect 463 54837 504 54913
rect 576 54837 626 54913
rect 698 54837 752 54913
rect 824 54837 947 54913
rect 463 54776 947 54837
rect 463 54700 504 54776
rect 576 54700 626 54776
rect 698 54700 752 54776
rect 824 54700 947 54776
rect 463 54650 947 54700
rect 463 53301 946 53350
rect 463 53225 504 53301
rect 576 53225 626 53301
rect 698 53225 752 53301
rect 824 53225 946 53301
rect 463 53154 946 53225
rect 463 53078 504 53154
rect 576 53078 626 53154
rect 698 53078 752 53154
rect 824 53078 946 53154
rect 463 53017 946 53078
rect 463 52941 504 53017
rect 576 52941 626 53017
rect 698 52941 752 53017
rect 824 52941 946 53017
rect 463 52891 946 52941
rect 464 51068 947 51109
rect 463 51060 947 51068
rect 463 50984 504 51060
rect 576 50984 626 51060
rect 698 50984 752 51060
rect 824 50984 947 51060
rect 463 50913 947 50984
rect 463 50837 504 50913
rect 576 50837 626 50913
rect 698 50837 752 50913
rect 824 50837 947 50913
rect 463 50776 947 50837
rect 463 50700 504 50776
rect 576 50700 626 50776
rect 698 50700 752 50776
rect 824 50700 947 50776
rect 463 50650 947 50700
rect 463 49299 946 49348
rect 463 49223 504 49299
rect 576 49223 626 49299
rect 698 49223 752 49299
rect 824 49223 946 49299
rect 463 49152 946 49223
rect 463 49076 504 49152
rect 576 49076 626 49152
rect 698 49076 752 49152
rect 824 49076 946 49152
rect 463 49015 946 49076
rect 463 48939 504 49015
rect 576 48939 626 49015
rect 698 48939 752 49015
rect 824 48939 946 49015
rect 463 48889 946 48939
rect 463 47060 946 47109
rect 463 46984 504 47060
rect 576 46984 626 47060
rect 698 46984 752 47060
rect 824 46984 946 47060
rect 463 46913 946 46984
rect 463 46837 504 46913
rect 576 46837 626 46913
rect 698 46837 752 46913
rect 824 46837 946 46913
rect 463 46776 946 46837
rect 463 46700 504 46776
rect 576 46700 626 46776
rect 698 46700 752 46776
rect 824 46700 946 46776
rect 463 46650 946 46700
rect 463 45301 946 45350
rect 463 45225 504 45301
rect 576 45225 626 45301
rect 698 45225 752 45301
rect 824 45225 946 45301
rect 463 45154 946 45225
rect 463 45078 504 45154
rect 576 45078 626 45154
rect 698 45078 752 45154
rect 824 45078 946 45154
rect 463 45017 946 45078
rect 463 44941 504 45017
rect 576 44941 626 45017
rect 698 44941 752 45017
rect 824 44941 946 45017
rect 463 44891 946 44941
rect 463 43060 946 43109
rect 463 42984 504 43060
rect 576 42984 626 43060
rect 698 42984 752 43060
rect 824 42984 946 43060
rect 463 42913 946 42984
rect 463 42837 504 42913
rect 576 42837 626 42913
rect 698 42837 752 42913
rect 824 42837 946 42913
rect 463 42776 946 42837
rect 463 42700 504 42776
rect 576 42700 626 42776
rect 698 42700 752 42776
rect 824 42700 946 42776
rect 463 42650 946 42700
rect 463 41301 946 41350
rect 463 41225 504 41301
rect 576 41225 626 41301
rect 698 41225 752 41301
rect 824 41225 946 41301
rect 463 41154 946 41225
rect 463 41078 504 41154
rect 576 41078 626 41154
rect 698 41078 752 41154
rect 824 41078 946 41154
rect 463 41017 946 41078
rect 463 40941 504 41017
rect 576 40941 626 41017
rect 698 40941 752 41017
rect 824 40941 946 41017
rect 463 40891 946 40941
rect 463 39060 946 39109
rect 463 38984 504 39060
rect 576 38984 626 39060
rect 698 38984 752 39060
rect 824 38984 946 39060
rect 463 38913 946 38984
rect 463 38837 504 38913
rect 576 38837 626 38913
rect 698 38837 752 38913
rect 824 38837 946 38913
rect 463 38776 946 38837
rect 463 38700 504 38776
rect 576 38700 626 38776
rect 698 38700 752 38776
rect 824 38700 946 38776
rect 463 38650 946 38700
rect 463 37300 946 37350
rect 463 37224 504 37300
rect 576 37224 626 37300
rect 698 37224 752 37300
rect 824 37224 946 37300
rect 463 37153 946 37224
rect 463 37077 504 37153
rect 576 37077 626 37153
rect 698 37077 752 37153
rect 824 37077 946 37153
rect 463 37016 946 37077
rect 463 36940 504 37016
rect 576 36940 626 37016
rect 698 36940 752 37016
rect 824 36940 946 37016
rect 463 36891 946 36940
rect 463 36890 836 36891
rect 944 35679 5768 35727
rect 944 35519 1306 35679
rect 1466 35519 1706 35679
rect 1866 35519 2106 35679
rect 2266 35519 2506 35679
rect 2666 35519 2906 35679
rect 3066 35519 3306 35679
rect 3466 35519 3706 35679
rect 3866 35519 4106 35679
rect 4266 35519 4506 35679
rect 4666 35519 4906 35679
rect 5066 35519 5306 35679
rect 5462 35519 5768 35679
rect 944 35496 5768 35519
rect 944 35336 1008 35496
rect 1168 35476 5547 35496
rect 1168 35336 1238 35476
rect 944 35138 1238 35336
rect 2468 35409 2935 35410
rect 2468 35395 3015 35409
rect 2012 35316 2160 35333
rect 2012 35315 2108 35316
rect 2012 35273 2020 35315
rect 2062 35274 2108 35315
rect 2150 35274 2160 35316
rect 2062 35273 2160 35274
rect 2012 35226 2160 35273
rect 2012 35225 2109 35226
rect 2012 35183 2021 35225
rect 2063 35184 2109 35225
rect 2151 35184 2160 35226
rect 2250 35321 2396 35329
rect 2250 35279 2262 35321
rect 2304 35279 2342 35321
rect 2384 35279 2396 35321
rect 2250 35241 2396 35279
rect 2468 35281 2485 35395
rect 2603 35281 2641 35395
rect 2759 35281 2797 35395
rect 2915 35281 3015 35395
rect 5478 35336 5547 35476
rect 5707 35336 5768 35496
rect 2468 35270 3015 35281
rect 2250 35199 2262 35241
rect 2304 35199 2342 35241
rect 2384 35223 2396 35241
rect 2384 35199 2527 35223
rect 2250 35189 2527 35199
rect 2063 35183 2160 35184
rect 2012 35169 2160 35183
rect 944 35137 1126 35138
rect 944 35062 969 35137
rect 1041 35096 1126 35137
rect 1198 35063 1238 35138
rect 944 35021 1008 35062
rect 1168 35024 1238 35063
rect 944 34946 972 35021
rect 1198 34949 1238 35024
rect 944 34936 1008 34946
rect 1168 34936 1238 34949
rect 944 34696 1238 34936
rect 1606 35085 1671 35086
rect 1606 34977 1736 35085
rect 2018 34977 2156 35169
rect 1606 34937 1640 34977
rect 1606 34850 1640 34896
rect 1864 34851 1898 34977
rect 2122 34937 2156 34977
rect 2122 34849 2156 34896
rect 2235 34977 2369 35085
rect 2493 35084 2527 35189
rect 2651 34977 3015 35270
rect 3139 35328 3285 35336
rect 3139 35286 3151 35328
rect 3193 35286 3231 35328
rect 3273 35286 3285 35328
rect 3139 35248 3285 35286
rect 3139 35206 3151 35248
rect 3193 35206 3231 35248
rect 3273 35206 3285 35248
rect 3139 35196 3285 35206
rect 3139 35085 3173 35196
rect 5478 35108 5768 35336
rect 5321 35096 5768 35108
rect 3297 34977 3431 35085
rect 5321 35074 5547 35096
rect 2235 34945 2269 34977
rect 2235 34851 2269 34890
rect 2493 34851 2527 34977
rect 2751 34945 2785 34977
rect 2751 34851 2785 34890
rect 2881 34949 2915 34977
rect 2881 34851 2915 34890
rect 3139 34851 3173 34977
rect 3397 34949 3431 34977
rect 3485 34981 3551 34982
rect 3485 34947 3501 34981
rect 3535 34947 3551 34981
rect 3485 34946 3551 34947
rect 5478 34936 5547 35074
rect 5707 34936 5768 35096
rect 3397 34851 3431 34890
rect 4915 34870 5157 34876
rect 3500 34836 3521 34870
rect 3555 34836 3573 34870
rect 4915 34836 4939 34870
rect 4973 34836 5157 34870
rect 4915 34828 5157 34836
rect 5191 34871 5263 34876
rect 5191 34836 5215 34871
rect 5250 34836 5263 34871
rect 5191 34829 5263 34836
rect 5191 34828 5238 34829
rect 944 34536 1008 34696
rect 1168 34536 1238 34696
rect 944 34296 1238 34536
rect 5478 34696 5768 34936
rect 5478 34536 5547 34696
rect 5707 34536 5768 34696
rect 944 34136 1008 34296
rect 1168 34136 1238 34296
rect 1939 34260 2123 34269
rect 1939 34225 2079 34260
rect 2115 34225 2123 34260
rect 1939 34217 2123 34225
rect 3418 34202 3542 34343
rect 4340 34202 4464 34343
rect 5478 34296 5768 34536
rect 5232 34258 5304 34262
rect 5232 34224 5262 34258
rect 5296 34224 5304 34258
rect 5232 34207 5304 34224
rect 944 33896 1238 34136
rect 5478 34136 5547 34296
rect 5707 34136 5768 34296
rect 5478 34020 5768 34136
rect 5412 33986 5768 34020
rect 944 33736 1008 33896
rect 1168 33736 1238 33896
rect 5478 33896 5768 33986
rect 24526 34392 25428 34442
rect 24526 34316 25069 34392
rect 25141 34316 25191 34392
rect 25263 34316 25317 34392
rect 25389 34316 25428 34392
rect 24526 34245 25428 34316
rect 24526 34169 25069 34245
rect 25141 34169 25191 34245
rect 25263 34169 25317 34245
rect 25389 34169 25428 34245
rect 24526 34108 25428 34169
rect 24526 34032 25069 34108
rect 25141 34032 25191 34108
rect 25263 34032 25317 34108
rect 25389 34032 25428 34108
rect 24526 33983 25428 34032
rect 24526 33982 25401 33983
rect 2173 33745 2369 33788
rect 944 33496 1238 33736
rect 3418 33663 3542 33804
rect 4340 33663 4464 33804
rect 5296 33748 5304 33780
rect 5275 33745 5304 33748
rect 5478 33736 5547 33896
rect 5707 33736 5768 33896
rect 944 33336 1008 33496
rect 1168 33336 1238 33496
rect 5478 33496 5768 33736
rect 944 33096 1238 33336
rect 2280 33358 2339 33375
rect 2563 33363 2597 33465
rect 2280 33310 2286 33358
rect 2332 33310 2339 33358
rect 2280 33245 2339 33310
rect 2280 33200 2286 33245
rect 2332 33200 2339 33245
rect 5478 33336 5547 33496
rect 5707 33336 5768 33496
rect 2280 33187 2339 33200
rect 944 33079 1008 33096
rect 1168 33079 1238 33096
rect 944 32991 975 33079
rect 1203 32991 1238 33079
rect 944 32949 1008 32991
rect 1168 32949 1238 32991
rect 944 32861 975 32949
rect 1070 32861 1109 32936
rect 1204 32861 1238 32949
rect 2305 33140 2339 33173
rect 2305 33029 2339 33092
rect 2563 33029 2597 33155
rect 2821 33140 2855 33173
rect 2821 33029 2855 33092
rect 2305 32921 2439 33029
rect 2721 32921 2855 33029
rect 2937 33140 2971 33173
rect 2937 33029 2971 33092
rect 3195 33029 3229 33155
rect 3453 33140 3487 33173
rect 3439 33092 3453 33138
rect 3544 33138 3562 33172
rect 3596 33138 3612 33172
rect 4915 33170 5157 33178
rect 4915 33136 5123 33170
rect 4915 33130 5157 33136
rect 5191 33170 5261 33178
rect 5191 33136 5215 33170
rect 5249 33136 5261 33170
rect 5191 33131 5261 33136
rect 5191 33130 5257 33131
rect 5478 33096 5768 33336
rect 3439 33029 3479 33092
rect 2937 32921 3071 33029
rect 944 32650 1238 32861
rect 3195 32838 3229 32921
rect 3353 32838 3479 33029
rect 3513 33038 3556 33058
rect 3513 33003 3516 33038
rect 3553 33003 3556 33038
rect 3513 32987 3556 33003
rect 5478 32936 5547 33096
rect 5707 32936 5768 33096
rect 5478 32932 5768 32936
rect 5321 32898 5768 32932
rect 3138 32830 3285 32838
rect 3138 32788 3151 32830
rect 3193 32788 3231 32830
rect 3273 32788 3285 32830
rect 3138 32750 3285 32788
rect 3138 32711 3151 32750
rect 3193 32711 3231 32750
rect 3273 32711 3285 32750
rect 3138 32703 3285 32711
rect 3352 32830 3499 32838
rect 3352 32788 3365 32830
rect 3407 32788 3445 32830
rect 3487 32788 3499 32830
rect 3352 32747 3499 32788
rect 3352 32713 3365 32747
rect 3407 32713 3445 32747
rect 3487 32713 3499 32747
rect 3352 32707 3499 32713
rect 5478 32650 5768 32898
rect 944 32614 5768 32650
rect 944 32454 1008 32614
rect 1168 32454 1408 32614
rect 1568 32454 1808 32614
rect 1968 32454 2208 32614
rect 2368 32454 2608 32614
rect 2768 32454 3008 32614
rect 3168 32454 3408 32614
rect 3568 32454 3808 32614
rect 3968 32454 4208 32614
rect 4368 32454 4608 32614
rect 4768 32454 5008 32614
rect 5168 32454 5547 32614
rect 5707 32454 5768 32614
rect 944 32449 5768 32454
rect 24526 32632 25428 32682
rect 24526 32556 25069 32632
rect 25141 32556 25191 32632
rect 25263 32556 25317 32632
rect 25389 32556 25428 32632
rect 24526 32485 25428 32556
rect 944 32411 5767 32449
rect 24526 32409 25069 32485
rect 25141 32409 25191 32485
rect 25263 32409 25317 32485
rect 25389 32409 25428 32485
rect 24526 32348 25428 32409
rect 24526 32272 25069 32348
rect 25141 32272 25191 32348
rect 25263 32272 25317 32348
rect 25389 32272 25428 32348
rect 24526 32223 25428 32272
rect 24526 32222 25401 32223
rect 485 27110 847 27111
rect 463 27061 1116 27110
rect 463 26985 504 27061
rect 576 26985 626 27061
rect 698 26985 752 27061
rect 824 26985 1116 27061
rect 463 26914 1116 26985
rect 463 26838 504 26914
rect 576 26838 626 26914
rect 698 26838 752 26914
rect 824 26838 1116 26914
rect 463 26777 1116 26838
rect 463 26701 504 26777
rect 576 26701 626 26777
rect 698 26701 752 26777
rect 824 26701 1116 26777
rect 463 26652 1116 26701
rect 463 26651 946 26652
rect 463 25294 1026 25350
rect 463 25218 504 25294
rect 576 25218 626 25294
rect 698 25218 752 25294
rect 824 25218 1026 25294
rect 463 25147 1026 25218
rect 463 25071 504 25147
rect 576 25071 626 25147
rect 698 25071 752 25147
rect 824 25071 1026 25147
rect 463 25010 1026 25071
rect 463 24934 504 25010
rect 576 24934 626 25010
rect 698 24934 752 25010
rect 824 24934 1026 25010
rect 463 24890 1026 24934
rect 463 24885 863 24890
rect 463 24884 862 24885
rect 463 23060 946 23109
rect 463 22984 504 23060
rect 576 22984 626 23060
rect 698 22984 752 23060
rect 824 22984 946 23060
rect 463 22913 946 22984
rect 463 22837 504 22913
rect 576 22837 626 22913
rect 698 22837 752 22913
rect 824 22837 946 22913
rect 463 22776 946 22837
rect 463 22700 504 22776
rect 576 22700 626 22776
rect 698 22700 752 22776
rect 824 22700 946 22776
rect 463 22650 946 22700
rect 463 21300 946 21349
rect 463 21224 504 21300
rect 576 21224 626 21300
rect 698 21224 752 21300
rect 824 21224 946 21300
rect 463 21153 946 21224
rect 463 21077 504 21153
rect 576 21077 626 21153
rect 698 21077 752 21153
rect 824 21077 946 21153
rect 463 21016 946 21077
rect 463 20940 504 21016
rect 576 20940 626 21016
rect 698 20940 752 21016
rect 824 20940 946 21016
rect 463 20890 946 20940
rect 463 19060 946 19109
rect 463 18984 504 19060
rect 576 18984 626 19060
rect 698 18984 752 19060
rect 824 18984 946 19060
rect 463 18913 946 18984
rect 463 18837 504 18913
rect 576 18837 626 18913
rect 698 18837 752 18913
rect 824 18837 946 18913
rect 463 18776 946 18837
rect 463 18700 504 18776
rect 576 18700 626 18776
rect 698 18700 752 18776
rect 824 18700 946 18776
rect 463 18650 946 18700
rect 463 17301 946 17350
rect 463 17225 504 17301
rect 576 17225 626 17301
rect 698 17225 752 17301
rect 824 17225 946 17301
rect 463 17154 946 17225
rect 463 17078 504 17154
rect 576 17078 626 17154
rect 698 17078 752 17154
rect 824 17078 946 17154
rect 463 17017 946 17078
rect 463 16941 504 17017
rect 576 16941 626 17017
rect 698 16941 752 17017
rect 824 16941 946 17017
rect 463 16891 946 16941
rect 463 15060 946 15109
rect 463 14984 504 15060
rect 576 14984 626 15060
rect 698 14984 752 15060
rect 824 14984 946 15060
rect 463 14913 946 14984
rect 463 14837 504 14913
rect 576 14837 626 14913
rect 698 14837 752 14913
rect 824 14837 946 14913
rect 463 14776 946 14837
rect 463 14700 504 14776
rect 576 14700 626 14776
rect 698 14700 752 14776
rect 824 14700 946 14776
rect 463 14650 946 14700
rect 463 13300 946 13349
rect 463 13224 504 13300
rect 576 13224 626 13300
rect 698 13224 752 13300
rect 824 13224 946 13300
rect 463 13153 946 13224
rect 463 13077 504 13153
rect 576 13077 626 13153
rect 698 13077 752 13153
rect 824 13077 946 13153
rect 463 13016 946 13077
rect 463 12940 504 13016
rect 576 12940 626 13016
rect 698 12940 752 13016
rect 824 12940 946 13016
rect 463 12890 946 12940
rect 463 11060 946 11109
rect 463 10984 504 11060
rect 576 10984 626 11060
rect 698 10984 752 11060
rect 824 10984 946 11060
rect 463 10913 946 10984
rect 463 10837 504 10913
rect 576 10837 626 10913
rect 698 10837 752 10913
rect 824 10837 946 10913
rect 463 10776 946 10837
rect 463 10700 504 10776
rect 576 10700 626 10776
rect 698 10700 752 10776
rect 824 10700 946 10776
rect 463 10650 946 10700
rect 463 9300 946 9349
rect 463 9224 504 9300
rect 576 9224 626 9300
rect 698 9224 752 9300
rect 824 9224 946 9300
rect 463 9153 946 9224
rect 463 9077 504 9153
rect 576 9077 626 9153
rect 698 9077 752 9153
rect 824 9077 946 9153
rect 463 9016 946 9077
rect 463 8940 504 9016
rect 576 8940 626 9016
rect 698 8940 752 9016
rect 824 8940 946 9016
rect 463 8890 946 8940
rect 463 7061 946 7110
rect 463 6985 504 7061
rect 576 6985 626 7061
rect 698 6985 752 7061
rect 824 6985 946 7061
rect 463 6914 946 6985
rect 463 6838 504 6914
rect 576 6838 626 6914
rect 698 6838 752 6914
rect 824 6838 946 6914
rect 463 6777 946 6838
rect 463 6701 504 6777
rect 576 6701 626 6777
rect 698 6701 752 6777
rect 824 6701 946 6777
rect 463 6651 946 6701
rect 463 5299 946 5348
rect 463 5223 504 5299
rect 576 5223 626 5299
rect 698 5223 752 5299
rect 824 5223 946 5299
rect 463 5152 946 5223
rect 463 5076 504 5152
rect 576 5076 626 5152
rect 698 5076 752 5152
rect 824 5076 946 5152
rect 463 5015 946 5076
rect 463 4939 504 5015
rect 576 4939 626 5015
rect 698 4939 752 5015
rect 824 4939 946 5015
rect 463 4889 946 4939
rect 463 3061 946 3110
rect 463 2985 504 3061
rect 576 2985 626 3061
rect 698 2985 752 3061
rect 824 2985 946 3061
rect 463 2914 946 2985
rect 463 2838 504 2914
rect 576 2838 626 2914
rect 698 2838 752 2914
rect 824 2838 946 2914
rect 463 2777 946 2838
rect 463 2701 504 2777
rect 576 2701 626 2777
rect 698 2701 752 2777
rect 824 2701 946 2777
rect 463 2651 946 2701
rect 463 1300 946 1349
rect 463 1224 504 1300
rect 576 1224 626 1300
rect 698 1224 752 1300
rect 824 1224 946 1300
rect 463 1153 946 1224
rect 463 1077 504 1153
rect 576 1077 626 1153
rect 698 1077 752 1153
rect 824 1077 946 1153
rect 463 1016 946 1077
rect 463 940 504 1016
rect 576 940 626 1016
rect 698 940 752 1016
rect 824 940 946 1016
rect 463 890 946 940
<< viali >>
rect 503 63376 575 63452
rect 629 63376 701 63452
rect 749 63376 821 63452
rect 25068 63416 25140 63492
rect 25194 63416 25266 63492
rect 25314 63416 25386 63492
rect 503 63258 575 63334
rect 629 63258 701 63334
rect 749 63258 821 63334
rect 25068 63298 25140 63374
rect 25194 63298 25266 63374
rect 25314 63298 25386 63374
rect 504 62984 576 63060
rect 626 62984 698 63060
rect 752 62984 824 63060
rect 504 62837 576 62913
rect 626 62837 698 62913
rect 752 62837 824 62913
rect 504 62700 576 62776
rect 626 62700 698 62776
rect 752 62700 824 62776
rect 26010 61995 26082 62071
rect 26136 61995 26208 62071
rect 26256 61995 26328 62071
rect 26010 61877 26082 61953
rect 26136 61877 26208 61953
rect 26256 61877 26328 61953
rect 504 61224 576 61300
rect 626 61224 698 61300
rect 752 61224 824 61300
rect 504 61077 576 61153
rect 626 61077 698 61153
rect 752 61077 824 61153
rect 504 60940 576 61016
rect 626 60940 698 61016
rect 752 60940 824 61016
rect 503 60703 575 60779
rect 629 60703 701 60779
rect 749 60703 821 60779
rect 503 60585 575 60661
rect 629 60585 701 60661
rect 749 60585 821 60661
rect 25068 60619 25140 60695
rect 25194 60619 25266 60695
rect 25314 60619 25386 60695
rect 25068 60501 25140 60577
rect 25194 60501 25266 60577
rect 25314 60501 25386 60577
rect 503 59374 575 59450
rect 629 59374 701 59450
rect 749 59374 821 59450
rect 25068 59416 25140 59492
rect 25194 59416 25266 59492
rect 25314 59416 25386 59492
rect 503 59256 575 59332
rect 629 59256 701 59332
rect 749 59256 821 59332
rect 25068 59298 25140 59374
rect 25194 59298 25266 59374
rect 25314 59298 25386 59374
rect 504 58984 576 59060
rect 626 58984 698 59060
rect 752 58984 824 59060
rect 504 58837 576 58913
rect 626 58837 698 58913
rect 752 58837 824 58913
rect 504 58700 576 58776
rect 626 58700 698 58776
rect 752 58700 824 58776
rect 26010 57982 26082 58058
rect 26136 57982 26208 58058
rect 26256 57982 26328 58058
rect 26010 57864 26082 57940
rect 26136 57864 26208 57940
rect 26256 57864 26328 57940
rect 504 57225 576 57301
rect 626 57225 698 57301
rect 752 57225 824 57301
rect 504 57078 576 57154
rect 626 57078 698 57154
rect 752 57078 824 57154
rect 504 56941 576 57017
rect 626 56941 698 57017
rect 752 56941 824 57017
rect 503 56634 575 56710
rect 629 56634 701 56710
rect 749 56634 821 56710
rect 25068 56619 25140 56695
rect 25194 56619 25266 56695
rect 25314 56619 25386 56695
rect 503 56516 575 56592
rect 629 56516 701 56592
rect 749 56516 821 56592
rect 25068 56501 25140 56577
rect 25194 56501 25266 56577
rect 25314 56501 25386 56577
rect 503 55456 575 55532
rect 629 55456 701 55532
rect 749 55456 821 55532
rect 25068 55416 25140 55492
rect 25194 55416 25266 55492
rect 25314 55416 25386 55492
rect 503 55338 575 55414
rect 629 55338 701 55414
rect 749 55338 821 55414
rect 25068 55298 25140 55374
rect 25194 55298 25266 55374
rect 25314 55298 25386 55374
rect 504 54984 576 55060
rect 626 54984 698 55060
rect 752 54984 824 55060
rect 504 54837 576 54913
rect 626 54837 698 54913
rect 752 54837 824 54913
rect 504 54700 576 54776
rect 626 54700 698 54776
rect 752 54700 824 54776
rect 26010 53981 26082 54057
rect 26136 53981 26208 54057
rect 26256 53981 26328 54057
rect 26010 53863 26082 53939
rect 26136 53863 26208 53939
rect 26256 53863 26328 53939
rect 504 53225 576 53301
rect 626 53225 698 53301
rect 752 53225 824 53301
rect 504 53078 576 53154
rect 626 53078 698 53154
rect 752 53078 824 53154
rect 504 52941 576 53017
rect 626 52941 698 53017
rect 752 52941 824 53017
rect 503 52608 575 52684
rect 629 52608 701 52684
rect 749 52608 821 52684
rect 25068 52619 25140 52695
rect 25194 52619 25266 52695
rect 25314 52619 25386 52695
rect 503 52490 575 52566
rect 629 52490 701 52566
rect 749 52490 821 52566
rect 25068 52501 25140 52577
rect 25194 52501 25266 52577
rect 25314 52501 25386 52577
rect 503 51405 575 51481
rect 629 51405 701 51481
rect 749 51405 821 51481
rect 25068 51470 25140 51546
rect 25194 51470 25266 51546
rect 25314 51470 25386 51546
rect 503 51287 575 51363
rect 629 51287 701 51363
rect 749 51287 821 51363
rect 25068 51352 25140 51428
rect 25194 51352 25266 51428
rect 25314 51352 25386 51428
rect 504 50984 576 51060
rect 626 50984 698 51060
rect 752 50984 824 51060
rect 504 50837 576 50913
rect 626 50837 698 50913
rect 752 50837 824 50913
rect 504 50700 576 50776
rect 626 50700 698 50776
rect 752 50700 824 50776
rect 26010 50020 26082 50096
rect 26136 50020 26208 50096
rect 26256 50020 26328 50096
rect 26010 49902 26082 49978
rect 26136 49902 26208 49978
rect 26256 49902 26328 49978
rect 504 49223 576 49299
rect 626 49223 698 49299
rect 752 49223 824 49299
rect 504 49076 576 49152
rect 626 49076 698 49152
rect 752 49076 824 49152
rect 504 48939 576 49015
rect 626 48939 698 49015
rect 752 48939 824 49015
rect 503 48628 575 48704
rect 629 48628 701 48704
rect 749 48628 821 48704
rect 503 48510 575 48586
rect 629 48510 701 48586
rect 749 48510 821 48586
rect 25068 48554 25140 48630
rect 25194 48554 25266 48630
rect 25314 48554 25386 48630
rect 25068 48436 25140 48512
rect 25194 48436 25266 48512
rect 25314 48436 25386 48512
rect 503 47421 575 47497
rect 629 47421 701 47497
rect 749 47421 821 47497
rect 503 47303 575 47379
rect 629 47303 701 47379
rect 749 47303 821 47379
rect 25068 47371 25140 47447
rect 25194 47371 25266 47447
rect 25314 47371 25386 47447
rect 25068 47253 25140 47329
rect 25194 47253 25266 47329
rect 25314 47253 25386 47329
rect 504 46984 576 47060
rect 626 46984 698 47060
rect 752 46984 824 47060
rect 504 46837 576 46913
rect 626 46837 698 46913
rect 752 46837 824 46913
rect 504 46700 576 46776
rect 626 46700 698 46776
rect 752 46700 824 46776
rect 26010 46003 26082 46079
rect 26136 46003 26208 46079
rect 26256 46003 26328 46079
rect 26010 45885 26082 45961
rect 26136 45885 26208 45961
rect 26256 45885 26328 45961
rect 504 45225 576 45301
rect 626 45225 698 45301
rect 752 45225 824 45301
rect 504 45078 576 45154
rect 626 45078 698 45154
rect 752 45078 824 45154
rect 504 44941 576 45017
rect 626 44941 698 45017
rect 752 44941 824 45017
rect 503 44655 575 44731
rect 629 44655 701 44731
rect 749 44655 821 44731
rect 503 44537 575 44613
rect 629 44537 701 44613
rect 749 44537 821 44613
rect 25068 44499 25140 44575
rect 25194 44499 25266 44575
rect 25314 44499 25386 44575
rect 25068 44381 25140 44457
rect 25194 44381 25266 44457
rect 25314 44381 25386 44457
rect 503 43468 575 43544
rect 629 43468 701 43544
rect 749 43468 821 43544
rect 503 43350 575 43426
rect 629 43350 701 43426
rect 749 43350 821 43426
rect 25068 43364 25140 43440
rect 25194 43364 25266 43440
rect 25314 43364 25386 43440
rect 25068 43246 25140 43322
rect 25194 43246 25266 43322
rect 25314 43246 25386 43322
rect 504 42984 576 43060
rect 626 42984 698 43060
rect 752 42984 824 43060
rect 504 42837 576 42913
rect 626 42837 698 42913
rect 752 42837 824 42913
rect 504 42700 576 42776
rect 626 42700 698 42776
rect 752 42700 824 42776
rect 26010 42082 26082 42158
rect 26136 42082 26208 42158
rect 26256 42082 26328 42158
rect 26010 41964 26082 42040
rect 26136 41964 26208 42040
rect 26256 41964 26328 42040
rect 504 41225 576 41301
rect 626 41225 698 41301
rect 752 41225 824 41301
rect 504 41078 576 41154
rect 626 41078 698 41154
rect 752 41078 824 41154
rect 504 40941 576 41017
rect 626 40941 698 41017
rect 752 40941 824 41017
rect 503 40646 575 40722
rect 629 40646 701 40722
rect 749 40646 821 40722
rect 25068 40605 25140 40681
rect 25194 40605 25266 40681
rect 25314 40605 25386 40681
rect 503 40528 575 40604
rect 629 40528 701 40604
rect 749 40528 821 40604
rect 25068 40487 25140 40563
rect 25194 40487 25266 40563
rect 25314 40487 25386 40563
rect 503 39493 575 39569
rect 629 39493 701 39569
rect 749 39493 821 39569
rect 25068 39452 25140 39528
rect 25194 39452 25266 39528
rect 25314 39452 25386 39528
rect 503 39375 575 39451
rect 629 39375 701 39451
rect 749 39375 821 39451
rect 25068 39334 25140 39410
rect 25194 39334 25266 39410
rect 25314 39334 25386 39410
rect 504 38984 576 39060
rect 626 38984 698 39060
rect 752 38984 824 39060
rect 504 38837 576 38913
rect 626 38837 698 38913
rect 752 38837 824 38913
rect 504 38700 576 38776
rect 626 38700 698 38776
rect 752 38700 824 38776
rect 26010 37824 26082 37900
rect 26136 37824 26208 37900
rect 26256 37824 26328 37900
rect 26010 37706 26082 37782
rect 26136 37706 26208 37782
rect 26256 37706 26328 37782
rect 504 37224 576 37300
rect 626 37224 698 37300
rect 752 37224 824 37300
rect 504 37077 576 37153
rect 626 37077 698 37153
rect 752 37077 824 37153
rect 504 36940 576 37016
rect 626 36940 698 37016
rect 752 36940 824 37016
rect 503 36433 575 36509
rect 629 36433 701 36509
rect 749 36433 821 36509
rect 503 36315 575 36391
rect 629 36315 701 36391
rect 749 36315 821 36391
rect 25068 36336 25140 36412
rect 25194 36336 25266 36412
rect 25314 36336 25386 36412
rect 25068 36218 25140 36294
rect 25194 36218 25266 36294
rect 25314 36218 25386 36294
rect 2020 35273 2062 35315
rect 2108 35274 2150 35316
rect 2021 35183 2063 35225
rect 2109 35184 2151 35226
rect 2262 35279 2304 35321
rect 2342 35279 2384 35321
rect 2485 35281 2603 35395
rect 2641 35281 2759 35395
rect 2797 35281 2915 35395
rect 2262 35199 2304 35241
rect 2342 35199 2384 35241
rect 969 35096 1041 35137
rect 1126 35096 1198 35138
rect 969 35062 1008 35096
rect 1008 35062 1041 35096
rect 1126 35063 1168 35096
rect 1168 35063 1198 35096
rect 972 34946 1008 35021
rect 1008 34946 1044 35021
rect 1126 34949 1168 35024
rect 1168 34949 1198 35024
rect 1864 34993 1898 35069
rect 1606 34896 1640 34937
rect 2122 34896 2156 34937
rect 3151 35286 3193 35328
rect 3231 35286 3273 35328
rect 3151 35206 3193 35248
rect 3231 35206 3273 35248
rect 2235 34890 2269 34945
rect 2751 34890 2785 34945
rect 2881 34890 2915 34949
rect 3397 34890 3431 34949
rect 3501 34947 3535 34981
rect 4851 34926 4885 34960
rect 3521 34836 3555 34870
rect 3853 34836 3888 34870
rect 4153 34836 4187 34870
rect 4705 34836 4739 34870
rect 4939 34836 4973 34870
rect 5215 34836 5250 34871
rect 4400 34779 4435 34813
rect 2079 34225 2115 34260
rect 2315 34224 2349 34258
rect 2407 34227 2441 34261
rect 2499 34224 2533 34258
rect 2629 34218 2663 34252
rect 5262 34224 5296 34258
rect 25069 34316 25141 34392
rect 25191 34316 25263 34392
rect 25317 34316 25389 34392
rect 25069 34169 25141 34245
rect 25191 34169 25263 34245
rect 25317 34169 25389 34245
rect 25069 34032 25141 34108
rect 25191 34032 25263 34108
rect 25317 34032 25389 34108
rect 2081 33748 2115 33782
rect 2405 33753 2439 33787
rect 2489 33754 2523 33788
rect 2586 33748 2620 33782
rect 5262 33748 5296 33782
rect 2286 33310 2332 33358
rect 2286 33200 2332 33245
rect 4407 33193 4441 33227
rect 975 32991 1008 33079
rect 1008 32991 1070 33079
rect 1108 32991 1168 33079
rect 1168 32991 1203 33079
rect 975 32936 1008 32949
rect 1008 32936 1070 32949
rect 1109 32936 1168 32949
rect 1168 32936 1204 32949
rect 975 32861 1070 32936
rect 1109 32861 1204 32936
rect 2305 33092 2339 33140
rect 2821 33092 2855 33140
rect 2937 33092 2971 33140
rect 3453 33092 3487 33140
rect 3562 33138 3596 33172
rect 3837 33137 3871 33171
rect 4153 33136 4187 33170
rect 4705 33136 4739 33170
rect 5123 33136 5157 33170
rect 5215 33136 5249 33170
rect 4851 33046 4885 33080
rect 3516 33003 3553 33038
rect 3151 32788 3193 32830
rect 3231 32788 3273 32830
rect 3151 32711 3193 32750
rect 3231 32711 3273 32750
rect 3365 32788 3407 32830
rect 3445 32788 3487 32830
rect 3365 32713 3407 32747
rect 3445 32713 3487 32747
rect 25069 32556 25141 32632
rect 25191 32556 25263 32632
rect 25317 32556 25389 32632
rect 25069 32409 25141 32485
rect 25191 32409 25263 32485
rect 25317 32409 25389 32485
rect 25069 32272 25141 32348
rect 25191 32272 25263 32348
rect 25317 32272 25389 32348
rect 503 28226 575 28302
rect 629 28226 701 28302
rect 749 28226 821 28302
rect 25068 28226 25140 28302
rect 25194 28226 25266 28302
rect 25314 28226 25386 28302
rect 503 28108 575 28184
rect 629 28108 701 28184
rect 749 28108 821 28184
rect 25068 28108 25140 28184
rect 25194 28108 25266 28184
rect 25314 28108 25386 28184
rect 503 27444 575 27520
rect 629 27444 701 27520
rect 749 27444 821 27520
rect 25068 27444 25140 27520
rect 25194 27444 25266 27520
rect 25314 27444 25386 27520
rect 503 27326 575 27402
rect 629 27326 701 27402
rect 749 27326 821 27402
rect 25068 27326 25140 27402
rect 25194 27326 25266 27402
rect 25314 27326 25386 27402
rect 504 26985 576 27061
rect 626 26985 698 27061
rect 752 26985 824 27061
rect 504 26838 576 26914
rect 626 26838 698 26914
rect 752 26838 824 26914
rect 504 26701 576 26777
rect 626 26701 698 26777
rect 752 26701 824 26777
rect 26010 26054 26082 26130
rect 26136 26054 26208 26130
rect 26256 26054 26328 26130
rect 26010 25936 26082 26012
rect 26136 25936 26208 26012
rect 26256 25936 26328 26012
rect 504 25218 576 25294
rect 626 25218 698 25294
rect 752 25218 824 25294
rect 504 25071 576 25147
rect 626 25071 698 25147
rect 752 25071 824 25147
rect 504 24934 576 25010
rect 626 24934 698 25010
rect 752 24934 824 25010
rect 503 24532 575 24608
rect 629 24532 701 24608
rect 749 24532 821 24608
rect 503 24414 575 24490
rect 629 24414 701 24490
rect 749 24414 821 24490
rect 25068 24483 25140 24559
rect 25194 24483 25266 24559
rect 25314 24483 25386 24559
rect 25068 24365 25140 24441
rect 25194 24365 25266 24441
rect 25314 24365 25386 24441
rect 503 23528 575 23604
rect 629 23528 701 23604
rect 749 23528 821 23604
rect 503 23410 575 23486
rect 629 23410 701 23486
rect 749 23410 821 23486
rect 25068 23366 25140 23442
rect 25194 23366 25266 23442
rect 25314 23366 25386 23442
rect 25068 23248 25140 23324
rect 25194 23248 25266 23324
rect 25314 23248 25386 23324
rect 504 22984 576 23060
rect 626 22984 698 23060
rect 752 22984 824 23060
rect 504 22837 576 22913
rect 626 22837 698 22913
rect 752 22837 824 22913
rect 504 22700 576 22776
rect 626 22700 698 22776
rect 752 22700 824 22776
rect 26010 21895 26082 21971
rect 26136 21895 26208 21971
rect 26256 21895 26328 21971
rect 26010 21777 26082 21853
rect 26136 21777 26208 21853
rect 26256 21777 26328 21853
rect 504 21224 576 21300
rect 626 21224 698 21300
rect 752 21224 824 21300
rect 504 21077 576 21153
rect 626 21077 698 21153
rect 752 21077 824 21153
rect 504 20940 576 21016
rect 626 20940 698 21016
rect 752 20940 824 21016
rect 503 20550 575 20626
rect 629 20550 701 20626
rect 749 20550 821 20626
rect 25068 20523 25140 20599
rect 25194 20523 25266 20599
rect 25314 20523 25386 20599
rect 503 20432 575 20508
rect 629 20432 701 20508
rect 749 20432 821 20508
rect 25068 20405 25140 20481
rect 25194 20405 25266 20481
rect 25314 20405 25386 20481
rect 503 19468 575 19544
rect 629 19468 701 19544
rect 749 19468 821 19544
rect 503 19350 575 19426
rect 629 19350 701 19426
rect 749 19350 821 19426
rect 25068 19348 25140 19424
rect 25194 19348 25266 19424
rect 25314 19348 25386 19424
rect 25068 19230 25140 19306
rect 25194 19230 25266 19306
rect 25314 19230 25386 19306
rect 504 18984 576 19060
rect 626 18984 698 19060
rect 752 18984 824 19060
rect 504 18837 576 18913
rect 626 18837 698 18913
rect 752 18837 824 18913
rect 504 18700 576 18776
rect 626 18700 698 18776
rect 752 18700 824 18776
rect 26010 18105 26082 18181
rect 26136 18105 26208 18181
rect 26256 18105 26328 18181
rect 26010 17987 26082 18063
rect 26136 17987 26208 18063
rect 26256 17987 26328 18063
rect 504 17225 576 17301
rect 626 17225 698 17301
rect 752 17225 824 17301
rect 504 17078 576 17154
rect 626 17078 698 17154
rect 752 17078 824 17154
rect 504 16941 576 17017
rect 626 16941 698 17017
rect 752 16941 824 17017
rect 503 16593 575 16669
rect 629 16593 701 16669
rect 749 16593 821 16669
rect 503 16475 575 16551
rect 629 16475 701 16551
rect 749 16475 821 16551
rect 25068 16507 25140 16583
rect 25194 16507 25266 16583
rect 25314 16507 25386 16583
rect 25068 16389 25140 16465
rect 25194 16389 25266 16465
rect 25314 16389 25386 16465
rect 503 15492 575 15568
rect 629 15492 701 15568
rect 749 15492 821 15568
rect 503 15374 575 15450
rect 629 15374 701 15450
rect 749 15374 821 15450
rect 25068 15336 25140 15412
rect 25194 15336 25266 15412
rect 25314 15336 25386 15412
rect 25068 15218 25140 15294
rect 25194 15218 25266 15294
rect 25314 15218 25386 15294
rect 504 14984 576 15060
rect 626 14984 698 15060
rect 752 14984 824 15060
rect 504 14837 576 14913
rect 626 14837 698 14913
rect 752 14837 824 14913
rect 504 14700 576 14776
rect 626 14700 698 14776
rect 752 14700 824 14776
rect 26010 13998 26082 14074
rect 26136 13998 26208 14074
rect 26256 13998 26328 14074
rect 26010 13880 26082 13956
rect 26136 13880 26208 13956
rect 26256 13880 26328 13956
rect 504 13224 576 13300
rect 626 13224 698 13300
rect 752 13224 824 13300
rect 504 13077 576 13153
rect 626 13077 698 13153
rect 752 13077 824 13153
rect 504 12940 576 13016
rect 626 12940 698 13016
rect 752 12940 824 13016
rect 503 12626 575 12702
rect 629 12626 701 12702
rect 749 12626 821 12702
rect 503 12508 575 12584
rect 629 12508 701 12584
rect 749 12508 821 12584
rect 25068 12575 25140 12651
rect 25194 12575 25266 12651
rect 25314 12575 25386 12651
rect 25068 12457 25140 12533
rect 25194 12457 25266 12533
rect 25314 12457 25386 12533
rect 503 11410 575 11486
rect 629 11410 701 11486
rect 749 11410 821 11486
rect 503 11292 575 11368
rect 629 11292 701 11368
rect 749 11292 821 11368
rect 25068 11361 25140 11437
rect 25194 11361 25266 11437
rect 25314 11361 25386 11437
rect 25068 11243 25140 11319
rect 25194 11243 25266 11319
rect 25314 11243 25386 11319
rect 504 10984 576 11060
rect 626 10984 698 11060
rect 752 10984 824 11060
rect 504 10837 576 10913
rect 626 10837 698 10913
rect 752 10837 824 10913
rect 504 10700 576 10776
rect 626 10700 698 10776
rect 752 10700 824 10776
rect 26010 10180 26082 10256
rect 26136 10180 26208 10256
rect 26256 10180 26328 10256
rect 26010 10062 26082 10138
rect 26136 10062 26208 10138
rect 26256 10062 26328 10138
rect 504 9224 576 9300
rect 626 9224 698 9300
rect 752 9224 824 9300
rect 504 9077 576 9153
rect 626 9077 698 9153
rect 752 9077 824 9153
rect 504 8940 576 9016
rect 626 8940 698 9016
rect 752 8940 824 9016
rect 503 8545 575 8621
rect 629 8545 701 8621
rect 749 8545 821 8621
rect 25068 8518 25140 8594
rect 25194 8518 25266 8594
rect 25314 8518 25386 8594
rect 503 8427 575 8503
rect 629 8427 701 8503
rect 749 8427 821 8503
rect 25068 8400 25140 8476
rect 25194 8400 25266 8476
rect 25314 8400 25386 8476
rect 503 7423 575 7499
rect 629 7423 701 7499
rect 749 7423 821 7499
rect 503 7305 575 7381
rect 629 7305 701 7381
rect 749 7305 821 7381
rect 25068 7361 25140 7437
rect 25194 7361 25266 7437
rect 25314 7361 25386 7437
rect 25068 7243 25140 7319
rect 25194 7243 25266 7319
rect 25314 7243 25386 7319
rect 504 6985 576 7061
rect 626 6985 698 7061
rect 752 6985 824 7061
rect 504 6838 576 6914
rect 626 6838 698 6914
rect 752 6838 824 6914
rect 504 6701 576 6777
rect 626 6701 698 6777
rect 752 6701 824 6777
rect 26010 6216 26082 6292
rect 26136 6216 26208 6292
rect 26256 6216 26328 6292
rect 26010 6098 26082 6174
rect 26136 6098 26208 6174
rect 26256 6098 26328 6174
rect 504 5223 576 5299
rect 626 5223 698 5299
rect 752 5223 824 5299
rect 504 5076 576 5152
rect 626 5076 698 5152
rect 752 5076 824 5152
rect 504 4939 576 5015
rect 626 4939 698 5015
rect 752 4939 824 5015
rect 503 4563 575 4639
rect 629 4563 701 4639
rect 749 4563 821 4639
rect 503 4445 575 4521
rect 629 4445 701 4521
rect 749 4445 821 4521
rect 25068 4518 25140 4594
rect 25194 4518 25266 4594
rect 25314 4518 25386 4594
rect 25068 4400 25140 4476
rect 25194 4400 25266 4476
rect 25314 4400 25386 4476
rect 503 3452 575 3528
rect 629 3452 701 3528
rect 749 3452 821 3528
rect 503 3334 575 3410
rect 629 3334 701 3410
rect 749 3334 821 3410
rect 25068 3361 25140 3437
rect 25194 3361 25266 3437
rect 25314 3361 25386 3437
rect 25068 3243 25140 3319
rect 25194 3243 25266 3319
rect 25314 3243 25386 3319
rect 504 2985 576 3061
rect 626 2985 698 3061
rect 752 2985 824 3061
rect 504 2838 576 2914
rect 626 2838 698 2914
rect 752 2838 824 2914
rect 504 2701 576 2777
rect 626 2701 698 2777
rect 752 2701 824 2777
rect 26010 2204 26082 2280
rect 26136 2204 26208 2280
rect 26256 2204 26328 2280
rect 26010 2086 26082 2162
rect 26136 2086 26208 2162
rect 26256 2086 26328 2162
rect 504 1224 576 1300
rect 626 1224 698 1300
rect 752 1224 824 1300
rect 504 1077 576 1153
rect 626 1077 698 1153
rect 752 1077 824 1153
rect 504 940 576 1016
rect 626 940 698 1016
rect 752 940 824 1016
rect 503 629 575 705
rect 629 629 701 705
rect 749 629 821 705
rect 503 511 575 587
rect 629 511 701 587
rect 749 511 821 587
rect 25068 518 25140 594
rect 25194 518 25266 594
rect 25314 518 25386 594
rect 25068 400 25140 476
rect 25194 400 25266 476
rect 25314 400 25386 476
<< metal1 >>
rect 24946 63492 25426 63517
rect 463 63452 947 63477
rect 463 63376 503 63452
rect 575 63376 629 63452
rect 701 63376 749 63452
rect 821 63376 947 63452
rect 463 63334 947 63376
rect 463 63258 503 63334
rect 575 63258 629 63334
rect 701 63258 749 63334
rect 821 63258 947 63334
rect 24946 63416 25068 63492
rect 25140 63416 25194 63492
rect 25266 63416 25314 63492
rect 25386 63416 25426 63492
rect 24946 63374 25426 63416
rect 24946 63298 25068 63374
rect 25140 63298 25194 63374
rect 25266 63298 25314 63374
rect 25386 63298 25426 63374
rect 24946 63262 25426 63298
rect 463 63222 947 63258
rect 463 63060 863 63109
rect 463 62984 504 63060
rect 576 62984 626 63060
rect 698 62984 752 63060
rect 824 62984 863 63060
rect 463 62913 863 62984
rect 463 62837 504 62913
rect 576 62837 626 62913
rect 698 62837 752 62913
rect 824 62837 863 62913
rect 463 62776 863 62837
rect 463 62700 504 62776
rect 576 62700 626 62776
rect 698 62700 752 62776
rect 824 62700 863 62776
rect 463 62650 863 62700
rect 24946 62071 26370 62096
rect 24946 61995 26010 62071
rect 26082 61995 26136 62071
rect 26208 61995 26256 62071
rect 26328 61995 26370 62071
rect 24946 61953 26370 61995
rect 24946 61877 26010 61953
rect 26082 61877 26136 61953
rect 26208 61877 26256 61953
rect 26328 61877 26370 61953
rect 24946 61841 26370 61877
rect 463 61300 863 61349
rect 463 61224 504 61300
rect 576 61224 626 61300
rect 698 61224 752 61300
rect 824 61224 863 61300
rect 463 61153 863 61224
rect 463 61077 504 61153
rect 576 61077 626 61153
rect 698 61077 752 61153
rect 824 61077 863 61153
rect 463 61016 863 61077
rect 463 60940 504 61016
rect 576 60940 626 61016
rect 698 60940 752 61016
rect 824 60940 863 61016
rect 463 60890 863 60940
rect 463 60779 947 60804
rect 463 60703 503 60779
rect 575 60703 629 60779
rect 701 60703 749 60779
rect 821 60703 947 60779
rect 463 60661 947 60703
rect 463 60585 503 60661
rect 575 60585 629 60661
rect 701 60585 749 60661
rect 821 60585 947 60661
rect 463 60549 947 60585
rect 24946 60695 25428 60720
rect 24946 60619 25068 60695
rect 25140 60619 25194 60695
rect 25266 60619 25314 60695
rect 25386 60619 25428 60695
rect 24946 60577 25428 60619
rect 24946 60501 25068 60577
rect 25140 60501 25194 60577
rect 25266 60501 25314 60577
rect 25386 60501 25428 60577
rect 24946 60465 25428 60501
rect 24945 59517 24946 59530
rect 24945 59492 25426 59517
rect 463 59450 947 59475
rect 463 59374 503 59450
rect 575 59374 629 59450
rect 701 59374 749 59450
rect 821 59374 947 59450
rect 463 59332 947 59374
rect 463 59256 503 59332
rect 575 59256 629 59332
rect 701 59256 749 59332
rect 821 59256 947 59332
rect 24945 59416 25068 59492
rect 25140 59416 25194 59492
rect 25266 59416 25314 59492
rect 25386 59416 25426 59492
rect 24945 59374 25426 59416
rect 24945 59298 25068 59374
rect 25140 59298 25194 59374
rect 25266 59298 25314 59374
rect 25386 59298 25426 59374
rect 24945 59275 25426 59298
rect 24946 59262 25426 59275
rect 463 59220 947 59256
rect 463 59060 863 59109
rect 463 58984 504 59060
rect 576 58984 626 59060
rect 698 58984 752 59060
rect 824 58984 863 59060
rect 463 58913 863 58984
rect 463 58837 504 58913
rect 576 58837 626 58913
rect 698 58837 752 58913
rect 824 58837 863 58913
rect 463 58776 863 58837
rect 463 58700 504 58776
rect 576 58700 626 58776
rect 698 58700 752 58776
rect 824 58700 863 58776
rect 463 58650 863 58700
rect 24946 58058 26370 58083
rect 24946 57982 26010 58058
rect 26082 57982 26136 58058
rect 26208 57982 26256 58058
rect 26328 57982 26370 58058
rect 24946 57940 26370 57982
rect 24946 57864 26010 57940
rect 26082 57864 26136 57940
rect 26208 57864 26256 57940
rect 26328 57864 26370 57940
rect 24946 57828 26370 57864
rect 463 57301 863 57350
rect 463 57225 504 57301
rect 576 57225 626 57301
rect 698 57225 752 57301
rect 824 57225 863 57301
rect 463 57154 863 57225
rect 463 57078 504 57154
rect 576 57078 626 57154
rect 698 57078 752 57154
rect 824 57078 863 57154
rect 463 57017 863 57078
rect 463 56941 504 57017
rect 576 56941 626 57017
rect 698 56941 752 57017
rect 824 56941 863 57017
rect 463 56891 863 56941
rect 463 56710 947 56735
rect 463 56634 503 56710
rect 575 56634 629 56710
rect 701 56634 749 56710
rect 821 56634 947 56710
rect 463 56592 947 56634
rect 463 56516 503 56592
rect 575 56516 629 56592
rect 701 56516 749 56592
rect 821 56516 947 56592
rect 463 56480 947 56516
rect 24945 56720 24946 56760
rect 24945 56695 25428 56720
rect 24945 56619 25068 56695
rect 25140 56619 25194 56695
rect 25266 56619 25314 56695
rect 25386 56619 25428 56695
rect 24945 56577 25428 56619
rect 24945 56505 25068 56577
rect 24946 56501 25068 56505
rect 25140 56501 25194 56577
rect 25266 56501 25314 56577
rect 25386 56501 25428 56577
rect 24946 56465 25428 56501
rect 463 55532 947 55557
rect 463 55456 503 55532
rect 575 55456 629 55532
rect 701 55456 749 55532
rect 821 55456 947 55532
rect 463 55414 947 55456
rect 463 55338 503 55414
rect 575 55338 629 55414
rect 701 55338 749 55414
rect 821 55338 947 55414
rect 463 55302 947 55338
rect 24944 55492 25426 55517
rect 24944 55416 25068 55492
rect 25140 55416 25194 55492
rect 25266 55416 25314 55492
rect 25386 55416 25426 55492
rect 24944 55374 25426 55416
rect 24944 55298 25068 55374
rect 25140 55298 25194 55374
rect 25266 55298 25314 55374
rect 25386 55298 25426 55374
rect 24944 55262 25426 55298
rect 464 55068 864 55109
rect 463 55060 864 55068
rect 463 54984 504 55060
rect 576 54984 626 55060
rect 698 54984 752 55060
rect 824 54984 864 55060
rect 463 54913 864 54984
rect 463 54837 504 54913
rect 576 54837 626 54913
rect 698 54837 752 54913
rect 824 54837 864 54913
rect 463 54776 864 54837
rect 463 54700 504 54776
rect 576 54700 626 54776
rect 698 54700 752 54776
rect 824 54700 864 54776
rect 463 54650 864 54700
rect 24946 54057 26370 54082
rect 24946 53981 26010 54057
rect 26082 53981 26136 54057
rect 26208 53981 26256 54057
rect 26328 53981 26370 54057
rect 24946 53939 26370 53981
rect 24946 53863 26010 53939
rect 26082 53863 26136 53939
rect 26208 53863 26256 53939
rect 26328 53863 26370 53939
rect 24946 53827 26370 53863
rect 463 53301 863 53350
rect 463 53225 504 53301
rect 576 53225 626 53301
rect 698 53225 752 53301
rect 824 53225 863 53301
rect 463 53154 863 53225
rect 463 53078 504 53154
rect 576 53078 626 53154
rect 698 53078 752 53154
rect 824 53078 863 53154
rect 463 53017 863 53078
rect 463 52941 504 53017
rect 576 52941 626 53017
rect 698 52941 752 53017
rect 824 52941 863 53017
rect 463 52891 863 52941
rect 463 52684 949 52709
rect 463 52608 503 52684
rect 575 52608 629 52684
rect 701 52608 749 52684
rect 821 52608 949 52684
rect 463 52566 949 52608
rect 463 52490 503 52566
rect 575 52490 629 52566
rect 701 52490 749 52566
rect 821 52490 949 52566
rect 463 52454 949 52490
rect 24946 52695 25428 52720
rect 24946 52619 25068 52695
rect 25140 52619 25194 52695
rect 25266 52619 25314 52695
rect 25386 52619 25428 52695
rect 24946 52577 25428 52619
rect 24946 52501 25068 52577
rect 25140 52501 25194 52577
rect 25266 52501 25314 52577
rect 25386 52501 25428 52577
rect 24946 52465 25428 52501
rect 24945 51546 25427 51571
rect 463 51481 947 51506
rect 463 51405 503 51481
rect 575 51405 629 51481
rect 701 51405 749 51481
rect 821 51405 947 51481
rect 463 51363 947 51405
rect 463 51287 503 51363
rect 575 51287 629 51363
rect 701 51287 749 51363
rect 821 51287 947 51363
rect 24945 51470 25068 51546
rect 25140 51470 25194 51546
rect 25266 51470 25314 51546
rect 25386 51470 25427 51546
rect 24945 51428 25427 51470
rect 24945 51352 25068 51428
rect 25140 51352 25194 51428
rect 25266 51352 25314 51428
rect 25386 51352 25427 51428
rect 24945 51316 25427 51352
rect 463 51251 947 51287
rect 464 51068 864 51109
rect 463 51060 864 51068
rect 463 50984 504 51060
rect 576 50984 626 51060
rect 698 50984 752 51060
rect 824 50984 864 51060
rect 463 50913 864 50984
rect 463 50837 504 50913
rect 576 50837 626 50913
rect 698 50837 752 50913
rect 824 50837 864 50913
rect 463 50776 864 50837
rect 463 50700 504 50776
rect 576 50700 626 50776
rect 698 50700 752 50776
rect 824 50700 864 50776
rect 463 50650 864 50700
rect 24946 50096 26370 50121
rect 24946 50020 26010 50096
rect 26082 50020 26136 50096
rect 26208 50020 26256 50096
rect 26328 50020 26370 50096
rect 24946 49978 26370 50020
rect 24946 49902 26010 49978
rect 26082 49902 26136 49978
rect 26208 49902 26256 49978
rect 26328 49902 26370 49978
rect 24946 49866 26370 49902
rect 463 49299 863 49348
rect 463 49223 504 49299
rect 576 49223 626 49299
rect 698 49223 752 49299
rect 824 49223 863 49299
rect 463 49152 863 49223
rect 463 49076 504 49152
rect 576 49076 626 49152
rect 698 49076 752 49152
rect 824 49076 863 49152
rect 463 49015 863 49076
rect 463 48939 504 49015
rect 576 48939 626 49015
rect 698 48939 752 49015
rect 824 48939 863 49015
rect 463 48889 863 48939
rect 463 48704 947 48729
rect 463 48628 503 48704
rect 575 48628 629 48704
rect 701 48628 749 48704
rect 821 48628 947 48704
rect 463 48586 947 48628
rect 463 48510 503 48586
rect 575 48510 629 48586
rect 701 48510 749 48586
rect 821 48510 947 48586
rect 463 48474 947 48510
rect 24946 48630 25428 48655
rect 24946 48554 25068 48630
rect 25140 48554 25194 48630
rect 25266 48554 25314 48630
rect 25386 48554 25428 48630
rect 24946 48512 25428 48554
rect 24946 48436 25068 48512
rect 25140 48436 25194 48512
rect 25266 48436 25314 48512
rect 25386 48436 25428 48512
rect 24946 48400 25428 48436
rect 463 47497 949 47522
rect 463 47421 503 47497
rect 575 47421 629 47497
rect 701 47421 749 47497
rect 821 47421 949 47497
rect 463 47379 949 47421
rect 463 47303 503 47379
rect 575 47303 629 47379
rect 701 47303 749 47379
rect 821 47303 949 47379
rect 463 47267 949 47303
rect 24945 47447 25427 47472
rect 24945 47371 25068 47447
rect 25140 47371 25194 47447
rect 25266 47371 25314 47447
rect 25386 47371 25427 47447
rect 24945 47329 25427 47371
rect 24945 47253 25068 47329
rect 25140 47253 25194 47329
rect 25266 47253 25314 47329
rect 25386 47253 25427 47329
rect 24945 47217 25427 47253
rect 463 47060 863 47109
rect 463 46984 504 47060
rect 576 46984 626 47060
rect 698 46984 752 47060
rect 824 46984 863 47060
rect 463 46913 863 46984
rect 463 46837 504 46913
rect 576 46837 626 46913
rect 698 46837 752 46913
rect 824 46837 863 46913
rect 463 46776 863 46837
rect 463 46700 504 46776
rect 576 46700 626 46776
rect 698 46700 752 46776
rect 824 46700 863 46776
rect 463 46650 863 46700
rect 24946 46079 26370 46104
rect 24946 46003 26010 46079
rect 26082 46003 26136 46079
rect 26208 46003 26256 46079
rect 26328 46003 26370 46079
rect 24946 45961 26370 46003
rect 24946 45885 26010 45961
rect 26082 45885 26136 45961
rect 26208 45885 26256 45961
rect 26328 45885 26370 45961
rect 24946 45849 26370 45885
rect 463 45301 863 45350
rect 463 45225 504 45301
rect 576 45225 626 45301
rect 698 45225 752 45301
rect 824 45225 863 45301
rect 463 45154 863 45225
rect 463 45078 504 45154
rect 576 45078 626 45154
rect 698 45078 752 45154
rect 824 45078 863 45154
rect 463 45017 863 45078
rect 463 44941 504 45017
rect 576 44941 626 45017
rect 698 44941 752 45017
rect 824 44941 863 45017
rect 463 44891 863 44941
rect 463 44731 947 44756
rect 463 44655 503 44731
rect 575 44655 629 44731
rect 701 44655 749 44731
rect 821 44655 947 44731
rect 463 44613 947 44655
rect 463 44537 503 44613
rect 575 44537 629 44613
rect 701 44537 749 44613
rect 821 44537 947 44613
rect 463 44501 947 44537
rect 24946 44575 25428 44600
rect 24946 44499 25068 44575
rect 25140 44499 25194 44575
rect 25266 44499 25314 44575
rect 25386 44499 25428 44575
rect 24946 44457 25428 44499
rect 24946 44381 25068 44457
rect 25140 44381 25194 44457
rect 25266 44381 25314 44457
rect 25386 44381 25428 44457
rect 24946 44345 25428 44381
rect 463 43544 947 43569
rect 463 43468 503 43544
rect 575 43468 629 43544
rect 701 43468 749 43544
rect 821 43468 947 43544
rect 463 43426 947 43468
rect 463 43350 503 43426
rect 575 43350 629 43426
rect 701 43350 749 43426
rect 821 43350 947 43426
rect 463 43314 947 43350
rect 24946 43440 25428 43465
rect 24946 43364 25068 43440
rect 25140 43364 25194 43440
rect 25266 43364 25314 43440
rect 25386 43364 25428 43440
rect 24946 43322 25428 43364
rect 24946 43246 25068 43322
rect 25140 43246 25194 43322
rect 25266 43246 25314 43322
rect 25386 43246 25428 43322
rect 24946 43210 25428 43246
rect 463 43060 863 43109
rect 463 42984 504 43060
rect 576 42984 626 43060
rect 698 42984 752 43060
rect 824 42984 863 43060
rect 463 42913 863 42984
rect 463 42837 504 42913
rect 576 42837 626 42913
rect 698 42837 752 42913
rect 824 42837 863 42913
rect 463 42776 863 42837
rect 463 42700 504 42776
rect 576 42700 626 42776
rect 698 42700 752 42776
rect 824 42700 863 42776
rect 463 42650 863 42700
rect 24946 42158 26370 42183
rect 24946 42082 26010 42158
rect 26082 42082 26136 42158
rect 26208 42082 26256 42158
rect 26328 42082 26370 42158
rect 24946 42040 26370 42082
rect 24946 41964 26010 42040
rect 26082 41964 26136 42040
rect 26208 41964 26256 42040
rect 26328 41964 26370 42040
rect 24946 41928 26370 41964
rect 463 41301 863 41350
rect 463 41225 504 41301
rect 576 41225 626 41301
rect 698 41225 752 41301
rect 824 41225 863 41301
rect 463 41154 863 41225
rect 463 41078 504 41154
rect 576 41078 626 41154
rect 698 41078 752 41154
rect 824 41078 863 41154
rect 463 41017 863 41078
rect 463 40941 504 41017
rect 576 40941 626 41017
rect 698 40941 752 41017
rect 824 40941 863 41017
rect 463 40891 863 40941
rect 463 40722 947 40747
rect 463 40646 503 40722
rect 575 40646 629 40722
rect 701 40646 749 40722
rect 821 40646 947 40722
rect 463 40604 947 40646
rect 463 40528 503 40604
rect 575 40528 629 40604
rect 701 40528 749 40604
rect 821 40528 947 40604
rect 463 40492 947 40528
rect 24946 40681 25428 40706
rect 24946 40605 25068 40681
rect 25140 40605 25194 40681
rect 25266 40605 25314 40681
rect 25386 40605 25428 40681
rect 24946 40563 25428 40605
rect 24946 40487 25068 40563
rect 25140 40487 25194 40563
rect 25266 40487 25314 40563
rect 25386 40487 25428 40563
rect 24946 40451 25428 40487
rect 463 39569 947 39594
rect 463 39493 503 39569
rect 575 39493 629 39569
rect 701 39493 749 39569
rect 821 39493 947 39569
rect 463 39451 947 39493
rect 463 39375 503 39451
rect 575 39375 629 39451
rect 701 39375 749 39451
rect 821 39375 947 39451
rect 463 39339 947 39375
rect 24946 39528 25428 39553
rect 24946 39452 25068 39528
rect 25140 39452 25194 39528
rect 25266 39452 25314 39528
rect 25386 39452 25428 39528
rect 24946 39410 25428 39452
rect 24946 39334 25068 39410
rect 25140 39334 25194 39410
rect 25266 39334 25314 39410
rect 25386 39334 25428 39410
rect 24946 39298 25428 39334
rect 463 39060 863 39109
rect 463 38984 504 39060
rect 576 38984 626 39060
rect 698 38984 752 39060
rect 824 38984 863 39060
rect 463 38913 863 38984
rect 463 38837 504 38913
rect 576 38837 626 38913
rect 698 38837 752 38913
rect 824 38837 863 38913
rect 463 38776 863 38837
rect 463 38700 504 38776
rect 576 38700 626 38776
rect 698 38700 752 38776
rect 824 38700 863 38776
rect 463 38650 863 38700
rect 24946 37900 26370 37925
rect 24946 37824 26010 37900
rect 26082 37824 26136 37900
rect 26208 37824 26256 37900
rect 26328 37824 26370 37900
rect 24946 37782 26370 37824
rect 24946 37706 26010 37782
rect 26082 37706 26136 37782
rect 26208 37706 26256 37782
rect 26328 37706 26370 37782
rect 24946 37670 26370 37706
rect 463 37300 863 37350
rect 463 37224 504 37300
rect 576 37224 626 37300
rect 698 37224 752 37300
rect 824 37224 863 37300
rect 463 37153 863 37224
rect 463 37077 504 37153
rect 576 37077 626 37153
rect 698 37077 752 37153
rect 824 37077 863 37153
rect 463 37016 863 37077
rect 463 36940 504 37016
rect 576 36940 626 37016
rect 698 36940 752 37016
rect 824 36940 863 37016
rect 463 36891 863 36940
rect 463 36890 836 36891
rect 463 36509 946 36534
rect 463 36433 503 36509
rect 575 36433 629 36509
rect 701 36433 749 36509
rect 821 36433 946 36509
rect 463 36391 946 36433
rect 463 36315 503 36391
rect 575 36315 629 36391
rect 701 36315 749 36391
rect 821 36315 946 36391
rect 463 36279 946 36315
rect 24946 36412 25428 36437
rect 24946 36336 25068 36412
rect 25140 36336 25194 36412
rect 25266 36336 25314 36412
rect 25386 36336 25428 36412
rect 24946 36294 25428 36336
rect 24946 36218 25068 36294
rect 25140 36218 25194 36294
rect 25266 36218 25314 36294
rect 25386 36218 25428 36294
rect 24946 36182 25428 36218
rect 3287 35752 4421 35753
rect 0 35741 25902 35752
rect 0 35661 32 35741
rect 112 35661 157 35741
rect 237 35661 282 35741
rect 362 35726 25902 35741
rect 362 35661 25535 35726
rect 0 35646 25535 35661
rect 25615 35646 25660 35726
rect 25740 35646 25785 35726
rect 25865 35646 25902 35726
rect 0 35635 25902 35646
rect 0 35555 32 35635
rect 112 35555 157 35635
rect 237 35555 282 35635
rect 362 35606 25902 35635
rect 362 35555 25534 35606
rect 0 35526 25534 35555
rect 25614 35526 25659 35606
rect 25739 35526 25784 35606
rect 25864 35526 25902 35606
rect 0 35497 25902 35526
rect 2468 35395 2935 35410
rect 2011 35316 2160 35333
rect 2011 35315 2098 35316
rect 2011 35263 2020 35315
rect 2072 35264 2098 35315
rect 2150 35264 2160 35316
rect 2072 35263 2160 35264
rect 2011 35236 2160 35263
rect 2011 35235 2099 35236
rect 2011 35183 2021 35235
rect 2073 35184 2099 35235
rect 2151 35184 2160 35236
rect 2250 35321 2396 35329
rect 2250 35269 2262 35321
rect 2314 35269 2332 35321
rect 2384 35269 2396 35321
rect 2468 35281 2485 35395
rect 2603 35281 2641 35395
rect 2759 35281 2797 35395
rect 2915 35281 2935 35395
rect 2468 35270 2935 35281
rect 3139 35328 3285 35336
rect 3139 35276 3151 35328
rect 3203 35276 3221 35328
rect 3273 35276 3285 35328
rect 2250 35251 2396 35269
rect 2250 35199 2262 35251
rect 2314 35199 2332 35251
rect 2384 35199 2396 35251
rect 2250 35189 2396 35199
rect 3139 35258 3285 35276
rect 3139 35206 3151 35258
rect 3203 35206 3221 35258
rect 3273 35206 3285 35258
rect 3139 35196 3285 35206
rect 2073 35183 2160 35184
rect 944 35139 1238 35173
rect 2011 35169 2160 35183
rect 463 35138 3573 35139
rect 463 35137 1126 35138
rect 463 35130 969 35137
rect 463 35052 479 35130
rect 561 35052 593 35130
rect 675 35052 707 35130
rect 789 35062 969 35130
rect 1041 35063 1126 35137
rect 1198 35069 3573 35138
rect 1198 35063 1864 35069
rect 1041 35062 1864 35063
rect 789 35052 1864 35062
rect 463 35043 1864 35052
rect 944 35024 1238 35043
rect 944 35021 1126 35024
rect 944 34946 972 35021
rect 1044 34949 1126 35021
rect 1198 34949 1238 35024
rect 1856 34993 1864 35043
rect 1898 35043 3573 35069
rect 1898 34993 1907 35043
rect 1856 34979 1907 34993
rect 3489 34982 3550 34987
rect 3489 34981 3970 34982
rect 1044 34946 1238 34949
rect 944 34923 1238 34946
rect 2223 34945 2797 34954
rect 1594 34937 2168 34944
rect 1594 34896 1606 34937
rect 1640 34896 2122 34937
rect 2156 34896 2168 34937
rect 1594 34887 2168 34896
rect 2223 34890 2235 34945
rect 2269 34890 2751 34945
rect 2785 34890 2797 34945
rect 2223 34882 2797 34890
rect 2869 34949 3443 34955
rect 2869 34890 2881 34949
rect 2915 34890 3397 34949
rect 3431 34890 3443 34949
rect 3489 34947 3501 34981
rect 3535 34947 3970 34981
rect 24527 34972 25428 34998
rect 3489 34946 3970 34947
rect 3489 34941 3550 34946
rect 2869 34883 3443 34890
rect 3500 34870 3901 34876
rect 3500 34836 3521 34870
rect 3555 34836 3853 34870
rect 3888 34836 3901 34870
rect 3500 34829 3901 34836
rect 3942 34772 3970 34946
rect 4215 34960 4897 34966
rect 4215 34926 4851 34960
rect 4885 34926 4897 34960
rect 4215 34920 4897 34926
rect 4123 34828 4129 34880
rect 4181 34876 4187 34880
rect 4215 34876 4250 34920
rect 24527 34892 25061 34972
rect 25141 34892 25186 34972
rect 25266 34892 25311 34972
rect 25391 34892 25428 34972
rect 5210 34879 5262 34885
rect 4692 34876 4756 34878
rect 4181 34870 4250 34876
rect 4187 34836 4250 34870
rect 4181 34830 4250 34836
rect 4675 34870 4985 34876
rect 4675 34836 4705 34870
rect 4739 34836 4939 34870
rect 4973 34836 4985 34870
rect 4675 34830 4985 34836
rect 4181 34828 4187 34830
rect 4692 34826 4756 34830
rect 5208 34829 5210 34877
rect 4392 34813 4441 34825
rect 5210 34821 5262 34827
rect 24527 34852 25428 34892
rect 4392 34779 4400 34813
rect 4435 34779 4441 34813
rect 4392 34772 4441 34779
rect 3941 34737 4441 34772
rect 24527 34772 25060 34852
rect 25140 34772 25185 34852
rect 25265 34772 25310 34852
rect 25390 34772 25428 34852
rect 24527 34743 25428 34772
rect 0 34586 2193 34595
rect 0 34508 16 34586
rect 98 34508 130 34586
rect 212 34508 244 34586
rect 326 34508 2193 34586
rect 0 34499 2193 34508
rect 25028 34392 25428 34442
rect 4208 34348 4260 34354
rect 2493 34305 4208 34334
rect 2065 34217 2071 34269
rect 2123 34268 2129 34269
rect 2123 34258 2373 34268
rect 2123 34224 2315 34258
rect 2349 34224 2373 34258
rect 2123 34218 2373 34224
rect 2401 34261 2447 34275
rect 2401 34227 2407 34261
rect 2441 34227 2447 34261
rect 2123 34217 2129 34218
rect 2401 34210 2447 34227
rect 2493 34258 2541 34305
rect 4208 34290 4260 34296
rect 25028 34316 25069 34392
rect 25141 34316 25191 34392
rect 25263 34316 25317 34392
rect 25389 34316 25428 34392
rect 2493 34224 2499 34258
rect 2533 34224 2541 34258
rect 2493 34212 2541 34224
rect 2619 34252 2676 34275
rect 2619 34218 2629 34252
rect 2663 34218 2676 34252
rect 2405 34184 2447 34210
rect 2619 34202 2676 34218
rect 5252 34267 5304 34273
rect 5252 34209 5304 34215
rect 25028 34245 25428 34316
rect 2619 34184 2663 34202
rect 2405 34155 2663 34184
rect 25028 34169 25069 34245
rect 25141 34169 25191 34245
rect 25263 34169 25317 34245
rect 25389 34169 25428 34245
rect 25028 34108 25428 34169
rect 463 34042 2656 34051
rect 463 33964 479 34042
rect 561 33964 593 34042
rect 675 33964 707 34042
rect 789 33964 2656 34042
rect 25028 34032 25069 34108
rect 25141 34032 25191 34108
rect 25263 34032 25317 34108
rect 25389 34032 25428 34108
rect 25028 33983 25428 34032
rect 25028 33982 25401 33983
rect 463 33955 2656 33964
rect 4117 33889 4123 33897
rect 2474 33854 4123 33889
rect 2057 33738 2063 33790
rect 2115 33738 2139 33790
rect 2399 33787 2445 33851
rect 2399 33753 2405 33787
rect 2439 33753 2445 33787
rect 2399 33708 2445 33753
rect 2474 33788 2540 33854
rect 4117 33845 4123 33854
rect 4175 33845 4181 33897
rect 2474 33754 2489 33788
rect 2523 33754 2540 33788
rect 2474 33738 2540 33754
rect 2580 33782 2632 33795
rect 2580 33748 2586 33782
rect 2620 33748 2632 33782
rect 2580 33708 2632 33748
rect 5252 33791 5304 33797
rect 5252 33733 5304 33739
rect 2399 33680 2632 33708
rect 0 33498 1917 33507
rect 0 33420 16 33498
rect 98 33420 130 33498
rect 212 33420 244 33498
rect 326 33420 1917 33498
rect 0 33411 1917 33420
rect 24526 33476 25902 33502
rect 24526 33396 24560 33476
rect 24640 33396 24685 33476
rect 24765 33396 24810 33476
rect 24890 33396 25535 33476
rect 25615 33396 25660 33476
rect 25740 33396 25785 33476
rect 25865 33396 25902 33476
rect 2280 33358 2339 33375
rect 2280 33306 2283 33358
rect 2335 33306 2339 33358
rect 2280 33252 2339 33306
rect 24526 33356 25902 33396
rect 2280 33200 2283 33252
rect 2335 33200 2339 33252
rect 2280 33187 2339 33200
rect 3932 33265 4441 33300
rect 3527 33172 3895 33178
rect 2293 33140 2867 33150
rect 944 33079 1238 33111
rect 2293 33092 2305 33140
rect 2339 33092 2821 33140
rect 2855 33092 2867 33140
rect 2293 33083 2867 33092
rect 2925 33140 3499 33152
rect 2925 33092 2937 33140
rect 2971 33092 3453 33140
rect 3487 33092 3499 33140
rect 3527 33138 3562 33172
rect 3596 33171 3895 33172
rect 3596 33138 3837 33171
rect 3527 33137 3837 33138
rect 3871 33137 3895 33171
rect 3527 33131 3895 33137
rect 2925 33085 3499 33092
rect 944 32991 975 33079
rect 1070 32991 1108 33079
rect 1203 32991 1238 33079
rect 3932 33069 3975 33265
rect 4406 33233 4441 33265
rect 24526 33276 24559 33356
rect 24639 33276 24684 33356
rect 24764 33276 24809 33356
rect 24889 33276 25534 33356
rect 25614 33276 25659 33356
rect 25739 33276 25784 33356
rect 25864 33276 25902 33356
rect 24526 33247 25902 33276
rect 4401 33227 4448 33233
rect 4401 33193 4407 33227
rect 4441 33193 4448 33227
rect 4147 33176 4153 33182
rect 4123 33130 4153 33176
rect 4205 33130 4246 33182
rect 4401 33181 4448 33193
rect 5209 33181 5261 33187
rect 3569 33058 3975 33069
rect 3510 33038 3975 33058
rect 4210 33086 4246 33130
rect 4675 33178 4756 33180
rect 4675 33170 5169 33178
rect 4675 33136 4705 33170
rect 4739 33136 5123 33170
rect 5157 33136 5169 33170
rect 4675 33130 5169 33136
rect 4675 33128 4756 33130
rect 5209 33123 5261 33129
rect 4210 33080 4897 33086
rect 4210 33046 4851 33080
rect 4885 33046 4897 33080
rect 4210 33038 4897 33046
rect 3510 33003 3516 33038
rect 3553 33034 3975 33038
rect 3553 33023 3587 33034
rect 3553 33003 3559 33023
rect 3510 32991 3559 33003
rect 944 32963 1238 32991
rect 463 32954 3573 32963
rect 463 32876 479 32954
rect 561 32876 593 32954
rect 675 32876 707 32954
rect 789 32949 3573 32954
rect 789 32876 975 32949
rect 463 32867 975 32876
rect 944 32861 975 32867
rect 1070 32861 1109 32949
rect 1204 32867 3573 32949
rect 1204 32861 1238 32867
rect 944 32835 1238 32861
rect 3138 32830 3285 32838
rect 3138 32778 3151 32830
rect 3203 32778 3221 32830
rect 3273 32778 3285 32830
rect 3138 32763 3285 32778
rect 3138 32711 3151 32763
rect 3203 32711 3221 32763
rect 3273 32711 3285 32763
rect 3138 32649 3285 32711
rect 3352 32830 3499 32838
rect 3352 32778 3365 32830
rect 3417 32778 3435 32830
rect 3487 32778 3499 32830
rect 3352 32765 3499 32778
rect 3352 32713 3365 32765
rect 3417 32713 3435 32765
rect 3487 32713 3499 32765
rect 3352 32707 3499 32713
rect 25028 32632 25428 32682
rect 25028 32556 25069 32632
rect 25141 32556 25191 32632
rect 25263 32556 25317 32632
rect 25389 32556 25428 32632
rect 25028 32485 25428 32556
rect 25028 32409 25069 32485
rect 25141 32409 25191 32485
rect 25263 32409 25317 32485
rect 25389 32409 25428 32485
rect 25028 32348 25428 32409
rect 25028 32272 25069 32348
rect 25141 32272 25191 32348
rect 25263 32272 25317 32348
rect 25389 32272 25428 32348
rect 25028 32223 25428 32272
rect 25028 32222 25401 32223
rect 24514 31917 25427 31943
rect 24514 31837 25060 31917
rect 25140 31837 25185 31917
rect 25265 31837 25310 31917
rect 25390 31837 25427 31917
rect 24514 31797 25427 31837
rect 24514 31717 25059 31797
rect 25139 31717 25184 31797
rect 25264 31717 25309 31797
rect 25389 31717 25427 31797
rect 24514 31688 25427 31717
rect 463 28302 25428 28360
rect 463 28226 503 28302
rect 575 28226 629 28302
rect 701 28226 749 28302
rect 821 28226 25068 28302
rect 25140 28226 25194 28302
rect 25266 28226 25314 28302
rect 25386 28226 25428 28302
rect 463 28184 25428 28226
rect 463 28108 503 28184
rect 575 28108 629 28184
rect 701 28108 749 28184
rect 821 28108 25068 28184
rect 25140 28108 25194 28184
rect 25266 28108 25314 28184
rect 25386 28108 25428 28184
rect 463 28072 25428 28108
rect 463 27520 946 27545
rect 463 27444 503 27520
rect 575 27444 629 27520
rect 701 27444 749 27520
rect 821 27444 946 27520
rect 463 27402 946 27444
rect 463 27326 503 27402
rect 575 27326 629 27402
rect 701 27326 749 27402
rect 821 27326 946 27402
rect 463 27290 946 27326
rect 24946 27520 25428 27545
rect 24946 27444 25068 27520
rect 25140 27444 25194 27520
rect 25266 27444 25314 27520
rect 25386 27444 25428 27520
rect 24946 27402 25428 27444
rect 24946 27326 25068 27402
rect 25140 27326 25194 27402
rect 25266 27326 25314 27402
rect 25386 27326 25428 27402
rect 24946 27290 25428 27326
rect 463 27061 863 27111
rect 463 26985 504 27061
rect 576 26985 626 27061
rect 698 26985 752 27061
rect 824 26985 863 27061
rect 463 26914 863 26985
rect 463 26838 504 26914
rect 576 26838 626 26914
rect 698 26838 752 26914
rect 824 26838 863 26914
rect 463 26777 863 26838
rect 463 26701 504 26777
rect 576 26701 626 26777
rect 698 26701 752 26777
rect 824 26701 863 26777
rect 463 26651 863 26701
rect 24946 26130 26370 26155
rect 24946 26054 26010 26130
rect 26082 26054 26136 26130
rect 26208 26054 26256 26130
rect 26328 26054 26370 26130
rect 24946 26012 26370 26054
rect 24946 25936 26010 26012
rect 26082 25936 26136 26012
rect 26208 25936 26256 26012
rect 26328 25936 26370 26012
rect 24946 25900 26370 25936
rect 463 25294 863 25350
rect 463 25218 504 25294
rect 576 25218 626 25294
rect 698 25218 752 25294
rect 824 25218 863 25294
rect 463 25147 863 25218
rect 463 25071 504 25147
rect 576 25071 626 25147
rect 698 25071 752 25147
rect 824 25071 863 25147
rect 463 25010 863 25071
rect 463 24934 504 25010
rect 576 24934 626 25010
rect 698 24934 752 25010
rect 824 24934 863 25010
rect 463 24885 863 24934
rect 463 24884 862 24885
rect 944 24681 946 24880
rect 463 24608 946 24633
rect 463 24532 503 24608
rect 575 24532 629 24608
rect 701 24532 749 24608
rect 821 24532 946 24608
rect 463 24490 946 24532
rect 463 24414 503 24490
rect 575 24414 629 24490
rect 701 24414 749 24490
rect 821 24414 946 24490
rect 463 24378 946 24414
rect 24946 24559 25428 24584
rect 24946 24483 25068 24559
rect 25140 24483 25194 24559
rect 25266 24483 25314 24559
rect 25386 24483 25428 24559
rect 24946 24441 25428 24483
rect 24946 24365 25068 24441
rect 25140 24365 25194 24441
rect 25266 24365 25314 24441
rect 25386 24365 25428 24441
rect 24946 24329 25428 24365
rect 463 23604 946 23629
rect 463 23528 503 23604
rect 575 23528 629 23604
rect 701 23528 749 23604
rect 821 23528 946 23604
rect 463 23486 946 23528
rect 463 23410 503 23486
rect 575 23410 629 23486
rect 701 23410 749 23486
rect 821 23410 946 23486
rect 463 23374 946 23410
rect 24945 23442 25427 23467
rect 24945 23366 25068 23442
rect 25140 23366 25194 23442
rect 25266 23366 25314 23442
rect 25386 23366 25427 23442
rect 24945 23324 25427 23366
rect 24945 23248 25068 23324
rect 25140 23248 25194 23324
rect 25266 23248 25314 23324
rect 25386 23248 25427 23324
rect 24945 23212 25427 23248
rect 463 23060 863 23109
rect 463 22984 504 23060
rect 576 22984 626 23060
rect 698 22984 752 23060
rect 824 22984 863 23060
rect 463 22913 863 22984
rect 463 22837 504 22913
rect 576 22837 626 22913
rect 698 22837 752 22913
rect 824 22837 863 22913
rect 463 22776 863 22837
rect 463 22700 504 22776
rect 576 22700 626 22776
rect 698 22700 752 22776
rect 824 22700 863 22776
rect 463 22650 863 22700
rect 24946 21971 26370 21996
rect 24946 21895 26010 21971
rect 26082 21895 26136 21971
rect 26208 21895 26256 21971
rect 26328 21895 26370 21971
rect 24946 21853 26370 21895
rect 24946 21777 26010 21853
rect 26082 21777 26136 21853
rect 26208 21777 26256 21853
rect 26328 21777 26370 21853
rect 24946 21741 26370 21777
rect 463 21300 863 21349
rect 463 21224 504 21300
rect 576 21224 626 21300
rect 698 21224 752 21300
rect 824 21224 863 21300
rect 463 21153 863 21224
rect 463 21077 504 21153
rect 576 21077 626 21153
rect 698 21077 752 21153
rect 824 21077 863 21153
rect 463 21016 863 21077
rect 463 20940 504 21016
rect 576 20940 626 21016
rect 698 20940 752 21016
rect 824 20940 863 21016
rect 463 20890 863 20940
rect 463 20626 947 20651
rect 463 20550 503 20626
rect 575 20550 629 20626
rect 701 20550 749 20626
rect 821 20550 947 20626
rect 463 20508 947 20550
rect 463 20432 503 20508
rect 575 20432 629 20508
rect 701 20432 749 20508
rect 821 20432 947 20508
rect 463 20396 947 20432
rect 24946 20599 25428 20624
rect 24946 20523 25068 20599
rect 25140 20523 25194 20599
rect 25266 20523 25314 20599
rect 25386 20523 25428 20599
rect 24946 20481 25428 20523
rect 24946 20405 25068 20481
rect 25140 20405 25194 20481
rect 25266 20405 25314 20481
rect 25386 20405 25428 20481
rect 24946 20369 25428 20405
rect 463 19544 947 19569
rect 463 19468 503 19544
rect 575 19468 629 19544
rect 701 19468 749 19544
rect 821 19468 947 19544
rect 463 19426 947 19468
rect 463 19350 503 19426
rect 575 19350 629 19426
rect 701 19350 749 19426
rect 821 19350 947 19426
rect 463 19314 947 19350
rect 24946 19424 25428 19449
rect 24946 19348 25068 19424
rect 25140 19348 25194 19424
rect 25266 19348 25314 19424
rect 25386 19348 25428 19424
rect 24946 19306 25428 19348
rect 24946 19230 25068 19306
rect 25140 19230 25194 19306
rect 25266 19230 25314 19306
rect 25386 19230 25428 19306
rect 24946 19194 25428 19230
rect 463 19060 863 19109
rect 463 18984 504 19060
rect 576 18984 626 19060
rect 698 18984 752 19060
rect 824 18984 863 19060
rect 463 18913 863 18984
rect 463 18837 504 18913
rect 576 18837 626 18913
rect 698 18837 752 18913
rect 824 18837 863 18913
rect 463 18776 863 18837
rect 463 18700 504 18776
rect 576 18700 626 18776
rect 698 18700 752 18776
rect 824 18700 863 18776
rect 463 18650 863 18700
rect 24946 18181 26370 18206
rect 24946 18105 26010 18181
rect 26082 18105 26136 18181
rect 26208 18105 26256 18181
rect 26328 18105 26370 18181
rect 24946 18063 26370 18105
rect 24946 17987 26010 18063
rect 26082 17987 26136 18063
rect 26208 17987 26256 18063
rect 26328 17987 26370 18063
rect 24946 17951 26370 17987
rect 463 17301 863 17350
rect 463 17225 504 17301
rect 576 17225 626 17301
rect 698 17225 752 17301
rect 824 17225 863 17301
rect 463 17154 863 17225
rect 463 17078 504 17154
rect 576 17078 626 17154
rect 698 17078 752 17154
rect 824 17078 863 17154
rect 463 17017 863 17078
rect 463 16941 504 17017
rect 576 16941 626 17017
rect 698 16941 752 17017
rect 824 16941 863 17017
rect 463 16891 863 16941
rect 463 16669 947 16694
rect 463 16593 503 16669
rect 575 16593 629 16669
rect 701 16593 749 16669
rect 821 16593 947 16669
rect 463 16551 947 16593
rect 463 16475 503 16551
rect 575 16475 629 16551
rect 701 16475 749 16551
rect 821 16475 947 16551
rect 463 16439 947 16475
rect 24945 16583 25427 16608
rect 24945 16507 25068 16583
rect 25140 16507 25194 16583
rect 25266 16507 25314 16583
rect 25386 16507 25427 16583
rect 24945 16465 25427 16507
rect 24945 16389 25068 16465
rect 25140 16389 25194 16465
rect 25266 16389 25314 16465
rect 25386 16389 25427 16465
rect 24945 16353 25427 16389
rect 463 15568 947 15593
rect 463 15492 503 15568
rect 575 15492 629 15568
rect 701 15492 749 15568
rect 821 15492 947 15568
rect 463 15450 947 15492
rect 463 15374 503 15450
rect 575 15374 629 15450
rect 701 15374 749 15450
rect 821 15374 947 15450
rect 463 15338 947 15374
rect 24945 15412 25427 15437
rect 24945 15336 25068 15412
rect 25140 15336 25194 15412
rect 25266 15336 25314 15412
rect 25386 15336 25427 15412
rect 24945 15294 25427 15336
rect 24945 15218 25068 15294
rect 25140 15218 25194 15294
rect 25266 15218 25314 15294
rect 25386 15218 25427 15294
rect 24945 15182 25427 15218
rect 463 15060 863 15109
rect 463 14984 504 15060
rect 576 14984 626 15060
rect 698 14984 752 15060
rect 824 14984 863 15060
rect 463 14913 863 14984
rect 463 14837 504 14913
rect 576 14837 626 14913
rect 698 14837 752 14913
rect 824 14837 863 14913
rect 463 14776 863 14837
rect 463 14700 504 14776
rect 576 14700 626 14776
rect 698 14700 752 14776
rect 824 14700 863 14776
rect 463 14650 863 14700
rect 24946 14074 26370 14099
rect 24946 13998 26010 14074
rect 26082 13998 26136 14074
rect 26208 13998 26256 14074
rect 26328 13998 26370 14074
rect 24946 13956 26370 13998
rect 24946 13880 26010 13956
rect 26082 13880 26136 13956
rect 26208 13880 26256 13956
rect 26328 13880 26370 13956
rect 24946 13844 26370 13880
rect 463 13300 863 13349
rect 463 13224 504 13300
rect 576 13224 626 13300
rect 698 13224 752 13300
rect 824 13224 863 13300
rect 463 13153 863 13224
rect 463 13077 504 13153
rect 576 13077 626 13153
rect 698 13077 752 13153
rect 824 13077 863 13153
rect 463 13016 863 13077
rect 463 12940 504 13016
rect 576 12940 626 13016
rect 698 12940 752 13016
rect 824 12940 863 13016
rect 463 12890 863 12940
rect 463 12702 948 12727
rect 463 12626 503 12702
rect 575 12626 629 12702
rect 701 12626 749 12702
rect 821 12626 948 12702
rect 463 12584 948 12626
rect 463 12508 503 12584
rect 575 12508 629 12584
rect 701 12508 749 12584
rect 821 12508 948 12584
rect 463 12472 948 12508
rect 24945 12651 25427 12676
rect 24945 12575 25068 12651
rect 25140 12575 25194 12651
rect 25266 12575 25314 12651
rect 25386 12575 25427 12651
rect 24945 12533 25427 12575
rect 24945 12457 25068 12533
rect 25140 12457 25194 12533
rect 25266 12457 25314 12533
rect 25386 12457 25427 12533
rect 24945 12421 25427 12457
rect 463 11486 949 11511
rect 463 11410 503 11486
rect 575 11410 629 11486
rect 701 11410 749 11486
rect 821 11410 949 11486
rect 463 11368 949 11410
rect 463 11292 503 11368
rect 575 11292 629 11368
rect 701 11292 749 11368
rect 821 11292 949 11368
rect 463 11256 949 11292
rect 24945 11437 25427 11462
rect 24945 11361 25068 11437
rect 25140 11361 25194 11437
rect 25266 11361 25314 11437
rect 25386 11361 25427 11437
rect 24945 11319 25427 11361
rect 24945 11243 25068 11319
rect 25140 11243 25194 11319
rect 25266 11243 25314 11319
rect 25386 11243 25427 11319
rect 24945 11207 25427 11243
rect 463 11060 863 11109
rect 463 10984 504 11060
rect 576 10984 626 11060
rect 698 10984 752 11060
rect 824 10984 863 11060
rect 463 10913 863 10984
rect 463 10837 504 10913
rect 576 10837 626 10913
rect 698 10837 752 10913
rect 824 10837 863 10913
rect 463 10776 863 10837
rect 463 10700 504 10776
rect 576 10700 626 10776
rect 698 10700 752 10776
rect 824 10700 863 10776
rect 463 10650 863 10700
rect 24946 10256 26370 10281
rect 24946 10180 26010 10256
rect 26082 10180 26136 10256
rect 26208 10180 26256 10256
rect 26328 10180 26370 10256
rect 24946 10138 26370 10180
rect 24946 10062 26010 10138
rect 26082 10062 26136 10138
rect 26208 10062 26256 10138
rect 26328 10062 26370 10138
rect 24946 10026 26370 10062
rect 463 9300 863 9349
rect 463 9224 504 9300
rect 576 9224 626 9300
rect 698 9224 752 9300
rect 824 9224 863 9300
rect 463 9153 863 9224
rect 463 9077 504 9153
rect 576 9077 626 9153
rect 698 9077 752 9153
rect 824 9077 863 9153
rect 463 9016 863 9077
rect 463 8940 504 9016
rect 576 8940 626 9016
rect 698 8940 752 9016
rect 824 8940 863 9016
rect 463 8890 863 8940
rect 463 8621 947 8646
rect 463 8545 503 8621
rect 575 8545 629 8621
rect 701 8545 749 8621
rect 821 8545 947 8621
rect 463 8503 947 8545
rect 463 8427 503 8503
rect 575 8427 629 8503
rect 701 8427 749 8503
rect 821 8427 947 8503
rect 463 8391 947 8427
rect 24946 8594 25428 8619
rect 24946 8518 25068 8594
rect 25140 8518 25194 8594
rect 25266 8518 25314 8594
rect 25386 8518 25428 8594
rect 24946 8476 25428 8518
rect 24946 8400 25068 8476
rect 25140 8400 25194 8476
rect 25266 8400 25314 8476
rect 25386 8400 25428 8476
rect 24946 8364 25428 8400
rect 463 7499 947 7524
rect 463 7423 503 7499
rect 575 7423 629 7499
rect 701 7423 749 7499
rect 821 7423 947 7499
rect 463 7381 947 7423
rect 463 7305 503 7381
rect 575 7305 629 7381
rect 701 7305 749 7381
rect 821 7305 947 7381
rect 463 7269 947 7305
rect 24946 7437 25427 7462
rect 24946 7361 25068 7437
rect 25140 7361 25194 7437
rect 25266 7361 25314 7437
rect 25386 7361 25427 7437
rect 24946 7319 25427 7361
rect 24946 7243 25068 7319
rect 25140 7243 25194 7319
rect 25266 7243 25314 7319
rect 25386 7243 25427 7319
rect 24946 7207 25427 7243
rect 463 7061 863 7110
rect 463 6985 504 7061
rect 576 6985 626 7061
rect 698 6985 752 7061
rect 824 6985 863 7061
rect 463 6914 863 6985
rect 463 6838 504 6914
rect 576 6838 626 6914
rect 698 6838 752 6914
rect 824 6838 863 6914
rect 463 6777 863 6838
rect 463 6701 504 6777
rect 576 6701 626 6777
rect 698 6701 752 6777
rect 824 6701 863 6777
rect 463 6651 863 6701
rect 24946 6292 26370 6317
rect 24946 6216 26010 6292
rect 26082 6216 26136 6292
rect 26208 6216 26256 6292
rect 26328 6216 26370 6292
rect 24946 6174 26370 6216
rect 24946 6098 26010 6174
rect 26082 6098 26136 6174
rect 26208 6098 26256 6174
rect 26328 6098 26370 6174
rect 24946 6062 26370 6098
rect 463 5299 863 5348
rect 463 5223 504 5299
rect 576 5223 626 5299
rect 698 5223 752 5299
rect 824 5223 863 5299
rect 463 5152 863 5223
rect 463 5076 504 5152
rect 576 5076 626 5152
rect 698 5076 752 5152
rect 824 5076 863 5152
rect 463 5015 863 5076
rect 463 4939 504 5015
rect 576 4939 626 5015
rect 698 4939 752 5015
rect 824 4939 863 5015
rect 463 4889 863 4939
rect 463 4639 946 4664
rect 463 4563 503 4639
rect 575 4563 629 4639
rect 701 4563 749 4639
rect 821 4563 946 4639
rect 463 4521 946 4563
rect 463 4445 503 4521
rect 575 4445 629 4521
rect 701 4445 749 4521
rect 821 4445 946 4521
rect 463 4409 946 4445
rect 24946 4594 25428 4619
rect 24946 4518 25068 4594
rect 25140 4518 25194 4594
rect 25266 4518 25314 4594
rect 25386 4518 25428 4594
rect 24946 4476 25428 4518
rect 24946 4400 25068 4476
rect 25140 4400 25194 4476
rect 25266 4400 25314 4476
rect 25386 4400 25428 4476
rect 24946 4364 25428 4400
rect 463 3528 946 3553
rect 463 3452 503 3528
rect 575 3452 629 3528
rect 701 3452 749 3528
rect 821 3452 946 3528
rect 463 3410 946 3452
rect 463 3334 503 3410
rect 575 3334 629 3410
rect 701 3334 749 3410
rect 821 3334 946 3410
rect 463 3298 946 3334
rect 24946 3437 25427 3462
rect 24946 3361 25068 3437
rect 25140 3361 25194 3437
rect 25266 3361 25314 3437
rect 25386 3361 25427 3437
rect 24946 3319 25427 3361
rect 24946 3243 25068 3319
rect 25140 3243 25194 3319
rect 25266 3243 25314 3319
rect 25386 3243 25427 3319
rect 24946 3207 25427 3243
rect 463 3061 863 3110
rect 463 2985 504 3061
rect 576 2985 626 3061
rect 698 2985 752 3061
rect 824 2985 863 3061
rect 463 2914 863 2985
rect 463 2838 504 2914
rect 576 2838 626 2914
rect 698 2838 752 2914
rect 824 2838 863 2914
rect 463 2777 863 2838
rect 463 2701 504 2777
rect 576 2701 626 2777
rect 698 2701 752 2777
rect 824 2701 863 2777
rect 463 2651 863 2701
rect 24946 2280 26370 2305
rect 24946 2204 26010 2280
rect 26082 2204 26136 2280
rect 26208 2204 26256 2280
rect 26328 2204 26370 2280
rect 24946 2162 26370 2204
rect 24946 2086 26010 2162
rect 26082 2086 26136 2162
rect 26208 2086 26256 2162
rect 26328 2086 26370 2162
rect 24946 2050 26370 2086
rect 463 1300 863 1349
rect 463 1224 504 1300
rect 576 1224 626 1300
rect 698 1224 752 1300
rect 824 1224 863 1300
rect 463 1153 863 1224
rect 463 1077 504 1153
rect 576 1077 626 1153
rect 698 1077 752 1153
rect 824 1077 863 1153
rect 463 1016 863 1077
rect 463 940 504 1016
rect 576 940 626 1016
rect 698 940 752 1016
rect 824 940 863 1016
rect 463 890 863 940
rect 463 705 948 730
rect 463 629 503 705
rect 575 629 629 705
rect 701 629 749 705
rect 821 629 948 705
rect 463 587 948 629
rect 463 511 503 587
rect 575 511 629 587
rect 701 511 749 587
rect 821 511 948 587
rect 463 475 948 511
rect 24946 594 25428 619
rect 24946 518 25068 594
rect 25140 518 25194 594
rect 25266 518 25314 594
rect 25386 518 25428 594
rect 24946 476 25428 518
rect 24946 400 25068 476
rect 25140 400 25194 476
rect 25266 400 25314 476
rect 25386 400 25428 476
rect 24946 364 25428 400
<< via1 >>
rect 503 63376 575 63452
rect 629 63376 701 63452
rect 749 63376 821 63452
rect 503 63258 575 63334
rect 629 63258 701 63334
rect 749 63258 821 63334
rect 25068 63416 25140 63492
rect 25194 63416 25266 63492
rect 25314 63416 25386 63492
rect 25068 63298 25140 63374
rect 25194 63298 25266 63374
rect 25314 63298 25386 63374
rect 504 62984 576 63060
rect 626 62984 698 63060
rect 752 62984 824 63060
rect 504 62837 576 62913
rect 626 62837 698 62913
rect 752 62837 824 62913
rect 504 62700 576 62776
rect 626 62700 698 62776
rect 752 62700 824 62776
rect 26010 61995 26082 62071
rect 26136 61995 26208 62071
rect 26256 61995 26328 62071
rect 26010 61877 26082 61953
rect 26136 61877 26208 61953
rect 26256 61877 26328 61953
rect 504 61224 576 61300
rect 626 61224 698 61300
rect 752 61224 824 61300
rect 504 61077 576 61153
rect 626 61077 698 61153
rect 752 61077 824 61153
rect 504 60940 576 61016
rect 626 60940 698 61016
rect 752 60940 824 61016
rect 503 60703 575 60779
rect 629 60703 701 60779
rect 749 60703 821 60779
rect 503 60585 575 60661
rect 629 60585 701 60661
rect 749 60585 821 60661
rect 25068 60619 25140 60695
rect 25194 60619 25266 60695
rect 25314 60619 25386 60695
rect 25068 60501 25140 60577
rect 25194 60501 25266 60577
rect 25314 60501 25386 60577
rect 503 59374 575 59450
rect 629 59374 701 59450
rect 749 59374 821 59450
rect 503 59256 575 59332
rect 629 59256 701 59332
rect 749 59256 821 59332
rect 25068 59416 25140 59492
rect 25194 59416 25266 59492
rect 25314 59416 25386 59492
rect 25068 59298 25140 59374
rect 25194 59298 25266 59374
rect 25314 59298 25386 59374
rect 504 58984 576 59060
rect 626 58984 698 59060
rect 752 58984 824 59060
rect 504 58837 576 58913
rect 626 58837 698 58913
rect 752 58837 824 58913
rect 504 58700 576 58776
rect 626 58700 698 58776
rect 752 58700 824 58776
rect 26010 57982 26082 58058
rect 26136 57982 26208 58058
rect 26256 57982 26328 58058
rect 26010 57864 26082 57940
rect 26136 57864 26208 57940
rect 26256 57864 26328 57940
rect 504 57225 576 57301
rect 626 57225 698 57301
rect 752 57225 824 57301
rect 504 57078 576 57154
rect 626 57078 698 57154
rect 752 57078 824 57154
rect 504 56941 576 57017
rect 626 56941 698 57017
rect 752 56941 824 57017
rect 503 56634 575 56710
rect 629 56634 701 56710
rect 749 56634 821 56710
rect 503 56516 575 56592
rect 629 56516 701 56592
rect 749 56516 821 56592
rect 25068 56619 25140 56695
rect 25194 56619 25266 56695
rect 25314 56619 25386 56695
rect 25068 56501 25140 56577
rect 25194 56501 25266 56577
rect 25314 56501 25386 56577
rect 503 55456 575 55532
rect 629 55456 701 55532
rect 749 55456 821 55532
rect 503 55338 575 55414
rect 629 55338 701 55414
rect 749 55338 821 55414
rect 25068 55416 25140 55492
rect 25194 55416 25266 55492
rect 25314 55416 25386 55492
rect 25068 55298 25140 55374
rect 25194 55298 25266 55374
rect 25314 55298 25386 55374
rect 504 54984 576 55060
rect 626 54984 698 55060
rect 752 54984 824 55060
rect 504 54837 576 54913
rect 626 54837 698 54913
rect 752 54837 824 54913
rect 504 54700 576 54776
rect 626 54700 698 54776
rect 752 54700 824 54776
rect 26010 53981 26082 54057
rect 26136 53981 26208 54057
rect 26256 53981 26328 54057
rect 26010 53863 26082 53939
rect 26136 53863 26208 53939
rect 26256 53863 26328 53939
rect 504 53225 576 53301
rect 626 53225 698 53301
rect 752 53225 824 53301
rect 504 53078 576 53154
rect 626 53078 698 53154
rect 752 53078 824 53154
rect 504 52941 576 53017
rect 626 52941 698 53017
rect 752 52941 824 53017
rect 503 52608 575 52684
rect 629 52608 701 52684
rect 749 52608 821 52684
rect 503 52490 575 52566
rect 629 52490 701 52566
rect 749 52490 821 52566
rect 25068 52619 25140 52695
rect 25194 52619 25266 52695
rect 25314 52619 25386 52695
rect 25068 52501 25140 52577
rect 25194 52501 25266 52577
rect 25314 52501 25386 52577
rect 503 51405 575 51481
rect 629 51405 701 51481
rect 749 51405 821 51481
rect 503 51287 575 51363
rect 629 51287 701 51363
rect 749 51287 821 51363
rect 25068 51470 25140 51546
rect 25194 51470 25266 51546
rect 25314 51470 25386 51546
rect 25068 51352 25140 51428
rect 25194 51352 25266 51428
rect 25314 51352 25386 51428
rect 504 50984 576 51060
rect 626 50984 698 51060
rect 752 50984 824 51060
rect 504 50837 576 50913
rect 626 50837 698 50913
rect 752 50837 824 50913
rect 504 50700 576 50776
rect 626 50700 698 50776
rect 752 50700 824 50776
rect 26010 50020 26082 50096
rect 26136 50020 26208 50096
rect 26256 50020 26328 50096
rect 26010 49902 26082 49978
rect 26136 49902 26208 49978
rect 26256 49902 26328 49978
rect 504 49223 576 49299
rect 626 49223 698 49299
rect 752 49223 824 49299
rect 504 49076 576 49152
rect 626 49076 698 49152
rect 752 49076 824 49152
rect 504 48939 576 49015
rect 626 48939 698 49015
rect 752 48939 824 49015
rect 503 48628 575 48704
rect 629 48628 701 48704
rect 749 48628 821 48704
rect 503 48510 575 48586
rect 629 48510 701 48586
rect 749 48510 821 48586
rect 25068 48554 25140 48630
rect 25194 48554 25266 48630
rect 25314 48554 25386 48630
rect 25068 48436 25140 48512
rect 25194 48436 25266 48512
rect 25314 48436 25386 48512
rect 503 47421 575 47497
rect 629 47421 701 47497
rect 749 47421 821 47497
rect 503 47303 575 47379
rect 629 47303 701 47379
rect 749 47303 821 47379
rect 25068 47371 25140 47447
rect 25194 47371 25266 47447
rect 25314 47371 25386 47447
rect 25068 47253 25140 47329
rect 25194 47253 25266 47329
rect 25314 47253 25386 47329
rect 504 46984 576 47060
rect 626 46984 698 47060
rect 752 46984 824 47060
rect 504 46837 576 46913
rect 626 46837 698 46913
rect 752 46837 824 46913
rect 504 46700 576 46776
rect 626 46700 698 46776
rect 752 46700 824 46776
rect 26010 46003 26082 46079
rect 26136 46003 26208 46079
rect 26256 46003 26328 46079
rect 26010 45885 26082 45961
rect 26136 45885 26208 45961
rect 26256 45885 26328 45961
rect 504 45225 576 45301
rect 626 45225 698 45301
rect 752 45225 824 45301
rect 504 45078 576 45154
rect 626 45078 698 45154
rect 752 45078 824 45154
rect 504 44941 576 45017
rect 626 44941 698 45017
rect 752 44941 824 45017
rect 503 44655 575 44731
rect 629 44655 701 44731
rect 749 44655 821 44731
rect 503 44537 575 44613
rect 629 44537 701 44613
rect 749 44537 821 44613
rect 25068 44499 25140 44575
rect 25194 44499 25266 44575
rect 25314 44499 25386 44575
rect 25068 44381 25140 44457
rect 25194 44381 25266 44457
rect 25314 44381 25386 44457
rect 503 43468 575 43544
rect 629 43468 701 43544
rect 749 43468 821 43544
rect 503 43350 575 43426
rect 629 43350 701 43426
rect 749 43350 821 43426
rect 25068 43364 25140 43440
rect 25194 43364 25266 43440
rect 25314 43364 25386 43440
rect 25068 43246 25140 43322
rect 25194 43246 25266 43322
rect 25314 43246 25386 43322
rect 504 42984 576 43060
rect 626 42984 698 43060
rect 752 42984 824 43060
rect 504 42837 576 42913
rect 626 42837 698 42913
rect 752 42837 824 42913
rect 504 42700 576 42776
rect 626 42700 698 42776
rect 752 42700 824 42776
rect 26010 42082 26082 42158
rect 26136 42082 26208 42158
rect 26256 42082 26328 42158
rect 26010 41964 26082 42040
rect 26136 41964 26208 42040
rect 26256 41964 26328 42040
rect 504 41225 576 41301
rect 626 41225 698 41301
rect 752 41225 824 41301
rect 504 41078 576 41154
rect 626 41078 698 41154
rect 752 41078 824 41154
rect 504 40941 576 41017
rect 626 40941 698 41017
rect 752 40941 824 41017
rect 503 40646 575 40722
rect 629 40646 701 40722
rect 749 40646 821 40722
rect 503 40528 575 40604
rect 629 40528 701 40604
rect 749 40528 821 40604
rect 25068 40605 25140 40681
rect 25194 40605 25266 40681
rect 25314 40605 25386 40681
rect 25068 40487 25140 40563
rect 25194 40487 25266 40563
rect 25314 40487 25386 40563
rect 503 39493 575 39569
rect 629 39493 701 39569
rect 749 39493 821 39569
rect 503 39375 575 39451
rect 629 39375 701 39451
rect 749 39375 821 39451
rect 25068 39452 25140 39528
rect 25194 39452 25266 39528
rect 25314 39452 25386 39528
rect 25068 39334 25140 39410
rect 25194 39334 25266 39410
rect 25314 39334 25386 39410
rect 504 38984 576 39060
rect 626 38984 698 39060
rect 752 38984 824 39060
rect 504 38837 576 38913
rect 626 38837 698 38913
rect 752 38837 824 38913
rect 504 38700 576 38776
rect 626 38700 698 38776
rect 752 38700 824 38776
rect 26010 37824 26082 37900
rect 26136 37824 26208 37900
rect 26256 37824 26328 37900
rect 26010 37706 26082 37782
rect 26136 37706 26208 37782
rect 26256 37706 26328 37782
rect 504 37224 576 37300
rect 626 37224 698 37300
rect 752 37224 824 37300
rect 504 37077 576 37153
rect 626 37077 698 37153
rect 752 37077 824 37153
rect 504 36940 576 37016
rect 626 36940 698 37016
rect 752 36940 824 37016
rect 503 36433 575 36509
rect 629 36433 701 36509
rect 749 36433 821 36509
rect 503 36315 575 36391
rect 629 36315 701 36391
rect 749 36315 821 36391
rect 25068 36336 25140 36412
rect 25194 36336 25266 36412
rect 25314 36336 25386 36412
rect 25068 36218 25140 36294
rect 25194 36218 25266 36294
rect 25314 36218 25386 36294
rect 32 35661 112 35741
rect 157 35661 237 35741
rect 282 35661 362 35741
rect 25535 35646 25615 35726
rect 25660 35646 25740 35726
rect 25785 35646 25865 35726
rect 32 35555 112 35635
rect 157 35555 237 35635
rect 282 35555 362 35635
rect 25534 35526 25614 35606
rect 25659 35526 25739 35606
rect 25784 35526 25864 35606
rect 2020 35273 2062 35315
rect 2062 35273 2072 35315
rect 2020 35263 2072 35273
rect 2098 35274 2108 35316
rect 2108 35274 2150 35316
rect 2098 35264 2150 35274
rect 2021 35225 2073 35235
rect 2021 35183 2063 35225
rect 2063 35183 2073 35225
rect 2099 35226 2151 35236
rect 2099 35184 2109 35226
rect 2109 35184 2151 35226
rect 2262 35279 2304 35321
rect 2304 35279 2314 35321
rect 2262 35269 2314 35279
rect 2332 35279 2342 35321
rect 2342 35279 2384 35321
rect 2332 35269 2384 35279
rect 2485 35281 2603 35395
rect 2641 35281 2759 35395
rect 2797 35281 2915 35395
rect 3151 35286 3193 35328
rect 3193 35286 3203 35328
rect 3151 35276 3203 35286
rect 3221 35286 3231 35328
rect 3231 35286 3273 35328
rect 3221 35276 3273 35286
rect 2262 35241 2314 35251
rect 2262 35199 2304 35241
rect 2304 35199 2314 35241
rect 2332 35241 2384 35251
rect 2332 35199 2342 35241
rect 2342 35199 2384 35241
rect 3151 35248 3203 35258
rect 3151 35206 3193 35248
rect 3193 35206 3203 35248
rect 3221 35248 3273 35258
rect 3221 35206 3231 35248
rect 3231 35206 3273 35248
rect 479 35052 561 35130
rect 593 35052 675 35130
rect 707 35052 789 35130
rect 4129 34870 4181 34880
rect 25061 34892 25141 34972
rect 25186 34892 25266 34972
rect 25311 34892 25391 34972
rect 4129 34836 4153 34870
rect 4153 34836 4181 34870
rect 4129 34828 4181 34836
rect 5210 34871 5262 34879
rect 5210 34836 5215 34871
rect 5215 34836 5250 34871
rect 5250 34836 5262 34871
rect 5210 34827 5262 34836
rect 25060 34772 25140 34852
rect 25185 34772 25265 34852
rect 25310 34772 25390 34852
rect 16 34508 98 34586
rect 130 34508 212 34586
rect 244 34508 326 34586
rect 2071 34260 2123 34269
rect 2071 34225 2079 34260
rect 2079 34225 2115 34260
rect 2115 34225 2123 34260
rect 2071 34217 2123 34225
rect 4208 34296 4260 34348
rect 25069 34316 25141 34392
rect 25191 34316 25263 34392
rect 25317 34316 25389 34392
rect 5252 34258 5304 34267
rect 5252 34224 5262 34258
rect 5262 34224 5296 34258
rect 5296 34224 5304 34258
rect 5252 34215 5304 34224
rect 25069 34169 25141 34245
rect 25191 34169 25263 34245
rect 25317 34169 25389 34245
rect 479 33964 561 34042
rect 593 33964 675 34042
rect 707 33964 789 34042
rect 25069 34032 25141 34108
rect 25191 34032 25263 34108
rect 25317 34032 25389 34108
rect 2063 33782 2115 33790
rect 2063 33748 2081 33782
rect 2081 33748 2115 33782
rect 2063 33738 2115 33748
rect 4123 33845 4175 33897
rect 5252 33782 5304 33791
rect 5252 33748 5262 33782
rect 5262 33748 5296 33782
rect 5296 33748 5304 33782
rect 5252 33739 5304 33748
rect 16 33420 98 33498
rect 130 33420 212 33498
rect 244 33420 326 33498
rect 24560 33396 24640 33476
rect 24685 33396 24765 33476
rect 24810 33396 24890 33476
rect 25535 33396 25615 33476
rect 25660 33396 25740 33476
rect 25785 33396 25865 33476
rect 2283 33310 2286 33358
rect 2286 33310 2332 33358
rect 2332 33310 2335 33358
rect 2283 33306 2335 33310
rect 2283 33245 2335 33252
rect 2283 33200 2286 33245
rect 2286 33200 2332 33245
rect 2332 33200 2335 33245
rect 24559 33276 24639 33356
rect 24684 33276 24764 33356
rect 24809 33276 24889 33356
rect 25534 33276 25614 33356
rect 25659 33276 25739 33356
rect 25784 33276 25864 33356
rect 4153 33170 4205 33182
rect 4153 33136 4187 33170
rect 4187 33136 4205 33170
rect 4153 33130 4205 33136
rect 5209 33170 5261 33181
rect 5209 33136 5215 33170
rect 5215 33136 5249 33170
rect 5249 33136 5261 33170
rect 5209 33129 5261 33136
rect 479 32876 561 32954
rect 593 32876 675 32954
rect 707 32876 789 32954
rect 3151 32788 3193 32830
rect 3193 32788 3203 32830
rect 3151 32778 3203 32788
rect 3221 32788 3231 32830
rect 3231 32788 3273 32830
rect 3221 32778 3273 32788
rect 3151 32750 3203 32763
rect 3151 32711 3193 32750
rect 3193 32711 3203 32750
rect 3221 32750 3273 32763
rect 3221 32711 3231 32750
rect 3231 32711 3273 32750
rect 3365 32788 3407 32830
rect 3407 32788 3417 32830
rect 3365 32778 3417 32788
rect 3435 32788 3445 32830
rect 3445 32788 3487 32830
rect 3435 32778 3487 32788
rect 3365 32747 3417 32765
rect 3365 32713 3407 32747
rect 3407 32713 3417 32747
rect 3435 32747 3487 32765
rect 3435 32713 3445 32747
rect 3445 32713 3487 32747
rect 25069 32556 25141 32632
rect 25191 32556 25263 32632
rect 25317 32556 25389 32632
rect 25069 32409 25141 32485
rect 25191 32409 25263 32485
rect 25317 32409 25389 32485
rect 25069 32272 25141 32348
rect 25191 32272 25263 32348
rect 25317 32272 25389 32348
rect 25060 31837 25140 31917
rect 25185 31837 25265 31917
rect 25310 31837 25390 31917
rect 25059 31717 25139 31797
rect 25184 31717 25264 31797
rect 25309 31717 25389 31797
rect 503 28226 575 28302
rect 629 28226 701 28302
rect 749 28226 821 28302
rect 25068 28226 25140 28302
rect 25194 28226 25266 28302
rect 25314 28226 25386 28302
rect 503 28108 575 28184
rect 629 28108 701 28184
rect 749 28108 821 28184
rect 25068 28108 25140 28184
rect 25194 28108 25266 28184
rect 25314 28108 25386 28184
rect 503 27444 575 27520
rect 629 27444 701 27520
rect 749 27444 821 27520
rect 503 27326 575 27402
rect 629 27326 701 27402
rect 749 27326 821 27402
rect 25068 27444 25140 27520
rect 25194 27444 25266 27520
rect 25314 27444 25386 27520
rect 25068 27326 25140 27402
rect 25194 27326 25266 27402
rect 25314 27326 25386 27402
rect 504 26985 576 27061
rect 626 26985 698 27061
rect 752 26985 824 27061
rect 504 26838 576 26914
rect 626 26838 698 26914
rect 752 26838 824 26914
rect 504 26701 576 26777
rect 626 26701 698 26777
rect 752 26701 824 26777
rect 26010 26054 26082 26130
rect 26136 26054 26208 26130
rect 26256 26054 26328 26130
rect 26010 25936 26082 26012
rect 26136 25936 26208 26012
rect 26256 25936 26328 26012
rect 504 25218 576 25294
rect 626 25218 698 25294
rect 752 25218 824 25294
rect 504 25071 576 25147
rect 626 25071 698 25147
rect 752 25071 824 25147
rect 504 24934 576 25010
rect 626 24934 698 25010
rect 752 24934 824 25010
rect 503 24532 575 24608
rect 629 24532 701 24608
rect 749 24532 821 24608
rect 503 24414 575 24490
rect 629 24414 701 24490
rect 749 24414 821 24490
rect 25068 24483 25140 24559
rect 25194 24483 25266 24559
rect 25314 24483 25386 24559
rect 25068 24365 25140 24441
rect 25194 24365 25266 24441
rect 25314 24365 25386 24441
rect 503 23528 575 23604
rect 629 23528 701 23604
rect 749 23528 821 23604
rect 503 23410 575 23486
rect 629 23410 701 23486
rect 749 23410 821 23486
rect 25068 23366 25140 23442
rect 25194 23366 25266 23442
rect 25314 23366 25386 23442
rect 25068 23248 25140 23324
rect 25194 23248 25266 23324
rect 25314 23248 25386 23324
rect 504 22984 576 23060
rect 626 22984 698 23060
rect 752 22984 824 23060
rect 504 22837 576 22913
rect 626 22837 698 22913
rect 752 22837 824 22913
rect 504 22700 576 22776
rect 626 22700 698 22776
rect 752 22700 824 22776
rect 26010 21895 26082 21971
rect 26136 21895 26208 21971
rect 26256 21895 26328 21971
rect 26010 21777 26082 21853
rect 26136 21777 26208 21853
rect 26256 21777 26328 21853
rect 504 21224 576 21300
rect 626 21224 698 21300
rect 752 21224 824 21300
rect 504 21077 576 21153
rect 626 21077 698 21153
rect 752 21077 824 21153
rect 504 20940 576 21016
rect 626 20940 698 21016
rect 752 20940 824 21016
rect 503 20550 575 20626
rect 629 20550 701 20626
rect 749 20550 821 20626
rect 503 20432 575 20508
rect 629 20432 701 20508
rect 749 20432 821 20508
rect 25068 20523 25140 20599
rect 25194 20523 25266 20599
rect 25314 20523 25386 20599
rect 25068 20405 25140 20481
rect 25194 20405 25266 20481
rect 25314 20405 25386 20481
rect 503 19468 575 19544
rect 629 19468 701 19544
rect 749 19468 821 19544
rect 503 19350 575 19426
rect 629 19350 701 19426
rect 749 19350 821 19426
rect 25068 19348 25140 19424
rect 25194 19348 25266 19424
rect 25314 19348 25386 19424
rect 25068 19230 25140 19306
rect 25194 19230 25266 19306
rect 25314 19230 25386 19306
rect 504 18984 576 19060
rect 626 18984 698 19060
rect 752 18984 824 19060
rect 504 18837 576 18913
rect 626 18837 698 18913
rect 752 18837 824 18913
rect 504 18700 576 18776
rect 626 18700 698 18776
rect 752 18700 824 18776
rect 26010 18105 26082 18181
rect 26136 18105 26208 18181
rect 26256 18105 26328 18181
rect 26010 17987 26082 18063
rect 26136 17987 26208 18063
rect 26256 17987 26328 18063
rect 504 17225 576 17301
rect 626 17225 698 17301
rect 752 17225 824 17301
rect 504 17078 576 17154
rect 626 17078 698 17154
rect 752 17078 824 17154
rect 504 16941 576 17017
rect 626 16941 698 17017
rect 752 16941 824 17017
rect 503 16593 575 16669
rect 629 16593 701 16669
rect 749 16593 821 16669
rect 503 16475 575 16551
rect 629 16475 701 16551
rect 749 16475 821 16551
rect 25068 16507 25140 16583
rect 25194 16507 25266 16583
rect 25314 16507 25386 16583
rect 25068 16389 25140 16465
rect 25194 16389 25266 16465
rect 25314 16389 25386 16465
rect 503 15492 575 15568
rect 629 15492 701 15568
rect 749 15492 821 15568
rect 503 15374 575 15450
rect 629 15374 701 15450
rect 749 15374 821 15450
rect 25068 15336 25140 15412
rect 25194 15336 25266 15412
rect 25314 15336 25386 15412
rect 25068 15218 25140 15294
rect 25194 15218 25266 15294
rect 25314 15218 25386 15294
rect 504 14984 576 15060
rect 626 14984 698 15060
rect 752 14984 824 15060
rect 504 14837 576 14913
rect 626 14837 698 14913
rect 752 14837 824 14913
rect 504 14700 576 14776
rect 626 14700 698 14776
rect 752 14700 824 14776
rect 26010 13998 26082 14074
rect 26136 13998 26208 14074
rect 26256 13998 26328 14074
rect 26010 13880 26082 13956
rect 26136 13880 26208 13956
rect 26256 13880 26328 13956
rect 504 13224 576 13300
rect 626 13224 698 13300
rect 752 13224 824 13300
rect 504 13077 576 13153
rect 626 13077 698 13153
rect 752 13077 824 13153
rect 504 12940 576 13016
rect 626 12940 698 13016
rect 752 12940 824 13016
rect 503 12626 575 12702
rect 629 12626 701 12702
rect 749 12626 821 12702
rect 503 12508 575 12584
rect 629 12508 701 12584
rect 749 12508 821 12584
rect 25068 12575 25140 12651
rect 25194 12575 25266 12651
rect 25314 12575 25386 12651
rect 25068 12457 25140 12533
rect 25194 12457 25266 12533
rect 25314 12457 25386 12533
rect 503 11410 575 11486
rect 629 11410 701 11486
rect 749 11410 821 11486
rect 503 11292 575 11368
rect 629 11292 701 11368
rect 749 11292 821 11368
rect 25068 11361 25140 11437
rect 25194 11361 25266 11437
rect 25314 11361 25386 11437
rect 25068 11243 25140 11319
rect 25194 11243 25266 11319
rect 25314 11243 25386 11319
rect 504 10984 576 11060
rect 626 10984 698 11060
rect 752 10984 824 11060
rect 504 10837 576 10913
rect 626 10837 698 10913
rect 752 10837 824 10913
rect 504 10700 576 10776
rect 626 10700 698 10776
rect 752 10700 824 10776
rect 26010 10180 26082 10256
rect 26136 10180 26208 10256
rect 26256 10180 26328 10256
rect 26010 10062 26082 10138
rect 26136 10062 26208 10138
rect 26256 10062 26328 10138
rect 504 9224 576 9300
rect 626 9224 698 9300
rect 752 9224 824 9300
rect 504 9077 576 9153
rect 626 9077 698 9153
rect 752 9077 824 9153
rect 504 8940 576 9016
rect 626 8940 698 9016
rect 752 8940 824 9016
rect 503 8545 575 8621
rect 629 8545 701 8621
rect 749 8545 821 8621
rect 503 8427 575 8503
rect 629 8427 701 8503
rect 749 8427 821 8503
rect 25068 8518 25140 8594
rect 25194 8518 25266 8594
rect 25314 8518 25386 8594
rect 25068 8400 25140 8476
rect 25194 8400 25266 8476
rect 25314 8400 25386 8476
rect 503 7423 575 7499
rect 629 7423 701 7499
rect 749 7423 821 7499
rect 503 7305 575 7381
rect 629 7305 701 7381
rect 749 7305 821 7381
rect 25068 7361 25140 7437
rect 25194 7361 25266 7437
rect 25314 7361 25386 7437
rect 25068 7243 25140 7319
rect 25194 7243 25266 7319
rect 25314 7243 25386 7319
rect 504 6985 576 7061
rect 626 6985 698 7061
rect 752 6985 824 7061
rect 504 6838 576 6914
rect 626 6838 698 6914
rect 752 6838 824 6914
rect 504 6701 576 6777
rect 626 6701 698 6777
rect 752 6701 824 6777
rect 26010 6216 26082 6292
rect 26136 6216 26208 6292
rect 26256 6216 26328 6292
rect 26010 6098 26082 6174
rect 26136 6098 26208 6174
rect 26256 6098 26328 6174
rect 504 5223 576 5299
rect 626 5223 698 5299
rect 752 5223 824 5299
rect 504 5076 576 5152
rect 626 5076 698 5152
rect 752 5076 824 5152
rect 504 4939 576 5015
rect 626 4939 698 5015
rect 752 4939 824 5015
rect 503 4563 575 4639
rect 629 4563 701 4639
rect 749 4563 821 4639
rect 503 4445 575 4521
rect 629 4445 701 4521
rect 749 4445 821 4521
rect 25068 4518 25140 4594
rect 25194 4518 25266 4594
rect 25314 4518 25386 4594
rect 25068 4400 25140 4476
rect 25194 4400 25266 4476
rect 25314 4400 25386 4476
rect 503 3452 575 3528
rect 629 3452 701 3528
rect 749 3452 821 3528
rect 503 3334 575 3410
rect 629 3334 701 3410
rect 749 3334 821 3410
rect 25068 3361 25140 3437
rect 25194 3361 25266 3437
rect 25314 3361 25386 3437
rect 25068 3243 25140 3319
rect 25194 3243 25266 3319
rect 25314 3243 25386 3319
rect 504 2985 576 3061
rect 626 2985 698 3061
rect 752 2985 824 3061
rect 504 2838 576 2914
rect 626 2838 698 2914
rect 752 2838 824 2914
rect 504 2701 576 2777
rect 626 2701 698 2777
rect 752 2701 824 2777
rect 26010 2204 26082 2280
rect 26136 2204 26208 2280
rect 26256 2204 26328 2280
rect 26010 2086 26082 2162
rect 26136 2086 26208 2162
rect 26256 2086 26328 2162
rect 504 1224 576 1300
rect 626 1224 698 1300
rect 752 1224 824 1300
rect 504 1077 576 1153
rect 626 1077 698 1153
rect 752 1077 824 1153
rect 504 940 576 1016
rect 626 940 698 1016
rect 752 940 824 1016
rect 503 629 575 705
rect 629 629 701 705
rect 749 629 821 705
rect 503 511 575 587
rect 629 511 701 587
rect 749 511 821 587
rect 25068 518 25140 594
rect 25194 518 25266 594
rect 25314 518 25386 594
rect 25068 400 25140 476
rect 25194 400 25266 476
rect 25314 400 25386 476
<< metal2 >>
rect 25026 63492 25426 63517
rect 463 63452 864 63477
rect 463 63376 503 63452
rect 575 63376 629 63452
rect 701 63376 749 63452
rect 821 63376 864 63452
rect 463 63334 864 63376
rect 463 63258 503 63334
rect 575 63258 629 63334
rect 701 63258 749 63334
rect 821 63258 864 63334
rect 25026 63416 25068 63492
rect 25140 63416 25194 63492
rect 25266 63416 25314 63492
rect 25386 63416 25426 63492
rect 25026 63374 25426 63416
rect 25026 63298 25068 63374
rect 25140 63298 25194 63374
rect 25266 63298 25314 63374
rect 25386 63298 25426 63374
rect 25026 63262 25426 63298
rect 463 63222 864 63258
rect 463 63060 863 63109
rect 463 62984 504 63060
rect 576 62984 626 63060
rect 698 62984 752 63060
rect 824 62984 863 63060
rect 463 62913 863 62984
rect 463 62837 504 62913
rect 576 62837 626 62913
rect 698 62837 752 62913
rect 824 62837 863 62913
rect 463 62776 863 62837
rect 463 62700 504 62776
rect 576 62700 626 62776
rect 698 62700 752 62776
rect 824 62700 863 62776
rect 463 62650 863 62700
rect 25970 62071 26370 62096
rect 25970 61995 26010 62071
rect 26082 61995 26136 62071
rect 26208 61995 26256 62071
rect 26328 61995 26370 62071
rect 25970 61953 26370 61995
rect 25970 61877 26010 61953
rect 26082 61877 26136 61953
rect 26208 61877 26256 61953
rect 26328 61877 26370 61953
rect 25970 61841 26370 61877
rect 463 61300 863 61349
rect 463 61224 504 61300
rect 576 61224 626 61300
rect 698 61224 752 61300
rect 824 61224 863 61300
rect 463 61153 863 61224
rect 463 61077 504 61153
rect 576 61077 626 61153
rect 698 61077 752 61153
rect 824 61077 863 61153
rect 463 61016 863 61077
rect 463 60940 504 61016
rect 576 60940 626 61016
rect 698 60940 752 61016
rect 824 60940 863 61016
rect 463 60890 863 60940
rect 463 60779 864 60804
rect 463 60703 503 60779
rect 575 60703 629 60779
rect 701 60703 749 60779
rect 821 60703 864 60779
rect 463 60661 864 60703
rect 463 60585 503 60661
rect 575 60585 629 60661
rect 701 60585 749 60661
rect 821 60585 864 60661
rect 463 60549 864 60585
rect 25028 60695 25428 60720
rect 25028 60619 25068 60695
rect 25140 60619 25194 60695
rect 25266 60619 25314 60695
rect 25386 60619 25428 60695
rect 25028 60577 25428 60619
rect 25028 60501 25068 60577
rect 25140 60501 25194 60577
rect 25266 60501 25314 60577
rect 25386 60501 25428 60577
rect 25028 60465 25428 60501
rect 25026 59492 25426 59517
rect 463 59450 864 59475
rect 463 59374 503 59450
rect 575 59374 629 59450
rect 701 59374 749 59450
rect 821 59374 864 59450
rect 463 59332 864 59374
rect 463 59256 503 59332
rect 575 59256 629 59332
rect 701 59256 749 59332
rect 821 59256 864 59332
rect 25026 59416 25068 59492
rect 25140 59416 25194 59492
rect 25266 59416 25314 59492
rect 25386 59416 25426 59492
rect 25026 59374 25426 59416
rect 25026 59298 25068 59374
rect 25140 59298 25194 59374
rect 25266 59298 25314 59374
rect 25386 59298 25426 59374
rect 25026 59262 25426 59298
rect 463 59220 864 59256
rect 463 59060 863 59109
rect 463 58984 504 59060
rect 576 58984 626 59060
rect 698 58984 752 59060
rect 824 58984 863 59060
rect 463 58913 863 58984
rect 463 58837 504 58913
rect 576 58837 626 58913
rect 698 58837 752 58913
rect 824 58837 863 58913
rect 463 58776 863 58837
rect 463 58700 504 58776
rect 576 58700 626 58776
rect 698 58700 752 58776
rect 824 58700 863 58776
rect 463 58650 863 58700
rect 25970 58058 26370 58083
rect 25970 57982 26010 58058
rect 26082 57982 26136 58058
rect 26208 57982 26256 58058
rect 26328 57982 26370 58058
rect 25970 57940 26370 57982
rect 25970 57864 26010 57940
rect 26082 57864 26136 57940
rect 26208 57864 26256 57940
rect 26328 57864 26370 57940
rect 25970 57828 26370 57864
rect 463 57301 863 57350
rect 463 57225 504 57301
rect 576 57225 626 57301
rect 698 57225 752 57301
rect 824 57225 863 57301
rect 463 57154 863 57225
rect 463 57078 504 57154
rect 576 57078 626 57154
rect 698 57078 752 57154
rect 824 57078 863 57154
rect 463 57017 863 57078
rect 463 56941 504 57017
rect 576 56941 626 57017
rect 698 56941 752 57017
rect 824 56941 863 57017
rect 463 56891 863 56941
rect 463 56710 864 56735
rect 463 56634 503 56710
rect 575 56634 629 56710
rect 701 56634 749 56710
rect 821 56634 864 56710
rect 463 56592 864 56634
rect 463 56516 503 56592
rect 575 56516 629 56592
rect 701 56516 749 56592
rect 821 56516 864 56592
rect 463 56480 864 56516
rect 25028 56695 25428 56720
rect 25028 56619 25068 56695
rect 25140 56619 25194 56695
rect 25266 56619 25314 56695
rect 25386 56619 25428 56695
rect 25028 56577 25428 56619
rect 25028 56501 25068 56577
rect 25140 56501 25194 56577
rect 25266 56501 25314 56577
rect 25386 56501 25428 56577
rect 25028 56465 25428 56501
rect 463 55532 864 55557
rect 463 55456 503 55532
rect 575 55456 629 55532
rect 701 55456 749 55532
rect 821 55456 864 55532
rect 463 55414 864 55456
rect 463 55338 503 55414
rect 575 55338 629 55414
rect 701 55338 749 55414
rect 821 55338 864 55414
rect 463 55302 864 55338
rect 25026 55492 25426 55517
rect 25026 55416 25068 55492
rect 25140 55416 25194 55492
rect 25266 55416 25314 55492
rect 25386 55416 25426 55492
rect 25026 55374 25426 55416
rect 25026 55298 25068 55374
rect 25140 55298 25194 55374
rect 25266 55298 25314 55374
rect 25386 55298 25426 55374
rect 25026 55262 25426 55298
rect 464 55068 864 55109
rect 463 55060 864 55068
rect 463 54984 504 55060
rect 576 54984 626 55060
rect 698 54984 752 55060
rect 824 54984 864 55060
rect 463 54913 864 54984
rect 463 54837 504 54913
rect 576 54837 626 54913
rect 698 54837 752 54913
rect 824 54837 864 54913
rect 463 54776 864 54837
rect 463 54700 504 54776
rect 576 54700 626 54776
rect 698 54700 752 54776
rect 824 54700 864 54776
rect 463 54650 864 54700
rect 25970 54057 26370 54082
rect 25970 53981 26010 54057
rect 26082 53981 26136 54057
rect 26208 53981 26256 54057
rect 26328 53981 26370 54057
rect 25970 53939 26370 53981
rect 25970 53863 26010 53939
rect 26082 53863 26136 53939
rect 26208 53863 26256 53939
rect 26328 53863 26370 53939
rect 25970 53827 26370 53863
rect 463 53301 863 53350
rect 463 53225 504 53301
rect 576 53225 626 53301
rect 698 53225 752 53301
rect 824 53225 863 53301
rect 463 53154 863 53225
rect 463 53078 504 53154
rect 576 53078 626 53154
rect 698 53078 752 53154
rect 824 53078 863 53154
rect 463 53017 863 53078
rect 463 52941 504 53017
rect 576 52941 626 53017
rect 698 52941 752 53017
rect 824 52941 863 53017
rect 463 52891 863 52941
rect 463 52684 866 52709
rect 463 52608 503 52684
rect 575 52608 629 52684
rect 701 52608 749 52684
rect 821 52608 866 52684
rect 463 52566 866 52608
rect 463 52490 503 52566
rect 575 52490 629 52566
rect 701 52490 749 52566
rect 821 52490 866 52566
rect 463 52454 866 52490
rect 25028 52695 25428 52720
rect 25028 52619 25068 52695
rect 25140 52619 25194 52695
rect 25266 52619 25314 52695
rect 25386 52619 25428 52695
rect 25028 52577 25428 52619
rect 25028 52501 25068 52577
rect 25140 52501 25194 52577
rect 25266 52501 25314 52577
rect 25386 52501 25428 52577
rect 25028 52465 25428 52501
rect 25027 51546 25427 51571
rect 463 51481 864 51506
rect 463 51405 503 51481
rect 575 51405 629 51481
rect 701 51405 749 51481
rect 821 51405 864 51481
rect 463 51363 864 51405
rect 463 51287 503 51363
rect 575 51287 629 51363
rect 701 51287 749 51363
rect 821 51287 864 51363
rect 25027 51470 25068 51546
rect 25140 51470 25194 51546
rect 25266 51470 25314 51546
rect 25386 51470 25427 51546
rect 25027 51428 25427 51470
rect 25027 51352 25068 51428
rect 25140 51352 25194 51428
rect 25266 51352 25314 51428
rect 25386 51352 25427 51428
rect 25027 51316 25427 51352
rect 463 51251 864 51287
rect 464 51068 864 51109
rect 463 51060 864 51068
rect 463 50984 504 51060
rect 576 50984 626 51060
rect 698 50984 752 51060
rect 824 50984 864 51060
rect 463 50913 864 50984
rect 463 50837 504 50913
rect 576 50837 626 50913
rect 698 50837 752 50913
rect 824 50837 864 50913
rect 463 50776 864 50837
rect 463 50700 504 50776
rect 576 50700 626 50776
rect 698 50700 752 50776
rect 824 50700 864 50776
rect 463 50650 864 50700
rect 25970 50096 26370 50121
rect 25970 50020 26010 50096
rect 26082 50020 26136 50096
rect 26208 50020 26256 50096
rect 26328 50020 26370 50096
rect 25970 49978 26370 50020
rect 25970 49902 26010 49978
rect 26082 49902 26136 49978
rect 26208 49902 26256 49978
rect 26328 49902 26370 49978
rect 25970 49866 26370 49902
rect 463 49299 863 49348
rect 463 49223 504 49299
rect 576 49223 626 49299
rect 698 49223 752 49299
rect 824 49223 863 49299
rect 463 49152 863 49223
rect 463 49076 504 49152
rect 576 49076 626 49152
rect 698 49076 752 49152
rect 824 49076 863 49152
rect 463 49015 863 49076
rect 463 48939 504 49015
rect 576 48939 626 49015
rect 698 48939 752 49015
rect 824 48939 863 49015
rect 463 48889 863 48939
rect 463 48704 864 48729
rect 463 48628 503 48704
rect 575 48628 629 48704
rect 701 48628 749 48704
rect 821 48628 864 48704
rect 463 48586 864 48628
rect 463 48510 503 48586
rect 575 48510 629 48586
rect 701 48510 749 48586
rect 821 48510 864 48586
rect 463 48474 864 48510
rect 25028 48630 25428 48655
rect 25028 48554 25068 48630
rect 25140 48554 25194 48630
rect 25266 48554 25314 48630
rect 25386 48554 25428 48630
rect 25028 48512 25428 48554
rect 25028 48436 25068 48512
rect 25140 48436 25194 48512
rect 25266 48436 25314 48512
rect 25386 48436 25428 48512
rect 25028 48400 25428 48436
rect 463 47497 866 47522
rect 463 47421 503 47497
rect 575 47421 629 47497
rect 701 47421 749 47497
rect 821 47421 866 47497
rect 463 47379 866 47421
rect 463 47303 503 47379
rect 575 47303 629 47379
rect 701 47303 749 47379
rect 821 47303 866 47379
rect 463 47267 866 47303
rect 25027 47447 25427 47472
rect 25027 47371 25068 47447
rect 25140 47371 25194 47447
rect 25266 47371 25314 47447
rect 25386 47371 25427 47447
rect 25027 47329 25427 47371
rect 25027 47253 25068 47329
rect 25140 47253 25194 47329
rect 25266 47253 25314 47329
rect 25386 47253 25427 47329
rect 25027 47217 25427 47253
rect 463 47060 863 47109
rect 463 46984 504 47060
rect 576 46984 626 47060
rect 698 46984 752 47060
rect 824 46984 863 47060
rect 463 46913 863 46984
rect 463 46837 504 46913
rect 576 46837 626 46913
rect 698 46837 752 46913
rect 824 46837 863 46913
rect 463 46776 863 46837
rect 463 46700 504 46776
rect 576 46700 626 46776
rect 698 46700 752 46776
rect 824 46700 863 46776
rect 463 46650 863 46700
rect 25970 46079 26370 46104
rect 25970 46003 26010 46079
rect 26082 46003 26136 46079
rect 26208 46003 26256 46079
rect 26328 46003 26370 46079
rect 25970 45961 26370 46003
rect 25970 45885 26010 45961
rect 26082 45885 26136 45961
rect 26208 45885 26256 45961
rect 26328 45885 26370 45961
rect 25970 45849 26370 45885
rect 463 45301 863 45350
rect 463 45225 504 45301
rect 576 45225 626 45301
rect 698 45225 752 45301
rect 824 45225 863 45301
rect 463 45154 863 45225
rect 463 45078 504 45154
rect 576 45078 626 45154
rect 698 45078 752 45154
rect 824 45078 863 45154
rect 463 45017 863 45078
rect 463 44941 504 45017
rect 576 44941 626 45017
rect 698 44941 752 45017
rect 824 44941 863 45017
rect 463 44891 863 44941
rect 463 44731 864 44756
rect 463 44655 503 44731
rect 575 44655 629 44731
rect 701 44655 749 44731
rect 821 44655 864 44731
rect 463 44613 864 44655
rect 463 44537 503 44613
rect 575 44537 629 44613
rect 701 44537 749 44613
rect 821 44537 864 44613
rect 463 44501 864 44537
rect 25028 44575 25428 44600
rect 25028 44499 25068 44575
rect 25140 44499 25194 44575
rect 25266 44499 25314 44575
rect 25386 44499 25428 44575
rect 25028 44457 25428 44499
rect 25028 44381 25068 44457
rect 25140 44381 25194 44457
rect 25266 44381 25314 44457
rect 25386 44381 25428 44457
rect 25028 44345 25428 44381
rect 463 43544 864 43569
rect 463 43468 503 43544
rect 575 43468 629 43544
rect 701 43468 749 43544
rect 821 43468 864 43544
rect 463 43426 864 43468
rect 463 43350 503 43426
rect 575 43350 629 43426
rect 701 43350 749 43426
rect 821 43350 864 43426
rect 463 43314 864 43350
rect 25028 43440 25428 43465
rect 25028 43364 25068 43440
rect 25140 43364 25194 43440
rect 25266 43364 25314 43440
rect 25386 43364 25428 43440
rect 25028 43322 25428 43364
rect 25028 43246 25068 43322
rect 25140 43246 25194 43322
rect 25266 43246 25314 43322
rect 25386 43246 25428 43322
rect 25028 43210 25428 43246
rect 463 43060 863 43109
rect 463 42984 504 43060
rect 576 42984 626 43060
rect 698 42984 752 43060
rect 824 42984 863 43060
rect 463 42913 863 42984
rect 463 42837 504 42913
rect 576 42837 626 42913
rect 698 42837 752 42913
rect 824 42837 863 42913
rect 463 42776 863 42837
rect 463 42700 504 42776
rect 576 42700 626 42776
rect 698 42700 752 42776
rect 824 42700 863 42776
rect 463 42650 863 42700
rect 25970 42158 26370 42183
rect 25970 42082 26010 42158
rect 26082 42082 26136 42158
rect 26208 42082 26256 42158
rect 26328 42082 26370 42158
rect 25970 42040 26370 42082
rect 25970 41964 26010 42040
rect 26082 41964 26136 42040
rect 26208 41964 26256 42040
rect 26328 41964 26370 42040
rect 25970 41928 26370 41964
rect 463 41301 863 41350
rect 463 41225 504 41301
rect 576 41225 626 41301
rect 698 41225 752 41301
rect 824 41225 863 41301
rect 463 41154 863 41225
rect 463 41078 504 41154
rect 576 41078 626 41154
rect 698 41078 752 41154
rect 824 41078 863 41154
rect 463 41017 863 41078
rect 463 40941 504 41017
rect 576 40941 626 41017
rect 698 40941 752 41017
rect 824 40941 863 41017
rect 463 40891 863 40941
rect 463 40722 864 40747
rect 463 40646 503 40722
rect 575 40646 629 40722
rect 701 40646 749 40722
rect 821 40646 864 40722
rect 463 40604 864 40646
rect 463 40528 503 40604
rect 575 40528 629 40604
rect 701 40528 749 40604
rect 821 40528 864 40604
rect 463 40492 864 40528
rect 25028 40681 25428 40706
rect 25028 40605 25068 40681
rect 25140 40605 25194 40681
rect 25266 40605 25314 40681
rect 25386 40605 25428 40681
rect 25028 40563 25428 40605
rect 25028 40487 25068 40563
rect 25140 40487 25194 40563
rect 25266 40487 25314 40563
rect 25386 40487 25428 40563
rect 25028 40451 25428 40487
rect 463 39569 864 39594
rect 463 39493 503 39569
rect 575 39493 629 39569
rect 701 39493 749 39569
rect 821 39493 864 39569
rect 463 39451 864 39493
rect 463 39375 503 39451
rect 575 39375 629 39451
rect 701 39375 749 39451
rect 821 39375 864 39451
rect 463 39339 864 39375
rect 25028 39528 25428 39553
rect 25028 39452 25068 39528
rect 25140 39452 25194 39528
rect 25266 39452 25314 39528
rect 25386 39452 25428 39528
rect 25028 39410 25428 39452
rect 25028 39334 25068 39410
rect 25140 39334 25194 39410
rect 25266 39334 25314 39410
rect 25386 39334 25428 39410
rect 25028 39298 25428 39334
rect 463 39060 863 39109
rect 463 38984 504 39060
rect 576 38984 626 39060
rect 698 38984 752 39060
rect 824 38984 863 39060
rect 463 38913 863 38984
rect 463 38837 504 38913
rect 576 38837 626 38913
rect 698 38837 752 38913
rect 824 38837 863 38913
rect 463 38776 863 38837
rect 463 38700 504 38776
rect 576 38700 626 38776
rect 698 38700 752 38776
rect 824 38700 863 38776
rect 463 38650 863 38700
rect 25970 37900 26370 37925
rect 25970 37824 26010 37900
rect 26082 37824 26136 37900
rect 26208 37824 26256 37900
rect 26328 37824 26370 37900
rect 25970 37782 26370 37824
rect 25970 37706 26010 37782
rect 26082 37706 26136 37782
rect 26208 37706 26256 37782
rect 26328 37706 26370 37782
rect 25970 37670 26370 37706
rect 463 37300 863 37350
rect 463 37224 504 37300
rect 576 37224 626 37300
rect 698 37224 752 37300
rect 824 37224 863 37300
rect 463 37153 863 37224
rect 463 37077 504 37153
rect 576 37077 626 37153
rect 698 37077 752 37153
rect 824 37077 863 37153
rect 463 37016 863 37077
rect 463 36940 504 37016
rect 576 36940 626 37016
rect 698 36940 752 37016
rect 824 36940 863 37016
rect 463 36891 863 36940
rect 463 36890 836 36891
rect 463 36509 863 36534
rect 463 36433 503 36509
rect 575 36433 629 36509
rect 701 36433 749 36509
rect 821 36433 863 36509
rect 463 36391 863 36433
rect 463 36315 503 36391
rect 575 36315 629 36391
rect 701 36315 749 36391
rect 821 36315 863 36391
rect 463 36279 863 36315
rect 25028 36412 25428 36437
rect 25028 36336 25068 36412
rect 25140 36336 25194 36412
rect 25266 36336 25314 36412
rect 25386 36336 25428 36412
rect 25028 36294 25428 36336
rect 25028 36218 25068 36294
rect 25140 36218 25194 36294
rect 25266 36218 25314 36294
rect 25386 36218 25428 36294
rect 25028 36182 25428 36218
rect 2248 35925 2398 35940
rect 2248 35869 2257 35925
rect 2313 35869 2337 35925
rect 2393 35869 2398 35925
rect 2248 35845 2398 35869
rect 2248 35789 2257 35845
rect 2313 35789 2337 35845
rect 2393 35789 2398 35845
rect 2248 35776 2398 35789
rect 0 35741 400 35752
rect 0 35661 32 35741
rect 112 35661 157 35741
rect 237 35661 282 35741
rect 362 35661 400 35741
rect 0 35635 400 35661
rect 0 35555 32 35635
rect 112 35555 157 35635
rect 237 35555 282 35635
rect 362 35555 400 35635
rect 0 35528 400 35555
rect 2011 35320 2160 35333
rect 2011 35319 2098 35320
rect 2011 35263 2016 35319
rect 2072 35264 2098 35319
rect 2154 35264 2160 35320
rect 2072 35263 2160 35264
rect 2011 35240 2160 35263
rect 2011 35239 2099 35240
rect 2011 35183 2017 35239
rect 2073 35184 2099 35239
rect 2155 35184 2160 35240
rect 2250 35321 2396 35776
rect 2468 35459 2867 36000
rect 2467 35410 2867 35459
rect 3352 35904 3502 35919
rect 3352 35848 3361 35904
rect 3417 35848 3441 35904
rect 3497 35848 3502 35904
rect 3352 35824 3502 35848
rect 3352 35768 3361 35824
rect 3417 35768 3441 35824
rect 3497 35768 3502 35824
rect 3352 35755 3502 35768
rect 3352 35754 3500 35755
rect 3352 35449 3499 35754
rect 25502 35726 25902 35752
rect 25502 35646 25535 35726
rect 25615 35646 25660 35726
rect 25740 35646 25785 35726
rect 25865 35646 25902 35726
rect 25502 35606 25902 35646
rect 25502 35526 25534 35606
rect 25614 35526 25659 35606
rect 25739 35526 25784 35606
rect 25864 35526 25902 35606
rect 25502 35497 25902 35526
rect 2250 35269 2262 35321
rect 2314 35269 2332 35321
rect 2384 35269 2396 35321
rect 2250 35251 2396 35269
rect 2250 35199 2262 35251
rect 2314 35199 2332 35251
rect 2384 35199 2396 35251
rect 2250 35189 2396 35199
rect 2468 35395 2935 35410
rect 2468 35281 2485 35395
rect 2603 35281 2641 35395
rect 2759 35281 2797 35395
rect 2915 35281 2935 35395
rect 2468 35270 2935 35281
rect 3138 35328 3285 35336
rect 3138 35276 3151 35328
rect 3203 35276 3221 35328
rect 3273 35276 3285 35328
rect 2073 35183 2160 35184
rect 2011 35169 2160 35183
rect 463 35130 805 35139
rect 463 35052 479 35130
rect 561 35052 593 35130
rect 675 35052 707 35130
rect 789 35052 805 35130
rect 463 35043 805 35052
rect 0 34586 342 34595
rect 0 34508 16 34586
rect 98 34508 130 34586
rect 212 34508 244 34586
rect 326 34508 342 34586
rect 0 34499 342 34508
rect 2071 34269 2123 34275
rect 2071 34211 2123 34217
rect 463 34042 805 34051
rect 463 33964 479 34042
rect 561 33964 593 34042
rect 675 33964 707 34042
rect 789 33964 805 34042
rect 463 33955 805 33964
rect 2071 33797 2104 34211
rect 2063 33790 2115 33797
rect 2063 33732 2115 33738
rect 0 33498 342 33507
rect 0 33420 16 33498
rect 98 33420 130 33498
rect 212 33420 244 33498
rect 326 33420 342 33498
rect 0 33411 342 33420
rect 2280 33358 2339 35189
rect 2280 33306 2283 33358
rect 2335 33306 2339 33358
rect 2280 33252 2339 33306
rect 2280 33200 2283 33252
rect 2335 33200 2339 33252
rect 2280 33187 2339 33200
rect 463 32954 805 32963
rect 463 32876 479 32954
rect 561 32876 593 32954
rect 675 32876 707 32954
rect 789 32876 805 32954
rect 463 32867 805 32876
rect 463 28302 866 28360
rect 463 28226 503 28302
rect 575 28226 629 28302
rect 701 28226 749 28302
rect 821 28226 866 28302
rect 463 28184 866 28226
rect 463 28108 503 28184
rect 575 28108 629 28184
rect 701 28108 749 28184
rect 821 28108 866 28184
rect 463 28072 866 28108
rect 2468 28000 2867 35270
rect 3138 35258 3285 35276
rect 3138 35206 3151 35258
rect 3203 35206 3221 35258
rect 3273 35206 3285 35258
rect 3351 35318 3499 35449
rect 3351 35262 3360 35318
rect 3416 35317 3499 35318
rect 3416 35262 3440 35317
rect 3351 35261 3440 35262
rect 3496 35261 3499 35317
rect 3351 35253 3499 35261
rect 3138 32830 3285 35206
rect 3138 32778 3151 32830
rect 3203 32778 3221 32830
rect 3273 32778 3285 32830
rect 3138 32763 3285 32778
rect 3138 32711 3151 32763
rect 3203 32711 3221 32763
rect 3273 32711 3285 32763
rect 3138 32476 3285 32711
rect 3352 35237 3499 35253
rect 3352 35181 3361 35237
rect 3417 35181 3441 35237
rect 3497 35181 3499 35237
rect 3352 32830 3499 35181
rect 25028 34972 25428 34998
rect 25028 34892 25061 34972
rect 25141 34892 25186 34972
rect 25266 34892 25311 34972
rect 25391 34892 25428 34972
rect 4123 34828 4129 34880
rect 4181 34828 4187 34880
rect 5210 34879 5304 34885
rect 4137 33897 4168 34828
rect 5262 34827 5304 34879
rect 5210 34821 5304 34827
rect 4208 34348 4260 34354
rect 4208 34290 4260 34296
rect 4117 33845 4123 33897
rect 4175 33845 4181 33897
rect 4220 33185 4249 34290
rect 5252 34267 5304 34821
rect 25028 34852 25428 34892
rect 25028 34772 25060 34852
rect 25140 34772 25185 34852
rect 25265 34772 25310 34852
rect 25390 34772 25428 34852
rect 25028 34743 25428 34772
rect 5252 34209 5304 34215
rect 25028 34392 25428 34442
rect 25028 34316 25069 34392
rect 25141 34316 25191 34392
rect 25263 34316 25317 34392
rect 25389 34316 25428 34392
rect 25028 34245 25428 34316
rect 25028 34169 25069 34245
rect 25141 34169 25191 34245
rect 25263 34169 25317 34245
rect 25389 34169 25428 34245
rect 25028 34108 25428 34169
rect 25028 34032 25069 34108
rect 25141 34032 25191 34108
rect 25263 34032 25317 34108
rect 25389 34032 25428 34108
rect 25028 33983 25428 34032
rect 25028 33982 25401 33983
rect 5252 33791 5304 33797
rect 5252 33187 5304 33739
rect 24527 33476 24927 33502
rect 24527 33396 24560 33476
rect 24640 33396 24685 33476
rect 24765 33396 24810 33476
rect 24890 33396 24927 33476
rect 24527 33356 24927 33396
rect 24527 33276 24559 33356
rect 24639 33276 24684 33356
rect 24764 33276 24809 33356
rect 24889 33276 24927 33356
rect 24527 33247 24927 33276
rect 25502 33476 25902 33502
rect 25502 33396 25535 33476
rect 25615 33396 25660 33476
rect 25740 33396 25785 33476
rect 25865 33396 25902 33476
rect 25502 33356 25902 33396
rect 25502 33276 25534 33356
rect 25614 33276 25659 33356
rect 25739 33276 25784 33356
rect 25864 33276 25902 33356
rect 25502 33247 25902 33276
rect 4136 33182 4249 33185
rect 4136 33130 4153 33182
rect 4205 33130 4249 33182
rect 4136 33126 4249 33130
rect 5209 33181 5304 33187
rect 5261 33129 5304 33181
rect 5209 33123 5304 33129
rect 3352 32778 3365 32830
rect 3417 32778 3435 32830
rect 3487 32778 3499 32830
rect 3352 32765 3499 32778
rect 3352 32713 3365 32765
rect 3417 32713 3435 32765
rect 3487 32713 3499 32765
rect 3352 32707 3499 32713
rect 3135 32475 3285 32476
rect 25028 32632 25428 32682
rect 25028 32556 25069 32632
rect 25141 32556 25191 32632
rect 25263 32556 25317 32632
rect 25389 32556 25428 32632
rect 25028 32485 25428 32556
rect 3135 32463 3289 32475
rect 3135 32401 3144 32463
rect 3200 32401 3224 32463
rect 3280 32401 3289 32463
rect 3135 32391 3289 32401
rect 25028 32409 25069 32485
rect 25141 32409 25191 32485
rect 25263 32409 25317 32485
rect 25389 32409 25428 32485
rect 25028 32348 25428 32409
rect 25028 32272 25069 32348
rect 25141 32272 25191 32348
rect 25263 32272 25317 32348
rect 25389 32272 25428 32348
rect 25028 32223 25428 32272
rect 25028 32222 25401 32223
rect 25027 31917 25427 31943
rect 25027 31837 25060 31917
rect 25140 31837 25185 31917
rect 25265 31837 25310 31917
rect 25390 31837 25427 31917
rect 25027 31797 25427 31837
rect 25027 31717 25059 31797
rect 25139 31717 25184 31797
rect 25264 31717 25309 31797
rect 25389 31717 25427 31797
rect 25027 31688 25427 31717
rect 25025 28302 25428 28360
rect 25025 28226 25068 28302
rect 25140 28226 25194 28302
rect 25266 28226 25314 28302
rect 25386 28226 25428 28302
rect 25025 28184 25428 28226
rect 25025 28108 25068 28184
rect 25140 28108 25194 28184
rect 25266 28108 25314 28184
rect 25386 28108 25428 28184
rect 25025 28072 25428 28108
rect 463 27520 863 27545
rect 463 27444 503 27520
rect 575 27444 629 27520
rect 701 27444 749 27520
rect 821 27444 863 27520
rect 463 27402 863 27444
rect 463 27326 503 27402
rect 575 27326 629 27402
rect 701 27326 749 27402
rect 821 27326 863 27402
rect 463 27290 863 27326
rect 25028 27520 25428 27545
rect 25028 27444 25068 27520
rect 25140 27444 25194 27520
rect 25266 27444 25314 27520
rect 25386 27444 25428 27520
rect 25028 27402 25428 27444
rect 25028 27326 25068 27402
rect 25140 27326 25194 27402
rect 25266 27326 25314 27402
rect 25386 27326 25428 27402
rect 25028 27290 25428 27326
rect 463 27061 863 27111
rect 463 26985 504 27061
rect 576 26985 626 27061
rect 698 26985 752 27061
rect 824 26985 863 27061
rect 463 26914 863 26985
rect 463 26838 504 26914
rect 576 26838 626 26914
rect 698 26838 752 26914
rect 824 26838 863 26914
rect 463 26777 863 26838
rect 463 26701 504 26777
rect 576 26701 626 26777
rect 698 26701 752 26777
rect 824 26701 863 26777
rect 463 26651 863 26701
rect 25970 26130 26370 26155
rect 25970 26054 26010 26130
rect 26082 26054 26136 26130
rect 26208 26054 26256 26130
rect 26328 26054 26370 26130
rect 25970 26012 26370 26054
rect 25970 25936 26010 26012
rect 26082 25936 26136 26012
rect 26208 25936 26256 26012
rect 26328 25936 26370 26012
rect 25970 25900 26370 25936
rect 463 25294 863 25349
rect 463 25218 504 25294
rect 576 25218 626 25294
rect 698 25218 752 25294
rect 824 25218 863 25294
rect 463 25147 863 25218
rect 463 25071 504 25147
rect 576 25071 626 25147
rect 698 25071 752 25147
rect 824 25071 863 25147
rect 463 25010 863 25071
rect 463 24934 504 25010
rect 576 24934 626 25010
rect 698 24934 752 25010
rect 824 24934 863 25010
rect 463 24885 863 24934
rect 463 24884 862 24885
rect 463 24608 863 24633
rect 463 24532 503 24608
rect 575 24532 629 24608
rect 701 24532 749 24608
rect 821 24532 863 24608
rect 463 24490 863 24532
rect 463 24414 503 24490
rect 575 24414 629 24490
rect 701 24414 749 24490
rect 821 24414 863 24490
rect 463 24378 863 24414
rect 25028 24559 25428 24584
rect 25028 24483 25068 24559
rect 25140 24483 25194 24559
rect 25266 24483 25314 24559
rect 25386 24483 25428 24559
rect 25028 24441 25428 24483
rect 25028 24365 25068 24441
rect 25140 24365 25194 24441
rect 25266 24365 25314 24441
rect 25386 24365 25428 24441
rect 25028 24329 25428 24365
rect 463 23604 863 23629
rect 463 23528 503 23604
rect 575 23528 629 23604
rect 701 23528 749 23604
rect 821 23528 863 23604
rect 463 23486 863 23528
rect 463 23410 503 23486
rect 575 23410 629 23486
rect 701 23410 749 23486
rect 821 23410 863 23486
rect 463 23374 863 23410
rect 25027 23442 25427 23467
rect 25027 23366 25068 23442
rect 25140 23366 25194 23442
rect 25266 23366 25314 23442
rect 25386 23366 25427 23442
rect 25027 23324 25427 23366
rect 25027 23248 25068 23324
rect 25140 23248 25194 23324
rect 25266 23248 25314 23324
rect 25386 23248 25427 23324
rect 25027 23212 25427 23248
rect 463 23060 863 23109
rect 463 22984 504 23060
rect 576 22984 626 23060
rect 698 22984 752 23060
rect 824 22984 863 23060
rect 463 22913 863 22984
rect 463 22837 504 22913
rect 576 22837 626 22913
rect 698 22837 752 22913
rect 824 22837 863 22913
rect 463 22776 863 22837
rect 463 22700 504 22776
rect 576 22700 626 22776
rect 698 22700 752 22776
rect 824 22700 863 22776
rect 463 22650 863 22700
rect 25970 21971 26370 21996
rect 25970 21895 26010 21971
rect 26082 21895 26136 21971
rect 26208 21895 26256 21971
rect 26328 21895 26370 21971
rect 25970 21853 26370 21895
rect 25970 21777 26010 21853
rect 26082 21777 26136 21853
rect 26208 21777 26256 21853
rect 26328 21777 26370 21853
rect 25970 21741 26370 21777
rect 463 21300 863 21349
rect 463 21224 504 21300
rect 576 21224 626 21300
rect 698 21224 752 21300
rect 824 21224 863 21300
rect 463 21153 863 21224
rect 463 21077 504 21153
rect 576 21077 626 21153
rect 698 21077 752 21153
rect 824 21077 863 21153
rect 463 21016 863 21077
rect 463 20940 504 21016
rect 576 20940 626 21016
rect 698 20940 752 21016
rect 824 20940 863 21016
rect 463 20890 863 20940
rect 463 20626 864 20651
rect 463 20550 503 20626
rect 575 20550 629 20626
rect 701 20550 749 20626
rect 821 20550 864 20626
rect 463 20508 864 20550
rect 463 20432 503 20508
rect 575 20432 629 20508
rect 701 20432 749 20508
rect 821 20432 864 20508
rect 463 20396 864 20432
rect 25028 20599 25428 20624
rect 25028 20523 25068 20599
rect 25140 20523 25194 20599
rect 25266 20523 25314 20599
rect 25386 20523 25428 20599
rect 25028 20481 25428 20523
rect 25028 20405 25068 20481
rect 25140 20405 25194 20481
rect 25266 20405 25314 20481
rect 25386 20405 25428 20481
rect 25028 20369 25428 20405
rect 463 19544 864 19569
rect 463 19468 503 19544
rect 575 19468 629 19544
rect 701 19468 749 19544
rect 821 19468 864 19544
rect 463 19426 864 19468
rect 463 19350 503 19426
rect 575 19350 629 19426
rect 701 19350 749 19426
rect 821 19350 864 19426
rect 463 19314 864 19350
rect 25028 19424 25428 19449
rect 25028 19348 25068 19424
rect 25140 19348 25194 19424
rect 25266 19348 25314 19424
rect 25386 19348 25428 19424
rect 25028 19306 25428 19348
rect 25028 19230 25068 19306
rect 25140 19230 25194 19306
rect 25266 19230 25314 19306
rect 25386 19230 25428 19306
rect 25028 19194 25428 19230
rect 463 19060 863 19109
rect 463 18984 504 19060
rect 576 18984 626 19060
rect 698 18984 752 19060
rect 824 18984 863 19060
rect 463 18913 863 18984
rect 463 18837 504 18913
rect 576 18837 626 18913
rect 698 18837 752 18913
rect 824 18837 863 18913
rect 463 18776 863 18837
rect 463 18700 504 18776
rect 576 18700 626 18776
rect 698 18700 752 18776
rect 824 18700 863 18776
rect 463 18650 863 18700
rect 25970 18181 26370 18206
rect 25970 18105 26010 18181
rect 26082 18105 26136 18181
rect 26208 18105 26256 18181
rect 26328 18105 26370 18181
rect 25970 18063 26370 18105
rect 25970 17987 26010 18063
rect 26082 17987 26136 18063
rect 26208 17987 26256 18063
rect 26328 17987 26370 18063
rect 25970 17951 26370 17987
rect 463 17301 863 17350
rect 463 17225 504 17301
rect 576 17225 626 17301
rect 698 17225 752 17301
rect 824 17225 863 17301
rect 463 17154 863 17225
rect 463 17078 504 17154
rect 576 17078 626 17154
rect 698 17078 752 17154
rect 824 17078 863 17154
rect 463 17017 863 17078
rect 463 16941 504 17017
rect 576 16941 626 17017
rect 698 16941 752 17017
rect 824 16941 863 17017
rect 463 16891 863 16941
rect 463 16669 864 16694
rect 463 16593 503 16669
rect 575 16593 629 16669
rect 701 16593 749 16669
rect 821 16593 864 16669
rect 463 16551 864 16593
rect 463 16475 503 16551
rect 575 16475 629 16551
rect 701 16475 749 16551
rect 821 16475 864 16551
rect 463 16439 864 16475
rect 25027 16583 25427 16608
rect 25027 16507 25068 16583
rect 25140 16507 25194 16583
rect 25266 16507 25314 16583
rect 25386 16507 25427 16583
rect 25027 16465 25427 16507
rect 25027 16389 25068 16465
rect 25140 16389 25194 16465
rect 25266 16389 25314 16465
rect 25386 16389 25427 16465
rect 25027 16353 25427 16389
rect 463 15568 864 15593
rect 463 15492 503 15568
rect 575 15492 629 15568
rect 701 15492 749 15568
rect 821 15492 864 15568
rect 463 15450 864 15492
rect 463 15374 503 15450
rect 575 15374 629 15450
rect 701 15374 749 15450
rect 821 15374 864 15450
rect 463 15338 864 15374
rect 25027 15412 25427 15437
rect 25027 15336 25068 15412
rect 25140 15336 25194 15412
rect 25266 15336 25314 15412
rect 25386 15336 25427 15412
rect 25027 15294 25427 15336
rect 25027 15218 25068 15294
rect 25140 15218 25194 15294
rect 25266 15218 25314 15294
rect 25386 15218 25427 15294
rect 25027 15182 25427 15218
rect 463 15060 863 15109
rect 463 14984 504 15060
rect 576 14984 626 15060
rect 698 14984 752 15060
rect 824 14984 863 15060
rect 463 14913 863 14984
rect 463 14837 504 14913
rect 576 14837 626 14913
rect 698 14837 752 14913
rect 824 14837 863 14913
rect 463 14776 863 14837
rect 463 14700 504 14776
rect 576 14700 626 14776
rect 698 14700 752 14776
rect 824 14700 863 14776
rect 463 14650 863 14700
rect 25970 14074 26370 14099
rect 25970 13998 26010 14074
rect 26082 13998 26136 14074
rect 26208 13998 26256 14074
rect 26328 13998 26370 14074
rect 25970 13956 26370 13998
rect 25970 13880 26010 13956
rect 26082 13880 26136 13956
rect 26208 13880 26256 13956
rect 26328 13880 26370 13956
rect 25970 13844 26370 13880
rect 463 13300 863 13349
rect 463 13224 504 13300
rect 576 13224 626 13300
rect 698 13224 752 13300
rect 824 13224 863 13300
rect 463 13153 863 13224
rect 463 13077 504 13153
rect 576 13077 626 13153
rect 698 13077 752 13153
rect 824 13077 863 13153
rect 463 13016 863 13077
rect 463 12940 504 13016
rect 576 12940 626 13016
rect 698 12940 752 13016
rect 824 12940 863 13016
rect 463 12890 863 12940
rect 463 12702 865 12727
rect 463 12626 503 12702
rect 575 12626 629 12702
rect 701 12626 749 12702
rect 821 12626 865 12702
rect 463 12584 865 12626
rect 463 12508 503 12584
rect 575 12508 629 12584
rect 701 12508 749 12584
rect 821 12508 865 12584
rect 463 12472 865 12508
rect 25027 12651 25427 12676
rect 25027 12575 25068 12651
rect 25140 12575 25194 12651
rect 25266 12575 25314 12651
rect 25386 12575 25427 12651
rect 25027 12533 25427 12575
rect 25027 12457 25068 12533
rect 25140 12457 25194 12533
rect 25266 12457 25314 12533
rect 25386 12457 25427 12533
rect 25027 12421 25427 12457
rect 463 11486 866 11511
rect 463 11410 503 11486
rect 575 11410 629 11486
rect 701 11410 749 11486
rect 821 11410 866 11486
rect 463 11368 866 11410
rect 463 11292 503 11368
rect 575 11292 629 11368
rect 701 11292 749 11368
rect 821 11292 866 11368
rect 463 11256 866 11292
rect 25027 11437 25427 11462
rect 25027 11361 25068 11437
rect 25140 11361 25194 11437
rect 25266 11361 25314 11437
rect 25386 11361 25427 11437
rect 25027 11319 25427 11361
rect 25027 11243 25068 11319
rect 25140 11243 25194 11319
rect 25266 11243 25314 11319
rect 25386 11243 25427 11319
rect 25027 11207 25427 11243
rect 463 11060 863 11109
rect 463 10984 504 11060
rect 576 10984 626 11060
rect 698 10984 752 11060
rect 824 10984 863 11060
rect 463 10913 863 10984
rect 463 10837 504 10913
rect 576 10837 626 10913
rect 698 10837 752 10913
rect 824 10837 863 10913
rect 463 10776 863 10837
rect 463 10700 504 10776
rect 576 10700 626 10776
rect 698 10700 752 10776
rect 824 10700 863 10776
rect 463 10650 863 10700
rect 25970 10256 26370 10281
rect 25970 10180 26010 10256
rect 26082 10180 26136 10256
rect 26208 10180 26256 10256
rect 26328 10180 26370 10256
rect 25970 10138 26370 10180
rect 25970 10062 26010 10138
rect 26082 10062 26136 10138
rect 26208 10062 26256 10138
rect 26328 10062 26370 10138
rect 25970 10026 26370 10062
rect 463 9300 863 9349
rect 463 9224 504 9300
rect 576 9224 626 9300
rect 698 9224 752 9300
rect 824 9224 863 9300
rect 463 9153 863 9224
rect 463 9077 504 9153
rect 576 9077 626 9153
rect 698 9077 752 9153
rect 824 9077 863 9153
rect 463 9016 863 9077
rect 463 8940 504 9016
rect 576 8940 626 9016
rect 698 8940 752 9016
rect 824 8940 863 9016
rect 463 8890 863 8940
rect 463 8621 864 8646
rect 463 8545 503 8621
rect 575 8545 629 8621
rect 701 8545 749 8621
rect 821 8545 864 8621
rect 463 8503 864 8545
rect 463 8427 503 8503
rect 575 8427 629 8503
rect 701 8427 749 8503
rect 821 8427 864 8503
rect 463 8391 864 8427
rect 25028 8594 25428 8619
rect 25028 8518 25068 8594
rect 25140 8518 25194 8594
rect 25266 8518 25314 8594
rect 25386 8518 25428 8594
rect 25028 8476 25428 8518
rect 25028 8400 25068 8476
rect 25140 8400 25194 8476
rect 25266 8400 25314 8476
rect 25386 8400 25428 8476
rect 25028 8364 25428 8400
rect 463 7499 864 7524
rect 463 7423 503 7499
rect 575 7423 629 7499
rect 701 7423 749 7499
rect 821 7423 864 7499
rect 463 7381 864 7423
rect 463 7305 503 7381
rect 575 7305 629 7381
rect 701 7305 749 7381
rect 821 7305 864 7381
rect 463 7269 864 7305
rect 25027 7437 25427 7462
rect 25027 7361 25068 7437
rect 25140 7361 25194 7437
rect 25266 7361 25314 7437
rect 25386 7361 25427 7437
rect 25027 7319 25427 7361
rect 25027 7243 25068 7319
rect 25140 7243 25194 7319
rect 25266 7243 25314 7319
rect 25386 7243 25427 7319
rect 25027 7207 25427 7243
rect 463 7061 863 7110
rect 463 6985 504 7061
rect 576 6985 626 7061
rect 698 6985 752 7061
rect 824 6985 863 7061
rect 463 6914 863 6985
rect 463 6838 504 6914
rect 576 6838 626 6914
rect 698 6838 752 6914
rect 824 6838 863 6914
rect 463 6777 863 6838
rect 463 6701 504 6777
rect 576 6701 626 6777
rect 698 6701 752 6777
rect 824 6701 863 6777
rect 463 6651 863 6701
rect 25970 6292 26370 6317
rect 25970 6216 26010 6292
rect 26082 6216 26136 6292
rect 26208 6216 26256 6292
rect 26328 6216 26370 6292
rect 25970 6174 26370 6216
rect 25970 6098 26010 6174
rect 26082 6098 26136 6174
rect 26208 6098 26256 6174
rect 26328 6098 26370 6174
rect 25970 6062 26370 6098
rect 463 5299 863 5348
rect 463 5223 504 5299
rect 576 5223 626 5299
rect 698 5223 752 5299
rect 824 5223 863 5299
rect 463 5152 863 5223
rect 463 5076 504 5152
rect 576 5076 626 5152
rect 698 5076 752 5152
rect 824 5076 863 5152
rect 463 5015 863 5076
rect 463 4939 504 5015
rect 576 4939 626 5015
rect 698 4939 752 5015
rect 824 4939 863 5015
rect 463 4889 863 4939
rect 463 4639 863 4664
rect 463 4563 503 4639
rect 575 4563 629 4639
rect 701 4563 749 4639
rect 821 4563 863 4639
rect 463 4521 863 4563
rect 463 4445 503 4521
rect 575 4445 629 4521
rect 701 4445 749 4521
rect 821 4445 863 4521
rect 463 4409 863 4445
rect 25028 4594 25428 4619
rect 25028 4518 25068 4594
rect 25140 4518 25194 4594
rect 25266 4518 25314 4594
rect 25386 4518 25428 4594
rect 25028 4476 25428 4518
rect 25028 4400 25068 4476
rect 25140 4400 25194 4476
rect 25266 4400 25314 4476
rect 25386 4400 25428 4476
rect 25028 4364 25428 4400
rect 463 3528 863 3553
rect 463 3452 503 3528
rect 575 3452 629 3528
rect 701 3452 749 3528
rect 821 3452 863 3528
rect 463 3410 863 3452
rect 463 3334 503 3410
rect 575 3334 629 3410
rect 701 3334 749 3410
rect 821 3334 863 3410
rect 463 3298 863 3334
rect 25027 3437 25427 3462
rect 25027 3361 25068 3437
rect 25140 3361 25194 3437
rect 25266 3361 25314 3437
rect 25386 3361 25427 3437
rect 25027 3319 25427 3361
rect 25027 3243 25068 3319
rect 25140 3243 25194 3319
rect 25266 3243 25314 3319
rect 25386 3243 25427 3319
rect 25027 3207 25427 3243
rect 463 3061 863 3110
rect 463 2985 504 3061
rect 576 2985 626 3061
rect 698 2985 752 3061
rect 824 2985 863 3061
rect 463 2914 863 2985
rect 463 2838 504 2914
rect 576 2838 626 2914
rect 698 2838 752 2914
rect 824 2838 863 2914
rect 463 2777 863 2838
rect 463 2701 504 2777
rect 576 2701 626 2777
rect 698 2701 752 2777
rect 824 2701 863 2777
rect 463 2651 863 2701
rect 25970 2280 26370 2305
rect 25970 2204 26010 2280
rect 26082 2204 26136 2280
rect 26208 2204 26256 2280
rect 26328 2204 26370 2280
rect 25970 2162 26370 2204
rect 25970 2086 26010 2162
rect 26082 2086 26136 2162
rect 26208 2086 26256 2162
rect 26328 2086 26370 2162
rect 25970 2050 26370 2086
rect 463 1300 863 1349
rect 463 1224 504 1300
rect 576 1224 626 1300
rect 698 1224 752 1300
rect 824 1224 863 1300
rect 463 1153 863 1224
rect 463 1077 504 1153
rect 576 1077 626 1153
rect 698 1077 752 1153
rect 824 1077 863 1153
rect 463 1016 863 1077
rect 463 940 504 1016
rect 576 940 626 1016
rect 698 940 752 1016
rect 824 940 863 1016
rect 463 890 863 940
rect 463 705 865 730
rect 463 629 503 705
rect 575 629 629 705
rect 701 629 749 705
rect 821 629 865 705
rect 463 587 865 629
rect 463 511 503 587
rect 575 511 629 587
rect 701 511 749 587
rect 821 511 865 587
rect 463 475 865 511
rect 25028 594 25428 619
rect 25028 518 25068 594
rect 25140 518 25194 594
rect 25266 518 25314 594
rect 25386 518 25428 594
rect 25028 476 25428 518
rect 25028 400 25068 476
rect 25140 400 25194 476
rect 25266 400 25314 476
rect 25386 400 25428 476
rect 25028 364 25428 400
<< via2 >>
rect 503 63376 575 63452
rect 629 63376 701 63452
rect 749 63376 821 63452
rect 503 63258 575 63334
rect 629 63258 701 63334
rect 749 63258 821 63334
rect 25068 63416 25140 63492
rect 25194 63416 25266 63492
rect 25314 63416 25386 63492
rect 25068 63298 25140 63374
rect 25194 63298 25266 63374
rect 25314 63298 25386 63374
rect 504 62984 576 63060
rect 626 62984 698 63060
rect 752 62984 824 63060
rect 504 62837 576 62913
rect 626 62837 698 62913
rect 752 62837 824 62913
rect 504 62700 576 62776
rect 626 62700 698 62776
rect 752 62700 824 62776
rect 26010 61995 26082 62071
rect 26136 61995 26208 62071
rect 26256 61995 26328 62071
rect 26010 61877 26082 61953
rect 26136 61877 26208 61953
rect 26256 61877 26328 61953
rect 504 61224 576 61300
rect 626 61224 698 61300
rect 752 61224 824 61300
rect 504 61077 576 61153
rect 626 61077 698 61153
rect 752 61077 824 61153
rect 504 60940 576 61016
rect 626 60940 698 61016
rect 752 60940 824 61016
rect 503 60703 575 60779
rect 629 60703 701 60779
rect 749 60703 821 60779
rect 503 60585 575 60661
rect 629 60585 701 60661
rect 749 60585 821 60661
rect 25068 60619 25140 60695
rect 25194 60619 25266 60695
rect 25314 60619 25386 60695
rect 25068 60501 25140 60577
rect 25194 60501 25266 60577
rect 25314 60501 25386 60577
rect 503 59374 575 59450
rect 629 59374 701 59450
rect 749 59374 821 59450
rect 503 59256 575 59332
rect 629 59256 701 59332
rect 749 59256 821 59332
rect 25068 59416 25140 59492
rect 25194 59416 25266 59492
rect 25314 59416 25386 59492
rect 25068 59298 25140 59374
rect 25194 59298 25266 59374
rect 25314 59298 25386 59374
rect 504 58984 576 59060
rect 626 58984 698 59060
rect 752 58984 824 59060
rect 504 58837 576 58913
rect 626 58837 698 58913
rect 752 58837 824 58913
rect 504 58700 576 58776
rect 626 58700 698 58776
rect 752 58700 824 58776
rect 26010 57982 26082 58058
rect 26136 57982 26208 58058
rect 26256 57982 26328 58058
rect 26010 57864 26082 57940
rect 26136 57864 26208 57940
rect 26256 57864 26328 57940
rect 504 57225 576 57301
rect 626 57225 698 57301
rect 752 57225 824 57301
rect 504 57078 576 57154
rect 626 57078 698 57154
rect 752 57078 824 57154
rect 504 56941 576 57017
rect 626 56941 698 57017
rect 752 56941 824 57017
rect 503 56634 575 56710
rect 629 56634 701 56710
rect 749 56634 821 56710
rect 503 56516 575 56592
rect 629 56516 701 56592
rect 749 56516 821 56592
rect 25068 56619 25140 56695
rect 25194 56619 25266 56695
rect 25314 56619 25386 56695
rect 25068 56501 25140 56577
rect 25194 56501 25266 56577
rect 25314 56501 25386 56577
rect 503 55456 575 55532
rect 629 55456 701 55532
rect 749 55456 821 55532
rect 503 55338 575 55414
rect 629 55338 701 55414
rect 749 55338 821 55414
rect 25068 55416 25140 55492
rect 25194 55416 25266 55492
rect 25314 55416 25386 55492
rect 25068 55298 25140 55374
rect 25194 55298 25266 55374
rect 25314 55298 25386 55374
rect 504 54984 576 55060
rect 626 54984 698 55060
rect 752 54984 824 55060
rect 504 54837 576 54913
rect 626 54837 698 54913
rect 752 54837 824 54913
rect 504 54700 576 54776
rect 626 54700 698 54776
rect 752 54700 824 54776
rect 26010 53981 26082 54057
rect 26136 53981 26208 54057
rect 26256 53981 26328 54057
rect 26010 53863 26082 53939
rect 26136 53863 26208 53939
rect 26256 53863 26328 53939
rect 504 53225 576 53301
rect 626 53225 698 53301
rect 752 53225 824 53301
rect 504 53078 576 53154
rect 626 53078 698 53154
rect 752 53078 824 53154
rect 504 52941 576 53017
rect 626 52941 698 53017
rect 752 52941 824 53017
rect 503 52608 575 52684
rect 629 52608 701 52684
rect 749 52608 821 52684
rect 503 52490 575 52566
rect 629 52490 701 52566
rect 749 52490 821 52566
rect 25068 52619 25140 52695
rect 25194 52619 25266 52695
rect 25314 52619 25386 52695
rect 25068 52501 25140 52577
rect 25194 52501 25266 52577
rect 25314 52501 25386 52577
rect 503 51405 575 51481
rect 629 51405 701 51481
rect 749 51405 821 51481
rect 503 51287 575 51363
rect 629 51287 701 51363
rect 749 51287 821 51363
rect 25068 51470 25140 51546
rect 25194 51470 25266 51546
rect 25314 51470 25386 51546
rect 25068 51352 25140 51428
rect 25194 51352 25266 51428
rect 25314 51352 25386 51428
rect 504 50984 576 51060
rect 626 50984 698 51060
rect 752 50984 824 51060
rect 504 50837 576 50913
rect 626 50837 698 50913
rect 752 50837 824 50913
rect 504 50700 576 50776
rect 626 50700 698 50776
rect 752 50700 824 50776
rect 26010 50020 26082 50096
rect 26136 50020 26208 50096
rect 26256 50020 26328 50096
rect 26010 49902 26082 49978
rect 26136 49902 26208 49978
rect 26256 49902 26328 49978
rect 504 49223 576 49299
rect 626 49223 698 49299
rect 752 49223 824 49299
rect 504 49076 576 49152
rect 626 49076 698 49152
rect 752 49076 824 49152
rect 504 48939 576 49015
rect 626 48939 698 49015
rect 752 48939 824 49015
rect 503 48628 575 48704
rect 629 48628 701 48704
rect 749 48628 821 48704
rect 503 48510 575 48586
rect 629 48510 701 48586
rect 749 48510 821 48586
rect 25068 48554 25140 48630
rect 25194 48554 25266 48630
rect 25314 48554 25386 48630
rect 25068 48436 25140 48512
rect 25194 48436 25266 48512
rect 25314 48436 25386 48512
rect 503 47421 575 47497
rect 629 47421 701 47497
rect 749 47421 821 47497
rect 503 47303 575 47379
rect 629 47303 701 47379
rect 749 47303 821 47379
rect 25068 47371 25140 47447
rect 25194 47371 25266 47447
rect 25314 47371 25386 47447
rect 25068 47253 25140 47329
rect 25194 47253 25266 47329
rect 25314 47253 25386 47329
rect 504 46984 576 47060
rect 626 46984 698 47060
rect 752 46984 824 47060
rect 504 46837 576 46913
rect 626 46837 698 46913
rect 752 46837 824 46913
rect 504 46700 576 46776
rect 626 46700 698 46776
rect 752 46700 824 46776
rect 26010 46003 26082 46079
rect 26136 46003 26208 46079
rect 26256 46003 26328 46079
rect 26010 45885 26082 45961
rect 26136 45885 26208 45961
rect 26256 45885 26328 45961
rect 504 45225 576 45301
rect 626 45225 698 45301
rect 752 45225 824 45301
rect 504 45078 576 45154
rect 626 45078 698 45154
rect 752 45078 824 45154
rect 504 44941 576 45017
rect 626 44941 698 45017
rect 752 44941 824 45017
rect 503 44655 575 44731
rect 629 44655 701 44731
rect 749 44655 821 44731
rect 503 44537 575 44613
rect 629 44537 701 44613
rect 749 44537 821 44613
rect 25068 44499 25140 44575
rect 25194 44499 25266 44575
rect 25314 44499 25386 44575
rect 25068 44381 25140 44457
rect 25194 44381 25266 44457
rect 25314 44381 25386 44457
rect 503 43468 575 43544
rect 629 43468 701 43544
rect 749 43468 821 43544
rect 503 43350 575 43426
rect 629 43350 701 43426
rect 749 43350 821 43426
rect 25068 43364 25140 43440
rect 25194 43364 25266 43440
rect 25314 43364 25386 43440
rect 25068 43246 25140 43322
rect 25194 43246 25266 43322
rect 25314 43246 25386 43322
rect 504 42984 576 43060
rect 626 42984 698 43060
rect 752 42984 824 43060
rect 504 42837 576 42913
rect 626 42837 698 42913
rect 752 42837 824 42913
rect 504 42700 576 42776
rect 626 42700 698 42776
rect 752 42700 824 42776
rect 26010 42082 26082 42158
rect 26136 42082 26208 42158
rect 26256 42082 26328 42158
rect 26010 41964 26082 42040
rect 26136 41964 26208 42040
rect 26256 41964 26328 42040
rect 504 41225 576 41301
rect 626 41225 698 41301
rect 752 41225 824 41301
rect 504 41078 576 41154
rect 626 41078 698 41154
rect 752 41078 824 41154
rect 504 40941 576 41017
rect 626 40941 698 41017
rect 752 40941 824 41017
rect 503 40646 575 40722
rect 629 40646 701 40722
rect 749 40646 821 40722
rect 503 40528 575 40604
rect 629 40528 701 40604
rect 749 40528 821 40604
rect 25068 40605 25140 40681
rect 25194 40605 25266 40681
rect 25314 40605 25386 40681
rect 25068 40487 25140 40563
rect 25194 40487 25266 40563
rect 25314 40487 25386 40563
rect 503 39493 575 39569
rect 629 39493 701 39569
rect 749 39493 821 39569
rect 503 39375 575 39451
rect 629 39375 701 39451
rect 749 39375 821 39451
rect 25068 39452 25140 39528
rect 25194 39452 25266 39528
rect 25314 39452 25386 39528
rect 25068 39334 25140 39410
rect 25194 39334 25266 39410
rect 25314 39334 25386 39410
rect 504 38984 576 39060
rect 626 38984 698 39060
rect 752 38984 824 39060
rect 504 38837 576 38913
rect 626 38837 698 38913
rect 752 38837 824 38913
rect 504 38700 576 38776
rect 626 38700 698 38776
rect 752 38700 824 38776
rect 26010 37824 26082 37900
rect 26136 37824 26208 37900
rect 26256 37824 26328 37900
rect 26010 37706 26082 37782
rect 26136 37706 26208 37782
rect 26256 37706 26328 37782
rect 504 37224 576 37300
rect 626 37224 698 37300
rect 752 37224 824 37300
rect 504 37077 576 37153
rect 626 37077 698 37153
rect 752 37077 824 37153
rect 504 36940 576 37016
rect 626 36940 698 37016
rect 752 36940 824 37016
rect 503 36433 575 36509
rect 629 36433 701 36509
rect 749 36433 821 36509
rect 503 36315 575 36391
rect 629 36315 701 36391
rect 749 36315 821 36391
rect 25068 36336 25140 36412
rect 25194 36336 25266 36412
rect 25314 36336 25386 36412
rect 25068 36218 25140 36294
rect 25194 36218 25266 36294
rect 25314 36218 25386 36294
rect 2257 35869 2313 35925
rect 2337 35869 2393 35925
rect 2257 35789 2313 35845
rect 2337 35789 2393 35845
rect 32 35661 112 35741
rect 157 35661 237 35741
rect 282 35661 362 35741
rect 32 35555 112 35635
rect 157 35555 237 35635
rect 282 35555 362 35635
rect 2016 35315 2072 35319
rect 2016 35263 2020 35315
rect 2020 35263 2072 35315
rect 2098 35316 2154 35320
rect 2098 35264 2150 35316
rect 2150 35264 2154 35316
rect 2017 35235 2073 35239
rect 2017 35183 2021 35235
rect 2021 35183 2073 35235
rect 2099 35236 2155 35240
rect 2099 35184 2151 35236
rect 2151 35184 2155 35236
rect 3361 35848 3417 35904
rect 3441 35848 3497 35904
rect 3361 35768 3417 35824
rect 3441 35768 3497 35824
rect 25535 35646 25615 35726
rect 25660 35646 25740 35726
rect 25785 35646 25865 35726
rect 25534 35526 25614 35606
rect 25659 35526 25739 35606
rect 25784 35526 25864 35606
rect 479 35052 561 35130
rect 593 35052 675 35130
rect 707 35052 789 35130
rect 16 34508 98 34586
rect 130 34508 212 34586
rect 244 34508 326 34586
rect 479 33964 561 34042
rect 593 33964 675 34042
rect 707 33964 789 34042
rect 16 33420 98 33498
rect 130 33420 212 33498
rect 244 33420 326 33498
rect 479 32876 561 32954
rect 593 32876 675 32954
rect 707 32876 789 32954
rect 503 28226 575 28302
rect 629 28226 701 28302
rect 749 28226 821 28302
rect 503 28108 575 28184
rect 629 28108 701 28184
rect 749 28108 821 28184
rect 3360 35262 3416 35318
rect 3440 35261 3496 35317
rect 3361 35181 3417 35237
rect 3441 35181 3497 35237
rect 25061 34892 25141 34972
rect 25186 34892 25266 34972
rect 25311 34892 25391 34972
rect 25060 34772 25140 34852
rect 25185 34772 25265 34852
rect 25310 34772 25390 34852
rect 25069 34316 25141 34392
rect 25191 34316 25263 34392
rect 25317 34316 25389 34392
rect 25069 34169 25141 34245
rect 25191 34169 25263 34245
rect 25317 34169 25389 34245
rect 25069 34032 25141 34108
rect 25191 34032 25263 34108
rect 25317 34032 25389 34108
rect 24560 33396 24640 33476
rect 24685 33396 24765 33476
rect 24810 33396 24890 33476
rect 24559 33276 24639 33356
rect 24684 33276 24764 33356
rect 24809 33276 24889 33356
rect 25535 33396 25615 33476
rect 25660 33396 25740 33476
rect 25785 33396 25865 33476
rect 25534 33276 25614 33356
rect 25659 33276 25739 33356
rect 25784 33276 25864 33356
rect 25069 32556 25141 32632
rect 25191 32556 25263 32632
rect 25317 32556 25389 32632
rect 3144 32401 3200 32463
rect 3224 32401 3280 32463
rect 25069 32409 25141 32485
rect 25191 32409 25263 32485
rect 25317 32409 25389 32485
rect 25069 32272 25141 32348
rect 25191 32272 25263 32348
rect 25317 32272 25389 32348
rect 25060 31837 25140 31917
rect 25185 31837 25265 31917
rect 25310 31837 25390 31917
rect 25059 31717 25139 31797
rect 25184 31717 25264 31797
rect 25309 31717 25389 31797
rect 25068 28226 25140 28302
rect 25194 28226 25266 28302
rect 25314 28226 25386 28302
rect 25068 28108 25140 28184
rect 25194 28108 25266 28184
rect 25314 28108 25386 28184
rect 503 27444 575 27520
rect 629 27444 701 27520
rect 749 27444 821 27520
rect 503 27326 575 27402
rect 629 27326 701 27402
rect 749 27326 821 27402
rect 25068 27444 25140 27520
rect 25194 27444 25266 27520
rect 25314 27444 25386 27520
rect 25068 27326 25140 27402
rect 25194 27326 25266 27402
rect 25314 27326 25386 27402
rect 504 26985 576 27061
rect 626 26985 698 27061
rect 752 26985 824 27061
rect 504 26838 576 26914
rect 626 26838 698 26914
rect 752 26838 824 26914
rect 504 26701 576 26777
rect 626 26701 698 26777
rect 752 26701 824 26777
rect 26010 26054 26082 26130
rect 26136 26054 26208 26130
rect 26256 26054 26328 26130
rect 26010 25936 26082 26012
rect 26136 25936 26208 26012
rect 26256 25936 26328 26012
rect 504 25218 576 25294
rect 626 25218 698 25294
rect 752 25218 824 25294
rect 504 25071 576 25147
rect 626 25071 698 25147
rect 752 25071 824 25147
rect 504 24934 576 25010
rect 626 24934 698 25010
rect 752 24934 824 25010
rect 503 24532 575 24608
rect 629 24532 701 24608
rect 749 24532 821 24608
rect 503 24414 575 24490
rect 629 24414 701 24490
rect 749 24414 821 24490
rect 25068 24483 25140 24559
rect 25194 24483 25266 24559
rect 25314 24483 25386 24559
rect 25068 24365 25140 24441
rect 25194 24365 25266 24441
rect 25314 24365 25386 24441
rect 503 23528 575 23604
rect 629 23528 701 23604
rect 749 23528 821 23604
rect 503 23410 575 23486
rect 629 23410 701 23486
rect 749 23410 821 23486
rect 25068 23366 25140 23442
rect 25194 23366 25266 23442
rect 25314 23366 25386 23442
rect 25068 23248 25140 23324
rect 25194 23248 25266 23324
rect 25314 23248 25386 23324
rect 504 22984 576 23060
rect 626 22984 698 23060
rect 752 22984 824 23060
rect 504 22837 576 22913
rect 626 22837 698 22913
rect 752 22837 824 22913
rect 504 22700 576 22776
rect 626 22700 698 22776
rect 752 22700 824 22776
rect 26010 21895 26082 21971
rect 26136 21895 26208 21971
rect 26256 21895 26328 21971
rect 26010 21777 26082 21853
rect 26136 21777 26208 21853
rect 26256 21777 26328 21853
rect 504 21224 576 21300
rect 626 21224 698 21300
rect 752 21224 824 21300
rect 504 21077 576 21153
rect 626 21077 698 21153
rect 752 21077 824 21153
rect 504 20940 576 21016
rect 626 20940 698 21016
rect 752 20940 824 21016
rect 503 20550 575 20626
rect 629 20550 701 20626
rect 749 20550 821 20626
rect 503 20432 575 20508
rect 629 20432 701 20508
rect 749 20432 821 20508
rect 25068 20523 25140 20599
rect 25194 20523 25266 20599
rect 25314 20523 25386 20599
rect 25068 20405 25140 20481
rect 25194 20405 25266 20481
rect 25314 20405 25386 20481
rect 503 19468 575 19544
rect 629 19468 701 19544
rect 749 19468 821 19544
rect 503 19350 575 19426
rect 629 19350 701 19426
rect 749 19350 821 19426
rect 25068 19348 25140 19424
rect 25194 19348 25266 19424
rect 25314 19348 25386 19424
rect 25068 19230 25140 19306
rect 25194 19230 25266 19306
rect 25314 19230 25386 19306
rect 504 18984 576 19060
rect 626 18984 698 19060
rect 752 18984 824 19060
rect 504 18837 576 18913
rect 626 18837 698 18913
rect 752 18837 824 18913
rect 504 18700 576 18776
rect 626 18700 698 18776
rect 752 18700 824 18776
rect 26010 18105 26082 18181
rect 26136 18105 26208 18181
rect 26256 18105 26328 18181
rect 26010 17987 26082 18063
rect 26136 17987 26208 18063
rect 26256 17987 26328 18063
rect 504 17225 576 17301
rect 626 17225 698 17301
rect 752 17225 824 17301
rect 504 17078 576 17154
rect 626 17078 698 17154
rect 752 17078 824 17154
rect 504 16941 576 17017
rect 626 16941 698 17017
rect 752 16941 824 17017
rect 503 16593 575 16669
rect 629 16593 701 16669
rect 749 16593 821 16669
rect 503 16475 575 16551
rect 629 16475 701 16551
rect 749 16475 821 16551
rect 25068 16507 25140 16583
rect 25194 16507 25266 16583
rect 25314 16507 25386 16583
rect 25068 16389 25140 16465
rect 25194 16389 25266 16465
rect 25314 16389 25386 16465
rect 503 15492 575 15568
rect 629 15492 701 15568
rect 749 15492 821 15568
rect 503 15374 575 15450
rect 629 15374 701 15450
rect 749 15374 821 15450
rect 25068 15336 25140 15412
rect 25194 15336 25266 15412
rect 25314 15336 25386 15412
rect 25068 15218 25140 15294
rect 25194 15218 25266 15294
rect 25314 15218 25386 15294
rect 504 14984 576 15060
rect 626 14984 698 15060
rect 752 14984 824 15060
rect 504 14837 576 14913
rect 626 14837 698 14913
rect 752 14837 824 14913
rect 504 14700 576 14776
rect 626 14700 698 14776
rect 752 14700 824 14776
rect 26010 13998 26082 14074
rect 26136 13998 26208 14074
rect 26256 13998 26328 14074
rect 26010 13880 26082 13956
rect 26136 13880 26208 13956
rect 26256 13880 26328 13956
rect 504 13224 576 13300
rect 626 13224 698 13300
rect 752 13224 824 13300
rect 504 13077 576 13153
rect 626 13077 698 13153
rect 752 13077 824 13153
rect 504 12940 576 13016
rect 626 12940 698 13016
rect 752 12940 824 13016
rect 503 12626 575 12702
rect 629 12626 701 12702
rect 749 12626 821 12702
rect 503 12508 575 12584
rect 629 12508 701 12584
rect 749 12508 821 12584
rect 25068 12575 25140 12651
rect 25194 12575 25266 12651
rect 25314 12575 25386 12651
rect 25068 12457 25140 12533
rect 25194 12457 25266 12533
rect 25314 12457 25386 12533
rect 503 11410 575 11486
rect 629 11410 701 11486
rect 749 11410 821 11486
rect 503 11292 575 11368
rect 629 11292 701 11368
rect 749 11292 821 11368
rect 25068 11361 25140 11437
rect 25194 11361 25266 11437
rect 25314 11361 25386 11437
rect 25068 11243 25140 11319
rect 25194 11243 25266 11319
rect 25314 11243 25386 11319
rect 504 10984 576 11060
rect 626 10984 698 11060
rect 752 10984 824 11060
rect 504 10837 576 10913
rect 626 10837 698 10913
rect 752 10837 824 10913
rect 504 10700 576 10776
rect 626 10700 698 10776
rect 752 10700 824 10776
rect 26010 10180 26082 10256
rect 26136 10180 26208 10256
rect 26256 10180 26328 10256
rect 26010 10062 26082 10138
rect 26136 10062 26208 10138
rect 26256 10062 26328 10138
rect 504 9224 576 9300
rect 626 9224 698 9300
rect 752 9224 824 9300
rect 504 9077 576 9153
rect 626 9077 698 9153
rect 752 9077 824 9153
rect 504 8940 576 9016
rect 626 8940 698 9016
rect 752 8940 824 9016
rect 503 8545 575 8621
rect 629 8545 701 8621
rect 749 8545 821 8621
rect 503 8427 575 8503
rect 629 8427 701 8503
rect 749 8427 821 8503
rect 25068 8518 25140 8594
rect 25194 8518 25266 8594
rect 25314 8518 25386 8594
rect 25068 8400 25140 8476
rect 25194 8400 25266 8476
rect 25314 8400 25386 8476
rect 503 7423 575 7499
rect 629 7423 701 7499
rect 749 7423 821 7499
rect 503 7305 575 7381
rect 629 7305 701 7381
rect 749 7305 821 7381
rect 25068 7361 25140 7437
rect 25194 7361 25266 7437
rect 25314 7361 25386 7437
rect 25068 7243 25140 7319
rect 25194 7243 25266 7319
rect 25314 7243 25386 7319
rect 504 6985 576 7061
rect 626 6985 698 7061
rect 752 6985 824 7061
rect 504 6838 576 6914
rect 626 6838 698 6914
rect 752 6838 824 6914
rect 504 6701 576 6777
rect 626 6701 698 6777
rect 752 6701 824 6777
rect 26010 6216 26082 6292
rect 26136 6216 26208 6292
rect 26256 6216 26328 6292
rect 26010 6098 26082 6174
rect 26136 6098 26208 6174
rect 26256 6098 26328 6174
rect 504 5223 576 5299
rect 626 5223 698 5299
rect 752 5223 824 5299
rect 504 5076 576 5152
rect 626 5076 698 5152
rect 752 5076 824 5152
rect 504 4939 576 5015
rect 626 4939 698 5015
rect 752 4939 824 5015
rect 503 4563 575 4639
rect 629 4563 701 4639
rect 749 4563 821 4639
rect 503 4445 575 4521
rect 629 4445 701 4521
rect 749 4445 821 4521
rect 25068 4518 25140 4594
rect 25194 4518 25266 4594
rect 25314 4518 25386 4594
rect 25068 4400 25140 4476
rect 25194 4400 25266 4476
rect 25314 4400 25386 4476
rect 503 3452 575 3528
rect 629 3452 701 3528
rect 749 3452 821 3528
rect 503 3334 575 3410
rect 629 3334 701 3410
rect 749 3334 821 3410
rect 25068 3361 25140 3437
rect 25194 3361 25266 3437
rect 25314 3361 25386 3437
rect 25068 3243 25140 3319
rect 25194 3243 25266 3319
rect 25314 3243 25386 3319
rect 504 2985 576 3061
rect 626 2985 698 3061
rect 752 2985 824 3061
rect 504 2838 576 2914
rect 626 2838 698 2914
rect 752 2838 824 2914
rect 504 2701 576 2777
rect 626 2701 698 2777
rect 752 2701 824 2777
rect 26010 2204 26082 2280
rect 26136 2204 26208 2280
rect 26256 2204 26328 2280
rect 26010 2086 26082 2162
rect 26136 2086 26208 2162
rect 26256 2086 26328 2162
rect 504 1224 576 1300
rect 626 1224 698 1300
rect 752 1224 824 1300
rect 504 1077 576 1153
rect 626 1077 698 1153
rect 752 1077 824 1153
rect 504 940 576 1016
rect 626 940 698 1016
rect 752 940 824 1016
rect 503 629 575 705
rect 629 629 701 705
rect 749 629 821 705
rect 503 511 575 587
rect 629 511 701 587
rect 749 511 821 587
rect 25068 518 25140 594
rect 25194 518 25266 594
rect 25314 518 25386 594
rect 25068 400 25140 476
rect 25194 400 25266 476
rect 25314 400 25386 476
<< metal3 >>
rect 25026 63492 25426 63517
rect 463 63452 864 63477
rect 463 63376 503 63452
rect 575 63376 629 63452
rect 701 63376 749 63452
rect 821 63376 864 63452
rect 463 63334 864 63376
rect 463 63258 503 63334
rect 575 63258 629 63334
rect 701 63258 749 63334
rect 821 63258 864 63334
rect 25026 63416 25068 63492
rect 25140 63416 25194 63492
rect 25266 63416 25314 63492
rect 25386 63416 25426 63492
rect 25026 63374 25426 63416
rect 25026 63298 25068 63374
rect 25140 63298 25194 63374
rect 25266 63298 25314 63374
rect 25386 63298 25426 63374
rect 25026 63262 25426 63298
rect 463 63222 864 63258
rect 463 63060 863 63109
rect 463 62984 504 63060
rect 576 62984 626 63060
rect 698 62984 752 63060
rect 824 62984 863 63060
rect 463 62913 863 62984
rect 463 62837 504 62913
rect 576 62837 626 62913
rect 698 62837 752 62913
rect 824 62837 863 62913
rect 463 62776 863 62837
rect 463 62700 504 62776
rect 576 62700 626 62776
rect 698 62700 752 62776
rect 824 62700 863 62776
rect 463 62650 863 62700
rect 25970 62071 26370 62096
rect 25970 61995 26010 62071
rect 26082 61995 26136 62071
rect 26208 61995 26256 62071
rect 26328 61995 26370 62071
rect 25970 61953 26370 61995
rect 25970 61877 26010 61953
rect 26082 61877 26136 61953
rect 26208 61877 26256 61953
rect 26328 61877 26370 61953
rect 25970 61841 26370 61877
rect 463 61300 863 61349
rect 463 61224 504 61300
rect 576 61224 626 61300
rect 698 61224 752 61300
rect 824 61224 863 61300
rect 463 61153 863 61224
rect 463 61077 504 61153
rect 576 61077 626 61153
rect 698 61077 752 61153
rect 824 61077 863 61153
rect 463 61016 863 61077
rect 463 60940 504 61016
rect 576 60940 626 61016
rect 698 60940 752 61016
rect 824 60940 863 61016
rect 463 60890 863 60940
rect 463 60779 864 60804
rect 463 60703 503 60779
rect 575 60703 629 60779
rect 701 60703 749 60779
rect 821 60703 864 60779
rect 463 60661 864 60703
rect 463 60585 503 60661
rect 575 60585 629 60661
rect 701 60585 749 60661
rect 821 60585 864 60661
rect 463 60549 864 60585
rect 25028 60695 25428 60720
rect 25028 60619 25068 60695
rect 25140 60619 25194 60695
rect 25266 60619 25314 60695
rect 25386 60619 25428 60695
rect 25028 60577 25428 60619
rect 25028 60501 25068 60577
rect 25140 60501 25194 60577
rect 25266 60501 25314 60577
rect 25386 60501 25428 60577
rect 25028 60465 25428 60501
rect 25026 59492 25426 59517
rect 463 59450 864 59475
rect 463 59374 503 59450
rect 575 59374 629 59450
rect 701 59374 749 59450
rect 821 59374 864 59450
rect 463 59332 864 59374
rect 463 59256 503 59332
rect 575 59256 629 59332
rect 701 59256 749 59332
rect 821 59256 864 59332
rect 25026 59416 25068 59492
rect 25140 59416 25194 59492
rect 25266 59416 25314 59492
rect 25386 59416 25426 59492
rect 25026 59374 25426 59416
rect 25026 59298 25068 59374
rect 25140 59298 25194 59374
rect 25266 59298 25314 59374
rect 25386 59298 25426 59374
rect 25026 59262 25426 59298
rect 463 59220 864 59256
rect 463 59060 863 59109
rect 463 58984 504 59060
rect 576 58984 626 59060
rect 698 58984 752 59060
rect 824 58984 863 59060
rect 463 58913 863 58984
rect 463 58837 504 58913
rect 576 58837 626 58913
rect 698 58837 752 58913
rect 824 58837 863 58913
rect 463 58776 863 58837
rect 463 58700 504 58776
rect 576 58700 626 58776
rect 698 58700 752 58776
rect 824 58700 863 58776
rect 463 58650 863 58700
rect 25970 58058 26370 58083
rect 25970 57982 26010 58058
rect 26082 57982 26136 58058
rect 26208 57982 26256 58058
rect 26328 57982 26370 58058
rect 25970 57940 26370 57982
rect 25970 57864 26010 57940
rect 26082 57864 26136 57940
rect 26208 57864 26256 57940
rect 26328 57864 26370 57940
rect 25970 57828 26370 57864
rect 463 57301 863 57350
rect 463 57225 504 57301
rect 576 57225 626 57301
rect 698 57225 752 57301
rect 824 57225 863 57301
rect 463 57154 863 57225
rect 463 57078 504 57154
rect 576 57078 626 57154
rect 698 57078 752 57154
rect 824 57078 863 57154
rect 463 57017 863 57078
rect 463 56941 504 57017
rect 576 56941 626 57017
rect 698 56941 752 57017
rect 824 56941 863 57017
rect 463 56891 863 56941
rect 463 56710 864 56735
rect 463 56634 503 56710
rect 575 56634 629 56710
rect 701 56634 749 56710
rect 821 56634 864 56710
rect 463 56592 864 56634
rect 463 56516 503 56592
rect 575 56516 629 56592
rect 701 56516 749 56592
rect 821 56516 864 56592
rect 463 56480 864 56516
rect 25028 56695 25428 56720
rect 25028 56619 25068 56695
rect 25140 56619 25194 56695
rect 25266 56619 25314 56695
rect 25386 56619 25428 56695
rect 25028 56577 25428 56619
rect 25028 56501 25068 56577
rect 25140 56501 25194 56577
rect 25266 56501 25314 56577
rect 25386 56501 25428 56577
rect 25028 56465 25428 56501
rect 463 55532 864 55557
rect 463 55456 503 55532
rect 575 55456 629 55532
rect 701 55456 749 55532
rect 821 55456 864 55532
rect 463 55414 864 55456
rect 463 55338 503 55414
rect 575 55338 629 55414
rect 701 55338 749 55414
rect 821 55338 864 55414
rect 463 55302 864 55338
rect 25026 55492 25426 55517
rect 25026 55416 25068 55492
rect 25140 55416 25194 55492
rect 25266 55416 25314 55492
rect 25386 55416 25426 55492
rect 25026 55374 25426 55416
rect 25026 55298 25068 55374
rect 25140 55298 25194 55374
rect 25266 55298 25314 55374
rect 25386 55298 25426 55374
rect 25026 55262 25426 55298
rect 464 55068 864 55109
rect 463 55060 864 55068
rect 463 54984 504 55060
rect 576 54984 626 55060
rect 698 54984 752 55060
rect 824 54984 864 55060
rect 463 54913 864 54984
rect 463 54837 504 54913
rect 576 54837 626 54913
rect 698 54837 752 54913
rect 824 54837 864 54913
rect 463 54776 864 54837
rect 463 54700 504 54776
rect 576 54700 626 54776
rect 698 54700 752 54776
rect 824 54700 864 54776
rect 463 54650 864 54700
rect 25970 54057 26370 54082
rect 25970 53981 26010 54057
rect 26082 53981 26136 54057
rect 26208 53981 26256 54057
rect 26328 53981 26370 54057
rect 25970 53939 26370 53981
rect 25970 53863 26010 53939
rect 26082 53863 26136 53939
rect 26208 53863 26256 53939
rect 26328 53863 26370 53939
rect 25970 53827 26370 53863
rect 463 53301 863 53350
rect 463 53225 504 53301
rect 576 53225 626 53301
rect 698 53225 752 53301
rect 824 53225 863 53301
rect 463 53154 863 53225
rect 463 53078 504 53154
rect 576 53078 626 53154
rect 698 53078 752 53154
rect 824 53078 863 53154
rect 463 53017 863 53078
rect 463 52941 504 53017
rect 576 52941 626 53017
rect 698 52941 752 53017
rect 824 52941 863 53017
rect 463 52891 863 52941
rect 463 52684 866 52709
rect 463 52608 503 52684
rect 575 52608 629 52684
rect 701 52608 749 52684
rect 821 52608 866 52684
rect 463 52566 866 52608
rect 463 52490 503 52566
rect 575 52490 629 52566
rect 701 52490 749 52566
rect 821 52490 866 52566
rect 463 52454 866 52490
rect 25028 52695 25428 52720
rect 25028 52619 25068 52695
rect 25140 52619 25194 52695
rect 25266 52619 25314 52695
rect 25386 52619 25428 52695
rect 25028 52577 25428 52619
rect 25028 52501 25068 52577
rect 25140 52501 25194 52577
rect 25266 52501 25314 52577
rect 25386 52501 25428 52577
rect 25028 52465 25428 52501
rect 25027 51546 25427 51571
rect 463 51481 864 51506
rect 463 51405 503 51481
rect 575 51405 629 51481
rect 701 51405 749 51481
rect 821 51405 864 51481
rect 463 51363 864 51405
rect 463 51287 503 51363
rect 575 51287 629 51363
rect 701 51287 749 51363
rect 821 51287 864 51363
rect 25027 51470 25068 51546
rect 25140 51470 25194 51546
rect 25266 51470 25314 51546
rect 25386 51470 25427 51546
rect 25027 51428 25427 51470
rect 25027 51352 25068 51428
rect 25140 51352 25194 51428
rect 25266 51352 25314 51428
rect 25386 51352 25427 51428
rect 25027 51316 25427 51352
rect 463 51251 864 51287
rect 464 51068 864 51109
rect 463 51060 864 51068
rect 463 50984 504 51060
rect 576 50984 626 51060
rect 698 50984 752 51060
rect 824 50984 864 51060
rect 463 50913 864 50984
rect 463 50837 504 50913
rect 576 50837 626 50913
rect 698 50837 752 50913
rect 824 50837 864 50913
rect 463 50776 864 50837
rect 463 50700 504 50776
rect 576 50700 626 50776
rect 698 50700 752 50776
rect 824 50700 864 50776
rect 463 50650 864 50700
rect 25970 50096 26370 50121
rect 25970 50020 26010 50096
rect 26082 50020 26136 50096
rect 26208 50020 26256 50096
rect 26328 50020 26370 50096
rect 25970 49978 26370 50020
rect 25970 49902 26010 49978
rect 26082 49902 26136 49978
rect 26208 49902 26256 49978
rect 26328 49902 26370 49978
rect 25970 49866 26370 49902
rect 463 49299 863 49348
rect 463 49223 504 49299
rect 576 49223 626 49299
rect 698 49223 752 49299
rect 824 49223 863 49299
rect 463 49152 863 49223
rect 463 49076 504 49152
rect 576 49076 626 49152
rect 698 49076 752 49152
rect 824 49076 863 49152
rect 463 49015 863 49076
rect 463 48939 504 49015
rect 576 48939 626 49015
rect 698 48939 752 49015
rect 824 48939 863 49015
rect 463 48889 863 48939
rect 463 48704 864 48729
rect 463 48628 503 48704
rect 575 48628 629 48704
rect 701 48628 749 48704
rect 821 48628 864 48704
rect 463 48586 864 48628
rect 463 48510 503 48586
rect 575 48510 629 48586
rect 701 48510 749 48586
rect 821 48510 864 48586
rect 463 48474 864 48510
rect 25028 48630 25428 48655
rect 25028 48554 25068 48630
rect 25140 48554 25194 48630
rect 25266 48554 25314 48630
rect 25386 48554 25428 48630
rect 25028 48512 25428 48554
rect 25028 48436 25068 48512
rect 25140 48436 25194 48512
rect 25266 48436 25314 48512
rect 25386 48436 25428 48512
rect 25028 48400 25428 48436
rect 463 47497 866 47522
rect 463 47421 503 47497
rect 575 47421 629 47497
rect 701 47421 749 47497
rect 821 47421 866 47497
rect 463 47379 866 47421
rect 463 47303 503 47379
rect 575 47303 629 47379
rect 701 47303 749 47379
rect 821 47303 866 47379
rect 463 47267 866 47303
rect 25027 47447 25427 47472
rect 25027 47371 25068 47447
rect 25140 47371 25194 47447
rect 25266 47371 25314 47447
rect 25386 47371 25427 47447
rect 25027 47329 25427 47371
rect 25027 47253 25068 47329
rect 25140 47253 25194 47329
rect 25266 47253 25314 47329
rect 25386 47253 25427 47329
rect 25027 47217 25427 47253
rect 463 47060 863 47109
rect 463 46984 504 47060
rect 576 46984 626 47060
rect 698 46984 752 47060
rect 824 46984 863 47060
rect 463 46913 863 46984
rect 463 46837 504 46913
rect 576 46837 626 46913
rect 698 46837 752 46913
rect 824 46837 863 46913
rect 463 46776 863 46837
rect 463 46700 504 46776
rect 576 46700 626 46776
rect 698 46700 752 46776
rect 824 46700 863 46776
rect 463 46650 863 46700
rect 25970 46079 26370 46104
rect 25970 46003 26010 46079
rect 26082 46003 26136 46079
rect 26208 46003 26256 46079
rect 26328 46003 26370 46079
rect 25970 45961 26370 46003
rect 25970 45885 26010 45961
rect 26082 45885 26136 45961
rect 26208 45885 26256 45961
rect 26328 45885 26370 45961
rect 25970 45849 26370 45885
rect 463 45301 863 45350
rect 463 45225 504 45301
rect 576 45225 626 45301
rect 698 45225 752 45301
rect 824 45225 863 45301
rect 463 45154 863 45225
rect 463 45078 504 45154
rect 576 45078 626 45154
rect 698 45078 752 45154
rect 824 45078 863 45154
rect 463 45017 863 45078
rect 463 44941 504 45017
rect 576 44941 626 45017
rect 698 44941 752 45017
rect 824 44941 863 45017
rect 463 44891 863 44941
rect 463 44731 864 44756
rect 463 44655 503 44731
rect 575 44655 629 44731
rect 701 44655 749 44731
rect 821 44655 864 44731
rect 463 44613 864 44655
rect 463 44537 503 44613
rect 575 44537 629 44613
rect 701 44537 749 44613
rect 821 44537 864 44613
rect 463 44501 864 44537
rect 25028 44575 25428 44600
rect 25028 44499 25068 44575
rect 25140 44499 25194 44575
rect 25266 44499 25314 44575
rect 25386 44499 25428 44575
rect 25028 44457 25428 44499
rect 25028 44381 25068 44457
rect 25140 44381 25194 44457
rect 25266 44381 25314 44457
rect 25386 44381 25428 44457
rect 25028 44345 25428 44381
rect 463 43544 864 43569
rect 463 43468 503 43544
rect 575 43468 629 43544
rect 701 43468 749 43544
rect 821 43468 864 43544
rect 463 43426 864 43468
rect 463 43350 503 43426
rect 575 43350 629 43426
rect 701 43350 749 43426
rect 821 43350 864 43426
rect 463 43314 864 43350
rect 25028 43440 25428 43465
rect 25028 43364 25068 43440
rect 25140 43364 25194 43440
rect 25266 43364 25314 43440
rect 25386 43364 25428 43440
rect 25028 43322 25428 43364
rect 25028 43246 25068 43322
rect 25140 43246 25194 43322
rect 25266 43246 25314 43322
rect 25386 43246 25428 43322
rect 25028 43210 25428 43246
rect 463 43060 863 43109
rect 463 42984 504 43060
rect 576 42984 626 43060
rect 698 42984 752 43060
rect 824 42984 863 43060
rect 463 42913 863 42984
rect 463 42837 504 42913
rect 576 42837 626 42913
rect 698 42837 752 42913
rect 824 42837 863 42913
rect 463 42776 863 42837
rect 463 42700 504 42776
rect 576 42700 626 42776
rect 698 42700 752 42776
rect 824 42700 863 42776
rect 463 42650 863 42700
rect 25970 42158 26370 42183
rect 25970 42082 26010 42158
rect 26082 42082 26136 42158
rect 26208 42082 26256 42158
rect 26328 42082 26370 42158
rect 25970 42040 26370 42082
rect 25970 41964 26010 42040
rect 26082 41964 26136 42040
rect 26208 41964 26256 42040
rect 26328 41964 26370 42040
rect 25970 41928 26370 41964
rect 463 41301 863 41350
rect 463 41225 504 41301
rect 576 41225 626 41301
rect 698 41225 752 41301
rect 824 41225 863 41301
rect 463 41154 863 41225
rect 463 41078 504 41154
rect 576 41078 626 41154
rect 698 41078 752 41154
rect 824 41078 863 41154
rect 463 41017 863 41078
rect 463 40941 504 41017
rect 576 40941 626 41017
rect 698 40941 752 41017
rect 824 40941 863 41017
rect 463 40891 863 40941
rect 463 40722 864 40747
rect 463 40646 503 40722
rect 575 40646 629 40722
rect 701 40646 749 40722
rect 821 40646 864 40722
rect 463 40604 864 40646
rect 463 40528 503 40604
rect 575 40528 629 40604
rect 701 40528 749 40604
rect 821 40528 864 40604
rect 463 40492 864 40528
rect 25028 40681 25428 40706
rect 25028 40605 25068 40681
rect 25140 40605 25194 40681
rect 25266 40605 25314 40681
rect 25386 40605 25428 40681
rect 25028 40563 25428 40605
rect 25028 40487 25068 40563
rect 25140 40487 25194 40563
rect 25266 40487 25314 40563
rect 25386 40487 25428 40563
rect 25028 40451 25428 40487
rect 463 39569 864 39594
rect 463 39493 503 39569
rect 575 39493 629 39569
rect 701 39493 749 39569
rect 821 39493 864 39569
rect 463 39451 864 39493
rect 463 39375 503 39451
rect 575 39375 629 39451
rect 701 39375 749 39451
rect 821 39375 864 39451
rect 463 39339 864 39375
rect 25028 39528 25428 39553
rect 25028 39452 25068 39528
rect 25140 39452 25194 39528
rect 25266 39452 25314 39528
rect 25386 39452 25428 39528
rect 25028 39410 25428 39452
rect 25028 39334 25068 39410
rect 25140 39334 25194 39410
rect 25266 39334 25314 39410
rect 25386 39334 25428 39410
rect 25028 39298 25428 39334
rect 463 39060 863 39109
rect 463 38984 504 39060
rect 576 38984 626 39060
rect 698 38984 752 39060
rect 824 38984 863 39060
rect 463 38913 863 38984
rect 463 38837 504 38913
rect 576 38837 626 38913
rect 698 38837 752 38913
rect 824 38837 863 38913
rect 463 38776 863 38837
rect 463 38700 504 38776
rect 576 38700 626 38776
rect 698 38700 752 38776
rect 824 38700 863 38776
rect 463 38650 863 38700
rect 25970 37900 26370 37925
rect 25970 37824 26010 37900
rect 26082 37824 26136 37900
rect 26208 37824 26256 37900
rect 26328 37824 26370 37900
rect 25970 37782 26370 37824
rect 25970 37706 26010 37782
rect 26082 37706 26136 37782
rect 26208 37706 26256 37782
rect 26328 37706 26370 37782
rect 25970 37670 26370 37706
rect 463 37300 863 37350
rect 463 37224 504 37300
rect 576 37224 626 37300
rect 698 37224 752 37300
rect 824 37224 863 37300
rect 463 37153 863 37224
rect 463 37077 504 37153
rect 576 37077 626 37153
rect 698 37077 752 37153
rect 824 37077 863 37153
rect 463 37016 863 37077
rect 463 36940 504 37016
rect 576 36940 626 37016
rect 698 36940 752 37016
rect 824 36940 863 37016
rect 463 36891 863 36940
rect 463 36890 836 36891
rect 463 36509 863 36534
rect 463 36433 503 36509
rect 575 36433 629 36509
rect 701 36433 749 36509
rect 821 36433 863 36509
rect 463 36391 863 36433
rect 463 36315 503 36391
rect 575 36315 629 36391
rect 701 36315 749 36391
rect 821 36315 863 36391
rect 463 36279 863 36315
rect 25028 36412 25428 36437
rect 25028 36336 25068 36412
rect 25140 36336 25194 36412
rect 25266 36336 25314 36412
rect 25386 36336 25428 36412
rect 25028 36294 25428 36336
rect 25028 36218 25068 36294
rect 25140 36218 25194 36294
rect 25266 36218 25314 36294
rect 25386 36218 25428 36294
rect 25028 36182 25428 36218
rect 2248 35925 2401 35940
rect 2248 35861 2249 35925
rect 2313 35861 2337 35925
rect 2248 35845 2401 35861
rect 2248 35781 2249 35845
rect 2313 35781 2337 35845
rect 2248 35775 2401 35781
rect 3352 35905 4345 35920
rect 3352 35904 4192 35905
rect 3352 35848 3361 35904
rect 3417 35848 3441 35904
rect 3497 35848 4192 35904
rect 3352 35841 4192 35848
rect 4256 35841 4280 35905
rect 4344 35841 4345 35905
rect 3352 35825 4345 35841
rect 3352 35824 4192 35825
rect 3352 35768 3361 35824
rect 3417 35768 3441 35824
rect 3497 35768 4192 35824
rect 3352 35761 4192 35768
rect 4256 35761 4280 35825
rect 4344 35761 4345 35825
rect 3352 35754 4345 35761
rect 0 35741 400 35752
rect 0 35661 32 35741
rect 112 35661 156 35741
rect 237 35661 282 35741
rect 362 35661 400 35741
rect 0 35635 400 35661
rect 0 35555 32 35635
rect 112 35555 156 35635
rect 237 35555 282 35635
rect 362 35555 400 35635
rect 0 35528 400 35555
rect 25502 35726 25902 35752
rect 25502 35646 25535 35726
rect 25615 35646 25660 35726
rect 25740 35646 25785 35726
rect 25865 35646 25902 35726
rect 25502 35606 25902 35646
rect 25502 35526 25534 35606
rect 25614 35526 25659 35606
rect 25739 35526 25784 35606
rect 25864 35526 25902 35606
rect 25502 35497 25902 35526
rect 2011 35320 3502 35333
rect 2011 35319 2098 35320
rect 2011 35263 2016 35319
rect 2072 35264 2098 35319
rect 2154 35318 3502 35320
rect 2154 35264 3360 35318
rect 2072 35263 3360 35264
rect 2011 35262 3360 35263
rect 3416 35317 3502 35318
rect 3416 35262 3440 35317
rect 2011 35261 3440 35262
rect 3496 35261 3502 35317
rect 2011 35240 3502 35261
rect 2011 35239 2099 35240
rect 2011 35183 2017 35239
rect 2073 35184 2099 35239
rect 2155 35237 3502 35240
rect 2155 35184 3361 35237
rect 2073 35183 3361 35184
rect 2011 35181 3361 35183
rect 3417 35181 3441 35237
rect 3497 35181 3502 35237
rect 2011 35169 3502 35181
rect 463 35131 805 35139
rect 463 35051 478 35131
rect 562 35051 592 35131
rect 676 35051 706 35131
rect 790 35051 805 35131
rect 463 35043 805 35051
rect 25028 34972 25428 34998
rect 25028 34892 25061 34972
rect 25141 34892 25186 34972
rect 25266 34892 25311 34972
rect 25391 34892 25428 34972
rect 25028 34852 25428 34892
rect 25028 34772 25060 34852
rect 25140 34772 25185 34852
rect 25265 34772 25310 34852
rect 25390 34772 25428 34852
rect 25028 34743 25428 34772
rect 0 34587 342 34595
rect 0 34507 15 34587
rect 99 34507 129 34587
rect 213 34507 243 34587
rect 327 34507 342 34587
rect 0 34499 342 34507
rect 25028 34392 25428 34442
rect 25028 34316 25069 34392
rect 25141 34316 25191 34392
rect 25263 34316 25317 34392
rect 25389 34316 25428 34392
rect 25028 34245 25428 34316
rect 25028 34169 25069 34245
rect 25141 34169 25191 34245
rect 25263 34169 25317 34245
rect 25389 34169 25428 34245
rect 25028 34108 25428 34169
rect 463 34043 805 34051
rect 463 33963 478 34043
rect 562 33963 592 34043
rect 676 33963 706 34043
rect 790 33963 805 34043
rect 25028 34032 25069 34108
rect 25141 34032 25191 34108
rect 25263 34032 25317 34108
rect 25389 34032 25428 34108
rect 25028 33983 25428 34032
rect 25028 33982 25401 33983
rect 463 33955 805 33963
rect 0 33499 342 33507
rect 0 33419 15 33499
rect 99 33419 129 33499
rect 213 33419 243 33499
rect 327 33419 342 33499
rect 0 33411 342 33419
rect 24527 33476 24927 33502
rect 24527 33396 24560 33476
rect 24640 33396 24685 33476
rect 24765 33396 24810 33476
rect 24890 33396 24927 33476
rect 24527 33356 24927 33396
rect 24527 33276 24559 33356
rect 24639 33276 24684 33356
rect 24764 33276 24809 33356
rect 24889 33276 24927 33356
rect 24527 33247 24927 33276
rect 25502 33476 25902 33502
rect 25502 33396 25535 33476
rect 25615 33396 25660 33476
rect 25740 33396 25785 33476
rect 25865 33396 25902 33476
rect 25502 33356 25902 33396
rect 25502 33276 25534 33356
rect 25614 33276 25659 33356
rect 25739 33276 25784 33356
rect 25864 33276 25902 33356
rect 25502 33247 25902 33276
rect 463 32955 805 32963
rect 463 32875 478 32955
rect 562 32875 592 32955
rect 676 32875 706 32955
rect 790 32875 805 32955
rect 463 32867 805 32875
rect 25028 32632 25428 32682
rect 25028 32556 25069 32632
rect 25141 32556 25191 32632
rect 25263 32556 25317 32632
rect 25389 32556 25428 32632
rect 25028 32485 25428 32556
rect 3135 32475 3288 32476
rect 3135 32463 3289 32475
rect 3135 32399 3136 32463
rect 3200 32399 3224 32463
rect 3288 32399 3289 32463
rect 3135 32391 3289 32399
rect 25028 32409 25069 32485
rect 25141 32409 25191 32485
rect 25263 32409 25317 32485
rect 25389 32409 25428 32485
rect 25028 32348 25428 32409
rect 25028 32272 25069 32348
rect 25141 32272 25191 32348
rect 25263 32272 25317 32348
rect 25389 32272 25428 32348
rect 25028 32223 25428 32272
rect 25028 32222 25401 32223
rect 25027 31917 25427 31943
rect 25027 31837 25060 31917
rect 25140 31837 25185 31917
rect 25265 31837 25310 31917
rect 25390 31837 25427 31917
rect 25027 31797 25427 31837
rect 25027 31717 25059 31797
rect 25139 31717 25184 31797
rect 25264 31717 25309 31797
rect 25389 31717 25427 31797
rect 25027 31688 25427 31717
rect 463 28302 866 28360
rect 463 28226 503 28302
rect 575 28226 629 28302
rect 701 28226 749 28302
rect 821 28226 866 28302
rect 463 28184 866 28226
rect 463 28108 503 28184
rect 575 28108 629 28184
rect 701 28108 749 28184
rect 821 28108 866 28184
rect 463 28072 866 28108
rect 25025 28302 25428 28360
rect 25025 28226 25068 28302
rect 25140 28226 25194 28302
rect 25266 28226 25314 28302
rect 25386 28226 25428 28302
rect 25025 28184 25428 28226
rect 25025 28108 25068 28184
rect 25140 28108 25194 28184
rect 25266 28108 25314 28184
rect 25386 28108 25428 28184
rect 25025 28072 25428 28108
rect 463 27520 863 27545
rect 463 27444 503 27520
rect 575 27444 629 27520
rect 701 27444 749 27520
rect 821 27444 863 27520
rect 463 27402 863 27444
rect 463 27326 503 27402
rect 575 27326 629 27402
rect 701 27326 749 27402
rect 821 27326 863 27402
rect 463 27290 863 27326
rect 25028 27520 25428 27545
rect 25028 27444 25068 27520
rect 25140 27444 25194 27520
rect 25266 27444 25314 27520
rect 25386 27444 25428 27520
rect 25028 27402 25428 27444
rect 25028 27326 25068 27402
rect 25140 27326 25194 27402
rect 25266 27326 25314 27402
rect 25386 27326 25428 27402
rect 25028 27290 25428 27326
rect 463 27061 863 27111
rect 463 26985 504 27061
rect 576 26985 626 27061
rect 698 26985 752 27061
rect 824 26985 863 27061
rect 463 26914 863 26985
rect 463 26838 504 26914
rect 576 26838 626 26914
rect 698 26838 752 26914
rect 824 26838 863 26914
rect 463 26777 863 26838
rect 463 26701 504 26777
rect 576 26701 626 26777
rect 698 26701 752 26777
rect 824 26701 863 26777
rect 463 26651 863 26701
rect 25970 26130 26370 26155
rect 25970 26054 26010 26130
rect 26082 26054 26136 26130
rect 26208 26054 26256 26130
rect 26328 26054 26370 26130
rect 25970 26012 26370 26054
rect 25970 25936 26010 26012
rect 26082 25936 26136 26012
rect 26208 25936 26256 26012
rect 26328 25936 26370 26012
rect 25970 25900 26370 25936
rect 463 25294 863 25349
rect 463 25218 504 25294
rect 576 25218 626 25294
rect 698 25218 752 25294
rect 824 25218 863 25294
rect 463 25147 863 25218
rect 463 25071 504 25147
rect 576 25071 626 25147
rect 698 25071 752 25147
rect 824 25071 863 25147
rect 463 25010 863 25071
rect 463 24934 504 25010
rect 576 24934 626 25010
rect 698 24934 752 25010
rect 824 24934 863 25010
rect 463 24885 863 24934
rect 463 24884 862 24885
rect 463 24608 863 24633
rect 463 24532 503 24608
rect 575 24532 629 24608
rect 701 24532 749 24608
rect 821 24532 863 24608
rect 463 24490 863 24532
rect 463 24414 503 24490
rect 575 24414 629 24490
rect 701 24414 749 24490
rect 821 24414 863 24490
rect 463 24378 863 24414
rect 25028 24559 25428 24584
rect 25028 24483 25068 24559
rect 25140 24483 25194 24559
rect 25266 24483 25314 24559
rect 25386 24483 25428 24559
rect 25028 24441 25428 24483
rect 25028 24365 25068 24441
rect 25140 24365 25194 24441
rect 25266 24365 25314 24441
rect 25386 24365 25428 24441
rect 25028 24329 25428 24365
rect 463 23604 863 23629
rect 463 23528 503 23604
rect 575 23528 629 23604
rect 701 23528 749 23604
rect 821 23528 863 23604
rect 463 23486 863 23528
rect 463 23410 503 23486
rect 575 23410 629 23486
rect 701 23410 749 23486
rect 821 23410 863 23486
rect 463 23374 863 23410
rect 25027 23442 25427 23467
rect 25027 23366 25068 23442
rect 25140 23366 25194 23442
rect 25266 23366 25314 23442
rect 25386 23366 25427 23442
rect 25027 23324 25427 23366
rect 25027 23248 25068 23324
rect 25140 23248 25194 23324
rect 25266 23248 25314 23324
rect 25386 23248 25427 23324
rect 25027 23212 25427 23248
rect 463 23060 863 23109
rect 463 22984 504 23060
rect 576 22984 626 23060
rect 698 22984 752 23060
rect 824 22984 863 23060
rect 463 22913 863 22984
rect 463 22837 504 22913
rect 576 22837 626 22913
rect 698 22837 752 22913
rect 824 22837 863 22913
rect 463 22776 863 22837
rect 463 22700 504 22776
rect 576 22700 626 22776
rect 698 22700 752 22776
rect 824 22700 863 22776
rect 463 22650 863 22700
rect 25970 21971 26370 21996
rect 25970 21895 26010 21971
rect 26082 21895 26136 21971
rect 26208 21895 26256 21971
rect 26328 21895 26370 21971
rect 25970 21853 26370 21895
rect 25970 21777 26010 21853
rect 26082 21777 26136 21853
rect 26208 21777 26256 21853
rect 26328 21777 26370 21853
rect 25970 21741 26370 21777
rect 463 21300 863 21349
rect 463 21224 504 21300
rect 576 21224 626 21300
rect 698 21224 752 21300
rect 824 21224 863 21300
rect 463 21153 863 21224
rect 463 21077 504 21153
rect 576 21077 626 21153
rect 698 21077 752 21153
rect 824 21077 863 21153
rect 463 21016 863 21077
rect 463 20940 504 21016
rect 576 20940 626 21016
rect 698 20940 752 21016
rect 824 20940 863 21016
rect 463 20890 863 20940
rect 463 20626 864 20651
rect 463 20550 503 20626
rect 575 20550 629 20626
rect 701 20550 749 20626
rect 821 20550 864 20626
rect 463 20508 864 20550
rect 463 20432 503 20508
rect 575 20432 629 20508
rect 701 20432 749 20508
rect 821 20432 864 20508
rect 463 20396 864 20432
rect 25028 20599 25428 20624
rect 25028 20523 25068 20599
rect 25140 20523 25194 20599
rect 25266 20523 25314 20599
rect 25386 20523 25428 20599
rect 25028 20481 25428 20523
rect 25028 20405 25068 20481
rect 25140 20405 25194 20481
rect 25266 20405 25314 20481
rect 25386 20405 25428 20481
rect 25028 20369 25428 20405
rect 463 19544 864 19569
rect 463 19468 503 19544
rect 575 19468 629 19544
rect 701 19468 749 19544
rect 821 19468 864 19544
rect 463 19426 864 19468
rect 463 19350 503 19426
rect 575 19350 629 19426
rect 701 19350 749 19426
rect 821 19350 864 19426
rect 463 19314 864 19350
rect 25028 19424 25428 19449
rect 25028 19348 25068 19424
rect 25140 19348 25194 19424
rect 25266 19348 25314 19424
rect 25386 19348 25428 19424
rect 25028 19306 25428 19348
rect 25028 19230 25068 19306
rect 25140 19230 25194 19306
rect 25266 19230 25314 19306
rect 25386 19230 25428 19306
rect 25028 19194 25428 19230
rect 463 19060 863 19109
rect 463 18984 504 19060
rect 576 18984 626 19060
rect 698 18984 752 19060
rect 824 18984 863 19060
rect 463 18913 863 18984
rect 463 18837 504 18913
rect 576 18837 626 18913
rect 698 18837 752 18913
rect 824 18837 863 18913
rect 463 18776 863 18837
rect 463 18700 504 18776
rect 576 18700 626 18776
rect 698 18700 752 18776
rect 824 18700 863 18776
rect 463 18650 863 18700
rect 25970 18181 26370 18206
rect 25970 18105 26010 18181
rect 26082 18105 26136 18181
rect 26208 18105 26256 18181
rect 26328 18105 26370 18181
rect 25970 18063 26370 18105
rect 25970 17987 26010 18063
rect 26082 17987 26136 18063
rect 26208 17987 26256 18063
rect 26328 17987 26370 18063
rect 25970 17951 26370 17987
rect 463 17301 863 17350
rect 463 17225 504 17301
rect 576 17225 626 17301
rect 698 17225 752 17301
rect 824 17225 863 17301
rect 463 17154 863 17225
rect 463 17078 504 17154
rect 576 17078 626 17154
rect 698 17078 752 17154
rect 824 17078 863 17154
rect 463 17017 863 17078
rect 463 16941 504 17017
rect 576 16941 626 17017
rect 698 16941 752 17017
rect 824 16941 863 17017
rect 463 16891 863 16941
rect 463 16669 864 16694
rect 463 16593 503 16669
rect 575 16593 629 16669
rect 701 16593 749 16669
rect 821 16593 864 16669
rect 463 16551 864 16593
rect 463 16475 503 16551
rect 575 16475 629 16551
rect 701 16475 749 16551
rect 821 16475 864 16551
rect 463 16439 864 16475
rect 25027 16583 25427 16608
rect 25027 16507 25068 16583
rect 25140 16507 25194 16583
rect 25266 16507 25314 16583
rect 25386 16507 25427 16583
rect 25027 16465 25427 16507
rect 25027 16389 25068 16465
rect 25140 16389 25194 16465
rect 25266 16389 25314 16465
rect 25386 16389 25427 16465
rect 25027 16353 25427 16389
rect 463 15568 864 15593
rect 463 15492 503 15568
rect 575 15492 629 15568
rect 701 15492 749 15568
rect 821 15492 864 15568
rect 463 15450 864 15492
rect 463 15374 503 15450
rect 575 15374 629 15450
rect 701 15374 749 15450
rect 821 15374 864 15450
rect 463 15338 864 15374
rect 25027 15412 25427 15437
rect 25027 15336 25068 15412
rect 25140 15336 25194 15412
rect 25266 15336 25314 15412
rect 25386 15336 25427 15412
rect 25027 15294 25427 15336
rect 25027 15218 25068 15294
rect 25140 15218 25194 15294
rect 25266 15218 25314 15294
rect 25386 15218 25427 15294
rect 25027 15182 25427 15218
rect 463 15060 863 15109
rect 463 14984 504 15060
rect 576 14984 626 15060
rect 698 14984 752 15060
rect 824 14984 863 15060
rect 463 14913 863 14984
rect 463 14837 504 14913
rect 576 14837 626 14913
rect 698 14837 752 14913
rect 824 14837 863 14913
rect 463 14776 863 14837
rect 463 14700 504 14776
rect 576 14700 626 14776
rect 698 14700 752 14776
rect 824 14700 863 14776
rect 463 14650 863 14700
rect 25970 14074 26370 14099
rect 25970 13998 26010 14074
rect 26082 13998 26136 14074
rect 26208 13998 26256 14074
rect 26328 13998 26370 14074
rect 25970 13956 26370 13998
rect 25970 13880 26010 13956
rect 26082 13880 26136 13956
rect 26208 13880 26256 13956
rect 26328 13880 26370 13956
rect 25970 13844 26370 13880
rect 463 13300 863 13349
rect 463 13224 504 13300
rect 576 13224 626 13300
rect 698 13224 752 13300
rect 824 13224 863 13300
rect 463 13153 863 13224
rect 463 13077 504 13153
rect 576 13077 626 13153
rect 698 13077 752 13153
rect 824 13077 863 13153
rect 463 13016 863 13077
rect 463 12940 504 13016
rect 576 12940 626 13016
rect 698 12940 752 13016
rect 824 12940 863 13016
rect 463 12890 863 12940
rect 463 12702 865 12727
rect 463 12626 503 12702
rect 575 12626 629 12702
rect 701 12626 749 12702
rect 821 12626 865 12702
rect 463 12584 865 12626
rect 463 12508 503 12584
rect 575 12508 629 12584
rect 701 12508 749 12584
rect 821 12508 865 12584
rect 463 12472 865 12508
rect 25027 12651 25427 12676
rect 25027 12575 25068 12651
rect 25140 12575 25194 12651
rect 25266 12575 25314 12651
rect 25386 12575 25427 12651
rect 25027 12533 25427 12575
rect 25027 12457 25068 12533
rect 25140 12457 25194 12533
rect 25266 12457 25314 12533
rect 25386 12457 25427 12533
rect 25027 12421 25427 12457
rect 463 11486 866 11511
rect 463 11410 503 11486
rect 575 11410 629 11486
rect 701 11410 749 11486
rect 821 11410 866 11486
rect 463 11368 866 11410
rect 463 11292 503 11368
rect 575 11292 629 11368
rect 701 11292 749 11368
rect 821 11292 866 11368
rect 463 11256 866 11292
rect 25027 11437 25427 11462
rect 25027 11361 25068 11437
rect 25140 11361 25194 11437
rect 25266 11361 25314 11437
rect 25386 11361 25427 11437
rect 25027 11319 25427 11361
rect 25027 11243 25068 11319
rect 25140 11243 25194 11319
rect 25266 11243 25314 11319
rect 25386 11243 25427 11319
rect 25027 11207 25427 11243
rect 463 11060 863 11109
rect 463 10984 504 11060
rect 576 10984 626 11060
rect 698 10984 752 11060
rect 824 10984 863 11060
rect 463 10913 863 10984
rect 463 10837 504 10913
rect 576 10837 626 10913
rect 698 10837 752 10913
rect 824 10837 863 10913
rect 463 10776 863 10837
rect 463 10700 504 10776
rect 576 10700 626 10776
rect 698 10700 752 10776
rect 824 10700 863 10776
rect 463 10650 863 10700
rect 25970 10256 26370 10281
rect 25970 10180 26010 10256
rect 26082 10180 26136 10256
rect 26208 10180 26256 10256
rect 26328 10180 26370 10256
rect 25970 10138 26370 10180
rect 25970 10062 26010 10138
rect 26082 10062 26136 10138
rect 26208 10062 26256 10138
rect 26328 10062 26370 10138
rect 25970 10026 26370 10062
rect 463 9300 863 9349
rect 463 9224 504 9300
rect 576 9224 626 9300
rect 698 9224 752 9300
rect 824 9224 863 9300
rect 463 9153 863 9224
rect 463 9077 504 9153
rect 576 9077 626 9153
rect 698 9077 752 9153
rect 824 9077 863 9153
rect 463 9016 863 9077
rect 463 8940 504 9016
rect 576 8940 626 9016
rect 698 8940 752 9016
rect 824 8940 863 9016
rect 463 8890 863 8940
rect 463 8621 864 8646
rect 463 8545 503 8621
rect 575 8545 629 8621
rect 701 8545 749 8621
rect 821 8545 864 8621
rect 463 8503 864 8545
rect 463 8427 503 8503
rect 575 8427 629 8503
rect 701 8427 749 8503
rect 821 8427 864 8503
rect 463 8391 864 8427
rect 25028 8594 25428 8619
rect 25028 8518 25068 8594
rect 25140 8518 25194 8594
rect 25266 8518 25314 8594
rect 25386 8518 25428 8594
rect 25028 8476 25428 8518
rect 25028 8400 25068 8476
rect 25140 8400 25194 8476
rect 25266 8400 25314 8476
rect 25386 8400 25428 8476
rect 25028 8364 25428 8400
rect 463 7499 864 7524
rect 463 7423 503 7499
rect 575 7423 629 7499
rect 701 7423 749 7499
rect 821 7423 864 7499
rect 463 7381 864 7423
rect 463 7305 503 7381
rect 575 7305 629 7381
rect 701 7305 749 7381
rect 821 7305 864 7381
rect 463 7269 864 7305
rect 25027 7437 25427 7462
rect 25027 7361 25068 7437
rect 25140 7361 25194 7437
rect 25266 7361 25314 7437
rect 25386 7361 25427 7437
rect 25027 7319 25427 7361
rect 25027 7243 25068 7319
rect 25140 7243 25194 7319
rect 25266 7243 25314 7319
rect 25386 7243 25427 7319
rect 25027 7207 25427 7243
rect 463 7061 863 7110
rect 463 6985 504 7061
rect 576 6985 626 7061
rect 698 6985 752 7061
rect 824 6985 863 7061
rect 463 6914 863 6985
rect 463 6838 504 6914
rect 576 6838 626 6914
rect 698 6838 752 6914
rect 824 6838 863 6914
rect 463 6777 863 6838
rect 463 6701 504 6777
rect 576 6701 626 6777
rect 698 6701 752 6777
rect 824 6701 863 6777
rect 463 6651 863 6701
rect 25970 6292 26370 6317
rect 25970 6216 26010 6292
rect 26082 6216 26136 6292
rect 26208 6216 26256 6292
rect 26328 6216 26370 6292
rect 25970 6174 26370 6216
rect 25970 6098 26010 6174
rect 26082 6098 26136 6174
rect 26208 6098 26256 6174
rect 26328 6098 26370 6174
rect 25970 6062 26370 6098
rect 463 5299 863 5348
rect 463 5223 504 5299
rect 576 5223 626 5299
rect 698 5223 752 5299
rect 824 5223 863 5299
rect 463 5152 863 5223
rect 463 5076 504 5152
rect 576 5076 626 5152
rect 698 5076 752 5152
rect 824 5076 863 5152
rect 463 5015 863 5076
rect 463 4939 504 5015
rect 576 4939 626 5015
rect 698 4939 752 5015
rect 824 4939 863 5015
rect 463 4889 863 4939
rect 463 4639 863 4664
rect 463 4563 503 4639
rect 575 4563 629 4639
rect 701 4563 749 4639
rect 821 4563 863 4639
rect 463 4521 863 4563
rect 463 4445 503 4521
rect 575 4445 629 4521
rect 701 4445 749 4521
rect 821 4445 863 4521
rect 463 4409 863 4445
rect 25028 4594 25428 4619
rect 25028 4518 25068 4594
rect 25140 4518 25194 4594
rect 25266 4518 25314 4594
rect 25386 4518 25428 4594
rect 25028 4476 25428 4518
rect 25028 4400 25068 4476
rect 25140 4400 25194 4476
rect 25266 4400 25314 4476
rect 25386 4400 25428 4476
rect 25028 4364 25428 4400
rect 463 3528 863 3553
rect 463 3452 503 3528
rect 575 3452 629 3528
rect 701 3452 749 3528
rect 821 3452 863 3528
rect 463 3410 863 3452
rect 463 3334 503 3410
rect 575 3334 629 3410
rect 701 3334 749 3410
rect 821 3334 863 3410
rect 463 3298 863 3334
rect 25027 3437 25427 3462
rect 25027 3361 25068 3437
rect 25140 3361 25194 3437
rect 25266 3361 25314 3437
rect 25386 3361 25427 3437
rect 25027 3319 25427 3361
rect 25027 3243 25068 3319
rect 25140 3243 25194 3319
rect 25266 3243 25314 3319
rect 25386 3243 25427 3319
rect 25027 3207 25427 3243
rect 463 3061 863 3110
rect 463 2985 504 3061
rect 576 2985 626 3061
rect 698 2985 752 3061
rect 824 2985 863 3061
rect 463 2914 863 2985
rect 463 2838 504 2914
rect 576 2838 626 2914
rect 698 2838 752 2914
rect 824 2838 863 2914
rect 463 2777 863 2838
rect 463 2701 504 2777
rect 576 2701 626 2777
rect 698 2701 752 2777
rect 824 2701 863 2777
rect 463 2651 863 2701
rect 25970 2280 26370 2305
rect 25970 2204 26010 2280
rect 26082 2204 26136 2280
rect 26208 2204 26256 2280
rect 26328 2204 26370 2280
rect 25970 2162 26370 2204
rect 25970 2086 26010 2162
rect 26082 2086 26136 2162
rect 26208 2086 26256 2162
rect 26328 2086 26370 2162
rect 25970 2050 26370 2086
rect 463 1300 863 1349
rect 463 1224 504 1300
rect 576 1224 626 1300
rect 698 1224 752 1300
rect 824 1224 863 1300
rect 463 1153 863 1224
rect 463 1077 504 1153
rect 576 1077 626 1153
rect 698 1077 752 1153
rect 824 1077 863 1153
rect 463 1016 863 1077
rect 463 940 504 1016
rect 576 940 626 1016
rect 698 940 752 1016
rect 824 940 863 1016
rect 463 890 863 940
rect 463 705 865 730
rect 463 629 503 705
rect 575 629 629 705
rect 701 629 749 705
rect 821 629 865 705
rect 463 587 865 629
rect 463 511 503 587
rect 575 511 629 587
rect 701 511 749 587
rect 821 511 865 587
rect 463 475 865 511
rect 25028 594 25428 619
rect 25028 518 25068 594
rect 25140 518 25194 594
rect 25266 518 25314 594
rect 25386 518 25428 594
rect 25028 476 25428 518
rect 25028 400 25068 476
rect 25140 400 25194 476
rect 25266 400 25314 476
rect 25386 400 25428 476
rect 25028 364 25428 400
<< via3 >>
rect 503 63376 575 63452
rect 629 63376 701 63452
rect 749 63376 821 63452
rect 503 63258 575 63334
rect 629 63258 701 63334
rect 749 63258 821 63334
rect 25068 63416 25140 63492
rect 25194 63416 25266 63492
rect 25314 63416 25386 63492
rect 25068 63298 25140 63374
rect 25194 63298 25266 63374
rect 25314 63298 25386 63374
rect 504 62984 576 63060
rect 626 62984 698 63060
rect 752 62984 824 63060
rect 504 62837 576 62913
rect 626 62837 698 62913
rect 752 62837 824 62913
rect 504 62700 576 62776
rect 626 62700 698 62776
rect 752 62700 824 62776
rect 26010 61995 26082 62071
rect 26136 61995 26208 62071
rect 26256 61995 26328 62071
rect 26010 61877 26082 61953
rect 26136 61877 26208 61953
rect 26256 61877 26328 61953
rect 504 61224 576 61300
rect 626 61224 698 61300
rect 752 61224 824 61300
rect 504 61077 576 61153
rect 626 61077 698 61153
rect 752 61077 824 61153
rect 504 60940 576 61016
rect 626 60940 698 61016
rect 752 60940 824 61016
rect 503 60703 575 60779
rect 629 60703 701 60779
rect 749 60703 821 60779
rect 503 60585 575 60661
rect 629 60585 701 60661
rect 749 60585 821 60661
rect 25068 60619 25140 60695
rect 25194 60619 25266 60695
rect 25314 60619 25386 60695
rect 25068 60501 25140 60577
rect 25194 60501 25266 60577
rect 25314 60501 25386 60577
rect 503 59374 575 59450
rect 629 59374 701 59450
rect 749 59374 821 59450
rect 503 59256 575 59332
rect 629 59256 701 59332
rect 749 59256 821 59332
rect 25068 59416 25140 59492
rect 25194 59416 25266 59492
rect 25314 59416 25386 59492
rect 25068 59298 25140 59374
rect 25194 59298 25266 59374
rect 25314 59298 25386 59374
rect 504 58984 576 59060
rect 626 58984 698 59060
rect 752 58984 824 59060
rect 504 58837 576 58913
rect 626 58837 698 58913
rect 752 58837 824 58913
rect 504 58700 576 58776
rect 626 58700 698 58776
rect 752 58700 824 58776
rect 26010 57982 26082 58058
rect 26136 57982 26208 58058
rect 26256 57982 26328 58058
rect 26010 57864 26082 57940
rect 26136 57864 26208 57940
rect 26256 57864 26328 57940
rect 504 57225 576 57301
rect 626 57225 698 57301
rect 752 57225 824 57301
rect 504 57078 576 57154
rect 626 57078 698 57154
rect 752 57078 824 57154
rect 504 56941 576 57017
rect 626 56941 698 57017
rect 752 56941 824 57017
rect 503 56634 575 56710
rect 629 56634 701 56710
rect 749 56634 821 56710
rect 503 56516 575 56592
rect 629 56516 701 56592
rect 749 56516 821 56592
rect 25068 56619 25140 56695
rect 25194 56619 25266 56695
rect 25314 56619 25386 56695
rect 25068 56501 25140 56577
rect 25194 56501 25266 56577
rect 25314 56501 25386 56577
rect 503 55456 575 55532
rect 629 55456 701 55532
rect 749 55456 821 55532
rect 503 55338 575 55414
rect 629 55338 701 55414
rect 749 55338 821 55414
rect 25068 55416 25140 55492
rect 25194 55416 25266 55492
rect 25314 55416 25386 55492
rect 25068 55298 25140 55374
rect 25194 55298 25266 55374
rect 25314 55298 25386 55374
rect 504 54984 576 55060
rect 626 54984 698 55060
rect 752 54984 824 55060
rect 504 54837 576 54913
rect 626 54837 698 54913
rect 752 54837 824 54913
rect 504 54700 576 54776
rect 626 54700 698 54776
rect 752 54700 824 54776
rect 26010 53981 26082 54057
rect 26136 53981 26208 54057
rect 26256 53981 26328 54057
rect 26010 53863 26082 53939
rect 26136 53863 26208 53939
rect 26256 53863 26328 53939
rect 504 53225 576 53301
rect 626 53225 698 53301
rect 752 53225 824 53301
rect 504 53078 576 53154
rect 626 53078 698 53154
rect 752 53078 824 53154
rect 504 52941 576 53017
rect 626 52941 698 53017
rect 752 52941 824 53017
rect 503 52608 575 52684
rect 629 52608 701 52684
rect 749 52608 821 52684
rect 503 52490 575 52566
rect 629 52490 701 52566
rect 749 52490 821 52566
rect 25068 52619 25140 52695
rect 25194 52619 25266 52695
rect 25314 52619 25386 52695
rect 25068 52501 25140 52577
rect 25194 52501 25266 52577
rect 25314 52501 25386 52577
rect 503 51405 575 51481
rect 629 51405 701 51481
rect 749 51405 821 51481
rect 503 51287 575 51363
rect 629 51287 701 51363
rect 749 51287 821 51363
rect 25068 51470 25140 51546
rect 25194 51470 25266 51546
rect 25314 51470 25386 51546
rect 25068 51352 25140 51428
rect 25194 51352 25266 51428
rect 25314 51352 25386 51428
rect 504 50984 576 51060
rect 626 50984 698 51060
rect 752 50984 824 51060
rect 504 50837 576 50913
rect 626 50837 698 50913
rect 752 50837 824 50913
rect 504 50700 576 50776
rect 626 50700 698 50776
rect 752 50700 824 50776
rect 26010 50020 26082 50096
rect 26136 50020 26208 50096
rect 26256 50020 26328 50096
rect 26010 49902 26082 49978
rect 26136 49902 26208 49978
rect 26256 49902 26328 49978
rect 504 49223 576 49299
rect 626 49223 698 49299
rect 752 49223 824 49299
rect 504 49076 576 49152
rect 626 49076 698 49152
rect 752 49076 824 49152
rect 504 48939 576 49015
rect 626 48939 698 49015
rect 752 48939 824 49015
rect 503 48628 575 48704
rect 629 48628 701 48704
rect 749 48628 821 48704
rect 503 48510 575 48586
rect 629 48510 701 48586
rect 749 48510 821 48586
rect 25068 48554 25140 48630
rect 25194 48554 25266 48630
rect 25314 48554 25386 48630
rect 25068 48436 25140 48512
rect 25194 48436 25266 48512
rect 25314 48436 25386 48512
rect 503 47421 575 47497
rect 629 47421 701 47497
rect 749 47421 821 47497
rect 503 47303 575 47379
rect 629 47303 701 47379
rect 749 47303 821 47379
rect 25068 47371 25140 47447
rect 25194 47371 25266 47447
rect 25314 47371 25386 47447
rect 25068 47253 25140 47329
rect 25194 47253 25266 47329
rect 25314 47253 25386 47329
rect 504 46984 576 47060
rect 626 46984 698 47060
rect 752 46984 824 47060
rect 504 46837 576 46913
rect 626 46837 698 46913
rect 752 46837 824 46913
rect 504 46700 576 46776
rect 626 46700 698 46776
rect 752 46700 824 46776
rect 26010 46003 26082 46079
rect 26136 46003 26208 46079
rect 26256 46003 26328 46079
rect 26010 45885 26082 45961
rect 26136 45885 26208 45961
rect 26256 45885 26328 45961
rect 504 45225 576 45301
rect 626 45225 698 45301
rect 752 45225 824 45301
rect 504 45078 576 45154
rect 626 45078 698 45154
rect 752 45078 824 45154
rect 504 44941 576 45017
rect 626 44941 698 45017
rect 752 44941 824 45017
rect 503 44655 575 44731
rect 629 44655 701 44731
rect 749 44655 821 44731
rect 503 44537 575 44613
rect 629 44537 701 44613
rect 749 44537 821 44613
rect 25068 44499 25140 44575
rect 25194 44499 25266 44575
rect 25314 44499 25386 44575
rect 25068 44381 25140 44457
rect 25194 44381 25266 44457
rect 25314 44381 25386 44457
rect 503 43468 575 43544
rect 629 43468 701 43544
rect 749 43468 821 43544
rect 503 43350 575 43426
rect 629 43350 701 43426
rect 749 43350 821 43426
rect 25068 43364 25140 43440
rect 25194 43364 25266 43440
rect 25314 43364 25386 43440
rect 25068 43246 25140 43322
rect 25194 43246 25266 43322
rect 25314 43246 25386 43322
rect 504 42984 576 43060
rect 626 42984 698 43060
rect 752 42984 824 43060
rect 504 42837 576 42913
rect 626 42837 698 42913
rect 752 42837 824 42913
rect 504 42700 576 42776
rect 626 42700 698 42776
rect 752 42700 824 42776
rect 26010 42082 26082 42158
rect 26136 42082 26208 42158
rect 26256 42082 26328 42158
rect 26010 41964 26082 42040
rect 26136 41964 26208 42040
rect 26256 41964 26328 42040
rect 504 41225 576 41301
rect 626 41225 698 41301
rect 752 41225 824 41301
rect 504 41078 576 41154
rect 626 41078 698 41154
rect 752 41078 824 41154
rect 504 40941 576 41017
rect 626 40941 698 41017
rect 752 40941 824 41017
rect 503 40646 575 40722
rect 629 40646 701 40722
rect 749 40646 821 40722
rect 503 40528 575 40604
rect 629 40528 701 40604
rect 749 40528 821 40604
rect 25068 40605 25140 40681
rect 25194 40605 25266 40681
rect 25314 40605 25386 40681
rect 25068 40487 25140 40563
rect 25194 40487 25266 40563
rect 25314 40487 25386 40563
rect 503 39493 575 39569
rect 629 39493 701 39569
rect 749 39493 821 39569
rect 503 39375 575 39451
rect 629 39375 701 39451
rect 749 39375 821 39451
rect 25068 39452 25140 39528
rect 25194 39452 25266 39528
rect 25314 39452 25386 39528
rect 25068 39334 25140 39410
rect 25194 39334 25266 39410
rect 25314 39334 25386 39410
rect 504 38984 576 39060
rect 626 38984 698 39060
rect 752 38984 824 39060
rect 504 38837 576 38913
rect 626 38837 698 38913
rect 752 38837 824 38913
rect 504 38700 576 38776
rect 626 38700 698 38776
rect 752 38700 824 38776
rect 26010 37824 26082 37900
rect 26136 37824 26208 37900
rect 26256 37824 26328 37900
rect 26010 37706 26082 37782
rect 26136 37706 26208 37782
rect 26256 37706 26328 37782
rect 504 37224 576 37300
rect 626 37224 698 37300
rect 752 37224 824 37300
rect 504 37077 576 37153
rect 626 37077 698 37153
rect 752 37077 824 37153
rect 504 36940 576 37016
rect 626 36940 698 37016
rect 752 36940 824 37016
rect 503 36433 575 36509
rect 629 36433 701 36509
rect 749 36433 821 36509
rect 503 36315 575 36391
rect 629 36315 701 36391
rect 749 36315 821 36391
rect 25068 36336 25140 36412
rect 25194 36336 25266 36412
rect 25314 36336 25386 36412
rect 25068 36218 25140 36294
rect 25194 36218 25266 36294
rect 25314 36218 25386 36294
rect 2249 35869 2257 35925
rect 2257 35869 2313 35925
rect 2249 35861 2313 35869
rect 2337 35869 2393 35925
rect 2393 35869 2401 35925
rect 2337 35861 2401 35869
rect 2249 35789 2257 35845
rect 2257 35789 2313 35845
rect 2249 35781 2313 35789
rect 2337 35789 2393 35845
rect 2393 35789 2401 35845
rect 2337 35781 2401 35789
rect 4192 35841 4256 35905
rect 4280 35841 4344 35905
rect 4192 35761 4256 35825
rect 4280 35761 4344 35825
rect 32 35661 111 35741
rect 156 35661 157 35741
rect 157 35661 236 35741
rect 282 35661 362 35741
rect 32 35555 111 35635
rect 156 35555 157 35635
rect 157 35555 236 35635
rect 282 35555 362 35635
rect 25535 35646 25615 35726
rect 25660 35646 25740 35726
rect 25785 35646 25865 35726
rect 25534 35526 25614 35606
rect 25659 35526 25739 35606
rect 25784 35526 25864 35606
rect 478 35130 562 35131
rect 478 35052 479 35130
rect 479 35052 561 35130
rect 561 35052 562 35130
rect 478 35051 562 35052
rect 592 35130 676 35131
rect 592 35052 593 35130
rect 593 35052 675 35130
rect 675 35052 676 35130
rect 592 35051 676 35052
rect 706 35130 790 35131
rect 706 35052 707 35130
rect 707 35052 789 35130
rect 789 35052 790 35130
rect 706 35051 790 35052
rect 25061 34892 25141 34972
rect 25186 34892 25266 34972
rect 25311 34892 25391 34972
rect 25060 34772 25140 34852
rect 25185 34772 25265 34852
rect 25310 34772 25390 34852
rect 15 34586 99 34587
rect 15 34508 16 34586
rect 16 34508 98 34586
rect 98 34508 99 34586
rect 15 34507 99 34508
rect 129 34586 213 34587
rect 129 34508 130 34586
rect 130 34508 212 34586
rect 212 34508 213 34586
rect 129 34507 213 34508
rect 243 34586 327 34587
rect 243 34508 244 34586
rect 244 34508 326 34586
rect 326 34508 327 34586
rect 243 34507 327 34508
rect 25069 34316 25141 34392
rect 25191 34316 25263 34392
rect 25317 34316 25389 34392
rect 25069 34169 25141 34245
rect 25191 34169 25263 34245
rect 25317 34169 25389 34245
rect 478 34042 562 34043
rect 478 33964 479 34042
rect 479 33964 561 34042
rect 561 33964 562 34042
rect 478 33963 562 33964
rect 592 34042 676 34043
rect 592 33964 593 34042
rect 593 33964 675 34042
rect 675 33964 676 34042
rect 592 33963 676 33964
rect 706 34042 790 34043
rect 706 33964 707 34042
rect 707 33964 789 34042
rect 789 33964 790 34042
rect 706 33963 790 33964
rect 25069 34032 25141 34108
rect 25191 34032 25263 34108
rect 25317 34032 25389 34108
rect 15 33498 99 33499
rect 15 33420 16 33498
rect 16 33420 98 33498
rect 98 33420 99 33498
rect 15 33419 99 33420
rect 129 33498 213 33499
rect 129 33420 130 33498
rect 130 33420 212 33498
rect 212 33420 213 33498
rect 129 33419 213 33420
rect 243 33498 327 33499
rect 243 33420 244 33498
rect 244 33420 326 33498
rect 326 33420 327 33498
rect 243 33419 327 33420
rect 24560 33396 24640 33476
rect 24685 33396 24765 33476
rect 24810 33396 24890 33476
rect 24559 33276 24639 33356
rect 24684 33276 24764 33356
rect 24809 33276 24889 33356
rect 25535 33396 25615 33476
rect 25660 33396 25740 33476
rect 25785 33396 25865 33476
rect 25534 33276 25614 33356
rect 25659 33276 25739 33356
rect 25784 33276 25864 33356
rect 478 32954 562 32955
rect 478 32876 479 32954
rect 479 32876 561 32954
rect 561 32876 562 32954
rect 478 32875 562 32876
rect 592 32954 676 32955
rect 592 32876 593 32954
rect 593 32876 675 32954
rect 675 32876 676 32954
rect 592 32875 676 32876
rect 706 32954 790 32955
rect 706 32876 707 32954
rect 707 32876 789 32954
rect 789 32876 790 32954
rect 706 32875 790 32876
rect 25069 32556 25141 32632
rect 25191 32556 25263 32632
rect 25317 32556 25389 32632
rect 3136 32401 3144 32463
rect 3144 32401 3200 32463
rect 3136 32399 3200 32401
rect 3224 32401 3280 32463
rect 3280 32401 3288 32463
rect 3224 32399 3288 32401
rect 25069 32409 25141 32485
rect 25191 32409 25263 32485
rect 25317 32409 25389 32485
rect 25069 32272 25141 32348
rect 25191 32272 25263 32348
rect 25317 32272 25389 32348
rect 25060 31837 25140 31917
rect 25185 31837 25265 31917
rect 25310 31837 25390 31917
rect 25059 31717 25139 31797
rect 25184 31717 25264 31797
rect 25309 31717 25389 31797
rect 503 28226 575 28302
rect 629 28226 701 28302
rect 749 28226 821 28302
rect 503 28108 575 28184
rect 629 28108 701 28184
rect 749 28108 821 28184
rect 25068 28226 25140 28302
rect 25194 28226 25266 28302
rect 25314 28226 25386 28302
rect 25068 28108 25140 28184
rect 25194 28108 25266 28184
rect 25314 28108 25386 28184
rect 503 27444 575 27520
rect 629 27444 701 27520
rect 749 27444 821 27520
rect 503 27326 575 27402
rect 629 27326 701 27402
rect 749 27326 821 27402
rect 25068 27444 25140 27520
rect 25194 27444 25266 27520
rect 25314 27444 25386 27520
rect 25068 27326 25140 27402
rect 25194 27326 25266 27402
rect 25314 27326 25386 27402
rect 504 26985 576 27061
rect 626 26985 698 27061
rect 752 26985 824 27061
rect 504 26838 576 26914
rect 626 26838 698 26914
rect 752 26838 824 26914
rect 504 26701 576 26777
rect 626 26701 698 26777
rect 752 26701 824 26777
rect 26010 26054 26082 26130
rect 26136 26054 26208 26130
rect 26256 26054 26328 26130
rect 26010 25936 26082 26012
rect 26136 25936 26208 26012
rect 26256 25936 26328 26012
rect 504 25218 576 25294
rect 626 25218 698 25294
rect 752 25218 824 25294
rect 504 25071 576 25147
rect 626 25071 698 25147
rect 752 25071 824 25147
rect 504 24934 576 25010
rect 626 24934 698 25010
rect 752 24934 824 25010
rect 503 24532 575 24608
rect 629 24532 701 24608
rect 749 24532 821 24608
rect 503 24414 575 24490
rect 629 24414 701 24490
rect 749 24414 821 24490
rect 25068 24483 25140 24559
rect 25194 24483 25266 24559
rect 25314 24483 25386 24559
rect 25068 24365 25140 24441
rect 25194 24365 25266 24441
rect 25314 24365 25386 24441
rect 503 23528 575 23604
rect 629 23528 701 23604
rect 749 23528 821 23604
rect 503 23410 575 23486
rect 629 23410 701 23486
rect 749 23410 821 23486
rect 25068 23366 25140 23442
rect 25194 23366 25266 23442
rect 25314 23366 25386 23442
rect 25068 23248 25140 23324
rect 25194 23248 25266 23324
rect 25314 23248 25386 23324
rect 504 22984 576 23060
rect 626 22984 698 23060
rect 752 22984 824 23060
rect 504 22837 576 22913
rect 626 22837 698 22913
rect 752 22837 824 22913
rect 504 22700 576 22776
rect 626 22700 698 22776
rect 752 22700 824 22776
rect 26010 21895 26082 21971
rect 26136 21895 26208 21971
rect 26256 21895 26328 21971
rect 26010 21777 26082 21853
rect 26136 21777 26208 21853
rect 26256 21777 26328 21853
rect 504 21224 576 21300
rect 626 21224 698 21300
rect 752 21224 824 21300
rect 504 21077 576 21153
rect 626 21077 698 21153
rect 752 21077 824 21153
rect 504 20940 576 21016
rect 626 20940 698 21016
rect 752 20940 824 21016
rect 503 20550 575 20626
rect 629 20550 701 20626
rect 749 20550 821 20626
rect 503 20432 575 20508
rect 629 20432 701 20508
rect 749 20432 821 20508
rect 25068 20523 25140 20599
rect 25194 20523 25266 20599
rect 25314 20523 25386 20599
rect 25068 20405 25140 20481
rect 25194 20405 25266 20481
rect 25314 20405 25386 20481
rect 503 19468 575 19544
rect 629 19468 701 19544
rect 749 19468 821 19544
rect 503 19350 575 19426
rect 629 19350 701 19426
rect 749 19350 821 19426
rect 25068 19348 25140 19424
rect 25194 19348 25266 19424
rect 25314 19348 25386 19424
rect 25068 19230 25140 19306
rect 25194 19230 25266 19306
rect 25314 19230 25386 19306
rect 504 18984 576 19060
rect 626 18984 698 19060
rect 752 18984 824 19060
rect 504 18837 576 18913
rect 626 18837 698 18913
rect 752 18837 824 18913
rect 504 18700 576 18776
rect 626 18700 698 18776
rect 752 18700 824 18776
rect 26010 18105 26082 18181
rect 26136 18105 26208 18181
rect 26256 18105 26328 18181
rect 26010 17987 26082 18063
rect 26136 17987 26208 18063
rect 26256 17987 26328 18063
rect 504 17225 576 17301
rect 626 17225 698 17301
rect 752 17225 824 17301
rect 504 17078 576 17154
rect 626 17078 698 17154
rect 752 17078 824 17154
rect 504 16941 576 17017
rect 626 16941 698 17017
rect 752 16941 824 17017
rect 503 16593 575 16669
rect 629 16593 701 16669
rect 749 16593 821 16669
rect 503 16475 575 16551
rect 629 16475 701 16551
rect 749 16475 821 16551
rect 25068 16507 25140 16583
rect 25194 16507 25266 16583
rect 25314 16507 25386 16583
rect 25068 16389 25140 16465
rect 25194 16389 25266 16465
rect 25314 16389 25386 16465
rect 503 15492 575 15568
rect 629 15492 701 15568
rect 749 15492 821 15568
rect 503 15374 575 15450
rect 629 15374 701 15450
rect 749 15374 821 15450
rect 25068 15336 25140 15412
rect 25194 15336 25266 15412
rect 25314 15336 25386 15412
rect 25068 15218 25140 15294
rect 25194 15218 25266 15294
rect 25314 15218 25386 15294
rect 504 14984 576 15060
rect 626 14984 698 15060
rect 752 14984 824 15060
rect 504 14837 576 14913
rect 626 14837 698 14913
rect 752 14837 824 14913
rect 504 14700 576 14776
rect 626 14700 698 14776
rect 752 14700 824 14776
rect 26010 13998 26082 14074
rect 26136 13998 26208 14074
rect 26256 13998 26328 14074
rect 26010 13880 26082 13956
rect 26136 13880 26208 13956
rect 26256 13880 26328 13956
rect 504 13224 576 13300
rect 626 13224 698 13300
rect 752 13224 824 13300
rect 504 13077 576 13153
rect 626 13077 698 13153
rect 752 13077 824 13153
rect 504 12940 576 13016
rect 626 12940 698 13016
rect 752 12940 824 13016
rect 503 12626 575 12702
rect 629 12626 701 12702
rect 749 12626 821 12702
rect 503 12508 575 12584
rect 629 12508 701 12584
rect 749 12508 821 12584
rect 25068 12575 25140 12651
rect 25194 12575 25266 12651
rect 25314 12575 25386 12651
rect 25068 12457 25140 12533
rect 25194 12457 25266 12533
rect 25314 12457 25386 12533
rect 503 11410 575 11486
rect 629 11410 701 11486
rect 749 11410 821 11486
rect 503 11292 575 11368
rect 629 11292 701 11368
rect 749 11292 821 11368
rect 25068 11361 25140 11437
rect 25194 11361 25266 11437
rect 25314 11361 25386 11437
rect 25068 11243 25140 11319
rect 25194 11243 25266 11319
rect 25314 11243 25386 11319
rect 504 10984 576 11060
rect 626 10984 698 11060
rect 752 10984 824 11060
rect 504 10837 576 10913
rect 626 10837 698 10913
rect 752 10837 824 10913
rect 504 10700 576 10776
rect 626 10700 698 10776
rect 752 10700 824 10776
rect 26010 10180 26082 10256
rect 26136 10180 26208 10256
rect 26256 10180 26328 10256
rect 26010 10062 26082 10138
rect 26136 10062 26208 10138
rect 26256 10062 26328 10138
rect 504 9224 576 9300
rect 626 9224 698 9300
rect 752 9224 824 9300
rect 504 9077 576 9153
rect 626 9077 698 9153
rect 752 9077 824 9153
rect 504 8940 576 9016
rect 626 8940 698 9016
rect 752 8940 824 9016
rect 503 8545 575 8621
rect 629 8545 701 8621
rect 749 8545 821 8621
rect 503 8427 575 8503
rect 629 8427 701 8503
rect 749 8427 821 8503
rect 25068 8518 25140 8594
rect 25194 8518 25266 8594
rect 25314 8518 25386 8594
rect 25068 8400 25140 8476
rect 25194 8400 25266 8476
rect 25314 8400 25386 8476
rect 503 7423 575 7499
rect 629 7423 701 7499
rect 749 7423 821 7499
rect 503 7305 575 7381
rect 629 7305 701 7381
rect 749 7305 821 7381
rect 25068 7361 25140 7437
rect 25194 7361 25266 7437
rect 25314 7361 25386 7437
rect 25068 7243 25140 7319
rect 25194 7243 25266 7319
rect 25314 7243 25386 7319
rect 504 6985 576 7061
rect 626 6985 698 7061
rect 752 6985 824 7061
rect 504 6838 576 6914
rect 626 6838 698 6914
rect 752 6838 824 6914
rect 504 6701 576 6777
rect 626 6701 698 6777
rect 752 6701 824 6777
rect 26010 6216 26082 6292
rect 26136 6216 26208 6292
rect 26256 6216 26328 6292
rect 26010 6098 26082 6174
rect 26136 6098 26208 6174
rect 26256 6098 26328 6174
rect 504 5223 576 5299
rect 626 5223 698 5299
rect 752 5223 824 5299
rect 504 5076 576 5152
rect 626 5076 698 5152
rect 752 5076 824 5152
rect 504 4939 576 5015
rect 626 4939 698 5015
rect 752 4939 824 5015
rect 503 4563 575 4639
rect 629 4563 701 4639
rect 749 4563 821 4639
rect 503 4445 575 4521
rect 629 4445 701 4521
rect 749 4445 821 4521
rect 25068 4518 25140 4594
rect 25194 4518 25266 4594
rect 25314 4518 25386 4594
rect 25068 4400 25140 4476
rect 25194 4400 25266 4476
rect 25314 4400 25386 4476
rect 503 3452 575 3528
rect 629 3452 701 3528
rect 749 3452 821 3528
rect 503 3334 575 3410
rect 629 3334 701 3410
rect 749 3334 821 3410
rect 25068 3361 25140 3437
rect 25194 3361 25266 3437
rect 25314 3361 25386 3437
rect 25068 3243 25140 3319
rect 25194 3243 25266 3319
rect 25314 3243 25386 3319
rect 504 2985 576 3061
rect 626 2985 698 3061
rect 752 2985 824 3061
rect 504 2838 576 2914
rect 626 2838 698 2914
rect 752 2838 824 2914
rect 504 2701 576 2777
rect 626 2701 698 2777
rect 752 2701 824 2777
rect 26010 2204 26082 2280
rect 26136 2204 26208 2280
rect 26256 2204 26328 2280
rect 26010 2086 26082 2162
rect 26136 2086 26208 2162
rect 26256 2086 26328 2162
rect 504 1224 576 1300
rect 626 1224 698 1300
rect 752 1224 824 1300
rect 504 1077 576 1153
rect 626 1077 698 1153
rect 752 1077 824 1153
rect 504 940 576 1016
rect 626 940 698 1016
rect 752 940 824 1016
rect 503 629 575 705
rect 629 629 701 705
rect 749 629 821 705
rect 503 511 575 587
rect 629 511 701 587
rect 749 511 821 587
rect 25068 518 25140 594
rect 25194 518 25266 594
rect 25314 518 25386 594
rect 25068 400 25140 476
rect 25194 400 25266 476
rect 25314 400 25386 476
<< metal4 >>
rect 0 35741 400 64000
rect 0 35661 32 35741
rect 111 35661 156 35741
rect 236 35661 282 35741
rect 362 35661 400 35741
rect 0 35635 400 35661
rect 0 35555 32 35635
rect 111 35555 156 35635
rect 236 35555 282 35635
rect 362 35555 400 35635
rect 0 34587 400 35555
rect 0 34507 15 34587
rect 99 34507 129 34587
rect 213 34507 243 34587
rect 327 34507 400 34587
rect 0 33499 400 34507
rect 0 33419 15 33499
rect 99 33419 129 33499
rect 213 33419 243 33499
rect 327 33419 400 33499
rect 0 0 400 33419
rect 463 63477 863 64000
rect 25028 63517 25428 64000
rect 25026 63492 25428 63517
rect 463 63452 864 63477
rect 463 63376 503 63452
rect 575 63376 629 63452
rect 701 63376 749 63452
rect 821 63376 864 63452
rect 463 63334 864 63376
rect 463 63258 503 63334
rect 575 63258 629 63334
rect 701 63258 749 63334
rect 821 63258 864 63334
rect 25026 63416 25068 63492
rect 25140 63416 25194 63492
rect 25266 63416 25314 63492
rect 25386 63416 25428 63492
rect 25026 63374 25428 63416
rect 25026 63298 25068 63374
rect 25140 63298 25194 63374
rect 25266 63298 25314 63374
rect 25386 63298 25428 63374
rect 25026 63262 25428 63298
rect 463 63222 864 63258
rect 463 63060 863 63222
rect 463 62984 504 63060
rect 576 62984 626 63060
rect 698 62984 752 63060
rect 824 62984 863 63060
rect 463 62913 863 62984
rect 463 62837 504 62913
rect 576 62837 626 62913
rect 698 62837 752 62913
rect 824 62837 863 62913
rect 463 62776 863 62837
rect 463 62700 504 62776
rect 576 62700 626 62776
rect 698 62700 752 62776
rect 824 62700 863 62776
rect 463 61300 863 62700
rect 463 61224 504 61300
rect 576 61224 626 61300
rect 698 61224 752 61300
rect 824 61224 863 61300
rect 463 61153 863 61224
rect 463 61077 504 61153
rect 576 61077 626 61153
rect 698 61077 752 61153
rect 824 61077 863 61153
rect 463 61016 863 61077
rect 463 60940 504 61016
rect 576 60940 626 61016
rect 698 60940 752 61016
rect 824 60940 863 61016
rect 463 60804 863 60940
rect 463 60779 864 60804
rect 463 60703 503 60779
rect 575 60703 629 60779
rect 701 60703 749 60779
rect 821 60703 864 60779
rect 463 60661 864 60703
rect 463 60585 503 60661
rect 575 60585 629 60661
rect 701 60585 749 60661
rect 821 60585 864 60661
rect 463 60549 864 60585
rect 25028 60695 25428 63262
rect 25028 60619 25068 60695
rect 25140 60619 25194 60695
rect 25266 60619 25314 60695
rect 25386 60619 25428 60695
rect 25028 60577 25428 60619
rect 463 59475 863 60549
rect 25028 60501 25068 60577
rect 25140 60501 25194 60577
rect 25266 60501 25314 60577
rect 25386 60501 25428 60577
rect 25028 59517 25428 60501
rect 25026 59492 25428 59517
rect 463 59450 864 59475
rect 463 59374 503 59450
rect 575 59374 629 59450
rect 701 59374 749 59450
rect 821 59374 864 59450
rect 463 59332 864 59374
rect 463 59256 503 59332
rect 575 59256 629 59332
rect 701 59256 749 59332
rect 821 59256 864 59332
rect 25026 59416 25068 59492
rect 25140 59416 25194 59492
rect 25266 59416 25314 59492
rect 25386 59416 25428 59492
rect 25026 59374 25428 59416
rect 25026 59298 25068 59374
rect 25140 59298 25194 59374
rect 25266 59298 25314 59374
rect 25386 59298 25428 59374
rect 25026 59262 25428 59298
rect 463 59220 864 59256
rect 463 59060 863 59220
rect 463 58984 504 59060
rect 576 58984 626 59060
rect 698 58984 752 59060
rect 824 58984 863 59060
rect 463 58913 863 58984
rect 463 58837 504 58913
rect 576 58837 626 58913
rect 698 58837 752 58913
rect 824 58837 863 58913
rect 463 58776 863 58837
rect 463 58700 504 58776
rect 576 58700 626 58776
rect 698 58700 752 58776
rect 824 58700 863 58776
rect 463 57301 863 58700
rect 463 57225 504 57301
rect 576 57225 626 57301
rect 698 57225 752 57301
rect 824 57225 863 57301
rect 463 57154 863 57225
rect 463 57078 504 57154
rect 576 57078 626 57154
rect 698 57078 752 57154
rect 824 57078 863 57154
rect 463 57017 863 57078
rect 463 56941 504 57017
rect 576 56941 626 57017
rect 698 56941 752 57017
rect 824 56941 863 57017
rect 463 56735 863 56941
rect 463 56710 864 56735
rect 463 56634 503 56710
rect 575 56634 629 56710
rect 701 56634 749 56710
rect 821 56634 864 56710
rect 463 56592 864 56634
rect 463 56516 503 56592
rect 575 56516 629 56592
rect 701 56516 749 56592
rect 821 56516 864 56592
rect 463 56480 864 56516
rect 25028 56695 25428 59262
rect 25028 56619 25068 56695
rect 25140 56619 25194 56695
rect 25266 56619 25314 56695
rect 25386 56619 25428 56695
rect 25028 56577 25428 56619
rect 25028 56501 25068 56577
rect 25140 56501 25194 56577
rect 25266 56501 25314 56577
rect 25386 56501 25428 56577
rect 463 55557 863 56480
rect 463 55532 864 55557
rect 463 55456 503 55532
rect 575 55456 629 55532
rect 701 55456 749 55532
rect 821 55456 864 55532
rect 25028 55517 25428 56501
rect 463 55414 864 55456
rect 463 55338 503 55414
rect 575 55338 629 55414
rect 701 55338 749 55414
rect 821 55338 864 55414
rect 463 55302 864 55338
rect 25026 55492 25428 55517
rect 25026 55416 25068 55492
rect 25140 55416 25194 55492
rect 25266 55416 25314 55492
rect 25386 55416 25428 55492
rect 25026 55374 25428 55416
rect 463 55109 863 55302
rect 25026 55298 25068 55374
rect 25140 55298 25194 55374
rect 25266 55298 25314 55374
rect 25386 55298 25428 55374
rect 25026 55262 25428 55298
rect 463 55060 864 55109
rect 463 54984 504 55060
rect 576 54984 626 55060
rect 698 54984 752 55060
rect 824 54984 864 55060
rect 463 54913 864 54984
rect 463 54837 504 54913
rect 576 54837 626 54913
rect 698 54837 752 54913
rect 824 54837 864 54913
rect 463 54776 864 54837
rect 463 54700 504 54776
rect 576 54700 626 54776
rect 698 54700 752 54776
rect 824 54700 864 54776
rect 463 54650 864 54700
rect 463 53301 863 54650
rect 463 53225 504 53301
rect 576 53225 626 53301
rect 698 53225 752 53301
rect 824 53225 863 53301
rect 463 53154 863 53225
rect 463 53078 504 53154
rect 576 53078 626 53154
rect 698 53078 752 53154
rect 824 53078 863 53154
rect 463 53017 863 53078
rect 463 52941 504 53017
rect 576 52941 626 53017
rect 698 52941 752 53017
rect 824 52941 863 53017
rect 463 52709 863 52941
rect 463 52684 866 52709
rect 463 52608 503 52684
rect 575 52608 629 52684
rect 701 52608 749 52684
rect 821 52608 866 52684
rect 463 52566 866 52608
rect 463 52490 503 52566
rect 575 52490 629 52566
rect 701 52490 749 52566
rect 821 52490 866 52566
rect 463 52454 866 52490
rect 25028 52695 25428 55262
rect 25028 52619 25068 52695
rect 25140 52619 25194 52695
rect 25266 52619 25314 52695
rect 25386 52619 25428 52695
rect 25028 52577 25428 52619
rect 25028 52501 25068 52577
rect 25140 52501 25194 52577
rect 25266 52501 25314 52577
rect 25386 52501 25428 52577
rect 463 51506 863 52454
rect 25028 51571 25428 52501
rect 25027 51546 25428 51571
rect 463 51481 864 51506
rect 463 51405 503 51481
rect 575 51405 629 51481
rect 701 51405 749 51481
rect 821 51405 864 51481
rect 463 51363 864 51405
rect 463 51287 503 51363
rect 575 51287 629 51363
rect 701 51287 749 51363
rect 821 51287 864 51363
rect 25027 51470 25068 51546
rect 25140 51470 25194 51546
rect 25266 51470 25314 51546
rect 25386 51470 25428 51546
rect 25027 51428 25428 51470
rect 25027 51352 25068 51428
rect 25140 51352 25194 51428
rect 25266 51352 25314 51428
rect 25386 51352 25428 51428
rect 25027 51316 25428 51352
rect 463 51251 864 51287
rect 463 51109 863 51251
rect 463 51060 864 51109
rect 463 50984 504 51060
rect 576 50984 626 51060
rect 698 50984 752 51060
rect 824 50984 864 51060
rect 463 50913 864 50984
rect 463 50837 504 50913
rect 576 50837 626 50913
rect 698 50837 752 50913
rect 824 50837 864 50913
rect 463 50776 864 50837
rect 463 50700 504 50776
rect 576 50700 626 50776
rect 698 50700 752 50776
rect 824 50700 864 50776
rect 463 50650 864 50700
rect 463 49299 863 50650
rect 463 49223 504 49299
rect 576 49223 626 49299
rect 698 49223 752 49299
rect 824 49223 863 49299
rect 463 49152 863 49223
rect 463 49076 504 49152
rect 576 49076 626 49152
rect 698 49076 752 49152
rect 824 49076 863 49152
rect 463 49015 863 49076
rect 463 48939 504 49015
rect 576 48939 626 49015
rect 698 48939 752 49015
rect 824 48939 863 49015
rect 463 48729 863 48939
rect 463 48704 864 48729
rect 463 48628 503 48704
rect 575 48628 629 48704
rect 701 48628 749 48704
rect 821 48628 864 48704
rect 463 48586 864 48628
rect 463 48510 503 48586
rect 575 48510 629 48586
rect 701 48510 749 48586
rect 821 48510 864 48586
rect 463 48474 864 48510
rect 25028 48630 25428 51316
rect 25028 48554 25068 48630
rect 25140 48554 25194 48630
rect 25266 48554 25314 48630
rect 25386 48554 25428 48630
rect 25028 48512 25428 48554
rect 463 47522 863 48474
rect 25028 48436 25068 48512
rect 25140 48436 25194 48512
rect 25266 48436 25314 48512
rect 25386 48436 25428 48512
rect 463 47497 866 47522
rect 463 47421 503 47497
rect 575 47421 629 47497
rect 701 47421 749 47497
rect 821 47421 866 47497
rect 25028 47472 25428 48436
rect 463 47379 866 47421
rect 463 47303 503 47379
rect 575 47303 629 47379
rect 701 47303 749 47379
rect 821 47303 866 47379
rect 463 47267 866 47303
rect 25027 47447 25428 47472
rect 25027 47371 25068 47447
rect 25140 47371 25194 47447
rect 25266 47371 25314 47447
rect 25386 47371 25428 47447
rect 25027 47329 25428 47371
rect 463 47060 863 47267
rect 25027 47253 25068 47329
rect 25140 47253 25194 47329
rect 25266 47253 25314 47329
rect 25386 47253 25428 47329
rect 25027 47217 25428 47253
rect 463 46984 504 47060
rect 576 46984 626 47060
rect 698 46984 752 47060
rect 824 46984 863 47060
rect 463 46913 863 46984
rect 463 46837 504 46913
rect 576 46837 626 46913
rect 698 46837 752 46913
rect 824 46837 863 46913
rect 463 46776 863 46837
rect 463 46700 504 46776
rect 576 46700 626 46776
rect 698 46700 752 46776
rect 824 46700 863 46776
rect 463 45301 863 46700
rect 463 45225 504 45301
rect 576 45225 626 45301
rect 698 45225 752 45301
rect 824 45225 863 45301
rect 463 45154 863 45225
rect 463 45078 504 45154
rect 576 45078 626 45154
rect 698 45078 752 45154
rect 824 45078 863 45154
rect 463 45017 863 45078
rect 463 44941 504 45017
rect 576 44941 626 45017
rect 698 44941 752 45017
rect 824 44941 863 45017
rect 463 44756 863 44941
rect 463 44731 864 44756
rect 463 44655 503 44731
rect 575 44655 629 44731
rect 701 44655 749 44731
rect 821 44655 864 44731
rect 463 44613 864 44655
rect 463 44537 503 44613
rect 575 44537 629 44613
rect 701 44537 749 44613
rect 821 44537 864 44613
rect 463 44501 864 44537
rect 25028 44575 25428 47217
rect 463 43569 863 44501
rect 25028 44499 25068 44575
rect 25140 44499 25194 44575
rect 25266 44499 25314 44575
rect 25386 44499 25428 44575
rect 25028 44457 25428 44499
rect 25028 44381 25068 44457
rect 25140 44381 25194 44457
rect 25266 44381 25314 44457
rect 25386 44381 25428 44457
rect 463 43544 864 43569
rect 463 43468 503 43544
rect 575 43468 629 43544
rect 701 43468 749 43544
rect 821 43468 864 43544
rect 463 43426 864 43468
rect 463 43350 503 43426
rect 575 43350 629 43426
rect 701 43350 749 43426
rect 821 43350 864 43426
rect 463 43314 864 43350
rect 25028 43440 25428 44381
rect 25028 43364 25068 43440
rect 25140 43364 25194 43440
rect 25266 43364 25314 43440
rect 25386 43364 25428 43440
rect 25028 43322 25428 43364
rect 463 43060 863 43314
rect 463 42984 504 43060
rect 576 42984 626 43060
rect 698 42984 752 43060
rect 824 42984 863 43060
rect 463 42913 863 42984
rect 463 42837 504 42913
rect 576 42837 626 42913
rect 698 42837 752 42913
rect 824 42837 863 42913
rect 463 42776 863 42837
rect 463 42700 504 42776
rect 576 42700 626 42776
rect 698 42700 752 42776
rect 824 42700 863 42776
rect 463 41301 863 42700
rect 463 41225 504 41301
rect 576 41225 626 41301
rect 698 41225 752 41301
rect 824 41225 863 41301
rect 463 41154 863 41225
rect 463 41078 504 41154
rect 576 41078 626 41154
rect 698 41078 752 41154
rect 824 41078 863 41154
rect 463 41017 863 41078
rect 463 40941 504 41017
rect 576 40941 626 41017
rect 698 40941 752 41017
rect 824 40941 863 41017
rect 463 40747 863 40941
rect 25028 43246 25068 43322
rect 25140 43246 25194 43322
rect 25266 43246 25314 43322
rect 25386 43246 25428 43322
rect 463 40722 864 40747
rect 463 40646 503 40722
rect 575 40646 629 40722
rect 701 40646 749 40722
rect 821 40646 864 40722
rect 463 40604 864 40646
rect 463 40528 503 40604
rect 575 40528 629 40604
rect 701 40528 749 40604
rect 821 40528 864 40604
rect 463 40492 864 40528
rect 25028 40681 25428 43246
rect 25028 40605 25068 40681
rect 25140 40605 25194 40681
rect 25266 40605 25314 40681
rect 25386 40605 25428 40681
rect 25028 40563 25428 40605
rect 463 39594 863 40492
rect 25028 40487 25068 40563
rect 25140 40487 25194 40563
rect 25266 40487 25314 40563
rect 25386 40487 25428 40563
rect 463 39569 864 39594
rect 463 39493 503 39569
rect 575 39493 629 39569
rect 701 39493 749 39569
rect 821 39493 864 39569
rect 463 39451 864 39493
rect 463 39375 503 39451
rect 575 39375 629 39451
rect 701 39375 749 39451
rect 821 39375 864 39451
rect 463 39339 864 39375
rect 25028 39528 25428 40487
rect 25028 39452 25068 39528
rect 25140 39452 25194 39528
rect 25266 39452 25314 39528
rect 25386 39452 25428 39528
rect 25028 39410 25428 39452
rect 463 39060 863 39339
rect 463 38984 504 39060
rect 576 38984 626 39060
rect 698 38984 752 39060
rect 824 38984 863 39060
rect 463 38913 863 38984
rect 463 38837 504 38913
rect 576 38837 626 38913
rect 698 38837 752 38913
rect 824 38837 863 38913
rect 463 38776 863 38837
rect 463 38700 504 38776
rect 576 38700 626 38776
rect 698 38700 752 38776
rect 824 38700 863 38776
rect 463 37300 863 38700
rect 463 37224 504 37300
rect 576 37224 626 37300
rect 698 37224 752 37300
rect 824 37224 863 37300
rect 463 37153 863 37224
rect 463 37077 504 37153
rect 576 37077 626 37153
rect 698 37077 752 37153
rect 824 37077 863 37153
rect 463 37016 863 37077
rect 463 36940 504 37016
rect 576 36940 626 37016
rect 698 36940 752 37016
rect 824 36940 863 37016
rect 463 36509 863 36940
rect 463 36433 503 36509
rect 575 36433 629 36509
rect 701 36433 749 36509
rect 821 36433 863 36509
rect 463 36391 863 36433
rect 463 36315 503 36391
rect 575 36315 629 36391
rect 701 36315 749 36391
rect 821 36315 863 36391
rect 463 35131 863 36315
rect 25028 39334 25068 39410
rect 25140 39334 25194 39410
rect 25266 39334 25314 39410
rect 25386 39334 25428 39410
rect 25028 36412 25428 39334
rect 25028 36336 25068 36412
rect 25140 36336 25194 36412
rect 25266 36336 25314 36412
rect 25386 36336 25428 36412
rect 25028 36294 25428 36336
rect 25028 36218 25068 36294
rect 25140 36218 25194 36294
rect 25266 36218 25314 36294
rect 25386 36218 25428 36294
rect 2306 35942 2467 36000
rect 2246 35925 2467 35942
rect 2246 35861 2249 35925
rect 2313 35861 2337 35925
rect 2401 35861 2467 35925
rect 2246 35845 2467 35861
rect 2246 35781 2249 35845
rect 2313 35781 2337 35845
rect 2401 35781 2467 35845
rect 2246 35775 2467 35781
rect 4190 35905 4348 36000
rect 4190 35841 4192 35905
rect 4256 35841 4280 35905
rect 4344 35841 4348 35905
rect 4190 35825 4348 35841
rect 4190 35761 4192 35825
rect 4256 35761 4280 35825
rect 4344 35761 4348 35825
rect 4190 35754 4348 35761
rect 463 35051 478 35131
rect 562 35051 592 35131
rect 676 35051 706 35131
rect 790 35051 863 35131
rect 463 34043 863 35051
rect 25028 34998 25428 36218
rect 24527 34972 25428 34998
rect 24527 34892 25061 34972
rect 25141 34892 25186 34972
rect 25266 34892 25311 34972
rect 25391 34892 25428 34972
rect 24527 34852 25428 34892
rect 24527 34772 25060 34852
rect 25140 34772 25185 34852
rect 25265 34772 25310 34852
rect 25390 34772 25428 34852
rect 24527 34743 25428 34772
rect 463 33963 478 34043
rect 562 33963 592 34043
rect 676 33963 706 34043
rect 790 33963 863 34043
rect 463 32955 863 33963
rect 25028 34392 25428 34743
rect 25028 34316 25069 34392
rect 25141 34316 25191 34392
rect 25263 34316 25317 34392
rect 25389 34316 25428 34392
rect 25028 34245 25428 34316
rect 25028 34169 25069 34245
rect 25141 34169 25191 34245
rect 25263 34169 25317 34245
rect 25389 34169 25428 34245
rect 25028 34108 25428 34169
rect 25028 34032 25069 34108
rect 25141 34032 25191 34108
rect 25263 34032 25317 34108
rect 25389 34032 25428 34108
rect 24527 33476 24927 33502
rect 24527 33396 24560 33476
rect 24640 33396 24685 33476
rect 24765 33396 24810 33476
rect 24890 33396 24927 33476
rect 24527 33356 24927 33396
rect 24527 33276 24559 33356
rect 24639 33276 24684 33356
rect 24764 33276 24809 33356
rect 24889 33276 24927 33356
rect 24527 33247 24927 33276
rect 463 32875 478 32955
rect 562 32875 592 32955
rect 676 32875 706 32955
rect 790 32875 863 32955
rect 463 28360 863 32875
rect 25028 32632 25428 34032
rect 25028 32556 25069 32632
rect 25141 32556 25191 32632
rect 25263 32556 25317 32632
rect 25389 32556 25428 32632
rect 25028 32485 25428 32556
rect 3093 32463 3338 32476
rect 3093 32399 3136 32463
rect 3200 32399 3224 32463
rect 3288 32399 3338 32463
rect 463 28302 866 28360
rect 463 28226 503 28302
rect 575 28226 629 28302
rect 701 28226 749 28302
rect 821 28226 866 28302
rect 463 28184 866 28226
rect 463 28108 503 28184
rect 575 28108 629 28184
rect 701 28108 749 28184
rect 821 28108 866 28184
rect 463 28072 866 28108
rect 463 28000 863 28072
rect 3093 28000 3338 32399
rect 25028 32409 25069 32485
rect 25141 32409 25191 32485
rect 25263 32409 25317 32485
rect 25389 32409 25428 32485
rect 25028 32348 25428 32409
rect 25028 32272 25069 32348
rect 25141 32272 25191 32348
rect 25263 32272 25317 32348
rect 25389 32272 25428 32348
rect 25028 31943 25428 32272
rect 24514 31917 25428 31943
rect 24514 31837 25060 31917
rect 25140 31837 25185 31917
rect 25265 31837 25310 31917
rect 25390 31837 25428 31917
rect 24514 31797 25428 31837
rect 24514 31717 25059 31797
rect 25139 31717 25184 31797
rect 25264 31717 25309 31797
rect 25389 31717 25428 31797
rect 24514 31688 25428 31717
rect 25028 28360 25428 31688
rect 25025 28302 25428 28360
rect 25025 28226 25068 28302
rect 25140 28226 25194 28302
rect 25266 28226 25314 28302
rect 25386 28226 25428 28302
rect 25025 28184 25428 28226
rect 25025 28108 25068 28184
rect 25140 28108 25194 28184
rect 25266 28108 25314 28184
rect 25386 28108 25428 28184
rect 25025 28072 25428 28108
rect 463 27760 946 28000
rect 463 27520 863 27760
rect 463 27444 503 27520
rect 575 27444 629 27520
rect 701 27444 749 27520
rect 821 27444 863 27520
rect 463 27402 863 27444
rect 463 27326 503 27402
rect 575 27326 629 27402
rect 701 27326 749 27402
rect 821 27326 863 27402
rect 463 27061 863 27326
rect 25028 27520 25428 28072
rect 25028 27444 25068 27520
rect 25140 27444 25194 27520
rect 25266 27444 25314 27520
rect 25386 27444 25428 27520
rect 25028 27402 25428 27444
rect 25028 27326 25068 27402
rect 25140 27326 25194 27402
rect 25266 27326 25314 27402
rect 25386 27326 25428 27402
rect 953 27120 1155 27121
rect 463 26985 504 27061
rect 576 26985 626 27061
rect 698 26985 752 27061
rect 824 26985 863 27061
rect 463 26914 863 26985
rect 463 26838 504 26914
rect 576 26838 626 26914
rect 698 26838 752 26914
rect 824 26838 863 26914
rect 463 26777 863 26838
rect 463 26701 504 26777
rect 576 26701 626 26777
rect 698 26701 752 26777
rect 824 26701 863 26777
rect 463 25294 863 26701
rect 463 25218 504 25294
rect 576 25218 626 25294
rect 698 25218 752 25294
rect 824 25218 863 25294
rect 463 25147 863 25218
rect 463 25071 504 25147
rect 576 25071 626 25147
rect 698 25071 752 25147
rect 824 25071 863 25147
rect 463 25010 863 25071
rect 463 24934 504 25010
rect 576 24934 626 25010
rect 698 24934 752 25010
rect 824 24934 863 25010
rect 463 24885 863 24934
rect 463 24668 862 24885
rect 944 24681 946 24880
rect 463 24608 863 24668
rect 463 24532 503 24608
rect 575 24532 629 24608
rect 701 24532 749 24608
rect 821 24532 863 24608
rect 463 24490 863 24532
rect 463 24414 503 24490
rect 575 24414 629 24490
rect 701 24414 749 24490
rect 821 24414 863 24490
rect 463 24238 863 24414
rect 25028 24559 25428 27326
rect 25028 24483 25068 24559
rect 25140 24483 25194 24559
rect 25266 24483 25314 24559
rect 25386 24483 25428 24559
rect 25028 24441 25428 24483
rect 25028 24365 25068 24441
rect 25140 24365 25194 24441
rect 25266 24365 25314 24441
rect 25386 24365 25428 24441
rect 463 24209 946 24238
rect 25028 24232 25428 24365
rect 462 23979 946 24209
rect 463 23760 946 23979
rect 24946 23766 25428 24232
rect 463 23604 863 23760
rect 463 23528 503 23604
rect 575 23528 629 23604
rect 701 23528 749 23604
rect 821 23528 863 23604
rect 463 23486 863 23528
rect 463 23410 503 23486
rect 575 23410 629 23486
rect 701 23410 749 23486
rect 821 23410 863 23486
rect 25028 23467 25428 23766
rect 463 23060 863 23410
rect 25027 23442 25428 23467
rect 25027 23366 25068 23442
rect 25140 23366 25194 23442
rect 25266 23366 25314 23442
rect 25386 23366 25428 23442
rect 25027 23324 25428 23366
rect 25027 23248 25068 23324
rect 25140 23248 25194 23324
rect 25266 23248 25314 23324
rect 25386 23248 25428 23324
rect 25027 23212 25428 23248
rect 463 22984 504 23060
rect 576 22984 626 23060
rect 698 22984 752 23060
rect 824 22984 863 23060
rect 463 22913 863 22984
rect 463 22837 504 22913
rect 576 22837 626 22913
rect 698 22837 752 22913
rect 824 22837 863 22913
rect 463 22776 863 22837
rect 463 22700 504 22776
rect 576 22700 626 22776
rect 698 22700 752 22776
rect 824 22700 863 22776
rect 463 21300 863 22700
rect 463 21224 504 21300
rect 576 21224 626 21300
rect 698 21224 752 21300
rect 824 21224 863 21300
rect 463 21153 863 21224
rect 463 21077 504 21153
rect 576 21077 626 21153
rect 698 21077 752 21153
rect 824 21077 863 21153
rect 463 21016 863 21077
rect 463 20940 504 21016
rect 576 20940 626 21016
rect 698 20940 752 21016
rect 824 20940 863 21016
rect 463 20651 863 20940
rect 463 20626 864 20651
rect 463 20550 503 20626
rect 575 20550 629 20626
rect 701 20550 749 20626
rect 821 20550 864 20626
rect 463 20508 864 20550
rect 463 20432 503 20508
rect 575 20432 629 20508
rect 701 20432 749 20508
rect 821 20432 864 20508
rect 463 20396 864 20432
rect 25028 20599 25428 23212
rect 25028 20523 25068 20599
rect 25140 20523 25194 20599
rect 25266 20523 25314 20599
rect 25386 20523 25428 20599
rect 25028 20481 25428 20523
rect 25028 20405 25068 20481
rect 25140 20405 25194 20481
rect 25266 20405 25314 20481
rect 25386 20405 25428 20481
rect 463 20239 863 20396
rect 463 19759 947 20239
rect 25028 20232 25428 20405
rect 24946 19767 25428 20232
rect 463 19569 863 19759
rect 463 19544 864 19569
rect 463 19468 503 19544
rect 575 19468 629 19544
rect 701 19468 749 19544
rect 821 19468 864 19544
rect 463 19426 864 19468
rect 463 19350 503 19426
rect 575 19350 629 19426
rect 701 19350 749 19426
rect 821 19350 864 19426
rect 463 19314 864 19350
rect 25028 19424 25428 19767
rect 25028 19348 25068 19424
rect 25140 19348 25194 19424
rect 25266 19348 25314 19424
rect 25386 19348 25428 19424
rect 463 19060 863 19314
rect 463 18984 504 19060
rect 576 18984 626 19060
rect 698 18984 752 19060
rect 824 18984 863 19060
rect 463 18913 863 18984
rect 463 18837 504 18913
rect 576 18837 626 18913
rect 698 18837 752 18913
rect 824 18837 863 18913
rect 463 18776 863 18837
rect 463 18700 504 18776
rect 576 18700 626 18776
rect 698 18700 752 18776
rect 824 18700 863 18776
rect 463 17301 863 18700
rect 463 17225 504 17301
rect 576 17225 626 17301
rect 698 17225 752 17301
rect 824 17225 863 17301
rect 463 17154 863 17225
rect 463 17078 504 17154
rect 576 17078 626 17154
rect 698 17078 752 17154
rect 824 17078 863 17154
rect 463 17017 863 17078
rect 463 16941 504 17017
rect 576 16941 626 17017
rect 698 16941 752 17017
rect 824 16941 863 17017
rect 463 16694 863 16941
rect 25028 19306 25428 19348
rect 25028 19230 25068 19306
rect 25140 19230 25194 19306
rect 25266 19230 25314 19306
rect 25386 19230 25428 19306
rect 463 16669 864 16694
rect 463 16593 503 16669
rect 575 16593 629 16669
rect 701 16593 749 16669
rect 821 16593 864 16669
rect 25028 16608 25428 19230
rect 463 16551 864 16593
rect 463 16475 503 16551
rect 575 16475 629 16551
rect 701 16475 749 16551
rect 821 16475 864 16551
rect 463 16439 864 16475
rect 25027 16583 25428 16608
rect 25027 16507 25068 16583
rect 25140 16507 25194 16583
rect 25266 16507 25314 16583
rect 25386 16507 25428 16583
rect 25027 16465 25428 16507
rect 463 16240 863 16439
rect 25027 16389 25068 16465
rect 25140 16389 25194 16465
rect 25266 16389 25314 16465
rect 25386 16389 25428 16465
rect 25027 16353 25428 16389
rect 463 15760 946 16240
rect 25028 16233 25428 16353
rect 24946 15768 25428 16233
rect 463 15593 863 15760
rect 463 15568 864 15593
rect 463 15492 503 15568
rect 575 15492 629 15568
rect 701 15492 749 15568
rect 821 15492 864 15568
rect 463 15450 864 15492
rect 463 15374 503 15450
rect 575 15374 629 15450
rect 701 15374 749 15450
rect 821 15374 864 15450
rect 25028 15437 25428 15768
rect 463 15338 864 15374
rect 25027 15412 25428 15437
rect 463 15060 863 15338
rect 25027 15336 25068 15412
rect 25140 15336 25194 15412
rect 25266 15336 25314 15412
rect 25386 15336 25428 15412
rect 25027 15294 25428 15336
rect 25027 15218 25068 15294
rect 25140 15218 25194 15294
rect 25266 15218 25314 15294
rect 25386 15218 25428 15294
rect 25027 15182 25428 15218
rect 463 14984 504 15060
rect 576 14984 626 15060
rect 698 14984 752 15060
rect 824 14984 863 15060
rect 463 14913 863 14984
rect 463 14837 504 14913
rect 576 14837 626 14913
rect 698 14837 752 14913
rect 824 14837 863 14913
rect 463 14776 863 14837
rect 463 14700 504 14776
rect 576 14700 626 14776
rect 698 14700 752 14776
rect 824 14700 863 14776
rect 463 13300 863 14700
rect 463 13224 504 13300
rect 576 13224 626 13300
rect 698 13224 752 13300
rect 824 13224 863 13300
rect 463 13153 863 13224
rect 463 13077 504 13153
rect 576 13077 626 13153
rect 698 13077 752 13153
rect 824 13077 863 13153
rect 463 13016 863 13077
rect 463 12940 504 13016
rect 576 12940 626 13016
rect 698 12940 752 13016
rect 824 12940 863 13016
rect 463 12727 863 12940
rect 463 12702 865 12727
rect 463 12626 503 12702
rect 575 12626 629 12702
rect 701 12626 749 12702
rect 821 12626 865 12702
rect 25028 12676 25428 15182
rect 463 12584 865 12626
rect 463 12508 503 12584
rect 575 12508 629 12584
rect 701 12508 749 12584
rect 821 12508 865 12584
rect 463 12472 865 12508
rect 25027 12651 25428 12676
rect 25027 12575 25068 12651
rect 25140 12575 25194 12651
rect 25266 12575 25314 12651
rect 25386 12575 25428 12651
rect 25027 12533 25428 12575
rect 463 12239 863 12472
rect 25027 12457 25068 12533
rect 25140 12457 25194 12533
rect 25266 12457 25314 12533
rect 25386 12457 25428 12533
rect 25027 12421 25428 12457
rect 463 11759 946 12239
rect 25028 12232 25428 12421
rect 24946 11766 25428 12232
rect 463 11511 863 11759
rect 463 11486 866 11511
rect 463 11410 503 11486
rect 575 11410 629 11486
rect 701 11410 749 11486
rect 821 11410 866 11486
rect 25028 11462 25428 11766
rect 463 11368 866 11410
rect 463 11292 503 11368
rect 575 11292 629 11368
rect 701 11292 749 11368
rect 821 11292 866 11368
rect 463 11256 866 11292
rect 25027 11437 25428 11462
rect 25027 11361 25068 11437
rect 25140 11361 25194 11437
rect 25266 11361 25314 11437
rect 25386 11361 25428 11437
rect 25027 11319 25428 11361
rect 463 11060 863 11256
rect 25027 11243 25068 11319
rect 25140 11243 25194 11319
rect 25266 11243 25314 11319
rect 25386 11243 25428 11319
rect 25027 11207 25428 11243
rect 463 10984 504 11060
rect 576 10984 626 11060
rect 698 10984 752 11060
rect 824 10984 863 11060
rect 463 10913 863 10984
rect 463 10837 504 10913
rect 576 10837 626 10913
rect 698 10837 752 10913
rect 824 10837 863 10913
rect 463 10776 863 10837
rect 463 10700 504 10776
rect 576 10700 626 10776
rect 698 10700 752 10776
rect 824 10700 863 10776
rect 463 9300 863 10700
rect 463 9224 504 9300
rect 576 9224 626 9300
rect 698 9224 752 9300
rect 824 9224 863 9300
rect 463 9153 863 9224
rect 463 9077 504 9153
rect 576 9077 626 9153
rect 698 9077 752 9153
rect 824 9077 863 9153
rect 463 9016 863 9077
rect 463 8940 504 9016
rect 576 8940 626 9016
rect 698 8940 752 9016
rect 824 8940 863 9016
rect 463 8646 863 8940
rect 463 8621 864 8646
rect 463 8545 503 8621
rect 575 8545 629 8621
rect 701 8545 749 8621
rect 821 8545 864 8621
rect 463 8503 864 8545
rect 463 8427 503 8503
rect 575 8427 629 8503
rect 701 8427 749 8503
rect 821 8427 864 8503
rect 463 8391 864 8427
rect 25028 8594 25428 11207
rect 25028 8518 25068 8594
rect 25140 8518 25194 8594
rect 25266 8518 25314 8594
rect 25386 8518 25428 8594
rect 25028 8476 25428 8518
rect 25028 8400 25068 8476
rect 25140 8400 25194 8476
rect 25266 8400 25314 8476
rect 25386 8400 25428 8476
rect 463 8238 863 8391
rect 463 7998 947 8238
rect 25028 8233 25428 8400
rect 463 7758 946 7998
rect 24946 7766 25428 8233
rect 463 7524 863 7758
rect 463 7499 864 7524
rect 463 7423 503 7499
rect 575 7423 629 7499
rect 701 7423 749 7499
rect 821 7423 864 7499
rect 25028 7462 25428 7766
rect 463 7381 864 7423
rect 463 7305 503 7381
rect 575 7305 629 7381
rect 701 7305 749 7381
rect 821 7305 864 7381
rect 463 7269 864 7305
rect 25027 7437 25428 7462
rect 25027 7361 25068 7437
rect 25140 7361 25194 7437
rect 25266 7361 25314 7437
rect 25386 7361 25428 7437
rect 25027 7319 25428 7361
rect 463 7061 863 7269
rect 25027 7243 25068 7319
rect 25140 7243 25194 7319
rect 25266 7243 25314 7319
rect 25386 7243 25428 7319
rect 25027 7207 25428 7243
rect 463 6985 504 7061
rect 576 6985 626 7061
rect 698 6985 752 7061
rect 824 6985 863 7061
rect 463 6914 863 6985
rect 463 6838 504 6914
rect 576 6838 626 6914
rect 698 6838 752 6914
rect 824 6838 863 6914
rect 463 6777 863 6838
rect 463 6701 504 6777
rect 576 6701 626 6777
rect 698 6701 752 6777
rect 824 6701 863 6777
rect 463 5299 863 6701
rect 463 5223 504 5299
rect 576 5223 626 5299
rect 698 5223 752 5299
rect 824 5223 863 5299
rect 463 5152 863 5223
rect 463 5076 504 5152
rect 576 5076 626 5152
rect 698 5076 752 5152
rect 824 5076 863 5152
rect 463 5015 863 5076
rect 463 4939 504 5015
rect 576 4939 626 5015
rect 698 4939 752 5015
rect 824 4939 863 5015
rect 463 4639 863 4939
rect 463 4563 503 4639
rect 575 4563 629 4639
rect 701 4563 749 4639
rect 821 4563 863 4639
rect 463 4521 863 4563
rect 463 4445 503 4521
rect 575 4445 629 4521
rect 701 4445 749 4521
rect 821 4445 863 4521
rect 463 4238 863 4445
rect 25028 4594 25428 7207
rect 25028 4518 25068 4594
rect 25140 4518 25194 4594
rect 25266 4518 25314 4594
rect 25386 4518 25428 4594
rect 25028 4476 25428 4518
rect 25028 4400 25068 4476
rect 25140 4400 25194 4476
rect 25266 4400 25314 4476
rect 25386 4400 25428 4476
rect 463 4000 946 4238
rect 25028 4233 25428 4400
rect 463 3760 947 4000
rect 24946 3766 25428 4233
rect 463 3528 863 3760
rect 463 3452 503 3528
rect 575 3452 629 3528
rect 701 3452 749 3528
rect 821 3452 863 3528
rect 25028 3462 25428 3766
rect 463 3410 863 3452
rect 463 3334 503 3410
rect 575 3334 629 3410
rect 701 3334 749 3410
rect 821 3334 863 3410
rect 463 3061 863 3334
rect 25027 3437 25428 3462
rect 25027 3361 25068 3437
rect 25140 3361 25194 3437
rect 25266 3361 25314 3437
rect 25386 3361 25428 3437
rect 25027 3319 25428 3361
rect 25027 3243 25068 3319
rect 25140 3243 25194 3319
rect 25266 3243 25314 3319
rect 25386 3243 25428 3319
rect 25027 3207 25428 3243
rect 463 2985 504 3061
rect 576 2985 626 3061
rect 698 2985 752 3061
rect 824 2985 863 3061
rect 463 2914 863 2985
rect 463 2838 504 2914
rect 576 2838 626 2914
rect 698 2838 752 2914
rect 824 2838 863 2914
rect 463 2777 863 2838
rect 463 2701 504 2777
rect 576 2701 626 2777
rect 698 2701 752 2777
rect 824 2701 863 2777
rect 463 1300 863 2701
rect 463 1224 504 1300
rect 576 1224 626 1300
rect 698 1224 752 1300
rect 824 1224 863 1300
rect 463 1153 863 1224
rect 463 1077 504 1153
rect 576 1077 626 1153
rect 698 1077 752 1153
rect 824 1077 863 1153
rect 463 1016 863 1077
rect 463 940 504 1016
rect 576 940 626 1016
rect 698 940 752 1016
rect 824 940 863 1016
rect 463 730 863 940
rect 463 705 865 730
rect 463 629 503 705
rect 575 629 629 705
rect 701 629 749 705
rect 821 629 865 705
rect 463 587 865 629
rect 463 511 503 587
rect 575 511 629 587
rect 701 511 749 587
rect 821 511 865 587
rect 463 475 865 511
rect 25028 594 25428 3207
rect 25028 518 25068 594
rect 25140 518 25194 594
rect 25266 518 25314 594
rect 25386 518 25428 594
rect 25028 476 25428 518
rect 463 239 863 475
rect 25028 400 25068 476
rect 25140 400 25194 476
rect 25266 400 25314 476
rect 25386 400 25428 476
rect 463 0 947 239
rect 25028 233 25428 400
rect 24946 0 25428 233
rect 25502 35726 25902 64000
rect 25502 35646 25535 35726
rect 25615 35646 25660 35726
rect 25740 35646 25785 35726
rect 25865 35646 25902 35726
rect 25502 35606 25902 35646
rect 25502 35526 25534 35606
rect 25614 35526 25659 35606
rect 25739 35526 25784 35606
rect 25864 35526 25902 35606
rect 25502 33476 25902 35526
rect 25502 33396 25535 33476
rect 25615 33396 25660 33476
rect 25740 33396 25785 33476
rect 25865 33396 25902 33476
rect 25502 33356 25902 33396
rect 25502 33276 25534 33356
rect 25614 33276 25659 33356
rect 25739 33276 25784 33356
rect 25864 33276 25902 33356
rect 25502 0 25902 33276
rect 25970 62071 26370 64000
rect 25970 61995 26010 62071
rect 26082 61995 26136 62071
rect 26208 61995 26256 62071
rect 26328 61995 26370 62071
rect 25970 61953 26370 61995
rect 25970 61877 26010 61953
rect 26082 61877 26136 61953
rect 26208 61877 26256 61953
rect 26328 61877 26370 61953
rect 25970 58058 26370 61877
rect 25970 57982 26010 58058
rect 26082 57982 26136 58058
rect 26208 57982 26256 58058
rect 26328 57982 26370 58058
rect 25970 57940 26370 57982
rect 25970 57864 26010 57940
rect 26082 57864 26136 57940
rect 26208 57864 26256 57940
rect 26328 57864 26370 57940
rect 25970 54057 26370 57864
rect 25970 53981 26010 54057
rect 26082 53981 26136 54057
rect 26208 53981 26256 54057
rect 26328 53981 26370 54057
rect 25970 53939 26370 53981
rect 25970 53863 26010 53939
rect 26082 53863 26136 53939
rect 26208 53863 26256 53939
rect 26328 53863 26370 53939
rect 25970 50096 26370 53863
rect 25970 50020 26010 50096
rect 26082 50020 26136 50096
rect 26208 50020 26256 50096
rect 26328 50020 26370 50096
rect 25970 49978 26370 50020
rect 25970 49902 26010 49978
rect 26082 49902 26136 49978
rect 26208 49902 26256 49978
rect 26328 49902 26370 49978
rect 25970 46079 26370 49902
rect 25970 46003 26010 46079
rect 26082 46003 26136 46079
rect 26208 46003 26256 46079
rect 26328 46003 26370 46079
rect 25970 45961 26370 46003
rect 25970 45885 26010 45961
rect 26082 45885 26136 45961
rect 26208 45885 26256 45961
rect 26328 45885 26370 45961
rect 25970 42158 26370 45885
rect 25970 42082 26010 42158
rect 26082 42082 26136 42158
rect 26208 42082 26256 42158
rect 26328 42082 26370 42158
rect 25970 42040 26370 42082
rect 25970 41964 26010 42040
rect 26082 41964 26136 42040
rect 26208 41964 26256 42040
rect 26328 41964 26370 42040
rect 25970 37900 26370 41964
rect 25970 37824 26010 37900
rect 26082 37824 26136 37900
rect 26208 37824 26256 37900
rect 26328 37824 26370 37900
rect 25970 37782 26370 37824
rect 25970 37706 26010 37782
rect 26082 37706 26136 37782
rect 26208 37706 26256 37782
rect 26328 37706 26370 37782
rect 25970 26130 26370 37706
rect 25970 26054 26010 26130
rect 26082 26054 26136 26130
rect 26208 26054 26256 26130
rect 26328 26054 26370 26130
rect 25970 26012 26370 26054
rect 25970 25936 26010 26012
rect 26082 25936 26136 26012
rect 26208 25936 26256 26012
rect 26328 25936 26370 26012
rect 25970 21971 26370 25936
rect 25970 21895 26010 21971
rect 26082 21895 26136 21971
rect 26208 21895 26256 21971
rect 26328 21895 26370 21971
rect 25970 21853 26370 21895
rect 25970 21777 26010 21853
rect 26082 21777 26136 21853
rect 26208 21777 26256 21853
rect 26328 21777 26370 21853
rect 25970 18181 26370 21777
rect 25970 18105 26010 18181
rect 26082 18105 26136 18181
rect 26208 18105 26256 18181
rect 26328 18105 26370 18181
rect 25970 18063 26370 18105
rect 25970 17987 26010 18063
rect 26082 17987 26136 18063
rect 26208 17987 26256 18063
rect 26328 17987 26370 18063
rect 25970 14074 26370 17987
rect 25970 13998 26010 14074
rect 26082 13998 26136 14074
rect 26208 13998 26256 14074
rect 26328 13998 26370 14074
rect 25970 13956 26370 13998
rect 25970 13880 26010 13956
rect 26082 13880 26136 13956
rect 26208 13880 26256 13956
rect 26328 13880 26370 13956
rect 25970 10256 26370 13880
rect 25970 10180 26010 10256
rect 26082 10180 26136 10256
rect 26208 10180 26256 10256
rect 26328 10180 26370 10256
rect 25970 10138 26370 10180
rect 25970 10062 26010 10138
rect 26082 10062 26136 10138
rect 26208 10062 26256 10138
rect 26328 10062 26370 10138
rect 25970 6292 26370 10062
rect 25970 6216 26010 6292
rect 26082 6216 26136 6292
rect 26208 6216 26256 6292
rect 26328 6216 26370 6292
rect 25970 6174 26370 6216
rect 25970 6098 26010 6174
rect 26082 6098 26136 6174
rect 26208 6098 26256 6174
rect 26328 6098 26370 6174
rect 25970 2280 26370 6098
rect 25970 2204 26010 2280
rect 26082 2204 26136 2280
rect 26208 2204 26256 2280
rect 26328 2204 26370 2280
rect 25970 2162 26370 2204
rect 25970 2086 26010 2162
rect 26082 2086 26136 2162
rect 26208 2086 26256 2162
rect 26328 2086 26370 2162
rect 25970 0 26370 2086
use adc_noise_decoup_cell1  adc_noise_decoup_cell1_0
array 0 3 4000 0 0 4000
timestamp 1663849571
transform 1 0 8527 0 1 31332
box 0 0 4000 4000
use adc_noise_decoup_cell1  adc_noise_decoup_cell1_1
array 0 5 4000 0 6 4000
timestamp 1663849571
transform 1 0 946 0 1 0
box 0 0 4000 4000
use adc_noise_decoup_cell1  adc_noise_decoup_cell1_3
array 0 5 4000 0 6 4000
timestamp 1663849571
transform 1 0 946 0 1 36000
box 0 0 4000 4000
use sky130_fd_pr__nfet_01v8_8PFHMD  sky130_fd_pr__nfet_01v8_8PFHMD_0
timestamp 1663599054
transform 1 0 3156 0 1 35031
box -187 -76 187 76
use sky130_fd_pr__nfet_01v8_8PFHMD  sky130_fd_pr__nfet_01v8_8PFHMD_1
timestamp 1663599054
transform 1 0 2510 0 1 35031
box -187 -76 187 76
use sky130_fd_pr__nfet_01v8_8PFHMD  sky130_fd_pr__nfet_01v8_8PFHMD_2
timestamp 1663599054
transform 1 0 3212 0 1 32975
box -187 -76 187 76
use sky130_fd_pr__nfet_01v8_8PFHMD  sky130_fd_pr__nfet_01v8_8PFHMD_3
timestamp 1663599054
transform 1 0 2580 0 1 32975
box -187 -76 187 76
use sky130_fd_pr__nfet_01v8_8PFHMD  sky130_fd_pr__nfet_01v8_8PFHMD_4
timestamp 1663599054
transform 1 0 1881 0 -1 35031
box -187 -76 187 76
use sky130_fd_pr__pfet_01v8_K25L97  sky130_fd_pr__pfet_01v8_K25L97_0
timestamp 1663599042
transform 1 0 3156 0 1 34747
box -323 -162 323 162
use sky130_fd_pr__pfet_01v8_K25L97  sky130_fd_pr__pfet_01v8_K25L97_1
timestamp 1663599042
transform 1 0 2510 0 1 34747
box -323 -162 323 162
use sky130_fd_pr__pfet_01v8_K25L97  sky130_fd_pr__pfet_01v8_K25L97_2
timestamp 1663599042
transform 1 0 3212 0 1 33259
box -323 -162 323 162
use sky130_fd_pr__pfet_01v8_K25L97  sky130_fd_pr__pfet_01v8_K25L97_3
timestamp 1663599042
transform 1 0 2580 0 1 33259
box -323 -162 323 162
use sky130_fd_pr__pfet_01v8_K25L97  sky130_fd_pr__pfet_01v8_K25L97_4
timestamp 1663599042
transform 1 0 1881 0 -1 34747
box -323 -162 323 162
use sky130_fd_sc_hd__buf_4  sky130_fd_sc_hd__buf_4_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform -1 0 4769 0 -1 35091
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  sky130_fd_sc_hd__buf_4_1
timestamp 1662439860
transform -1 0 4217 0 -1 35091
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  sky130_fd_sc_hd__buf_4_2
timestamp 1662439860
transform -1 0 4769 0 1 32915
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  sky130_fd_sc_hd__buf_4_3
timestamp 1662439860
transform -1 0 4217 0 1 32915
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s6s_1  sky130_fd_sc_hd__dlymetal6s6s_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 2561 0 1 34003
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s6s_1  sky130_fd_sc_hd__dlymetal6s6s_1_1
timestamp 1662439860
transform 1 0 2561 0 -1 34003
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s6s_1  sky130_fd_sc_hd__dlymetal6s6s_1_2
timestamp 1662439860
transform 1 0 3481 0 1 34003
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s6s_1  sky130_fd_sc_hd__dlymetal6s6s_1_3
timestamp 1662439860
transform 1 0 4401 0 1 34003
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s6s_1  sky130_fd_sc_hd__dlymetal6s6s_1_4
timestamp 1662439860
transform 1 0 3481 0 -1 34003
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s6s_1  sky130_fd_sc_hd__dlymetal6s6s_1_5
timestamp 1662439860
transform 1 0 4401 0 -1 34003
box -38 -48 958 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform -1 0 5321 0 -1 35091
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_1
timestamp 1662439860
transform -1 0 5321 0 1 32915
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_2
timestamp 1662439860
transform -1 0 5045 0 -1 35091
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_3
timestamp 1662439860
transform -1 0 5045 0 1 32915
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_4
timestamp 1662439860
transform 1 0 2009 0 -1 34003
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  sky130_fd_sc_hd__nand2_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform -1 0 2561 0 1 34003
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  sky130_fd_sc_hd__nand2_1_1
timestamp 1662439860
transform 1 0 2285 0 -1 34003
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 2193 0 1 34003
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_1
timestamp 1662439860
transform -1 0 3665 0 -1 35091
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_2
timestamp 1662439860
transform -1 0 3665 0 1 32915
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_3
timestamp 1662439860
transform 1 0 1917 0 -1 34003
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_4
timestamp 1662439860
transform 1 0 2101 0 1 32915
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_5
timestamp 1662439860
transform 1 0 1428 0 -1 35092
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_6
timestamp 1662439860
transform 1 0 5321 0 1 34003
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_7
timestamp 1662439860
transform 1 0 5321 0 -1 34003
box -38 -48 130 592
<< labels >>
flabel metal4 s 0 0 400 64000 0 FreeSans 1600 90 0 0 VDD
port 1 nsew power bidirectional
flabel metal4 s 463 0 863 64000 0 FreeSans 1600 90 0 0 VSS
port 2 nsew power bidirectional
flabel locali 1939 34217 1973 34269 0 FreeSans 800 0 0 0 clk
port 3 nsew signal input
flabel metal1 3519 33023 3556 33058 0 FreeSans 320 180 0 0 phi2
flabel metal1 3500 34829 3537 34876 0 FreeSans 320 180 0 0 phi1_n
flabel metal1 3527 33131 3564 33178 0 FreeSans 320 180 0 0 phi2_n
flabel metal1 3499 34946 3535 34981 0 FreeSans 320 180 0 0 phi1
flabel metal2 2468 28000 2867 36000 0 FreeSans 1600 90 0 0 vcm
port 4 nsew analog output
flabel metal4 2306 35775 2467 36000 0 FreeSans 480 90 0 0 mimtop1
flabel space 4189 35754 4348 36000 0 FreeSans 480 90 0 0 mimbot1
flabel metal4 3093 28001 3337 28321 0 FreeSans 480 90 0 0 mimtop2
flabel metal4 25502 0 25902 64000 0 FreeSans 1600 90 0 0 VDD
port 1 nsew power bidirectional
flabel metal4 25028 0 25428 64000 0 FreeSans 1600 90 0 0 VSS
port 2 nsew power bidirectional
flabel metal4 s 25970 0 26370 64000 0 FreeSans 1600 90 0 0 vcm
port 4 nsew analog output
<< properties >>
string LEFclass CORE
string LEForigin 0 0
string LEFsource USER
<< end >>
