magic
tech sky130A
magscale 1 2
timestamp 1659713046
<< error_p >>
rect 22 1206 2296 1234
rect 22 994 28 1000
rect 60 994 82 1052
rect 2296 1000 2318 1052
rect 2290 994 2318 1000
rect 16 992 23 994
rect 0 932 23 992
rect 16 930 23 932
rect 54 930 86 994
rect 2295 930 2328 994
rect 22 924 28 930
rect 22 754 28 760
rect 60 754 82 930
rect 2290 924 2318 930
rect 2296 760 2318 924
rect 2290 754 2318 760
rect 16 752 23 754
rect 0 692 23 752
rect 16 690 23 692
rect 54 690 86 754
rect 2295 690 2328 754
rect 22 684 28 690
rect 22 514 28 520
rect 60 514 82 690
rect 2290 684 2318 690
rect 2296 520 2318 684
rect 2290 514 2318 520
rect 16 512 23 514
rect 0 452 23 512
rect 16 450 23 452
rect 54 450 86 514
rect 2295 450 2328 514
rect 22 444 28 450
rect 22 274 28 280
rect 60 274 82 450
rect 2290 444 2318 450
rect 2296 280 2318 444
rect 2290 274 2318 280
rect 16 272 23 274
rect 0 212 23 272
rect 16 210 23 212
rect 54 210 86 274
rect 2295 210 2328 274
rect 22 204 28 210
rect 60 60 82 210
rect 2290 204 2318 210
rect 60 32 742 60
rect 818 32 1500 60
rect 1576 32 2258 60
rect 2296 32 2318 204
rect 90 26 144 32
rect 240 26 294 32
rect 506 26 560 32
rect 656 26 710 32
rect 848 26 902 32
rect 998 26 1052 32
rect 1264 26 1318 32
rect 1414 26 1468 32
rect 1606 26 1660 32
rect 1756 26 1810 32
rect 2022 26 2076 32
rect 2172 26 2226 32
<< metal1 >>
rect 22 1180 90 1206
rect 144 1180 240 1206
rect 294 1180 506 1206
rect 560 1180 656 1206
rect 710 1180 742 1206
rect 22 1176 742 1180
rect 780 1180 848 1206
rect 902 1180 998 1206
rect 1052 1180 1264 1206
rect 1318 1180 1414 1206
rect 1468 1180 1500 1206
rect 780 1176 1500 1180
rect 1538 1180 1606 1206
rect 1660 1180 1756 1206
rect 1810 1180 2022 1206
rect 2076 1180 2172 1206
rect 2226 1180 2258 1206
rect 1538 1176 2258 1180
rect 22 26 742 32
rect 22 0 90 26
rect 144 0 240 26
rect 294 0 506 26
rect 560 0 656 26
rect 710 0 742 26
rect 780 26 1500 32
rect 780 0 848 26
rect 902 0 998 26
rect 1052 0 1264 26
rect 1318 0 1414 26
rect 1468 0 1500 26
rect 1538 26 2258 32
rect 1538 0 1606 26
rect 1660 0 1756 26
rect 1810 0 2022 26
rect 2076 0 2172 26
rect 2226 0 2258 26
<< via1 >>
rect 90 1180 144 1206
rect 240 1180 294 1206
rect 506 1180 560 1206
rect 656 1180 710 1206
rect 848 1180 902 1206
rect 998 1180 1052 1206
rect 1264 1180 1318 1206
rect 1414 1180 1468 1206
rect 1606 1180 1660 1206
rect 1756 1180 1810 1206
rect 2022 1180 2076 1206
rect 2172 1180 2226 1206
rect 90 0 144 26
rect 240 0 294 26
rect 506 0 560 26
rect 656 0 710 26
rect 848 0 902 26
rect 998 0 1052 26
rect 1264 0 1318 26
rect 1414 0 1468 26
rect 1606 0 1660 26
rect 1756 0 1810 26
rect 2022 0 2076 26
rect 2172 0 2226 26
<< metal2 >>
rect 22 1180 90 1206
rect 144 1180 240 1206
rect 294 1180 506 1206
rect 560 1180 656 1206
rect 710 1180 848 1206
rect 902 1180 998 1206
rect 1052 1180 1264 1206
rect 1318 1180 1414 1206
rect 1468 1180 1606 1206
rect 1660 1180 1756 1206
rect 1810 1180 2022 1206
rect 2076 1180 2172 1206
rect 2226 1180 2296 1206
rect 22 1174 2296 1180
rect 22 1152 344 1174
rect 456 1152 1102 1174
rect 1214 1152 1860 1174
rect 1972 1152 2296 1174
rect 22 1016 314 1152
rect 372 1122 428 1146
rect 344 1116 456 1122
rect 344 1054 354 1116
rect 446 1054 456 1116
rect 344 1046 456 1054
rect 22 910 344 1016
rect 22 774 314 910
rect 372 880 428 1046
rect 486 1016 1072 1152
rect 1130 1122 1186 1146
rect 1102 1116 1214 1122
rect 1102 1054 1112 1116
rect 1204 1054 1214 1116
rect 1102 1046 1214 1054
rect 456 910 1102 1016
rect 344 874 456 880
rect 344 812 354 874
rect 446 812 456 874
rect 344 804 456 812
rect 22 670 344 774
rect 22 534 314 670
rect 372 640 428 804
rect 486 774 1072 910
rect 1130 880 1186 1046
rect 1244 1016 1830 1152
rect 1888 1122 1944 1146
rect 1860 1116 1972 1122
rect 1860 1054 1870 1116
rect 1962 1054 1972 1116
rect 1860 1046 1972 1054
rect 1214 910 1860 1016
rect 1102 874 1214 880
rect 1102 812 1112 874
rect 1204 812 1214 874
rect 1102 804 1214 812
rect 456 670 1102 774
rect 344 634 456 640
rect 344 572 354 634
rect 446 572 456 634
rect 344 564 456 572
rect 22 430 344 534
rect 22 294 314 430
rect 372 400 428 564
rect 486 534 1072 670
rect 1130 640 1186 804
rect 1244 774 1830 910
rect 1888 880 1944 1046
rect 2002 1016 2296 1152
rect 1972 910 2296 1016
rect 1860 874 1972 880
rect 1860 812 1870 874
rect 1962 812 1972 874
rect 1860 804 1972 812
rect 1214 670 1860 774
rect 1102 634 1214 640
rect 1102 572 1112 634
rect 1204 572 1214 634
rect 1102 564 1214 572
rect 456 430 1102 534
rect 344 394 456 400
rect 344 332 354 394
rect 446 332 456 394
rect 344 324 456 332
rect 22 190 344 294
rect 22 56 314 190
rect 372 160 428 324
rect 486 294 1072 430
rect 1130 400 1186 564
rect 1244 534 1830 670
rect 1888 640 1944 804
rect 2002 774 2296 910
rect 1972 670 2296 774
rect 1860 634 1972 640
rect 1860 572 1870 634
rect 1962 572 1972 634
rect 1860 564 1972 572
rect 1214 430 1860 534
rect 1102 394 1214 400
rect 1102 332 1112 394
rect 1204 332 1214 394
rect 1102 324 1214 332
rect 456 190 1102 294
rect 344 154 456 160
rect 344 92 354 154
rect 446 92 456 154
rect 344 84 456 92
rect 372 60 428 84
rect 486 56 1072 190
rect 1130 160 1186 324
rect 1244 294 1830 430
rect 1888 400 1944 564
rect 2002 534 2296 670
rect 1972 430 2296 534
rect 1860 394 1972 400
rect 1860 332 1870 394
rect 1962 332 1972 394
rect 1860 324 1972 332
rect 1214 190 1860 294
rect 1102 154 1214 160
rect 1102 92 1112 154
rect 1204 92 1214 154
rect 1102 84 1214 92
rect 1130 60 1186 84
rect 1244 56 1830 190
rect 1888 160 1944 324
rect 2002 294 2296 430
rect 1972 190 2296 294
rect 1860 154 1972 160
rect 1860 92 1870 154
rect 1962 92 1972 154
rect 1860 84 1972 92
rect 1888 60 1944 84
rect 2002 56 2296 190
rect 22 32 344 56
rect 456 32 1102 56
rect 1214 32 1860 56
rect 1972 32 2296 56
rect 22 26 2296 32
rect 22 0 90 26
rect 144 0 240 26
rect 294 0 506 26
rect 560 0 656 26
rect 710 0 848 26
rect 902 0 998 26
rect 1052 0 1264 26
rect 1318 0 1414 26
rect 1468 0 1606 26
rect 1660 0 1756 26
rect 1810 0 2022 26
rect 2076 0 2172 26
rect 2226 0 2296 26
<< via2 >>
rect 354 1054 446 1116
rect 1112 1054 1204 1116
rect 354 812 446 874
rect 1870 1054 1962 1116
rect 1112 812 1204 874
rect 354 572 446 634
rect 1870 812 1962 874
rect 1112 572 1204 634
rect 354 332 446 394
rect 1870 572 1962 634
rect 1112 332 1204 394
rect 354 92 446 154
rect 1870 332 1962 394
rect 1112 92 1204 154
rect 1870 92 1962 154
<< metal3 >>
rect 344 1116 456 1122
rect 344 1114 354 1116
rect 128 1054 354 1114
rect 446 1114 456 1116
rect 1102 1116 1214 1122
rect 1102 1114 1112 1116
rect 446 1054 674 1114
rect 886 1054 1112 1114
rect 1204 1114 1214 1116
rect 1860 1116 1972 1122
rect 1860 1114 1870 1116
rect 1204 1054 1432 1114
rect 1644 1054 1870 1114
rect 1962 1114 1972 1116
rect 1962 1054 2190 1114
rect 344 1046 456 1054
rect 1102 1046 1214 1054
rect 1860 1046 1972 1054
rect 54 992 60 994
rect 742 992 748 994
rect 54 932 314 992
rect 486 932 748 992
rect 54 930 60 932
rect 742 930 748 932
rect 812 992 818 994
rect 1500 992 1506 994
rect 812 932 1072 992
rect 1244 932 1506 992
rect 812 930 818 932
rect 1500 930 1506 932
rect 1570 992 1576 994
rect 2258 992 2264 994
rect 1570 932 1830 992
rect 2002 932 2264 992
rect 1570 930 1576 932
rect 2258 930 2264 932
rect 344 874 456 880
rect 344 872 354 874
rect 128 812 354 872
rect 446 872 456 874
rect 1102 874 1214 880
rect 1102 872 1112 874
rect 446 812 674 872
rect 886 812 1112 872
rect 1204 872 1214 874
rect 1860 874 1972 880
rect 1860 872 1870 874
rect 1204 812 1432 872
rect 1644 812 1870 872
rect 1962 872 1972 874
rect 1962 812 2190 872
rect 344 804 456 812
rect 1102 804 1214 812
rect 1860 804 1972 812
rect 54 752 60 754
rect 742 752 748 754
rect 54 692 314 752
rect 486 692 748 752
rect 54 690 60 692
rect 742 690 748 692
rect 812 752 818 754
rect 1500 752 1506 754
rect 812 692 1072 752
rect 1244 692 1506 752
rect 812 690 818 692
rect 1500 690 1506 692
rect 1570 752 1576 754
rect 2258 752 2264 754
rect 1570 692 1830 752
rect 2002 692 2264 752
rect 1570 690 1576 692
rect 2258 690 2264 692
rect 344 634 456 640
rect 344 632 354 634
rect 128 572 354 632
rect 446 632 456 634
rect 1102 634 1214 640
rect 1102 632 1112 634
rect 446 572 674 632
rect 886 572 1112 632
rect 1204 632 1214 634
rect 1860 634 1972 640
rect 1860 632 1870 634
rect 1204 572 1432 632
rect 1644 572 1870 632
rect 1962 632 1972 634
rect 1962 572 2190 632
rect 344 564 456 572
rect 1102 564 1214 572
rect 1860 564 1972 572
rect 54 512 60 514
rect 742 512 748 514
rect 54 452 314 512
rect 486 452 748 512
rect 54 450 60 452
rect 742 450 748 452
rect 812 512 818 514
rect 1500 512 1506 514
rect 812 452 1072 512
rect 1244 452 1506 512
rect 812 450 818 452
rect 1500 450 1506 452
rect 1570 512 1576 514
rect 2258 512 2264 514
rect 1570 452 1830 512
rect 2002 452 2264 512
rect 1570 450 1576 452
rect 2258 450 2264 452
rect 344 394 456 400
rect 344 392 354 394
rect 128 332 354 392
rect 446 392 456 394
rect 1102 394 1214 400
rect 1102 392 1112 394
rect 446 332 674 392
rect 886 332 1112 392
rect 1204 392 1214 394
rect 1860 394 1972 400
rect 1860 392 1870 394
rect 1204 332 1432 392
rect 1644 332 1870 392
rect 1962 392 1972 394
rect 1962 332 2190 392
rect 344 324 456 332
rect 1102 324 1214 332
rect 1860 324 1972 332
rect 54 272 60 274
rect 742 272 748 274
rect 54 212 314 272
rect 486 212 748 272
rect 54 210 60 212
rect 742 210 748 212
rect 812 272 818 274
rect 1500 272 1506 274
rect 812 212 1072 272
rect 1244 212 1506 272
rect 812 210 818 212
rect 1500 210 1506 212
rect 1570 272 1576 274
rect 2258 272 2264 274
rect 1570 212 1830 272
rect 2002 212 2264 272
rect 1570 210 1576 212
rect 2258 210 2264 212
rect 344 154 456 160
rect 344 152 354 154
rect 128 92 354 152
rect 446 152 456 154
rect 1102 154 1214 160
rect 1102 152 1112 154
rect 446 92 674 152
rect 886 92 1112 152
rect 1204 152 1214 154
rect 1860 154 1972 160
rect 1860 152 1870 154
rect 1204 92 1432 152
rect 1644 92 1870 152
rect 1962 152 1972 154
rect 1962 92 2190 152
rect 344 84 456 92
rect 1102 84 1214 92
rect 1860 84 1972 92
<< via3 >>
rect 22 930 54 994
rect 748 930 812 994
rect 1506 930 1570 994
rect 2264 930 2296 994
rect 22 690 54 754
rect 748 690 812 754
rect 1506 690 1570 754
rect 2264 690 2296 754
rect 22 450 54 514
rect 748 450 812 514
rect 1506 450 1570 514
rect 2264 450 2296 514
rect 22 210 54 274
rect 748 210 812 274
rect 1506 210 1570 274
rect 2264 210 2296 274
<< metal4 >>
rect 22 1174 2296 1206
rect 22 994 60 1052
rect 54 930 60 994
rect 22 754 60 930
rect 54 690 60 754
rect 22 514 60 690
rect 742 994 818 1174
rect 742 930 748 994
rect 812 930 818 994
rect 742 754 818 930
rect 742 690 748 754
rect 812 690 818 754
rect 742 598 818 690
rect 1500 994 1576 1174
rect 1500 930 1506 994
rect 1570 930 1576 994
rect 1500 754 1576 930
rect 1500 690 1506 754
rect 1570 690 1576 754
rect 1500 600 1576 690
rect 2258 994 2296 1052
rect 2258 930 2264 994
rect 2258 754 2296 930
rect 2258 690 2264 754
rect 54 450 60 514
rect 22 274 60 450
rect 54 210 60 274
rect 22 32 60 210
rect 742 514 818 518
rect 742 450 748 514
rect 812 450 818 514
rect 742 274 818 450
rect 742 210 748 274
rect 812 210 818 274
rect 742 32 818 210
rect 1500 514 1576 520
rect 1500 450 1506 514
rect 1570 450 1576 514
rect 1500 274 1576 450
rect 1500 210 1506 274
rect 1570 210 1576 274
rect 1500 32 1576 210
rect 2258 514 2296 690
rect 2258 450 2264 514
rect 2258 274 2296 450
rect 2258 210 2264 274
rect 2258 32 2296 210
rect 22 0 2296 32
<< end >>
