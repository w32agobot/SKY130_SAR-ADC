magic
tech sky130A
magscale 1 2
timestamp 1662367448
<< nwell >>
rect 2402 226 2858 230
rect 44 16 2858 226
rect 44 -178 2570 16
rect 44 -196 2336 -178
rect 570 -198 812 -196
rect 1178 -546 2336 -196
<< nmos >>
rect 144 -910 174 -510
rect 240 -910 270 -510
rect 336 -910 366 -510
rect 432 -910 462 -510
rect 528 -910 558 -510
rect 624 -910 654 -510
rect 720 -910 750 -510
rect 816 -910 846 -510
rect 144 -1170 174 -1070
rect 240 -1170 270 -1070
rect 336 -1170 366 -1070
rect 432 -1170 462 -1070
rect 528 -1170 558 -1070
rect 624 -1170 654 -1070
rect 720 -1170 750 -1070
rect 816 -1170 846 -1070
rect 1598 -1176 1628 -776
rect 1694 -1176 1724 -776
rect 1790 -1176 1820 -776
rect 1886 -1176 1916 -776
<< pmos >>
rect 144 -96 174 4
rect 240 -96 270 4
rect 336 -96 366 4
rect 432 -96 462 4
rect 528 -96 558 4
rect 624 -96 654 4
rect 720 -96 750 4
rect 816 -96 846 4
rect 1276 -446 1306 -46
rect 1372 -446 1402 -46
rect 1598 -446 1628 -46
rect 1694 -446 1724 -46
rect 1790 -446 1820 -46
rect 1886 -446 1916 -46
rect 2112 -446 2142 -46
rect 2208 -446 2238 -46
<< ndiff >>
rect 82 -522 144 -510
rect 82 -898 94 -522
rect 128 -898 144 -522
rect 82 -910 144 -898
rect 174 -522 240 -510
rect 174 -898 190 -522
rect 224 -898 240 -522
rect 174 -910 240 -898
rect 270 -522 336 -510
rect 270 -898 286 -522
rect 320 -898 336 -522
rect 270 -910 336 -898
rect 366 -522 432 -510
rect 366 -898 382 -522
rect 416 -898 432 -522
rect 366 -910 432 -898
rect 462 -522 528 -510
rect 462 -898 478 -522
rect 512 -898 528 -522
rect 462 -910 528 -898
rect 558 -522 624 -510
rect 558 -898 574 -522
rect 608 -898 624 -522
rect 558 -910 624 -898
rect 654 -522 720 -510
rect 654 -898 670 -522
rect 704 -898 720 -522
rect 654 -910 720 -898
rect 750 -522 816 -510
rect 750 -898 766 -522
rect 800 -898 816 -522
rect 750 -910 816 -898
rect 846 -522 908 -510
rect 846 -898 862 -522
rect 896 -898 908 -522
rect 846 -910 908 -898
rect 1536 -788 1598 -776
rect 82 -1082 144 -1070
rect 82 -1158 94 -1082
rect 128 -1158 144 -1082
rect 82 -1170 144 -1158
rect 174 -1082 240 -1070
rect 174 -1158 190 -1082
rect 224 -1158 240 -1082
rect 174 -1170 240 -1158
rect 270 -1082 336 -1070
rect 270 -1158 286 -1082
rect 320 -1158 336 -1082
rect 270 -1170 336 -1158
rect 366 -1082 432 -1070
rect 366 -1158 382 -1082
rect 416 -1158 432 -1082
rect 366 -1170 432 -1158
rect 462 -1082 528 -1070
rect 462 -1158 478 -1082
rect 512 -1158 528 -1082
rect 462 -1170 528 -1158
rect 558 -1082 624 -1070
rect 558 -1158 574 -1082
rect 608 -1158 624 -1082
rect 558 -1170 624 -1158
rect 654 -1082 720 -1070
rect 654 -1158 670 -1082
rect 704 -1158 720 -1082
rect 654 -1170 720 -1158
rect 750 -1082 816 -1070
rect 750 -1158 766 -1082
rect 800 -1158 816 -1082
rect 750 -1170 816 -1158
rect 846 -1082 908 -1070
rect 846 -1158 862 -1082
rect 896 -1158 908 -1082
rect 846 -1170 908 -1158
rect 1536 -1164 1548 -788
rect 1582 -1164 1598 -788
rect 1536 -1176 1598 -1164
rect 1628 -788 1694 -776
rect 1628 -1164 1644 -788
rect 1678 -1164 1694 -788
rect 1628 -1176 1694 -1164
rect 1724 -788 1790 -776
rect 1724 -1164 1740 -788
rect 1774 -1164 1790 -788
rect 1724 -1176 1790 -1164
rect 1820 -788 1886 -776
rect 1820 -1164 1836 -788
rect 1870 -1164 1886 -788
rect 1820 -1176 1886 -1164
rect 1916 -788 1978 -776
rect 1916 -1164 1932 -788
rect 1966 -1164 1978 -788
rect 1916 -1176 1978 -1164
<< pdiff >>
rect 82 -8 144 4
rect 82 -84 94 -8
rect 128 -84 144 -8
rect 82 -96 144 -84
rect 174 -8 240 4
rect 174 -84 190 -8
rect 224 -84 240 -8
rect 174 -96 240 -84
rect 270 -8 336 4
rect 270 -84 286 -8
rect 320 -84 336 -8
rect 270 -96 336 -84
rect 366 -8 432 4
rect 366 -84 382 -8
rect 416 -84 432 -8
rect 366 -96 432 -84
rect 462 -8 528 4
rect 462 -84 478 -8
rect 512 -84 528 -8
rect 462 -96 528 -84
rect 558 -8 624 4
rect 558 -84 574 -8
rect 608 -84 624 -8
rect 558 -96 624 -84
rect 654 -8 720 4
rect 654 -84 670 -8
rect 704 -84 720 -8
rect 654 -96 720 -84
rect 750 -8 816 4
rect 750 -84 766 -8
rect 800 -84 816 -8
rect 750 -96 816 -84
rect 846 -8 908 4
rect 846 -84 862 -8
rect 896 -84 908 -8
rect 846 -96 908 -84
rect 1214 -58 1276 -46
rect 1214 -434 1226 -58
rect 1260 -434 1276 -58
rect 1214 -446 1276 -434
rect 1306 -58 1372 -46
rect 1306 -434 1322 -58
rect 1356 -434 1372 -58
rect 1306 -446 1372 -434
rect 1402 -58 1464 -46
rect 1402 -434 1418 -58
rect 1452 -434 1464 -58
rect 1402 -446 1464 -434
rect 1536 -58 1598 -46
rect 1536 -434 1548 -58
rect 1582 -434 1598 -58
rect 1536 -446 1598 -434
rect 1628 -58 1694 -46
rect 1628 -434 1644 -58
rect 1678 -434 1694 -58
rect 1628 -446 1694 -434
rect 1724 -58 1790 -46
rect 1724 -434 1740 -58
rect 1774 -434 1790 -58
rect 1724 -446 1790 -434
rect 1820 -58 1886 -46
rect 1820 -434 1836 -58
rect 1870 -434 1886 -58
rect 1820 -446 1886 -434
rect 1916 -58 1978 -46
rect 1916 -434 1932 -58
rect 1966 -434 1978 -58
rect 1916 -446 1978 -434
rect 2050 -58 2112 -46
rect 2050 -434 2062 -58
rect 2096 -434 2112 -58
rect 2050 -446 2112 -434
rect 2142 -58 2208 -46
rect 2142 -434 2158 -58
rect 2192 -434 2208 -58
rect 2142 -446 2208 -434
rect 2238 -58 2300 -46
rect 2238 -434 2254 -58
rect 2288 -434 2300 -58
rect 2238 -446 2300 -434
<< ndiffc >>
rect 94 -898 128 -522
rect 190 -898 224 -522
rect 286 -898 320 -522
rect 382 -898 416 -522
rect 478 -898 512 -522
rect 574 -898 608 -522
rect 670 -898 704 -522
rect 766 -898 800 -522
rect 862 -898 896 -522
rect 94 -1158 128 -1082
rect 190 -1158 224 -1082
rect 286 -1158 320 -1082
rect 382 -1158 416 -1082
rect 478 -1158 512 -1082
rect 574 -1158 608 -1082
rect 670 -1158 704 -1082
rect 766 -1158 800 -1082
rect 862 -1158 896 -1082
rect 1548 -1164 1582 -788
rect 1644 -1164 1678 -788
rect 1740 -1164 1774 -788
rect 1836 -1164 1870 -788
rect 1932 -1164 1966 -788
<< pdiffc >>
rect 94 -84 128 -8
rect 190 -84 224 -8
rect 286 -84 320 -8
rect 382 -84 416 -8
rect 478 -84 512 -8
rect 574 -84 608 -8
rect 670 -84 704 -8
rect 766 -84 800 -8
rect 862 -84 896 -8
rect 1226 -434 1260 -58
rect 1322 -434 1356 -58
rect 1418 -434 1452 -58
rect 1548 -434 1582 -58
rect 1644 -434 1678 -58
rect 1740 -434 1774 -58
rect 1836 -434 1870 -58
rect 1932 -434 1966 -58
rect 2062 -434 2096 -58
rect 2158 -434 2192 -58
rect 2254 -434 2288 -58
<< psubdiff >>
rect -286 3918 -164 3944
rect -286 3844 -262 3918
rect -188 3844 -164 3918
rect -286 3820 -164 3844
rect 262 3918 384 3944
rect 262 3844 286 3918
rect 360 3844 384 3918
rect 262 3820 384 3844
rect 810 3918 932 3944
rect 810 3844 834 3918
rect 908 3844 932 3918
rect 810 3820 932 3844
rect 1358 3918 1480 3944
rect 1358 3844 1382 3918
rect 1456 3844 1480 3918
rect 1358 3820 1480 3844
rect 1906 3918 2028 3944
rect 1906 3844 1930 3918
rect 2004 3844 2028 3918
rect 1906 3820 2028 3844
rect 2436 3918 2558 3944
rect 2436 3844 2460 3918
rect 2534 3844 2558 3918
rect 2436 3820 2558 3844
rect 2984 3918 3106 3944
rect 2984 3844 3008 3918
rect 3082 3844 3106 3918
rect 2984 3820 3106 3844
rect 3534 3918 3656 3944
rect 3534 3844 3558 3918
rect 3632 3844 3656 3918
rect 3534 3820 3656 3844
rect -652 3442 -530 3468
rect -652 3368 -628 3442
rect -554 3368 -530 3442
rect -652 3344 -530 3368
rect 4030 3374 4152 3400
rect 4030 3300 4054 3374
rect 4128 3300 4152 3374
rect 4030 3276 4152 3300
rect -652 2968 -530 2994
rect -652 2894 -628 2968
rect -554 2894 -530 2968
rect -652 2870 -530 2894
rect 4030 2900 4152 2926
rect 4030 2826 4054 2900
rect 4128 2826 4152 2900
rect 4030 2802 4152 2826
rect -652 2494 -530 2520
rect -652 2420 -628 2494
rect -554 2420 -530 2494
rect -652 2396 -530 2420
rect 4030 2426 4152 2452
rect 4030 2352 4054 2426
rect 4128 2352 4152 2426
rect 4030 2328 4152 2352
rect -652 2020 -530 2046
rect -652 1946 -628 2020
rect -554 1946 -530 2020
rect -652 1922 -530 1946
rect 4030 1950 4152 1976
rect 4030 1876 4054 1950
rect 4128 1876 4152 1950
rect 4030 1852 4152 1876
rect -652 1546 -530 1572
rect -652 1472 -628 1546
rect -554 1472 -530 1546
rect -652 1448 -530 1472
rect 4030 1474 4152 1500
rect 4030 1400 4054 1474
rect 4128 1400 4152 1474
rect 4030 1376 4152 1400
rect -652 1072 -530 1098
rect -652 998 -628 1072
rect -554 998 -530 1072
rect -652 974 -530 998
rect 4030 1000 4152 1026
rect 4030 926 4054 1000
rect 4128 926 4152 1000
rect 4030 902 4152 926
rect -652 598 -530 624
rect -652 524 -628 598
rect -554 524 -530 598
rect -652 500 -530 524
rect 4028 526 4150 552
rect 4028 452 4052 526
rect 4126 452 4150 526
rect 4028 434 4150 452
rect -652 -88 -530 -62
rect -652 -162 -628 -88
rect -554 -162 -530 -88
rect -652 -186 -530 -162
rect 4028 -86 4150 -60
rect 4028 -160 4052 -86
rect 4126 -160 4150 -86
rect 4028 -184 4150 -160
rect -660 -614 -538 -588
rect -660 -688 -636 -614
rect -562 -688 -538 -614
rect -660 -712 -538 -688
rect 4028 -560 4150 -534
rect 4028 -634 4052 -560
rect 4126 -634 4150 -560
rect 4028 -658 4150 -634
rect -660 -1088 -538 -1062
rect -660 -1162 -636 -1088
rect -562 -1162 -538 -1088
rect -660 -1186 -538 -1162
rect 4028 -1034 4150 -1008
rect 4028 -1108 4052 -1034
rect 4126 -1108 4150 -1034
rect 4028 -1132 4150 -1108
rect 1542 -1324 1566 -1288
rect 1602 -1324 1658 -1288
rect 1694 -1324 1750 -1288
rect 1786 -1324 1842 -1288
rect 1878 -1324 1934 -1288
rect 1970 -1324 1994 -1288
rect 1542 -1326 1994 -1324
rect 76 -1332 894 -1330
rect 76 -1368 100 -1332
rect 136 -1368 218 -1332
rect 254 -1368 336 -1332
rect 372 -1368 454 -1332
rect 490 -1368 572 -1332
rect 608 -1368 690 -1332
rect 726 -1368 808 -1332
rect 844 -1368 894 -1332
rect 76 -1372 894 -1368
rect -646 -1740 -524 -1714
rect -646 -1814 -622 -1740
rect -548 -1814 -524 -1740
rect -646 -1838 -524 -1814
rect 4028 -1770 4150 -1744
rect 4028 -1844 4052 -1770
rect 4126 -1844 4150 -1770
rect 4028 -1868 4150 -1844
rect -646 -2214 -524 -2188
rect -646 -2288 -622 -2214
rect -548 -2288 -524 -2214
rect -646 -2312 -524 -2288
rect 4028 -2244 4150 -2218
rect 4028 -2318 4052 -2244
rect 4126 -2318 4150 -2244
rect 4028 -2342 4150 -2318
rect -646 -2688 -524 -2662
rect -646 -2762 -622 -2688
rect -548 -2762 -524 -2688
rect -646 -2786 -524 -2762
rect 4028 -2718 4150 -2692
rect 4028 -2792 4052 -2718
rect 4126 -2792 4150 -2718
rect 4028 -2816 4150 -2792
rect -646 -3164 -524 -3138
rect -646 -3238 -622 -3164
rect -548 -3238 -524 -3164
rect -646 -3262 -524 -3238
rect 4028 -3192 4150 -3166
rect 4028 -3266 4052 -3192
rect 4126 -3266 4150 -3192
rect 4028 -3290 4150 -3266
rect -646 -3638 -524 -3612
rect -646 -3712 -622 -3638
rect -548 -3712 -524 -3638
rect -646 -3736 -524 -3712
rect 4028 -3666 4150 -3640
rect 4028 -3740 4052 -3666
rect 4126 -3740 4150 -3666
rect 4028 -3764 4150 -3740
rect -646 -4112 -524 -4086
rect -646 -4186 -622 -4112
rect -548 -4186 -524 -4112
rect -646 -4210 -524 -4186
rect 4028 -4140 4150 -4114
rect 4028 -4214 4052 -4140
rect 4126 -4214 4150 -4140
rect 4028 -4238 4150 -4214
rect -646 -4586 -524 -4560
rect -646 -4660 -622 -4586
rect -548 -4660 -524 -4586
rect -646 -4684 -524 -4660
rect 4030 -4614 4152 -4588
rect 4030 -4688 4054 -4614
rect 4128 -4688 4152 -4614
rect 4030 -4712 4152 -4688
rect -116 -5000 6 -4974
rect -116 -5074 -92 -5000
rect -18 -5074 6 -5000
rect -116 -5098 6 -5074
rect 432 -5000 554 -4974
rect 432 -5074 456 -5000
rect 530 -5074 554 -5000
rect 432 -5098 554 -5074
rect 980 -5000 1102 -4974
rect 980 -5074 1004 -5000
rect 1078 -5074 1102 -5000
rect 980 -5098 1102 -5074
rect 1528 -5000 1650 -4974
rect 1528 -5074 1552 -5000
rect 1626 -5074 1650 -5000
rect 1528 -5098 1650 -5074
rect 2076 -5000 2198 -4974
rect 2076 -5074 2100 -5000
rect 2174 -5074 2198 -5000
rect 2076 -5098 2198 -5074
rect 2624 -5000 2746 -4974
rect 2624 -5074 2648 -5000
rect 2722 -5074 2746 -5000
rect 2624 -5098 2746 -5074
rect 3174 -5000 3296 -4974
rect 3174 -5074 3198 -5000
rect 3272 -5074 3296 -5000
rect 3174 -5098 3296 -5074
<< nsubdiff >>
rect 1382 110 2106 118
rect 82 100 938 108
rect 82 66 112 100
rect 146 66 196 100
rect 230 66 280 100
rect 314 66 364 100
rect 398 66 448 100
rect 482 66 532 100
rect 566 66 616 100
rect 650 66 700 100
rect 734 66 784 100
rect 818 66 874 100
rect 908 66 938 100
rect 1382 76 1420 110
rect 1454 76 1504 110
rect 1538 76 1588 110
rect 1622 76 1672 110
rect 1706 76 1756 110
rect 1790 76 1840 110
rect 1874 76 1924 110
rect 1958 76 2008 110
rect 2042 76 2106 110
rect 1382 70 2106 76
rect 82 60 938 66
<< psubdiffcont >>
rect -262 3844 -188 3918
rect 286 3844 360 3918
rect 834 3844 908 3918
rect 1382 3844 1456 3918
rect 1930 3844 2004 3918
rect 2460 3844 2534 3918
rect 3008 3844 3082 3918
rect 3558 3844 3632 3918
rect -628 3368 -554 3442
rect 4054 3300 4128 3374
rect -628 2894 -554 2968
rect 4054 2826 4128 2900
rect -628 2420 -554 2494
rect 4054 2352 4128 2426
rect -628 1946 -554 2020
rect 4054 1876 4128 1950
rect -628 1472 -554 1546
rect 4054 1400 4128 1474
rect -628 998 -554 1072
rect 4054 926 4128 1000
rect -628 524 -554 598
rect 4052 452 4126 526
rect -628 -162 -554 -88
rect 4052 -160 4126 -86
rect -636 -688 -562 -614
rect 4052 -634 4126 -560
rect -636 -1162 -562 -1088
rect 4052 -1108 4126 -1034
rect 1566 -1324 1602 -1288
rect 1658 -1324 1694 -1288
rect 1750 -1324 1786 -1288
rect 1842 -1324 1878 -1288
rect 1934 -1324 1970 -1288
rect 100 -1368 136 -1332
rect 218 -1368 254 -1332
rect 336 -1368 372 -1332
rect 454 -1368 490 -1332
rect 572 -1368 608 -1332
rect 690 -1368 726 -1332
rect 808 -1368 844 -1332
rect -622 -1814 -548 -1740
rect 4052 -1844 4126 -1770
rect -622 -2288 -548 -2214
rect 4052 -2318 4126 -2244
rect -622 -2762 -548 -2688
rect 4052 -2792 4126 -2718
rect -622 -3238 -548 -3164
rect 4052 -3266 4126 -3192
rect -622 -3712 -548 -3638
rect 4052 -3740 4126 -3666
rect -622 -4186 -548 -4112
rect 4052 -4214 4126 -4140
rect -622 -4660 -548 -4586
rect 4054 -4688 4128 -4614
rect -92 -5074 -18 -5000
rect 456 -5074 530 -5000
rect 1004 -5074 1078 -5000
rect 1552 -5074 1626 -5000
rect 2100 -5074 2174 -5000
rect 2648 -5074 2722 -5000
rect 3198 -5074 3272 -5000
<< nsubdiffcont >>
rect 112 66 146 100
rect 196 66 230 100
rect 280 66 314 100
rect 364 66 398 100
rect 448 66 482 100
rect 532 66 566 100
rect 616 66 650 100
rect 700 66 734 100
rect 784 66 818 100
rect 874 66 908 100
rect 1420 76 1454 110
rect 1504 76 1538 110
rect 1588 76 1622 110
rect 1672 76 1706 110
rect 1756 76 1790 110
rect 1840 76 1874 110
rect 1924 76 1958 110
rect 2008 76 2042 110
<< poly >>
rect 144 4 174 30
rect 240 4 270 30
rect 336 4 366 30
rect 432 4 462 30
rect 528 4 558 30
rect 624 4 654 30
rect 720 4 750 30
rect 816 4 846 30
rect 1276 -46 1306 -20
rect 1372 -46 1402 -20
rect 1598 -46 1628 -20
rect 1694 -46 1724 -20
rect 1790 -46 1820 -20
rect 1886 -46 1916 -20
rect 2112 -46 2142 -20
rect 2208 -46 2238 -20
rect 144 -122 174 -96
rect 240 -122 270 -96
rect 336 -122 366 -96
rect 432 -122 462 -96
rect 528 -122 558 -96
rect 624 -122 654 -96
rect 720 -122 750 -96
rect 816 -122 846 -96
rect 144 -154 846 -122
rect 466 -196 524 -154
rect -14 -206 524 -196
rect -14 -240 2 -206
rect 36 -232 524 -206
rect 36 -240 52 -232
rect -14 -254 52 -240
rect 652 -284 724 -274
rect 652 -324 668 -284
rect 708 -324 724 -284
rect 260 -334 332 -324
rect 652 -334 724 -324
rect 1100 -294 1168 -284
rect 1100 -330 1116 -294
rect 1152 -330 1168 -294
rect 260 -374 276 -334
rect 316 -374 332 -334
rect 260 -384 332 -374
rect 284 -454 322 -384
rect 668 -454 706 -334
rect 1100 -368 1168 -330
rect 1100 -404 1116 -368
rect 1152 -404 1168 -368
rect 1100 -442 1168 -404
rect 144 -484 462 -454
rect 144 -510 174 -484
rect 240 -510 270 -484
rect 336 -510 366 -484
rect 432 -510 462 -484
rect 528 -484 846 -454
rect 528 -510 558 -484
rect 624 -510 654 -484
rect 720 -510 750 -484
rect 816 -510 846 -484
rect 1100 -478 1116 -442
rect 1152 -462 1168 -442
rect 2396 -204 2470 -188
rect 2396 -238 2410 -204
rect 2446 -238 2470 -204
rect 2396 -276 2470 -238
rect 2396 -310 2410 -276
rect 2446 -310 2470 -276
rect 2396 -326 2470 -310
rect 1276 -462 1306 -446
rect 1372 -462 1402 -446
rect 1152 -478 1402 -462
rect 1100 -492 1402 -478
rect 1598 -462 1628 -446
rect 1694 -462 1724 -446
rect 1598 -492 1724 -462
rect 1690 -558 1724 -492
rect 1658 -568 1724 -558
rect 1658 -602 1674 -568
rect 1708 -602 1724 -568
rect 1658 -612 1724 -602
rect 1598 -776 1628 -750
rect 1694 -776 1724 -612
rect 1790 -462 1820 -446
rect 1886 -462 1916 -446
rect 1790 -492 1916 -462
rect 2112 -462 2142 -446
rect 2208 -462 2238 -446
rect 2112 -492 2238 -462
rect 1790 -626 1824 -492
rect 1790 -636 2050 -626
rect 1790 -670 1808 -636
rect 1842 -670 2050 -636
rect 2204 -668 2238 -492
rect 1790 -680 2050 -670
rect 1790 -776 1820 -680
rect 1886 -776 1916 -750
rect 144 -938 174 -910
rect 240 -938 270 -910
rect 336 -938 366 -910
rect 432 -938 462 -910
rect 528 -938 558 -910
rect 624 -938 654 -910
rect 720 -938 750 -910
rect 816 -938 846 -910
rect -6 -1004 60 -994
rect -6 -1038 10 -1004
rect 44 -1014 60 -1004
rect 44 -1038 846 -1014
rect -6 -1044 846 -1038
rect -6 -1048 60 -1044
rect 144 -1070 174 -1044
rect 240 -1070 270 -1044
rect 336 -1070 366 -1044
rect 432 -1070 462 -1044
rect 528 -1070 558 -1044
rect 624 -1070 654 -1044
rect 720 -1070 750 -1044
rect 816 -1070 846 -1044
rect 144 -1196 174 -1170
rect 240 -1196 270 -1170
rect 336 -1196 366 -1170
rect 432 -1196 462 -1170
rect 528 -1196 558 -1170
rect 624 -1196 654 -1170
rect 720 -1196 750 -1170
rect 816 -1196 846 -1170
rect 1994 -796 2050 -680
rect 2108 -684 2238 -668
rect 2108 -720 2118 -684
rect 2154 -720 2192 -684
rect 2228 -720 2238 -684
rect 2108 -736 2238 -720
rect 1994 -852 2466 -796
rect 1598 -1244 1628 -1176
rect 1694 -1202 1724 -1176
rect 1790 -1202 1820 -1176
rect 1886 -1244 1916 -1176
rect 1440 -1254 1916 -1244
rect 1440 -1288 1456 -1254
rect 1490 -1274 1916 -1254
rect 1490 -1288 1506 -1274
rect 1440 -1298 1506 -1288
<< polycont >>
rect 2 -240 36 -206
rect 668 -324 708 -284
rect 1116 -330 1152 -294
rect 276 -374 316 -334
rect 1116 -404 1152 -368
rect 1116 -478 1152 -442
rect 2410 -238 2446 -204
rect 2410 -310 2446 -276
rect 1674 -602 1708 -568
rect 1808 -670 1842 -636
rect 10 -1038 44 -1004
rect 2118 -720 2154 -684
rect 2192 -720 2228 -684
rect 1456 -1288 1490 -1254
<< locali >>
rect -686 3918 4192 3974
rect -686 3844 -262 3918
rect -188 3844 286 3918
rect 360 3844 834 3918
rect 908 3844 1382 3918
rect 1456 3844 1930 3918
rect 2004 3844 2460 3918
rect 2534 3844 3008 3918
rect 3082 3844 3558 3918
rect 3632 3844 4192 3918
rect -686 3776 4192 3844
rect -686 3442 -488 3776
rect -686 3368 -628 3442
rect -554 3368 -488 3442
rect -686 2968 -488 3368
rect -686 2894 -628 2968
rect -554 2894 -488 2968
rect -686 2494 -488 2894
rect -686 2420 -628 2494
rect -554 2420 -488 2494
rect -686 2020 -488 2420
rect -686 1946 -628 2020
rect -554 1946 -488 2020
rect -686 1546 -488 1946
rect -686 1472 -628 1546
rect -554 1472 -488 1546
rect -686 1072 -488 1472
rect -686 998 -628 1072
rect -554 998 -488 1072
rect -686 604 -488 998
rect 3994 3374 4192 3776
rect 3994 3300 4054 3374
rect 4128 3300 4192 3374
rect 3994 2900 4192 3300
rect 3994 2826 4054 2900
rect 4128 2826 4192 2900
rect 3994 2426 4192 2826
rect 3994 2352 4054 2426
rect 4128 2352 4192 2426
rect 3994 1950 4192 2352
rect 3994 1876 4054 1950
rect 4128 1876 4192 1950
rect 3994 1474 4192 1876
rect 3994 1400 4054 1474
rect 4128 1400 4192 1474
rect 3994 1000 4192 1400
rect 3994 926 4054 1000
rect 4128 926 4192 1000
rect 3994 604 4192 926
rect -686 598 566 604
rect -686 524 -628 598
rect -554 564 566 598
rect -554 524 -372 564
rect -686 498 -372 524
rect -308 498 -264 564
rect -200 498 -156 564
rect -92 498 -48 564
rect 16 498 60 564
rect 124 498 168 564
rect 232 498 276 564
rect 340 498 384 564
rect 448 498 492 564
rect 556 498 566 564
rect 2996 564 4192 604
rect -686 476 566 498
rect 938 506 1050 522
rect -686 -88 -488 476
rect 938 440 950 506
rect 1032 440 1050 506
rect 938 420 1050 440
rect 82 100 938 108
rect 82 66 112 100
rect 146 66 196 100
rect 230 66 280 100
rect 314 66 364 100
rect 398 66 448 100
rect 482 66 532 100
rect 566 66 616 100
rect 650 66 700 100
rect 734 66 784 100
rect 818 66 874 100
rect 908 66 938 100
rect 82 60 938 66
rect -686 -162 -628 -88
rect -554 -162 -488 -88
rect 94 42 896 60
rect 94 -8 128 42
rect 94 -100 128 -84
rect 190 -8 224 8
rect -686 -614 -488 -162
rect 190 -160 224 -84
rect 286 -8 320 42
rect 286 -100 320 -84
rect 382 -8 416 8
rect 382 -160 416 -84
rect 478 -8 512 42
rect 478 -100 512 -84
rect 574 -8 608 8
rect 190 -194 416 -160
rect 574 -160 608 -84
rect 670 -8 704 42
rect 670 -100 704 -84
rect 766 -8 800 8
rect 766 -160 800 -84
rect 862 -8 896 42
rect 862 -100 896 -84
rect 574 -194 800 -160
rect -14 -206 52 -196
rect -14 -240 2 -206
rect 36 -240 52 -206
rect -14 -254 52 -240
rect -686 -688 -636 -614
rect -562 -688 -488 -614
rect -686 -1088 -488 -688
rect 6 -994 52 -254
rect 190 -418 224 -194
rect 260 -334 332 -324
rect 260 -374 276 -334
rect 316 -374 332 -334
rect 260 -384 332 -374
rect 368 -364 416 -358
rect 368 -400 374 -364
rect 410 -400 416 -364
rect 368 -418 416 -400
rect 190 -452 416 -418
rect 94 -522 128 -506
rect 94 -948 128 -898
rect 190 -522 224 -452
rect 190 -914 224 -898
rect 286 -522 320 -506
rect 286 -948 320 -898
rect 382 -522 416 -452
rect 574 -416 608 -194
rect 652 -284 724 -274
rect 652 -324 668 -284
rect 708 -324 724 -284
rect 652 -334 724 -324
rect 974 -416 1050 420
rect 574 -450 1050 -416
rect 382 -914 416 -898
rect 478 -522 512 -506
rect 478 -948 512 -898
rect 574 -522 608 -450
rect 574 -914 608 -898
rect 670 -522 704 -506
rect 670 -948 704 -898
rect 766 -522 800 -450
rect 766 -914 800 -898
rect 862 -522 896 -506
rect 974 -540 1050 -450
rect 1096 508 1222 524
rect 1096 442 1134 508
rect 1204 442 1222 508
rect 2996 498 3008 564
rect 3072 498 3116 564
rect 3180 498 3224 564
rect 3288 498 3336 564
rect 3400 498 3444 564
rect 3508 498 3552 564
rect 3616 498 3660 564
rect 3724 498 3768 564
rect 3832 498 3876 564
rect 3940 526 4192 564
rect 3940 498 4052 526
rect 2996 474 4052 498
rect 1096 420 1222 442
rect 3994 452 4052 474
rect 4126 452 4192 526
rect 1096 -294 1172 420
rect 2404 230 2952 250
rect 2404 194 2498 230
rect 2534 194 2574 230
rect 2610 194 2650 230
rect 2686 194 2726 230
rect 2762 194 2802 230
rect 2838 194 2878 230
rect 2914 194 2952 230
rect 2404 152 2952 194
rect 1382 110 2106 118
rect 1382 76 1420 110
rect 1454 76 1504 110
rect 1538 76 1588 110
rect 1622 76 1672 110
rect 1706 76 1756 110
rect 1790 76 1840 110
rect 1874 76 1924 110
rect 1958 76 2008 110
rect 2042 76 2106 110
rect 1382 70 2106 76
rect 1718 36 1808 70
rect 1096 -330 1116 -294
rect 1152 -330 1172 -294
rect 1096 -368 1172 -330
rect 1096 -404 1116 -368
rect 1152 -404 1172 -368
rect 1096 -442 1172 -404
rect 1096 -478 1116 -442
rect 1152 -478 1172 -442
rect 1096 -506 1172 -478
rect 1226 -8 1452 26
rect 1226 -58 1260 -8
rect 974 -552 1172 -540
rect 974 -588 1116 -552
rect 1152 -588 1172 -552
rect 1226 -568 1260 -434
rect 1322 -58 1356 -42
rect 1322 -500 1356 -434
rect 1418 -58 1452 -8
rect 1418 -450 1452 -434
rect 1548 2 1966 36
rect 1548 -58 1582 2
rect 1548 -450 1582 -434
rect 1644 -58 1678 -42
rect 1644 -500 1678 -434
rect 1740 -58 1774 2
rect 1740 -450 1774 -434
rect 1836 -58 1870 -42
rect 1322 -534 1678 -500
rect 1836 -500 1870 -434
rect 1932 -58 1966 2
rect 1932 -450 1966 -434
rect 2062 -8 2288 26
rect 2062 -58 2096 -8
rect 2062 -450 2096 -434
rect 2158 -58 2192 -42
rect 2158 -500 2192 -434
rect 1836 -534 2192 -500
rect 2254 -58 2288 -8
rect 2288 -204 2452 -188
rect 2288 -238 2410 -204
rect 2446 -238 2452 -204
rect 2288 -276 2452 -238
rect 2288 -310 2410 -276
rect 2446 -310 2452 -276
rect 2786 -234 2846 -224
rect 2786 -236 2860 -234
rect 2786 -272 2792 -236
rect 2828 -272 2860 -236
rect 2786 -284 2846 -272
rect 2288 -326 2452 -310
rect 2254 -568 2288 -434
rect 974 -628 1172 -588
rect 1210 -602 1622 -568
rect 1658 -602 1674 -568
rect 1708 -602 2300 -568
rect 2338 -582 2436 -514
rect 974 -664 1116 -628
rect 1152 -664 1172 -628
rect 974 -702 1172 -664
rect 1588 -636 1622 -602
rect 1588 -670 1808 -636
rect 1842 -670 1858 -636
rect 974 -738 1116 -702
rect 1152 -738 1172 -702
rect 974 -750 1172 -738
rect 862 -948 896 -898
rect 94 -984 896 -948
rect -6 -1004 60 -994
rect -6 -1038 10 -1004
rect 44 -1038 60 -1004
rect -6 -1048 60 -1038
rect -686 -1162 -636 -1088
rect -562 -1162 -488 -1088
rect -686 -1222 -488 -1162
rect 94 -1082 128 -984
rect 94 -1174 128 -1158
rect 190 -1082 224 -1064
rect -686 -1256 -670 -1222
rect -636 -1256 -598 -1222
rect -564 -1256 -526 -1222
rect -492 -1256 -488 -1222
rect -686 -1294 -488 -1256
rect -686 -1328 -670 -1294
rect -636 -1328 -598 -1294
rect -564 -1328 -526 -1294
rect -492 -1328 -488 -1294
rect -686 -1366 -488 -1328
rect 190 -1316 224 -1158
rect 286 -1082 320 -984
rect 286 -1174 320 -1158
rect 382 -1082 416 -1066
rect 382 -1316 416 -1158
rect 478 -1082 512 -984
rect 478 -1174 512 -1158
rect 574 -1082 608 -1066
rect 574 -1316 608 -1158
rect 670 -1082 704 -984
rect 670 -1174 704 -1158
rect 766 -1082 800 -1066
rect 766 -1316 800 -1158
rect 862 -1082 896 -984
rect 862 -1174 896 -1158
rect 974 -858 1050 -834
rect 974 -894 994 -858
rect 1030 -894 1050 -858
rect 974 -932 1050 -894
rect 974 -968 994 -932
rect 1030 -968 1050 -932
rect 974 -1006 1050 -968
rect 974 -1042 994 -1006
rect 1030 -1042 1050 -1006
rect 190 -1330 800 -1316
rect -686 -1400 -670 -1366
rect -636 -1400 -598 -1366
rect -564 -1400 -526 -1366
rect -492 -1400 -488 -1366
rect 76 -1332 894 -1330
rect 76 -1368 100 -1332
rect 136 -1368 218 -1332
rect 254 -1368 336 -1332
rect 372 -1368 454 -1332
rect 490 -1368 572 -1332
rect 608 -1368 690 -1332
rect 726 -1368 808 -1332
rect 844 -1368 894 -1332
rect 76 -1372 894 -1368
rect -686 -1438 -488 -1400
rect -686 -1472 -670 -1438
rect -636 -1472 -598 -1438
rect -564 -1472 -526 -1438
rect -492 -1472 -488 -1438
rect -686 -1510 -488 -1472
rect -686 -1544 -672 -1510
rect -638 -1544 -600 -1510
rect -566 -1544 -528 -1510
rect -494 -1544 -488 -1510
rect -686 -1700 -488 -1544
rect 974 -1586 1050 -1042
rect 954 -1602 1050 -1586
rect 954 -1668 968 -1602
rect 1042 -1668 1050 -1602
rect 954 -1680 1050 -1668
rect 1096 -1586 1172 -750
rect 1548 -788 1582 -772
rect 1440 -1254 1506 -1244
rect 1440 -1288 1456 -1254
rect 1490 -1288 1506 -1254
rect 1548 -1288 1582 -1164
rect 1644 -788 1678 -670
rect 1902 -704 1936 -602
rect 1836 -738 1936 -704
rect 2112 -684 2234 -668
rect 2112 -720 2118 -684
rect 2154 -720 2192 -684
rect 2228 -720 2234 -684
rect 2112 -736 2234 -720
rect 1644 -1180 1678 -1164
rect 1740 -788 1774 -772
rect 1740 -1288 1774 -1164
rect 1836 -788 1870 -738
rect 1836 -1180 1870 -1164
rect 1932 -788 1966 -772
rect 2338 -908 2406 -582
rect 2790 -824 2850 -814
rect 2790 -826 2862 -824
rect 2790 -862 2796 -826
rect 2832 -862 2862 -826
rect 2790 -874 2850 -862
rect 1932 -1288 1966 -1164
rect 2268 -976 2406 -908
rect 1440 -1298 1506 -1288
rect 1542 -1324 1566 -1288
rect 1602 -1324 1658 -1288
rect 1694 -1324 1750 -1288
rect 1786 -1324 1842 -1288
rect 1878 -1324 1934 -1288
rect 1970 -1324 1994 -1288
rect 1542 -1326 1994 -1324
rect 2268 -1326 2348 -976
rect 2896 -1248 2952 152
rect 2406 -1286 2952 -1248
rect 3994 -86 4192 452
rect 3994 -160 4052 -86
rect 4126 -160 4192 -86
rect 3994 -560 4192 -160
rect 3994 -634 4052 -560
rect 4126 -634 4192 -560
rect 3994 -1034 4192 -634
rect 3994 -1108 4052 -1034
rect 4126 -1108 4192 -1034
rect 3994 -1222 4192 -1108
rect 3994 -1256 4008 -1222
rect 4042 -1256 4080 -1222
rect 4114 -1256 4152 -1222
rect 4186 -1256 4192 -1222
rect 3994 -1294 4192 -1256
rect 2268 -1344 2632 -1326
rect 2268 -1346 2350 -1344
rect 2268 -1382 2276 -1346
rect 2312 -1380 2350 -1346
rect 2386 -1380 2430 -1344
rect 2466 -1380 2510 -1344
rect 2546 -1380 2590 -1344
rect 2626 -1380 2632 -1344
rect 2312 -1382 2632 -1380
rect 2268 -1396 2632 -1382
rect 3994 -1328 4008 -1294
rect 4042 -1328 4080 -1294
rect 4114 -1328 4152 -1294
rect 4186 -1328 4192 -1294
rect 3994 -1366 4192 -1328
rect 3994 -1400 4008 -1366
rect 4042 -1400 4080 -1366
rect 4114 -1400 4152 -1366
rect 4186 -1400 4192 -1366
rect 3994 -1438 4192 -1400
rect 3994 -1472 4008 -1438
rect 4042 -1472 4080 -1438
rect 4114 -1472 4152 -1438
rect 4186 -1472 4192 -1438
rect 3994 -1510 4192 -1472
rect 3994 -1544 4008 -1510
rect 4042 -1544 4080 -1510
rect 4114 -1544 4152 -1510
rect 4186 -1544 4192 -1510
rect 1096 -1602 1214 -1586
rect 1096 -1668 1120 -1602
rect 1196 -1668 1214 -1602
rect 1096 -1680 1214 -1668
rect 3994 -1698 4192 -1544
rect -686 -1740 526 -1700
rect -686 -1814 -622 -1740
rect -548 -1806 -354 -1740
rect -290 -1806 -220 -1740
rect -156 -1806 -86 -1740
rect -22 -1806 22 -1740
rect 86 -1806 130 -1740
rect 194 -1806 238 -1740
rect 302 -1806 346 -1740
rect 410 -1806 454 -1740
rect 518 -1806 526 -1740
rect -548 -1814 526 -1806
rect -686 -1828 526 -1814
rect 3006 -1738 4192 -1698
rect 3006 -1804 3028 -1738
rect 3092 -1804 3136 -1738
rect 3200 -1804 3244 -1738
rect 3308 -1804 3356 -1738
rect 3420 -1804 3464 -1738
rect 3528 -1804 3572 -1738
rect 3642 -1804 3686 -1738
rect 3756 -1804 3800 -1738
rect 3870 -1770 4192 -1738
rect 3870 -1804 4052 -1770
rect 3006 -1826 4052 -1804
rect -686 -2214 -488 -1828
rect -686 -2288 -622 -2214
rect -548 -2288 -488 -2214
rect -686 -2688 -488 -2288
rect -686 -2762 -622 -2688
rect -548 -2762 -488 -2688
rect -686 -3164 -488 -2762
rect -686 -3238 -622 -3164
rect -548 -3238 -488 -3164
rect -686 -3638 -488 -3238
rect -686 -3712 -622 -3638
rect -548 -3712 -488 -3638
rect -686 -4112 -488 -3712
rect -686 -4186 -622 -4112
rect -548 -4186 -488 -4112
rect -686 -4586 -488 -4186
rect -686 -4660 -622 -4586
rect -548 -4660 -488 -4586
rect -686 -4932 -488 -4660
rect 3994 -1844 4052 -1826
rect 4126 -1844 4192 -1770
rect 3994 -2244 4192 -1844
rect 3994 -2318 4052 -2244
rect 4126 -2318 4192 -2244
rect 3994 -2718 4192 -2318
rect 3994 -2792 4052 -2718
rect 4126 -2792 4192 -2718
rect 3994 -3192 4192 -2792
rect 3994 -3266 4052 -3192
rect 4126 -3266 4192 -3192
rect 3994 -3666 4192 -3266
rect 3994 -3740 4052 -3666
rect 4126 -3740 4192 -3666
rect 3994 -4140 4192 -3740
rect 3994 -4214 4052 -4140
rect 4126 -4214 4192 -4140
rect 3994 -4614 4192 -4214
rect 3994 -4688 4054 -4614
rect 4128 -4688 4192 -4614
rect 3994 -4932 4192 -4688
rect -686 -5000 4192 -4932
rect -686 -5074 -92 -5000
rect -18 -5074 456 -5000
rect 530 -5074 1004 -5000
rect 1078 -5074 1552 -5000
rect 1626 -5074 2100 -5000
rect 2174 -5074 2648 -5000
rect 2722 -5074 3198 -5000
rect 3272 -5074 4192 -5000
rect -686 -5130 4192 -5074
<< viali >>
rect -372 498 -308 564
rect -264 498 -200 564
rect -156 498 -92 564
rect -48 498 16 564
rect 60 498 124 564
rect 168 498 232 564
rect 276 498 340 564
rect 384 498 448 564
rect 492 498 556 564
rect 950 440 1032 506
rect 112 66 146 100
rect 196 66 230 100
rect 280 66 314 100
rect 364 66 398 100
rect 448 66 482 100
rect 532 66 566 100
rect 616 66 650 100
rect 700 66 734 100
rect 784 66 818 100
rect 874 66 908 100
rect 276 -374 316 -334
rect 374 -400 410 -364
rect 668 -324 708 -284
rect 1134 442 1204 508
rect 3008 498 3072 564
rect 3116 498 3180 564
rect 3224 498 3288 564
rect 3336 498 3400 564
rect 3444 498 3508 564
rect 3552 498 3616 564
rect 3660 498 3724 564
rect 3768 498 3832 564
rect 3876 498 3940 564
rect 2498 194 2534 230
rect 2574 194 2610 230
rect 2650 194 2686 230
rect 2726 194 2762 230
rect 2802 194 2838 230
rect 2878 194 2914 230
rect 1420 76 1454 110
rect 1504 76 1538 110
rect 1588 76 1622 110
rect 1672 76 1706 110
rect 1756 76 1790 110
rect 1840 76 1874 110
rect 1924 76 1958 110
rect 2008 76 2042 110
rect 1116 -330 1152 -294
rect 1116 -404 1152 -368
rect 1116 -478 1152 -442
rect 1116 -588 1152 -552
rect 2410 -238 2446 -204
rect 2410 -310 2446 -276
rect 2792 -272 2828 -236
rect 1116 -664 1152 -628
rect 1116 -738 1152 -702
rect -670 -1256 -636 -1222
rect -598 -1256 -564 -1222
rect -526 -1256 -492 -1222
rect -670 -1328 -636 -1294
rect -598 -1328 -564 -1294
rect -526 -1328 -492 -1294
rect 994 -894 1030 -858
rect 994 -968 1030 -932
rect 994 -1042 1030 -1006
rect -670 -1400 -636 -1366
rect -598 -1400 -564 -1366
rect -526 -1400 -492 -1366
rect 100 -1368 136 -1332
rect 218 -1368 254 -1332
rect 336 -1368 372 -1332
rect 454 -1368 490 -1332
rect 572 -1368 608 -1332
rect 690 -1368 726 -1332
rect 808 -1368 844 -1332
rect -670 -1472 -636 -1438
rect -598 -1472 -564 -1438
rect -526 -1472 -492 -1438
rect -672 -1544 -638 -1510
rect -600 -1544 -566 -1510
rect -528 -1544 -494 -1510
rect 968 -1668 1042 -1602
rect 2118 -720 2154 -684
rect 2192 -720 2228 -684
rect 2796 -862 2832 -826
rect 1566 -1324 1602 -1288
rect 1658 -1324 1694 -1288
rect 1750 -1324 1786 -1288
rect 1842 -1324 1878 -1288
rect 1934 -1324 1970 -1288
rect 4008 -1256 4042 -1222
rect 4080 -1256 4114 -1222
rect 4152 -1256 4186 -1222
rect 2276 -1382 2312 -1346
rect 2350 -1380 2386 -1344
rect 2430 -1380 2466 -1344
rect 2510 -1380 2546 -1344
rect 2590 -1380 2626 -1344
rect 4008 -1328 4042 -1294
rect 4080 -1328 4114 -1294
rect 4152 -1328 4186 -1294
rect 4008 -1400 4042 -1366
rect 4080 -1400 4114 -1366
rect 4152 -1400 4186 -1366
rect 4008 -1472 4042 -1438
rect 4080 -1472 4114 -1438
rect 4152 -1472 4186 -1438
rect 4008 -1544 4042 -1510
rect 4080 -1544 4114 -1510
rect 4152 -1544 4186 -1510
rect 1120 -1668 1196 -1602
rect -354 -1806 -290 -1740
rect -220 -1806 -156 -1740
rect -86 -1806 -22 -1740
rect 22 -1806 86 -1740
rect 130 -1806 194 -1740
rect 238 -1806 302 -1740
rect 346 -1806 410 -1740
rect 454 -1806 518 -1740
rect 3028 -1804 3092 -1738
rect 3136 -1804 3200 -1738
rect 3244 -1804 3308 -1738
rect 3356 -1804 3420 -1738
rect 3464 -1804 3528 -1738
rect 3572 -1804 3642 -1738
rect 3686 -1804 3756 -1738
rect 3800 -1804 3870 -1738
<< metal1 >>
rect -488 564 566 604
rect -488 498 -372 564
rect -308 498 -264 564
rect -200 498 -156 564
rect -92 498 -48 564
rect 16 498 60 564
rect 124 498 168 564
rect 232 498 276 564
rect 340 498 384 564
rect 448 498 492 564
rect 556 498 566 564
rect 2996 564 3974 604
rect -488 476 566 498
rect 938 506 1050 522
rect 938 440 950 506
rect 1032 440 1050 506
rect 938 420 1050 440
rect 1110 508 1222 524
rect 1110 442 1134 508
rect 1204 442 1222 508
rect 2996 498 3008 564
rect 3076 498 3116 564
rect 3184 498 3224 564
rect 3292 498 3336 564
rect 3400 498 3444 564
rect 3508 498 3552 564
rect 3616 498 3660 564
rect 3724 498 3768 564
rect 3832 498 3876 564
rect 3940 498 3974 564
rect 2996 476 3974 498
rect 1110 430 1222 442
rect -838 230 4360 392
rect -838 194 2498 230
rect 2534 194 2574 230
rect 2610 194 2650 230
rect 2686 194 2726 230
rect 2762 194 2802 230
rect 2838 194 2878 230
rect 2914 194 4360 230
rect -838 162 4360 194
rect 82 100 938 162
rect 82 66 112 100
rect 146 66 196 100
rect 230 66 280 100
rect 314 66 364 100
rect 398 66 448 100
rect 482 66 532 100
rect 566 66 616 100
rect 650 66 700 100
rect 734 66 784 100
rect 818 66 874 100
rect 908 66 938 100
rect 1382 110 2106 162
rect 1382 76 1420 110
rect 1454 76 1504 110
rect 1538 76 1588 110
rect 1622 76 1672 110
rect 1706 76 1756 110
rect 1790 76 1840 110
rect 1874 76 1924 110
rect 1958 76 2008 110
rect 2042 76 2106 110
rect 1382 70 2106 76
rect 82 60 938 66
rect 2396 -204 2452 -188
rect 2396 -238 2410 -204
rect 2446 -238 2452 -204
rect -838 -284 724 -268
rect 2396 -276 2452 -238
rect -838 -296 668 -284
rect 652 -324 668 -296
rect 708 -324 724 -284
rect -838 -334 332 -324
rect 652 -334 724 -324
rect 1104 -294 1164 -284
rect 1104 -330 1116 -294
rect 1152 -330 1164 -294
rect 2396 -310 2410 -276
rect 2446 -310 2452 -276
rect 2786 -236 2846 -224
rect 2786 -272 2792 -236
rect 2828 -272 2846 -236
rect 2786 -284 2846 -272
rect 2396 -328 2452 -310
rect -838 -352 276 -334
rect 260 -374 276 -352
rect 316 -374 332 -334
rect 260 -384 332 -374
rect 362 -362 416 -358
rect 1104 -362 1164 -330
rect 362 -364 1164 -362
rect 362 -376 374 -364
rect 360 -400 374 -376
rect 410 -368 1164 -364
rect 410 -400 1116 -368
rect 360 -404 1116 -400
rect 1152 -404 1164 -368
rect 360 -414 1164 -404
rect 974 -858 1050 -414
rect 1104 -442 1164 -414
rect 1104 -478 1116 -442
rect 1152 -478 1164 -442
rect 1104 -484 1164 -478
rect 1104 -552 1164 -546
rect 1104 -588 1116 -552
rect 1152 -588 1164 -552
rect 1104 -628 1164 -588
rect 1104 -664 1116 -628
rect 1152 -664 1164 -628
rect 1104 -700 1164 -664
rect 2108 -684 2238 -668
rect 2108 -700 2118 -684
rect 1104 -702 2118 -700
rect 1104 -738 1116 -702
rect 1152 -720 2118 -702
rect 2154 -720 2192 -684
rect 2228 -720 2238 -684
rect 1152 -736 2238 -720
rect 1152 -738 1164 -736
rect 1104 -744 1164 -738
rect 974 -894 994 -858
rect 1030 -894 1050 -858
rect 2790 -826 2850 -814
rect 2790 -862 2796 -826
rect 2832 -862 2850 -826
rect 2790 -874 2850 -862
rect 974 -932 1050 -894
rect 974 -968 994 -932
rect 1030 -968 1050 -932
rect 974 -1006 1050 -968
rect 974 -1042 994 -1006
rect 1030 -1042 1050 -1006
rect 974 -1070 1050 -1042
rect -686 -1222 -486 -1202
rect -686 -1256 -670 -1222
rect -636 -1256 -598 -1222
rect -564 -1256 -526 -1222
rect -492 -1256 -486 -1222
rect -686 -1294 -486 -1256
rect 3994 -1222 4192 -1202
rect 3994 -1256 4008 -1222
rect 4042 -1256 4080 -1222
rect 4114 -1256 4152 -1222
rect 4186 -1256 4192 -1222
rect -686 -1326 -670 -1294
rect -838 -1328 -670 -1326
rect -636 -1328 -598 -1294
rect -564 -1328 -526 -1294
rect -492 -1326 -486 -1294
rect 1542 -1288 1994 -1282
rect 1542 -1324 1566 -1288
rect 1602 -1324 1658 -1288
rect 1694 -1324 1750 -1288
rect 1786 -1324 1842 -1288
rect 1878 -1324 1934 -1288
rect 1970 -1324 1994 -1288
rect 1542 -1326 1994 -1324
rect 3994 -1294 4192 -1256
rect 3994 -1326 4008 -1294
rect -492 -1328 4008 -1326
rect 4042 -1328 4080 -1294
rect 4114 -1328 4152 -1294
rect 4186 -1326 4192 -1294
rect 4186 -1328 4360 -1326
rect -838 -1332 4360 -1328
rect -838 -1366 100 -1332
rect -838 -1400 -670 -1366
rect -636 -1400 -598 -1366
rect -564 -1400 -526 -1366
rect -492 -1368 100 -1366
rect 136 -1368 218 -1332
rect 254 -1368 336 -1332
rect 372 -1368 454 -1332
rect 490 -1368 572 -1332
rect 608 -1368 690 -1332
rect 726 -1368 808 -1332
rect 844 -1344 4360 -1332
rect 844 -1346 2350 -1344
rect 844 -1368 2276 -1346
rect -492 -1382 2276 -1368
rect 2312 -1380 2350 -1346
rect 2386 -1380 2430 -1344
rect 2466 -1380 2510 -1344
rect 2546 -1380 2590 -1344
rect 2626 -1366 4360 -1344
rect 2626 -1380 4008 -1366
rect 2312 -1382 4008 -1380
rect -492 -1400 4008 -1382
rect 4042 -1400 4080 -1366
rect 4114 -1400 4152 -1366
rect 4186 -1400 4360 -1366
rect -838 -1438 4360 -1400
rect -838 -1472 -670 -1438
rect -636 -1472 -598 -1438
rect -564 -1472 -526 -1438
rect -492 -1472 4008 -1438
rect 4042 -1472 4080 -1438
rect 4114 -1472 4152 -1438
rect 4186 -1472 4360 -1438
rect -838 -1510 4360 -1472
rect -838 -1544 -672 -1510
rect -638 -1544 -600 -1510
rect -566 -1544 -528 -1510
rect -494 -1544 4008 -1510
rect 4042 -1544 4080 -1510
rect 4114 -1544 4152 -1510
rect 4186 -1544 4360 -1510
rect -838 -1558 4360 -1544
rect 942 -1602 1050 -1586
rect 942 -1668 968 -1602
rect 1042 -1668 1050 -1602
rect 942 -1680 1050 -1668
rect 1110 -1602 1214 -1586
rect 1110 -1668 1120 -1602
rect 1196 -1668 1214 -1602
rect 1110 -1680 1214 -1668
rect -380 -1740 526 -1700
rect -380 -1806 -354 -1740
rect -290 -1806 -220 -1740
rect -156 -1806 -86 -1740
rect -22 -1806 22 -1740
rect 86 -1806 130 -1740
rect 194 -1806 238 -1740
rect 302 -1806 346 -1740
rect 410 -1806 454 -1740
rect 518 -1806 526 -1740
rect -380 -1828 526 -1806
rect 3006 -1738 3994 -1698
rect 3006 -1804 3028 -1738
rect 3096 -1804 3136 -1738
rect 3204 -1804 3244 -1738
rect 3312 -1804 3356 -1738
rect 3420 -1804 3464 -1738
rect 3528 -1804 3572 -1738
rect 3642 -1804 3686 -1738
rect 3756 -1804 3800 -1738
rect 3870 -1804 3994 -1738
rect 3006 -1826 3994 -1804
<< via1 >>
rect -372 498 -308 564
rect -264 498 -200 564
rect -156 498 -92 564
rect -48 498 16 564
rect 60 498 124 564
rect 168 498 232 564
rect 276 498 340 564
rect 384 498 448 564
rect 492 498 556 564
rect 950 440 1032 506
rect 1134 442 1204 508
rect 3008 498 3072 564
rect 3072 498 3076 564
rect 3116 498 3180 564
rect 3180 498 3184 564
rect 3224 498 3288 564
rect 3288 498 3292 564
rect 3336 498 3400 564
rect 3444 498 3508 564
rect 3552 498 3616 564
rect 3660 498 3724 564
rect 3768 498 3832 564
rect 3876 498 3940 564
rect 968 -1668 1042 -1602
rect 1120 -1668 1196 -1602
rect -354 -1806 -290 -1740
rect -220 -1806 -156 -1740
rect -86 -1806 -22 -1740
rect 22 -1806 86 -1740
rect 130 -1806 194 -1740
rect 238 -1806 302 -1740
rect 346 -1806 410 -1740
rect 454 -1806 518 -1740
rect 3028 -1804 3092 -1738
rect 3092 -1804 3096 -1738
rect 3136 -1804 3200 -1738
rect 3200 -1804 3204 -1738
rect 3244 -1804 3308 -1738
rect 3308 -1804 3312 -1738
rect 3356 -1804 3420 -1738
rect 3464 -1804 3528 -1738
rect 3572 -1804 3642 -1738
rect 3686 -1804 3756 -1738
rect 3800 -1804 3870 -1738
<< metal2 >>
rect -488 564 566 604
rect -488 498 -372 564
rect -308 498 -264 564
rect -200 498 -156 564
rect -92 498 -48 564
rect 16 498 60 564
rect 124 498 168 564
rect 232 498 276 564
rect 340 498 384 564
rect 448 498 492 564
rect 556 498 566 564
rect 2996 564 3974 604
rect -488 476 566 498
rect 938 506 1050 522
rect 938 440 950 506
rect 1032 440 1050 506
rect 938 420 1050 440
rect 1110 508 1222 524
rect 1110 442 1134 508
rect 1204 442 1222 508
rect 2996 498 3008 564
rect 3076 498 3116 564
rect 3184 498 3224 564
rect 3292 498 3336 564
rect 3400 498 3444 564
rect 3508 498 3552 564
rect 3616 498 3660 564
rect 3724 498 3768 564
rect 3832 498 3876 564
rect 3940 498 3974 564
rect 2996 476 3974 498
rect 1110 430 1222 442
rect 942 -1602 1050 -1586
rect 942 -1668 968 -1602
rect 1042 -1668 1050 -1602
rect 942 -1680 1050 -1668
rect 1110 -1602 1214 -1586
rect 1110 -1668 1120 -1602
rect 1196 -1668 1214 -1602
rect 1110 -1680 1214 -1668
rect -380 -1740 526 -1700
rect -380 -1806 -354 -1740
rect -290 -1806 -220 -1740
rect -156 -1806 -86 -1740
rect -22 -1806 22 -1740
rect 86 -1806 130 -1740
rect 194 -1806 238 -1740
rect 302 -1806 346 -1740
rect 410 -1806 454 -1740
rect 518 -1806 526 -1740
rect -380 -1828 526 -1806
rect 3006 -1738 3994 -1698
rect 3006 -1804 3028 -1738
rect 3096 -1804 3136 -1738
rect 3204 -1804 3244 -1738
rect 3312 -1804 3356 -1738
rect 3420 -1804 3464 -1738
rect 3528 -1804 3572 -1738
rect 3642 -1804 3686 -1738
rect 3756 -1804 3800 -1738
rect 3870 -1804 3994 -1738
rect 3006 -1826 3994 -1804
<< via2 >>
rect -372 498 -308 564
rect -264 498 -200 564
rect -156 498 -92 564
rect -48 498 16 564
rect 60 498 124 564
rect 168 498 232 564
rect 276 498 340 564
rect 384 498 448 564
rect 492 498 556 564
rect 950 440 1032 506
rect 1134 442 1204 508
rect 3008 498 3076 564
rect 3116 498 3184 564
rect 3224 498 3292 564
rect 3336 498 3400 564
rect 3444 498 3508 564
rect 3552 498 3616 564
rect 3660 498 3724 564
rect 3768 498 3832 564
rect 3876 498 3940 564
rect 968 -1668 1042 -1602
rect 1120 -1668 1196 -1602
rect -354 -1806 -290 -1740
rect -220 -1806 -156 -1740
rect -86 -1806 -22 -1740
rect 22 -1806 86 -1740
rect 130 -1806 194 -1740
rect 238 -1806 302 -1740
rect 346 -1806 410 -1740
rect 454 -1806 518 -1740
rect 3028 -1804 3096 -1738
rect 3136 -1804 3204 -1738
rect 3244 -1804 3312 -1738
rect 3356 -1804 3420 -1738
rect 3464 -1804 3528 -1738
rect 3572 -1804 3642 -1738
rect 3686 -1804 3756 -1738
rect 3800 -1804 3870 -1738
<< metal3 >>
rect -372 604 -156 606
rect 3616 604 3940 606
rect -488 564 566 604
rect -488 498 -372 564
rect -308 498 -264 564
rect -200 498 -156 564
rect -92 498 -48 564
rect 16 498 60 564
rect 124 498 168 564
rect 232 498 276 564
rect 340 498 384 564
rect 448 498 492 564
rect 556 498 566 564
rect 2996 564 3974 604
rect -488 474 566 498
rect 938 506 1050 522
rect 938 440 950 506
rect 1032 440 1050 506
rect 938 420 1050 440
rect 1110 508 1222 524
rect 1110 442 1134 508
rect 1204 442 1222 508
rect 2996 498 3008 564
rect 3076 498 3116 564
rect 3184 498 3224 564
rect 3292 498 3336 564
rect 3400 498 3444 564
rect 3508 498 3552 564
rect 3616 498 3660 564
rect 3724 498 3768 564
rect 3832 498 3876 564
rect 3940 498 3974 564
rect 2996 474 3974 498
rect 1110 430 1222 442
rect 942 -1602 1050 -1586
rect 942 -1668 968 -1602
rect 1042 -1668 1050 -1602
rect 942 -1680 1050 -1668
rect 1110 -1602 1214 -1586
rect 1110 -1668 1120 -1602
rect 1196 -1668 1214 -1602
rect 1110 -1680 1214 -1668
rect -380 -1740 526 -1700
rect -380 -1806 -354 -1740
rect -290 -1806 -220 -1740
rect -156 -1806 -86 -1740
rect -22 -1806 22 -1740
rect 86 -1806 130 -1740
rect 194 -1806 238 -1740
rect 302 -1806 346 -1740
rect 410 -1806 454 -1740
rect 518 -1806 526 -1740
rect -380 -1828 526 -1806
rect 3006 -1738 3994 -1698
rect 3006 -1804 3028 -1738
rect 3096 -1804 3136 -1738
rect 3204 -1804 3244 -1738
rect 3312 -1804 3356 -1738
rect 3420 -1804 3464 -1738
rect 3528 -1804 3572 -1738
rect 3642 -1804 3686 -1738
rect 3756 -1804 3800 -1738
rect 3870 -1804 3994 -1738
rect 3006 -1828 3994 -1804
<< via3 >>
rect 950 440 1032 506
rect 1134 442 1204 508
rect 968 -1668 1042 -1602
rect 1120 -1668 1196 -1602
<< metal4 >>
rect 568 522 674 580
rect 2888 524 2992 640
rect 568 506 1050 522
rect 568 440 950 506
rect 1032 440 1050 506
rect 568 420 1050 440
rect 1110 508 2992 524
rect 1110 442 1134 508
rect 1204 442 2992 508
rect 1110 420 2992 442
rect 942 -1596 1050 -1586
rect 534 -1602 1050 -1596
rect 534 -1668 968 -1602
rect 1042 -1668 1050 -1602
rect 534 -1680 1050 -1668
rect 1110 -1596 1214 -1586
rect 1110 -1602 2960 -1596
rect 1110 -1668 1120 -1602
rect 1196 -1668 2960 -1602
rect 1110 -1680 2960 -1668
rect 534 -1832 640 -1680
rect 2854 -1830 2960 -1680
<< comment >>
rect 94 -58 126 -16
rect 290 -62 322 -20
rect 480 -64 512 -22
rect 672 -64 704 -22
rect 864 -62 896 -20
rect 1332 -350 1350 -146
rect 1554 -338 1574 -118
rect 1748 -366 1768 -146
rect 1942 -308 1962 -88
rect 2168 -350 2186 -146
rect 100 -752 132 -710
rect 288 -738 320 -696
rect 476 -736 508 -694
rect 680 -732 712 -690
rect 868 -724 900 -682
rect 1548 -1056 1576 -888
rect 1742 -1058 1770 -890
rect 1934 -1072 1962 -904
rect 192 -1140 224 -1098
rect 390 -1142 422 -1100
rect 578 -1140 610 -1098
rect 766 -1140 798 -1098
use adc_comp_buffer  adc_comp_buffer_0 ../adc_comp_buffer
timestamp 1662367448
transform 1 0 2448 0 1 -226
box -42 -326 408 452
use adc_comp_buffer  adc_comp_buffer_1
timestamp 1662367448
transform 1 0 2448 0 -1 -870
box -42 -326 408 452
use cap_64_92  cap_64_92_0
timestamp 1661518684
transform 1 0 1750 0 1 2134
box -2149 -1580 2210 1580
use cap_64_92  cap_64_92_1
timestamp 1661518684
transform 1 0 1717 0 -1 -3358
box -2149 -1580 2210 1580
<< labels >>
rlabel locali 1210 -602 1210 -568 7 bn
rlabel locali 2300 -602 2300 -568 3 bp
rlabel locali 2862 -862 2862 -824 3 outn
port 7 e
rlabel locali 2860 -272 2860 -234 3 outp
port 8 e
rlabel locali 574 -450 574 -418 7 on
rlabel locali 190 -450 190 -418 7 op
rlabel metal1 -838 -296 -838 -268 7 inp
port 5 w
rlabel metal1 -838 -352 -838 -324 7 inn
port 6 w
rlabel metal1 -838 -1484 -838 -1326 7 VSS
port 2 w
rlabel metal1 -838 162 -838 300 7 VDD
port 1 w
rlabel locali 1440 -1298 1440 -1244 7 nclk
port 10 w
rlabel locali -6 -1044 -6 -1014 7 clk
port 9 w
<< end >>
