* NGSPICE file created from adc_array_matrix_12bit.ext - technology: sky130A

.subckt adc_array_matrix_12bit_ext VDD VSS vcm sample sample_n row_n[0] row_n[1] row_n[2] row_n[3]
+ row_n[4] row_n[5] row_n[6] row_n[7] row_n[8] row_n[9] row_n[10] row_n[11] row_n[12] row_n[13] row_n[14]
+ row_n[15] rowon_n[0] rowon_n[1] rowon_n[2] rowon_n[3] rowon_n[4] rowon_n[5] rowon_n[6] rowon_n[7] rowon_n[8]
+ rowon_n[9] rowon_n[10] rowon_n[11] rowon_n[12] rowon_n[13] rowon_n[14] rowon_n[15] col_n[0] col_n[1] col_n[2]
+ col_n[3] col_n[4] col_n[5] col_n[6] col_n[7] col_n[8] col_n[9] col_n[10] col_n[11] col_n[12] col_n[13]
+ col_n[14] col_n[15] col_n[16] col_n[17] col_n[18] col_n[19] col_n[20] col_n[21] col_n[22] col_n[23] col_n[24]
+ col_n[25] col_n[26] col_n[27] col_n[28] col_n[29] col_n[30] col_n[31] en_bit_n[0] en_bit_n[1] en_bit_n[2] en_C0_n sw sw_n analog_in ctop rowoff_n[0] rowoff_n[1] rowoff_n[2]
+ rowoff_n[3] rowoff_n[4] rowoff_n[5] rowoff_n[6] rowoff_n[7] rowoff_n[8] rowoff_n[9] rowoff_n[10] rowoff_n[11]
+ rowoff_n[12] rowoff_n[13] rowoff_n[14] rowoff_n[15] col[0] col[1] col[2] col[3] col[4] col[5] col[6] col[7] col[8] col[9]
+ col[10] col[11] col[12] col[13] col[14] col[15] col[16] col[17] col[18] col[19] col[20] col[21] col[22]
+ col[23] col[24] col[25] col[26] col[27] col[28] col[29] col[30] col[31] 
X0 a_3970_15182# a_2475_15206# a_3878_15182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1 a_3878_9158# a_2275_9182# a_3970_9158# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2 VDD rowon_n[5] a_18938_7150# VDD sky130_fd_pr__pfet_01v8 ad=1.71672e+14p pd=1.45178e+09u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3 a_30986_7150# row_n[5] a_31478_7512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4 vcm a_2275_18218# a_32082_18194# VSS sky130_fd_pr__nfet_01v8 ad=7.72086e+13p pd=8.6578e+08u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5 a_12002_2130# a_2475_2154# a_11910_2130# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X6 a_5374_4500# col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7 a_14410_15544# col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X8 a_10906_12170# row_n[10] a_11398_12532# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X9 a_35398_9198# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=4.3415e+14p ps=1.9839e+09u w=420000u l=150000u
X10 a_17422_7512# col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X11 a_18026_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=1.47064e+14p ps=1.31646e+09u w=800000u l=150000u
X12 VSS row_n[4] a_9294_6186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X13 a_4370_15544# col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X14 a_23046_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X15 a_22346_10202# rowon_n[8] a_21950_10162# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X16 a_14922_11166# row_n[9] a_15414_11528# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X17 a_15414_2492# col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X18 a_4882_11166# row_n[9] a_5374_11528# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X19 a_34394_2170# col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X20 a_27062_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X21 VSS row_n[6] a_26362_8194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X22 a_1957_14202# VSS sample VDD sky130_fd_pr__pfet_01v8 ad=3.42e+11p pd=2.97e+06u as=6.156e+12p ps=5.346e+07u w=1.2e+06u l=150000u
X23 a_34090_3134# a_2475_3158# a_33998_3134# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X24 a_1957_4162# VDD sample VSS sky130_fd_pr__nfet_01v8 ad=1.71e+11p pd=1.77e+06u as=3.078e+12p ps=3.186e+07u w=600000u l=150000u
X25 a_26058_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X26 a_21342_2170# rowon_n[0] a_20946_2130# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X27 a_35002_9158# row_n[7] a_35494_9520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X28 a_23350_18234# VDD a_22954_18194# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X29 VSS row_n[13] a_20338_15222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X30 a_26970_14178# a_2275_14202# a_27062_14178# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X31 a_11302_8194# rowon_n[6] a_10906_8154# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X32 a_29982_4138# a_2275_4162# a_30074_4138# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X33 a_12306_4178# rowon_n[2] a_11910_4138# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X34 vcm a_2275_2154# a_13006_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X35 VDD rowon_n[3] a_22954_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X36 VSS row_n[12] a_24354_14218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X37 a_21342_11206# col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X38 a_34394_10202# col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X39 a_24962_17190# a_2275_17214# a_25054_17190# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X40 a_18938_7150# a_2275_7174# a_19030_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X41 a_4274_13214# rowon_n[11] a_3878_13174# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X42 a_14314_13214# rowon_n[11] a_13918_13174# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X43 VSS row_n[8] a_11302_10202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X44 a_20034_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X45 a_21038_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X46 a_19430_18556# col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X47 a_19030_14178# a_2475_14202# a_18938_14178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X48 a_11910_11166# a_2275_11190# a_12002_11166# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X49 VDD VSS VSS sky130_fd_pr__cap_var_lvt w=1.64e+07u l=1.6e+07u
X50 VDD rowon_n[14] a_22954_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X51 a_28978_14178# row_n[12] a_29470_14540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X52 a_20434_13536# col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X53 a_33486_12532# col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X54 vcm a_2275_10186# a_29070_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X55 a_20338_6186# col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X56 a_15926_12170# a_2275_12194# a_16018_12170# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X57 a_3270_7190# rowon_n[5] a_2874_7150# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X58 VSS row_n[4] a_30378_6186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X59 a_4274_3174# rowon_n[1] a_3878_3134# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X60 VDD rowon_n[2] a_11910_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X61 a_5886_12170# a_2275_12194# a_5978_12170# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X62 VDD rowon_n[10] a_9902_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X63 a_16322_6186# rowon_n[4] a_15926_6146# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X64 vcm a_2275_6170# a_24050_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X65 a_35398_18234# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X66 VDD rowon_n[9] a_3878_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X67 VDD rowon_n[9] a_13918_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X68 VDD rowon_n[4] a_5886_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X69 VSS VDD a_12306_18234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X70 a_30074_17190# a_2475_17214# a_29982_17190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X71 a_16018_7150# a_2475_7174# a_15926_7150# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X72 a_26058_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X73 a_25054_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X74 a_13310_14218# col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X75 VDD en_C0_n a_3878_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X76 a_30986_17190# row_n[15] a_31478_17552# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X77 a_12002_16186# a_2475_16210# a_11910_16186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X78 a_34090_16186# a_2475_16210# a_33998_16186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X79 a_3270_14218# col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X80 vcm a_2275_13198# a_31078_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X81 a_25358_4178# col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X82 a_35002_16186# row_n[14] a_35494_16548# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X83 a_10906_8154# row_n[6] a_11398_8516# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X84 VSS row_n[6] a_34394_8194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X85 a_8290_5182# rowon_n[3] a_7894_5142# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X86 a_9294_1166# VSS a_8898_1126# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X87 VSS row_n[2] a_35398_4178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X88 a_9994_9158# a_2475_9182# a_9902_9158# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X89 a_12402_16548# col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X90 a_19334_16226# rowon_n[14] a_18938_16186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X91 a_20338_11206# rowon_n[9] a_19942_11166# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X92 vcm a_2275_8178# a_28066_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X93 vcm a_2275_4162# a_29070_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X94 VSS a_2161_13198# a_2275_13198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.71e+11p ps=1.77e+06u w=600000u l=150000u
X95 a_25358_7190# rowon_n[5] a_24962_7150# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X96 a_25054_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X97 a_13310_7190# col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X98 a_29070_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X99 a_14314_3174# col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X100 a_16018_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X101 a_33998_9158# a_2275_9182# a_34090_9158# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X102 VDD rowon_n[1] a_7894_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X103 a_24962_4138# row_n[2] a_25454_4500# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X104 a_5978_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X105 a_2874_7150# row_n[5] a_3366_7512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X106 vcm a_2275_7174# a_17022_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X107 a_35494_4500# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X108 a_19942_11166# a_2275_11190# a_20034_11166# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X109 a_32994_10162# a_2275_10186# a_33086_10162# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X110 a_15926_6146# row_n[4] a_16418_6508# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X111 a_34394_18234# VDD a_33998_18194# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X112 a_27366_17230# col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X113 VSS row_n[13] a_31382_15222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X114 a_13918_1126# VDD a_14410_1488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X115 VSS row_n[12] a_35398_14218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X116 a_32386_11206# col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X117 a_6282_2170# col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X118 a_22954_18194# a_2275_18218# a_23046_18194# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X119 a_12306_14218# rowon_n[12] a_11910_14178# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X120 a_18330_5182# col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X121 a_19334_1166# en_bit_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X122 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X123 VDD rowon_n[15] a_29982_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X124 a_26058_15182# a_2475_15206# a_25966_15182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X125 VSS en_bit_n[0] a_20338_1166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X126 vcm a_2275_11190# a_27062_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X127 a_7894_5142# row_n[3] a_8386_5504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X128 a_30378_1166# VSS a_29982_1126# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X129 VDD rowon_n[14] a_33998_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X130 a_26970_15182# row_n[13] a_27462_15544# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X131 a_31478_13536# col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X132 a_3878_13174# a_2275_13198# a_3970_13174# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X133 a_13918_13174# a_2275_13198# a_14010_13174# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X134 a_23046_5142# a_2475_5166# a_22954_5142# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X135 VDD rowon_n[6] a_30986_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X136 a_17934_3134# row_n[1] a_18426_3496# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X137 a_29374_9198# col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X138 a_29982_12170# row_n[10] a_30474_12532# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X139 VSS row_n[1] a_24354_3174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X140 a_10394_7512# col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X141 a_33390_7190# rowon_n[5] a_32994_7150# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X142 a_34394_3174# rowon_n[1] a_33998_3134# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X143 a_18330_11206# rowon_n[9] a_17934_11166# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X144 a_10998_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X145 VSS row_n[7] a_14314_9198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X146 a_27062_7150# a_2475_7174# a_26970_7150# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X147 a_28066_3134# a_2475_3158# a_27974_3134# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X148 vcm a_2275_9182# a_32082_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X149 a_18938_18194# VDD a_19430_18556# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X150 vcm a_2275_14202# a_8990_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X151 vcm a_2275_14202# a_19030_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X152 a_4974_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X153 a_28978_9158# row_n[7] a_29470_9520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X154 a_8898_18194# VDD a_9390_18556# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X155 a_22954_8154# a_2275_8178# a_23046_8154# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X156 a_24450_1488# col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X157 a_19030_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X158 VSS row_n[0] a_13310_2170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X159 a_23958_4138# a_2275_4162# a_24050_4138# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X160 a_33086_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X161 a_23046_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X162 VSS VDD a_29374_1166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X163 a_14410_9520# col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X164 a_15414_5504# col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X165 VSS row_n[13] a_29374_15222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X166 a_33390_13214# rowon_n[11] a_32994_13174# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X167 a_26362_12210# col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X168 VSS row_n[8] a_30378_10202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X169 a_16018_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X170 VSS row_n[2] a_7286_4178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X171 a_30986_11166# a_2275_11190# a_31078_11166# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X172 a_11910_7150# a_2275_7174# a_12002_7150# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X173 VDD rowon_n[15] a_27974_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X174 a_25454_14540# col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X175 a_35002_12170# a_2275_12194# a_35094_12170# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X176 a_25054_10162# a_2475_10186# a_24962_10162# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X177 a_27974_6146# a_2275_6170# a_28066_6146# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X178 a_32082_1126# a_2475_1150# a_31990_1126# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X179 a_5886_9158# a_2275_9182# a_5978_9158# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X180 a_33998_18194# a_2275_18218# a_34090_18194# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X181 a_29470_13536# col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X182 VDD rowon_n[9] a_32994_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X183 a_25966_10162# row_n[8] a_26458_10524# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X184 a_32994_7150# row_n[5] a_33486_7512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X185 a_7382_4500# col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X186 a_14010_2130# a_2475_2154# a_13918_2130# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X187 a_30986_2130# row_n[0] a_31478_2492# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X188 VDD rowon_n[0] a_18938_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X189 a_11910_14178# a_2275_14202# a_12002_14178# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X190 VDD rowon_n[10] a_8898_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X191 a_16930_5142# a_2275_5166# a_17022_5142# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X192 a_17422_2492# col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X193 vcm a_2275_15206# a_23046_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X194 VSS row_n[6] a_28370_8194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X195 a_17022_17190# a_2475_17214# a_16930_17190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X196 a_8290_15222# col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X197 a_18330_15222# col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X198 a_6982_17190# a_2475_17214# a_6890_17190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X199 a_9902_17190# a_2275_17214# a_9994_17190# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X200 a_1957_8178# VSS sample VDD sky130_fd_pr__pfet_01v8 ad=3.42e+11p pd=2.97e+06u as=0p ps=0u w=1.2e+06u l=150000u
X201 a_23350_2170# rowon_n[0] a_22954_2130# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X202 vcm a_2275_10186# a_14010_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X203 a_2966_9158# a_2475_9182# a_2874_9158# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X204 a_2161_6170# sample VSS VSS sky130_fd_pr__nfet_01v8 ad=1.71e+11p pd=1.77e+06u as=0p ps=0u w=600000u l=150000u
X205 a_7382_17552# col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X206 a_17422_17552# col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X207 a_3878_14178# row_n[12] a_4370_14540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X208 a_13918_14178# row_n[12] a_14410_14540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X209 a_25358_12210# rowon_n[10] a_24962_12170# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X210 vcm a_2275_10186# a_3970_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X211 a_13310_8194# rowon_n[6] a_12914_8154# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X212 vcm a_2275_8178# a_21038_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X213 vcm a_2275_4162# a_22042_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X214 a_14314_4178# rowon_n[2] a_13918_4138# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X215 a_17934_13174# row_n[11] a_18426_13536# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X216 a_29374_11206# rowon_n[9] a_28978_11166# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X217 a_31078_8154# a_2475_8178# a_30986_8154# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X218 vcm a_2275_2154# a_15014_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X219 a_7894_13174# row_n[11] a_8386_13536# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X220 VDD rowon_n[6] a_2874_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X221 a_23046_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X222 a_22042_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X223 VDD rowon_n[8] a_24962_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X224 VDD rowon_n[2] a_13918_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X225 vcm a_2275_18218# a_4974_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X226 vcm a_2275_18218# a_15014_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X227 VSS row_n[15] a_23350_17230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X228 VSS row_n[4] a_32386_6186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X229 a_6282_3174# rowon_n[1] a_5886_3134# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X230 vcm a_2275_6170# a_26058_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X231 VSS row_n[14] a_27366_16226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X232 a_31382_14218# rowon_n[12] a_30986_14178# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X233 a_24354_13214# col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X234 vcm a_2275_9182# a_3970_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X235 VDD rowon_n[4] a_7894_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X236 a_2475_4162# a_1957_4162# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.71e+11p pd=1.77e+06u as=0p ps=0u w=600000u l=150000u
X237 a_32082_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X238 a_17326_15222# rowon_n[13] a_16930_15182# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X239 a_11302_5182# col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X240 a_12306_1166# col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X241 a_28066_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X242 a_7286_15222# rowon_n[13] a_6890_15182# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X243 a_19942_14178# a_2275_14202# a_20034_14178# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X244 a_32994_13174# a_2275_13198# a_33086_13174# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X245 a_18026_7150# a_2475_7174# a_17934_7150# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X246 a_27062_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X247 VDD VDD a_25966_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X248 a_3970_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X249 a_14010_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X250 a_23446_15544# col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X251 VSS row_n[9] a_8290_11206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X252 VSS row_n[9] a_18330_11206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X253 a_23046_11166# a_2475_11190# a_22954_11166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X254 VDD VSS a_5886_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X255 a_23958_11166# row_n[9] a_24450_11528# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X256 a_12914_8154# row_n[6] a_13406_8516# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X257 VDD rowon_n[6] a_24962_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X258 VDD rowon_n[11] a_6890_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X259 VDD rowon_n[11] a_16930_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X260 a_10906_3134# row_n[1] a_11398_3496# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X261 a_12306_17230# col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X262 a_22346_9198# col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X263 a_27366_7190# rowon_n[5] a_26970_7150# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X264 a_16322_3174# col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X265 vcm a_2275_4162# a_30074_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X266 a_16322_16226# col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X267 vcm a_2275_16210# a_21038_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X268 a_15318_7190# col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X269 a_15014_18194# a_2475_18218# a_14922_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X270 a_6282_16226# col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X271 vcm a_2275_15206# a_34090_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X272 a_4882_7150# row_n[5] a_5374_7512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X273 a_4974_18194# a_2475_18218# a_4882_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X274 vcm a_2275_7174# a_19030_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X275 a_17934_6146# row_n[4] a_18426_6508# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X276 a_21038_3134# a_2475_3158# a_20946_3134# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X277 a_15414_18556# col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X278 a_11910_15182# row_n[13] a_12402_15544# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X279 vcm a_2275_11190# a_12002_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X280 a_20034_7150# a_2475_7174# a_19942_7150# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X281 a_2874_2130# row_n[0] a_3366_2492# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X282 a_5374_18556# col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X283 a_21950_9158# row_n[7] a_22442_9520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X284 a_15926_1126# VDD a_16418_1488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X285 a_8290_2170# col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X286 a_28066_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X287 a_9902_2130# a_2275_2154# a_9994_2130# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X288 VSS row_n[10] a_22346_12210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X289 VSS VDD a_22346_1166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X290 a_32386_1166# VSS a_31990_1126# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X291 a_31382_5182# rowon_n[3] a_30986_5142# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X292 a_26058_1126# a_2475_1150# a_25966_1126# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X293 VSS VDD a_21342_18234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X294 a_25054_5142# a_2475_5166# a_24962_5142# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X295 VDD rowon_n[12] a_20946_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X296 a_22346_14218# col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X297 a_16322_10202# rowon_n[8] a_15926_10162# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X298 VDD rowon_n[6] a_32994_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X299 a_26970_7150# row_n[5] a_27462_7512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X300 a_6282_10202# rowon_n[8] a_5886_10162# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X301 a_30074_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X302 a_22442_10524# col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X303 a_20946_6146# a_2275_6170# a_21038_6146# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X304 a_5278_16226# rowon_n[14] a_4882_16186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X305 a_15318_16226# rowon_n[14] a_14922_16186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X306 a_31078_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X307 VDD rowon_n[1] a_30986_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X308 a_20338_17230# col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X309 a_21438_16548# col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X310 a_30986_14178# a_2275_14202# a_31078_14178# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X311 a_18330_9198# rowon_n[7] a_17934_9158# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X312 a_30378_9198# col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X313 a_12402_7512# col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X314 a_13006_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X315 VSS row_n[4] a_4274_6186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X316 a_6890_15182# a_2275_15206# a_6982_15182# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X317 a_16930_15182# a_2275_15206# a_17022_15182# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X318 vcm a_2275_9182# a_34090_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X319 a_29070_7150# a_2475_7174# a_28978_7150# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X320 a_10394_2492# col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X321 VSS row_n[13] a_4274_15222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X322 VSS row_n[13] a_14314_15222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X323 a_11302_12210# col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X324 a_19942_15182# row_n[13] a_20434_15544# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X325 a_15318_11206# col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X326 vcm a_2275_11190# a_20034_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X327 a_6982_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X328 VSS row_n[6] a_21342_8194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X329 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X330 a_32994_14178# row_n[12] a_33486_14540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X331 a_14010_13174# a_2475_13198# a_13918_13174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X332 a_5278_11206# col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X333 vcm a_2275_10186# a_33086_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X334 a_24962_8154# a_2275_8178# a_25054_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X335 VSS row_n[0] a_15318_2170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X336 a_25966_4138# a_2275_4162# a_26058_4138# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X337 a_3970_13174# a_2475_13198# a_3878_13174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X338 VDD rowon_n[7] a_17934_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X339 a_29982_9158# row_n[7] a_30474_9520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X340 a_35094_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X341 VDD rowon_n[3] a_18938_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X342 a_30986_5142# row_n[3] a_31478_5504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X343 VDD rowon_n[15] a_2874_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X344 VDD rowon_n[15] a_12914_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X345 vcm a_2275_16210# a_32082_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X346 a_10394_14540# col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X347 a_5978_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X348 a_14410_13536# col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X349 a_10906_10162# row_n[8] a_11398_10524# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X350 a_17422_5504# col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X351 a_18026_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X352 VSS row_n[2] a_9294_4178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X353 a_4370_13536# col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X354 VDD a_2161_7174# a_2275_7174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.42e+11p ps=2.97e+06u w=1.2e+06u l=150000u
X355 a_13918_7150# a_2275_7174# a_14010_7150# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X356 VSS row_n[4] a_26362_6186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X357 a_1957_2154# VDD sample VSS sky130_fd_pr__nfet_01v8 ad=1.71e+11p pd=1.77e+06u as=0p ps=0u w=600000u l=150000u
X358 a_26058_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X359 a_7894_9158# a_2275_9182# a_7986_9158# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X360 a_35002_7150# row_n[5] a_35494_7512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X361 a_9390_4500# col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X362 VSS VDD a_19334_18234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X363 a_23350_16226# rowon_n[14] a_22954_16186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X364 VSS row_n[11] a_20338_13214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X365 a_11302_6186# rowon_n[4] a_10906_6146# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X366 VSS row_n[10] a_33390_12210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X367 a_32994_2130# row_n[0] a_33486_2492# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X368 a_6890_2130# a_2275_2154# a_6982_2130# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X369 a_10298_12210# rowon_n[10] a_9902_12170# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X370 a_24962_15182# a_2275_15206# a_25054_15182# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X371 a_18938_5142# a_2275_5166# a_19030_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X372 a_28066_12170# a_2475_12194# a_27974_12170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X373 a_4274_11206# rowon_n[9] a_3878_11166# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X374 a_14314_11206# rowon_n[9] a_13918_11166# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X375 a_10998_7150# a_2475_7174# a_10906_7150# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X376 a_21038_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X377 a_20034_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X378 a_8990_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X379 a_19430_16548# col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X380 VDD rowon_n[12] a_31990_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X381 a_28978_12170# row_n[10] a_29470_12532# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X382 a_20434_11528# col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X383 a_33486_10524# col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X384 a_20338_4178# col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X385 a_3270_5182# rowon_n[3] a_2874_5142# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X386 a_4274_1166# en_C0_n a_3878_1126# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X387 VSS row_n[2] a_30378_4178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X388 a_31382_17230# col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X389 VDD rowon_n[8] a_9902_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X390 a_4974_9158# a_2475_9182# a_4882_9158# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X391 a_19030_2130# a_2475_2154# a_18938_2130# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X392 a_16322_4178# rowon_n[2] a_15926_4138# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X393 vcm a_2275_8178# a_23046_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X394 vcm a_2275_4162# a_24050_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X395 a_35398_16226# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X396 a_33086_8154# a_2475_8178# a_32994_8154# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X397 VSS row_n[14] a_12306_16226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X398 a_20338_7190# rowon_n[5] a_19942_7150# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X399 vcm a_2275_17214# a_26058_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X400 a_30074_15182# a_2475_15206# a_29982_15182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X401 a_24050_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X402 a_16018_5142# a_2475_5166# a_15926_5142# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X403 a_25054_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X404 a_34090_14178# a_2475_14202# a_33998_14178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X405 VDD rowon_n[1] a_2874_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X406 a_19942_4138# row_n[2] a_20434_4500# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X407 a_34490_18556# col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X408 a_30986_15182# row_n[13] a_31478_15544# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X409 a_12002_14178# a_2475_14202# a_11910_14178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X410 vcm a_2275_11190# a_31078_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X411 vcm a_2275_7174# a_12002_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X412 a_30474_4500# col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X413 VDD VDD a_10906_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X414 vcm a_2275_12194# a_17022_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X415 a_10906_6146# row_n[4] a_11398_6508# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X416 VSS row_n[4] a_34394_6186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X417 a_8290_3174# rowon_n[1] a_7894_3134# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X418 VDD rowon_n[2] a_15926_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X419 vcm a_2275_12194# a_6982_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X420 a_19334_14218# rowon_n[12] a_18938_14178# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X421 vcm a_2275_6170# a_28066_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X422 vcm a_2275_9182# a_5978_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X423 a_21038_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X424 a_2475_8178# a_1957_8178# VDD VDD sky130_fd_pr__pfet_01v8 ad=3.42e+11p pd=2.97e+06u as=0p ps=0u w=1.2e+06u l=150000u
X425 a_25358_5182# rowon_n[3] a_24962_5142# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X426 a_13310_5182# col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X427 a_14314_1166# col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X428 a_29070_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X429 VDD VSS a_7894_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X430 VDD rowon_n[6] a_26970_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X431 a_2874_5142# row_n[3] a_3366_5504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X432 vcm a_2275_5166# a_17022_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X433 a_30378_17230# rowon_n[15] a_29982_17190# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X434 a_14922_8154# row_n[6] a_15414_8516# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X435 a_3970_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X436 a_14010_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X437 a_34394_16226# rowon_n[14] a_33998_16186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X438 a_27366_15222# col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X439 VSS row_n[11] a_31382_13214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X440 VDD rowon_n[1] a_24962_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X441 a_12914_3134# row_n[1] a_13406_3496# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X442 a_24354_9198# col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X443 VSS row_n[5] a_19334_7190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X444 a_29374_7190# rowon_n[5] a_28978_7150# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X445 a_22954_16186# a_2275_16210# a_23046_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X446 a_18330_3174# col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X447 a_6982_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X448 a_17022_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X449 a_26458_17552# col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X450 VDD rowon_n[13] a_29982_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X451 a_26058_13174# a_2475_13198# a_25966_13174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X452 VDD VSS VSS sky130_fd_pr__cap_var_lvt w=1.64e+07u l=1.6e+07u
X453 a_30378_12210# col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X454 a_26970_13174# row_n[11] a_27462_13536# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X455 a_31478_11528# col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X456 a_22042_7150# a_2475_7174# a_21950_7150# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X457 a_23046_3134# a_2475_3158# a_22954_3134# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X458 VDD rowon_n[4] a_30986_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X459 a_4882_2130# row_n[0] a_5374_2492# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X460 vcm a_2275_12194# a_25054_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X461 a_23958_9158# row_n[7] a_24450_9520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X462 a_17934_1126# en_bit_n[1] a_18426_1488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X463 a_19334_18234# col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X464 vcm a_2275_18218# a_24050_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X465 a_29982_10162# row_n[8] a_30474_10524# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X466 a_9294_18234# col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X467 VSS VDD a_24354_1166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X468 a_9390_14540# col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X469 a_10394_5504# col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X470 a_33390_5182# rowon_n[3] a_32994_5142# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X471 a_28066_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X472 a_10998_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X473 a_28066_1126# a_2475_1150# a_27974_1126# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X474 a_27062_5142# a_2475_5166# a_26970_5142# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X475 a_19030_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X476 a_18938_16186# row_n[14] a_19430_16548# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X477 a_28978_7150# row_n[5] a_29470_7512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X478 a_8898_16186# row_n[14] a_9390_16548# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X479 a_22954_6146# a_2275_6170# a_23046_6146# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X480 a_33086_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X481 a_26970_2130# row_n[0] a_27462_2492# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X482 VDD rowon_n[1] a_32994_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X483 a_28370_17230# rowon_n[15] a_27974_17190# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X484 a_14410_7512# col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X485 VSS row_n[11] a_29374_13214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X486 a_33390_11206# rowon_n[9] a_32994_11166# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X487 a_26362_10202# col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X488 a_15014_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X489 VSS a_2161_1150# a_2275_1150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.71e+11p ps=1.77e+06u w=600000u l=150000u
X490 a_16018_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X491 a_11910_5142# a_2275_5166# a_12002_5142# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X492 a_12402_2492# col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X493 a_9294_12210# rowon_n[10] a_8898_12170# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X494 a_16930_10162# a_2275_10186# a_17022_10162# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X495 a_8990_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X496 VSS row_n[6] a_23350_8194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X497 a_31382_2170# col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X498 a_19334_2170# rowon_n[0] a_18938_2130# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X499 VDD rowon_n[13] a_27974_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X500 a_25454_12532# col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X501 a_6890_10162# a_2275_10186# a_6982_10162# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X502 VSS row_n[0] a_17326_2170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X503 a_27974_4138# a_2275_4162# a_28066_4138# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X504 a_33998_16186# a_2275_16210# a_34090_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X505 a_29470_11528# col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X506 a_32994_5142# row_n[3] a_33486_5504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X507 a_7986_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X508 VDD rowon_n[8] a_8898_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X509 vcm a_2275_2154# a_9994_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X510 VSS row_n[15] a_7286_17230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X511 VSS row_n[15] a_17326_17230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X512 a_22042_17190# a_2475_17214# a_21950_17190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X513 a_15926_7150# a_2275_7174# a_16018_7150# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X514 a_16930_3134# a_2275_3158# a_17022_3134# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X515 a_18330_13214# col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X516 vcm a_2275_13198# a_23046_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X517 VSS row_n[4] a_28370_6186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X518 a_22954_17190# row_n[15] a_23446_17552# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X519 a_17022_15182# a_2475_15206# a_16930_15182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X520 a_8290_13214# col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X521 VSS row_n[7] a_6282_9198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X522 a_6982_15182# a_2475_15206# a_6890_15182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X523 a_9902_15182# a_2275_15206# a_9994_15182# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X524 a_1957_6170# VSS sample VDD sky130_fd_pr__pfet_01v8 ad=3.42e+11p pd=2.97e+06u as=0p ps=0u w=1.2e+06u l=150000u
X525 a_17422_15544# col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X526 a_2161_4162# sample VSS VSS sky130_fd_pr__nfet_01v8 ad=1.71e+11p pd=1.77e+06u as=0p ps=0u w=600000u l=150000u
X527 a_7382_15544# col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X528 a_3878_12170# row_n[10] a_4370_12532# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X529 a_13918_12170# row_n[10] a_14410_12532# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X530 a_26058_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X531 a_25358_10202# rowon_n[8] a_24962_10162# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X532 a_13310_6186# rowon_n[4] a_12914_6146# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X533 vcm a_2275_6170# a_21038_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X534 a_17934_11166# row_n[9] a_18426_11528# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X535 a_31078_6146# a_2475_6170# a_30986_6146# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X536 a_35002_2130# row_n[0] a_35494_2492# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X537 a_8898_2130# a_2275_2154# a_8990_2130# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X538 a_7894_11166# row_n[9] a_8386_11528# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X539 VDD rowon_n[4] a_2874_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X540 a_6378_9520# col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X541 a_23046_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X542 a_13006_7150# a_2475_7174# a_12914_7150# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X543 a_22042_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X544 vcm a_2275_17214# a_10998_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X545 a_24962_10162# a_2275_10186# a_25054_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X546 VDD rowon_n[6] a_19942_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X547 a_26362_18234# VDD a_25966_18194# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X548 vcm a_2275_16210# a_4974_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X549 vcm a_2275_16210# a_15014_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X550 VSS row_n[13] a_23350_15222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X551 a_6982_9158# a_2475_9182# a_6890_9158# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X552 a_6282_1166# VSS a_5886_1126# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X553 VSS row_n[2] a_32386_4178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X554 vcm a_2275_8178# a_25054_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X555 vcm a_2275_4162# a_26058_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X556 VSS row_n[12] a_27366_14218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X557 a_24354_11206# col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X558 a_35094_8154# a_2475_8178# a_35002_8154# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X559 a_27974_17190# a_2275_17214# a_28066_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X560 a_5978_2130# a_2475_2154# a_5886_2130# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X561 a_2475_2154# a_1957_2154# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.71e+11p pd=1.77e+06u as=0p ps=0u w=600000u l=150000u
X562 VDD rowon_n[15] a_21950_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X563 a_32082_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X564 a_17326_13214# rowon_n[11] a_16930_13174# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X565 a_22346_7190# rowon_n[5] a_21950_7150# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X566 a_11302_3174# col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X567 a_7286_13214# rowon_n[11] a_6890_13174# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X568 a_30986_9158# a_2275_9182# a_31078_9158# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X569 a_10298_7190# col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X570 a_18026_5142# a_2475_5166# a_17934_5142# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X571 a_27062_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X572 VDD rowon_n[14] a_25966_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X573 a_3970_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X574 a_14010_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X575 a_23446_13536# col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X576 a_32482_4500# col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X577 a_18938_12170# a_2275_12194# a_19030_12170# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X578 vcm a_2275_7174# a_14010_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X579 a_12914_6146# row_n[4] a_13406_6508# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X580 VDD rowon_n[4] a_24962_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X581 a_8898_12170# a_2275_12194# a_8990_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X582 VDD rowon_n[9] a_6890_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X583 VDD rowon_n[9] a_16930_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X584 a_10906_1126# VDD a_11398_1488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X585 VSS VDD a_15318_18234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X586 a_20034_18194# a_2475_18218# a_19942_18194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X587 a_12306_15222# col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X588 vcm a_2275_9182# a_7986_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X589 a_3270_2170# col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X590 VSS VDD a_5278_18234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X591 a_10998_17190# a_2475_17214# a_10906_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X592 a_33086_17190# a_2475_17214# a_32994_17190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X593 a_16322_1166# col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X594 a_27366_5182# rowon_n[3] a_26970_5142# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X595 a_20946_18194# VDD a_21438_18556# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X596 a_16322_14218# col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X597 vcm a_2275_14202# a_21038_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X598 a_5278_8194# rowon_n[6] a_4882_8154# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X599 a_15318_5182# col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X600 a_33998_17190# row_n[15] a_34490_17552# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X601 a_15014_16186# a_2475_16210# a_14922_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X602 a_6282_14218# col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X603 vcm a_2275_13198# a_34090_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X604 a_19430_8516# col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X605 a_4882_5142# row_n[3] a_5374_5504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X606 vcm a_2275_2154# a_6982_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X607 a_11398_17552# col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X608 a_4974_16186# a_2475_16210# a_4882_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X609 VDD rowon_n[6] a_28978_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X610 vcm a_2275_5166# a_19030_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X611 a_21038_1126# a_2475_1150# a_20946_1126# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X612 a_20034_5142# a_2475_5166# a_19942_5142# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X613 a_15414_16548# col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X614 a_11910_13174# row_n[11] a_12402_13536# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X615 VDD rowon_n[1] a_26970_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X616 a_5374_16548# col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X617 a_21950_7150# row_n[5] a_22442_7512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X618 a_14922_3134# row_n[1] a_15414_3496# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X619 a_2475_16210# a_1957_16210# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.71e+11p pd=1.77e+06u as=0p ps=0u w=600000u l=150000u
X620 a_28066_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X621 vcm a_2275_12194# a_9994_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X622 a_26362_9198# col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X623 VSS row_n[8] a_22346_10202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X624 a_22954_11166# a_2275_11190# a_23046_11166# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X625 a_31382_3174# rowon_n[1] a_30986_3134# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X626 a_25054_3134# a_2475_3158# a_24962_3134# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X627 VSS row_n[14] a_21342_16226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X628 a_24050_7150# a_2475_7174# a_23958_7150# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X629 VDD rowon_n[10] a_20946_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X630 a_25966_9158# row_n[7] a_26458_9520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X631 VDD rowon_n[4] a_32994_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X632 a_26970_5142# row_n[3] a_27462_5504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X633 a_25966_18194# a_2275_18218# a_26058_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X634 a_30074_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X635 a_19942_8154# a_2275_8178# a_20034_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X636 VDD VSS a_30986_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X637 VSS row_n[0] a_10298_2170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X638 a_31078_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X639 a_20946_4138# a_2275_4162# a_21038_4138# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X640 VDD VDD a_19942_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X641 a_5278_14218# rowon_n[12] a_4882_14178# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X642 a_15318_14218# rowon_n[12] a_14922_14178# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X643 a_30074_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X644 a_20338_15222# col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X645 a_2475_17214# a_1957_17214# VDD VDD sky130_fd_pr__pfet_01v8 ad=3.42e+11p pd=2.97e+06u as=0p ps=0u w=1.2e+06u l=150000u
X646 a_12402_5504# col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X647 a_13006_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X648 VSS row_n[2] a_4274_4178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X649 a_13310_17230# rowon_n[15] a_12914_17190# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X650 a_6890_13174# a_2275_13198# a_6982_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X651 a_16930_13174# a_2275_13198# a_17022_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X652 a_7286_7190# col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X653 a_3270_17230# rowon_n[15] a_2874_17190# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X654 a_29070_5142# a_2475_5166# a_28978_5142# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X655 VSS row_n[11] a_4274_13214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X656 VSS row_n[11] a_14314_13214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X657 a_32082_12170# a_2475_12194# a_31990_12170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X658 a_11302_10202# col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X659 a_19942_13174# row_n[11] a_20434_13536# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X660 VSS row_n[4] a_21342_6186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X661 a_32994_12170# row_n[10] a_33486_12532# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X662 a_14010_11166# a_2475_11190# a_13918_11166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X663 a_24962_6146# a_2275_6170# a_25054_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X664 a_31078_18194# a_2475_18218# a_30986_18194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X665 a_3970_11166# a_2475_11190# a_3878_11166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X666 a_2874_9158# a_2275_9182# a_2966_9158# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X667 VDD rowon_n[5] a_17934_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X668 a_29982_7150# row_n[5] a_30474_7512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X669 a_35094_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X670 a_28978_2130# row_n[0] a_29470_2492# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X671 a_31990_18194# VDD a_32482_18556# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X672 VDD rowon_n[13] a_2874_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X673 VDD rowon_n[13] a_12914_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X674 vcm a_2275_14202# a_32082_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X675 a_10394_12532# col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X676 a_4370_4500# col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X677 a_14410_11528# col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X678 a_18026_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X679 a_4370_11528# col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X680 a_17022_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X681 VDD a_2161_5166# a_2275_5166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.42e+11p ps=2.97e+06u w=1.2e+06u l=150000u
X682 vcm a_2275_17214# a_30074_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X683 a_13918_5142# a_2275_5166# a_14010_5142# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X684 a_33390_2170# col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X685 a_14410_2492# col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X686 VSS row_n[6] a_25358_8194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X687 VSS row_n[2] a_26362_4178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X688 a_35398_8194# rowon_n[6] a_35002_8154# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X689 a_26058_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X690 a_35002_5142# row_n[3] a_35494_5504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X691 a_9994_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X692 VSS row_n[14] a_19334_16226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X693 a_23350_14218# rowon_n[12] a_22954_14178# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X694 a_29374_12210# col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X695 VSS row_n[9] a_20338_11206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X696 VSS row_n[8] a_33390_10202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X697 a_11302_4178# rowon_n[2] a_10906_4138# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X698 a_24050_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X699 a_33998_11166# a_2275_11190# a_34090_11166# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X700 a_10298_10202# rowon_n[8] a_9902_10162# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X701 a_26458_4500# col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X702 a_24962_13174# a_2275_13198# a_25054_13174# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X703 a_17934_7150# a_2275_7174# a_18026_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X704 a_18938_3134# a_2275_3158# a_19030_3134# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X705 VDD VDD a_17934_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X706 a_28466_14540# col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X707 VDD rowon_n[10] a_31990_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X708 a_28066_10162# a_2475_10186# a_27974_10162# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X709 a_10998_5142# a_2475_5166# a_10906_5142# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X710 a_20034_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X711 a_8990_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X712 VSS row_n[7] a_8290_9198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X713 a_28978_10162# row_n[8] a_29470_10524# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X714 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X715 a_3270_3174# rowon_n[1] a_2874_3134# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X716 VDD rowon_n[2] a_10906_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X717 VSS VDD a_34394_18234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X718 a_31382_15222# col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X719 a_9902_10162# a_2275_10186# a_9994_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X720 a_2161_8178# sample VDD VDD sky130_fd_pr__pfet_01v8 ad=3.42e+11p pd=2.97e+06u as=0p ps=0u w=1.2e+06u l=150000u
X721 vcm a_2275_6170# a_23046_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X722 a_11302_18234# VDD a_10906_18194# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X723 a_35398_14218# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X724 a_33086_6146# a_2475_6170# a_32994_6146# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X725 a_29070_18194# a_2475_18218# a_28978_18194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X726 VSS row_n[12] a_12306_14218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X727 a_20338_5182# rowon_n[3] a_19942_5142# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X728 a_30474_17552# col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X729 vcm a_2275_15206# a_26058_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X730 a_30074_13174# a_2475_13198# a_29982_13174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X731 a_8386_9520# col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X732 a_15014_7150# a_2475_7174# a_14922_7150# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X733 a_25054_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X734 a_16018_3134# a_2475_3158# a_15926_3134# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X735 a_24050_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X736 a_2874_17190# a_2275_17214# a_2966_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X737 a_9994_17190# a_2475_17214# a_9902_17190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X738 a_12914_17190# a_2275_17214# a_13006_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X739 VDD VSS a_2874_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X740 a_34490_16548# col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X741 a_30986_13174# row_n[11] a_31478_13536# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X742 VDD rowon_n[6] a_21950_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X743 vcm a_2275_5166# a_12002_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X744 VDD rowon_n[14] a_10906_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X745 vcm a_2275_10186# a_17022_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X746 a_9902_8154# row_n[6] a_10394_8516# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X747 a_8290_1166# VSS a_7894_1126# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X748 VSS row_n[2] a_34394_4178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X749 a_6890_14178# row_n[12] a_7382_14540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X750 a_16930_14178# row_n[12] a_17422_14540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X751 vcm a_2275_10186# a_6982_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X752 a_8990_9158# a_2475_9182# a_8898_9158# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X753 VDD rowon_n[1] a_19942_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X754 vcm a_2275_4162# a_28066_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X755 a_24354_7190# rowon_n[5] a_23958_7150# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X756 a_2475_6170# a_1957_6170# VDD VDD sky130_fd_pr__pfet_01v8 ad=3.42e+11p pd=2.97e+06u as=0p ps=0u w=1.2e+06u l=150000u
X757 a_7986_2130# a_2475_2154# a_7894_2130# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X758 a_25358_3174# rowon_n[1] a_24962_3134# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X759 a_29070_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X760 a_13310_3174# col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X761 a_15318_9198# rowon_n[7] a_14922_9158# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X762 a_32994_9158# a_2275_9182# a_33086_9158# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X763 a_32082_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X764 VDD rowon_n[4] a_26970_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X765 vcm a_2275_3158# a_17022_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X766 a_34490_4500# col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X767 vcm a_2275_18218# a_7986_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X768 vcm a_2275_18218# a_18026_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X769 VSS row_n[15] a_26362_17230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X770 a_30378_15222# rowon_n[13] a_29982_15182# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X771 vcm a_2275_7174# a_16018_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X772 a_14922_6146# row_n[4] a_15414_6508# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X773 a_31990_2130# a_2275_2154# a_32082_2130# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X774 a_34394_14218# rowon_n[12] a_33998_14178# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X775 a_27366_13214# col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X776 VSS row_n[9] a_31382_11206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X777 VDD VSS a_24962_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X778 a_22042_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X779 a_12914_1126# VDD a_13406_1488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X780 VSS row_n[3] a_19334_5182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X781 a_13006_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X782 a_35094_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X783 a_5278_2170# col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X784 a_29374_5182# rowon_n[3] a_28978_5142# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X785 a_2966_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X786 a_22954_14178# a_2275_14202# a_23046_14178# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X787 VDD rowon_n[7] a_14922_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X788 a_7286_8194# rowon_n[6] a_6890_8154# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X789 a_18330_1166# en_bit_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X790 VDD VDD a_28978_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X791 a_6982_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X792 a_17022_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X793 a_26458_15544# col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X794 VDD rowon_n[11] a_29982_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X795 a_26058_11166# a_2475_11190# a_25966_11166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X796 vcm a_2275_2154# a_8990_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X797 a_30378_10202# col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X798 VDD a_2161_12194# a_2275_12194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.42e+11p ps=2.97e+06u w=1.2e+06u l=150000u
X799 a_26970_11166# row_n[9] a_27462_11528# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X800 a_23046_1126# a_2475_1150# a_22954_1126# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X801 a_19430_3496# col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X802 a_22042_5142# a_2475_5166# a_21950_5142# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X803 VDD rowon_n[1] a_28978_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X804 a_24962_14178# row_n[12] a_25454_14540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X805 vcm a_2275_10186# a_25054_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X806 a_23958_7150# row_n[5] a_24450_7512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X807 a_8990_12170# a_2475_12194# a_8898_12170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X808 a_28370_9198# col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X809 a_19334_16226# col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X810 vcm a_2275_16210# a_24050_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X811 a_21950_2130# row_n[0] a_22442_2492# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X812 a_10906_18194# a_2275_18218# a_10998_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X813 a_18026_18194# a_2475_18218# a_17934_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X814 a_9294_16226# col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X815 a_7986_18194# a_2475_18218# a_7894_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X816 a_9390_12532# col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X817 a_2475_11190# a_1957_11190# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.71e+11p pd=1.77e+06u as=0p ps=0u w=600000u l=150000u
X818 a_27366_2170# col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X819 a_33390_3174# rowon_n[1] a_32994_3134# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X820 a_10998_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X821 a_18426_18556# col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X822 a_27062_3134# a_2475_3158# a_26970_3134# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X823 a_8386_18556# col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X824 vcm a_2275_9182# a_31078_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X825 a_17326_8194# col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X826 a_3970_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X827 a_27974_9158# row_n[7] a_28466_9520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X828 a_28978_5142# row_n[3] a_29470_5504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X829 a_6890_8154# row_n[6] a_7382_8516# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X830 VSS row_n[0] a_12306_2170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X831 a_22954_4138# a_2275_4162# a_23046_4138# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X832 a_32082_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X833 VDD VSS a_32994_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X834 a_33086_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X835 a_2161_17214# sample VSS VSS sky130_fd_pr__nfet_01v8 ad=1.71e+11p pd=1.77e+06u as=0p ps=0u w=600000u l=150000u
X836 a_28370_15222# rowon_n[13] a_27974_15182# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X837 VSS row_n[10] a_25358_12210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X838 a_30074_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X839 a_14410_5504# col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X840 a_2966_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X841 VSS row_n[9] a_29374_11206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X842 a_15014_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X843 a_16018_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X844 a_9294_7190# col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X845 VDD rowon_n[12] a_23958_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X846 a_12002_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X847 a_34090_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X848 a_10906_7150# a_2275_7174# a_10998_7150# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X849 a_11910_3134# a_2275_3158# a_12002_3134# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X850 a_9294_10202# rowon_n[8] a_8898_10162# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X851 VSS row_n[4] a_23350_6186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X852 a_33086_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X853 VDD rowon_n[11] a_27974_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X854 a_25454_10524# col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X855 a_10998_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X856 a_23350_17230# col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X857 a_33998_14178# a_2275_14202# a_34090_14178# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X858 a_4882_9158# a_2275_9182# a_4974_9158# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X859 VDD rowon_n[0] a_17934_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X860 a_2161_18218# sample VDD VDD sky130_fd_pr__pfet_01v8 ad=3.42e+11p pd=2.97e+06u as=0p ps=0u w=1.2e+06u l=150000u
X861 a_29982_2130# row_n[0] a_30474_2492# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X862 a_3878_2130# a_2275_2154# a_3970_2130# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X863 VSS row_n[13] a_7286_15222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X864 VSS row_n[13] a_17326_15222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X865 a_22042_15182# a_2475_15206# a_21950_15182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X866 a_4274_12210# col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X867 a_14314_12210# col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X868 a_15926_5142# a_2275_5166# a_16018_5142# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X869 a_16930_1126# a_2275_1150# a_17022_1126# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X870 a_18330_11206# col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X871 vcm a_2275_11190# a_23046_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X872 a_35398_2170# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X873 VSS row_n[2] a_28370_4178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X874 a_22954_15182# row_n[13] a_23446_15544# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X875 a_17022_13174# a_2475_13198# a_16930_13174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X876 a_8290_11206# col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X877 VSS row_n[6] a_27366_8194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X878 a_6982_13174# a_2475_13198# a_6890_13174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X879 a_9902_13174# a_2275_13198# a_9994_13174# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X880 a_1957_4162# VSS sample VDD sky130_fd_pr__pfet_01v8 ad=3.42e+11p pd=2.97e+06u as=0p ps=0u w=1.2e+06u l=150000u
X881 VDD rowon_n[15] a_5886_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X882 VDD rowon_n[15] a_15926_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X883 a_3366_14540# col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X884 a_13406_14540# col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X885 a_17422_13536# col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X886 a_13918_10162# row_n[8] a_14410_10524# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X887 a_2161_2154# sample VSS VSS sky130_fd_pr__nfet_01v8 ad=1.71e+11p pd=1.77e+06u as=0p ps=0u w=600000u l=150000u
X888 a_7382_13536# col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X889 a_3878_10162# row_n[8] a_4370_10524# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X890 vcm a_2275_8178# a_20034_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X891 vcm a_2275_4162# a_21038_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X892 a_13310_4178# rowon_n[2] a_12914_4138# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X893 a_26970_9158# a_2275_9182# a_27062_9158# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X894 a_30074_8154# a_2475_8178# a_29982_8154# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X895 VSS row_n[5] a_16322_7190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X896 a_31078_4138# a_2475_4162# a_30986_4138# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X897 a_28466_4500# col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X898 a_6378_7512# col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X899 a_13006_5142# a_2475_5166# a_12914_5142# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X900 a_22042_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X901 a_22346_17230# rowon_n[15] a_21950_17190# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X902 vcm a_2275_15206# a_10998_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X903 VDD rowon_n[4] a_19942_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X904 a_4882_18194# VDD a_5374_18556# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X905 a_14922_18194# VDD a_15414_18556# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X906 a_26362_16226# rowon_n[14] a_25966_16186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X907 vcm a_2275_14202# a_4974_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X908 vcm a_2275_14202# a_15014_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X909 VSS row_n[11] a_23350_13214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X910 a_8990_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X911 VDD rowon_n[2] a_12914_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X912 vcm a_2275_6170# a_25054_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X913 a_35094_6146# a_2475_6170# a_35002_6146# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X914 a_27974_15182# a_2275_15206# a_28066_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X915 a_32082_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X916 vcm a_2275_9182# a_2966_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X917 VDD rowon_n[13] a_21950_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X918 a_17326_11206# rowon_n[9] a_16930_11166# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X919 a_11302_1166# col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X920 a_22346_5182# rowon_n[3] a_21950_5142# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X921 VDD rowon_n[12] a_35002_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X922 a_7286_11206# rowon_n[9] a_6890_11166# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X923 a_17022_7150# a_2475_7174# a_16930_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X924 a_10298_5182# col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X925 a_27062_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X926 a_18026_3134# a_2475_3158# a_17934_3134# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X927 a_23446_11528# col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X928 VDD VSS VSS sky130_fd_pr__cap_var_lvt w=1.64e+07u l=1.6e+07u
X929 a_21342_18234# col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X930 VDD rowon_n[6] a_23958_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X931 vcm a_2275_5166# a_14010_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X932 a_34394_17230# col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X933 VDD rowon_n[1] a_21950_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X934 VSS row_n[15] a_11302_17230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X935 a_9902_3134# row_n[1] a_10394_3496# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X936 a_29982_18194# a_2275_18218# a_30074_18194# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X937 VSS row_n[14] a_15318_16226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X938 a_20034_16186# a_2475_16210# a_19942_16186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X939 a_12306_13214# col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X940 vcm a_2275_17214# a_29070_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X941 VSS row_n[14] a_5278_16226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X942 a_10998_15182# a_2475_15206# a_10906_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X943 a_33086_15182# a_2475_15206# a_32994_15182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X944 a_21342_9198# col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X945 VSS row_n[7] a_31382_9198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X946 a_26362_7190# rowon_n[5] a_25966_7150# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X947 a_9994_2130# a_2475_2154# a_9902_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X948 a_27366_3174# rowon_n[1] a_26970_3134# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X949 a_15318_3174# col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X950 a_20946_16186# row_n[14] a_21438_16548# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X951 a_5278_6186# rowon_n[4] a_4882_6146# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X952 a_33998_15182# row_n[13] a_34490_15544# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X953 a_15014_14178# a_2475_14202# a_14922_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X954 vcm a_2275_11190# a_34090_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X955 a_17326_9198# rowon_n[7] a_16930_9158# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X956 a_35002_9158# a_2275_9182# a_35094_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X957 a_19430_6508# col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X958 VDD VDD a_13918_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X959 a_11398_15544# col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X960 a_4974_14178# a_2475_14202# a_4882_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X961 vcm a_2275_7174# a_18026_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X962 VDD rowon_n[4] a_28978_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X963 vcm a_2275_3158# a_19030_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X964 VDD VDD a_3878_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X965 a_20034_3134# a_2475_3158# a_19942_3134# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X966 a_11910_11166# row_n[9] a_12402_11528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X967 a_33998_2130# a_2275_2154# a_34090_2130# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X968 VDD VSS a_26970_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X969 a_20946_9158# row_n[7] a_21438_9520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X970 a_26058_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X971 a_14922_1126# VDD a_15414_1488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X972 a_21950_5142# row_n[3] a_22442_5504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X973 a_31478_9520# col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X974 a_2475_14202# a_1957_14202# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.71e+11p pd=1.77e+06u as=0p ps=0u w=600000u l=150000u
X975 a_9902_14178# row_n[12] a_10394_14540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X976 vcm a_2275_10186# a_9994_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X977 a_21342_12210# rowon_n[10] a_20946_12170# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X978 VDD rowon_n[7] a_16930_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X979 a_9294_8194# rowon_n[6] a_8898_8154# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X980 a_20338_18234# VDD a_19942_18194# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X981 a_31382_1166# VSS a_30986_1126# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X982 a_17022_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X983 a_25054_1126# a_2475_1150# a_24962_1126# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X984 VSS row_n[12] a_21342_14218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X985 a_6982_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X986 a_24050_5142# a_2475_5166# a_23958_5142# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X987 a_21950_17190# a_2275_17214# a_22042_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X988 VDD rowon_n[8] a_20946_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X989 a_25966_7150# row_n[5] a_26458_7512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X990 VDD VSS VSS sky130_fd_pr__cap_var_lvt w=1.64e+07u l=1.6e+07u
X991 a_25966_16186# a_2275_16210# a_26058_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X992 a_30074_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X993 a_19942_6146# a_2275_6170# a_20034_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X994 a_9994_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X995 VDD rowon_n[14] a_19942_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X996 a_30074_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X997 a_23958_2130# row_n[0] a_24450_2492# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X998 a_20338_13214# col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X999 a_33390_12210# col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1000 a_2475_15206# a_1957_15206# VDD VDD sky130_fd_pr__pfet_01v8 ad=3.42e+11p pd=2.97e+06u as=0p ps=0u w=1.2e+06u l=150000u
X1001 a_12002_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1002 a_29374_2170# col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1003 a_13006_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1004 a_3270_15222# rowon_n[13] a_2874_15182# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1005 a_13310_15222# rowon_n[13] a_12914_15182# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1006 VSS row_n[10] a_10298_12210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1007 a_7286_5182# col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1008 a_32386_18234# col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1009 a_19334_8194# col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1010 a_29070_3134# a_2475_3158# a_28978_3134# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1011 a_32482_14540# col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1012 vcm a_2275_12194# a_28066_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1013 VSS row_n[9] a_4274_11206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1014 VSS row_n[9] a_14314_11206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1015 a_32082_10162# a_2475_10186# a_31990_10162# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1016 vcm a_2275_9182# a_33086_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1017 a_19942_11166# row_n[9] a_20434_11528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1018 a_8898_8154# row_n[6] a_9390_8516# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1019 VSS row_n[6] a_20338_8194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1020 VSS row_n[2] a_21342_4178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1021 vcm a_2275_18218# a_27062_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1022 a_31078_16186# a_2475_16210# a_30986_16186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1023 a_32994_10162# row_n[8] a_33486_10524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1024 a_30378_8194# rowon_n[6] a_29982_8154# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1025 VSS row_n[0] a_14314_2170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1026 a_24962_4138# a_2275_4162# a_25054_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1027 a_34090_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1028 VDD rowon_n[3] a_17934_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1029 vcm a_2275_2154# a_32082_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1030 a_35094_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1031 a_29982_5142# row_n[3] a_30474_5504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1032 a_31990_16186# row_n[14] a_32482_16548# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1033 VDD rowon_n[11] a_2874_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1034 VDD rowon_n[11] a_12914_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1035 a_10394_10524# col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1036 a_4974_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1037 a_6890_3134# row_n[1] a_7382_3496# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1038 a_17022_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1039 a_18026_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1040 a_2161_12194# sample VSS VSS sky130_fd_pr__nfet_01v8 ad=1.71e+11p pd=1.77e+06u as=0p ps=0u w=600000u l=150000u
X1041 VDD a_2161_3158# a_2275_3158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.42e+11p ps=2.97e+06u w=1.2e+06u l=150000u
X1042 a_13918_3134# a_2275_3158# a_14010_3134# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1043 a_21438_4500# col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1044 vcm a_2275_15206# a_30074_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1045 a_12914_7150# a_2275_7174# a_13006_7150# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1046 VSS row_n[4] a_25358_6186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1047 VSS row_n[7] a_3270_9198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1048 a_35398_6186# rowon_n[4] a_35002_6146# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1049 a_18330_18234# VDD a_17934_18194# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1050 a_32386_12210# rowon_n[10] a_31990_12170# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1051 VSS row_n[12] a_19334_14218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1052 a_29374_10202# col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1053 ctop sw ctop VDD sky130_fd_pr__pfet_01v8 ad=2.7075e+12p pd=2.185e+07u as=0p ps=0u w=1.9e+06u l=220000u
X1054 a_24050_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1055 a_20946_12170# a_2275_12194# a_21038_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1056 a_5886_2130# a_2275_2154# a_5978_2130# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1057 a_18938_1126# a_2275_1150# a_19030_1126# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1058 a_17934_5142# a_2275_5166# a_18026_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1059 VDD rowon_n[14] a_17934_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1060 a_28466_12532# col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1061 VDD rowon_n[8] a_31990_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1062 a_3366_9520# col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1063 VSS row_n[6] a_29374_8194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1064 a_20034_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1065 a_10998_3134# a_2475_3158# a_10906_3134# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1066 a_8990_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1067 a_16418_8516# col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1068 VSS row_n[15] a_30378_17230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1069 a_3270_1166# VSS a_2874_1126# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1070 VSS row_n[14] a_34394_16226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1071 a_31382_13214# col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1072 a_3970_9158# a_2475_9182# a_3878_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1073 a_32386_7190# col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1074 a_2161_6170# sample VDD VDD sky130_fd_pr__pfet_01v8 ad=3.42e+11p pd=2.97e+06u as=0p ps=0u w=1.2e+06u l=150000u
X1075 a_11302_16226# rowon_n[14] a_10906_16186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1076 vcm a_2275_4162# a_23046_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1077 a_25054_17190# a_2475_17214# a_24962_17190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1078 a_28978_9158# a_2275_9182# a_29070_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1079 a_32082_8154# a_2475_8178# a_31990_8154# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1080 VSS row_n[5] a_18330_7190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1081 a_33086_4138# a_2475_4162# a_32994_4138# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1082 a_29070_16186# a_2475_16210# a_28978_16186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1083 vcm a_2275_13198# a_26058_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1084 a_2966_2130# a_2475_2154# a_2874_2130# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1085 a_20338_3174# rowon_n[1] a_19942_3134# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1086 VDD VDD a_32994_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1087 a_25966_17190# row_n[15] a_26458_17552# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1088 a_30474_15544# col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1089 a_30074_11166# a_2475_11190# a_29982_11166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1090 a_8386_7512# col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1091 a_15014_5142# a_2475_5166# a_14922_5142# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1092 a_16018_1126# a_2475_1150# a_15926_1126# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1093 a_24050_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1094 a_2874_15182# a_2275_15206# a_2966_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1095 a_9994_15182# a_2475_15206# a_9902_15182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1096 a_12914_15182# a_2275_15206# a_13006_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1097 a_10298_9198# rowon_n[7] a_9902_9158# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1098 a_30986_11166# row_n[9] a_31478_11528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1099 VDD rowon_n[4] a_21950_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1100 a_6378_2492# col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1101 vcm a_2275_3158# a_12002_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1102 vcm a_2275_7174# a_10998_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1103 a_9902_6146# row_n[4] a_10394_6508# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1104 a_6890_12170# row_n[10] a_7382_12532# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1105 a_16930_12170# row_n[10] a_17422_12532# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1106 VDD en_bit_n[0] a_19942_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1107 vcm a_2275_9182# a_4974_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1108 a_25358_1166# VSS a_24962_1126# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1109 a_2475_4162# a_1957_4162# VDD VDD sky130_fd_pr__pfet_01v8 ad=3.42e+11p pd=2.97e+06u as=0p ps=0u w=1.2e+06u l=150000u
X1110 a_24354_5182# rowon_n[3] a_23958_5142# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1111 VDD rowon_n[7] a_9902_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1112 a_13310_1166# col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1113 a_29070_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1114 vcm a_2275_17214# a_14010_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1115 a_27974_10162# a_2275_10186# a_28066_10162# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1116 vcm a_2275_2154# a_3970_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1117 vcm a_2275_17214# a_3970_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1118 VDD rowon_n[6] a_25966_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1119 vcm a_2275_1150# a_17022_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1120 a_29374_18234# VDD a_28978_18194# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1121 vcm a_2275_16210# a_7986_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1122 vcm a_2275_16210# a_18026_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1123 VSS row_n[13] a_26362_15222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1124 a_30378_13214# rowon_n[11] a_29982_13174# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1125 vcm a_2275_5166# a_16018_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1126 a_27366_11206# col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1127 VDD rowon_n[1] a_23958_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1128 a_22042_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1129 VSS row_n[1] a_19334_3174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1130 VDD rowon_n[15] a_24962_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1131 a_13006_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1132 a_35094_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1133 a_31990_12170# a_2275_12194# a_32082_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1134 a_23350_9198# col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1135 a_28370_7190# rowon_n[5] a_27974_7150# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1136 a_29374_3174# rowon_n[1] a_28978_3134# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1137 a_2966_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1138 VSS row_n[7] a_33390_9198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1139 VDD rowon_n[5] a_14922_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1140 a_7286_6186# rowon_n[4] a_6890_6146# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1141 VDD rowon_n[14] a_28978_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1142 a_6982_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1143 a_17022_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1144 a_26458_13536# col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1145 VDD rowon_n[9] a_29982_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1146 vcm a_2275_9182# a_27062_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1147 a_22346_2170# col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1148 VDD a_2161_10186# a_2275_10186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.42e+11p ps=2.97e+06u w=1.2e+06u l=150000u
X1149 a_24050_12170# a_2475_12194# a_23958_12170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1150 a_19430_1488# en_bit_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1151 a_22042_3134# a_2475_3158# a_21950_3134# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1152 VSS row_n[10] a_9294_12210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1153 a_12306_8194# col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1154 a_28066_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1155 VDD VSS a_28978_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1156 VSS VDD a_18330_18234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1157 a_23046_18194# a_2475_18218# a_22954_18194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1158 a_24962_12170# row_n[10] a_25454_12532# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1159 a_22954_9158# row_n[7] a_23446_9520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1160 a_23958_5142# row_n[3] a_24450_5504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1161 VSS VDD a_8290_18234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1162 a_8990_10162# a_2475_10186# a_8898_10162# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1163 a_33486_9520# col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1164 a_23958_18194# VDD a_24450_18556# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1165 a_19334_14218# col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1166 vcm a_2275_14202# a_24050_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1167 a_10906_16186# a_2275_16210# a_10998_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1168 a_18026_16186# a_2475_16210# a_17934_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1169 VDD rowon_n[12] a_7894_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1170 a_9294_14218# col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1171 a_7986_16186# a_2475_16210# a_7894_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1172 a_9390_10524# col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1173 a_33390_1166# VSS a_32994_1126# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1174 a_10998_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1175 a_18426_16548# col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1176 a_4274_7190# col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1177 a_27062_1126# a_2475_1150# a_26970_1126# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1178 a_8386_16548# col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1179 a_17326_6186# col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1180 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X1181 a_27974_7150# row_n[5] a_28466_7512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1182 vcm a_2275_12194# a_13006_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1183 a_6890_6146# row_n[4] a_7382_6508# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1184 vcm a_2275_12194# a_2966_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1185 a_32082_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1186 a_25966_2130# row_n[0] a_26458_2492# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1187 a_2161_15206# sample VSS VSS sky130_fd_pr__nfet_01v8 ad=1.71e+11p pd=1.77e+06u as=0p ps=0u w=600000u l=150000u
X1188 a_28370_13214# rowon_n[11] a_27974_13174# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1189 VSS row_n[8] a_25358_10202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1190 vcm a_2275_18218# a_12002_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1191 a_25966_11166# a_2275_11190# a_26058_11166# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1192 a_14010_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1193 a_15014_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1194 a_9294_5182# col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1195 VDD rowon_n[10] a_23958_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1196 vcm a_2275_9182# a_35094_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1197 a_10906_5142# a_2275_5166# a_10998_5142# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1198 a_11910_1126# a_2275_1150# a_12002_1126# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1199 a_30378_2170# col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1200 a_18330_2170# rowon_n[0] a_17934_2130# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1201 VSS row_n[2] a_23350_4178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1202 a_28978_18194# a_2275_18218# a_29070_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1203 a_33086_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1204 VDD rowon_n[9] a_27974_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1205 VSS row_n[6] a_22346_8194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1206 a_32386_8194# rowon_n[6] a_31990_8154# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1207 a_10998_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1208 vcm a_2275_2154# a_34090_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1209 a_23350_15222# col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1210 a_26058_8154# a_2475_8178# a_25966_8154# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1211 a_8898_3134# row_n[1] a_9390_3496# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1212 a_6982_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1213 a_16322_17230# rowon_n[15] a_15926_17190# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1214 a_6282_17230# rowon_n[15] a_5886_17190# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1215 a_2161_16210# sample VDD VDD sky130_fd_pr__pfet_01v8 ad=3.42e+11p pd=2.97e+06u as=0p ps=0u w=1.2e+06u l=150000u
X1216 a_21950_9158# a_2275_9182# a_22042_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1217 VSS row_n[5] a_11302_7190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1218 a_22442_17552# col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1219 VSS row_n[11] a_7286_13214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1220 VSS row_n[11] a_17326_13214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1221 a_22042_13174# a_2475_13198# a_21950_13174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1222 a_35094_12170# a_2475_12194# a_35002_12170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1223 a_4274_10202# col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1224 a_14314_10202# col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1225 a_14922_7150# a_2275_7174# a_15014_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1226 a_15926_3134# a_2275_3158# a_16018_3134# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1227 a_23446_4500# col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1228 a_2966_12170# a_2475_12194# a_2874_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1229 a_13006_12170# a_2475_12194# a_12914_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1230 a_22954_13174# row_n[11] a_23446_13536# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1231 a_17022_11166# a_2475_11190# a_16930_11166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1232 VSS row_n[4] a_27366_6186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1233 a_6982_11166# a_2475_11190# a_6890_11166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1234 VSS row_n[7] a_5278_9198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1235 a_1957_18218# VDD sample VSS sky130_fd_pr__nfet_01v8 ad=1.71e+11p pd=1.77e+06u as=0p ps=0u w=600000u l=150000u
X1236 VDD rowon_n[13] a_5886_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1237 VDD rowon_n[13] a_15926_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1238 a_3366_12532# col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1239 a_13406_12532# col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1240 a_17422_11528# col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1241 a_7382_11528# col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1242 vcm a_2275_6170# a_20034_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1243 a_15318_18234# col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1244 vcm a_2275_18218# a_20034_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1245 a_30074_6146# a_2475_6170# a_29982_6146# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1246 VSS row_n[3] a_16322_5182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1247 a_7894_2130# a_2275_2154# a_7986_2130# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1248 a_5278_18234# col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1249 vcm a_2275_17214# a_33086_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1250 a_5374_9520# col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1251 a_31990_8154# row_n[6] a_32482_8516# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1252 a_6378_5504# col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1253 a_24050_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1254 a_18426_8516# col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1255 a_12002_7150# a_2475_7174# a_11910_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1256 a_22042_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1257 a_13006_3134# a_2475_3158# a_12914_3134# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1258 a_10906_17190# row_n[15] a_11398_17552# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1259 a_22346_15222# rowon_n[13] a_21950_15182# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1260 vcm a_2275_13198# a_10998_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1261 a_4882_16186# row_n[14] a_5374_16548# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1262 a_14922_16186# row_n[14] a_15414_16548# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1263 a_26362_14218# rowon_n[12] a_25966_14178# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1264 VSS row_n[9] a_23350_11206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1265 a_16418_3496# col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1266 a_34394_7190# col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1267 vcm a_2275_4162# a_25054_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1268 a_27062_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1269 a_34090_8154# a_2475_8178# a_33998_8154# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1270 a_35094_4138# a_2475_4162# a_35002_4138# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1271 a_27974_13174# a_2275_13198# a_28066_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1272 a_1957_9182# VDD sample VSS sky130_fd_pr__nfet_01v8 ad=1.71e+11p pd=1.77e+06u as=0p ps=0u w=600000u l=150000u
X1273 VDD rowon_n[11] a_21950_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1274 a_21342_7190# rowon_n[5] a_20946_7150# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1275 a_4974_2130# a_2475_2154# a_4882_2130# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1276 a_22346_3174# rowon_n[1] a_21950_3134# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1277 a_10298_3174# col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1278 VDD rowon_n[10] a_35002_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1279 a_17022_5142# a_2475_5166# a_16930_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1280 a_18026_1126# a_2475_1150# a_17934_1126# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1281 a_12306_9198# rowon_n[7] a_11910_9158# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1282 a_29982_9158# a_2275_9182# a_30074_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1283 a_21342_16226# col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1284 vcm a_2275_7174# a_13006_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1285 VDD rowon_n[4] a_23958_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1286 a_8386_2492# col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1287 vcm a_2275_3158# a_14010_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1288 a_34394_15222# col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1289 a_12914_10162# a_2275_10186# a_13006_10162# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1290 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X1291 a_2874_10162# a_2275_10186# a_2966_10162# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1292 VDD VSS a_21950_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1293 a_4274_18234# VDD a_3878_18194# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1294 a_14314_18234# VDD a_13918_18194# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1295 VSS row_n[13] a_11302_15222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1296 a_21038_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1297 a_9902_1126# VDD a_10394_1488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1298 a_20434_18556# col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1299 a_29982_16186# a_2275_16210# a_30074_16186# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1300 VSS row_n[12] a_15318_14218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1301 a_20034_14178# a_2475_14202# a_19942_14178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1302 a_12306_11206# col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1303 a_33486_17552# col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1304 vcm a_2275_15206# a_29070_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1305 VSS row_n[12] a_5278_14218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1306 a_10998_13174# a_2475_13198# a_10906_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1307 a_33086_13174# a_2475_13198# a_32994_13174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1308 a_15318_1166# col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1309 a_27366_1166# VSS a_26970_1126# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1310 a_26362_5182# rowon_n[3] a_25966_5142# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1311 a_5886_17190# a_2275_17214# a_5978_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1312 a_15926_17190# a_2275_17214# a_16018_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1313 VDD rowon_n[7] a_11910_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1314 a_4274_8194# rowon_n[6] a_3878_8154# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1315 a_5278_4178# rowon_n[2] a_4882_4138# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1316 VDD rowon_n[15] a_9902_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1317 a_33998_13174# row_n[11] a_34490_13536# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1318 vcm a_2275_2154# a_5978_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1319 VDD rowon_n[14] a_13918_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1320 a_11398_13536# col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1321 VDD rowon_n[6] a_27974_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1322 vcm a_2275_5166# a_18026_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1323 vcm a_2275_1150# a_19030_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1324 VDD rowon_n[14] a_3878_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1325 a_20034_1126# a_2475_1150# a_19942_1126# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1326 a_20946_7150# row_n[5] a_21438_7512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1327 a_26058_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1328 VDD rowon_n[1] a_25966_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1329 vcm a_2275_18218# a_31078_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1330 a_31478_7512# col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1331 VDD rowon_n[2] a_4882_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1332 a_9902_12170# row_n[10] a_10394_12532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1333 a_21342_10202# rowon_n[8] a_20946_10162# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1334 a_25358_9198# col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1335 a_22042_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1336 VSS row_n[7] a_35398_9198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1337 VDD rowon_n[5] a_16930_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1338 a_9294_6186# rowon_n[4] a_8898_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1339 a_13006_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1340 a_35094_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1341 vcm a_2275_9182# a_29070_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1342 a_20338_16226# rowon_n[14] a_19942_16186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1343 a_2966_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1344 a_24354_2170# col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1345 VDD rowon_n[0] a_14922_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1346 a_14314_8194# col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1347 a_24050_3134# a_2475_3158# a_23958_3134# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1348 a_25054_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1349 a_21950_15182# a_2275_15206# a_22042_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1350 a_24962_9158# row_n[7] a_25454_9520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1351 a_25966_5142# row_n[3] a_26458_5504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1352 a_16018_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1353 a_35494_9520# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1354 a_3878_8154# row_n[6] a_4370_8516# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1355 a_5978_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1356 a_25966_14178# a_2275_14202# a_26058_14178# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1357 a_19942_4138# a_2275_4162# a_20034_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1358 a_9994_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1359 a_30074_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1360 a_20338_11206# col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1361 a_33390_10202# col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1362 a_2475_13198# a_1957_13198# VDD VDD sky130_fd_pr__pfet_01v8 ad=3.42e+11p pd=2.97e+06u as=0p ps=0u w=1.2e+06u l=150000u
X1363 a_12002_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1364 a_13006_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1365 a_3270_13214# rowon_n[11] a_2874_13174# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1366 a_13310_13214# rowon_n[11] a_12914_13174# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1367 VSS row_n[8] a_10298_10202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1368 a_6282_7190# col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1369 a_7286_3174# col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1370 a_32386_16226# col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1371 a_10906_11166# a_2275_11190# a_10998_11166# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1372 a_19334_6186# col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1373 a_29070_1126# a_2475_1150# a_28978_1126# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1374 a_27974_14178# row_n[12] a_28466_14540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1375 a_32482_12532# col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1376 vcm a_2275_10186# a_28066_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1377 a_14922_12170# a_2275_12194# a_15014_12170# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1378 a_8898_6146# row_n[4] a_9390_6508# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1379 VSS row_n[4] a_20338_6186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1380 vcm a_2275_16210# a_27062_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1381 a_31078_14178# a_2475_14202# a_30986_14178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1382 a_4882_12170# a_2275_12194# a_4974_12170# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1383 a_30378_6186# rowon_n[4] a_29982_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1384 a_13918_18194# a_2275_18218# a_14010_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1385 a_31478_18556# col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1386 a_34090_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1387 a_27974_2130# row_n[0] a_28466_2492# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1388 a_3878_18194# a_2275_18218# a_3970_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1389 VDD rowon_n[9] a_2874_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1390 VDD rowon_n[9] a_12914_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1391 a_6890_1126# VDD a_7382_1488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1392 a_17022_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1393 a_2161_10186# sample VSS VSS sky130_fd_pr__nfet_01v8 ad=1.71e+11p pd=1.77e+06u as=0p ps=0u w=600000u l=150000u
X1394 VDD a_2161_1150# a_2275_1150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.42e+11p ps=2.97e+06u w=1.2e+06u l=150000u
X1395 a_13918_1126# a_2275_1150# a_14010_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1396 a_29982_17190# row_n[15] a_30474_17552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1397 vcm a_2275_13198# a_30074_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1398 a_12914_5142# a_2275_5166# a_13006_5142# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1399 VSS row_n[6] a_24354_8194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1400 VSS row_n[2] a_25358_4178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1401 a_11398_8516# col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1402 a_34394_8194# rowon_n[6] a_33998_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1403 a_35398_4178# rowon_n[2] a_35002_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1404 a_18330_16226# rowon_n[14] a_17934_16186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1405 VSS row_n[10] a_28370_12210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1406 a_33086_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1407 a_32386_10202# rowon_n[8] a_31990_10162# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1408 a_28066_8154# a_2475_8178# a_27974_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1409 a_8990_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1410 a_10998_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1411 a_24050_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1412 a_19030_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1413 VDD rowon_n[12] a_26970_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1414 a_15014_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1415 a_23958_9158# a_2275_9182# a_24050_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1416 VSS row_n[5] a_13310_7190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1417 a_4974_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1418 a_17934_3134# a_2275_3158# a_18026_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1419 VDD rowon_n[2] a_35002_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1420 a_25454_4500# col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1421 a_28466_10524# col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1422 a_3366_7512# col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1423 VSS row_n[4] a_29374_6186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1424 a_10998_1126# a_2475_1150# a_10906_1126# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1425 VSS row_n[7] a_7286_9198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1426 a_16418_6508# col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1427 a_33390_18234# VDD a_32994_18194# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1428 a_26362_17230# col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1429 VSS row_n[13] a_30378_15222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1430 VSS row_n[12] a_34394_14218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1431 a_31382_11206# col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1432 VSS row_n[0] a_6282_2170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1433 a_2161_4162# sample VDD VDD sky130_fd_pr__pfet_01v8 ad=3.42e+11p pd=2.97e+06u as=0p ps=0u w=1.2e+06u l=150000u
X1434 a_32386_5182# col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1435 a_35002_17190# a_2275_17214# a_35094_17190# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1436 a_11302_14218# rowon_n[12] a_10906_14178# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1437 a_1957_13198# VDD sample VSS sky130_fd_pr__nfet_01v8 ad=1.71e+11p pd=1.77e+06u as=0p ps=0u w=600000u l=150000u
X1438 a_25054_15182# a_2475_15206# a_24962_15182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1439 a_7286_12210# col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1440 a_17326_12210# col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1441 vcm a_2275_12194# a_22042_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1442 a_32082_6146# a_2475_6170# a_31990_6146# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1443 VSS row_n[3] a_18330_5182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1444 a_29070_14178# a_2475_14202# a_28978_14178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1445 vcm a_2275_11190# a_26058_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1446 a_33998_8154# row_n[6] a_34490_8516# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1447 a_20338_1166# en_bit_n[0] a_19942_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1448 a_29470_18556# col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1449 VDD rowon_n[14] a_32994_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1450 a_25966_15182# row_n[13] a_26458_15544# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1451 a_30474_13536# col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1452 a_7382_9520# col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1453 a_8386_5504# col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1454 a_24050_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1455 a_15014_3134# a_2475_3158# a_14922_3134# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1456 a_2874_13174# a_2275_13198# a_2966_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1457 a_9994_13174# a_2475_13198# a_9902_13174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1458 a_12914_13174# a_2275_13198# a_13006_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1459 a_14010_7150# a_2475_7174# a_13918_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1460 VDD rowon_n[15] a_8898_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1461 a_6378_14540# col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1462 a_16418_14540# col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1463 VDD rowon_n[6] a_20946_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1464 vcm a_2275_1150# a_12002_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1465 a_31990_3134# row_n[1] a_32482_3496# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1466 vcm a_2275_5166# a_10998_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1467 a_18426_3496# col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1468 a_6890_10162# row_n[8] a_7382_10524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1469 a_16930_10162# row_n[8] a_17422_10524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1470 a_23350_7190# rowon_n[5] a_22954_7150# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1471 a_6982_2130# a_2475_2154# a_6890_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1472 a_24354_3174# rowon_n[1] a_23958_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1473 VDD rowon_n[5] a_9902_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1474 a_25358_17230# rowon_n[15] a_24962_17190# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1475 vcm a_2275_15206# a_14010_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1476 vcm a_2275_15206# a_3970_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1477 a_14314_9198# rowon_n[7] a_13918_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1478 vcm a_2275_9182# a_22042_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1479 VDD rowon_n[4] a_25966_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1480 a_17934_18194# VDD a_18426_18556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1481 a_29374_16226# rowon_n[14] a_28978_16186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1482 vcm a_2275_14202# a_7986_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1483 vcm a_2275_14202# a_18026_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1484 VSS row_n[11] a_26362_13214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1485 a_30378_11206# rowon_n[9] a_29982_11166# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1486 vcm a_2275_7174# a_15014_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1487 vcm a_2275_3158# a_16018_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1488 a_7894_18194# VDD a_8386_18556# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1489 a_30986_2130# a_2275_2154# a_31078_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1490 a_23046_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1491 VDD VSS a_23958_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1492 a_22042_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1493 VSS en_bit_n[2] a_19334_1166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1494 VDD rowon_n[13] a_24962_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1495 a_13006_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1496 a_35094_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1497 a_29374_1166# VSS a_28978_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1498 a_28370_5182# rowon_n[3] a_27974_5142# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1499 a_2966_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1500 a_25358_12210# col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1501 VDD rowon_n[7] a_13918_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1502 VDD rowon_n[3] a_14922_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1503 a_7286_4178# rowon_n[2] a_6890_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1504 a_26458_11528# col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1505 a_29982_11166# a_2275_11190# a_30074_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1506 a_6282_8194# rowon_n[6] a_5886_8154# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1507 vcm a_2275_2154# a_7986_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1508 a_24354_18234# col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1509 a_24450_14540# col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1510 a_24050_10162# a_2475_10186# a_23958_10162# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1511 a_2475_9182# a_1957_9182# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.71e+11p pd=1.77e+06u as=0p ps=0u w=600000u l=150000u
X1512 a_22042_1126# a_2475_1150# a_21950_1126# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1513 VSS row_n[8] a_9294_10202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1514 a_12306_6186# col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1515 a_28066_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1516 VDD rowon_n[1] a_27974_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1517 a_32994_18194# a_2275_18218# a_33086_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1518 VSS row_n[14] a_18330_16226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1519 a_23046_16186# a_2475_16210# a_22954_16186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1520 a_24962_10162# row_n[8] a_25454_10524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1521 a_22954_7150# row_n[5] a_23446_7512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1522 VSS row_n[14] a_8290_16226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1523 a_33486_7512# col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1524 VDD rowon_n[2] a_6890_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1525 a_23958_16186# row_n[14] a_24450_16548# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1526 a_20946_2130# row_n[0] a_21438_2492# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1527 a_10906_14178# a_2275_14202# a_10998_14178# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1528 a_18026_14178# a_2475_14202# a_17934_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1529 VDD rowon_n[10] a_7894_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1530 a_31478_2492# col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1531 VDD VDD a_16930_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1532 a_7986_14178# a_2475_14202# a_7894_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1533 VDD VDD a_6890_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1534 a_26362_2170# col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1535 VDD rowon_n[0] a_16930_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1536 a_4274_5182# col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1537 vcm a_2275_9182# a_30074_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1538 a_16322_8194# col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1539 a_17326_4178# col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1540 a_27974_5142# row_n[3] a_28466_5504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1541 vcm a_2275_10186# a_13006_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1542 a_5886_8154# row_n[6] a_6378_8516# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1543 a_2874_14178# row_n[12] a_3366_14540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1544 a_12914_14178# row_n[12] a_13406_14540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1545 a_24354_12210# rowon_n[10] a_23958_12170# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1546 vcm a_2275_10186# a_2966_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1547 a_21950_10162# a_2275_10186# a_22042_10162# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1548 a_32082_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1549 a_28370_11206# rowon_n[9] a_27974_11166# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1550 a_21038_8154# a_2475_8178# a_20946_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1551 a_3878_3134# row_n[1] a_4370_3496# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1552 vcm a_2275_16210# a_12002_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1553 a_14010_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1554 a_15014_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1555 a_16930_4138# row_n[2] a_17422_4500# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1556 a_9994_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1557 a_8290_7190# col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1558 a_9294_3174# col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1559 VDD rowon_n[8] a_23958_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1560 a_9902_7150# a_2275_7174# a_9994_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1561 a_10906_3134# a_2275_3158# a_10998_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1562 VSS row_n[15] a_22346_17230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1563 a_28978_16186# a_2275_16210# a_29070_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1564 a_33086_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1565 VSS row_n[4] a_22346_6186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1566 a_32386_6186# rowon_n[4] a_31990_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1567 a_10998_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1568 a_23350_13214# col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1569 a_26058_6146# a_2475_6170# a_25966_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1570 a_8898_1126# VDD a_9390_1488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1571 a_16322_15222# rowon_n[13] a_15926_15182# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1572 VSS row_n[10] a_13310_12210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1573 a_6282_15222# rowon_n[13] a_5886_15182# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1574 a_2161_14202# sample VDD VDD sky130_fd_pr__pfet_01v8 ad=3.42e+11p pd=2.97e+06u as=0p ps=0u w=1.2e+06u l=150000u
X1575 VSS row_n[10] a_3270_12210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1576 VSS row_n[3] a_11302_5182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1577 a_2874_2130# a_2275_2154# a_2966_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1578 a_22442_15544# col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1579 a_35494_14540# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1580 VSS row_n[9] a_7286_11206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1581 VSS row_n[9] a_17326_11206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1582 a_22042_11166# a_2475_11190# a_21950_11166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1583 a_35094_10162# a_2475_10186# a_35002_10162# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1584 a_14922_5142# a_2275_5166# a_15014_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1585 a_15926_1126# a_2275_1150# a_16018_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1586 a_22954_11166# row_n[9] a_23446_11528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1587 a_2966_10162# a_2475_10186# a_2874_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1588 a_13006_10162# a_2475_10186# a_12914_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1589 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X1590 VSS row_n[2] a_27366_4178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1591 VDD rowon_n[12] a_11910_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1592 a_13406_8516# col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1593 VDD rowon_n[11] a_5886_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1594 VDD rowon_n[11] a_15926_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1595 a_3366_10524# col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1596 a_13406_10524# col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1597 a_11302_17230# col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1598 a_11398_3496# col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1599 vcm a_2275_4162# a_20034_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1600 a_15318_16226# col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1601 vcm a_2275_16210# a_20034_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1602 a_25966_9158# a_2275_9182# a_26058_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1603 VSS row_n[5] a_15318_7190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1604 VSS row_n[1] a_16322_3174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1605 a_30074_4138# a_2475_4162# a_29982_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1606 a_14010_18194# a_2475_18218# a_13918_18194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1607 a_5278_16226# col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1608 vcm a_2275_15206# a_33086_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1609 a_27462_4500# col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1610 a_3970_18194# a_2475_18218# a_3878_18194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1611 a_5374_7512# col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1612 a_31990_6146# row_n[4] a_32482_6508# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1613 a_5978_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1614 a_18426_6508# col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1615 a_12002_5142# a_2475_5166# a_11910_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1616 a_13006_1126# a_2475_1150# a_12914_1126# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1617 a_14410_18556# col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1618 a_10906_15182# row_n[13] a_11398_15544# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1619 a_22346_13214# rowon_n[11] a_21950_13174# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1620 vcm a_2275_11190# a_10998_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1621 VSS row_n[7] a_9294_9198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1622 a_4370_18556# col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1623 a_35398_12210# rowon_n[10] a_35002_12170# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1624 a_3366_2492# col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1625 a_16418_1488# col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1626 a_27062_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1627 a_23958_12170# a_2275_12194# a_24050_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1628 VSS row_n[0] a_8290_2170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1629 a_34394_5182# col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1630 a_34090_6146# a_2475_6170# a_33998_6146# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1631 a_1957_7174# VDD sample VSS sky130_fd_pr__nfet_01v8 ad=1.71e+11p pd=1.77e+06u as=0p ps=0u w=600000u l=150000u
X1632 VDD rowon_n[9] a_21950_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1633 a_9390_9520# col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1634 a_10298_1166# col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1635 a_22346_1166# VSS a_21950_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1636 a_21342_5182# rowon_n[3] a_20946_5142# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1637 VDD rowon_n[8] a_35002_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1638 a_17022_3134# a_2475_3158# a_16930_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1639 VSS VDD a_20338_18234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1640 VSS row_n[15] a_33390_17230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1641 a_33998_3134# row_n[1] a_34490_3496# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1642 a_21342_14218# col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1643 VDD rowon_n[6] a_22954_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1644 a_6890_7150# a_2275_7174# a_6982_7150# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1645 vcm a_2275_5166# a_13006_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1646 vcm a_2275_1150# a_14010_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1647 a_10298_17230# rowon_n[15] a_9902_17190# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1648 a_34394_13214# col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1649 a_28066_17190# a_2475_17214# a_27974_17190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1650 a_4274_16226# rowon_n[14] a_3878_16186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1651 a_14314_16226# rowon_n[14] a_13918_16186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1652 VSS row_n[11] a_11302_13214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1653 a_21038_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1654 VDD rowon_n[1] a_20946_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1655 a_20434_16548# col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1656 a_29982_14178# a_2275_14202# a_30074_14178# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1657 a_28978_17190# row_n[15] a_29470_17552# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1658 a_33486_15544# col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1659 vcm a_2275_13198# a_29070_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1660 a_10998_11166# a_2475_11190# a_10906_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1661 a_33086_11166# a_2475_11190# a_32994_11166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1662 a_20338_9198# col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1663 a_8990_2130# a_2475_2154# a_8898_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1664 a_26362_3174# rowon_n[1] a_25966_3134# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1665 a_5886_15182# a_2275_15206# a_5978_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1666 a_15926_15182# a_2275_15206# a_16018_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1667 VSS row_n[7] a_30378_9198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1668 VDD rowon_n[5] a_11910_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1669 a_4274_6186# rowon_n[4] a_3878_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1670 VDD rowon_n[13] a_9902_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1671 a_33998_11166# row_n[9] a_34490_11528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1672 a_16322_9198# rowon_n[7] a_15926_9158# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1673 vcm a_2275_9182# a_24050_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1674 a_19030_7150# a_2475_7174# a_18938_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1675 a_10298_12210# col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1676 a_11398_11528# col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1677 VDD rowon_n[4] a_27974_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1678 VDD rowon_n[0] a_9902_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1679 vcm a_2275_3158# a_18026_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1680 VDD VSS a_25966_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1681 a_32994_2130# a_2275_2154# a_33086_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1682 a_15318_2170# rowon_n[0] a_14922_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1683 a_26058_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1684 a_19942_9158# row_n[7] a_20434_9520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1685 a_25054_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1686 a_20946_5142# row_n[3] a_21438_5504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1687 vcm a_2275_16210# a_31078_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1688 a_30474_9520# col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1689 a_31478_5504# col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1690 a_9902_10162# row_n[8] a_10394_10524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1691 vcm a_2275_17214# a_17022_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1692 VDD rowon_n[7] a_15926_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1693 a_8290_8194# rowon_n[6] a_7894_8154# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1694 VDD rowon_n[3] a_16930_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1695 a_9294_4178# rowon_n[2] a_8898_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1696 vcm a_2275_17214# a_6982_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1697 a_20338_14218# rowon_n[12] a_19942_14178# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1698 a_21038_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1699 a_14314_6186# col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1700 a_24050_1126# a_2475_1150# a_23958_1126# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1701 a_25054_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1702 a_21950_13174# a_2275_13198# a_22042_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1703 a_24962_7150# row_n[5] a_25454_7512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1704 a_16018_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1705 a_35494_7512# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1706 a_3878_6146# row_n[4] a_4370_6508# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1707 a_5978_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1708 VDD rowon_n[2] a_8898_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1709 a_9994_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1710 VSS row_n[10] a_32386_12210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1711 a_22954_2130# row_n[0] a_23446_2492# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1712 a_33486_2492# col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1713 VSS VDD a_31382_18234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1714 a_2475_11190# a_1957_11190# VDD VDD sky130_fd_pr__pfet_01v8 ad=3.42e+11p pd=2.97e+06u as=0p ps=0u w=1.2e+06u l=150000u
X1715 a_28370_2170# col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1716 a_12002_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1717 VDD rowon_n[12] a_30986_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1718 a_27062_12170# a_2475_12194# a_26970_12170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1719 a_3270_11206# rowon_n[9] a_2874_11166# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1720 a_13310_11206# rowon_n[9] a_12914_11166# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1721 a_6282_5182# col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1722 a_7286_1166# col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1723 a_32386_14218# col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1724 a_19334_4178# col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1725 a_26058_18194# a_2475_18218# a_25966_18194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1726 a_27974_12170# row_n[10] a_28466_12532# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1727 a_32482_10524# col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1728 a_18330_8194# col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1729 VSS row_n[2] a_20338_4178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1730 a_26970_18194# VDD a_27462_18556# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1731 a_30378_17230# col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1732 vcm a_2275_14202# a_27062_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1733 a_7894_8154# row_n[6] a_8386_8516# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1734 a_30378_4178# rowon_n[2] a_29982_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1735 a_13918_16186# a_2275_16210# a_14010_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1736 a_31478_16548# col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1737 vcm a_2275_2154# a_31078_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1738 a_34090_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1739 a_3878_16186# a_2275_16210# a_3970_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1740 a_23046_8154# a_2475_8178# a_22954_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1741 a_3970_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1742 a_5886_3134# row_n[1] a_6378_3496# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1743 a_17022_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1744 vcm a_2275_17214# a_25054_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1745 a_18938_4138# row_n[2] a_19430_4500# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1746 vcm a_2275_11190# a_30074_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1747 a_20434_4500# col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1748 a_29982_15182# row_n[13] a_30474_15544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1749 a_12914_3134# a_2275_3158# a_13006_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1750 VDD rowon_n[2] a_29982_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1751 vcm a_2275_12194# a_16018_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1752 VSS row_n[4] a_24354_6186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1753 vcm a_2275_12194# a_5978_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1754 a_11398_6508# col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1755 a_34394_6186# rowon_n[4] a_33998_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1756 a_18330_14218# rowon_n[12] a_17934_14178# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1757 VSS row_n[8] a_28370_10202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1758 a_19030_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1759 a_28978_11166# a_2275_11190# a_29070_11166# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1760 a_28066_6146# a_2475_6170# a_27974_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1761 a_20034_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1762 a_19030_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1763 VDD rowon_n[10] a_26970_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1764 VSS row_n[3] a_13310_5182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1765 a_4882_2130# a_2275_2154# a_4974_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1766 a_17934_1126# a_2275_1150# a_18026_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1767 a_3366_5504# col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1768 VSS row_n[2] a_29374_4178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1769 a_15414_8516# col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1770 a_16018_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1771 VSS VDD a_29374_18234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1772 a_33390_16226# rowon_n[14] a_32994_16186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1773 a_26362_15222# col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1774 VSS row_n[11] a_30378_13214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1775 VSS a_2161_6170# a_2275_6170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.71e+11p ps=1.77e+06u w=600000u l=150000u
X1776 a_13406_3496# col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1777 a_19334_7190# rowon_n[5] a_18938_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1778 a_31382_7190# col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1779 a_32386_3174# col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1780 a_9294_17230# rowon_n[15] a_8898_17190# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1781 a_35002_15182# a_2275_15206# a_35094_15182# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1782 a_25454_17552# col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1783 a_21950_14178# row_n[12] a_22442_14540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1784 a_25054_13174# a_2475_13198# a_24962_13174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1785 a_7286_10202# col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1786 a_17326_10202# col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1787 vcm a_2275_10186# a_22042_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1788 a_27974_9158# a_2275_9182# a_28066_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1789 VSS row_n[5] a_17326_7190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1790 VSS row_n[1] a_18330_3174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1791 a_32082_4138# a_2475_4162# a_31990_4138# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1792 a_5978_12170# a_2475_12194# a_5886_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1793 a_16018_12170# a_2475_12194# a_15926_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1794 a_33998_6146# row_n[4] a_34490_6508# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1795 a_29470_4500# col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1796 a_29470_16548# col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1797 a_25966_13174# row_n[11] a_26458_13536# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1798 a_30474_11528# col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1799 a_7382_7512# col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1800 a_7986_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1801 a_14010_5142# a_2475_5166# a_13918_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1802 a_15014_1126# a_2475_1150# a_14922_1126# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1803 a_9994_11166# a_2475_11190# a_9902_11166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1804 a_26970_2130# a_2275_2154# a_27062_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1805 VDD rowon_n[13] a_8898_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1806 a_6378_12532# col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1807 a_16418_12532# col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1808 VDD rowon_n[4] a_20946_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1809 a_31990_1126# VDD a_32482_1488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1810 a_5374_2492# col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1811 vcm a_2275_3158# a_10998_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1812 vcm a_2275_7174# a_9994_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1813 a_18426_1488# en_bit_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1814 a_16930_8154# a_2275_8178# a_17022_8154# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1815 a_18330_18234# col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1816 vcm a_2275_18218# a_23046_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1817 VDD VSS VSS sky130_fd_pr__cap_var_lvt w=1.64e+07u l=1.6e+07u
X1818 a_8290_18234# col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1819 a_24354_1166# VSS a_23958_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1820 a_23350_5182# rowon_n[3] a_22954_5142# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1821 a_27062_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1822 VDD rowon_n[3] a_9902_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1823 a_13918_17190# row_n[15] a_14410_17552# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1824 a_25358_15222# rowon_n[13] a_24962_15182# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1825 vcm a_2275_13198# a_14010_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1826 a_2161_9182# sample VSS VSS sky130_fd_pr__nfet_01v8 ad=1.71e+11p pd=1.77e+06u as=0p ps=0u w=600000u l=150000u
X1827 vcm a_2275_2154# a_2966_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1828 a_3878_17190# row_n[15] a_4370_17552# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1829 vcm a_2275_13198# a_3970_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1830 vcm a_2275_1150# a_16018_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1831 a_17934_16186# row_n[14] a_18426_16548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1832 a_29374_14218# rowon_n[12] a_28978_14178# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1833 VSS row_n[9] a_26362_11206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1834 a_8898_7150# a_2275_7174# a_8990_7150# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1835 vcm a_2275_5166# a_15014_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1836 a_7894_16186# row_n[14] a_8386_16548# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1837 a_31078_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1838 a_23046_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1839 VDD rowon_n[1] a_22954_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1840 VDD rowon_n[11] a_24962_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1841 a_28370_3174# rowon_n[1] a_27974_3134# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1842 a_25358_10202# col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1843 VSS row_n[7] a_32386_9198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1844 VDD rowon_n[5] a_13918_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1845 a_6282_6186# rowon_n[4] a_5886_6146# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1846 a_24354_16226# col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1847 vcm a_2275_9182# a_26058_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1848 a_8290_12210# rowon_n[10] a_7894_12170# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1849 a_15926_10162# a_2275_10186# a_16018_10162# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1850 VSS row_n[0] a_31382_2170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1851 a_21342_2170# col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1852 VDD rowon_n[0] a_11910_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1853 a_24450_12532# col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1854 a_5886_10162# a_2275_10186# a_5978_10162# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1855 a_2475_7174# a_1957_7174# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.71e+11p pd=1.77e+06u as=0p ps=0u w=600000u l=150000u
X1856 a_5978_7150# a_2475_7174# a_5886_7150# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1857 a_7286_18234# VDD a_6890_18194# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1858 a_17326_18234# VDD a_16930_18194# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1859 a_11302_8194# col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1860 a_27062_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1861 a_35002_2130# a_2275_2154# a_35094_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1862 VDD VSS a_27974_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1863 a_17326_2170# rowon_n[0] a_16930_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1864 a_28066_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1865 a_12306_4178# col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1866 a_23446_18556# col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1867 a_32994_16186# a_2275_16210# a_33086_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1868 VSS row_n[12] a_18330_14218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1869 a_23046_14178# a_2475_14202# a_22954_14178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1870 a_22954_5142# row_n[3] a_23446_5504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1871 VSS row_n[12] a_8290_14218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1872 a_32482_9520# col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1873 a_33486_5504# col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1874 a_18938_17190# a_2275_17214# a_19030_17190# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1875 a_8898_17190# a_2275_17214# a_8990_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1876 VDD rowon_n[8] a_7894_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1877 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X1878 VDD rowon_n[14] a_16930_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1879 VDD rowon_n[14] a_6890_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1880 a_11910_4138# row_n[2] a_12402_4500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1881 vcm a_2275_12194# a_35094_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1882 a_3270_7190# col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1883 a_4274_3174# col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1884 a_16322_6186# col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1885 vcm a_2275_18218# a_34090_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1886 vcm a_2275_7174# a_6982_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1887 a_12914_12170# row_n[10] a_13406_12532# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1888 a_5886_6146# row_n[4] a_6378_6508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1889 a_2874_12170# row_n[10] a_3366_12532# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1890 a_25054_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1891 a_24354_10202# rowon_n[8] a_23958_10162# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1892 a_16018_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1893 a_21038_6146# a_2475_6170# a_20946_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1894 a_35494_2492# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1895 a_3878_1126# en_C0_n a_4370_1488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1896 a_24962_2130# row_n[0] a_25454_2492# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1897 a_11910_18194# VDD a_12402_18556# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1898 vcm a_2275_14202# a_12002_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1899 a_5978_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1900 VDD rowon_n[12] a_18938_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1901 a_29070_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1902 a_14010_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1903 a_8290_5182# col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1904 a_9294_1166# col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1905 a_28066_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1906 vcm a_2275_17214# a_9994_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1907 a_9902_5142# a_2275_5166# a_9994_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1908 a_10906_1126# a_2275_1150# a_10998_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1909 VSS row_n[2] a_22346_4178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1910 VSS row_n[13] a_22346_15222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1911 a_28978_14178# a_2275_14202# a_29070_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1912 a_32386_4178# rowon_n[2] a_31990_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1913 a_31382_8194# rowon_n[6] a_30986_8154# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1914 vcm a_2275_2154# a_33086_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1915 a_23350_11206# col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1916 a_25054_8154# a_2475_8178# a_24962_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1917 a_26058_4138# a_2475_4162# a_25966_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1918 a_7894_3134# row_n[1] a_8386_3496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1919 VDD rowon_n[15] a_20946_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1920 a_16322_13214# rowon_n[11] a_15926_13174# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1921 VSS row_n[8] a_13310_10202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1922 a_6282_13214# rowon_n[11] a_5886_13174# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1923 a_3878_11166# a_2275_11190# a_3970_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1924 a_13918_11166# a_2275_11190# a_14010_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1925 VSS row_n[8] a_3270_10202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1926 a_20946_9158# a_2275_9182# a_21038_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1927 VSS row_n[5] a_10298_7190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1928 VSS row_n[1] a_11302_3174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1929 a_22442_13536# col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1930 a_35494_12532# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1931 a_31078_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1932 a_14922_3134# a_2275_3158# a_15014_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1933 a_22442_4500# col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1934 a_17934_12170# a_2275_12194# a_18026_12170# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1935 VDD rowon_n[2] a_31990_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1936 a_7894_12170# a_2275_12194# a_7986_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1937 VDD rowon_n[10] a_11910_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1938 a_13406_6508# col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1939 VSS row_n[7] a_4274_9198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1940 a_6890_18194# a_2275_18218# a_6982_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1941 a_16930_18194# a_2275_18218# a_17022_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1942 VDD rowon_n[9] a_5886_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1943 VDD rowon_n[9] a_15926_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1944 VSS VDD a_14314_18234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1945 a_11302_15222# col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1946 a_11398_1488# col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1947 VSS VDD a_4274_18234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1948 a_32082_17190# a_2475_17214# a_31990_17190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1949 VSS row_n[0] a_3270_2170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1950 a_19942_18194# VDD a_20434_18556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1951 a_15318_14218# col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1952 vcm a_2275_14202# a_20034_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1953 VSS row_n[3] a_15318_5182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1954 VSS VDD a_16322_1166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1955 a_32994_17190# row_n[15] a_33486_17552# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1956 a_14010_16186# a_2475_16210# a_13918_16186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1957 a_5278_14218# col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1958 vcm a_2275_13198# a_33086_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1959 a_10394_17552# col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1960 a_3970_16186# a_2475_16210# a_3878_16186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1961 a_4370_9520# col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1962 VDD rowon_n[6] a_18938_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1963 a_30986_8154# row_n[6] a_31478_8516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1964 a_5374_5504# col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1965 a_17422_8516# col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1966 a_5978_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1967 a_12002_3134# a_2475_3158# a_11910_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1968 a_14410_16548# col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1969 a_10906_13174# row_n[11] a_11398_13536# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1970 a_22346_11206# rowon_n[9] a_21950_11166# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1971 a_18026_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1972 analog_in sw ctop VSS sky130_fd_pr__nfet_01v8 ad=1.102e+12p pd=8.76e+06u as=2.7645e+12p ps=2.191e+07u w=1.9e+06u l=220000u
X1973 a_4370_16548# col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1974 a_35398_10202# rowon_n[8] a_35002_10162# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1975 a_15414_3496# col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1976 a_27062_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1977 VSS row_n[7] a_26362_9198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1978 a_33390_7190# col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1979 a_34394_3174# col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1980 a_18026_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1981 a_34090_4138# a_2475_4162# a_33998_4138# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1982 a_7986_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1983 a_1957_5166# VDD sample VSS sky130_fd_pr__nfet_01v8 ad=1.71e+11p pd=1.77e+06u as=0p ps=0u w=600000u l=150000u
X1984 a_9390_7512# col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1985 a_3970_2130# a_2475_2154# a_3878_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1986 a_21342_3174# rowon_n[1] a_20946_3134# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1987 a_35002_10162# a_2275_10186# a_35094_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1988 a_9994_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1989 a_17022_1126# a_2475_1150# a_16930_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1990 a_29374_17230# col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1991 VSS row_n[14] a_20338_16226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1992 VSS row_n[13] a_33390_15222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1993 a_11302_9198# rowon_n[7] a_10906_9158# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1994 a_28978_2130# a_2275_2154# a_29070_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1995 VDD rowon_n[4] a_22954_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1996 a_6890_5142# a_2275_5166# a_6982_5142# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1997 a_7382_2492# col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1998 vcm a_2275_3158# a_13006_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1999 a_10298_15222# rowon_n[13] a_9902_15182# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2000 a_34394_11206# col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2001 a_26458_9520# col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2002 a_18938_8154# a_2275_8178# a_19030_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2003 a_24962_18194# a_2275_18218# a_25054_18194# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2004 VDD VSS a_20946_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2005 a_10298_2170# rowon_n[0] a_9902_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2006 a_21038_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2007 VDD rowon_n[15] a_31990_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2008 a_28066_15182# a_2475_15206# a_27974_15182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2009 a_4274_14218# rowon_n[12] a_3878_14178# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2010 a_14314_14218# rowon_n[12] a_13918_14178# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2011 VSS row_n[9] a_11302_11206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2012 a_20034_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2013 a_28978_15182# row_n[13] a_29470_15544# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2014 a_33486_13536# col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2015 vcm a_2275_11190# a_29070_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2016 VDD rowon_n[3] a_11910_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2017 a_26362_1166# VSS a_25966_1126# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2018 a_5886_13174# a_2275_13198# a_5978_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2019 a_15926_13174# a_2275_13198# a_16018_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2020 VDD rowon_n[7] a_10906_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2021 a_3270_8194# rowon_n[6] a_2874_8154# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2022 a_4274_4178# rowon_n[2] a_3878_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2023 VDD rowon_n[11] a_9902_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2024 vcm a_2275_2154# a_4974_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2025 a_19030_5142# a_2475_5166# a_18938_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2026 a_10298_10202# col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2027 vcm a_2275_1150# a_18026_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2028 a_30074_18194# a_2475_18218# a_29982_18194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2029 a_16018_8154# a_2475_8178# a_15926_8154# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2030 a_19942_7150# row_n[5] a_20434_7512# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2031 a_25054_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2032 a_30986_18194# VDD a_31478_18556# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2033 vcm a_2275_14202# a_31078_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2034 a_30474_7512# col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2035 VDD rowon_n[2] a_3878_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2036 vcm a_2275_15206# a_17022_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2037 VSS row_n[7] a_34394_9198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2038 VDD rowon_n[5] a_15926_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2039 a_8290_6186# rowon_n[4] a_7894_6146# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2040 vcm a_2275_15206# a_6982_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2041 vcm a_2275_9182# a_28066_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2042 a_23350_2170# col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2043 VDD rowon_n[0] a_13918_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2044 a_21038_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2045 VSS row_n[0] a_33390_2170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2046 a_25358_8194# rowon_n[6] a_24962_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2047 a_7986_7150# a_2475_7174# a_7894_7150# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2048 a_14314_4178# col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2049 VSS a_2161_16210# a_2275_16210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.71e+11p ps=1.77e+06u w=600000u l=150000u
X2050 a_25054_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2051 a_13310_8194# col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2052 a_29070_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2053 vcm a_2275_2154# a_27062_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2054 a_24962_5142# row_n[3] a_25454_5504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2055 a_16018_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2056 a_34490_9520# col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2057 a_35494_5504# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2058 a_5978_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2059 a_28370_12210# col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2060 VSS row_n[8] a_32386_10202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2061 a_2874_8154# row_n[6] a_3366_8516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2062 vcm a_2275_8178# a_17022_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2063 a_32994_11166# a_2275_11190# a_33086_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2064 a_31990_7150# a_2275_7174# a_32082_7150# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2065 a_27366_18234# col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2066 VSS row_n[14] a_31382_16226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2067 a_12002_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2068 a_27462_14540# col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2069 VDD rowon_n[10] a_30986_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2070 a_27062_10162# a_2475_10186# a_26970_10162# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2071 a_6282_3174# col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2072 a_13918_4138# row_n[2] a_14410_4500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2073 a_5278_7190# col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2074 a_26058_16186# a_2475_16210# a_25966_16186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2075 a_27974_10162# row_n[8] a_28466_10524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2076 a_18330_6186# col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2077 VDD VDD a_29982_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2078 vcm a_2275_7174# a_8990_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2079 a_26970_16186# row_n[14] a_27462_16548# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2080 a_30378_15222# col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2081 a_7894_6146# row_n[4] a_8386_6508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2082 VDD a_2161_17214# a_2275_17214# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.42e+11p ps=2.97e+06u w=1.2e+06u l=150000u
X2083 a_13918_14178# a_2275_14202# a_14010_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2084 a_3878_14178# a_2275_14202# a_3970_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2085 a_23046_6146# a_2475_6170# a_22954_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2086 a_5886_1126# VDD a_6378_1488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2087 vcm a_2275_15206# a_25054_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2088 a_8990_17190# a_2475_17214# a_8898_17190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2089 a_29982_13174# row_n[11] a_30474_13536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2090 a_12914_1126# a_2275_1150# a_13006_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2091 vcm a_2275_10186# a_16018_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2092 VSS row_n[2] a_24354_4178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2093 a_9390_17552# col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2094 a_5886_14178# row_n[12] a_6378_14540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2095 a_15926_14178# row_n[12] a_16418_14540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2096 a_27366_12210# rowon_n[10] a_26970_12170# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2097 vcm a_2275_10186# a_5978_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2098 a_10394_8516# col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2099 a_10998_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2100 a_33390_8194# rowon_n[6] a_32994_8154# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2101 a_27366_7190# col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2102 a_34394_4178# rowon_n[2] a_33998_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2103 vcm a_2275_2154# a_35094_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2104 a_19030_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2105 a_27062_8154# a_2475_8178# a_26970_8154# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2106 a_28066_4138# a_2475_4162# a_27974_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2107 a_19030_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2108 VDD rowon_n[8] a_26970_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2109 a_22954_9158# a_2275_9182# a_23046_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2110 VSS row_n[5] a_12306_7190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2111 VSS row_n[1] a_13310_3174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2112 a_33086_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2113 VDD rowon_n[2] a_33998_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2114 a_24450_4500# col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2115 VSS row_n[15] a_25358_17230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2116 a_2966_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2117 a_15414_6508# col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2118 a_16018_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2119 a_21950_2130# a_2275_2154# a_22042_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2120 VSS row_n[14] a_29374_16226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2121 a_33390_14218# rowon_n[12] a_32994_14178# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2122 a_26362_13214# col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2123 VSS row_n[9] a_30378_11206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2124 VSS a_2161_4162# a_2275_4162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.71e+11p ps=1.77e+06u w=600000u l=150000u
X2125 a_13406_1488# col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2126 a_12002_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2127 a_34090_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2128 VSS row_n[10] a_16322_12210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2129 a_21038_12170# a_2475_12194# a_20946_12170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2130 a_11910_8154# a_2275_8178# a_12002_8154# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2131 a_32386_1166# col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2132 a_31382_5182# col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2133 a_19334_5182# rowon_n[3] a_18938_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2134 a_9294_15222# rowon_n[13] a_8898_15182# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2135 a_35002_13174# a_2275_13198# a_35094_13174# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2136 VSS row_n[10] a_6282_12210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2137 VSS row_n[0] a_5278_2170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2138 VDD VDD a_27974_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2139 a_25454_15544# col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2140 a_21950_12170# row_n[10] a_22442_12532# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2141 a_25054_11166# a_2475_11190# a_24962_11166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2142 VSS row_n[3] a_17326_5182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2143 VSS en_bit_n[1] a_18330_1166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2144 a_5978_10162# a_2475_10186# a_5886_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2145 a_16018_10162# a_2475_10186# a_15926_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2146 VDD rowon_n[12] a_14922_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2147 a_25966_11166# row_n[9] a_26458_11528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2148 a_32994_8154# row_n[6] a_33486_8516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2149 a_7382_5504# col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2150 a_7986_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2151 a_14010_3134# a_2475_3158# a_13918_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2152 VDD rowon_n[12] a_4882_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2153 VDD rowon_n[11] a_8898_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2154 a_6378_10524# col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2155 a_16418_10524# col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2156 vcm a_2275_1150# a_10998_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2157 a_30986_3134# row_n[1] a_31478_3496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2158 VDD rowon_n[1] a_18938_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2159 a_14314_17230# col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2160 a_3878_7150# a_2275_7174# a_3970_7150# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2161 vcm a_2275_5166# a_9994_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2162 a_4274_17230# col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2163 a_16930_6146# a_2275_6170# a_17022_6146# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2164 a_17422_3496# col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2165 a_18330_16226# col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2166 vcm a_2275_16210# a_23046_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2167 VSS row_n[7] a_28370_9198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2168 a_35398_7190# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2169 a_9902_18194# a_2275_18218# a_9994_18194# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2170 a_17022_18194# a_2475_18218# a_16930_18194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2171 a_8290_16226# col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2172 a_1957_9182# VSS sample VDD sky130_fd_pr__pfet_01v8 ad=3.42e+11p pd=2.97e+06u as=0p ps=0u w=1.2e+06u l=150000u
X2173 a_6982_18194# a_2475_18218# a_6890_18194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2174 a_23350_3174# rowon_n[1] a_22954_3134# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2175 a_17422_18556# col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2176 a_13918_15182# row_n[13] a_14410_15544# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2177 a_25358_13214# rowon_n[11] a_24962_13174# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2178 a_1957_12194# VSS sample VDD sky130_fd_pr__pfet_01v8 ad=3.42e+11p pd=2.97e+06u as=0p ps=0u w=1.2e+06u l=150000u
X2179 vcm a_2275_11190# a_14010_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2180 a_2161_7174# sample VSS VSS sky130_fd_pr__nfet_01v8 ad=1.71e+11p pd=1.77e+06u as=0p ps=0u w=600000u l=150000u
X2181 a_7382_18556# col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2182 a_3878_15182# row_n[13] a_4370_15544# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2183 vcm a_2275_11190# a_3970_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2184 a_13310_9198# rowon_n[7] a_12914_9158# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2185 vcm a_2275_9182# a_21038_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2186 a_31078_9158# a_2475_9182# a_30986_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2187 a_8898_5142# a_2275_5166# a_8990_5142# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2188 a_9390_2492# col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2189 vcm a_2275_3158# a_15014_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2190 a_28466_9520# col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2191 a_26970_12170# a_2275_12194# a_27062_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2192 a_22042_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2193 VDD VSS a_22954_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2194 a_29982_2130# a_2275_2154# a_30074_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2195 a_12306_2170# rowon_n[0] a_11910_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2196 a_23046_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2197 VSS row_n[10] a_24354_12210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2198 VDD rowon_n[9] a_24962_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2199 a_28370_1166# VSS a_27974_1126# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2200 VDD rowon_n[7] a_12914_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2201 VDD rowon_n[3] a_13918_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2202 a_6282_4178# rowon_n[2] a_5886_4138# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2203 VSS VDD a_23350_18234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2204 VDD rowon_n[12] a_22954_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2205 a_24354_14218# col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2206 a_19030_12170# a_2475_12194# a_18938_12170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2207 a_8290_10202# rowon_n[8] a_7894_10162# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2208 a_32082_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2209 a_24450_10524# col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2210 a_2475_5166# a_1957_5166# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.71e+11p pd=1.77e+06u as=0p ps=0u w=600000u l=150000u
X2211 a_5978_5142# a_2475_5166# a_5886_5142# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2212 a_7286_16226# rowon_n[14] a_6890_16186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2213 a_17326_16226# rowon_n[14] a_16930_16186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2214 a_18026_8154# a_2475_8178# a_17934_8154# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2215 a_11302_6186# col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2216 a_27062_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2217 a_23446_16548# col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2218 a_32994_14178# a_2275_14202# a_33086_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2219 a_32482_7512# col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2220 VDD rowon_n[2] a_5886_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2221 a_18938_15182# a_2275_15206# a_19030_15182# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2222 a_8898_15182# a_2275_15206# a_8990_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2223 a_30474_2492# col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2224 a_19942_2130# row_n[0] a_20434_2492# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2225 a_3270_12210# col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2226 a_13310_12210# col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2227 a_25358_2170# col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2228 VDD rowon_n[0] a_15926_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2229 a_12306_18234# col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2230 a_35002_14178# row_n[12] a_35494_14540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2231 vcm a_2275_10186# a_35094_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2232 a_27366_8194# rowon_n[6] a_26970_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2233 a_9994_7150# a_2475_7174# a_9902_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2234 a_3270_5182# col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2235 VSS row_n[0] a_35398_2170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2236 a_4274_1166# en_C0_n VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2237 a_15318_8194# col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2238 vcm a_2275_2154# a_29070_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2239 a_16322_4178# col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2240 vcm a_2275_16210# a_34090_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2241 a_12402_14540# col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2242 a_21038_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2243 vcm a_2275_5166# a_6982_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2244 a_12914_10162# row_n[8] a_13406_10524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2245 a_4882_8154# row_n[6] a_5374_8516# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2246 VSS a_2161_11190# a_2275_11190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.71e+11p ps=1.77e+06u w=600000u l=150000u
X2247 a_2874_10162# row_n[8] a_3366_10524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2248 vcm a_2275_8178# a_19030_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2249 a_20034_8154# a_2475_8178# a_19942_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2250 a_21038_4138# a_2475_4162# a_20946_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2251 a_11910_16186# row_n[14] a_12402_16548# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2252 a_33998_7150# a_2275_7174# a_34090_7150# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2253 a_2874_3134# row_n[1] a_3366_3496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2254 VDD rowon_n[10] a_18938_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2255 a_14010_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2256 a_8290_3174# col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2257 a_15926_4138# row_n[2] a_16418_4500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2258 a_21342_17230# rowon_n[15] a_20946_17190# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2259 a_28066_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2260 vcm a_2275_15206# a_9994_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2261 a_9902_3134# a_2275_3158# a_9994_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2262 VSS row_n[11] a_22346_13214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2263 a_31382_6186# rowon_n[4] a_30986_6146# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2264 VSS row_n[10] a_35398_12210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2265 a_12306_12210# rowon_n[10] a_11910_12170# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2266 a_25054_6146# a_2475_6170# a_24962_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2267 a_7894_1126# VDD a_8386_1488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2268 VDD rowon_n[13] a_20946_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2269 a_6282_11206# rowon_n[9] a_5886_11166# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2270 a_16322_11206# rowon_n[9] a_15926_11166# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2271 a_26970_8154# row_n[6] a_27462_8516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2272 VDD rowon_n[12] a_33998_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2273 VSS row_n[3] a_10298_5182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2274 VSS VDD a_11302_1166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2275 a_22442_11528# col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2276 a_35494_10524# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2277 a_14922_1126# a_2275_1150# a_15014_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2278 a_20338_18234# col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2279 a_33390_17230# col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2280 VDD rowon_n[8] a_11910_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2281 a_12402_8516# col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2282 a_13006_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2283 a_29374_7190# col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2284 VSS row_n[15] a_10298_17230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2285 a_6890_16186# a_2275_16210# a_6982_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2286 a_16930_16186# a_2275_16210# a_17022_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2287 a_29070_8154# a_2475_8178# a_28978_8154# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2288 VSS row_n[14] a_14314_16226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2289 a_11302_13214# col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2290 a_10394_3496# col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2291 vcm a_2275_17214# a_28066_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2292 VSS row_n[14] a_4274_16226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2293 a_32082_15182# a_2475_15206# a_31990_15182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2294 VSS row_n[7] a_21342_9198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2295 a_19942_16186# row_n[14] a_20434_16548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2296 a_19030_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2297 VSS row_n[1] a_15318_3174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2298 a_32994_15182# row_n[13] a_33486_15544# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2299 a_14010_14178# a_2475_14202# a_13918_14178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2300 vcm a_2275_11190# a_33086_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2301 a_24962_9158# a_2275_9182# a_25054_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2302 a_35094_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2303 VSS row_n[5] a_14314_7190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2304 vcm a_2275_7174# a_32082_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2305 VDD VDD a_12914_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2306 a_10394_15544# col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2307 a_3970_14178# a_2475_14202# a_3878_14178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2308 a_4370_7512# col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2309 VDD rowon_n[4] a_18938_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2310 a_30986_6146# row_n[4] a_31478_6508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2311 VDD VDD a_2874_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2312 vcm a_2275_12194# a_8990_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2313 vcm a_2275_12194# a_19030_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2314 a_4974_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2315 a_17422_6508# col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2316 a_12002_1126# a_2475_1150# a_11910_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2317 a_5978_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2318 a_10906_11166# row_n[9] a_11398_11528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2319 VDD a_2161_8178# a_2275_8178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.42e+11p ps=2.97e+06u w=1.2e+06u l=150000u
X2320 a_18026_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2321 a_23958_2130# a_2275_2154# a_24050_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2322 ctop sw analog_in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.9e+06u l=220000u
X2323 a_23046_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2324 a_21438_9520# col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2325 a_13918_8154# a_2275_8178# a_14010_8154# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2326 a_15414_1488# col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2327 VSS row_n[0] a_7286_2170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2328 a_33390_5182# col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2329 a_1957_3158# VDD sample VSS sky130_fd_pr__nfet_01v8 ad=1.71e+11p pd=1.77e+06u as=0p ps=0u w=600000u l=150000u
X2330 a_32386_17230# rowon_n[15] a_31990_17190# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2331 a_35002_8154# row_n[6] a_35494_8516# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2332 a_9390_5504# col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2333 a_21342_1166# VSS a_20946_1126# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2334 a_9994_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2335 a_29374_15222# col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2336 VSS row_n[12] a_20338_14218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2337 VSS row_n[11] a_33390_13214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2338 a_20946_17190# a_2275_17214# a_21038_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2339 a_5886_7150# a_2275_7174# a_5978_7150# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2340 vcm a_2275_1150# a_13006_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2341 a_32994_3134# row_n[1] a_33486_3496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2342 a_6890_3134# a_2275_3158# a_6982_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2343 a_10298_13214# rowon_n[11] a_9902_13174# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2344 a_26458_7512# col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2345 a_18938_6146# a_2275_6170# a_19030_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2346 a_24962_16186# a_2275_16210# a_25054_16186# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2347 a_8990_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2348 a_28466_17552# col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2349 VDD rowon_n[13] a_31990_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2350 a_28066_13174# a_2475_13198# a_27974_13174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2351 a_10998_8154# a_2475_8178# a_10906_8154# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2352 a_20034_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2353 a_11910_12170# a_2275_12194# a_12002_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2354 a_28978_13174# row_n[11] a_29470_13536# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2355 a_33486_11528# col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2356 VDD rowon_n[9] a_9902_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2357 VDD rowon_n[5] a_10906_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2358 a_3270_6186# rowon_n[4] a_2874_6146# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2359 a_31382_18234# col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2360 vcm a_2275_9182# a_23046_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2361 a_19030_3134# a_2475_3158# a_18938_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2362 a_33086_9158# a_2475_9182# a_32994_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2363 vcm a_2275_18218# a_26058_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2364 a_30074_16186# a_2475_16210# a_29982_16186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2365 a_20338_8194# rowon_n[6] a_19942_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2366 a_2966_7150# a_2475_7174# a_2874_7150# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2367 a_24050_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2368 a_16018_6146# a_2475_6170# a_15926_6146# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2369 vcm a_2275_2154# a_22042_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2370 a_14314_2170# rowon_n[0] a_13918_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2371 a_25054_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2372 a_19942_5142# row_n[3] a_20434_5504# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2373 a_30986_16186# row_n[14] a_31478_16548# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2374 a_30474_5504# col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2375 vcm a_2275_8178# a_12002_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2376 a_16930_17190# row_n[15] a_17422_17552# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2377 vcm a_2275_13198# a_17022_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2378 VDD rowon_n[3] a_15926_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2379 a_8290_4178# rowon_n[2] a_7894_4138# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2380 a_6890_17190# row_n[15] a_7382_17552# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2381 vcm a_2275_13198# a_6982_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2382 a_21038_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2383 a_2475_9182# a_1957_9182# VDD VDD sky130_fd_pr__pfet_01v8 ad=3.42e+11p pd=2.97e+06u as=0p ps=0u w=1.2e+06u l=150000u
X2384 a_25358_6186# rowon_n[4] a_24962_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2385 a_7986_5142# a_2475_5166# a_7894_5142# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2386 VSS a_2161_14202# a_2275_14202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.71e+11p ps=1.77e+06u w=600000u l=150000u
X2387 a_13310_6186# col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2388 a_29070_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2389 a_31382_12210# rowon_n[10] a_30986_12170# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2390 vcm a_2275_7174# a_3970_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2391 a_34490_7512# col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2392 a_2874_6146# row_n[4] a_3366_6508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2393 a_28370_10202# col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2394 vcm a_2275_6170# a_17022_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2395 VDD rowon_n[2] a_7894_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2396 a_30378_18234# VDD a_29982_18194# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2397 a_19942_12170# a_2275_12194# a_20034_12170# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2398 a_32482_2492# col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2399 a_31990_5142# a_2275_5166# a_32082_5142# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2400 a_27366_16226# col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2401 VSS row_n[12] a_31382_14218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2402 a_18938_10162# a_2275_10186# a_19030_10162# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2403 a_31990_17190# a_2275_17214# a_32082_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2404 a_27462_12532# col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2405 a_8898_10162# a_2275_10186# a_8990_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2406 VDD rowon_n[8] a_30986_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2407 VSS row_n[6] a_19334_8194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2408 a_6282_1166# col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2409 a_29374_8194# rowon_n[6] a_28978_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2410 a_5278_5182# col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2411 a_26058_14178# a_2475_14202# a_25966_14178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2412 a_18330_4178# col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2413 a_26458_18556# col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2414 VDD rowon_n[14] a_29982_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2415 vcm a_2275_5166# a_8990_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2416 a_30378_13214# col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2417 a_22346_7190# col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2418 VDD a_2161_15206# a_2275_15206# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.42e+11p ps=2.97e+06u w=1.2e+06u l=150000u
X2419 vcm a_2275_2154# a_30074_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2420 VSS row_n[15] a_9294_17230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2421 a_24050_17190# a_2475_17214# a_23958_17190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2422 a_22042_8154# a_2475_8178# a_21950_8154# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2423 a_4882_3134# row_n[1] a_5374_3496# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2424 a_23046_4138# a_2475_4162# a_22954_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2425 vcm a_2275_13198# a_25054_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2426 a_24962_17190# row_n[15] a_25454_17552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2427 a_17934_4138# row_n[2] a_18426_4500# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2428 a_8990_15182# a_2475_15206# a_8898_15182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2429 a_29982_11166# row_n[9] a_30474_11528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2430 a_9390_15544# col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2431 a_5886_12170# row_n[10] a_6378_12532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2432 a_15926_12170# row_n[10] a_16418_12532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2433 a_28066_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2434 a_27366_10202# rowon_n[8] a_26970_10162# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2435 a_10394_6508# col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2436 a_10998_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2437 a_33390_6186# rowon_n[4] a_32994_6146# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2438 a_27366_5182# col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2439 a_19030_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2440 a_27062_6146# a_2475_6170# a_26970_6146# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2441 a_28978_8154# row_n[6] a_29470_8516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2442 a_19030_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2443 vcm a_2275_17214# a_13006_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2444 VSS row_n[3] a_12306_5182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2445 VSS VDD a_13310_1166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2446 vcm a_2275_17214# a_2966_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2447 a_26970_3134# row_n[1] a_27462_3496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2448 a_28370_18234# VDD a_27974_18194# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2449 VSS row_n[13] a_25358_15222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2450 a_22346_12210# col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2451 a_2966_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2452 a_14410_8516# col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2453 a_16018_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2454 VSS row_n[12] a_29374_14218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2455 a_26362_11206# col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2456 a_15014_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2457 VSS a_2161_2154# a_2275_2154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.71e+11p ps=1.77e+06u w=600000u l=150000u
X2458 VDD rowon_n[15] a_23958_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2459 a_12002_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2460 a_34090_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2461 a_21438_14540# col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2462 a_30986_12170# a_2275_12194# a_31078_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2463 VSS row_n[8] a_16322_10202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2464 a_21038_10162# a_2475_10186# a_20946_10162# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2465 a_18330_7190# rowon_n[5] a_17934_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2466 a_11910_6146# a_2275_6170# a_12002_6146# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2467 a_31382_3174# col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2468 a_19334_3174# rowon_n[1] a_18938_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2469 a_12402_3496# col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2470 a_9294_13214# rowon_n[11] a_8898_13174# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2471 a_6890_11166# a_2275_11190# a_6982_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2472 a_16930_11166# a_2275_11190# a_17022_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2473 VSS row_n[8] a_6282_10202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2474 VSS row_n[7] a_23350_9198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2475 a_30378_7190# col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2476 VDD rowon_n[14] a_27974_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2477 a_25454_13536# col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2478 a_21950_10162# row_n[8] a_22442_10524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2479 VSS row_n[1] a_17326_3174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2480 vcm a_2275_7174# a_34090_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2481 a_32994_6146# row_n[4] a_33486_6508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2482 VDD rowon_n[10] a_14922_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2483 a_14010_1126# a_2475_1150# a_13918_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2484 a_7986_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2485 VDD rowon_n[10] a_4882_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2486 a_6982_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2487 a_25966_2130# a_2275_2154# a_26058_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2488 VDD rowon_n[9] a_8898_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2489 VDD en_bit_n[2] a_18938_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2490 a_30986_1126# VDD a_31478_1488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2491 VSS VDD a_17326_18234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2492 a_22042_18194# a_2475_18218# a_21950_18194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2493 a_14314_15222# col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2494 a_3878_5142# a_2275_5166# a_3970_5142# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2495 a_4370_2492# col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2496 vcm a_2275_3158# a_9994_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2497 VSS VDD a_7286_18234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2498 a_13006_17190# a_2475_17214# a_12914_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2499 a_35094_17190# a_2475_17214# a_35002_17190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2500 a_4274_15222# col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2501 a_23446_9520# col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2502 a_15926_8154# a_2275_8178# a_16018_8154# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2503 a_17422_1488# col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2504 a_16930_4138# a_2275_4162# a_17022_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2505 a_22954_18194# VDD a_23446_18556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2506 a_2966_17190# a_2475_17214# a_2874_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2507 a_18330_14218# col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2508 vcm a_2275_14202# a_23046_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2509 VSS row_n[0] a_9294_2170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2510 a_35398_5182# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2511 a_9902_16186# a_2275_16210# a_9994_16186# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2512 a_17022_16186# a_2475_16210# a_16930_16186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2513 a_8290_14218# col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2514 a_13406_17552# col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2515 a_6982_16186# a_2475_16210# a_6890_16186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2516 a_23350_1166# VSS a_22954_1126# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2517 a_3366_17552# col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2518 a_17422_16548# col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2519 a_13918_13174# row_n[11] a_14410_13536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2520 a_25358_11206# rowon_n[9] a_24962_11166# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2521 a_1957_10186# VSS sample VDD sky130_fd_pr__pfet_01v8 ad=3.42e+11p pd=2.97e+06u as=0p ps=0u w=1.2e+06u l=150000u
X2522 a_2161_5166# sample VSS VSS sky130_fd_pr__nfet_01v8 ad=1.71e+11p pd=1.77e+06u as=0p ps=0u w=600000u l=150000u
X2523 a_7382_16548# col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2524 a_3878_13174# row_n[11] a_4370_13536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2525 a_35002_3134# row_n[1] a_35494_3496# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2526 a_7894_7150# a_2275_7174# a_7986_7150# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2527 vcm a_2275_1150# a_15014_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2528 a_8898_3134# a_2275_3158# a_8990_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2529 a_28466_7512# col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2530 a_13006_8154# a_2475_8178# a_12914_8154# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2531 a_22042_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2532 ctop sw_n analog_in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.102e+12p ps=8.76e+06u w=1.9e+06u l=220000u
X2533 VSS row_n[8] a_24354_10202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2534 a_26458_2492# col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2535 vcm a_2275_18218# a_10998_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2536 a_24962_11166# a_2275_11190# a_25054_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2537 VDD rowon_n[5] a_12914_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2538 VSS row_n[14] a_23350_16226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2539 a_19430_14540# col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2540 VDD rowon_n[10] a_22954_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2541 a_19030_10162# a_2475_10186# a_18938_10162# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2542 vcm a_2275_9182# a_25054_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2543 a_35094_9158# a_2475_9182# a_35002_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2544 a_20338_2170# col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2545 VDD rowon_n[0] a_10906_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2546 a_27974_18194# a_2275_18218# a_28066_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2547 a_32082_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2548 a_22346_8194# rowon_n[6] a_21950_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2549 a_4974_7150# a_2475_7174# a_4882_7150# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2550 VSS row_n[0] a_30378_2170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2551 a_5978_3134# a_2475_3158# a_5886_3134# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2552 a_2475_3158# a_1957_3158# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.71e+11p pd=1.77e+06u as=0p ps=0u w=600000u l=150000u
X2553 VDD VDD a_21950_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2554 VDD rowon_n[15] a_35002_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2555 a_7286_14218# rowon_n[12] a_6890_14178# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2556 a_17326_14218# rowon_n[12] a_16930_14178# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2557 a_10298_8194# col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2558 a_18026_6146# a_2475_6170# a_17934_6146# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2559 vcm a_2275_2154# a_24050_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2560 a_16322_2170# rowon_n[0] a_15926_2130# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2561 a_27062_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2562 a_11302_4178# col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2563 analog_in sw_n ctop VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.9e+06u l=220000u
X2564 a_32482_5504# col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2565 a_8898_13174# a_2275_13198# a_8990_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2566 a_18938_13174# a_2275_13198# a_19030_13174# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2567 vcm a_2275_8178# a_14010_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2568 a_34090_12170# a_2475_12194# a_33998_12170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2569 a_3270_10202# col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2570 a_13310_10202# col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2571 a_12002_12170# a_2475_12194# a_11910_12170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2572 a_12306_16226# col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2573 a_35002_12170# row_n[10] a_35494_12532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2574 a_27366_6186# rowon_n[4] a_26970_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2575 a_9994_5142# a_2475_5166# a_9902_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2576 a_3270_3174# col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2577 a_10906_4138# row_n[2] a_11398_4500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2578 a_10998_18194# a_2475_18218# a_10906_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2579 a_33086_18194# a_2475_18218# a_32994_18194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2580 a_5278_9198# rowon_n[7] a_4882_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2581 a_15318_6186# col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2582 a_33998_18194# VDD a_34490_18556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2583 vcm a_2275_14202# a_34090_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2584 a_12402_12532# col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2585 a_19334_12210# rowon_n[10] a_18938_12170# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2586 vcm a_2275_3158# a_6982_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2587 vcm a_2275_7174# a_5978_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2588 a_4882_6146# row_n[4] a_5374_6508# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2589 a_11398_18556# col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2590 vcm a_2275_6170# a_19030_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2591 a_20034_6146# a_2475_6170# a_19942_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2592 a_34490_2492# col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2593 a_2874_1126# VDD a_3366_1488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2594 a_33998_5142# a_2275_5166# a_34090_5142# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2595 VDD rowon_n[8] a_18938_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2596 a_21950_8154# row_n[6] a_22442_8516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2597 a_2475_17214# a_1957_17214# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.71e+11p pd=1.77e+06u as=0p ps=0u w=600000u l=150000u
X2598 VDD rowon_n[7] a_4882_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2599 a_8290_1166# col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2600 a_9902_17190# row_n[15] a_10394_17552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2601 a_21342_15222# rowon_n[13] a_20946_15182# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2602 a_28066_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2603 vcm a_2275_13198# a_9994_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2604 a_9902_1126# a_2275_1150# a_9994_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2605 VSS row_n[9] a_22346_11206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2606 a_31382_4178# rowon_n[2] a_30986_4138# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2607 VSS row_n[8] a_35398_10202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2608 a_24354_7190# col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2609 a_12306_10202# rowon_n[8] a_11910_10162# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2610 a_24050_8154# a_2475_8178# a_23958_8154# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2611 a_25054_4138# a_2475_4162# a_24962_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2612 VDD rowon_n[11] a_20946_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2613 a_26970_6146# row_n[4] a_27462_6508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2614 VDD rowon_n[10] a_33998_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2615 VSS row_n[1] a_10298_3174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2616 a_19942_9158# a_2275_9182# a_20034_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2617 a_30074_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2618 a_20338_16226# col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2619 VDD rowon_n[2] a_30986_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2620 a_2475_18218# a_1957_18218# VDD VDD sky130_fd_pr__pfet_01v8 ad=3.42e+11p pd=2.97e+06u as=0p ps=0u w=1.2e+06u l=150000u
X2621 a_33390_15222# col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2622 a_12402_6508# col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2623 a_16930_14178# a_2275_14202# a_17022_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2624 a_13006_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2625 a_29374_5182# col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2626 a_3270_18234# VDD a_2874_18194# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2627 a_13310_18234# VDD a_12914_18194# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2628 VSS row_n[13] a_10298_15222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2629 a_6890_14178# a_2275_14202# a_6982_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2630 a_7286_8194# col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2631 a_29070_6146# a_2475_6170# a_28978_6146# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2632 VSS row_n[12] a_14314_14218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2633 a_11302_11206# col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2634 a_10394_1488# col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2635 a_32482_17552# col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2636 vcm a_2275_15206# a_28066_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2637 VSS row_n[12] a_4274_14218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2638 a_32082_13174# a_2475_13198# a_31990_13174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2639 a_4882_17190# a_2275_17214# a_4974_17190# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2640 a_14922_17190# a_2275_17214# a_15014_17190# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2641 VSS row_n[3] a_14314_5182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2642 VSS VDD a_15318_1166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2643 a_32994_13174# row_n[11] a_33486_13536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2644 a_28978_3134# row_n[1] a_29470_3496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2645 vcm a_2275_5166# a_32082_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2646 VDD rowon_n[14] a_12914_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2647 a_10394_13536# col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2648 vcm a_2275_10186# a_19030_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2649 VDD rowon_n[6] a_17934_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2650 a_29982_8154# row_n[6] a_30474_8516# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2651 a_4370_5504# col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2652 VDD rowon_n[14] a_2874_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2653 a_8898_14178# row_n[12] a_9390_14540# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2654 a_18938_14178# row_n[12] a_19430_14540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2655 vcm a_2275_10186# a_8990_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2656 a_4974_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2657 a_5978_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2658 a_17022_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2659 VDD a_2161_6170# a_2275_6170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.42e+11p ps=2.97e+06u w=1.2e+06u l=150000u
X2660 a_18026_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2661 vcm a_2275_18218# a_30074_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2662 a_21438_7512# col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2663 a_13918_6146# a_2275_6170# a_14010_6146# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2664 analog_in sw ctop VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.9e+06u l=220000u
X2665 a_14410_3496# col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2666 a_33390_3174# col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2667 VSS row_n[7] a_25358_9198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2668 a_35398_9198# rowon_n[7] a_35002_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2669 a_12002_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2670 a_34090_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2671 VSS row_n[15] a_28370_17230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2672 a_32386_15222# rowon_n[13] a_31990_15182# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2673 a_35002_6146# row_n[4] a_35494_6508# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2674 a_8990_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2675 a_9994_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2676 a_29374_13214# col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2677 VSS row_n[9] a_33390_11206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2678 a_27974_2130# a_2275_2154# a_28066_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2679 a_24050_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2680 a_20946_15182# a_2275_15206# a_21038_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2681 a_5886_5142# a_2275_5166# a_5978_5142# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2682 a_6890_1126# a_2275_1150# a_6982_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2683 a_32994_1126# VDD a_33486_1488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2684 a_15014_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2685 a_10298_11206# rowon_n[9] a_9902_11166# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2686 a_25454_9520# col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2687 a_17934_8154# a_2275_8178# a_18026_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2688 a_18938_4138# a_2275_4162# a_19030_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2689 a_26458_5504# col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2690 a_4974_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2691 a_24962_14178# a_2275_14202# a_25054_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2692 VDD rowon_n[7] a_35002_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2693 a_8990_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2694 a_28466_15544# col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2695 VDD rowon_n[11] a_31990_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2696 a_28066_11166# a_2475_11190# a_27974_11166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2697 a_10998_6146# a_2475_6170# a_10906_6146# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2698 a_20034_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2699 a_28978_11166# row_n[9] a_29470_11528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2700 a_9902_11166# a_2275_11190# a_9994_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2701 a_2161_9182# sample VDD VDD sky130_fd_pr__pfet_01v8 ad=3.42e+11p pd=2.97e+06u as=0p ps=0u w=1.2e+06u l=150000u
X2702 VDD rowon_n[3] a_10906_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2703 a_3270_4178# rowon_n[2] a_2874_4138# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2704 a_31382_16226# col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2705 VSS row_n[5] a_6282_7190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2706 a_19030_1126# a_2475_1150# a_18938_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2707 vcm a_2275_17214# a_22042_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2708 a_7286_17230# col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2709 a_17326_17230# col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2710 vcm a_2275_16210# a_26058_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2711 a_30074_14178# a_2475_14202# a_29982_14178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2712 a_20338_6186# rowon_n[4] a_19942_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2713 a_2966_5142# a_2475_5166# a_2874_5142# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2714 a_12914_18194# a_2275_18218# a_13006_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2715 a_30474_18556# col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2716 a_15014_8154# a_2475_8178# a_14922_8154# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2717 a_24050_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2718 a_16018_4138# a_2475_4162# a_15926_4138# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2719 a_2874_18194# a_2275_18218# a_2966_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2720 a_9994_18194# a_2475_18218# a_9902_18194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2721 a_28466_2492# col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2722 vcm a_2275_6170# a_12002_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2723 VDD rowon_n[2] a_2874_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2724 a_16930_15182# row_n[13] a_17422_15544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2725 vcm a_2275_11190# a_17022_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2726 a_6890_15182# row_n[13] a_7382_15544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2727 vcm a_2275_11190# a_6982_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2728 VDD rowon_n[0] a_12914_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2729 VSS row_n[0] a_32386_2170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2730 a_24354_8194# rowon_n[6] a_23958_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2731 a_6982_7150# a_2475_7174# a_6890_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2732 a_7986_3134# a_2475_3158# a_7894_3134# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2733 a_25358_4178# rowon_n[2] a_24962_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2734 VSS row_n[10] a_27366_12210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2735 vcm a_2275_2154# a_26058_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2736 a_29070_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2737 a_13310_4178# col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2738 a_32082_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2739 a_31382_10202# rowon_n[8] a_30986_10162# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2740 vcm a_2275_5166# a_3970_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2741 a_34490_5504# col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2742 vcm a_2275_8178# a_16018_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2743 vcm a_2275_4162# a_17022_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2744 VSS VDD a_26362_18234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2745 a_30378_16226# rowon_n[14] a_29982_16186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2746 VDD rowon_n[12] a_25966_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2747 a_14010_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2748 a_30986_7150# a_2275_7174# a_31078_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2749 a_31990_3134# a_2275_3158# a_32082_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2750 a_27366_14218# col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2751 a_3970_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2752 VDD rowon_n[2] a_24962_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2753 a_35094_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2754 a_31990_15182# a_2275_15206# a_32082_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2755 a_27462_10524# col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2756 VSS row_n[4] a_19334_6186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2757 a_12914_4138# row_n[2] a_13406_4500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2758 a_2966_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2759 a_13006_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2760 a_29374_6186# rowon_n[4] a_28978_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2761 a_5278_3174# col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2762 a_25358_17230# col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2763 a_26458_16548# col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2764 a_7286_9198# rowon_n[7] a_6890_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2765 vcm a_2275_7174# a_7986_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2766 vcm a_2275_3158# a_8990_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2767 a_30378_11206# col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2768 ctop sw analog_in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.9e+06u l=220000u
X2769 a_22346_5182# col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2770 VDD a_2161_13198# a_2275_13198# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.42e+11p ps=2.97e+06u w=1.2e+06u l=150000u
X2771 VSS row_n[13] a_9294_15222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2772 a_24050_15182# a_2475_15206# a_23958_15182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2773 a_6282_12210# col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2774 a_16322_12210# col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2775 vcm a_2275_12194# a_21038_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2776 a_22042_6146# a_2475_6170# a_21950_6146# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2777 a_4882_1126# VDD a_5374_1488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2778 vcm a_2275_11190# a_25054_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2779 a_23958_8154# row_n[6] a_24450_8516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2780 a_24962_15182# row_n[13] a_25454_15544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2781 a_8990_13174# a_2475_13198# a_8898_13174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2782 VDD rowon_n[7] a_6890_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2783 VDD rowon_n[15] a_7894_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2784 a_5374_14540# col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2785 a_15414_14540# col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2786 a_21950_3134# row_n[1] a_22442_3496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2787 a_9390_13536# col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2788 a_2475_12194# a_1957_12194# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.71e+11p pd=1.77e+06u as=0p ps=0u w=600000u l=150000u
X2789 a_5886_10162# row_n[8] a_6378_10524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2790 a_15926_10162# row_n[8] a_16418_10524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2791 a_26362_7190# col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2792 a_27366_3174# col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2793 a_33390_4178# rowon_n[2] a_32994_4138# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2794 a_10998_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2795 a_17326_9198# col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2796 a_27062_4138# a_2475_4162# a_26970_4138# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2797 a_28978_6146# row_n[4] a_29470_6508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2798 a_24354_17230# rowon_n[15] a_23958_17190# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2799 vcm a_2275_15206# a_13006_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2800 VDD VSS VSS sky130_fd_pr__cap_var_lvt w=1.64e+07u l=1.6e+07u
X2801 VSS row_n[1] a_12306_3174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2802 vcm a_2275_15206# a_2966_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2803 a_32082_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2804 a_26970_1126# VDD a_27462_1488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2805 a_2161_18218# sample VSS VSS sky130_fd_pr__nfet_01v8 ad=1.71e+11p pd=1.77e+06u as=0p ps=0u w=600000u l=150000u
X2806 a_28370_16226# rowon_n[14] a_27974_16186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2807 VSS row_n[11] a_25358_13214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2808 a_22346_10202# col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2809 a_2966_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2810 VDD rowon_n[2] a_32994_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2811 a_14410_6508# col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2812 a_20946_2130# a_2275_2154# a_21038_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2813 a_15318_12210# rowon_n[10] a_14922_12170# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2814 a_16930_9158# row_n[7] a_17422_9520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2815 a_9294_8194# col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2816 a_15014_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2817 a_31078_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2818 a_5278_12210# rowon_n[10] a_4882_12170# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2819 VDD rowon_n[13] a_23958_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2820 a_12002_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2821 a_34090_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2822 a_21438_12532# col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2823 a_10906_8154# a_2275_8178# a_10998_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2824 a_18330_5182# rowon_n[3] a_17934_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2825 a_12402_1488# col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2826 a_19334_1166# en_bit_n[2] a_18938_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2827 a_31382_1166# col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2828 a_11910_4138# a_2275_4162# a_12002_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2829 a_9294_11206# rowon_n[9] a_8898_11166# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2830 VSS row_n[0] a_4274_2170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2831 a_30378_5182# col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2832 a_25454_11528# col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2833 VSS VDD a_17326_1166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2834 a_23350_18234# col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2835 vcm a_2275_5166# a_34090_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2836 VDD rowon_n[8] a_14922_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2837 a_7986_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2838 VDD rowon_n[8] a_4882_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2839 a_6982_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2840 VSS row_n[15] a_3270_17230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2841 VSS row_n[15] a_13310_17230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2842 a_29982_3134# row_n[1] a_30474_3496# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2843 VDD rowon_n[1] a_17934_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2844 VSS row_n[14] a_17326_16226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2845 a_22042_16186# a_2475_16210# a_21950_16186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2846 a_14314_13214# col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2847 a_2874_7150# a_2275_7174# a_2966_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2848 vcm a_2275_1150# a_9994_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2849 a_3878_3134# a_2275_3158# a_3970_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2850 VSS row_n[14] a_7286_16226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2851 a_13006_15182# a_2475_15206# a_12914_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2852 a_35094_15182# a_2475_15206# a_35002_15182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2853 a_4274_13214# col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2854 vcm a_2275_12194# a_32082_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2855 a_23446_7512# col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2856 a_15926_6146# a_2275_6170# a_16018_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2857 a_22954_16186# row_n[14] a_23446_16548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2858 a_2966_15182# a_2475_15206# a_2874_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2859 VSS row_n[7] a_27366_9198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2860 a_35398_3174# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2861 a_9902_14178# a_2275_14202# a_9994_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2862 a_17022_14178# a_2475_14202# a_16930_14178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2863 a_21438_2492# col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2864 VDD VDD a_15926_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2865 a_13406_15544# col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2866 a_6982_14178# a_2475_14202# a_6890_14178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2867 VDD VDD a_5886_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2868 a_3366_15544# col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2869 VSS row_n[0] a_26362_2170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2870 a_2161_3158# sample VSS VSS sky130_fd_pr__nfet_01v8 ad=1.71e+11p pd=1.77e+06u as=0p ps=0u w=600000u l=150000u
X2871 a_13918_11166# row_n[9] a_14410_11528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2872 a_3878_11166# row_n[9] a_4370_11528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2873 vcm a_2275_9182# a_20034_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2874 a_35002_1126# VDD a_35494_1488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2875 a_26058_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2876 a_30074_9158# a_2475_9182# a_29982_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2877 VSS row_n[6] a_16322_8194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2878 a_7894_5142# a_2275_5166# a_7986_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2879 a_8898_1126# a_2275_1150# a_8990_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2880 a_27462_9520# col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2881 a_28466_5504# col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2882 a_23350_12210# rowon_n[10] a_22954_12170# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2883 a_20946_10162# a_2275_10186# a_21038_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2884 a_6378_8516# col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2885 a_13006_6146# a_2475_6170# a_12914_6146# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2886 a_11302_2170# rowon_n[0] a_10906_2130# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2887 a_22042_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2888 a_22346_18234# VDD a_21950_18194# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2889 vcm a_2275_16210# a_10998_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2890 a_35398_17230# rowon_n[15] a_35002_17190# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2891 VDD rowon_n[3] a_12914_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2892 VSS row_n[12] a_23350_14218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2893 a_8990_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2894 a_23958_17190# a_2275_17214# a_24050_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2895 a_19430_12532# col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2896 VDD rowon_n[8] a_22954_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2897 VSS row_n[5] a_8290_7190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2898 a_27974_16186# a_2275_16210# a_28066_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2899 a_32082_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2900 a_22346_6186# rowon_n[4] a_21950_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2901 a_4974_5142# a_2475_5166# a_4882_5142# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2902 a_5978_1126# a_2475_1150# a_5886_1126# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2903 VDD rowon_n[14] a_21950_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2904 VDD rowon_n[13] a_35002_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2905 a_10298_6186# col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2906 a_18026_4138# a_2475_4162# a_17934_4138# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2907 a_35398_12210# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2908 a_17022_8154# a_2475_8178# a_16930_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2909 VSS row_n[10] a_12306_12210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2910 vcm a_2275_6170# a_14010_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2911 a_34394_18234# col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2912 VSS VDD a_11302_18234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2913 a_34490_14540# col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2914 a_34090_10162# a_2475_10186# a_33998_10162# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2915 a_12002_10162# a_2475_10186# a_11910_10162# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2916 vcm a_2275_18218# a_29070_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2917 VDD rowon_n[12] a_10906_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2918 a_12306_14218# col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2919 a_35002_10162# row_n[8] a_35494_10524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2920 VSS row_n[0] a_34394_2170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2921 a_3270_1166# col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2922 a_9994_3134# a_2475_3158# a_9902_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2923 a_27366_4178# rowon_n[2] a_26970_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2924 a_10998_16186# a_2475_16210# a_10906_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2925 a_33086_16186# a_2475_16210# a_32994_16186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2926 a_19334_10202# rowon_n[8] a_18938_10162# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2927 a_26362_8194# rowon_n[6] a_25966_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2928 a_8990_7150# a_2475_7174# a_8898_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2929 vcm a_2275_2154# a_28066_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2930 a_15318_4178# col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2931 a_33998_16186# row_n[14] a_34490_16548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2932 a_12402_10524# col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2933 vcm a_2275_1150# a_6982_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2934 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X2935 a_10298_17230# col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2936 vcm a_2275_5166# a_5978_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2937 a_11398_16548# col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2938 vcm a_2275_8178# a_18026_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2939 vcm a_2275_4162# a_19030_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2940 a_20034_4138# a_2475_4162# a_19942_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2941 a_26058_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2942 a_15318_7190# rowon_n[5] a_14922_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2943 a_32994_7150# a_2275_7174# a_33086_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2944 a_33998_3134# a_2275_3158# a_34090_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2945 a_21950_6146# row_n[4] a_22442_6508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2946 VDD rowon_n[2] a_26970_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2947 a_2475_15206# a_1957_15206# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.71e+11p pd=1.77e+06u as=0p ps=0u w=600000u l=150000u
X2948 VDD rowon_n[5] a_4882_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2949 a_14922_4138# row_n[2] a_15414_4500# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2950 a_9902_15182# row_n[13] a_10394_15544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2951 a_21342_13214# rowon_n[11] a_20946_13174# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2952 vcm a_2275_11190# a_9994_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2953 a_34394_12210# rowon_n[10] a_33998_12170# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2954 a_31990_10162# a_2275_10186# a_32082_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2955 a_9294_9198# rowon_n[7] a_8898_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2956 a_22954_12170# a_2275_12194# a_23046_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2957 a_24354_5182# col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2958 a_24050_6146# a_2475_6170# a_23958_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2959 a_21950_18194# a_2275_18218# a_22042_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2960 VDD rowon_n[9] a_20946_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2961 VDD rowon_n[8] a_33998_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2962 a_25966_8154# row_n[6] a_26458_8516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2963 VDD rowon_n[7] a_8898_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2964 VSS VDD a_10298_1166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2965 VSS row_n[15] a_32386_17230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2966 a_23958_3134# row_n[1] a_24450_3496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2967 a_20338_14218# col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2968 a_2475_16210# a_1957_16210# VDD VDD sky130_fd_pr__pfet_01v8 ad=3.42e+11p pd=2.97e+06u as=0p ps=0u w=1.2e+06u l=150000u
X2969 a_33390_13214# col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2970 a_12002_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2971 a_28370_7190# col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2972 a_29374_3174# col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2973 a_13006_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2974 a_27062_17190# a_2475_17214# a_26970_17190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2975 a_3270_16226# rowon_n[14] a_2874_16186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2976 a_13310_16226# rowon_n[14] a_12914_16186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2977 VSS row_n[11] a_10298_13214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2978 a_7286_6186# col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2979 a_29070_4138# a_2475_4162# a_28978_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2980 a_19334_9198# col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2981 a_27974_17190# row_n[15] a_28466_17552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2982 a_32482_15544# col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2983 vcm a_2275_13198# a_28066_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2984 a_32082_11166# a_2475_11190# a_31990_11166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2985 a_4882_15182# a_2275_15206# a_4974_15182# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2986 a_14922_15182# a_2275_15206# a_15014_15182# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2987 VSS row_n[7] a_20338_9198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2988 a_30378_9198# rowon_n[7] a_29982_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2989 VSS row_n[1] a_14314_3174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2990 a_32994_11166# row_n[9] a_33486_11528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2991 a_28978_1126# VDD a_29470_1488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2992 vcm a_2275_3158# a_32082_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2993 a_10394_11528# col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2994 a_34090_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2995 vcm a_2275_7174# a_31078_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2996 VDD rowon_n[4] a_17934_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2997 a_29982_6146# row_n[4] a_30474_6508# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2998 a_8898_12170# row_n[10] a_9390_12532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2999 a_18938_12170# row_n[10] a_19430_12532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3000 a_3970_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3001 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X3002 a_4974_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3003 a_17022_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3004 a_22954_2130# a_2275_2154# a_23046_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3005 VDD a_2161_4162# a_2275_4162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.42e+11p ps=2.97e+06u w=1.2e+06u l=150000u
X3006 a_2161_13198# sample VSS VSS sky130_fd_pr__nfet_01v8 ad=1.71e+11p pd=1.77e+06u as=0p ps=0u w=600000u l=150000u
X3007 a_18938_9158# row_n[7] a_19430_9520# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3008 a_33086_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3009 vcm a_2275_16210# a_30074_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3010 a_20434_9520# col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3011 a_12914_8154# a_2275_8178# a_13006_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3012 a_14410_1488# col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3013 a_13918_4138# a_2275_4162# a_14010_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3014 a_21438_5504# col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3015 VDD rowon_n[7] a_29982_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3016 a_33390_1166# col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3017 vcm a_2275_17214# a_16018_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3018 vcm a_2275_17214# a_5978_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3019 VSS row_n[13] a_28370_15222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3020 a_32386_13214# rowon_n[11] a_31990_13174# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3021 a_20034_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3022 a_8990_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3023 a_9994_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3024 a_29374_11206# col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3025 a_24050_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3026 a_20946_13174# a_2275_13198# a_21038_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3027 a_4882_7150# a_2275_7174# a_4974_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3028 a_5886_3134# a_2275_3158# a_5978_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3029 VDD rowon_n[15] a_26970_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3030 a_15014_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3031 a_33998_12170# a_2275_12194# a_34090_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3032 a_25454_7512# col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3033 a_17934_6146# a_2275_6170# a_18026_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3034 a_4974_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3035 VDD rowon_n[5] a_35002_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3036 a_8990_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3037 a_28466_13536# col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3038 VDD rowon_n[9] a_31990_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3039 VSS row_n[7] a_29374_9198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3040 a_10998_4138# a_2475_4162# a_10906_4138# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3041 a_23446_2492# col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3042 VSS VDD a_30378_18234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3043 VSS row_n[0] a_28370_2170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3044 a_31382_14218# col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3045 a_32386_8194# col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3046 VSS row_n[3] a_6282_5182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3047 a_1957_2154# VSS sample VDD sky130_fd_pr__pfet_01v8 ad=3.42e+11p pd=2.97e+06u as=0p ps=0u w=1.2e+06u l=150000u
X3048 a_25054_18194# a_2475_18218# a_24962_18194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3049 vcm a_2275_15206# a_22042_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3050 a_32082_9158# a_2475_9182# a_31990_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3051 VSS row_n[6] a_18330_8194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3052 a_16018_17190# a_2475_17214# a_15926_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3053 a_7286_15222# col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3054 a_17326_15222# col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3055 a_29470_9520# col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3056 a_25966_18194# VDD a_26458_18556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3057 a_5978_17190# a_2475_17214# a_5886_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3058 vcm a_2275_14202# a_26058_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3059 a_8386_8516# col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3060 a_2966_3134# a_2475_3158# a_2874_3134# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3061 a_20338_4178# rowon_n[2] a_19942_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3062 a_12914_16186# a_2275_16210# a_13006_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3063 a_30474_16548# col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3064 a_15014_6146# a_2475_6170# a_14922_6146# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3065 vcm a_2275_2154# a_21038_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3066 a_13310_2170# rowon_n[0] a_12914_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3067 a_24050_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3068 a_2874_16186# a_2275_16210# a_2966_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3069 a_9994_16186# a_2475_16210# a_9902_16186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3070 a_26970_7150# a_2275_7174# a_27062_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3071 a_31078_2130# a_2475_2154# a_30986_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3072 a_6378_17552# col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3073 a_16418_17552# col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3074 vcm a_2275_8178# a_10998_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3075 a_6378_3496# col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3076 vcm a_2275_4162# a_12002_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3077 a_16930_13174# row_n[11] a_17422_13536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3078 a_6890_13174# row_n[11] a_7382_13536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3079 VDD rowon_n[2] a_19942_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3080 vcm a_2275_12194# a_15014_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3081 vcm a_2275_12194# a_4974_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3082 a_24354_6186# rowon_n[4] a_23958_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3083 a_6982_5142# a_2475_5166# a_6890_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3084 a_7986_1126# a_2475_1150# a_7894_1126# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3085 VSS row_n[8] a_27366_10202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3086 vcm a_2275_18218# a_3970_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3087 vcm a_2275_18218# a_14010_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3088 a_27974_11166# a_2275_11190# a_28066_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3089 vcm a_2275_7174# a_2966_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3090 vcm a_2275_3158# a_3970_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3091 vcm a_2275_6170# a_16018_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3092 VSS row_n[14] a_26362_16226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3093 a_30378_14218# rowon_n[12] a_29982_14178# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3094 VDD rowon_n[10] a_25966_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3095 a_31990_1126# a_2275_1150# a_32082_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3096 a_30986_5142# a_2275_5166# a_31078_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3097 a_31078_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3098 a_35094_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3099 a_31990_13174# a_2275_13198# a_32082_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3100 a_5278_1166# col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3101 VSS row_n[2] a_19334_4178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3102 VDD VDD a_24962_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3103 a_2966_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3104 a_13006_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3105 a_28370_8194# rowon_n[6] a_27974_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3106 a_29374_4178# rowon_n[2] a_28978_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3107 a_25358_15222# col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3108 VDD rowon_n[6] a_14922_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3109 vcm a_2275_5166# a_7986_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3110 vcm a_2275_1150# a_8990_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3111 a_21342_7190# col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3112 a_22346_3174# col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3113 a_8290_17230# rowon_n[15] a_7894_17190# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3114 VDD a_2161_11190# a_2275_11190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.42e+11p ps=2.97e+06u w=1.2e+06u l=150000u
X3115 VSS row_n[5] a_31382_7190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3116 ctop sw_n ctop VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.9e+06u l=220000u
X3117 a_24450_17552# col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3118 a_20946_14178# row_n[12] a_21438_14540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3119 VSS row_n[11] a_9294_13214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3120 a_24050_13174# a_2475_13198# a_23958_13174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3121 a_6282_10202# col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3122 a_16322_10202# col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3123 vcm a_2275_10186# a_21038_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3124 a_12306_9198# col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3125 a_35002_7150# a_2275_7174# a_35094_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3126 a_22042_4138# a_2475_4162# a_21950_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3127 a_4974_12170# a_2475_12194# a_4882_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3128 a_15014_12170# a_2475_12194# a_14922_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3129 a_28066_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3130 a_17326_7190# rowon_n[5] a_16930_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3131 a_23958_6146# row_n[4] a_24450_6508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3132 VDD rowon_n[2] a_28978_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3133 a_19430_4500# col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3134 a_24962_13174# row_n[11] a_25454_13536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3135 a_8990_11166# a_2475_11190# a_8898_11166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3136 VDD rowon_n[5] a_6890_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3137 VDD rowon_n[13] a_7894_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3138 a_5374_12532# col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3139 a_15414_12532# col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3140 a_21950_1126# VDD a_22442_1488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3141 VDD rowon_n[0] a_4882_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3142 a_9390_11528# col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3143 a_2475_10186# a_1957_10186# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.71e+11p pd=1.77e+06u as=0p ps=0u w=600000u l=150000u
X3144 a_27366_1166# col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3145 a_26362_5182# col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3146 a_11910_9158# row_n[7] a_12402_9520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3147 a_4274_8194# col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3148 vcm a_2275_17214# a_35094_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3149 a_27974_8154# row_n[6] a_28466_8516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3150 a_12914_17190# row_n[15] a_13406_17552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3151 a_24354_15222# rowon_n[13] a_23958_15182# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3152 vcm a_2275_13198# a_13006_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3153 VSS row_n[10] a_21342_12210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3154 VSS VDD a_12306_1166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3155 a_2874_17190# row_n[15] a_3366_17552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3156 vcm a_2275_13198# a_2966_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3157 a_25966_3134# row_n[1] a_26458_3496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3158 a_28370_14218# rowon_n[12] a_27974_14178# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3159 VSS row_n[9] a_25358_11206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3160 a_2966_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3161 a_15014_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3162 a_29070_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3163 VDD rowon_n[12] a_19942_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3164 a_30074_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3165 a_15318_10202# rowon_n[8] a_14922_10162# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3166 a_14010_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3167 a_16930_7150# row_n[5] a_17422_7512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3168 a_9294_6186# col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3169 a_5278_10202# rowon_n[8] a_4882_10162# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3170 VDD rowon_n[11] a_23958_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3171 a_21438_10524# col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3172 a_10906_6146# a_2275_6170# a_10998_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3173 a_18330_3174# rowon_n[1] a_17934_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3174 VSS row_n[7] a_22346_9198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3175 a_30378_3174# col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3176 a_32386_9198# rowon_n[7] a_31990_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3177 a_23350_16226# col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3178 vcm a_2275_7174# a_33086_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3179 vcm a_2275_3158# a_34090_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3180 a_14922_10162# a_2275_10186# a_15014_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3181 a_26058_9158# a_2475_9182# a_25966_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3182 VSS row_n[0] a_21342_2170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3183 a_6982_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3184 a_4882_10162# a_2275_10186# a_4974_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3185 a_6282_18234# VDD a_5886_18194# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3186 a_16322_18234# VDD a_15926_18194# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3187 VSS row_n[13] a_3270_15222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3188 VSS row_n[13] a_13310_15222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3189 a_35094_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3190 a_3878_1126# a_2275_1150# a_3970_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3191 VDD en_bit_n[1] a_17934_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3192 a_29982_1126# VDD a_30474_1488# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3193 a_24962_2130# a_2275_2154# a_25054_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3194 a_22442_18556# col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3195 VSS row_n[12] a_17326_14218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3196 a_22042_14178# a_2475_14202# a_21950_14178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3197 a_14314_11206# col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3198 VSS row_n[6] a_11302_8194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3199 a_2874_5142# a_2275_5166# a_2966_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3200 a_35494_17552# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3201 VSS row_n[12] a_7286_14218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3202 a_31990_14178# row_n[12] a_32482_14540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3203 a_13006_13174# a_2475_13198# a_12914_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3204 a_35094_13174# a_2475_13198# a_35002_13174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3205 a_4274_11206# col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3206 vcm a_2275_10186# a_32082_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3207 a_22442_9520# col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3208 a_14922_8154# a_2275_8178# a_15014_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3209 a_35398_1166# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3210 a_15926_4138# a_2275_4162# a_16018_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3211 a_23446_5504# col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3212 a_17934_17190# a_2275_17214# a_18026_17190# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3213 a_2966_13174# a_2475_13198# a_2874_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3214 VDD rowon_n[7] a_31990_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3215 a_7894_17190# a_2275_17214# a_7986_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3216 VDD rowon_n[15] a_11910_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3217 VDD rowon_n[14] a_15926_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3218 a_13406_13536# col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3219 VDD rowon_n[14] a_5886_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3220 a_3366_13536# col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3221 VSS row_n[5] a_3270_7190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3222 vcm a_2275_18218# a_33086_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3223 VSS row_n[4] a_16322_6186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3224 a_7894_3134# a_2275_3158# a_7986_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3225 VSS row_n[10] a_19334_12210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3226 a_27462_7512# col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3227 a_24050_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3228 a_23350_10202# rowon_n[8] a_22954_10162# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3229 a_6378_6508# col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3230 a_13006_4138# a_2475_4162# a_12914_4138# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3231 a_15014_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3232 a_12002_8154# a_2475_8178# a_11910_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3233 a_25454_2492# col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3234 a_10906_18194# VDD a_11398_18556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3235 a_22346_16226# rowon_n[14] a_21950_16186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3236 a_35398_15222# rowon_n[13] a_35002_15182# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3237 vcm a_2275_14202# a_10998_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3238 a_4974_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3239 VDD rowon_n[0] a_35002_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3240 VDD rowon_n[12] a_17934_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3241 a_34394_8194# col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3242 a_27062_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3243 a_23958_15182# a_2275_15206# a_24050_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3244 a_19430_10524# col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3245 VSS row_n[3] a_8290_5182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3246 a_18026_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3247 a_34090_9158# a_2475_9182# a_33998_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3248 a_7986_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3249 a_27974_14178# a_2275_14202# a_28066_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3250 a_21342_8194# rowon_n[6] a_20946_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3251 a_4974_3134# a_2475_3158# a_4882_3134# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3252 a_22346_4178# rowon_n[2] a_21950_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3253 VDD rowon_n[11] a_35002_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3254 a_3970_7150# a_2475_7174# a_3878_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3255 vcm a_2275_2154# a_23046_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3256 a_10298_4178# col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3257 a_35398_10202# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3258 a_17022_6146# a_2475_6170# a_16930_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3259 a_33086_2130# a_2475_2154# a_32994_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3260 a_28978_7150# a_2275_7174# a_29070_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3261 a_8386_3496# col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3262 VSS row_n[8] a_12306_10202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3263 vcm a_2275_8178# a_13006_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3264 vcm a_2275_4162# a_14010_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3265 a_34394_16226# col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3266 a_2874_11166# a_2275_11190# a_2966_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3267 a_12914_11166# a_2275_11190# a_13006_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3268 VSS row_n[14] a_11302_16226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3269 a_34490_12532# col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3270 a_21038_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3271 a_10298_7190# rowon_n[5] a_9902_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3272 VDD rowon_n[2] a_21950_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3273 vcm a_2275_16210# a_29070_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3274 a_33086_14178# a_2475_14202# a_32994_14178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3275 VDD rowon_n[10] a_10906_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3276 a_26362_6186# rowon_n[4] a_25966_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3277 a_9994_1126# a_2475_1150# a_9902_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3278 a_9902_4138# row_n[2] a_10394_4500# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3279 a_33486_18556# col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3280 a_10998_14178# a_2475_14202# a_10906_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3281 a_8990_5142# a_2475_5166# a_8898_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3282 a_5886_18194# a_2275_18218# a_5978_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3283 VDD VDD a_9902_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3284 a_15926_18194# a_2275_18218# a_16018_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3285 a_4274_9198# rowon_n[7] a_3878_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3286 a_10298_15222# col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3287 vcm a_2275_7174# a_4974_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3288 vcm a_2275_3158# a_5978_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3289 vcm a_2275_6170# a_18026_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3290 a_2475_2154# a_1957_2154# VDD VDD sky130_fd_pr__pfet_01v8 ad=3.42e+11p pd=2.97e+06u as=0p ps=0u w=1.2e+06u l=150000u
X3291 a_15318_5182# rowon_n[3] a_14922_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3292 a_32994_5142# a_2275_5166# a_33086_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3293 a_20946_8154# row_n[6] a_21438_8516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3294 VDD rowon_n[7] a_3878_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3295 a_31478_8516# col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3296 VDD rowon_n[3] a_4882_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3297 a_9902_13174# row_n[11] a_10394_13536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3298 a_21342_11206# rowon_n[9] a_20946_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3299 VDD rowon_n[6] a_16930_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3300 a_35094_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3301 a_34394_10202# rowon_n[8] a_33998_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3302 a_2966_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3303 a_13006_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3304 a_23350_7190# col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3305 a_24354_3174# col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3306 VDD rowon_n[1] a_14922_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3307 VDD rowon_n[12] a_28978_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3308 a_17022_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3309 VSS row_n[5] a_33390_7190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3310 a_24050_4138# a_2475_4162# a_23958_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3311 a_6982_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3312 a_14314_9198# col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3313 vcm a_2275_7174# a_27062_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3314 a_21950_16186# a_2275_16210# a_22042_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3315 a_25966_6146# row_n[4] a_26458_6508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3316 a_5978_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3317 a_16018_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3318 VDD rowon_n[5] a_8898_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3319 a_28370_17230# col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3320 VSS row_n[13] a_32386_15222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3321 a_23958_1126# VDD a_24450_1488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3322 a_2475_14202# a_1957_14202# VDD VDD sky130_fd_pr__pfet_01v8 ad=3.42e+11p pd=2.97e+06u as=0p ps=0u w=1.2e+06u l=150000u
X3323 a_33390_11206# col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3324 VDD rowon_n[0] a_6890_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3325 a_13310_14218# rowon_n[12] a_12914_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3326 a_12002_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3327 a_29374_1166# col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3328 a_28370_5182# col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3329 VDD rowon_n[15] a_30986_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3330 a_27062_15182# a_2475_15206# a_26970_15182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3331 a_3270_14218# rowon_n[12] a_2874_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3332 a_9294_12210# col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3333 a_19334_12210# col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3334 vcm a_2275_12194# a_24050_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3335 VSS row_n[9] a_10298_11206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3336 a_13918_9158# row_n[7] a_14410_9520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3337 a_6282_8194# col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3338 a_7286_4178# col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3339 vcm a_2275_11190# a_28066_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3340 a_27974_15182# row_n[13] a_28466_15544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3341 a_32482_13536# col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3342 a_4882_13174# a_2275_13198# a_4974_13174# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3343 a_14922_13174# a_2275_13198# a_15014_13174# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3344 VSS VDD a_14314_1166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3345 a_8386_14540# col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3346 a_18426_14540# col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3347 vcm a_2275_1150# a_32082_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3348 a_27974_3134# row_n[1] a_28466_3496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3349 vcm a_2275_5166# a_31078_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3350 a_8898_10162# row_n[8] a_9390_10524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3351 a_18938_10162# row_n[8] a_19430_10524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3352 a_3970_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3353 a_4974_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3354 a_6890_4138# row_n[2] a_7382_4500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3355 a_17022_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3356 a_18938_7150# row_n[5] a_19430_7512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3357 a_29982_18194# VDD a_30474_18556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3358 vcm a_2275_14202# a_30074_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3359 a_20434_7512# col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3360 a_12914_6146# a_2275_6170# a_13006_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3361 VDD rowon_n[5] a_29982_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3362 a_16930_2130# row_n[0] a_17422_2492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3363 a_27366_17230# rowon_n[15] a_26970_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3364 vcm a_2275_15206# a_16018_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3365 VSS row_n[7] a_24354_9198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3366 vcm a_2275_15206# a_5978_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3367 a_34394_9198# rowon_n[7] a_33998_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3368 VSS row_n[11] a_28370_13214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3369 a_32386_11206# rowon_n[9] a_31990_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3370 a_28066_9158# a_2475_9182# a_27974_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3371 vcm a_2275_7174# a_35094_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3372 a_20034_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3373 VSS row_n[0] a_23350_2170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3374 a_8990_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3375 a_24050_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3376 VSS row_n[6] a_13310_8194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3377 a_19030_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3378 a_4882_5142# a_2275_5166# a_4974_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3379 a_5886_1126# a_2275_1150# a_5978_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3380 VDD rowon_n[13] a_26970_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3381 a_15014_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3382 a_24450_9520# col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3383 a_17934_4138# a_2275_4162# a_18026_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3384 a_25454_5504# col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3385 a_4974_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3386 VDD rowon_n[7] a_33998_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3387 a_3366_8516# col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3388 VDD rowon_n[3] a_35002_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3389 a_28466_11528# col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3390 VSS a_2161_9182# a_2275_9182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.71e+11p ps=1.77e+06u w=600000u l=150000u
X3391 a_21950_7150# a_2275_7174# a_22042_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3392 a_26362_18234# col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3393 VSS row_n[14] a_30378_16226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3394 VSS row_n[15] a_6282_17230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3395 VSS row_n[15] a_16322_17230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3396 a_21038_17190# a_2475_17214# a_20946_17190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3397 VSS row_n[5] a_5278_7190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3398 a_32386_6186# col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3399 VSS row_n[1] a_6282_3174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3400 a_35002_18194# a_2275_18218# a_35094_18194# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X3401 a_25054_16186# a_2475_16210# a_24962_16186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3402 a_17326_13214# col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3403 vcm a_2275_13198# a_22042_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3404 VSS row_n[4] a_18330_6186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3405 a_21950_17190# row_n[15] a_22442_17552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3406 a_1957_16210# VDD sample VSS sky130_fd_pr__nfet_01v8 ad=1.71e+11p pd=1.77e+06u as=0p ps=0u w=600000u l=150000u
X3407 a_16018_15182# a_2475_15206# a_15926_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3408 a_7286_13214# col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3409 a_29470_7512# col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3410 a_25966_16186# row_n[14] a_26458_16548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3411 a_5978_15182# a_2475_15206# a_5886_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3412 a_8386_6508# col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3413 a_2966_1126# a_2475_1150# a_2874_1126# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3414 a_12914_14178# a_2275_14202# a_13006_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3415 a_14010_8154# a_2475_8178# a_13918_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3416 a_15014_4138# a_2475_4162# a_14922_4138# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3417 a_16418_15544# col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3418 a_2874_14178# a_2275_14202# a_2966_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3419 a_9994_14178# a_2475_14202# a_9902_14178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3420 a_27462_2492# col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3421 a_26970_5142# a_2275_5166# a_27062_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3422 VDD VDD a_8898_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3423 a_6378_15544# col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3424 vcm a_2275_6170# a_10998_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3425 a_6378_1488# col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3426 a_16930_11166# row_n[9] a_17422_11528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3427 a_6890_11166# row_n[9] a_7382_11528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3428 vcm a_2275_10186# a_15014_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3429 a_4882_14178# row_n[12] a_5374_14540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3430 a_14922_14178# row_n[12] a_15414_14540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3431 a_26362_12210# rowon_n[10] a_25966_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3432 vcm a_2275_10186# a_4974_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3433 a_23958_10162# a_2275_10186# a_24050_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3434 a_23350_8194# rowon_n[6] a_22954_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3435 a_6982_3134# a_2475_3158# a_6890_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3436 a_24354_4178# rowon_n[2] a_23958_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3437 VDD rowon_n[6] a_9902_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3438 vcm a_2275_2154# a_25054_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3439 a_25358_18234# VDD a_24962_18194# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3440 a_1957_17214# VSS sample VDD sky130_fd_pr__pfet_01v8 ad=3.42e+11p pd=2.97e+06u as=0p ps=0u w=1.2e+06u l=150000u
X3441 vcm a_2275_16210# a_3970_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3442 vcm a_2275_16210# a_14010_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3443 vcm a_2275_5166# a_2966_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3444 a_35094_2130# a_2475_2154# a_35002_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3445 vcm a_2275_1150# a_3970_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3446 vcm a_2275_8178# a_15014_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3447 vcm a_2275_4162# a_16018_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3448 VSS row_n[12] a_26362_14218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3449 a_26970_17190# a_2275_17214# a_27062_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3450 VDD rowon_n[8] a_25966_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3451 a_29982_7150# a_2275_7174# a_30074_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3452 a_30986_3134# a_2275_3158# a_31078_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3453 a_31078_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3454 a_23046_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3455 a_12306_7190# rowon_n[5] a_11910_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3456 VDD rowon_n[2] a_23958_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3457 VSS row_n[15] a_24354_17230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3458 a_35094_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3459 VDD rowon_n[14] a_24962_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3460 a_2966_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3461 a_13006_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3462 a_28370_6186# rowon_n[4] a_27974_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3463 a_25358_13214# col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3464 a_6282_9198# rowon_n[7] a_5886_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3465 VDD rowon_n[4] a_14922_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3466 vcm a_2275_3158# a_7986_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3467 a_19030_17190# a_2475_17214# a_18938_17190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3468 VSS row_n[10] a_15318_12210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3469 a_20034_12170# a_2475_12194# a_19942_12170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3470 a_22346_1166# col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3471 a_21342_5182# col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3472 a_8290_15222# rowon_n[13] a_7894_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3473 VSS row_n[10] a_5278_12210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3474 a_5278_2170# rowon_n[0] a_4882_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3475 VSS row_n[3] a_31382_5182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3476 a_24450_15544# col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3477 a_20946_12170# row_n[10] a_21438_12532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3478 VSS row_n[9] a_9294_11206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3479 a_24050_11166# a_2475_11190# a_23958_11166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3480 ctop sw_n ctop VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.9e+06u l=220000u
X3481 a_35002_5142# a_2275_5166# a_35094_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3482 a_4974_10162# a_2475_10186# a_4882_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3483 a_15014_10162# a_2475_10186# a_14922_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3484 a_22954_8154# row_n[6] a_23446_8516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3485 a_17326_5182# rowon_n[3] a_16930_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3486 VDD rowon_n[12] a_13918_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3487 a_24962_11166# row_n[9] a_25454_11528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3488 a_33486_8516# col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3489 VDD rowon_n[12] a_3878_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3490 VDD rowon_n[7] a_5886_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3491 VDD rowon_n[3] a_6890_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3492 VDD rowon_n[11] a_7894_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3493 a_5374_10524# col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3494 a_15414_10524# col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3495 a_20946_3134# row_n[1] a_21438_3496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3496 a_13310_17230# col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3497 a_31478_3496# col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3498 a_3270_17230# col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3499 a_26362_3174# col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3500 VDD rowon_n[1] a_16930_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3501 a_11910_7150# row_n[5] a_12402_7512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3502 a_25358_7190# col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3503 VSS row_n[5] a_35398_7190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3504 a_4274_6186# col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3505 vcm a_2275_15206# a_35094_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3506 a_16322_9198# col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3507 vcm a_2275_7174# a_29070_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3508 a_27974_6146# row_n[4] a_28466_6508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3509 a_12914_15182# row_n[13] a_13406_15544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3510 a_24354_13214# rowon_n[11] a_23958_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3511 vcm a_2275_11190# a_13006_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3512 VSS row_n[8] a_21342_10202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3513 a_2874_15182# row_n[13] a_3366_15544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3514 vcm a_2275_11190# a_2966_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3515 a_21950_11166# a_2275_11190# a_22042_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3516 a_25966_1126# VDD a_26458_1488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3517 a_21038_9158# a_2475_9182# a_20946_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3518 VDD rowon_n[0] a_8898_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3519 VDD rowon_n[15] a_18938_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3520 a_29070_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3521 VDD rowon_n[10] a_19942_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3522 a_25966_12170# a_2275_12194# a_26058_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3523 a_15926_9158# row_n[7] a_16418_9520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3524 a_14010_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3525 a_16930_5142# row_n[3] a_17422_5504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3526 a_30074_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3527 a_19942_2130# a_2275_2154# a_20034_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3528 a_9294_4178# col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3529 a_8290_8194# col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3530 VDD rowon_n[9] a_23958_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3531 a_9902_8154# a_2275_8178# a_9994_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3532 a_18330_1166# en_bit_n[1] a_17934_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3533 a_30378_1166# col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3534 a_10906_4138# a_2275_4162# a_10998_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3535 VSS VDD a_22346_18234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3536 VSS row_n[15] a_35398_17230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3537 a_23350_14218# col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3538 vcm a_2275_5166# a_33086_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3539 a_12306_17230# rowon_n[15] a_11910_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3540 a_6982_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3541 a_8898_4138# row_n[2] a_9390_4500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3542 a_6282_16226# rowon_n[14] a_5886_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3543 a_16322_16226# rowon_n[14] a_15926_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3544 VSS row_n[11] a_3270_13214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3545 VSS row_n[11] a_13310_13214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3546 a_31078_12170# a_2475_12194# a_30986_12170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3547 a_22442_16548# col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3548 VSS row_n[4] a_11302_6186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3549 a_2874_3134# a_2275_3158# a_2966_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3550 a_35494_15544# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3551 a_31990_12170# row_n[10] a_32482_12532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3552 a_13006_11166# a_2475_11190# a_12914_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3553 a_35094_11166# a_2475_11190# a_35002_11166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3554 a_22442_7512# col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3555 a_14922_6146# a_2275_6170# a_15014_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3556 a_7894_15182# a_2275_15206# a_7986_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3557 a_17934_15182# a_2275_15206# a_18026_15182# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3558 a_2966_11166# a_2475_11190# a_2874_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3559 VDD rowon_n[5] a_31990_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3560 a_18938_2130# row_n[0] a_19430_2492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3561 VDD rowon_n[13] a_11910_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3562 a_20434_2492# col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3563 a_13406_11528# col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3564 VDD rowon_n[0] a_29982_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3565 a_3366_11528# col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3566 a_11302_18234# col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3567 a_35398_2170# rowon_n[0] a_35002_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3568 VSS row_n[0] a_25358_2170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3569 VSS row_n[3] a_3270_5182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3570 vcm a_2275_16210# a_33086_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3571 a_20034_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3572 VSS row_n[6] a_15318_8194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3573 a_7894_1126# a_2275_1150# a_7986_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3574 VSS row_n[2] a_16322_4178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3575 VSS row_n[8] a_19334_10202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3576 a_27462_5504# col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3577 vcm a_2275_17214# a_19030_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3578 a_5374_8516# col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3579 a_5978_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3580 vcm a_2275_17214# a_8990_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3581 a_12002_6146# a_2475_6170# a_11910_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3582 a_10906_16186# row_n[14] a_11398_16548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3583 a_22346_14218# rowon_n[12] a_21950_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3584 a_35398_13214# rowon_n[11] a_35002_13174# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3585 a_23958_7150# a_2275_7174# a_24050_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3586 a_3366_3496# col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3587 a_23046_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3588 VDD rowon_n[10] a_17934_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3589 a_34394_6186# col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3590 a_16418_4500# col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3591 a_27062_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3592 a_23958_13174# a_2275_13198# a_24050_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3593 VSS row_n[5] a_7286_7190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3594 VSS row_n[1] a_8290_3174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3595 a_18026_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3596 a_1957_8178# VDD sample VSS sky130_fd_pr__nfet_01v8 ad=1.71e+11p pd=1.77e+06u as=0p ps=0u w=600000u l=150000u
X3597 a_7986_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3598 a_21342_6186# rowon_n[4] a_20946_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3599 a_4974_1126# a_2475_1150# a_4882_1126# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3600 a_2161_2154# sample VDD VDD sky130_fd_pr__pfet_01v8 ad=3.42e+11p pd=2.97e+06u as=0p ps=0u w=1.2e+06u l=150000u
X3601 VSS row_n[10] a_34394_12210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3602 VDD rowon_n[9] a_35002_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3603 a_3970_5142# a_2475_5166# a_3878_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3604 a_11302_12210# rowon_n[10] a_10906_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3605 a_1957_11190# VDD sample VSS sky130_fd_pr__nfet_01v8 ad=1.71e+11p pd=1.77e+06u as=0p ps=0u w=600000u l=150000u
X3606 a_17022_4138# a_2475_4162# a_16930_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3607 VSS VDD a_33390_18234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3608 a_8386_1488# col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3609 a_29470_2492# col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3610 a_28978_5142# a_2275_5166# a_29070_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3611 a_29070_12170# a_2475_12194# a_28978_12170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3612 a_6890_8154# a_2275_8178# a_6982_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3613 vcm a_2275_6170# a_13006_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3614 a_10298_18234# VDD a_9902_18194# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3615 VDD rowon_n[12] a_32994_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3616 a_34394_14218# col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3617 a_28066_18194# a_2475_18218# a_27974_18194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3618 VSS row_n[12] a_11302_14218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3619 a_34490_10524# col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3620 a_10298_5182# rowon_n[3] a_9902_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3621 a_28978_18194# VDD a_29470_18556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3622 a_11910_17190# a_2275_17214# a_12002_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3623 vcm a_2275_14202# a_29070_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3624 VDD rowon_n[8] a_10906_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3625 a_26362_4178# rowon_n[2] a_25966_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3626 a_15926_16186# a_2275_16210# a_16018_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3627 a_33486_16548# col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3628 VDD rowon_n[6] a_11910_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3629 a_8990_3134# a_2475_3158# a_8898_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3630 a_5886_16186# a_2275_16210# a_5978_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3631 VDD rowon_n[14] a_9902_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3632 a_19030_8154# a_2475_8178# a_18938_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3633 a_10298_13214# col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3634 vcm a_2275_5166# a_4974_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3635 vcm a_2275_1150# a_5978_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3636 VDD rowon_n[1] a_9902_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3637 vcm a_2275_4162# a_18026_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3638 a_25054_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3639 a_14314_7190# rowon_n[5] a_13918_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3640 vcm a_2275_7174# a_22042_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3641 a_32994_3134# a_2275_3158# a_33086_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3642 a_15318_3174# rowon_n[1] a_14922_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3643 vcm a_2275_12194# a_18026_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3644 a_20946_6146# row_n[4] a_21438_6508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3645 VDD rowon_n[2] a_25966_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3646 vcm a_2275_12194# a_7986_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3647 VDD rowon_n[5] a_3878_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3648 a_31478_6508# col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3649 a_9902_11166# row_n[9] a_10394_11528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3650 a_31078_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3651 VDD rowon_n[4] a_16930_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3652 vcm a_2275_18218# a_6982_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3653 vcm a_2275_18218# a_17022_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3654 a_8290_9198# rowon_n[7] a_7894_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3655 a_22042_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3656 VDD VSS a_14922_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3657 a_24354_1166# col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3658 a_23350_5182# col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3659 a_21038_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3660 VDD rowon_n[10] a_28978_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3661 a_7286_2170# rowon_n[0] a_6890_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3662 VSS row_n[3] a_33390_5182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3663 vcm a_2275_5166# a_27062_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3664 a_31382_17230# rowon_n[15] a_30986_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3665 a_21950_14178# a_2275_14202# a_22042_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3666 a_24962_8154# row_n[6] a_25454_8516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3667 a_5978_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3668 a_16018_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3669 VDD rowon_n[7] a_7894_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3670 a_35494_8516# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3671 VDD rowon_n[3] a_8898_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3672 a_28370_15222# col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3673 VSS row_n[11] a_32386_13214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3674 a_19942_17190# a_2275_17214# a_20034_17190# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X3675 a_33486_3496# col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3676 a_22954_3134# row_n[1] a_23446_3496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3677 a_28370_3174# col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3678 a_12002_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3679 a_27462_17552# col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3680 VDD rowon_n[13] a_30986_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3681 a_23958_14178# row_n[12] a_24450_14540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3682 a_27062_13174# a_2475_13198# a_26970_13174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3683 a_9294_10202# col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3684 a_19334_10202# col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3685 vcm a_2275_10186# a_24050_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3686 a_13918_7150# row_n[5] a_14410_7512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3687 a_6282_6186# col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3688 a_7986_12170# a_2475_12194# a_7894_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3689 a_10906_12170# a_2275_12194# a_10998_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3690 a_18026_12170# a_2475_12194# a_17934_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3691 a_18330_9198# col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3692 a_27974_13174# row_n[11] a_28466_13536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3693 a_32482_11528# col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3694 a_11910_2130# row_n[0] a_12402_2492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3695 a_30378_18234# col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3696 a_8386_12532# col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3697 a_18426_12532# col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3698 a_17326_2170# col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3699 a_23046_9158# a_2475_9182# a_22954_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3700 vcm a_2275_7174# a_30074_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3701 a_27974_1126# VDD a_28466_1488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3702 vcm a_2275_3158# a_31078_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3703 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X3704 a_3970_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3705 vcm a_2275_18218# a_25054_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3706 a_17934_9158# row_n[7] a_18426_9520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3707 a_18938_5142# row_n[3] a_19430_5504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3708 a_32082_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3709 a_29982_16186# row_n[14] a_30474_16548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3710 a_12914_4138# a_2275_4162# a_13006_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3711 a_20434_5504# col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3712 a_29070_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3713 VDD rowon_n[3] a_29982_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3714 a_15926_17190# row_n[15] a_16418_17552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3715 a_27366_15222# rowon_n[13] a_26970_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3716 vcm a_2275_13198# a_16018_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3717 a_5886_17190# row_n[15] a_6378_17552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3718 vcm a_2275_13198# a_5978_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3719 VSS row_n[9] a_28370_11206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3720 vcm a_2275_5166# a_35094_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3721 a_19030_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3722 a_20034_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3723 a_8990_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3724 a_10998_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3725 a_33086_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3726 VSS row_n[4] a_13310_6186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3727 a_19030_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3728 a_4882_3134# a_2275_3158# a_4974_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3729 VDD rowon_n[11] a_26970_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3730 a_24450_7512# col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3731 VDD rowon_n[5] a_33998_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3732 a_3366_6508# col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3733 a_22346_17230# col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3734 a_2161_12194# sample VDD VDD sky130_fd_pr__pfet_01v8 ad=3.42e+11p pd=2.97e+06u as=0p ps=0u w=1.2e+06u l=150000u
X3735 a_16018_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3736 VSS a_2161_7174# a_2275_7174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.71e+11p ps=1.77e+06u w=600000u l=150000u
X3737 a_22442_2492# col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3738 a_21950_5142# a_2275_5166# a_22042_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3739 a_26362_16226# col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3740 VSS row_n[12] a_30378_14218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3741 a_17934_10162# a_2275_10186# a_18026_10162# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3742 VDD rowon_n[0] a_31990_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3743 a_30986_17190# a_2275_17214# a_31078_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3744 a_7894_10162# a_2275_10186# a_7986_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3745 VSS row_n[0] a_27366_2170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3746 a_9294_18234# VDD a_8898_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3747 VSS row_n[13] a_6282_15222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3748 VSS row_n[13] a_16322_15222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3749 a_21038_15182# a_2475_15206# a_20946_15182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3750 a_19334_8194# rowon_n[6] a_18938_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3751 a_31382_8194# col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3752 VSS row_n[3] a_5278_5182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3753 VSS VDD a_6282_1166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3754 a_32386_4178# col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3755 a_35002_16186# a_2275_16210# a_35094_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3756 a_25054_14178# a_2475_14202# a_24962_14178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3757 a_17326_11206# col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3758 vcm a_2275_11190# a_22042_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3759 VSS row_n[2] a_18330_4178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3760 a_25454_18556# col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3761 a_21950_15182# row_n[13] a_22442_15544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3762 a_1957_14202# VDD sample VSS sky130_fd_pr__nfet_01v8 ad=1.71e+11p pd=1.77e+06u as=0p ps=0u w=600000u l=150000u
X3763 a_16018_13174# a_2475_13198# a_15926_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3764 a_7286_11206# col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3765 VSS row_n[6] a_17326_8194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3766 a_29470_5504# col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3767 a_5978_13174# a_2475_13198# a_5886_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3768 a_7382_8516# col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3769 VDD rowon_n[15] a_4882_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3770 VDD rowon_n[15] a_14922_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3771 a_7986_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3772 a_14010_6146# a_2475_6170# a_13918_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3773 vcm a_2275_2154# a_20034_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3774 a_16418_13536# col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3775 a_25966_7150# a_2275_7174# a_26058_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3776 a_30074_2130# a_2475_2154# a_29982_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3777 a_26970_3134# a_2275_3158# a_27062_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3778 VDD rowon_n[14] a_8898_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3779 a_6378_13536# col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3780 vcm a_2275_8178# a_9994_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3781 a_5374_3496# col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3782 a_31990_4138# row_n[2] a_32482_4500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3783 vcm a_2275_4162# a_10998_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3784 a_16930_9158# a_2275_9182# a_17022_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3785 a_18426_4500# col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3786 VSS row_n[5] a_9294_7190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3787 a_4882_12170# row_n[10] a_5374_12532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3788 a_14922_12170# row_n[10] a_15414_12532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3789 a_27062_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3790 a_26362_10202# rowon_n[8] a_25966_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3791 a_23350_6186# rowon_n[4] a_22954_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3792 a_6982_1126# a_2475_1150# a_6890_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3793 a_18026_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3794 VDD rowon_n[4] a_9902_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3795 a_3878_18194# VDD a_4370_18556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3796 a_13918_18194# VDD a_14410_18556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3797 a_25358_16226# rowon_n[14] a_24962_16186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3798 a_1957_15206# VSS sample VDD sky130_fd_pr__pfet_01v8 ad=3.42e+11p pd=2.97e+06u as=0p ps=0u w=1.2e+06u l=150000u
X3799 vcm a_2275_14202# a_3970_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3800 vcm a_2275_14202# a_14010_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3801 a_7986_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3802 vcm a_2275_3158# a_2966_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3803 a_8898_8154# a_2275_8178# a_8990_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3804 vcm a_2275_6170# a_15014_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3805 a_26970_15182# a_2275_15206# a_27062_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3806 a_31078_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3807 a_30986_1126# a_2275_1150# a_31078_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3808 a_29982_5142# a_2275_5166# a_30074_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3809 a_12306_5182# rowon_n[3] a_11910_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3810 VSS row_n[13] a_24354_15222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3811 a_21342_12210# col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3812 a_28370_4178# rowon_n[2] a_27974_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3813 a_25358_11206# col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3814 VDD rowon_n[6] a_13918_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3815 vcm a_2275_1150# a_7986_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3816 VDD rowon_n[15] a_22954_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3817 a_19030_15182# a_2475_15206# a_18938_15182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3818 a_20434_14540# col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3819 a_29982_12170# a_2275_12194# a_30074_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3820 VSS row_n[8] a_15318_10202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3821 a_20034_10162# a_2475_10186# a_19942_10162# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3822 a_21342_3174# col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3823 VDD rowon_n[1] a_11910_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3824 a_8290_13214# rowon_n[11] a_7894_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3825 a_5886_11166# a_2275_11190# a_5978_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3826 a_15926_11166# a_2275_11190# a_16018_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3827 VSS row_n[8] a_5278_10202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3828 a_20338_7190# col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3829 VSS row_n[5] a_30378_7190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3830 VSS row_n[1] a_31382_3174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3831 a_24450_13536# col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3832 a_20946_10162# row_n[8] a_21438_10524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3833 a_2475_8178# a_1957_8178# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.71e+11p pd=1.77e+06u as=0p ps=0u w=600000u l=150000u
X3834 a_5978_8154# a_2475_8178# a_5886_8154# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3835 a_35002_3134# a_2275_3158# a_35094_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3836 a_11302_9198# col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3837 a_27062_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3838 a_16322_7190# rowon_n[5] a_15926_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3839 vcm a_2275_7174# a_24050_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3840 a_22954_6146# row_n[4] a_23446_6508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3841 a_17326_3174# rowon_n[1] a_16930_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3842 VDD rowon_n[10] a_13918_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3843 a_33486_6508# col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3844 VDD rowon_n[2] a_27974_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3845 VDD rowon_n[10] a_3878_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3846 VDD rowon_n[5] a_5886_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3847 a_8898_18194# a_2275_18218# a_8990_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3848 a_18938_18194# a_2275_18218# a_19030_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3849 VDD rowon_n[9] a_7894_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3850 a_20946_1126# VDD a_21438_1488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3851 a_26058_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3852 a_13310_15222# col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3853 a_31478_1488# col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3854 VDD rowon_n[0] a_3878_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3855 a_12002_17190# a_2475_17214# a_11910_17190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3856 a_34090_17190# a_2475_17214# a_33998_17190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3857 a_3270_15222# col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3858 VDD VSS a_16930_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3859 a_26362_1166# col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3860 a_10906_9158# row_n[7] a_11398_9520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3861 a_11910_5142# row_n[3] a_12402_5504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3862 a_4274_4178# col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3863 VSS row_n[3] a_35398_5182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3864 a_25358_5182# col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3865 a_35002_17190# row_n[15] a_35494_17552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3866 vcm a_2275_13198# a_35094_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3867 a_3270_8194# col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3868 a_9294_2170# rowon_n[0] a_8898_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3869 a_12402_17552# col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3870 a_19334_17230# rowon_n[15] a_18938_17190# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3871 vcm a_2275_5166# a_29070_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3872 a_20338_12210# rowon_n[10] a_19942_12170# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3873 vcm a_2275_8178# a_6982_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3874 a_12914_13174# row_n[11] a_13406_13536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3875 a_24354_11206# rowon_n[9] a_23958_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3876 a_2874_13174# row_n[11] a_3366_13536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3877 a_24962_3134# row_n[1] a_25454_3496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3878 a_5978_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3879 a_16018_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3880 a_35494_3496# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3881 a_29070_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3882 a_3878_4138# row_n[2] a_4370_4500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3883 VDD rowon_n[13] a_18938_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3884 VDD rowon_n[8] a_19942_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3885 a_15926_7150# row_n[5] a_16418_7512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3886 a_14010_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3887 a_9994_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3888 a_8290_6186# col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3889 vcm a_2275_18218# a_9994_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3890 a_9902_6146# a_2275_6170# a_9994_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3891 a_13918_2130# row_n[0] a_14410_2492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3892 VSS row_n[14] a_22346_16226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3893 VSS row_n[13] a_35398_15222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3894 a_32386_12210# col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3895 a_31382_9198# rowon_n[7] a_30986_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3896 a_19334_2170# col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3897 vcm a_2275_3158# a_33086_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3898 a_12306_15222# rowon_n[13] a_11910_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3899 a_25054_9158# a_2475_9182# a_24962_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3900 a_30378_2170# rowon_n[0] a_29982_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3901 VSS row_n[0] a_20338_2170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3902 VDD VDD a_20946_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3903 VDD rowon_n[15] a_33998_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3904 a_6282_14218# rowon_n[12] a_5886_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3905 a_16322_14218# rowon_n[12] a_15926_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3906 a_31478_14540# col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3907 vcm a_2275_12194# a_27062_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3908 VSS row_n[9] a_3270_11206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3909 VSS row_n[9] a_13310_11206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3910 a_31078_10162# a_2475_10186# a_30986_10162# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3911 VSS row_n[6] a_10298_8194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3912 a_34090_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3913 a_2874_1126# a_2275_1150# a_2966_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3914 VSS row_n[2] a_11302_4178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3915 a_35494_13536# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3916 a_31990_10162# row_n[8] a_32482_10524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3917 a_14922_4138# a_2275_4162# a_15014_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3918 a_22442_5504# col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3919 a_7894_13174# a_2275_13198# a_7986_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3920 a_17934_13174# a_2275_13198# a_18026_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3921 VDD rowon_n[7] a_30986_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3922 VDD rowon_n[3] a_31990_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3923 VDD rowon_n[11] a_11910_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3924 a_11302_16226# col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3925 a_11398_4500# col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3926 a_32082_18194# a_2475_18218# a_31990_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3927 VSS row_n[1] a_3270_3174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3928 a_32994_18194# VDD a_33486_18556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3929 vcm a_2275_14202# a_33086_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3930 a_18330_12210# rowon_n[10] a_17934_12170# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3931 VSS row_n[4] a_15318_6186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3932 a_10394_18556# col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3933 vcm a_2275_15206# a_19030_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3934 a_5374_6508# col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3935 a_5978_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3936 a_12002_4138# a_2475_4162# a_11910_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3937 vcm a_2275_15206# a_8990_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3938 a_35398_11206# rowon_n[9] a_35002_11166# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3939 a_18026_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3940 VDD rowon_n[0] a_33998_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3941 a_3366_1488# col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3942 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X3943 a_24450_2492# col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3944 a_23958_5142# a_2275_5166# a_24050_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3945 a_23046_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3946 VDD rowon_n[8] a_17934_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3947 VSS row_n[0] a_29374_2170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3948 a_34394_4178# col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3949 a_27062_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3950 a_33390_8194# col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3951 VSS row_n[3] a_7286_5182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3952 VSS VDD a_8290_1166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3953 a_18026_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3954 a_7986_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3955 a_3970_3134# a_2475_3158# a_3878_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3956 a_21342_4178# rowon_n[2] a_20946_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3957 a_35002_11166# a_2275_11190# a_35094_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3958 VSS row_n[8] a_34394_10202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3959 a_9390_8516# col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3960 a_11302_10202# rowon_n[8] a_10906_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3961 a_9994_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3962 a_32082_2130# a_2475_2154# a_31990_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3963 a_29374_18234# col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3964 VSS row_n[14] a_33390_16226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3965 a_27974_7150# a_2275_7174# a_28066_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3966 a_28978_3134# a_2275_3158# a_29070_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3967 a_10298_16226# rowon_n[14] a_9902_16186# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3968 a_29470_14540# col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3969 VDD rowon_n[10] a_32994_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3970 a_29070_10162# a_2475_10186# a_28978_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3971 a_6890_6146# a_2275_6170# a_6982_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3972 a_7382_3496# col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3973 a_33998_4138# row_n[2] a_34490_4500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3974 vcm a_2275_4162# a_13006_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3975 a_18938_9158# a_2275_9182# a_19030_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3976 a_28066_16186# a_2475_16210# a_27974_16186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3977 a_20034_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3978 a_10298_3174# rowon_n[1] a_9902_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3979 VDD VDD a_31990_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3980 VDD rowon_n[2] a_20946_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3981 a_28978_16186# row_n[14] a_29470_16548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3982 a_11910_15182# a_2275_15206# a_12002_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3983 a_8990_1126# a_2475_1150# a_8898_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3984 VDD VSS VSS sky130_fd_pr__cap_var_lvt w=1.64e+07u l=1.6e+07u
X3985 a_15926_14178# a_2275_14202# a_16018_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3986 VDD rowon_n[4] a_11910_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3987 a_5886_14178# a_2275_14202# a_5978_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3988 a_3270_9198# rowon_n[7] a_2874_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3989 a_19030_6146# a_2475_6170# a_18938_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3990 a_10298_11206# col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3991 vcm a_2275_3158# a_4974_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3992 VDD VSS a_9902_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3993 a_16018_9158# a_2475_9182# a_15926_9158# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3994 a_14314_5182# rowon_n[3] a_13918_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3995 a_15318_1166# VSS a_14922_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3996 a_32994_1126# a_2275_1150# a_33086_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3997 vcm a_2275_5166# a_22042_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3998 vcm a_2275_10186# a_18026_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3999 a_19942_8154# row_n[6] a_20434_8516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4000 a_7894_14178# row_n[12] a_8386_14540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4001 a_17934_14178# row_n[12] a_18426_14540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4002 a_29374_12210# rowon_n[10] a_28978_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4003 vcm a_2275_10186# a_7986_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4004 a_26970_10162# a_2275_10186# a_27062_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4005 VDD rowon_n[7] a_2874_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4006 a_30474_8516# col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4007 VDD rowon_n[3] a_3878_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4008 VDD rowon_n[6] a_15926_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4009 vcm a_2275_16210# a_6982_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4010 vcm a_2275_16210# a_17022_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4011 a_23350_3174# col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4012 VDD rowon_n[1] a_13918_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4013 a_21038_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4014 VDD rowon_n[8] a_28978_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4015 a_25358_9198# rowon_n[7] a_24962_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4016 a_7986_8154# a_2475_8178# a_7894_8154# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4017 VSS row_n[5] a_32386_7190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4018 VSS row_n[1] a_33390_3174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4019 a_13310_9198# col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4020 vcm a_2275_3158# a_27062_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4021 VSS a_2161_17214# a_2275_17214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.71e+11p ps=1.77e+06u w=600000u l=150000u
X4022 VSS row_n[15] a_27366_17230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4023 a_31382_15222# rowon_n[13] a_30986_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4024 a_29070_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4025 vcm a_2275_7174# a_26058_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4026 a_24962_6146# row_n[4] a_25454_6508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4027 a_5978_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4028 a_16018_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4029 VDD rowon_n[5] a_7894_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4030 a_35494_6508# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4031 a_28370_13214# col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4032 VSS row_n[9] a_32386_11206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4033 vcm a_2275_9182# a_17022_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4034 a_12306_2170# col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4035 a_19942_15182# a_2275_15206# a_20034_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4036 a_22954_1126# VDD a_23446_1488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4037 a_33486_1488# col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4038 a_28066_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4039 a_14010_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4040 VSS row_n[10] a_18330_12210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4041 a_23046_12170# a_2475_12194# a_22954_12170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4042 a_31990_8154# a_2275_8178# a_32082_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4043 VDD rowon_n[0] a_5886_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4044 a_3970_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4045 VSS row_n[10] a_8290_12210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4046 VDD rowon_n[7] a_24962_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4047 a_28370_1166# col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4048 a_27462_15544# col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4049 VDD rowon_n[11] a_30986_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4050 a_23958_12170# row_n[10] a_24450_12532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4051 a_27062_11166# a_2475_11190# a_26970_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4052 a_12914_9158# row_n[7] a_13406_9520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4053 a_5278_8194# col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4054 a_13918_5142# row_n[3] a_14410_5504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4055 a_6282_4178# col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4056 a_7986_10162# a_2475_10186# a_7894_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4057 a_18026_10162# a_2475_10186# a_17934_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4058 VDD rowon_n[12] a_16930_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4059 a_27974_11166# row_n[9] a_28466_11528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4060 VDD rowon_n[12] a_6890_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4061 vcm a_2275_8178# a_8990_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4062 a_30378_16226# col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4063 a_8386_10524# col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4064 a_18426_10524# col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4065 vcm a_2275_1150# a_31078_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4066 VDD a_2161_18218# a_2275_18218# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.42e+11p ps=2.97e+06u w=1.2e+06u l=150000u
X4067 vcm a_2275_17214# a_21038_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4068 vcm a_2275_5166# a_30074_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4069 a_6282_17230# col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4070 a_16322_17230# col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4071 a_3970_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4072 vcm a_2275_16210# a_25054_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4073 a_5886_4138# row_n[2] a_6378_4500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4074 a_17934_7150# row_n[5] a_18426_7512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4075 ctop sw_n analog_in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.9e+06u l=220000u
X4076 a_8990_18194# a_2475_18218# a_8898_18194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4077 vcm a_2275_12194# a_12002_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4078 a_15926_2130# row_n[0] a_16418_2492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4079 a_15926_15182# row_n[13] a_16418_15544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4080 a_27366_13214# rowon_n[11] a_26970_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4081 vcm a_2275_11190# a_16018_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4082 a_9390_18556# col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4083 a_5886_15182# row_n[13] a_6378_15544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4084 vcm a_2275_11190# a_5978_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4085 a_10998_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4086 a_33390_9198# rowon_n[7] a_32994_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4087 a_27366_8194# col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4088 a_27062_9158# a_2475_9182# a_26970_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4089 vcm a_2275_3158# a_35094_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4090 VDD VSS VSS sky130_fd_pr__cap_var_lvt w=1.64e+07u l=1.6e+07u
X4091 a_19030_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4092 VSS row_n[0] a_22346_2170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4093 a_28978_12170# a_2275_12194# a_29070_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4094 a_32386_2170# rowon_n[0] a_31990_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4095 a_4882_1126# a_2275_1150# a_4974_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4096 a_19030_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4097 VSS row_n[2] a_13310_4178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4098 VDD rowon_n[9] a_26970_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4099 VSS row_n[6] a_12306_8194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4100 a_26058_2130# a_2475_2154# a_25966_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4101 a_24450_5504# col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4102 VDD rowon_n[7] a_32994_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4103 VDD rowon_n[3] a_33998_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4104 VSS VDD a_25358_18234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4105 a_22346_15222# col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4106 a_2966_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4107 a_26362_14218# col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4108 a_2161_10186# sample VDD VDD sky130_fd_pr__pfet_01v8 ad=3.42e+11p pd=2.97e+06u as=0p ps=0u w=1.2e+06u l=150000u
X4109 a_20946_7150# a_2275_7174# a_21038_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4110 VSS a_2161_5166# a_2275_5166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.71e+11p ps=1.77e+06u w=600000u l=150000u
X4111 a_21950_3134# a_2275_3158# a_22042_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4112 a_15318_17230# rowon_n[15] a_14922_17190# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4113 a_31078_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4114 a_34090_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4115 a_5278_17230# rowon_n[15] a_4882_17190# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4116 a_30986_15182# a_2275_15206# a_31078_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4117 a_11910_9158# a_2275_9182# a_12002_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4118 a_12002_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4119 a_21438_17552# col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4120 a_9294_16226# rowon_n[14] a_8898_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4121 VSS row_n[11] a_6282_13214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4122 VSS row_n[11] a_16322_13214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4123 a_21038_13174# a_2475_13198# a_20946_13174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4124 a_19334_6186# rowon_n[4] a_18938_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4125 a_31382_6186# col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4126 VSS row_n[1] a_5278_3174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4127 a_13406_4500# col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4128 a_25454_16548# col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4129 a_35002_14178# a_2275_14202# a_35094_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4130 a_21950_13174# row_n[11] a_22442_13536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4131 VSS row_n[5] a_4274_7190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4132 a_16018_11166# a_2475_11190# a_15926_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4133 VSS row_n[4] a_17326_6186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4134 a_5978_11166# a_2475_11190# a_5886_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4135 a_7382_6508# col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4136 VDD rowon_n[13] a_4882_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4137 VDD rowon_n[13] a_14922_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4138 a_7986_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4139 a_14010_4138# a_2475_4162# a_13918_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4140 a_5278_12210# col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4141 a_15318_12210# col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4142 vcm a_2275_12194# a_20034_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4143 a_16418_11528# col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4144 a_26970_1126# a_2275_1150# a_27062_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4145 a_25966_5142# a_2275_5166# a_26058_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4146 a_6378_11528# col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4147 a_3878_8154# a_2275_8178# a_3970_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4148 vcm a_2275_6170# a_9994_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4149 a_5374_1488# col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4150 a_14314_18234# col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4151 a_4274_18234# col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4152 vcm a_2275_17214# a_32082_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4153 a_35398_8194# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4154 a_4370_14540# col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4155 a_14410_14540# col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4156 VSS row_n[3] a_9294_5182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4157 a_14922_10162# row_n[8] a_15414_10524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4158 a_23046_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4159 a_4882_10162# row_n[8] a_5374_10524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4160 a_23350_4178# rowon_n[2] a_22954_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4161 a_2161_8178# sample VSS VSS sky130_fd_pr__nfet_01v8 ad=1.71e+11p pd=1.77e+06u as=0p ps=0u w=600000u l=150000u
X4162 VSS row_n[5] a_26362_7190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4163 a_3878_16186# row_n[14] a_4370_16548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4164 a_13918_16186# row_n[14] a_14410_16548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4165 a_25358_14218# rowon_n[12] a_24962_14178# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X4166 a_1957_13198# VSS sample VDD sky130_fd_pr__pfet_01v8 ad=3.42e+11p pd=2.97e+06u as=0p ps=0u w=1.2e+06u l=150000u
X4167 a_34090_2130# a_2475_2154# a_33998_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4168 vcm a_2275_1150# a_2966_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4169 a_8898_6146# a_2275_6170# a_8990_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4170 a_9390_3496# col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4171 vcm a_2275_4162# a_15014_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4172 a_26058_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4173 a_23350_17230# rowon_n[15] a_22954_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4174 a_26970_13174# a_2275_13198# a_27062_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4175 a_29982_3134# a_2275_3158# a_30074_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4176 a_22042_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4177 a_11302_7190# rowon_n[5] a_10906_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4178 a_12306_3174# rowon_n[1] a_11910_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4179 VSS row_n[11] a_24354_13214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4180 a_21342_10202# col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4181 VDD rowon_n[2] a_22954_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4182 a_14314_12210# rowon_n[10] a_13918_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4183 VDD rowon_n[4] a_13918_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4184 a_21038_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4185 a_4274_12210# rowon_n[10] a_3878_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4186 a_11910_10162# a_2275_10186# a_12002_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4187 a_19430_17552# col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4188 VDD VSS VSS sky130_fd_pr__cap_var_lvt w=1.64e+07u l=1.6e+07u
X4189 VDD rowon_n[13] a_22954_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4190 a_19030_13174# a_2475_13198# a_18938_13174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4191 a_20434_12532# col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4192 VDD VSS a_11910_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4193 a_21342_1166# col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4194 a_8290_11206# rowon_n[9] a_7894_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4195 VSS VDD a_31382_1166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4196 VSS row_n[3] a_30378_5182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4197 a_20338_5182# col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4198 a_24450_11528# col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4199 a_5978_6146# a_2475_6170# a_5886_6146# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4200 a_35002_1126# a_2275_1150# a_35094_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4201 a_4274_2170# rowon_n[0] a_3878_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4202 a_18026_9158# a_2475_9182# a_17934_9158# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4203 a_16322_5182# rowon_n[3] a_15926_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4204 a_17326_1166# VSS a_16930_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4205 vcm a_2275_5166# a_24050_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4206 a_35398_17230# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4207 VDD rowon_n[8] a_13918_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4208 a_32482_8516# col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4209 VDD rowon_n[8] a_3878_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4210 VDD rowon_n[3] a_5886_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4211 VSS row_n[15] a_12306_17230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4212 a_8898_16186# a_2275_16210# a_8990_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4213 a_18938_16186# a_2275_16210# a_19030_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4214 a_19942_3134# row_n[1] a_20434_3496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4215 a_13310_13214# col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4216 a_30474_3496# col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4217 a_12002_15182# a_2475_15206# a_11910_15182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4218 a_34090_15182# a_2475_15206# a_33998_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4219 a_3270_13214# col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4220 vcm a_2275_12194# a_31078_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4221 a_25358_3174# col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4222 a_10906_7150# row_n[5] a_11398_7512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4223 VSS row_n[1] a_35398_3174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4224 VDD rowon_n[1] a_15926_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4225 a_35002_15182# row_n[13] a_35494_15544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4226 vcm a_2275_11190# a_35094_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4227 a_27366_9198# rowon_n[7] a_26970_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4228 a_9994_8154# a_2475_8178# a_9902_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4229 VSS row_n[5] a_34394_7190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4230 a_3270_6186# col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4231 a_12402_15544# col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4232 a_19334_15222# rowon_n[13] a_18938_15182# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X4233 a_20338_10202# rowon_n[8] a_19942_10162# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X4234 a_15318_9198# col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4235 vcm a_2275_7174# a_28066_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4236 vcm a_2275_3158# a_29070_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4237 a_21038_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4238 vcm a_2275_6170# a_6982_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4239 a_12914_11166# row_n[9] a_13406_11528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4240 vcm a_2275_9182# a_19030_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4241 VSS a_2161_12194# a_2275_12194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.71e+11p ps=1.77e+06u w=600000u l=150000u
X4242 a_2874_11166# row_n[9] a_3366_11528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4243 a_24962_1126# VDD a_25454_1488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4244 a_14314_2170# col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4245 a_25054_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4246 a_20034_9158# a_2475_9182# a_19942_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4247 a_33998_8154# a_2275_8178# a_34090_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4248 a_35494_1488# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4249 VDD rowon_n[0] a_7894_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4250 VDD rowon_n[11] a_18938_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4251 a_19942_10162# a_2275_10186# a_20034_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4252 a_14922_9158# row_n[7] a_15414_9520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4253 VDD rowon_n[7] a_26970_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4254 a_15926_5142# row_n[3] a_16418_5504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4255 a_8290_4178# col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4256 a_21342_18234# VDD a_20946_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4257 vcm a_2275_16210# a_9994_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4258 a_9902_4138# a_2275_4162# a_9994_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4259 a_34394_17230# rowon_n[15] a_33998_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4260 VSS row_n[12] a_22346_14218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4261 VSS row_n[11] a_35398_13214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4262 a_32386_10202# col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4263 a_22954_17190# a_2275_17214# a_23046_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4264 vcm a_2275_1150# a_33086_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4265 a_12306_13214# rowon_n[11] a_11910_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4266 a_7894_4138# row_n[2] a_8386_4500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4267 VDD rowon_n[14] a_20946_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4268 VDD rowon_n[13] a_33998_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4269 a_26970_14178# row_n[12] a_27462_14540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4270 a_31478_12532# col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4271 vcm a_2275_10186# a_27062_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4272 a_13918_12170# a_2275_12194# a_14010_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4273 VSS row_n[4] a_10298_6186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4274 a_3878_12170# a_2275_12194# a_3970_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4275 a_35494_11528# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4276 VDD rowon_n[5] a_30986_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4277 a_17934_2130# row_n[0] a_18426_2492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4278 a_33390_18234# col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4279 VDD rowon_n[9] a_11910_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4280 a_29374_8194# col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4281 VSS VDD a_10298_18234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4282 a_13006_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4283 a_29070_9158# a_2475_9182# a_28978_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4284 vcm a_2275_18218# a_28066_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4285 a_32082_16186# a_2475_16210# a_31990_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4286 a_11302_14218# col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4287 VSS row_n[0] a_24354_2170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4288 a_18330_10202# rowon_n[8] a_17934_10162# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X4289 a_34394_2170# rowon_n[0] a_33998_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4290 VSS VDD a_3270_1166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4291 a_32994_16186# row_n[14] a_33486_16548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4292 a_19030_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4293 VSS row_n[6] a_14314_8194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4294 a_28066_2130# a_2475_2154# a_27974_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4295 VSS row_n[2] a_15318_4178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4296 vcm a_2275_8178# a_32082_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4297 a_18938_17190# row_n[15] a_19430_17552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4298 a_10394_16548# col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4299 vcm a_2275_13198# a_19030_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4300 a_4370_8516# col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4301 a_5978_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4302 a_8898_17190# row_n[15] a_9390_17552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4303 vcm a_2275_13198# a_8990_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4304 a_4974_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4305 a_23958_3134# a_2275_3158# a_24050_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4306 VDD a_2161_9182# a_2275_9182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.42e+11p ps=2.97e+06u w=1.2e+06u l=150000u
X4307 a_22954_7150# a_2275_7174# a_23046_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4308 a_23046_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4309 a_33086_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4310 a_13918_9158# a_2275_9182# a_14010_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4311 a_33390_6186# col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4312 VSS row_n[1] a_7286_3174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4313 a_15414_4500# col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4314 a_33390_12210# rowon_n[10] a_32994_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4315 a_30986_10162# a_2275_10186# a_31078_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4316 a_3970_1126# a_2475_1150# a_3878_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4317 a_32386_18234# VDD a_31990_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4318 a_9390_6508# col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4319 a_9994_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4320 a_28978_1126# a_2275_1150# a_29070_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4321 a_29374_16226# col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4322 VSS row_n[12] a_33390_14218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4323 a_27974_5142# a_2275_5166# a_28066_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4324 a_20946_18194# a_2275_18218# a_21038_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4325 a_33998_17190# a_2275_17214# a_34090_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4326 a_10298_14218# rowon_n[12] a_9902_14178# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X4327 a_29470_12532# col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4328 VDD rowon_n[8] a_32994_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4329 a_5886_8154# a_2275_8178# a_5978_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4330 a_7382_1488# col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4331 a_6890_4138# a_2275_4162# a_6982_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4332 a_26458_8516# col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4333 a_28066_14178# a_2475_14202# a_27974_14178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4334 a_10998_9158# a_2475_9182# a_10906_9158# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4335 a_10298_1166# VSS a_9902_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4336 a_28466_18556# col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4337 VDD rowon_n[14] a_31990_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4338 a_11910_13174# a_2275_13198# a_12002_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4339 VDD rowon_n[6] a_10906_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4340 VSS row_n[5] a_28370_7190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4341 a_19030_4138# a_2475_4162# a_18938_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4342 a_1957_7174# VSS sample VDD sky130_fd_pr__pfet_01v8 ad=3.42e+11p pd=2.97e+06u as=0p ps=0u w=1.2e+06u l=150000u
X4343 vcm a_2275_1150# a_4974_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4344 a_20338_9198# rowon_n[7] a_19942_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4345 a_2966_8154# a_2475_8178# a_2874_8154# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4346 a_13310_7190# rowon_n[5] a_12914_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4347 vcm a_2275_3158# a_22042_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4348 a_14314_3174# rowon_n[1] a_13918_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4349 a_24050_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4350 vcm a_2275_7174# a_21038_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4351 a_31078_7150# a_2475_7174# a_30986_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4352 a_19942_6146# row_n[4] a_20434_6508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4353 a_7894_12170# row_n[10] a_8386_12532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4354 a_17934_12170# row_n[10] a_18426_12532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4355 a_29374_10202# rowon_n[8] a_28978_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4356 VDD rowon_n[5] a_2874_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4357 a_30474_6508# col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4358 vcm a_2275_9182# a_12002_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4359 VDD rowon_n[4] a_15926_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4360 a_16930_18194# VDD a_17422_18556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4361 vcm a_2275_14202# a_6982_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4362 vcm a_2275_14202# a_17022_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4363 a_23046_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4364 a_6890_18194# VDD a_7382_18556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4365 VDD rowon_n[7] a_19942_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4366 VDD VSS a_13918_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4367 a_23350_1166# col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4368 vcm a_2275_17214# a_15014_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4369 a_21038_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4370 a_7986_6146# a_2475_6170# a_7894_6146# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4371 VSS VDD a_33390_1166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4372 a_6282_2170# rowon_n[0] a_5886_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4373 VSS row_n[3] a_32386_5182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4374 vcm a_2275_17214# a_4974_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4375 vcm a_2275_1150# a_27062_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4376 VSS a_2161_15206# a_2275_15206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.71e+11p ps=1.77e+06u w=600000u l=150000u
X4377 VSS row_n[13] a_27366_15222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4378 a_31382_13214# rowon_n[11] a_30986_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4379 a_24354_12210# col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4380 vcm a_2275_5166# a_26058_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4381 vcm a_2275_8178# a_3970_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4382 a_34490_8516# col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4383 VDD rowon_n[3] a_7894_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4384 a_28370_11206# col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4385 a_19942_13174# a_2275_13198# a_20034_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4386 VDD rowon_n[15] a_25966_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4387 a_14010_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4388 a_23446_14540# col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4389 a_32994_12170# a_2275_12194# a_33086_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4390 VSS row_n[8] a_18330_10202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4391 a_23046_10162# a_2475_10186# a_22954_10162# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4392 a_31990_6146# a_2275_6170# a_32082_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4393 a_32482_3496# col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4394 a_3970_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4395 a_8898_11166# a_2275_11190# a_8990_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4396 a_18938_11166# a_2275_11190# a_19030_11166# VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X4397 VSS row_n[8] a_8290_10202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4398 VDD rowon_n[5] a_24962_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4399 a_31990_18194# a_2275_18218# a_32082_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4400 a_27462_13536# col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4401 VDD rowon_n[9] a_30986_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4402 a_23958_10162# row_n[8] a_24450_10524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4403 VSS row_n[7] a_19334_9198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4404 a_12914_7150# row_n[5] a_13406_7512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4405 a_5278_6186# col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4406 a_29374_9198# rowon_n[7] a_28978_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4407 VDD rowon_n[10] a_16930_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4408 a_10906_2130# row_n[0] a_11398_2492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4409 VDD rowon_n[10] a_6890_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4410 vcm a_2275_6170# a_8990_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4411 a_30378_14218# col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4412 a_22346_8194# col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4413 a_24050_18194# a_2475_18218# a_23958_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4414 VDD a_2161_16210# a_2275_16210# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.42e+11p ps=2.97e+06u w=1.2e+06u l=150000u
X4415 a_16322_15222# col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4416 vcm a_2275_15206# a_21038_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4417 a_22042_9158# a_2475_9182# a_21950_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4418 a_16322_2170# col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4419 vcm a_2275_3158# a_30074_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4420 VSS VDD a_9294_18234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4421 a_15014_17190# a_2475_17214# a_14922_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4422 a_6282_15222# col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4423 a_19430_9520# col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4424 a_24962_18194# VDD a_25454_18556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4425 a_4974_17190# a_2475_17214# a_4882_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4426 vcm a_2275_14202# a_25054_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4427 VDD rowon_n[7] a_28978_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4428 a_17934_5142# row_n[3] a_18426_5504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4429 a_15414_17552# col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4430 a_8990_16186# a_2475_16210# a_8898_16186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4431 vcm a_2275_10186# a_12002_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4432 a_21038_2130# a_2475_2154# a_20946_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4433 a_5374_17552# col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4434 a_11910_14178# row_n[12] a_12402_14540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4435 a_15926_13174# row_n[11] a_16418_13536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4436 a_27366_11206# rowon_n[9] a_26970_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4437 a_9390_16548# col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4438 a_5886_13174# row_n[11] a_6378_13536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4439 a_27366_6186# col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4440 vcm a_2275_1150# a_35094_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4441 a_19030_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4442 vcm a_2275_18218# a_2966_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4443 vcm a_2275_18218# a_13006_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4444 VSS row_n[15] a_21342_17230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4445 VSS row_n[4] a_12306_6186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4446 VDD rowon_n[5] a_32994_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4447 VSS row_n[14] a_25358_16226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4448 a_22346_13214# col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4449 a_2966_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4450 a_15014_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4451 a_21950_1126# a_2275_1150# a_22042_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4452 VSS a_2161_3158# a_2275_3158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.71e+11p ps=1.77e+06u w=600000u l=150000u
X4453 a_20946_5142# a_2275_5166# a_21038_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4454 a_30074_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4455 a_15318_15222# rowon_n[13] a_14922_15182# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4456 VDD rowon_n[0] a_30986_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4457 a_31078_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4458 a_34090_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4459 a_5278_15222# rowon_n[13] a_4882_15182# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4460 a_30986_13174# a_2275_13198# a_31078_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4461 VDD VDD a_23958_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4462 a_12002_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4463 a_21438_15544# col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4464 a_9294_14218# rowon_n[12] a_8898_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4465 VSS row_n[9] a_6282_11206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4466 VSS row_n[9] a_16322_11206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4467 a_21038_11166# a_2475_11190# a_20946_11166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4468 a_18330_8194# rowon_n[6] a_17934_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4469 a_30378_8194# col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4470 VSS VDD a_5278_1166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4471 a_31382_4178# col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4472 a_19334_4178# rowon_n[2] a_18938_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4473 a_21950_11166# row_n[9] a_22442_11528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4474 VSS row_n[3] a_4274_5182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4475 VSS row_n[2] a_17326_4178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4476 vcm a_2275_8178# a_34090_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4477 VDD rowon_n[11] a_4882_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4478 VDD rowon_n[11] a_14922_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4479 a_6982_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4480 VSS row_n[5] a_21342_7190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4481 a_7986_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4482 a_19942_14178# row_n[12] a_20434_14540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4483 a_5278_10202# col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4484 a_15318_10202# col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4485 vcm a_2275_10186# a_20034_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4486 a_24962_7150# a_2275_7174# a_25054_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4487 a_25966_3134# a_2275_3158# a_26058_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4488 a_3970_12170# a_2475_12194# a_3878_12170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4489 a_14010_12170# a_2475_12194# a_13918_12170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4490 a_35094_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4491 a_3878_6146# a_2275_6170# a_3970_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4492 a_4370_3496# col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4493 VDD rowon_n[2] a_18938_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4494 vcm a_2275_4162# a_9994_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4495 a_14314_16226# col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4496 a_15926_9158# a_2275_9182# a_16018_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4497 a_30986_4138# row_n[2] a_31478_4500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4498 a_13006_18194# a_2475_18218# a_12914_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4499 a_35094_18194# a_2475_18218# a_35002_18194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4500 a_4274_16226# col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4501 vcm a_2275_15206# a_32082_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4502 a_35398_6186# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4503 VSS row_n[1] a_9294_3174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4504 a_17422_4500# col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4505 a_2966_18194# a_2475_18218# a_2874_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4506 a_4370_12532# col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4507 a_14410_12532# col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4508 a_13406_18556# col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4509 a_3366_18556# col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4510 VSS row_n[3] a_26362_5182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4511 a_1957_11190# VSS sample VDD sky130_fd_pr__pfet_01v8 ad=3.42e+11p pd=2.97e+06u as=0p ps=0u w=1.2e+06u l=150000u
X4512 a_1957_1150# VDD sample VSS sky130_fd_pr__nfet_01v8 ad=1.71e+11p pd=1.77e+06u as=0p ps=0u w=600000u l=150000u
X4513 a_26058_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4514 a_7894_8154# a_2275_8178# a_7986_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4515 a_9390_1488# col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4516 a_8898_4138# a_2275_4162# a_8990_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4517 a_28466_8516# col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4518 VSS row_n[15] a_19334_17230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4519 a_23350_15222# rowon_n[13] a_22954_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4520 VSS row_n[10] a_20338_12210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4521 a_29982_1126# a_2275_1150# a_30074_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4522 a_13006_9158# a_2475_9182# a_12914_9158# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4523 a_11302_5182# rowon_n[3] a_10906_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4524 a_12306_1166# VSS a_11910_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4525 VSS row_n[9] a_24354_11206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4526 a_26458_3496# col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4527 a_14314_10202# rowon_n[8] a_13918_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4528 VDD rowon_n[6] a_12914_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4529 a_4274_10202# rowon_n[8] a_3878_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4530 a_19430_15544# col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4531 VDD rowon_n[11] a_22954_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4532 a_19030_11166# a_2475_11190# a_18938_11166# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4533 a_20434_10524# col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4534 a_20338_3174# col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4535 VSS row_n[1] a_30378_3174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4536 VDD rowon_n[1] a_10906_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4537 VDD VSS VSS sky130_fd_pr__cap_var_lvt w=1.64e+07u l=1.6e+07u
X4538 a_22346_9198# rowon_n[7] a_21950_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4539 a_4974_8154# a_2475_8178# a_4882_8154# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4540 a_5978_4138# a_2475_4162# a_5886_4138# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4541 VDD VDD a_35002_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4542 a_10298_9198# col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4543 vcm a_2275_7174# a_23046_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4544 vcm a_2275_3158# a_24050_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4545 a_16322_3174# rowon_n[1] a_15926_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4546 a_35398_15222# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4547 a_33086_7150# a_2475_7174# a_32994_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4548 a_32482_6508# col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4549 vcm a_2275_9182# a_14010_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4550 VSS row_n[13] a_12306_15222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4551 a_8898_14178# a_2275_14202# a_8990_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4552 a_18938_14178# a_2275_14202# a_19030_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4553 a_19942_1126# en_bit_n[0] a_20434_1488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4554 a_25054_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4555 a_13310_11206# col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4556 a_30474_1488# col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4557 a_34490_17552# col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4558 a_30986_14178# row_n[12] a_31478_14540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4559 a_12002_13174# a_2475_13198# a_11910_13174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4560 a_34090_13174# a_2475_13198# a_33998_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4561 a_3270_11206# col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4562 vcm a_2275_10186# a_31078_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4563 VDD VSS a_15926_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4564 a_25358_1166# col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4565 VDD rowon_n[0] a_2874_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4566 a_9902_9158# row_n[7] a_10394_9520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4567 VDD rowon_n[7] a_21950_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4568 a_10906_5142# row_n[3] a_11398_5504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4569 VSS VDD a_35398_1166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4570 VDD rowon_n[15] a_10906_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4571 a_35002_13174# row_n[11] a_35494_13536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4572 a_9994_6146# a_2475_6170# a_9902_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4573 a_8290_2170# rowon_n[0] a_7894_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4574 a_3270_4178# col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4575 VSS row_n[3] a_34394_5182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4576 a_12402_13536# col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4577 a_19334_13214# rowon_n[11] a_18938_13174# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X4578 vcm a_2275_1150# a_29070_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4579 vcm a_2275_5166# a_28066_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4580 vcm a_2275_8178# a_5978_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4581 vcm a_2275_4162# a_6982_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4582 a_2475_7174# a_1957_7174# VDD VDD sky130_fd_pr__pfet_01v8 ad=3.42e+11p pd=2.97e+06u as=0p ps=0u w=1.2e+06u l=150000u
X4583 VSS a_2161_10186# a_2275_10186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.71e+11p ps=1.77e+06u w=600000u l=150000u
X4584 a_33998_6146# a_2275_6170# a_34090_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4585 a_34490_3496# col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4586 a_2874_4138# row_n[2] a_3366_4500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4587 VDD rowon_n[9] a_18938_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4588 a_14922_7150# row_n[5] a_15414_7512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4589 VDD rowon_n[5] a_26970_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4590 a_2475_18218# a_1957_18218# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.71e+11p pd=1.77e+06u as=0p ps=0u w=600000u l=150000u
X4591 a_14010_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4592 a_9902_18194# VDD a_10394_18556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4593 a_21342_16226# rowon_n[14] a_20946_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4594 a_34394_15222# rowon_n[13] a_33998_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4595 vcm a_2275_14202# a_9994_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4596 VSS row_n[10] a_31382_12210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4597 a_3970_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4598 VDD rowon_n[0] a_24962_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4599 a_12914_2130# row_n[0] a_13406_2492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4600 VSS row_n[9] a_35398_11206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4601 a_24354_8194# col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4602 a_22954_15182# a_2275_15206# a_23046_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4603 a_18330_2170# col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4604 a_17022_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4605 VDD rowon_n[12] a_29982_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4606 a_26058_12170# a_2475_12194# a_25966_12170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4607 a_12306_11206# rowon_n[9] a_11910_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4608 a_24050_9158# a_2475_9182# a_23958_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4609 a_6982_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4610 VDD rowon_n[11] a_33998_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4611 a_26970_12170# row_n[10] a_27462_12532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4612 a_31478_10524# col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4613 a_23046_2130# a_2475_2154# a_22954_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4614 VSS row_n[2] a_10298_4178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4615 VDD rowon_n[3] a_30986_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4616 a_33390_16226# col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4617 a_29374_6186# col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4618 VSS row_n[14] a_10298_16226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4619 a_9294_17230# col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4620 a_19334_17230# col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4621 vcm a_2275_17214# a_24050_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4622 a_7286_9198# col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4623 vcm a_2275_16210# a_28066_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4624 a_32082_14178# a_2475_14202# a_31990_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4625 a_10394_4500# col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4626 a_14922_18194# a_2275_18218# a_15014_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4627 a_32482_18556# col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4628 a_4882_18194# a_2275_18218# a_4974_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4629 VSS row_n[4] a_14314_6186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4630 VDD VSS VSS sky130_fd_pr__cap_var_lvt w=1.64e+07u l=1.6e+07u
X4631 vcm a_2275_6170# a_32082_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4632 a_18938_15182# row_n[13] a_19430_15544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4633 vcm a_2275_11190# a_19030_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4634 a_4370_6508# col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4635 a_8898_15182# row_n[13] a_9390_15544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4636 vcm a_2275_11190# a_8990_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4637 a_6890_9158# row_n[7] a_7382_9520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4638 a_4974_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4639 a_23958_1126# a_2275_1150# a_24050_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4640 a_17022_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4641 a_33086_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4642 a_22954_5142# a_2275_5166# a_23046_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4643 VDD rowon_n[0] a_32994_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4644 a_21438_8516# col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4645 VSS row_n[10] a_29374_12210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4646 VSS VDD a_7286_1166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4647 a_16018_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4648 a_33390_4178# col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4649 a_34090_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4650 a_33390_10202# rowon_n[8] a_32994_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4651 a_12002_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4652 VSS VDD a_28370_18234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4653 a_32386_16226# rowon_n[14] a_31990_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4654 VDD rowon_n[12] a_27974_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4655 a_8990_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4656 VSS row_n[5] a_23350_7190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4657 a_9994_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4658 a_29374_14218# col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4659 a_27974_3134# a_2275_3158# a_28066_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4660 a_20946_16186# a_2275_16210# a_21038_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4661 a_33998_15182# a_2275_15206# a_34090_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4662 a_29470_10524# col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4663 a_5886_6146# a_2275_6170# a_5978_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4664 a_32994_4138# row_n[2] a_33486_4500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4665 a_4974_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4666 a_15014_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4667 a_17934_9158# a_2275_9182# a_18026_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4668 a_26458_6508# col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4669 a_28466_16548# col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4670 a_16930_2130# a_2275_2154# a_17022_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4671 VDD rowon_n[4] a_10906_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4672 a_8290_12210# col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4673 a_18330_12210# col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4674 vcm a_2275_12194# a_23046_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4675 VSS row_n[3] a_28370_5182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4676 VSS row_n[6] a_6282_8194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4677 a_1957_5166# VSS sample VDD sky130_fd_pr__pfet_01v8 ad=3.42e+11p pd=2.97e+06u as=0p ps=0u w=1.2e+06u l=150000u
X4678 a_17326_18234# col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4679 vcm a_2275_18218# a_22042_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4680 a_7286_18234# col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4681 a_2966_6146# a_2475_6170# a_2874_6146# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4682 a_7382_14540# col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4683 a_17422_14540# col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4684 a_13310_5182# rowon_n[3] a_12914_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4685 a_14314_1166# VSS a_13918_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4686 vcm a_2275_1150# a_22042_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4687 a_26058_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4688 a_15014_9158# a_2475_9182# a_14922_9158# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4689 a_28466_3496# col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4690 a_31078_5142# a_2475_5166# a_30986_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4691 vcm a_2275_5166# a_21038_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4692 a_7894_10162# row_n[8] a_8386_10524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4693 a_17934_10162# row_n[8] a_18426_10524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4694 VDD rowon_n[3] a_2874_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4695 a_16930_16186# row_n[14] a_17422_16548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4696 a_6890_16186# row_n[14] a_7382_16548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4697 VDD rowon_n[5] a_19942_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4698 VDD rowon_n[1] a_12914_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4699 a_26362_17230# rowon_n[15] a_25966_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4700 vcm a_2275_15206# a_15014_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4701 VSS row_n[1] a_32386_3174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4702 a_7986_4138# a_2475_4162# a_7894_4138# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4703 vcm a_2275_15206# a_4974_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4704 a_24354_9198# rowon_n[7] a_23958_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4705 a_6982_8154# a_2475_8178# a_6890_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4706 VSS row_n[11] a_27366_13214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4707 a_31382_11206# rowon_n[9] a_30986_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4708 a_24354_10202# col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4709 vcm a_2275_7174# a_25054_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4710 vcm a_2275_3158# a_26058_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4711 a_35094_7150# a_2475_7174# a_35002_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4712 vcm a_2275_6170# a_3970_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4713 a_34490_6508# col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4714 a_17326_12210# rowon_n[10] a_16930_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4715 vcm a_2275_9182# a_16018_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4716 a_2475_1150# a_1957_1150# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.71e+11p pd=1.77e+06u as=0p ps=0u w=600000u l=150000u
X4717 a_7286_12210# rowon_n[10] a_6890_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4718 a_27062_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4719 a_11302_2170# col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4720 VDD rowon_n[13] a_25966_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4721 a_14010_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4722 a_23446_12532# col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4723 a_30986_8154# a_2275_8178# a_31078_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4724 a_32482_1488# col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4725 a_31990_4138# a_2275_4162# a_32082_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4726 a_3970_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4727 VDD rowon_n[7] a_23958_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4728 VDD rowon_n[3] a_24962_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4729 a_31990_16186# a_2275_16210# a_32082_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4730 a_27462_11528# col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4731 a_12914_5142# row_n[3] a_13406_5504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4732 a_5278_4178# col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4733 a_25358_18234# col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4734 VDD rowon_n[8] a_16930_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4735 VDD rowon_n[8] a_6890_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4736 vcm a_2275_8178# a_7986_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4737 vcm a_2275_4162# a_8990_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4738 VSS row_n[15] a_5278_17230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4739 VSS row_n[15] a_15318_17230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4740 a_20034_17190# a_2475_17214# a_19942_17190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4741 a_22346_6186# col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4742 a_24050_16186# a_2475_16210# a_23958_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4743 VDD a_2161_14202# a_2275_14202# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.42e+11p ps=2.97e+06u w=1.2e+06u l=150000u
X4744 a_16322_13214# col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4745 vcm a_2275_13198# a_21038_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4746 a_5278_7190# rowon_n[5] a_4882_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4747 vcm a_2275_1150# a_30074_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4748 a_20946_17190# row_n[15] a_21438_17552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4749 VSS row_n[14] a_9294_16226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4750 a_15014_15182# a_2475_15206# a_14922_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4751 a_6282_13214# col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4752 vcm a_2275_12194# a_34090_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4753 a_19430_7512# col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4754 a_24962_16186# row_n[14] a_25454_16548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4755 a_4974_15182# a_2475_15206# a_4882_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4756 VDD rowon_n[5] a_28978_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4757 a_4882_4138# row_n[2] a_5374_4500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4758 a_15414_15544# col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4759 a_8990_14178# a_2475_14202# a_8898_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4760 a_11910_12170# row_n[10] a_12402_12532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4761 VDD VDD a_7894_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4762 a_5374_15544# col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4763 VDD rowon_n[0] a_26970_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4764 a_2475_13198# a_1957_13198# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.71e+11p pd=1.77e+06u as=0p ps=0u w=600000u l=150000u
X4765 a_15926_11166# row_n[9] a_16418_11528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4766 a_14922_2130# row_n[0] a_15414_2492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4767 a_5886_11166# row_n[9] a_6378_11528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4768 a_26362_8194# col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4769 a_27366_4178# col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4770 a_28066_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4771 a_22954_10162# a_2275_10186# a_23046_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4772 a_31382_2170# rowon_n[0] a_30986_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4773 VSS row_n[2] a_12306_4178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4774 a_24354_18234# VDD a_23958_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4775 vcm a_2275_16210# a_2966_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4776 vcm a_2275_16210# a_13006_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4777 VSS row_n[13] a_21342_15222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4778 a_25054_2130# a_2475_2154# a_24962_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4779 a_26970_4138# row_n[2] a_27462_4500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4780 VDD rowon_n[3] a_32994_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4781 VSS row_n[12] a_25358_14218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4782 a_22346_11206# col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4783 a_2966_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4784 a_25966_17190# a_2275_17214# a_26058_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4785 a_30074_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4786 a_19942_7150# a_2275_7174# a_20034_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4787 a_20946_3134# a_2275_3158# a_21038_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4788 VDD rowon_n[15] a_19942_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4789 a_15318_13214# rowon_n[11] a_14922_13174# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4790 a_9294_9198# col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4791 a_30074_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4792 a_31078_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4793 a_34090_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4794 a_5278_13214# rowon_n[11] a_4882_13174# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4795 a_10906_9158# a_2275_9182# a_10998_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4796 VDD rowon_n[14] a_23958_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4797 a_12002_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4798 a_21438_13536# col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4799 a_18330_6186# rowon_n[4] a_17934_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4800 a_30378_6186# col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4801 VSS row_n[1] a_4274_3174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4802 a_12402_4500# col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4803 a_16930_12170# a_2275_12194# a_17022_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4804 a_6890_12170# a_2275_12194# a_6982_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4805 VSS row_n[10] a_14314_12210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4806 vcm a_2275_6170# a_34090_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4807 VSS row_n[10] a_4274_12210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4808 VDD rowon_n[9] a_4882_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4809 VDD rowon_n[9] a_14922_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4810 a_6982_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4811 VSS row_n[3] a_21342_5182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4812 VSS VDD a_13310_18234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4813 a_19942_12170# row_n[10] a_20434_12532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4814 a_8898_9158# row_n[7] a_9390_9520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4815 a_25966_1126# a_2275_1150# a_26058_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4816 a_24962_5142# a_2275_5166# a_25054_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4817 VSS VDD a_3270_18234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4818 a_31078_17190# a_2475_17214# a_30986_17190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4819 a_3970_10162# a_2475_10186# a_3878_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4820 a_14010_10162# a_2475_10186# a_13918_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4821 a_2874_8154# a_2275_8178# a_2966_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4822 a_4370_1488# en_C0_n VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4823 a_3878_4138# a_2275_4162# a_3970_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4824 a_35094_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4825 VDD rowon_n[12] a_12914_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4826 a_14314_14218# col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4827 a_23446_8516# col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4828 a_31990_17190# row_n[15] a_32482_17552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4829 a_13006_16186# a_2475_16210# a_12914_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4830 a_35094_16186# a_2475_16210# a_35002_16186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4831 VDD rowon_n[12] a_2874_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4832 a_4274_14218# col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4833 vcm a_2275_13198# a_32082_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4834 VSS VDD a_9294_1166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4835 a_35398_4178# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4836 a_2966_16186# a_2475_16210# a_2874_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4837 a_4370_10524# col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4838 a_14410_10524# col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4839 a_18026_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4840 a_21438_3496# col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4841 a_13406_16548# col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4842 a_3366_16548# col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4843 VSS row_n[5] a_25358_7190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4844 VSS row_n[1] a_26362_3174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4845 a_35398_7190# rowon_n[5] a_35002_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4846 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X4847 a_26058_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4848 VSS row_n[7] a_16322_9198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4849 a_7894_6146# a_2275_6170# a_7986_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4850 a_28466_6508# col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4851 a_35002_4138# row_n[2] a_35494_4500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4852 VSS row_n[13] a_19334_15222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4853 a_23350_13214# rowon_n[11] a_22954_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4854 VSS row_n[8] a_20338_10202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4855 a_20946_11166# a_2275_11190# a_21038_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4856 a_11302_3174# rowon_n[1] a_10906_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4857 a_33998_10162# a_2275_10186# a_34090_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4858 a_26458_1488# col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4859 a_35398_18234# VDD a_35002_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4860 a_18938_2130# a_2275_2154# a_19030_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4861 VDD rowon_n[15] a_17934_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4862 a_24962_12170# a_2275_12194# a_25054_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4863 VDD rowon_n[4] a_12914_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4864 a_20034_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4865 a_16418_9520# col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4866 VSS row_n[6] a_8290_8194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4867 a_23958_18194# a_2275_18218# a_24050_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4868 a_19430_13536# col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4869 VDD rowon_n[9] a_22954_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4870 VDD VSS a_10906_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4871 a_20338_1166# en_bit_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4872 VSS VDD a_30378_1166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4873 VSS row_n[15] a_34394_17230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4874 a_2161_7174# sample VDD VDD sky130_fd_pr__pfet_01v8 ad=3.42e+11p pd=2.97e+06u as=0p ps=0u w=1.2e+06u l=150000u
X4875 a_4974_6146# a_2475_6170# a_4882_6146# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4876 a_3270_2170# rowon_n[0] a_2874_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4877 VDD rowon_n[14] a_35002_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4878 a_17022_9158# a_2475_9182# a_16930_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4879 a_16322_1166# VSS a_15926_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4880 vcm a_2275_1150# a_24050_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4881 vcm a_2275_5166# a_23046_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4882 a_11302_17230# rowon_n[15] a_10906_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4883 a_35398_13214# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4884 a_33086_5142# a_2475_5166# a_32994_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4885 a_29070_17190# a_2475_17214# a_28978_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4886 VSS row_n[11] a_12306_13214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4887 a_30074_12170# a_2475_12194# a_29982_12170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4888 a_16018_2130# a_2475_2154# a_15926_2130# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4889 a_34490_15544# col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4890 a_30986_12170# row_n[10] a_31478_12532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4891 a_12002_11166# a_2475_11190# a_11910_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4892 a_34090_11166# a_2475_11190# a_33998_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4893 a_9902_7150# row_n[5] a_10394_7512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4894 VDD rowon_n[5] a_21950_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4895 VSS row_n[1] a_34394_3174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4896 VDD rowon_n[13] a_10906_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4897 a_35002_11166# row_n[9] a_35494_11528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4898 a_26362_9198# rowon_n[7] a_25966_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4899 a_8990_8154# a_2475_8178# a_8898_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4900 a_9994_4138# a_2475_4162# a_9902_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4901 a_12402_11528# col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4902 a_19334_11206# rowon_n[9] a_18938_11166# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X4903 VDD rowon_n[0] a_19942_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4904 vcm a_2275_3158# a_28066_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4905 vcm a_2275_6170# a_5978_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4906 a_10298_18234# col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4907 vcm a_2275_9182# a_18026_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4908 a_2475_5166# a_1957_5166# VDD VDD sky130_fd_pr__pfet_01v8 ad=3.42e+11p pd=2.97e+06u as=0p ps=0u w=1.2e+06u l=150000u
X4909 a_25358_2170# rowon_n[0] a_24962_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4910 a_13310_2170# col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4911 a_32994_8154# a_2275_8178# a_33086_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4912 a_29070_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4913 a_33998_4138# a_2275_4162# a_34090_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4914 a_15318_8194# rowon_n[6] a_14922_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4915 vcm a_2275_17214# a_18026_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4916 VDD rowon_n[7] a_25966_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4917 a_14922_5142# row_n[3] a_15414_5504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4918 vcm a_2275_2154# a_17022_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4919 VDD rowon_n[3] a_26970_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4920 vcm a_2275_17214# a_7986_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4921 VDD rowon_n[6] a_4882_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4922 a_9902_16186# row_n[14] a_10394_16548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4923 a_21342_14218# rowon_n[12] a_20946_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4924 a_34394_13214# rowon_n[11] a_33998_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4925 a_27366_12210# col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4926 VSS row_n[8] a_31382_10202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4927 a_22042_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4928 a_31990_11166# a_2275_11190# a_32082_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4929 a_24354_6186# col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4930 a_22954_13174# a_2275_13198# a_23046_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4931 VDD rowon_n[15] a_28978_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4932 a_17022_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4933 a_26458_14540# col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4934 VDD rowon_n[10] a_29982_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4935 a_26058_10162# a_2475_10186# a_25966_10162# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4936 a_7286_7190# rowon_n[5] a_6890_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4937 a_6982_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4938 VDD rowon_n[9] a_33998_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4939 a_26970_10162# row_n[8] a_27462_10524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4940 VSS VDD a_32386_18234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4941 VDD rowon_n[0] a_28978_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4942 a_19430_2492# col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4943 a_33390_14218# col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4944 a_29374_4178# col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4945 a_27062_18194# a_2475_18218# a_26970_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4946 vcm a_2275_15206# a_24050_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4947 VSS row_n[12] a_10298_14218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4948 a_12002_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4949 a_28370_8194# col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4950 a_18026_17190# a_2475_17214# a_17934_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4951 a_9294_15222# col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4952 a_19334_15222# col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4953 a_27974_18194# VDD a_28466_18556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4954 a_7986_17190# a_2475_17214# a_7894_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4955 a_10906_17190# a_2275_17214# a_10998_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4956 vcm a_2275_14202# a_28066_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4957 a_14922_16186# a_2275_16210# a_15014_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4958 a_32482_16548# col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4959 a_33390_2170# rowon_n[0] a_32994_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4960 a_10998_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4961 a_4882_16186# a_2275_16210# a_4974_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4962 a_27062_2130# a_2475_2154# a_26970_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4963 VSS row_n[2] a_14314_4178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4964 a_8386_17552# col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4965 a_18426_17552# col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4966 vcm a_2275_8178# a_31078_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4967 a_17326_7190# col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4968 vcm a_2275_4162# a_32082_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4969 a_18938_13174# row_n[11] a_19430_13536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4970 a_28978_4138# row_n[2] a_29470_4500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4971 a_8898_13174# row_n[11] a_9390_13536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4972 a_3970_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4973 a_6890_7150# row_n[5] a_7382_7512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4974 a_4974_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4975 a_33086_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4976 a_22954_3134# a_2275_3158# a_23046_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4977 a_2161_16210# sample VSS VSS sky130_fd_pr__nfet_01v8 ad=1.71e+11p pd=1.77e+06u as=0p ps=0u w=600000u l=150000u
X4978 a_32082_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4979 a_12914_9158# a_2275_9182# a_13006_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4980 a_21438_6508# col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4981 a_30074_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4982 VSS row_n[8] a_29374_10202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4983 a_14410_4500# col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4984 vcm a_2275_18218# a_5978_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4985 vcm a_2275_18218# a_16018_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4986 a_11910_2130# a_2275_2154# a_12002_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4987 VSS row_n[14] a_28370_16226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4988 a_32386_14218# rowon_n[12] a_31990_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4989 a_20034_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4990 VDD rowon_n[10] a_27974_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4991 a_8990_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4992 VSS row_n[3] a_23350_5182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4993 a_10998_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4994 a_33086_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4995 a_27974_1126# a_2275_1150# a_28066_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4996 a_20946_14178# a_2275_14202# a_21038_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4997 a_33998_13174# a_2275_13198# a_34090_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4998 a_4882_8154# a_2275_8178# a_4974_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4999 a_5886_4138# a_2275_4162# a_5978_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5000 VDD VDD a_26970_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5001 a_4974_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5002 a_15014_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5003 a_25454_8516# col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5004 VDD rowon_n[6] a_35002_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5005 a_2161_17214# sample VDD VDD sky130_fd_pr__pfet_01v8 ad=3.42e+11p pd=2.97e+06u as=0p ps=0u w=1.2e+06u l=150000u
X5006 a_23446_3496# col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5007 a_22954_14178# row_n[12] a_23446_14540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5008 a_8290_10202# col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5009 a_18330_10202# col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5010 vcm a_2275_10186# a_23046_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5011 a_32386_9198# col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5012 VSS row_n[5] a_27366_7190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5013 VSS row_n[1] a_28370_3174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5014 a_6982_12170# a_2475_12194# a_6890_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5015 a_9902_12170# a_2275_12194# a_9994_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5016 a_17022_12170# a_2475_12194# a_16930_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5017 VSS row_n[4] a_6282_6186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5018 a_1957_3158# VSS sample VDD sky130_fd_pr__pfet_01v8 ad=3.42e+11p pd=2.97e+06u as=0p ps=0u w=1.2e+06u l=150000u
X5019 a_17326_16226# col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5020 vcm a_2275_16210# a_22042_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5021 VSS row_n[7] a_18330_9198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5022 a_16018_18194# a_2475_18218# a_15926_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5023 a_7286_16226# col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5024 a_2161_1150# sample VSS VSS sky130_fd_pr__nfet_01v8 ad=1.71e+11p pd=1.77e+06u as=0p ps=0u w=600000u l=150000u
X5025 a_2966_4138# a_2475_4162# a_2874_4138# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5026 a_5978_18194# a_2475_18218# a_5886_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5027 a_7382_12532# col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5028 a_17422_12532# col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5029 VDD VSS VSS sky130_fd_pr__cap_var_lvt w=1.64e+07u l=1.6e+07u
X5030 a_13310_3174# rowon_n[1] a_12914_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5031 vcm a_2275_7174# a_20034_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5032 a_28466_1488# col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5033 a_31078_3134# a_2475_3158# a_30986_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5034 vcm a_2275_3158# a_21038_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5035 a_16418_18556# col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5036 a_26970_8154# a_2275_8178# a_27062_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5037 a_30074_7150# a_2475_7174# a_29982_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5038 VDD VSS VSS sky130_fd_pr__cap_var_lvt w=1.64e+07u l=1.6e+07u
X5039 a_6378_18556# col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5040 vcm a_2275_9182# a_10998_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5041 a_31990_9158# row_n[7] a_32482_9520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5042 a_22042_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5043 a_18426_9520# col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5044 VDD VSS a_12914_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5045 VDD rowon_n[3] a_19942_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5046 a_14922_17190# row_n[15] a_15414_17552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5047 a_26362_15222# rowon_n[13] a_25966_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5048 vcm a_2275_13198# a_15014_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5049 VSS row_n[10] a_23350_12210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5050 VSS VDD a_32386_1166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5051 a_4882_17190# row_n[15] a_5374_17552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5052 vcm a_2275_13198# a_4974_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5053 a_6982_6146# a_2475_6170# a_6890_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5054 vcm a_2275_1150# a_26058_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5055 VSS row_n[9] a_27366_11206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5056 vcm a_2275_5166# a_25054_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5057 vcm a_2275_8178# a_2966_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5058 vcm a_2275_4162# a_3970_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5059 a_35094_5142# a_2475_5166# a_35002_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5060 VDD VSS VSS sky130_fd_pr__cap_var_lvt w=1.64e+07u l=1.6e+07u
X5061 VDD rowon_n[12] a_21950_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5062 a_32082_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5063 a_17326_10202# rowon_n[8] a_16930_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5064 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X5065 a_7286_10202# rowon_n[8] a_6890_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5066 a_18026_2130# a_2475_2154# a_17934_2130# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5067 a_31078_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5068 VDD rowon_n[11] a_25966_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5069 a_23446_10524# col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5070 a_30986_6146# a_2275_6170# a_31078_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5071 VDD rowon_n[5] a_23958_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5072 a_21342_17230# col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5073 a_31990_14178# a_2275_14202# a_32082_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5074 a_25358_16226# col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5075 a_28370_9198# rowon_n[7] a_27974_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5076 VDD rowon_n[0] a_21950_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5077 a_29982_17190# a_2275_17214# a_30074_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5078 vcm a_2275_6170# a_7986_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5079 a_9902_2130# row_n[0] a_10394_2492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5080 a_8290_18234# VDD a_7894_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5081 VSS row_n[13] a_5278_15222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5082 VSS row_n[13] a_15318_15222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5083 a_20034_15182# a_2475_15206# a_19942_15182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5084 a_12306_12210# col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5085 a_21342_8194# col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5086 a_27366_2170# rowon_n[0] a_26970_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5087 a_22346_4178# col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5088 a_24450_18556# col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5089 a_24050_14178# a_2475_14202# a_23958_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5090 a_16322_11206# col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5091 vcm a_2275_11190# a_21038_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5092 VSS row_n[6] a_31382_8194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5093 a_5278_5182# rowon_n[3] a_4882_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5094 a_15318_2170# col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5095 a_20946_15182# row_n[13] a_21438_15544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5096 VSS row_n[12] a_9294_14218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5097 a_33998_14178# row_n[12] a_34490_14540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5098 a_15014_13174# a_2475_13198# a_14922_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5099 a_6282_11206# col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5100 vcm a_2275_10186# a_34090_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5101 a_17326_8194# rowon_n[6] a_16930_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5102 a_35002_8154# a_2275_8178# a_35094_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5103 a_19430_5504# col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5104 a_4974_13174# a_2475_13198# a_4882_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5105 VDD rowon_n[7] a_27974_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5106 vcm a_2275_2154# a_19030_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5107 VDD rowon_n[3] a_28978_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5108 VDD rowon_n[15] a_3878_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5109 VDD rowon_n[15] a_13918_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5110 a_11398_14540# col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5111 VDD rowon_n[6] a_6890_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5112 a_15414_13536# col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5113 a_11910_10162# row_n[8] a_12402_10524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5114 a_20034_2130# a_2475_2154# a_19942_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5115 VDD rowon_n[14] a_7894_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5116 a_5374_13536# col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5117 a_26058_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5118 a_21950_4138# row_n[2] a_22442_4500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5119 VDD rowon_n[1] a_4882_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5120 a_26362_6186# col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5121 vcm a_2275_18218# a_35094_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5122 a_4274_9198# col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5123 a_9294_7190# rowon_n[5] a_8898_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5124 a_20338_17230# rowon_n[15] a_19942_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5125 a_17022_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5126 a_2874_18194# VDD a_3366_18556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5127 a_12914_18194# VDD a_13406_18556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5128 a_24354_16226# rowon_n[14] a_23958_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5129 vcm a_2275_14202# a_2966_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5130 vcm a_2275_14202# a_13006_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5131 VSS row_n[11] a_21342_13214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5132 a_6982_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5133 a_29070_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5134 a_25966_15182# a_2275_15206# a_26058_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5135 a_30074_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5136 a_3878_9158# row_n[7] a_4370_9520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5137 a_14010_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5138 a_20946_1126# a_2275_1150# a_21038_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5139 a_19942_5142# a_2275_5166# a_20034_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5140 VDD rowon_n[13] a_19942_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5141 a_5278_11206# rowon_n[9] a_4882_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5142 a_15318_11206# rowon_n[9] a_14922_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5143 a_16930_8154# row_n[6] a_17422_8516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5144 a_31078_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5145 a_30074_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5146 a_9994_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5147 a_20338_12210# col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5148 a_21438_11528# col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5149 VSS en_C0_n a_4274_1166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5150 a_30378_4178# col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5151 a_18330_4178# rowon_n[2] a_17934_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5152 a_13006_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5153 a_32386_17230# col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5154 a_29070_2130# a_2475_2154# a_28978_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5155 VSS row_n[8] a_14314_10202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5156 vcm a_2275_8178# a_33086_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5157 a_19334_7190# col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5158 vcm a_2275_4162# a_34090_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5159 a_4882_11166# a_2275_11190# a_4974_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5160 a_14922_11166# a_2275_11190# a_15014_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5161 VSS row_n[8] a_4274_10202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5162 VSS row_n[5] a_20338_7190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5163 VSS row_n[1] a_21342_3174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5164 a_6982_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5165 VSS row_n[14] a_13310_16226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5166 a_19942_10162# row_n[8] a_20434_10524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5167 a_8898_7150# row_n[5] a_9390_7512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5168 a_30378_7190# rowon_n[5] a_29982_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5169 a_24962_3134# a_2275_3158# a_25054_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5170 vcm a_2275_17214# a_27062_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5171 VSS row_n[14] a_3270_16226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5172 a_31078_15182# a_2475_15206# a_30986_15182# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5173 VSS row_n[7] a_11302_9198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5174 a_34090_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5175 a_2874_6146# a_2275_6170# a_2966_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5176 a_35094_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5177 VDD rowon_n[10] a_12914_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5178 a_23446_6508# col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5179 a_6890_2130# row_n[0] a_7382_2492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5180 a_29982_4138# row_n[2] a_30474_4500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5181 VDD rowon_n[2] a_17934_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5182 a_35494_18556# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5183 a_31990_15182# row_n[13] a_32482_15544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5184 a_13006_14178# a_2475_14202# a_12914_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5185 a_35094_14178# a_2475_14202# a_35002_14178# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5186 VDD rowon_n[10] a_2874_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5187 vcm a_2275_11190# a_32082_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5188 a_14922_9158# a_2275_9182# a_15014_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5189 a_7894_18194# a_2275_18218# a_7986_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5190 VDD VDD a_11910_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5191 a_17934_18194# a_2275_18218# a_18026_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5192 a_2966_14178# a_2475_14202# a_2874_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5193 a_2161_11190# sample VSS VSS sky130_fd_pr__nfet_01v8 ad=1.71e+11p pd=1.77e+06u as=0p ps=0u w=600000u l=150000u
X5194 VDD a_2161_2154# a_2275_2154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.42e+11p ps=2.97e+06u w=1.2e+06u l=150000u
X5195 a_21438_1488# col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5196 a_13918_2130# a_2275_2154# a_14010_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5197 VSS VDD a_26362_1166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5198 VSS row_n[3] a_25358_5182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5199 a_11398_9520# col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5200 VSS row_n[6] a_3270_8194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5201 a_35398_5182# rowon_n[3] a_35002_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5202 a_18330_17230# rowon_n[15] a_17934_17190# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X5203 a_7894_4138# a_2275_4162# a_7986_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5204 a_27462_8516# col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5205 VSS row_n[11] a_19334_13214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5206 a_23350_11206# rowon_n[9] a_22954_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5207 a_12002_9158# a_2475_9182# a_11910_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5208 a_11302_1166# VSS a_10906_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5209 a_4974_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5210 a_15014_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5211 a_25454_3496# col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5212 a_35398_16226# rowon_n[14] a_35002_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5213 VDD rowon_n[1] a_35002_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5214 VDD rowon_n[13] a_17934_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5215 a_10998_2130# a_2475_2154# a_10906_2130# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5216 a_8990_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5217 a_34394_9198# col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5218 a_16418_7512# col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5219 VSS row_n[5] a_29374_7190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5220 VSS row_n[4] a_8290_6186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5221 a_23958_16186# a_2275_16210# a_24050_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5222 a_19430_11528# col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5223 a_7986_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5224 a_18026_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5225 VSS row_n[13] a_34394_15222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5226 a_31382_12210# col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5227 a_21342_9198# rowon_n[7] a_20946_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5228 a_3970_8154# a_2475_8178# a_3878_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5229 a_2161_5166# sample VDD VDD sky130_fd_pr__pfet_01v8 ad=3.42e+11p pd=2.97e+06u as=0p ps=0u w=1.2e+06u l=150000u
X5230 a_4974_4138# a_2475_4162# a_4882_4138# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5231 vcm a_2275_3158# a_23046_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5232 a_11302_15222# rowon_n[13] a_10906_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5233 a_35398_11206# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5234 a_28978_8154# a_2275_8178# a_29070_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5235 a_32082_7150# a_2475_7174# a_31990_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5236 a_33086_3134# a_2475_3158# a_32994_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5237 vcm a_2275_9182# a_13006_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5238 a_20338_2170# rowon_n[0] a_19942_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5239 VDD rowon_n[15] a_32994_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5240 a_29070_15182# a_2475_15206# a_28978_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5241 a_30474_14540# col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5242 vcm a_2275_12194# a_26058_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5243 VSS row_n[9] a_12306_11206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5244 a_30074_10162# a_2475_10186# a_29982_10162# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5245 a_33998_9158# row_n[7] a_34490_9520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5246 a_24050_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5247 a_34490_13536# col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5248 a_30986_10162# row_n[8] a_31478_10524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5249 a_10298_8194# rowon_n[6] a_9902_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5250 VDD rowon_n[3] a_21950_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5251 VDD rowon_n[7] a_20946_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5252 a_9902_5142# row_n[3] a_10394_5504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5253 vcm a_2275_2154# a_12002_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5254 VDD rowon_n[11] a_10906_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5255 a_8990_6146# a_2475_6170# a_8898_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5256 vcm a_2275_1150# a_28066_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5257 vcm a_2275_8178# a_4974_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5258 vcm a_2275_4162# a_5978_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5259 a_10298_16226# col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5260 a_2475_3158# a_1957_3158# VDD VDD sky130_fd_pr__pfet_01v8 ad=3.42e+11p pd=2.97e+06u as=0p ps=0u w=1.2e+06u l=150000u
X5261 a_32994_6146# a_2275_6170# a_33086_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5262 a_15318_6186# rowon_n[4] a_14922_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5263 a_29374_17230# rowon_n[15] a_28978_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5264 vcm a_2275_15206# a_18026_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5265 VDD rowon_n[5] a_25966_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5266 vcm a_2275_15206# a_7986_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5267 a_30378_12210# rowon_n[10] a_29982_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5268 VDD rowon_n[4] a_4882_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5269 a_34394_11206# rowon_n[9] a_33998_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5270 a_27366_10202# col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5271 VDD rowon_n[0] a_23958_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5272 a_22042_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5273 VSS row_n[0] a_19334_2170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5274 a_24354_4178# col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5275 a_23350_8194# col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5276 VSS row_n[6] a_33390_8194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5277 a_29374_2170# rowon_n[0] a_28978_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5278 VDD rowon_n[13] a_28978_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5279 a_17022_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5280 a_26458_12532# col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5281 VDD rowon_n[8] a_29982_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5282 a_7286_5182# rowon_n[3] a_6890_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5283 a_6982_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5284 vcm a_2275_8178# a_27062_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5285 VDD rowon_n[6] a_8898_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5286 a_22042_2130# a_2475_2154# a_21950_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5287 a_28370_18234# col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5288 VSS row_n[14] a_32386_16226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5289 a_12306_7190# col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5290 a_28066_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5291 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X5292 VDD rowon_n[1] a_6890_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5293 a_23958_4138# row_n[2] a_24450_4500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5294 VSS row_n[15] a_8290_17230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5295 VSS row_n[15] a_18330_17230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5296 a_23046_17190# a_2475_17214# a_22954_17190# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5297 a_27062_16186# a_2475_16210# a_26970_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5298 vcm a_2275_13198# a_24050_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5299 a_28370_6186# col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5300 VDD VDD a_30986_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5301 a_23958_17190# row_n[15] a_24450_17552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5302 a_18026_15182# a_2475_15206# a_17934_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5303 a_9294_13214# col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5304 a_19334_13214# col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5305 a_6282_9198# col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5306 a_27974_16186# row_n[14] a_28466_16548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5307 a_7986_15182# a_2475_15206# a_7894_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5308 a_10906_15182# a_2275_15206# a_10998_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5309 a_14922_14178# a_2275_14202# a_15014_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5310 a_4882_14178# a_2275_14202# a_4974_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5311 a_8386_15544# col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5312 a_18426_15544# col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5313 vcm a_2275_6170# a_31078_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5314 a_17326_5182# col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5315 a_18938_11166# row_n[9] a_19430_11528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5316 a_8898_11166# row_n[9] a_9390_11528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5317 a_5886_9158# row_n[7] a_6378_9520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5318 a_3970_6146# a_2475_6170# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5319 a_6890_5142# row_n[3] a_7382_5504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5320 a_18938_8154# row_n[6] a_19430_8516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5321 a_22954_1126# a_2275_1150# a_23046_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5322 a_33086_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5323 a_2161_14202# sample VSS VSS sky130_fd_pr__nfet_01v8 ad=1.71e+11p pd=1.77e+06u as=0p ps=0u w=600000u l=150000u
X5324 a_32082_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5325 vcm a_2275_17214# a_12002_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5326 a_28370_12210# rowon_n[10] a_27974_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5327 a_25966_10162# a_2275_10186# a_26058_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5328 a_20434_8516# col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5329 VDD rowon_n[6] a_29982_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5330 a_15014_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5331 a_16930_3134# row_n[1] a_17422_3496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5332 a_27366_18234# VDD a_26970_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5333 vcm a_2275_16210# a_5978_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5334 vcm a_2275_16210# a_16018_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5335 vcm a_2275_8178# a_35094_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5336 VSS row_n[12] a_28370_14218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5337 a_28978_17190# a_2275_17214# a_29070_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5338 a_20034_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5339 VDD rowon_n[8] a_27974_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5340 VSS row_n[5] a_22346_7190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5341 VSS row_n[1] a_23350_3174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5342 a_8990_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5343 a_10998_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5344 a_33086_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5345 a_32386_7190# rowon_n[5] a_31990_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5346 VSS row_n[7] a_13310_9198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5347 a_19030_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5348 a_26058_7150# a_2475_7174# a_25966_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5349 a_4882_6146# a_2275_6170# a_4974_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5350 VDD rowon_n[14] a_26970_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5351 a_4974_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5352 a_15014_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5353 a_25454_6508# col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5354 a_8898_2130# row_n[0] a_9390_2492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5355 VDD rowon_n[4] a_35002_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5356 a_2161_15206# sample VDD VDD sky130_fd_pr__pfet_01v8 ad=3.42e+11p pd=2.97e+06u as=0p ps=0u w=1.2e+06u l=150000u
X5357 a_23446_1488# col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5358 VSS row_n[10] a_17326_12210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5359 a_22042_12170# a_2475_12194# a_21950_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5360 a_21950_8154# a_2275_8178# a_22042_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5361 a_15926_2130# a_2275_2154# a_16018_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5362 VSS row_n[10] a_7286_12210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5363 VSS VDD a_16322_18234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5364 a_21038_18194# a_2475_18218# a_20946_18194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5365 a_22954_12170# row_n[10] a_23446_12532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5366 VSS VDD a_28370_1166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5367 VSS row_n[3] a_27366_5182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5368 VSS VDD a_6282_18234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5369 a_6982_10162# a_2475_10186# a_6890_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5370 a_17022_10162# a_2475_10186# a_16930_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5371 a_13406_9520# col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5372 VSS row_n[6] a_5278_8194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5373 a_1957_1150# VSS sample VDD sky130_fd_pr__pfet_01v8 ad=3.42e+11p pd=2.97e+06u as=0p ps=0u w=1.2e+06u l=150000u
X5374 VSS row_n[2] a_6282_4178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5375 a_21950_18194# VDD a_22442_18556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5376 VDD rowon_n[12] a_15926_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5377 a_17326_14218# col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5378 vcm a_2275_14202# a_22042_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5379 a_1957_17214# VDD sample VSS sky130_fd_pr__nfet_01v8 ad=1.71e+11p pd=1.77e+06u as=0p ps=0u w=600000u l=150000u
X5380 a_16018_16186# a_2475_16210# a_15926_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5381 VDD rowon_n[12] a_5886_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5382 a_7286_14218# col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5383 a_29470_8516# col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5384 a_5978_16186# a_2475_16210# a_5886_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5385 a_7382_10524# col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5386 a_17422_10524# col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5387 a_13310_1166# VSS a_12914_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5388 vcm a_2275_1150# a_21038_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5389 a_15318_17230# col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5390 vcm a_2275_17214# a_20034_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5391 a_14010_9158# a_2475_9182# a_13918_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5392 a_31078_1126# a_2475_1150# a_30986_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5393 vcm a_2275_5166# a_20034_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5394 a_5278_17230# col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5395 a_16418_16548# col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5396 a_26970_6146# a_2275_6170# a_27062_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5397 a_27462_3496# col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5398 a_30074_5142# a_2475_5166# a_29982_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5399 a_6378_16548# col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5400 a_31990_7150# row_n[5] a_32482_7512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5401 a_6378_4500# col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5402 a_13006_2130# a_2475_2154# a_12914_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5403 vcm a_2275_12194# a_10998_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5404 a_18426_7512# col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5405 a_14922_15182# row_n[13] a_15414_15544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5406 a_26362_13214# rowon_n[11] a_25966_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5407 vcm a_2275_11190# a_15014_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5408 VSS row_n[8] a_23350_10202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5409 a_16418_2492# col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5410 a_4882_15182# row_n[13] a_5374_15544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5411 vcm a_2275_11190# a_4974_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5412 a_23958_11166# a_2275_11190# a_24050_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5413 a_23350_9198# rowon_n[7] a_22954_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5414 a_6982_4138# a_2475_4162# a_6890_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5415 a_35094_3134# a_2475_3158# a_35002_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5416 vcm a_2275_3158# a_25054_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5417 a_1957_18218# VSS sample VDD sky130_fd_pr__pfet_01v8 ad=3.42e+11p pd=2.97e+06u as=0p ps=0u w=1.2e+06u l=150000u
X5418 a_34090_7150# a_2475_7174# a_33998_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5419 vcm a_2275_6170# a_2966_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5420 VDD rowon_n[10] a_21950_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5421 a_27974_12170# a_2275_12194# a_28066_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5422 vcm a_2275_9182# a_15014_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5423 a_22346_2170# rowon_n[0] a_21950_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5424 a_10298_2170# col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5425 a_26970_18194# a_2275_18218# a_27062_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5426 a_31078_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5427 VDD rowon_n[9] a_25966_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5428 a_12306_8194# rowon_n[6] a_11910_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5429 a_29982_8154# a_2275_8178# a_30074_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5430 a_30986_4138# a_2275_4162# a_31078_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5431 VDD rowon_n[7] a_22954_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5432 vcm a_2275_2154# a_14010_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5433 VDD rowon_n[3] a_23958_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5434 VSS VDD a_24354_18234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5435 a_21342_15222# col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5436 a_25358_14218# col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5437 a_14314_17230# rowon_n[15] a_13918_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5438 a_21038_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5439 a_19030_18194# a_2475_18218# a_18938_18194# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5440 a_4274_17230# rowon_n[15] a_3878_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5441 a_29982_15182# a_2275_15206# a_30074_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5442 vcm a_2275_4162# a_7986_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5443 a_20434_17552# col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5444 a_8290_16226# rowon_n[14] a_7894_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5445 VSS row_n[11] a_5278_13214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5446 VSS row_n[11] a_15318_13214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5447 a_20034_13174# a_2475_13198# a_19942_13174# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5448 a_33086_12170# a_2475_12194# a_32994_12170# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5449 a_12306_10202# col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5450 a_21342_6186# col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5451 a_24450_16548# col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5452 a_20946_13174# row_n[11] a_21438_13536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5453 a_10998_12170# a_2475_12194# a_10906_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5454 a_4274_7190# rowon_n[5] a_3878_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5455 VSS row_n[4] a_31382_6186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5456 a_5278_3174# rowon_n[1] a_4882_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5457 a_33998_12170# row_n[10] a_34490_12532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5458 a_15014_11166# a_2475_11190# a_14922_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5459 a_17326_6186# rowon_n[4] a_16930_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5460 a_35002_6146# a_2275_6170# a_35094_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5461 a_4974_11166# a_2475_11190# a_4882_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5462 VDD rowon_n[5] a_27974_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5463 VDD rowon_n[13] a_3878_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5464 VDD rowon_n[13] a_13918_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5465 a_11398_12532# col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5466 VDD rowon_n[4] a_6890_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5467 a_15414_11528# col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5468 a_5374_11528# col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5469 VDD rowon_n[0] a_25966_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5470 a_26058_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5471 a_13310_18234# col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5472 VDD VSS a_4882_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5473 a_3270_18234# col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5474 vcm a_2275_17214# a_31078_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5475 a_25358_8194# col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5476 a_26362_4178# col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5477 vcm a_2275_16210# a_35094_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5478 a_11910_8154# row_n[6] a_12402_8516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5479 VSS row_n[6] a_35398_8194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5480 a_9294_5182# rowon_n[3] a_8898_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5481 a_22042_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5482 a_20338_15222# rowon_n[13] a_19942_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5483 vcm a_2275_8178# a_29070_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5484 a_2874_16186# row_n[14] a_3366_16548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5485 a_12914_16186# row_n[14] a_13406_16548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5486 a_24354_14218# rowon_n[12] a_23958_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5487 VSS row_n[9] a_21342_11206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5488 a_24050_2130# a_2475_2154# a_23958_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5489 a_25054_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5490 a_14314_7190# col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5491 VDD rowon_n[1] a_8898_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5492 a_25966_4138# row_n[2] a_26458_4500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5493 a_29070_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5494 a_25966_13174# a_2275_13198# a_26058_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5495 a_3878_7150# row_n[5] a_4370_7512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5496 a_19942_3134# a_2275_3158# a_20034_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5497 VDD VDD a_18938_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5498 VDD rowon_n[11] a_19942_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5499 a_8290_9198# col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5500 a_16930_6146# row_n[4] a_17422_6508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5501 a_30074_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5502 a_9994_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5503 a_20338_10202# col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5504 a_2475_12194# a_1957_12194# VDD VDD sky130_fd_pr__pfet_01v8 ad=3.42e+11p pd=2.97e+06u as=0p ps=0u w=1.2e+06u l=150000u
X5505 a_9902_9158# a_2275_9182# a_9994_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5506 a_13310_12210# rowon_n[10] a_12914_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5507 VSS VDD a_35398_18234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5508 a_32386_15222# col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5509 a_3270_12210# rowon_n[10] a_2874_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5510 a_10906_10162# a_2275_10186# a_10998_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5511 a_7286_2170# col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5512 vcm a_2275_6170# a_33086_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5513 a_19334_5182# col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5514 a_12306_18234# VDD a_11910_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5515 VSS VDD a_21342_1166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5516 VSS row_n[3] a_20338_5182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5517 VSS row_n[12] a_13310_14218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5518 a_7894_9158# row_n[7] a_8386_9520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5519 a_8898_5142# row_n[3] a_9390_5504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5520 a_24962_1126# a_2275_1150# a_25054_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5521 a_30378_5182# rowon_n[3] a_29982_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5522 a_31478_17552# col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5523 vcm a_2275_15206# a_27062_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5524 VSS row_n[12] a_3270_14218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5525 a_31078_13174# a_2475_13198# a_30986_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5526 a_35094_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5527 a_2874_4138# a_2275_4162# a_2966_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5528 a_34090_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5529 a_3878_17190# a_2275_17214# a_3970_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5530 a_13918_17190# a_2275_17214# a_14010_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5531 VDD rowon_n[8] a_12914_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5532 a_22442_8516# col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5533 a_35494_16548# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5534 a_31990_13174# row_n[11] a_32482_13536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5535 VDD rowon_n[8] a_2874_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5536 VDD rowon_n[6] a_31990_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5537 a_18938_3134# row_n[1] a_19430_3496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5538 a_7894_16186# a_2275_16210# a_7986_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5539 VDD rowon_n[14] a_11910_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5540 a_17934_16186# a_2275_16210# a_18026_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5541 a_17022_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5542 a_20434_3496# col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5543 vcm a_2275_12194# a_30074_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5544 VDD rowon_n[1] a_29982_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5545 VSS row_n[1] a_25358_3174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5546 a_11398_7512# col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5547 VSS row_n[5] a_24354_7190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5548 a_34394_7190# rowon_n[5] a_33998_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5549 VSS row_n[4] a_3270_6186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5550 a_35398_3174# rowon_n[1] a_35002_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5551 a_18330_15222# rowon_n[13] a_17934_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5552 a_20034_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5553 VSS row_n[7] a_15318_9198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5554 a_28066_7150# a_2475_7174# a_27974_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5555 a_27462_6508# col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5556 VSS row_n[9] a_19334_11206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5557 a_10998_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5558 a_33086_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5559 vcm a_2275_18218# a_19030_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5560 a_5978_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5561 vcm a_2275_18218# a_8990_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5562 a_24050_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5563 a_23958_8154# a_2275_8178# a_24050_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5564 a_25454_1488# col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5565 a_35398_14218# rowon_n[12] a_35002_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5566 VDD VSS a_35002_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5567 analog_in sw_n ctop VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.9e+06u l=220000u
X5568 a_17934_2130# a_2275_2154# a_18026_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5569 a_23046_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5570 VDD rowon_n[11] a_17934_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5571 VSS row_n[3] a_29374_5182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5572 a_15414_9520# col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5573 a_16418_5504# col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5574 VSS row_n[2] a_8290_4178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5575 a_33390_17230# rowon_n[15] a_32994_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5576 a_23958_14178# a_2275_14202# a_24050_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5577 VSS row_n[6] a_7286_8194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5578 a_7986_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5579 a_18026_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5580 VSS row_n[11] a_34394_13214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5581 a_31382_10202# col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5582 a_3970_6146# a_2475_6170# a_3878_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5583 a_2161_3158# sample VDD VDD sky130_fd_pr__pfet_01v8 ad=3.42e+11p pd=2.97e+06u as=0p ps=0u w=1.2e+06u l=150000u
X5584 vcm a_2275_1150# a_23046_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5585 a_11302_13214# rowon_n[11] a_10906_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5586 a_1957_12194# VDD sample VSS sky130_fd_pr__nfet_01v8 ad=1.71e+11p pd=1.77e+06u as=0p ps=0u w=600000u l=150000u
X5587 a_28978_6146# a_2275_6170# a_29070_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5588 a_33086_1126# a_2475_1150# a_32994_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5589 a_29470_3496# col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5590 a_32082_5142# a_2475_5166# a_31990_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5591 a_6890_9158# a_2275_9182# a_6982_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5592 a_29470_17552# col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5593 VDD rowon_n[13] a_32994_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5594 a_25966_14178# row_n[12] a_26458_14540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5595 a_29070_13174# a_2475_13198# a_28978_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5596 a_30474_12532# col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5597 vcm a_2275_10186# a_26058_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5598 a_33998_7150# row_n[5] a_34490_7512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5599 a_8386_4500# col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5600 a_9994_12170# a_2475_12194# a_9902_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5601 a_12914_12170# a_2275_12194# a_13006_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5602 a_15014_2130# a_2475_2154# a_14922_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5603 a_2874_12170# a_2275_12194# a_2966_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5604 a_34490_11528# col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5605 a_10298_6186# rowon_n[4] a_9902_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5606 a_31990_2130# row_n[0] a_32482_2492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5607 VDD VSS VSS sky130_fd_pr__cap_var_lvt w=1.64e+07u l=1.6e+07u
X5608 a_11910_18194# a_2275_18218# a_12002_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5609 VDD rowon_n[9] a_10906_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5610 VDD rowon_n[5] a_20946_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5611 a_18426_2492# col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5612 a_8990_4138# a_2475_4162# a_8898_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5613 a_19030_9158# a_2475_9182# a_18938_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5614 vcm a_2275_6170# a_4974_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5615 a_10298_14218# col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5616 a_2475_1150# a_1957_1150# VDD VDD sky130_fd_pr__pfet_01v8 ad=3.42e+11p pd=2.97e+06u as=0p ps=0u w=1.2e+06u l=150000u
X5617 a_24354_2170# rowon_n[0] a_23958_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5618 a_32994_4138# a_2275_4162# a_33086_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5619 a_14314_8194# rowon_n[6] a_13918_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5620 vcm a_2275_8178# a_22042_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5621 a_15318_4178# rowon_n[2] a_14922_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5622 a_17934_17190# row_n[15] a_18426_17552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5623 a_29374_15222# rowon_n[13] a_28978_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5624 vcm a_2275_13198# a_18026_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5625 VSS row_n[10] a_26362_12210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5626 vcm a_2275_2154# a_16018_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5627 VDD rowon_n[3] a_25966_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5628 a_7894_17190# row_n[15] a_8386_17552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5629 vcm a_2275_13198# a_7986_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5630 a_31078_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5631 a_30378_10202# rowon_n[8] a_29982_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5632 VDD rowon_n[6] a_3878_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5633 a_22042_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5634 a_23046_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5635 VDD rowon_n[12] a_24962_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5636 a_13006_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5637 a_35094_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5638 a_2966_12170# a_2475_12194# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5639 a_23350_6186# col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5640 VSS row_n[4] a_33390_6186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5641 VDD rowon_n[2] a_14922_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5642 VDD rowon_n[11] a_28978_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5643 a_26458_10524# col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5644 a_29982_10162# a_2275_10186# a_30074_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5645 a_6282_7190# rowon_n[5] a_5886_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5646 a_7286_3174# rowon_n[1] a_6890_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5647 vcm a_2275_6170# a_27062_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5648 a_31382_18234# VDD a_30986_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5649 a_24354_17230# col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5650 VDD rowon_n[4] a_8898_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5651 a_28370_16226# col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5652 VSS row_n[12] a_32386_14218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5653 a_12306_5182# col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5654 VDD rowon_n[0] a_27974_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5655 a_28066_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5656 a_19942_18194# a_2275_18218# a_20034_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5657 a_32994_17190# a_2275_17214# a_33086_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5658 VDD VSS a_6890_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5659 VSS row_n[13] a_8290_15222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5660 VSS row_n[13] a_18330_15222# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5661 a_23046_15182# a_2475_15206# a_22954_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5662 a_27062_14178# a_2475_14202# a_26970_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5663 a_19334_11206# col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5664 vcm a_2275_11190# a_24050_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5665 a_13918_8154# row_n[6] a_14410_8516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5666 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X5667 a_28370_4178# col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5668 a_27462_18556# col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5669 VDD rowon_n[14] a_30986_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5670 a_23958_15182# row_n[13] a_24450_15544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5671 a_18026_13174# a_2475_13198# a_17934_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5672 a_9294_11206# col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5673 a_7986_13174# a_2475_13198# a_7894_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5674 a_10906_13174# a_2275_13198# a_10998_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5675 VDD rowon_n[15] a_6890_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5676 VDD rowon_n[15] a_16930_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5677 a_11910_3134# row_n[1] a_12402_3496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5678 a_18426_13536# col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5679 a_8386_13536# col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5680 vcm a_2275_8178# a_30074_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5681 a_16322_7190# col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5682 a_17326_3174# col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5683 vcm a_2275_4162# a_31078_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5684 ctop sw ctop VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.9e+06u l=220000u
X5685 a_27974_4138# row_n[2] a_28466_4500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5686 a_5886_7150# row_n[5] a_6378_7512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5687 a_3970_4138# a_2475_4162# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5688 a_18938_6146# row_n[4] a_19430_6508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5689 a_21038_7150# a_2475_7174# a_20946_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5690 a_32082_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5691 vcm a_2275_15206# a_12002_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5692 a_29070_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5693 a_28370_10202# rowon_n[8] a_27974_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5694 a_20434_6508# col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5695 a_3878_2130# row_n[0] a_4370_2492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5696 VDD rowon_n[4] a_29982_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5697 a_16930_1126# VDD a_17422_1488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5698 a_15926_18194# VDD a_16418_18556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5699 a_27366_16226# rowon_n[14] a_26970_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5700 vcm a_2275_14202# a_5978_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5701 vcm a_2275_14202# a_16018_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5702 a_9994_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5703 a_9294_2170# col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5704 a_5886_18194# VDD a_6378_18556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5705 vcm a_2275_6170# a_35094_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5706 a_10906_2130# a_2275_2154# a_10998_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5707 a_28978_15182# a_2275_15206# a_29070_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5708 a_20034_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5709 VSS VDD a_23350_1166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5710 VSS row_n[3] a_22346_5182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5711 a_10998_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5712 a_33086_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5713 a_32386_5182# rowon_n[3] a_31990_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5714 a_23350_12210# col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5715 a_4882_4138# a_2275_4162# a_4974_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5716 a_26058_5142# a_2475_5166# a_25966_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5717 a_24450_8516# col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5718 a_22346_18234# col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5719 VDD rowon_n[6] a_33998_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5720 a_2161_13198# sample VDD VDD sky130_fd_pr__pfet_01v8 ad=3.42e+11p pd=2.97e+06u as=0p ps=0u w=1.2e+06u l=150000u
X5721 a_22442_14540# col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5722 VSS row_n[8] a_17326_10202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5723 a_22042_10162# a_2475_10186# a_21950_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5724 VSS a_2161_8178# a_2275_8178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.71e+11p ps=1.77e+06u w=600000u l=150000u
X5725 a_21950_6146# a_2275_6170# a_22042_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5726 VDD rowon_n[1] a_31990_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5727 a_22442_3496# col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5728 a_7894_11166# a_2275_11190# a_7986_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5729 a_17934_11166# a_2275_11190# a_18026_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5730 VSS row_n[8] a_7286_10202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5731 a_30986_18194# a_2275_18218# a_31078_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5732 VSS row_n[14] a_16322_16226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5733 a_21038_16186# a_2475_16210# a_20946_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5734 a_22954_10162# row_n[8] a_23446_10524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5735 VSS row_n[1] a_27366_3174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5736 VSS row_n[14] a_6282_16226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5737 a_19334_9198# rowon_n[7] a_18938_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5738 a_31382_9198# col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5739 a_13406_7512# col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5740 VSS row_n[4] a_5278_6186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5741 a_21950_16186# row_n[14] a_22442_16548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5742 VDD rowon_n[10] a_15926_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5743 VSS row_n[7] a_17326_9198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5744 a_1957_15206# VDD sample VSS sky130_fd_pr__nfet_01v8 ad=1.71e+11p pd=1.77e+06u as=0p ps=0u w=600000u l=150000u
X5745 a_16018_14178# a_2475_14202# a_15926_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5746 VDD rowon_n[10] a_5886_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5747 a_29470_6508# col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5748 a_11398_2492# col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5749 VDD VDD a_14922_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5750 a_5978_14178# a_2475_14202# a_5886_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5751 VDD VDD a_4882_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5752 a_15318_15222# col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5753 vcm a_2275_15206# a_20034_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5754 a_7986_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5755 VSS row_n[0] a_16322_2170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5756 a_30074_3134# a_2475_3158# a_29982_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5757 vcm a_2275_3158# a_20034_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5758 a_14010_17190# a_2475_17214# a_13918_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5759 a_5278_15222# col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5760 a_25966_8154# a_2275_8178# a_26058_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5761 a_27462_1488# col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5762 a_26970_4138# a_2275_4162# a_27062_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5763 a_3970_17190# a_2475_17214# a_3878_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5764 vcm a_2275_9182# a_9994_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5765 VDD rowon_n[7] a_18938_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5766 a_30986_9158# row_n[7] a_31478_9520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5767 a_31990_5142# row_n[3] a_32482_5504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5768 a_14410_17552# col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5769 a_10906_14178# row_n[12] a_11398_14540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5770 vcm a_2275_10186# a_10998_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5771 a_17422_9520# col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5772 VSS row_n[6] a_9294_8194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5773 a_18426_5504# col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5774 a_4370_17552# col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5775 a_22346_12210# rowon_n[10] a_21950_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5776 a_14922_13174# row_n[11] a_15414_13536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5777 a_26362_11206# rowon_n[9] a_25966_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5778 a_4882_13174# row_n[11] a_5374_13536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5779 a_18026_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5780 vcm a_2275_1150# a_25054_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5781 a_35094_1126# a_2475_1150# a_35002_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5782 a_1957_16210# VSS sample VDD sky130_fd_pr__pfet_01v8 ad=3.42e+11p pd=2.97e+06u as=0p ps=0u w=1.2e+06u l=150000u
X5783 a_7986_11166# a_2475_11190# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5784 a_1957_6170# VDD sample VSS sky130_fd_pr__nfet_01v8 ad=1.71e+11p pd=1.77e+06u as=0p ps=0u w=600000u l=150000u
X5785 vcm a_2275_4162# a_2966_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5786 a_34090_5142# a_2475_5166# a_33998_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5787 VDD rowon_n[8] a_21950_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5788 a_8898_9158# a_2275_9182# a_8990_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5789 a_17022_2130# a_2475_2154# a_16930_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5790 VSS row_n[15] a_20338_17230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5791 a_26970_16186# a_2275_16210# a_27062_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5792 a_31078_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5793 a_12306_6186# rowon_n[4] a_11910_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5794 a_29982_6146# a_2275_6170# a_30074_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5795 VDD rowon_n[5] a_22954_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5796 a_33998_2130# row_n[0] a_34490_2492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5797 VSS row_n[14] a_24354_16226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5798 a_21342_13214# col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5799 a_34394_12210# col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5800 a_14314_15222# rowon_n[13] a_13918_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5801 VSS row_n[10] a_11302_12210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5802 VDD rowon_n[0] a_20946_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5803 a_21038_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5804 a_19030_16186# a_2475_16210# a_18938_16186# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5805 a_4274_15222# rowon_n[13] a_3878_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5806 a_29982_13174# a_2275_13198# a_30074_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5807 VDD VDD a_22954_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5808 a_20434_15544# col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5809 a_8290_14218# rowon_n[12] a_7894_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5810 a_33486_14540# col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5811 vcm a_2275_12194# a_29070_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5812 VSS row_n[9] a_5278_11206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5813 VSS row_n[9] a_15318_11206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5814 a_20034_11166# a_2475_11190# a_19942_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5815 a_33086_10162# a_2475_10186# a_32994_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5816 a_20338_8194# col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5817 a_26362_2170# rowon_n[0] a_25966_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5818 a_21342_4178# col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5819 a_20946_11166# row_n[9] a_21438_11528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5820 a_10998_10162# a_2475_10186# a_10906_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5821 a_5978_9158# a_2475_9182# a_5886_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5822 VSS row_n[6] a_30378_8194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5823 a_4274_5182# rowon_n[3] a_3878_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5824 a_5278_1166# VSS a_4882_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5825 VSS row_n[2] a_31382_4178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5826 VDD rowon_n[12] a_9902_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5827 a_33998_10162# row_n[8] a_34490_10524# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5828 a_35002_4138# a_2275_4162# a_35094_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5829 a_17326_4178# rowon_n[2] a_16930_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5830 a_16322_8194# rowon_n[6] a_15926_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5831 vcm a_2275_8178# a_24050_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5832 vcm a_2275_2154# a_18026_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5833 VDD rowon_n[3] a_27974_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5834 VDD rowon_n[11] a_3878_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5835 VDD rowon_n[11] a_13918_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5836 a_11398_10524# col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5837 VDD rowon_n[6] a_5886_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5838 a_25054_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5839 a_26058_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5840 a_13310_16226# col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5841 VDD rowon_n[1] a_3878_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5842 a_31478_4500# col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5843 a_20946_4138# row_n[2] a_21438_4500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5844 a_12002_18194# a_2475_18218# a_11910_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5845 a_34090_18194# a_2475_18218# a_33998_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5846 a_3270_16226# col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5847 vcm a_2275_15206# a_31078_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5848 a_25358_6186# col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5849 a_35002_18194# VDD a_35494_18556# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5850 vcm a_2275_14202# a_35094_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5851 a_3270_9198# col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5852 a_11910_6146# row_n[4] a_12402_6508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5853 VSS row_n[4] a_35398_6186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5854 a_9294_3174# rowon_n[1] a_8898_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5855 VDD rowon_n[2] a_16930_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5856 a_8290_7190# rowon_n[5] a_7894_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5857 a_12402_18556# col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5858 a_19334_18234# VDD a_18938_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5859 a_20338_13214# rowon_n[11] a_19942_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5860 vcm a_2275_6170# a_29070_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5861 vcm a_2275_9182# a_6982_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5862 a_25054_15182# a_2475_15206# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5863 a_21950_12170# a_2275_12194# a_22042_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5864 a_14314_5182# col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5865 VDD VSS a_8898_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5866 a_29070_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5867 a_2874_9158# row_n[7] a_3366_9520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5868 a_3878_5142# row_n[3] a_4370_5504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5869 a_19942_1126# a_2275_1150# a_20034_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5870 VDD rowon_n[14] a_18938_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5871 VDD rowon_n[9] a_19942_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5872 a_15926_8154# row_n[6] a_16418_8516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5873 a_30074_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5874 a_9994_13174# a_2475_13198# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5875 VSS row_n[15] a_31382_17230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5876 a_2475_10186# a_1957_10186# VDD VDD sky130_fd_pr__pfet_01v8 ad=3.42e+11p pd=2.97e+06u as=0p ps=0u w=1.2e+06u l=150000u
X5877 a_13918_3134# row_n[1] a_14410_3496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5878 a_13310_10202# rowon_n[8] a_12914_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5879 a_12002_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5880 VSS row_n[14] a_35398_16226# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5881 a_32386_13214# col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5882 a_3270_10202# rowon_n[8] a_2874_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5883 a_18330_7190# col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5884 a_19334_3174# col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5885 vcm a_2275_4162# a_33086_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5886 a_26058_17190# a_2475_17214# a_25966_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5887 a_12306_16226# rowon_n[14] a_11910_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5888 VSS row_n[1] a_20338_3174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5889 a_7894_7150# row_n[5] a_8386_7512# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5890 a_30378_3174# rowon_n[1] a_29982_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5891 VDD VDD a_33998_18194# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5892 a_26970_17190# row_n[15] a_27462_17552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5893 a_31478_15544# col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5894 vcm a_2275_13198# a_27062_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5895 a_31078_11166# a_2475_11190# a_30986_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5896 a_34090_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5897 a_3878_15182# a_2275_15206# a_3970_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5898 a_13918_15182# a_2275_15206# a_14010_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5899 VSS row_n[7] a_10298_9198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5900 a_23046_7150# a_2475_7174# a_22954_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5901 a_22442_6508# col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5902 a_5886_2130# row_n[0] a_6378_2492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5903 a_17934_14178# a_2275_14202# a_18026_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5904 a_31990_11166# row_n[9] a_32482_11528# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5905 VDD rowon_n[4] a_31990_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5906 a_18938_1126# en_bit_n[2] a_19430_1488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5907 a_7894_14178# a_2275_14202# a_7986_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5908 a_20434_1488# en_bit_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5909 a_29982_14178# row_n[12] a_30474_14540# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5910 vcm a_2275_10186# a_30074_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5911 VDD VSS a_29982_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5912 a_12914_2130# a_2275_2154# a_13006_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5913 VSS VDD a_25358_1166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5914 VSS row_n[3] a_24354_5182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5915 a_10394_9520# col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5916 a_11398_5504# col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5917 a_35398_1166# VSS a_35002_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5918 VSS row_n[2] a_3270_4178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5919 a_34394_5182# rowon_n[3] a_33998_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5920 a_18330_13214# rowon_n[11] a_17934_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5921 a_28978_10162# a_2275_10186# a_29070_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5922 a_28066_5142# a_2475_5166# a_27974_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5923 vcm a_2275_16210# a_8990_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5924 vcm a_2275_16210# a_19030_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5925 a_23958_6146# a_2275_6170# a_24050_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5926 a_24450_3496# col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5927 VDD rowon_n[1] a_33998_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5928 a_23046_16186# a_2475_16210# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5929 VDD rowon_n[9] a_17934_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5930 VSS row_n[1] a_29374_3174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5931 a_3366_4500# col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5932 a_33390_9198# col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5933 a_15414_7512# col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5934 VSS row_n[15] a_29374_17230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5935 a_33390_15222# rowon_n[13] a_32994_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5936 VSS row_n[10] a_30378_12210# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5937 a_16018_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5938 VSS row_n[4] a_7286_6186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5939 a_7986_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5940 a_18026_14178# a_2475_14202# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5941 VSS row_n[9] a_34394_11206# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5942 a_32386_2170# col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5943 a_2161_1150# sample VDD VDD sky130_fd_pr__pfet_01v8 ad=3.42e+11p pd=2.97e+06u as=0p ps=0u w=1.2e+06u l=150000u
X5944 a_13406_2492# col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5945 a_3970_4138# a_2475_4162# a_3878_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5946 a_9994_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5947 a_25054_12170# a_2475_12194# a_24962_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5948 a_11302_11206# rowon_n[9] a_10906_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5949 a_1957_10186# VDD sample VSS sky130_fd_pr__nfet_01v8 ad=1.71e+11p pd=1.77e+06u as=0p ps=0u w=600000u l=150000u
X5950 a_27974_8154# a_2275_8178# a_28066_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5951 a_29470_1488# col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5952 VSS row_n[0] a_18330_2170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5953 a_32082_3134# a_2475_3158# a_31990_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5954 a_28978_4138# a_2275_4162# a_29070_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5955 a_29470_15544# col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5956 VDD rowon_n[11] a_32994_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5957 a_25966_12170# row_n[10] a_26458_12532# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5958 a_29070_11166# a_2475_11190# a_28978_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5959 a_30474_10524# col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5960 a_32994_9158# row_n[7] a_33486_9520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5961 a_33998_5142# row_n[3] a_34490_5504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5962 a_9994_10162# a_2475_10186# a_9902_10162# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5963 a_10298_4178# rowon_n[2] a_9902_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5964 a_11910_16186# a_2275_16210# a_12002_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5965 VDD rowon_n[12] a_8898_14178# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5966 vcm a_2275_2154# a_10998_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5967 VDD rowon_n[3] a_20946_5142# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5968 a_16930_7150# a_2275_7174# a_17022_7150# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5969 vcm a_2275_17214# a_23046_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5970 a_8290_17230# col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5971 a_18330_17230# col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5972 vcm a_2275_4162# a_4974_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5973 VDD rowon_n[2] a_9902_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5974 vcm a_2275_12194# a_14010_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5975 vcm a_2275_12194# a_3970_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5976 a_14314_6186# rowon_n[4] a_13918_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5977 vcm a_2275_6170# a_22042_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5978 a_17934_15182# row_n[13] a_18426_15544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5979 a_29374_13214# rowon_n[11] a_28978_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5980 vcm a_2275_11190# a_18026_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5981 VSS row_n[8] a_26362_10202# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5982 a_7894_15182# row_n[13] a_8386_15544# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5983 vcm a_2275_11190# a_7986_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5984 a_26970_11166# a_2275_11190# a_27062_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5985 VDD rowon_n[4] a_3878_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5986 VDD rowon_n[0] a_22954_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5987 a_23046_5142# a_2475_5166# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5988 VDD rowon_n[10] a_24962_12170# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5989 a_28370_2170# rowon_n[0] a_27974_2130# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5990 VSS row_n[2] a_33390_4178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5991 a_23350_4178# col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5992 VDD rowon_n[9] a_28978_11166# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5993 a_7986_9158# a_2475_9182# a_7894_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5994 VSS row_n[6] a_32386_8194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5995 a_6282_5182# rowon_n[3] a_5886_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5996 a_7286_1166# VSS a_6890_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5997 VSS a_2161_18218# a_2275_18218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.71e+11p ps=1.77e+06u w=600000u l=150000u
X5998 vcm a_2275_8178# a_26058_8154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5999 vcm a_2275_4162# a_27062_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6000 VSS VDD a_27366_18234# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6001 a_31382_16226# rowon_n[14] a_30986_16186# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6002 a_24354_15222# col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6003 VDD rowon_n[6] a_7894_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6004 a_2475_6170# a_1957_6170# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.71e+11p pd=1.77e+06u as=0p ps=0u w=600000u l=150000u
X6005 a_17326_17230# rowon_n[15] a_16930_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6006 a_28370_14218# col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6007 a_11302_7190# col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6008 a_28066_3134# a_2475_3158# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6009 a_12306_3174# col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6010 a_7286_17230# rowon_n[15] a_6890_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6011 a_19942_16186# a_2275_16210# a_20034_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6012 a_32994_15182# a_2275_15206# a_33086_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6013 a_31990_9158# a_2275_9182# a_32082_9158# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6014 a_27062_7150# a_2475_7174# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6015 a_22954_4138# row_n[2] a_23446_4500# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6016 a_3970_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6017 a_14010_18194# a_2475_18218# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6018 a_23446_17552# col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6019 VSS row_n[11] a_8290_13214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6020 VSS row_n[11] a_18330_13214# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6021 a_23046_13174# a_2475_13198# a_22954_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6022 VDD rowon_n[1] a_5886_3134# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6023 a_33486_4500# col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6024 a_13918_6146# row_n[4] a_14410_6508# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6025 a_27462_16548# col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6026 a_23958_13174# row_n[11] a_24450_13536# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6027 a_18026_11166# a_2475_11190# a_17934_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6028 a_5278_9198# col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6029 a_7986_11166# a_2475_11190# a_7894_11166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6030 VDD rowon_n[13] a_6890_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6031 VDD rowon_n[13] a_16930_15182# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6032 vcm a_2275_9182# a_8990_9158# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6033 a_11910_1126# VDD a_12402_1488# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6034 a_18426_11528# col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6035 a_4274_2170# col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6036 a_8386_11528# col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6037 vcm a_2275_6170# a_30074_6146# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6038 a_16322_5182# col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6039 a_17326_1166# col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6040 a_16322_18234# col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6041 vcm a_2275_18218# a_21038_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6042 a_6282_18234# col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6043 vcm a_2275_17214# a_34090_17190# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6044 a_5886_5142# row_n[3] a_6378_5504# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6045 a_4882_9158# row_n[7] a_5374_9520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6046 a_17934_8154# row_n[6] a_18426_8516# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6047 a_25054_10162# a_2475_10186# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6048 a_32082_1126# a_2475_1150# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6049 a_21038_5142# a_2475_5166# a_20946_5142# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6050 a_11910_17190# row_n[15] a_12402_17552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6051 vcm a_2275_13198# a_12002_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6052 a_14010_2130# a_2475_2154# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6053 a_15926_3134# row_n[1] a_16418_3496# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6054 a_5886_16186# row_n[14] a_6378_16548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6055 a_15926_16186# row_n[14] a_16418_16548# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6056 a_27366_14218# rowon_n[12] a_26970_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6057 a_27366_9198# col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6058 vcm a_2275_4162# a_35094_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6059 a_28066_17190# a_2475_17214# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6060 a_28978_13174# a_2275_13198# a_29070_13174# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6061 VSS row_n[1] a_22346_3174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6062 a_31382_7190# rowon_n[5] a_30986_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6063 a_32386_3174# rowon_n[1] a_31990_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6064 a_23350_10202# col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6065 VSS row_n[7] a_12306_9198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6066 a_26058_3134# a_2475_3158# a_25966_3134# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6067 a_25054_7150# a_2475_7174# a_24962_7150# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6068 a_24450_6508# col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6069 a_7894_2130# row_n[0] a_8386_2492# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6070 a_22346_16226# col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6071 a_16322_12210# rowon_n[10] a_15926_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6072 a_26970_9158# row_n[7] a_27462_9520# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6073 VDD rowon_n[4] a_33998_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6074 a_6282_12210# rowon_n[10] a_5886_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6075 a_2161_11190# sample VDD VDD sky130_fd_pr__pfet_01v8 ad=3.42e+11p pd=2.97e+06u as=0p ps=0u w=1.2e+06u l=150000u
X6076 a_13918_10162# a_2275_10186# a_14010_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6077 a_2966_9158# a_2475_9182# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6078 VSS row_n[0] a_11302_2170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6079 a_22442_12532# col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6080 a_3878_10162# a_2275_10186# a_3970_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6081 a_20946_8154# a_2275_8178# a_21038_8154# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6082 a_22442_1488# col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6083 VDD VSS a_31990_1126# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6084 a_21950_4138# a_2275_4162# a_22042_4138# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6085 a_5278_18234# VDD a_4882_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6086 a_15318_18234# VDD a_14922_18194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6087 a_31078_8154# a_2475_8178# vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6088 a_14922_2130# a_2275_2154# a_15014_2130# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6089 a_21438_18556# col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6090 a_30986_16186# a_2275_16210# a_31078_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6091 VSS row_n[12] a_16322_14218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6092 a_21038_14178# a_2475_14202# a_20946_14178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6093 VSS VDD a_27366_1166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6094 VSS row_n[12] a_6282_14218# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6095 a_12402_9520# col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6096 VSS row_n[6] a_4274_8194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6097 a_13406_5504# col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6098 VSS row_n[2] a_5278_4178# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6099 a_16930_17190# a_2275_17214# a_17022_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6100 VDD rowon_n[8] a_15926_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6101 a_6890_17190# a_2275_17214# a_6982_17190# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6102 VDD rowon_n[8] a_5886_10162# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6103 VSS row_n[15] a_4274_17230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6104 VSS row_n[15] a_14314_17230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6105 VDD rowon_n[14] a_14922_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6106 VDD rowon_n[14] a_4882_16186# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6107 a_15318_13214# col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6108 vcm a_2275_13198# a_20034_13174# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6109 vcm a_2275_1150# a_20034_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6110 a_30074_1126# a_2475_1150# a_29982_1126# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6111 a_19942_17190# row_n[15] a_20434_17552# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6112 a_14010_15182# a_2475_15206# a_13918_15182# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6113 a_5278_13214# col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6114 vcm a_2275_12194# a_33086_12170# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6115 a_25966_6146# a_2275_6170# a_26058_6146# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
C0 a_27974_10162# rowoff_n[8] 0.46fF
C1 a_2275_5166# vcm 7.71fF
C2 a_31078_13174# rowoff_n[11] 1.25fF
C3 a_25054_4138# col[22] 0.38fF
C4 a_2275_1150# a_18938_1126# 0.17fF
C5 a_26058_15182# vcm 0.89fF
C6 a_22954_5142# VDD 0.29fF
C7 m2_25828_946# VDD 3.85fF
C8 a_2966_9158# ctop 4.82fF
C9 col[14] rowoff_n[12] 0.25fF
C10 a_2275_2154# rowon_n[0] 1.99fF
C11 a_10998_15182# a_12002_15182# 0.86fF
C12 a_2475_15206# a_21038_15182# 0.68fF
C13 a_20338_4178# col_n[17] 0.11fF
C14 a_16322_9198# vcm 0.24fF
C15 a_3970_15182# col_n[1] 0.34fF
C16 a_30378_16226# col_n[27] 0.11fF
C17 a_2475_12194# col[5] 0.22fF
C18 a_2275_3158# a_33998_3134# 0.17fF
C19 a_6982_18194# vcm 0.15fF
C20 a_29070_4138# ctop 4.91fF
C21 a_2475_1150# col[10] 0.22fF
C22 a_25054_9158# row_n[7] 0.43fF
C23 a_26058_16186# m2_26256_16434# 0.19fF
C24 a_29982_8154# a_30074_8154# 0.45fF
C25 a_24962_13174# rowon_n[11] 0.14fF
C26 a_2275_12194# a_12002_12170# 0.71fF
C27 a_9902_3134# vcm 0.18fF
C28 a_35002_3134# rowon_n[1] 0.14fF
C29 a_2275_7174# col_n[17] 0.17fF
C30 m2_26832_18014# m2_27836_18014# 0.86fF
C31 a_31382_13214# vcm 0.24fF
C32 a_14010_2130# col[11] 0.38fF
C33 a_9994_7150# ctop 4.91fF
C34 a_24050_14178# col[21] 0.38fF
C35 a_18938_12170# VDD 0.29fF
C36 m2_31852_946# m2_32280_1374# 0.19fF
C37 a_2475_17214# rowon_n[15] 0.40fF
C38 a_2475_9182# a_4882_9158# 0.41fF
C39 a_2275_9182# a_3878_9158# 0.17fF
C40 a_2275_15206# col[2] 0.17fF
C41 a_2275_4162# col[7] 0.17fF
C42 a_2275_14202# a_27062_14178# 0.71fF
C43 a_12002_7150# rowon_n[5] 0.45fF
C44 a_24962_7150# vcm 0.18fF
C45 a_19030_14178# rowoff_n[12] 1.84fF
C46 a_21038_2130# a_22042_2130# 0.86fF
C47 a_9294_2170# col_n[6] 0.11fF
C48 a_12306_16226# vcm 0.24fF
C49 a_2475_14202# col[22] 0.22fF
C50 a_19334_14218# col_n[16] 0.11fF
C51 a_17022_14178# m2_17220_14426# 0.19fF
C52 a_2475_3158# col[27] 0.22fF
C53 a_25054_11166# ctop 4.91fF
C54 a_33998_16186# VDD 0.29fF
C55 a_2475_11190# a_19942_11166# 0.41fF
C56 a_2275_11190# a_17326_11206# 0.15fF
C57 a_10906_11166# a_10998_11166# 0.45fF
C58 a_2475_18218# col[13] 0.22fF
C59 a_14010_2130# m2_14208_2378# 0.19fF
C60 a_5886_10162# vcm 0.18fF
C61 a_23046_16186# row_n[14] 0.43fF
C62 a_12002_4138# a_12002_3134# 0.84fF
C63 a_1957_18218# a_2275_18218# 0.19fF
C64 a_2275_8178# a_10906_8154# 0.17fF
C65 a_5978_14178# ctop 4.91fF
C66 a_33086_6146# row_n[4] 0.43fF
C67 a_13006_12170# col[10] 0.38fF
C68 a_2275_13198# a_32386_13214# 0.15fF
C69 a_2475_13198# a_35002_13174# 0.41fF
C70 a_32994_10162# rowon_n[8] 0.14fF
C71 a_2275_17214# col[19] 0.17fF
C72 a_2275_6170# col[24] 0.17fF
C73 a_2275_18218# col[4] 0.17fF
C74 a_28066_8154# col_n[25] 0.34fF
C75 a_20946_14178# vcm 0.18fF
C76 a_17022_4138# VDD 2.99fF
C77 a_7986_12170# m2_8184_12418# 0.19fF
C78 a_2475_5166# a_2874_5142# 0.41fF
C79 a_1957_5166# a_2275_5166# 0.19fF
C80 a_8290_12210# col_n[5] 0.11fF
C81 a_2275_10186# a_25966_10162# 0.17fF
C82 a_9994_14178# rowon_n[12] 0.45fF
C83 a_25966_15182# a_26058_15182# 0.45fF
C84 row_n[12] sample_n 0.16fF
C85 ctop col[5] 0.13fF
C86 a_6982_15182# rowoff_n[13] 2.42fF
C87 a_20034_4138# rowon_n[2] 0.45fF
C88 a_27062_8154# m2_27260_8402# 0.19fF
C89 a_34394_18234# vcm 0.25fF
C90 a_32082_8154# VDD 1.44fF
C91 a_8990_7150# rowoff_n[5] 2.33fF
C92 a_2475_7174# a_18026_7150# 0.68fF
C93 a_27062_8154# a_27062_7150# 0.84fF
C94 m2_2736_1950# col_n[0] 0.33fF
C95 a_3970_2130# vcm 0.89fF
C96 a_18026_5142# rowoff_n[3] 1.89fF
C97 a_2275_4162# a_8990_4138# 0.71fF
C98 a_17022_6146# col_n[14] 0.34fF
C99 a_31078_13174# row_n[11] 0.43fF
C100 a_13006_11166# VDD 3.40fF
C101 a_2275_16210# col_n[6] 0.17fF
C102 a_2475_9182# a_33086_9158# 0.68fF
C103 a_30986_17190# rowon_n[15] 0.14fF
C104 a_17022_9158# a_18026_9158# 0.86fF
C105 a_2275_5166# col_n[11] 0.17fF
C106 a_27062_3134# rowoff_n[1] 1.45fF
C107 a_19030_6146# vcm 0.89fF
C108 a_6890_18194# a_6982_18194# 0.11fF
C109 a_18026_6146# m2_18224_6394# 0.19fF
C110 col[25] rowoff_n[12] 0.18fF
C111 m2_16792_18014# col_n[14] 0.33fF
C112 a_2275_6170# a_24050_6146# 0.71fF
C113 a_2275_2154# col[1] 0.17fF
C114 a_28066_15182# VDD 1.85fF
C115 a_7986_11166# a_7986_10162# 0.84fF
C116 m2_20808_18014# vcm 0.71fF
C117 a_2475_15206# a_2966_15182# 0.65fF
C118 a_2161_15206# a_2275_15206# 0.17fF
C119 a_2475_12194# col[16] 0.22fF
C120 m2_2736_946# m3_2868_1078# 4.41fF
C121 a_18026_11166# rowon_n[9] 0.45fF
C122 a_34090_10162# vcm 0.89fF
C123 a_2475_1150# col[21] 0.22fF
C124 a_2275_3158# a_14314_3174# 0.15fF
C125 a_2475_3158# a_16930_3134# 0.41fF
C126 a_2275_1150# m2_10768_946# 0.51fF
C127 m3_5880_1078# ctop 0.21fF
C128 a_5978_4138# col_n[3] 0.34fF
C129 a_32386_5182# col_n[29] 0.11fF
C130 a_16018_16186# col_n[13] 0.34fF
C131 a_32082_13174# a_33086_13174# 0.86fF
C132 a_2275_7174# col_n[28] 0.17fF
C133 a_24354_4178# vcm 0.24fF
C134 a_19942_11166# rowoff_n[9] 0.55fF
C135 a_2275_17214# a_17934_17190# 0.17fF
C136 col[9] rowoff_n[13] 0.29fF
C137 a_8990_4138# m2_9188_4386# 0.19fF
C138 a_15014_13174# vcm 0.89fF
C139 a_11910_3134# VDD 0.29fF
C140 a_16930_5142# a_17022_5142# 0.45fF
C141 a_2475_5166# a_31990_5142# 0.41fF
C142 a_2275_5166# a_29374_5182# 0.15fF
C143 a_2275_15206# col[13] 0.17fF
C144 a_5886_5142# rowon_n[3] 0.14fF
C145 a_2275_18218# a_27974_18194# 0.17fF
C146 a_2275_4162# col[18] 0.17fF
C147 a_28978_9158# rowoff_n[7] 0.44fF
C148 a_23046_15182# a_23046_14178# 0.84fF
C149 a_2475_14202# a_9994_14178# 0.68fF
C150 a_26058_3134# col[23] 0.38fF
C151 a_5278_7190# vcm 0.24fF
C152 a_2275_2154# a_22954_2130# 0.17fF
C153 a_30074_17190# vcm 0.89fF
C154 a_18026_2130# ctop 4.95fF
C155 a_26970_7150# VDD 0.29fF
C156 a_2475_18218# col[24] 0.22fF
C157 a_2966_14178# m2_1732_13998# 0.86fF
C158 a_21342_3174# col_n[18] 0.11fF
C159 a_32994_2130# vcm 0.18fF
C160 a_13006_16186# a_14010_16186# 0.86fF
C161 a_2475_16210# a_25054_16186# 0.68fF
C162 a_4974_14178# col_n[2] 0.34fF
C163 a_31382_15222# col_n[28] 0.11fF
C164 a_20338_11206# vcm 0.24fF
C165 a_18426_1488# VDD 0.15fF
C166 a_26058_8154# rowon_n[6] 0.45fF
C167 a_33086_6146# ctop 4.91fF
C168 a_7894_10162# VDD 0.29fF
C169 a_2275_17214# col[30] 0.17fF
C170 a_2275_17214# m2_34864_17010# 0.51fF
C171 a_31990_9158# a_32082_9158# 0.45fF
C172 m2_1732_3958# sample_n 0.12fF
C173 a_2275_18218# col[15] 0.17fF
C174 a_2275_13198# a_16018_13174# 0.71fF
C175 a_13918_5142# vcm 0.18fF
C176 a_7894_12170# rowoff_n[10] 0.68fF
C177 a_2275_18218# m2_4744_18014# 0.51fF
C178 a_3970_8154# row_n[6] 0.43fF
C179 a_2275_14202# vcm 7.71fF
C180 a_25054_13174# col[22] 0.38fF
C181 a_2275_3158# col_n[5] 0.17fF
C182 a_14010_9158# ctop 4.91fF
C183 a_22954_14178# VDD 0.29fF
C184 a_2475_10186# a_8898_10162# 0.41fF
C185 a_2275_10186# a_6282_10202# 0.15fF
C186 a_13918_2130# rowon_n[0] 0.14fF
C187 ctop col[16] 0.13fF
C188 rowon_n[6] sample_n 0.15fF
C189 a_2275_15206# a_31078_15182# 0.71fF
C190 a_10298_1166# col_n[7] 0.11fF
C191 a_28978_9158# vcm 0.18fF
C192 a_23958_16186# rowoff_n[14] 0.50fF
C193 a_20338_13214# col_n[17] 0.11fF
C194 a_23046_3134# a_24050_3134# 0.86fF
C195 a_16322_18234# vcm 0.25fF
C196 a_35002_16186# m2_34864_16006# 0.33fF
C197 m2_34864_9982# rowoff_n[8] 1.01fF
C198 a_29070_13174# ctop 4.91fF
C199 a_2475_10186# col[10] 0.22fF
C200 a_2475_12194# a_23958_12170# 0.41fF
C201 a_2275_12194# a_21342_12210# 0.15fF
C202 a_12914_12170# a_13006_12170# 0.45fF
C203 a_24050_15182# rowon_n[13] 0.45fF
C204 a_9902_12170# vcm 0.18fF
C205 a_5978_2130# VDD 4.13fF
C206 a_2275_16210# col_n[17] 0.17fF
C207 a_14010_5142# a_14010_4138# 0.84fF
C208 a_2275_5166# col_n[22] 0.17fF
C209 a_34090_5142# rowon_n[3] 0.45fF
C210 a_14010_11166# col[11] 0.38fF
C211 a_2275_9182# a_14922_9158# 0.17fF
C212 a_9994_16186# ctop 4.91fF
C213 a_2475_18218# m2_30848_18014# 0.62fF
C214 a_2966_14178# a_2966_13174# 0.84fF
C215 a_2475_15206# row_n[13] 0.48fF
C216 a_29070_7150# col_n[26] 0.34fF
C217 a_2275_13198# col[7] 0.17fF
C218 a_2275_2154# col[12] 0.17fF
C219 a_24962_16186# vcm 0.18fF
C220 a_21038_6146# VDD 2.58fF
C221 a_12002_5142# row_n[3] 0.43fF
C222 a_9294_11206# col_n[6] 0.11fF
C223 a_3970_6146# a_4974_6146# 0.86fF
C224 a_2475_6170# a_6982_6146# 0.68fF
C225 a_11910_9158# rowon_n[7] 0.14fF
C226 a_2275_11190# a_29982_11166# 0.17fF
C227 a_2475_12194# col[27] 0.22fF
C228 a_27062_1126# vcm 0.15fF
C229 a_27974_16186# a_28066_16186# 0.45fF
C230 m2_1732_7974# rowon_n[6] 0.43fF
C231 a_11910_17190# rowoff_n[15] 0.64fF
C232 m2_24824_18014# VDD 2.96fF
C233 a_9994_6146# rowoff_n[4] 2.28fF
C234 a_2475_9182# VDD 41.96fF
C235 a_32082_17190# m2_32280_17438# 0.19fF
C236 a_2475_8178# a_22042_8154# 0.68fF
C237 a_29070_9158# a_29070_8154# 0.84fF
C238 col[20] rowoff_n[13] 0.21fF
C239 a_7986_4138# vcm 0.89fF
C240 a_19030_4138# rowoff_n[2] 1.84fF
C241 col_n[2] rowoff_n[8] 0.32fF
C242 sample rowoff_n[4] 0.22fF
C243 col_n[3] rowoff_n[9] 0.32fF
C244 col_n[1] rowoff_n[7] 0.33fF
C245 VDD rowoff_n[3] 87.22fF
C246 vcm rowoff_n[6] 2.43fF
C247 col_n[0] rowoff_n[5] 0.34fF
C248 a_2275_15206# col[24] 0.17fF
C249 a_18026_5142# col_n[15] 0.34fF
C250 a_2275_4162# col[29] 0.17fF
C251 a_32082_12170# rowon_n[10] 0.45fF
C252 a_28066_17190# col_n[25] 0.34fF
C253 a_2275_5166# a_13006_5142# 0.71fF
C254 a_17022_13174# VDD 2.99fF
C255 a_2275_18218# a_8290_18234# 0.15fF
C256 a_19030_10162# a_20034_10162# 0.86fF
C257 a_28066_2130# rowoff_n[0] 1.40fF
C258 a_2275_1150# col_n[0] 0.17fF
C259 a_23046_8154# vcm 0.89fF
C260 a_9994_12170# row_n[10] 0.43fF
C261 a_2275_2154# a_3270_2170# 0.15fF
C262 a_2475_2154# a_5886_2130# 0.41fF
C263 m2_18800_18014# m3_18932_18146# 4.43fF
C264 a_9902_16186# rowon_n[14] 0.14fF
C265 a_23046_15182# m2_23244_15430# 0.19fF
C266 a_2275_7174# a_28066_7150# 0.71fF
C267 a_20034_2130# row_n[0] 0.43fF
C268 a_32082_17190# VDD 1.44fF
C269 col[4] rowoff_n[14] 0.32fF
C270 a_9994_12170# a_9994_11166# 0.84fF
C271 a_19942_6146# rowon_n[4] 0.14fF
C272 a_13310_2170# vcm 0.24fF
C273 a_2275_16210# a_6890_16186# 0.17fF
C274 a_3970_11166# vcm 0.89fF
C275 a_35002_2130# VDD 0.36fF
C276 a_2475_8178# col[4] 0.22fF
C277 a_2475_4162# a_20946_4138# 0.41fF
C278 a_2275_4162# a_18330_4178# 0.15fF
C279 a_6982_3134# col_n[4] 0.34fF
C280 a_33390_4178# col_n[30] 0.11fF
C281 a_2275_18218# col[26] 0.17fF
C282 a_17022_15182# col_n[14] 0.34fF
C283 a_20946_10162# rowoff_n[8] 0.54fF
C284 a_2275_14202# col_n[11] 0.17fF
C285 a_28370_6186# vcm 0.24fF
C286 a_24050_13174# rowoff_n[11] 1.59fF
C287 a_2275_3158# col_n[16] 0.17fF
C288 a_2275_1150# a_11910_1126# 0.17fF
C289 a_19030_15182# vcm 0.89fF
C290 a_15926_5142# VDD 0.29fF
C291 a_14010_13174# m2_14208_13422# 0.19fF
C292 a_2275_6170# a_33390_6186# 0.15fF
C293 a_18938_6146# a_19030_6146# 0.45fF
C294 vcm col_n[1] 3.19fF
C295 VDD col_n[4] 15.44fF
C296 row_n[1] sample_n 0.16fF
C297 ctop col[27] 0.13fF
C298 a_29982_8154# rowoff_n[6] 0.43fF
C299 a_2275_11190# col[1] 0.17fF
C300 a_27062_2130# col[24] 0.38fF
C301 a_2475_15206# a_14010_15182# 0.68fF
C302 a_25054_16186# a_25054_15182# 0.84fF
C303 a_9294_9198# vcm 0.24fF
C304 m2_31852_18014# col[29] 0.37fF
C305 a_33086_9158# m2_33284_9406# 0.19fF
C306 a_2275_3158# a_26970_3134# 0.17fF
C307 a_22042_4138# ctop 4.91fF
C308 a_2275_1150# m2_33860_946# 0.34fF
C309 a_12914_1126# m2_12776_946# 0.31fF
C310 a_2475_10186# col[21] 0.22fF
C311 a_30986_9158# VDD 0.29fF
C312 a_18026_9158# row_n[7] 0.43fF
C313 a_17934_13174# rowon_n[11] 0.14fF
C314 a_22346_2170# col_n[19] 0.11fF
C315 a_2275_12194# a_4974_12170# 0.71fF
C316 a_3878_12170# a_3970_12170# 0.45fF
C317 a_32386_14218# col_n[29] 0.11fF
C318 a_5978_13174# col_n[3] 0.34fF
C319 a_27974_3134# rowon_n[1] 0.14fF
C320 a_15014_17190# a_16018_17190# 0.86fF
C321 a_2475_17214# a_29070_17190# 0.68fF
C322 a_2275_16210# col_n[28] 0.17fF
C323 m2_19804_18014# m2_20808_18014# 0.86fF
C324 a_24354_13214# vcm 0.24fF
C325 a_4974_11166# m2_5172_11414# 0.19fF
C326 a_11910_12170# VDD 0.29fF
C327 m2_24824_946# m2_25252_1374# 0.19fF
C328 a_33998_10162# a_34090_10162# 0.45fF
C329 a_2275_13198# col[18] 0.17fF
C330 a_2275_14202# a_20034_14178# 0.71fF
C331 a_2275_2154# col[23] 0.17fF
C332 m2_1732_6970# m2_2160_7398# 0.19fF
C333 a_4974_7150# rowon_n[5] 0.45fF
C334 a_17934_7150# vcm 0.18fF
C335 a_12002_14178# rowoff_n[12] 2.18fF
C336 a_26058_12170# col[23] 0.38fF
C337 a_24050_7150# m2_24248_7398# 0.19fF
C338 a_2475_2154# a_34090_2130# 0.68fF
C339 a_5278_16226# vcm 0.24fF
C340 a_2966_6146# VDD 4.45fF
C341 a_18026_11166# ctop 4.91fF
C342 a_26970_16186# VDD 0.29fF
C343 a_2475_11190# a_12914_11166# 0.41fF
C344 a_2275_11190# a_10298_11206# 0.15fF
C345 a_2275_16210# a_35094_16186# 0.14fF
C346 a_21342_12210# col_n[18] 0.11fF
C347 a_32994_11166# vcm 0.18fF
C348 a_16018_16186# row_n[14] 0.43fF
C349 a_25054_4138# a_26058_4138# 0.86fF
C350 col[31] rowoff_n[13] 0.14fF
C351 a_2874_8154# a_2966_8154# 0.45fF
C352 a_33086_15182# ctop 4.91fF
C353 a_26058_6146# row_n[4] 0.43fF
C354 a_25966_10162# rowon_n[8] 0.14fF
C355 a_2275_13198# a_25358_13214# 0.15fF
C356 a_2475_13198# a_27974_13174# 0.41fF
C357 a_14922_13174# a_15014_13174# 0.45fF
C358 col_n[11] rowoff_n[6] 0.26fF
C359 col_n[14] rowoff_n[9] 0.24fF
C360 col_n[7] rowoff_n[2] 0.29fF
C361 col_n[10] rowoff_n[5] 0.27fF
C362 col_n[5] rowoff_n[0] 0.30fF
C363 col_n[8] rowoff_n[3] 0.28fF
C364 col_n[12] rowoff_n[7] 0.25fF
C365 col_n[9] rowoff_n[4] 0.27fF
C366 col_n[6] rowoff_n[1] 0.29fF
C367 col_n[13] rowoff_n[8] 0.24fF
C368 a_15014_5142# m2_15212_5390# 0.19fF
C369 a_13918_14178# vcm 0.18fF
C370 a_9994_4138# VDD 3.71fF
C371 a_2275_12194# m2_1732_11990# 0.27fF
C372 a_15014_10162# col[12] 0.38fF
C373 a_16018_6146# a_16018_5142# 0.84fF
C374 a_2275_12194# col_n[5] 0.17fF
C375 a_2275_10186# a_18938_10162# 0.17fF
C376 a_2275_1150# col_n[10] 0.17fF
C377 a_2874_14178# rowon_n[12] 0.14fF
C378 a_30074_6146# col_n[27] 0.34fF
C379 m2_34864_10986# m2_34864_9982# 0.84fF
C380 a_13006_4138# rowon_n[2] 0.45fF
C381 a_10298_10202# col_n[7] 0.11fF
C382 a_28978_18194# vcm 0.18fF
C383 col[15] rowoff_n[14] 0.25fF
C384 a_25054_8154# VDD 2.16fF
C385 a_2475_7174# rowoff_n[5] 4.75fF
C386 a_2475_7174# a_10998_7150# 0.68fF
C387 a_5978_7150# a_6982_7150# 0.86fF
C388 a_1957_2154# row_n[0] 0.29fF
C389 sample rowoff_n[10] 0.22fF
C390 a_2275_12194# a_33998_12170# 0.17fF
C391 a_31078_3134# vcm 0.89fF
C392 a_29982_17190# a_30074_17190# 0.45fF
C393 a_2475_8178# col[15] 0.22fF
C394 a_5978_3134# m2_6176_3382# 0.19fF
C395 a_10998_5142# rowoff_n[3] 2.23fF
C396 a_2475_4162# a_2275_4162# 2.96fF
C397 a_1957_4162# a_2161_4162# 0.11fF
C398 a_24050_13174# row_n[11] 0.43fF
C399 a_5978_11166# VDD 4.13fF
C400 m2_25828_946# m3_25960_1078# 4.41fF
C401 a_2475_9182# a_26058_9158# 0.68fF
C402 a_31078_10162# a_31078_9158# 0.84fF
C403 a_23958_17190# rowon_n[15] 0.14fF
C404 a_3970_8154# col[1] 0.38fF
C405 a_2275_14202# col_n[22] 0.17fF
C406 a_2275_3158# col_n[27] 0.17fF
C407 a_34090_3134# row_n[1] 0.43fF
C408 a_20034_3134# rowoff_n[1] 1.79fF
C409 a_2275_10186# rowoff_n[8] 0.81fF
C410 a_33998_7150# rowon_n[5] 0.14fF
C411 a_12002_6146# vcm 0.89fF
C412 a_19030_4138# col_n[16] 0.34fF
C413 VDD col_n[15] 12.25fF
C414 vcm col_n[12] 3.22fF
C415 a_29070_16186# col_n[26] 0.34fF
C416 a_2275_11190# col[12] 0.17fF
C417 a_2275_6170# a_17022_6146# 0.71fF
C418 a_34090_14178# m2_34864_13998# 0.86fF
C419 a_21038_15182# VDD 2.58fF
C420 a_21038_11166# a_22042_11166# 0.86fF
C421 m2_6752_18014# vcm 0.71fF
C422 a_10998_11166# rowon_n[9] 0.45fF
C423 a_27062_10162# vcm 0.89fF
C424 a_5886_3134# a_5978_3134# 0.45fF
C425 a_2475_3158# a_9902_3134# 0.41fF
C426 a_2275_3158# a_7286_3174# 0.15fF
C427 a_24050_2130# m2_23820_946# 0.84fF
C428 m3_34996_13126# ctop 0.22fF
C429 a_2275_8178# a_32082_8154# 0.71fF
C430 a_12002_13174# a_12002_12170# 0.84fF
C431 a_17326_4178# vcm 0.24fF
C432 a_12914_11166# rowoff_n[9] 0.63fF
C433 a_2275_17214# a_10906_17190# 0.17fF
C434 a_7986_13174# vcm 0.89fF
C435 a_4882_3134# VDD 0.29fF
C436 a_7986_2130# col_n[5] 0.34fF
C437 a_2475_5166# a_24962_5142# 0.41fF
C438 a_2275_5166# a_22346_5182# 0.15fF
C439 a_18026_14178# col_n[15] 0.34fF
C440 a_2275_13198# col[29] 0.17fF
C441 a_2275_18218# a_20946_18194# 0.17fF
C442 a_32082_10162# row_n[8] 0.43fF
C443 a_21950_9158# rowoff_n[7] 0.52fF
C444 a_31990_14178# rowon_n[12] 0.14fF
C445 a_1957_14202# a_2275_14202# 0.19fF
C446 a_2475_14202# a_2874_14178# 0.41fF
C447 m2_29844_946# col_n[27] 0.48fF
C448 a_32386_8194# vcm 0.24fF
C449 a_28978_15182# rowoff_n[13] 0.44fF
C450 a_2275_10186# col_n[0] 0.17fF
C451 a_2275_2154# a_15926_2130# 0.17fF
C452 a_23046_17190# vcm 0.89fF
C453 a_10998_2130# ctop 4.93fF
C454 a_19942_7150# VDD 0.29fF
C455 a_30986_7150# rowoff_n[5] 0.42fF
C456 a_20946_7150# a_21038_7150# 0.45fF
C457 a_25966_2130# vcm 0.18fF
C458 a_27062_17190# a_27062_16186# 0.84fF
C459 a_2475_16210# a_18026_16186# 0.68fF
C460 a_13310_11206# vcm 0.24fF
C461 a_11398_1488# VDD 0.17fF
C462 a_19030_8154# rowon_n[6] 0.45fF
C463 a_2275_4162# a_30986_4138# 0.17fF
C464 a_26058_6146# ctop 4.91fF
C465 a_35002_11166# VDD 0.36fF
C466 a_2475_17214# col[4] 0.22fF
C467 m3_26964_1078# m3_27968_1078# 0.21fF
C468 col_n[16] rowoff_n[0] 0.22fF
C469 col_n[19] rowoff_n[3] 0.20fF
C470 col_n[22] rowoff_n[6] 0.18fF
C471 col_n[25] rowoff_n[9] 0.16fF
C472 col_n[20] rowoff_n[4] 0.19fF
C473 col_n[23] rowoff_n[7] 0.17fF
C474 col_n[17] rowoff_n[1] 0.21fF
C475 col_n[24] rowoff_n[8] 0.16fF
C476 col_n[21] rowoff_n[5] 0.19fF
C477 a_23350_1166# col_n[20] 0.11fF
C478 col_n[18] rowoff_n[2] 0.21fF
C479 a_2475_6170# col[9] 0.22fF
C480 a_6982_12170# col_n[4] 0.34fF
C481 a_33390_13214# col_n[30] 0.11fF
C482 m2_1732_1950# vcm 1.11fF
C483 a_2275_13198# a_8990_13174# 0.71fF
C484 a_6890_5142# vcm 0.18fF
C485 a_28370_15222# vcm 0.24fF
C486 a_2475_18218# a_33998_18194# 0.41fF
C487 a_2275_12194# col_n[16] 0.17fF
C488 a_30074_17190# row_n[15] 0.43fF
C489 a_2275_1150# col_n[21] 0.17fF
C490 a_6982_9158# ctop 4.91fF
C491 a_15926_14178# VDD 0.29fF
C492 a_6890_2130# rowon_n[0] 0.14fF
C493 a_2275_15206# a_24050_15182# 0.71fF
C494 a_27062_11166# col[24] 0.38fF
C495 a_21950_9158# vcm 0.18fF
C496 a_2275_9182# col[6] 0.17fF
C497 a_16930_16186# rowoff_n[14] 0.58fF
C498 col[26] rowoff_n[14] 0.17fF
C499 a_9294_18234# vcm 0.25fF
C500 a_20034_1126# m2_20808_946# 0.86fF
C501 col_n[9] rowoff_n[10] 0.27fF
C502 a_29070_16186# m2_29268_16434# 0.19fF
C503 a_22042_13174# ctop 4.91fF
C504 a_30986_18194# VDD 0.50fF
C505 a_2475_8178# col[26] 0.22fF
C506 a_2275_12194# a_14314_12210# 0.15fF
C507 a_2475_12194# a_16930_12170# 0.41fF
C508 a_22346_11206# col_n[19] 0.11fF
C509 a_17022_15182# rowon_n[13] 0.45fF
C510 m2_30848_18014# m2_31276_18442# 0.19fF
C511 a_33086_3134# VDD 1.34fF
C512 a_27062_5142# a_28066_5142# 0.86fF
C513 a_27062_5142# rowon_n[3] 0.45fF
C514 a_6890_18194# m2_6752_18014# 0.34fF
C515 a_2275_9182# a_7894_9158# 0.17fF
C516 a_2475_18218# m2_16792_18014# 0.62fF
C517 a_2475_14202# a_31990_14178# 0.41fF
C518 a_2275_14202# a_29374_14218# 0.15fF
C519 a_16930_14178# a_17022_14178# 0.45fF
C520 a_1957_3158# rowoff_n[1] 0.14fF
C521 vcm col_n[23] 3.22fF
C522 VDD col_n[26] 9.99fF
C523 col[10] rowoff_n[15] 0.28fF
C524 a_2275_11190# col[23] 0.17fF
C525 a_17934_16186# vcm 0.18fF
C526 a_16018_9158# col[13] 0.38fF
C527 a_14010_6146# VDD 3.30fF
C528 a_4974_5142# row_n[3] 0.43fF
C529 a_18026_7150# a_18026_6146# 0.84fF
C530 a_20034_14178# m2_20232_14426# 0.19fF
C531 a_4882_9158# rowon_n[7] 0.14fF
C532 a_2966_15182# VDD 4.45fF
C533 a_2275_11190# a_22954_11166# 0.17fF
C534 a_31078_5142# col_n[28] 0.34fF
C535 a_20034_1126# vcm 0.89fF
C536 a_17022_2130# m2_17220_2378# 0.19fF
C537 a_4882_17190# rowoff_n[15] 0.72fF
C538 a_11302_9198# col_n[8] 0.11fF
C539 m2_10768_18014# VDD 4.49fF
C540 a_2874_6146# rowoff_n[4] 0.74fF
C541 a_29070_10162# VDD 1.75fF
C542 a_2475_8178# a_15014_8154# 0.68fF
C543 a_7986_8154# a_8990_8154# 0.86fF
C544 a_35094_5142# vcm 0.15fF
C545 a_12002_4138# rowoff_n[2] 2.18fF
C546 a_29070_12170# rowoff_n[10] 1.35fF
C547 a_31990_18194# a_32082_18194# 0.11fF
C548 a_26970_1126# a_27062_1126# 0.11fF
C549 a_25054_12170# rowon_n[10] 0.45fF
C550 a_2475_4162# col[3] 0.22fF
C551 a_2275_5166# a_5978_5142# 0.71fF
C552 a_10998_12170# m2_11196_12418# 0.19fF
C553 a_4974_7150# col[2] 0.38fF
C554 a_9994_13174# VDD 3.71fF
C555 a_33086_11166# a_33086_10162# 0.84fF
C556 a_2475_10186# a_30074_10162# 0.68fF
C557 a_3878_9158# rowoff_n[7] 0.73fF
C558 a_21038_2130# rowoff_n[0] 1.74fF
C559 a_20034_3134# col_n[17] 0.34fF
C560 a_2275_10186# col_n[10] 0.17fF
C561 a_16018_8154# vcm 0.89fF
C562 a_30074_15182# col_n[27] 0.34fF
C563 m2_34864_1950# m2_34864_946# 0.84fF
C564 a_30074_8154# m2_30272_8402# 0.19fF
C565 a_35398_8194# VDD 0.12fF
C566 a_2275_7174# a_21038_7150# 0.71fF
C567 a_13006_2130# row_n[0] 0.43fF
C568 a_25054_17190# VDD 2.16fF
C569 a_23046_12170# a_24050_12170# 0.86fF
C570 a_2275_7174# col[0] 0.16fF
C571 a_12914_6146# rowon_n[4] 0.14fF
C572 a_6282_2170# vcm 0.24fF
C573 a_31078_12170# vcm 0.89fF
C574 a_27974_2130# VDD 0.29fF
C575 a_2475_17214# col[15] 0.22fF
C576 col_n[28] rowoff_n[1] 0.14fF
C577 col_n[31] rowoff_n[4] 0.11fF
C578 col_n[27] rowoff_n[0] 0.14fF
C579 col_n[29] rowoff_n[2] 0.13fF
C580 col_n[30] rowoff_n[3] 0.12fF
C581 a_1957_10186# m2_1732_9982# 0.33fF
C582 a_2475_4162# a_13918_4138# 0.41fF
C583 a_2275_4162# a_11302_4178# 0.15fF
C584 a_7894_4138# a_7986_4138# 0.45fF
C585 a_2475_6170# col[20] 0.22fF
C586 m3_1864_6098# m3_1864_5094# 0.20fF
C587 a_25966_18194# m2_25828_18014# 0.34fF
C588 a_14010_14178# a_14010_13174# 0.84fF
C589 a_3970_17190# col[1] 0.38fF
C590 a_13918_10162# rowoff_n[8] 0.61fF
C591 a_21342_6186# vcm 0.24fF
C592 a_2275_12194# col_n[27] 0.17fF
C593 a_17022_13174# rowoff_n[11] 1.94fF
C594 a_2275_1150# a_4882_1126# 0.17fF
C595 a_21038_6146# m2_21236_6394# 0.19fF
C596 a_12002_15182# vcm 0.89fF
C597 a_8898_5142# VDD 0.29fF
C598 a_19030_13174# col_n[16] 0.34fF
C599 a_2475_6170# a_28978_6146# 0.41fF
C600 a_2275_6170# a_26362_6186# 0.15fF
C601 a_33086_9158# rowon_n[7] 0.45fF
C602 a_22954_8154# rowoff_n[6] 0.51fF
C603 a_2275_9182# col[17] 0.17fF
C604 a_3970_15182# a_4974_15182# 0.86fF
C605 a_2475_15206# a_6982_15182# 0.68fF
C606 a_3878_9158# vcm 0.18fF
C607 col_n[20] rowoff_n[10] 0.19fF
C608 a_33086_17190# rowoff_n[15] 1.15fF
C609 a_31990_6146# rowoff_n[4] 0.41fF
C610 a_2275_3158# a_19942_3134# 0.17fF
C611 a_15014_4138# ctop 4.91fF
C612 m3_20940_1078# ctop 0.21fF
C613 a_23958_9158# VDD 0.29fF
C614 a_10998_9158# row_n[7] 0.43fF
C615 a_22954_8154# a_23046_8154# 0.45fF
C616 a_10906_13174# rowon_n[11] 0.14fF
C617 a_29982_4138# vcm 0.18fF
C618 a_20946_3134# rowon_n[1] 0.14fF
C619 a_2475_17214# a_22042_17190# 0.68fF
C620 m2_12776_18014# m2_13780_18014# 0.86fF
C621 a_12002_4138# m2_12200_4386# 0.19fF
C622 a_17326_13214# vcm 0.24fF
C623 a_2275_5166# a_35002_5142# 0.17fF
C624 a_30074_8154# ctop 4.91fF
C625 a_4882_12170# VDD 0.29fF
C626 a_7986_11166# col_n[5] 0.34fF
C627 VDD row_n[13] 4.64fF
C628 col_n[2] rowon_n[15] 0.17fF
C629 sample rowon_n[13] 0.10fF
C630 vcm rowon_n[14] 0.91fF
C631 col_n[0] row_n[14] 0.37fF
C632 col_n[1] row_n[15] 0.37fF
C633 col[21] rowoff_n[15] 0.21fF
C634 a_2275_14202# a_13006_14178# 0.71fF
C635 col_n[4] rowoff_n[11] 0.31fF
C636 a_10906_7150# vcm 0.18fF
C637 a_4974_14178# rowoff_n[12] 2.52fF
C638 a_2475_2154# a_27062_2130# 0.68fF
C639 a_14010_2130# a_15014_2130# 0.86fF
C640 a_32386_17230# vcm 0.24fF
C641 m2_34864_17010# m3_34996_17142# 4.42fF
C642 a_31078_16186# rowon_n[14] 0.45fF
C643 a_10998_11166# ctop 4.91fF
C644 a_2275_8178# col_n[4] 0.17fF
C645 a_19942_16186# VDD 0.29fF
C646 a_2275_11190# a_3270_11206# 0.15fF
C647 a_2475_11190# a_5886_11166# 0.41fF
C648 a_1957_1150# vcm 0.16fF
C649 a_28066_10162# col[25] 0.38fF
C650 m2_10768_18014# col_n[8] 0.32fF
C651 a_2275_16210# a_28066_16186# 0.71fF
C652 a_2874_2130# m2_2736_1950# 0.34fF
C653 a_25966_11166# vcm 0.18fF
C654 a_8990_16186# row_n[14] 0.43fF
C655 a_22042_1126# VDD 0.11fF
C656 a_4974_4138# a_4974_3134# 0.84fF
C657 a_2275_5166# ctop 0.14fF
C658 a_22042_17190# m2_21812_18014# 0.84fF
C659 a_26058_15182# ctop 4.91fF
C660 a_19030_6146# row_n[4] 0.43fF
C661 a_18938_10162# rowon_n[8] 0.14fF
C662 a_2275_13198# a_18330_13214# 0.15fF
C663 a_2475_13198# a_20946_13174# 0.41fF
C664 a_23350_10202# col_n[20] 0.11fF
C665 a_2475_15206# col[9] 0.22fF
C666 a_2475_4162# col[14] 0.22fF
C667 m2_13780_946# vcm 0.71fF
C668 a_2275_1150# a_33086_1126# 0.14fF
C669 a_6890_14178# vcm 0.18fF
C670 a_2874_4138# VDD 0.29fF
C671 a_29070_6146# a_30074_6146# 0.86fF
C672 a_2275_10186# a_11910_10162# 0.17fF
C673 a_2275_10186# col_n[21] 0.17fF
C674 a_2966_2130# rowoff_n[0] 0.11fF
C675 a_18938_15182# a_19030_15182# 0.45fF
C676 a_2275_15206# a_33390_15222# 0.15fF
C677 a_17022_8154# col[14] 0.38fF
C678 m2_34864_12994# VDD 1.58fF
C679 a_5978_4138# rowon_n[2] 0.45fF
C680 a_21950_18194# vcm 0.18fF
C681 a_18026_8154# VDD 2.89fF
C682 a_2275_7174# col[11] 0.17fF
C683 a_2966_15182# m2_3164_15430# 0.19fF
C684 a_2275_7174# a_2966_7150# 0.67fF
C685 a_2475_7174# a_3970_7150# 0.68fF
C686 a_20034_8154# a_20034_7150# 0.84fF
C687 a_32082_4138# col_n[29] 0.34fF
C688 a_2275_12194# a_26970_12170# 0.17fF
C689 a_24050_3134# vcm 0.89fF
C690 a_2475_17214# col[26] 0.22fF
C691 rowon_n[8] rowoff_n[8] 20.66fF
C692 a_12306_8194# col_n[9] 0.11fF
C693 a_2475_6170# col[31] 0.22fF
C694 a_3970_5142# rowoff_n[3] 2.57fF
C695 a_17022_13174# row_n[11] 0.43fF
C696 a_33086_12170# VDD 1.34fF
C697 m3_22948_18146# m3_23952_18146# 0.21fF
C698 a_16930_17190# rowon_n[15] 0.14fF
C699 a_2475_9182# a_19030_9158# 0.68fF
C700 a_9994_9158# a_10998_9158# 0.86fF
C701 a_13006_3134# rowoff_n[1] 2.13fF
C702 a_27062_3134# row_n[1] 0.43fF
C703 a_4974_6146# vcm 0.89fF
C704 a_26970_7150# rowon_n[5] 0.14fF
C705 a_33998_14178# rowoff_n[12] 0.39fF
C706 a_28978_2130# a_29070_2130# 0.45fF
C707 m2_34864_13998# m3_34996_14130# 4.42fF
C708 a_5978_6146# col[3] 0.38fF
C709 a_2275_6170# a_9994_6146# 0.71fF
C710 a_2275_9182# col[28] 0.17fF
C711 a_14010_15182# VDD 3.30fF
C712 a_2475_11190# a_34090_11166# 0.68fF
C713 a_21038_2130# col_n[18] 0.34fF
C714 a_29374_1166# vcm 0.25fF
C715 col_n[31] rowoff_n[10] 0.11fF
C716 a_31078_14178# col_n[28] 0.34fF
C717 a_3970_11166# rowon_n[9] 0.45fF
C718 a_20034_10162# vcm 0.89fF
C719 a_11302_18234# col_n[8] 0.11fF
C720 m3_16924_18146# ctop 0.21fF
C721 a_2275_8178# a_25054_8154# 0.71fF
C722 a_25054_13174# a_26058_13174# 0.86fF
C723 a_10298_4178# vcm 0.24fF
C724 a_2275_3158# rowon_n[1] 1.99fF
C725 a_2874_17190# a_2966_17190# 0.45fF
C726 a_5886_11166# rowoff_n[9] 0.70fF
C727 a_35094_14178# vcm 0.15fF
C728 a_31990_4138# VDD 0.29fF
C729 col_n[11] rowon_n[14] 0.17fF
C730 col_n[9] rowon_n[13] 0.17fF
C731 col_n[1] rowon_n[9] 0.17fF
C732 col_n[4] row_n[11] 0.37fF
C733 col_n[0] rowon_n[8] 0.17fF
C734 col_n[12] row_n[15] 0.37fF
C735 col_n[10] row_n[14] 0.37fF
C736 col_n[8] row_n[13] 0.37fF
C737 col_n[5] rowon_n[11] 0.17fF
C738 sample row_n[8] 0.92fF
C739 VDD rowon_n[7] 4.61fF
C740 col_n[13] rowon_n[15] 0.17fF
C741 col_n[2] row_n[10] 0.37fF
C742 col_n[6] row_n[12] 0.37fF
C743 vcm row_n[9] 1.08fF
C744 a_2475_5166# a_17934_5142# 0.41fF
C745 a_2275_5166# a_15318_5182# 0.15fF
C746 col_n[3] rowon_n[10] 0.17fF
C747 a_9902_5142# a_9994_5142# 0.45fF
C748 col_n[7] rowon_n[12] 0.17fF
C749 sample_n rowoff_n[15] 0.55fF
C750 a_2475_13198# col[3] 0.22fF
C751 a_2275_18218# a_13918_18194# 0.17fF
C752 a_2475_2154# col[8] 0.22fF
C753 a_25054_10162# row_n[8] 0.43fF
C754 a_14922_9158# rowoff_n[7] 0.60fF
C755 a_4974_16186# col[2] 0.38fF
C756 col_n[15] rowoff_n[11] 0.23fF
C757 a_24962_14178# rowon_n[12] 0.14fF
C758 a_16018_15182# a_16018_14178# 0.84fF
C759 a_25358_8194# vcm 0.24fF
C760 a_21950_15182# rowoff_n[13] 0.52fF
C761 a_20034_12170# col_n[17] 0.34fF
C762 a_35002_4138# rowon_n[2] 0.14fF
C763 a_2275_2154# a_8898_2130# 0.17fF
C764 a_16018_17190# vcm 0.89fF
C765 a_3970_2130# ctop 4.87fF
C766 a_2275_8178# col_n[15] 0.17fF
C767 m2_23820_18014# m3_23952_18146# 4.41fF
C768 a_12914_7150# VDD 0.29fF
C769 a_23958_7150# rowoff_n[5] 0.50fF
C770 a_26058_15182# m2_26256_15430# 0.19fF
C771 a_2275_7174# a_30378_7190# 0.15fF
C772 a_2475_7174# a_32994_7150# 0.41fF
C773 a_35398_17230# VDD 0.12fF
C774 a_18938_2130# vcm 0.18fF
C775 a_2275_16210# col[0] 0.16fF
C776 a_5978_16186# a_6982_16186# 0.86fF
C777 a_2475_16210# a_10998_16186# 0.68fF
C778 a_2275_5166# col[5] 0.17fF
C779 a_6282_11206# vcm 0.24fF
C780 a_32994_5142# rowoff_n[3] 0.40fF
C781 a_4370_1488# VDD 0.18fF
C782 a_12002_8154# rowon_n[6] 0.45fF
C783 a_2275_4162# a_23958_4138# 0.17fF
C784 a_19030_6146# ctop 4.91fF
C785 a_27974_11166# VDD 0.29fF
C786 m3_12908_1078# m3_13912_1078# 0.21fF
C787 a_24962_9158# a_25054_9158# 0.45fF
C788 col_n[0] rowoff_n[12] 0.34fF
C789 a_2475_15206# col[20] 0.22fF
C790 a_2475_4162# col[25] 0.22fF
C791 m2_13780_946# col_n[11] 0.45fF
C792 a_1957_13198# a_2161_13198# 0.11fF
C793 a_2475_13198# a_2275_13198# 2.96fF
C794 a_33998_6146# vcm 0.18fF
C795 a_21342_15222# vcm 0.24fF
C796 m2_34864_10986# m3_34996_11118# 4.42fF
C797 a_2475_18218# a_26970_18194# 0.41fF
C798 a_17022_13174# m2_17220_13422# 0.19fF
C799 a_8990_10162# col_n[6] 0.34fF
C800 a_34090_10162# ctop 4.80fF
C801 a_23046_17190# row_n[15] 0.43fF
C802 a_8898_14178# VDD 0.29fF
C803 a_33086_7150# row_n[5] 0.43fF
C804 a_2275_15206# a_17022_15182# 0.71fF
C805 a_32994_11166# rowon_n[9] 0.14fF
C806 a_14922_9158# vcm 0.18fF
C807 a_9902_16186# rowoff_n[14] 0.66fF
C808 a_2275_7174# col[22] 0.17fF
C809 a_2475_3158# a_31078_3134# 0.68fF
C810 a_16018_3134# a_17022_3134# 0.86fF
C811 a_3878_18194# vcm 0.18fF
C812 a_15014_13174# ctop 4.91fF
C813 a_23958_18194# VDD 0.50fF
C814 a_2275_12194# a_7286_12210# 0.15fF
C815 a_2475_12194# a_9902_12170# 0.41fF
C816 a_29070_9158# col[26] 0.38fF
C817 a_5886_12170# a_5978_12170# 0.45fF
C818 a_34090_11166# rowoff_n[9] 1.10fF
C819 a_2275_17214# a_32082_17190# 0.71fF
C820 a_9994_15182# rowon_n[13] 0.45fF
C821 m2_23820_18014# m2_24248_18442# 0.19fF
C822 a_29982_13174# vcm 0.18fF
C823 a_26058_3134# VDD 2.06fF
C824 a_7986_11166# m2_8184_11414# 0.19fF
C825 a_6982_5142# a_6982_4138# 0.84fF
C826 a_20034_5142# rowon_n[3] 0.45fF
C827 a_30074_17190# ctop 4.93fF
C828 a_24354_9198# col_n[21] 0.11fF
C829 a_2475_18218# m2_2736_18014# 0.59fF
C830 a_2275_14202# a_22346_14218# 0.15fF
C831 a_2475_14202# a_24962_14178# 0.41fF
C832 a_27062_7150# m2_27260_7398# 0.19fF
C833 a_10906_16186# vcm 0.18fF
C834 a_6982_6146# VDD 4.02fF
C835 a_31078_7150# a_32082_7150# 0.86fF
C836 rowon_n[10] rowoff_n[10] 20.66fF
C837 a_31078_14178# row_n[12] 0.43fF
C838 a_2275_11190# a_15926_11166# 0.17fF
C839 a_2275_17214# col_n[4] 0.17fF
C840 a_13006_1126# vcm 0.15fF
C841 a_20946_16186# a_21038_16186# 0.45fF
C842 a_18026_7150# col[15] 0.38fF
C843 a_2275_6170# col_n[9] 0.17fF
C844 m2_1732_13998# m2_1732_12994# 0.84fF
C845 a_1957_10186# vcm 0.16fF
C846 a_6982_2130# m2_6752_946# 0.84fF
C847 a_33086_3134# col_n[30] 0.34fF
C848 a_22042_10162# VDD 2.47fF
C849 a_2475_8178# a_7986_8154# 0.68fF
C850 a_22042_9158# a_22042_8154# 0.84fF
C851 a_2275_14202# ctop 0.14fF
C852 a_2275_13198# a_30986_13174# 0.17fF
C853 m2_25828_18014# col[23] 0.39fF
C854 a_13310_7190# col_n[10] 0.11fF
C855 a_28066_5142# vcm 0.89fF
C856 a_4974_4138# rowoff_n[2] 2.52fF
C857 a_22042_12170# rowoff_n[10] 1.69fF
C858 a_2275_18218# m2_33860_18014# 0.51fF
C859 col_n[10] rowon_n[8] 0.17fF
C860 col_n[1] row_n[4] 0.37fF
C861 col_n[17] row_n[12] 0.37fF
C862 col_n[16] rowon_n[11] 0.17fF
C863 col_n[0] row_n[3] 0.37fF
C864 col_n[8] rowon_n[7] 0.17fF
C865 col_n[24] rowon_n[15] 0.17fF
C866 vcm rowon_n[3] 0.91fF
C867 col_n[6] rowon_n[6] 0.17fF
C868 col_n[13] row_n[10] 0.37fF
C869 col_n[22] rowon_n[14] 0.17fF
C870 sample rowon_n[2] 0.10fF
C871 col_n[4] rowon_n[5] 0.17fF
C872 col_n[11] row_n[9] 0.37fF
C873 col_n[20] rowon_n[13] 0.17fF
C874 col_n[2] rowon_n[4] 0.17fF
C875 col_n[9] row_n[8] 0.37fF
C876 col_n[15] row_n[11] 0.37fF
C877 col_n[14] rowon_n[10] 0.17fF
C878 col_n[12] rowon_n[9] 0.17fF
C879 VDD row_n[2] 4.64fF
C880 col_n[18] rowon_n[12] 0.17fF
C881 col_n[19] row_n[13] 0.37fF
C882 col_n[3] row_n[5] 0.37fF
C883 col_n[21] row_n[14] 0.37fF
C884 col_n[5] row_n[6] 0.37fF
C885 col_n[23] row_n[15] 0.37fF
C886 col_n[7] row_n[7] 0.37fF
C887 a_18026_5142# m2_18224_5390# 0.19fF
C888 m2_34864_7974# m3_34996_8106# 4.47fF
C889 a_2475_13198# col[14] 0.22fF
C890 a_18026_12170# rowon_n[10] 0.45fF
C891 a_2475_2154# col[19] 0.22fF
C892 col_n[26] rowoff_n[11] 0.15fF
C893 a_2874_13174# VDD 0.29fF
C894 a_2475_10186# a_23046_10162# 0.68fF
C895 a_12002_10162# a_13006_10162# 0.86fF
C896 a_28066_2130# rowon_n[0] 0.45fF
C897 a_14010_2130# rowoff_n[0] 2.08fF
C898 m2_34864_13998# vcm 0.74fF
C899 a_2275_8178# col_n[26] 0.17fF
C900 a_8990_8154# vcm 0.89fF
C901 a_3878_15182# rowoff_n[13] 0.73fF
C902 a_6982_5142# col[4] 0.38fF
C903 a_30986_3134# a_31078_3134# 0.45fF
C904 a_17022_17190# col[14] 0.38fF
C905 a_2275_7174# a_14010_7150# 0.71fF
C906 a_5978_2130# row_n[0] 0.43fF
C907 a_18026_17190# VDD 2.89fF
C908 a_2275_16210# col[11] 0.17fF
C909 a_5886_6146# rowon_n[4] 0.14fF
C910 a_32082_13174# col_n[29] 0.34fF
C911 a_2275_5166# col[16] 0.17fF
C912 a_33390_3174# vcm 0.24fF
C913 a_8990_3134# m2_9188_3382# 0.19fF
C914 a_24050_12170# vcm 0.89fF
C915 a_12306_17230# col_n[9] 0.11fF
C916 a_20946_2130# VDD 0.29fF
C917 col_n[10] rowoff_n[12] 0.27fF
C918 a_2475_15206# col[31] 0.22fF
C919 a_2475_4162# a_6890_4138# 0.41fF
C920 a_2275_4162# a_4274_4178# 0.15fF
C921 m2_30848_946# m3_30980_1078# 4.41fF
C922 m3_1864_13126# m3_1864_12122# 0.20fF
C923 a_2275_9182# a_29070_9158# 0.71fF
C924 a_27062_14178# a_28066_14178# 0.86fF
C925 a_6890_10162# rowoff_n[8] 0.69fF
C926 a_14314_6186# vcm 0.24fF
C927 a_9994_13174# rowoff_n[11] 2.28fF
C928 a_4974_15182# vcm 0.89fF
C929 a_2475_6170# a_21950_6146# 0.41fF
C930 a_2275_6170# a_19334_6186# 0.15fF
C931 a_11910_6146# a_12002_6146# 0.45fF
C932 a_2966_13174# m2_1732_12994# 0.86fF
C933 a_26058_9158# rowon_n[7] 0.45fF
C934 a_5978_15182# col[3] 0.38fF
C935 a_15926_8154# rowoff_n[6] 0.59fF
C936 a_18026_16186# a_18026_15182# 0.84fF
C937 m2_1732_4962# sample 0.31fF
C938 a_21038_11166# col_n[18] 0.34fF
C939 a_29374_10202# vcm 0.24fF
C940 a_26058_17190# rowoff_n[15] 1.50fF
C941 m2_1732_16006# VDD 5.46fF
C942 a_24962_6146# rowoff_n[4] 0.49fF
C943 a_2275_3158# a_12914_3134# 0.17fF
C944 a_7986_4138# ctop 4.91fF
C945 a_2475_1150# m2_5748_946# 0.62fF
C946 a_3970_9158# row_n[7] 0.43fF
C947 m3_1864_5094# ctop 0.22fF
C948 a_16930_9158# VDD 0.29fF
C949 ctop rowoff_n[6] 0.28fF
C950 row_n[1] rowoff_n[1] 0.64fF
C951 a_2275_8178# a_35398_8194# 0.15fF
C952 a_2275_16210# m2_34864_16006# 0.51fF
C953 a_2275_4162# col_n[3] 0.17fF
C954 a_22954_4138# vcm 0.18fF
C955 a_13918_3134# rowon_n[1] 0.14fF
C956 a_33998_4138# rowoff_n[2] 0.39fF
C957 a_2475_17214# a_15014_17190# 0.68fF
C958 a_7986_17190# a_8990_17190# 0.86fF
C959 m2_5748_18014# m2_6752_18014# 0.86fF
C960 a_10298_13214# vcm 0.24fF
C961 m2_34864_4962# m3_34996_5094# 4.42fF
C962 a_2275_5166# a_27974_5142# 0.17fF
C963 a_23046_8154# ctop 4.91fF
C964 a_31990_13174# VDD 0.29fF
C965 a_26970_10162# a_27062_10162# 0.45fF
C966 a_2275_14202# a_5978_14178# 0.71fF
C967 a_2475_11190# col[8] 0.22fF
C968 a_2475_2154# a_20034_2130# 0.68fF
C969 a_28066_3134# a_28066_2130# 0.84fF
C970 a_25358_17230# vcm 0.24fF
C971 a_9994_9158# col_n[7] 0.34fF
C972 a_24050_16186# rowon_n[14] 0.45fF
C973 a_35002_15182# m2_34864_15002# 0.33fF
C974 a_3970_11166# ctop 4.91fF
C975 a_2275_17214# col_n[15] 0.17fF
C976 a_12914_16186# VDD 0.29fF
C977 a_2275_6170# col_n[20] 0.17fF
C978 a_34090_6146# rowon_n[4] 0.45fF
C979 a_2275_18218# vcm 8.30fF
C980 a_2275_16210# a_21038_16186# 0.71fF
C981 a_18938_11166# vcm 0.18fF
C982 a_15014_1126# VDD 0.13fF
C983 a_2475_16210# row_n[14] 0.48fF
C984 a_2275_14202# col[5] 0.17fF
C985 a_18026_4138# a_19030_4138# 0.86fF
C986 a_2275_3158# col[10] 0.17fF
C987 a_34394_10202# col_n[31] 0.11fF
C988 a_30074_8154# col[27] 0.38fF
C989 a_19030_15182# ctop 4.91fF
C990 a_12002_6146# row_n[4] 0.43fF
C991 a_11910_10162# rowon_n[8] 0.14fF
C992 a_2475_13198# a_13918_13174# 0.41fF
C993 a_2275_13198# a_11302_13214# 0.15fF
C994 a_7894_13174# a_7986_13174# 0.45fF
C995 col_n[8] row_n[2] 0.37fF
C996 col_n[6] row_n[1] 0.37fF
C997 col_n[25] rowon_n[10] 0.17fF
C998 col_n[4] row_n[0] 0.37fF
C999 col_n[23] rowon_n[9] 0.17fF
C1000 col_n[21] rowon_n[8] 0.17fF
C1001 col_n[28] row_n[12] 0.37fF
C1002 col_n[27] rowon_n[11] 0.17fF
C1003 col_n[19] rowon_n[7] 0.17fF
C1004 col_n[17] rowon_n[6] 0.17fF
C1005 col_n[30] row_n[13] 0.37fF
C1006 col_n[12] row_n[4] 0.37fF
C1007 col_n[10] row_n[3] 0.37fF
C1008 col_n[29] rowon_n[12] 0.17fF
C1009 col_n[5] rowon_n[0] 0.17fF
C1010 col_n[14] row_n[5] 0.37fF
C1011 col_n[7] rowon_n[1] 0.17fF
C1012 VDD en_bit_n[0] 0.34fF
C1013 col_n[16] row_n[6] 0.37fF
C1014 col_n[9] rowon_n[2] 0.17fF
C1015 col_n[18] row_n[7] 0.37fF
C1016 col_n[11] rowon_n[3] 0.17fF
C1017 col_n[26] row_n[11] 0.37fF
C1018 col_n[20] row_n[8] 0.37fF
C1019 col_n[13] rowon_n[4] 0.17fF
C1020 col_n[31] rowon_n[13] 0.17fF
C1021 col_n[22] row_n[9] 0.37fF
C1022 col_n[15] rowon_n[5] 0.17fF
C1023 col_n[24] row_n[10] 0.37fF
C1024 a_2475_13198# col[25] 0.22fF
C1025 a_2475_2154# col[30] 0.22fF
C1026 a_2275_1150# a_26058_1126# 0.14fF
C1027 a_33998_15182# vcm 0.18fF
C1028 a_30074_5142# VDD 1.65fF
C1029 a_8990_6146# a_8990_5142# 0.84fF
C1030 a_25358_8194# col_n[22] 0.11fF
C1031 a_2275_10186# a_4882_10162# 0.17fF
C1032 a_2966_10162# a_3970_10162# 0.86fF
C1033 a_2475_15206# a_28978_15182# 0.41fF
C1034 a_2275_15206# a_26362_15222# 0.15fF
C1035 a_14922_18194# vcm 0.18fF
C1036 a_2275_16210# col[22] 0.17fF
C1037 a_10998_8154# VDD 3.61fF
C1038 a_33086_8154# a_34090_8154# 0.86fF
C1039 a_32082_16186# m2_32280_16434# 0.19fF
C1040 a_2275_5166# col[27] 0.17fF
C1041 a_32082_13174# rowon_n[11] 0.45fF
C1042 m2_23820_946# col_n[21] 0.45fF
C1043 a_2275_12194# a_19942_12170# 0.17fF
C1044 a_19030_6146# col[16] 0.38fF
C1045 a_17022_3134# vcm 0.89fF
C1046 a_22954_17190# a_23046_17190# 0.45fF
C1047 col_n[21] rowoff_n[12] 0.19fF
C1048 a_2275_2154# VDD 3.18fF
C1049 a_34090_2130# col_n[31] 0.46fF
C1050 a_9994_13174# row_n[11] 0.43fF
C1051 a_26058_12170# VDD 2.06fF
C1052 m3_8892_18146# m3_9896_18146# 0.21fF
C1053 a_9902_17190# rowon_n[15] 0.14fF
C1054 a_24050_10162# a_24050_9158# 0.84fF
C1055 a_2475_9182# a_12002_9158# 0.68fF
C1056 a_14314_6186# col_n[11] 0.11fF
C1057 a_2275_14202# a_35002_14178# 0.17fF
C1058 a_5978_3134# rowoff_n[1] 2.47fF
C1059 a_20034_3134# row_n[1] 0.43fF
C1060 a_24354_18234# col_n[21] 0.11fF
C1061 a_19942_7150# rowon_n[5] 0.14fF
C1062 a_32082_7150# vcm 0.89fF
C1063 a_26970_14178# rowoff_n[12] 0.47fF
C1064 a_2475_6170# a_3878_6146# 0.41fF
C1065 a_2275_6170# a_2874_6146# 0.17fF
C1066 a_23046_14178# m2_23244_14426# 0.19fF
C1067 a_2475_9182# col[2] 0.22fF
C1068 a_6982_15182# VDD 4.02fF
C1069 m2_34864_12994# rowoff_n[11] 1.01fF
C1070 a_14010_11166# a_15014_11166# 0.86fF
C1071 a_2475_11190# a_27062_11166# 0.68fF
C1072 col_n[5] rowoff_n[13] 0.30fF
C1073 a_22346_1166# vcm 0.25fF
C1074 a_7986_4138# col[5] 0.38fF
C1075 a_13006_10162# vcm 0.89fF
C1076 col[8] rowoff_n[9] 0.29fF
C1077 col[7] rowoff_n[8] 0.30fF
C1078 col[6] rowoff_n[7] 0.31fF
C1079 col[5] rowoff_n[6] 0.31fF
C1080 col[0] rowoff_n[1] 0.34fF
C1081 col[1] rowoff_n[2] 0.34fF
C1082 col[2] rowoff_n[3] 0.33fF
C1083 col[3] rowoff_n[4] 0.33fF
C1084 col[4] rowoff_n[5] 0.32fF
C1085 a_18026_16186# col[15] 0.38fF
C1086 a_2275_15206# col_n[9] 0.17fF
C1087 a_32994_4138# a_33086_4138# 0.45fF
C1088 a_2275_4162# col_n[14] 0.17fF
C1089 a_2275_8178# a_18026_8154# 0.71fF
C1090 a_33086_12170# col_n[30] 0.34fF
C1091 a_4974_13174# a_4974_12170# 0.84fF
C1092 a_3270_4178# vcm 0.24fF
C1093 a_2275_1150# col[4] 0.17fF
C1094 a_13310_16226# col_n[10] 0.11fF
C1095 a_28066_14178# vcm 0.89fF
C1096 a_24962_4138# VDD 0.29fF
C1097 a_14010_12170# m2_14208_12418# 0.19fF
C1098 a_2475_5166# a_10906_5142# 0.41fF
C1099 a_2275_5166# a_8290_5182# 0.15fF
C1100 a_2275_18218# a_6890_18194# 0.17fF
C1101 a_2275_10186# a_33086_10162# 0.71fF
C1102 a_2475_11190# col[19] 0.22fF
C1103 a_18026_10162# row_n[8] 0.43fF
C1104 a_7894_9158# rowoff_n[7] 0.68fF
C1105 a_17934_14178# rowon_n[12] 0.14fF
C1106 a_29070_15182# a_30074_15182# 0.86fF
C1107 a_18330_8194# vcm 0.24fF
C1108 a_14922_15182# rowoff_n[13] 0.60fF
C1109 a_33086_8154# m2_33284_8402# 0.19fF
C1110 a_27974_4138# rowon_n[2] 0.14fF
C1111 a_31078_3134# ctop 4.91fF
C1112 a_8990_17190# vcm 0.89fF
C1113 a_2275_17214# col_n[26] 0.17fF
C1114 a_5886_7150# VDD 0.29fF
C1115 a_16930_7150# rowoff_n[5] 0.58fF
C1116 a_2275_6170# col_n[31] 0.17fF
C1117 a_6982_14178# col[4] 0.38fF
C1118 a_2275_7174# a_23350_7190# 0.15fF
C1119 a_2475_7174# a_25966_7150# 0.41fF
C1120 a_13918_7150# a_14010_7150# 0.45fF
C1121 a_2275_18218# col_n[11] 0.17fF
C1122 a_22042_10162# col_n[19] 0.34fF
C1123 a_11910_2130# vcm 0.18fF
C1124 a_2475_16210# a_3970_16186# 0.68fF
C1125 a_2275_16210# a_2966_16186# 0.67fF
C1126 a_20034_17190# a_20034_16186# 0.84fF
C1127 a_2275_14202# col[16] 0.17fF
C1128 a_25966_5142# rowoff_n[3] 0.48fF
C1129 a_33390_12210# vcm 0.24fF
C1130 a_2275_3158# col[21] 0.17fF
C1131 a_4974_8154# rowon_n[6] 0.45fF
C1132 a_4974_10162# m2_5172_10410# 0.19fF
C1133 a_2275_4162# a_16930_4138# 0.17fF
C1134 a_12002_6146# ctop 4.91fF
C1135 a_20946_11166# VDD 0.29fF
C1136 m3_1864_2082# m3_2868_2082# 0.21fF
C1137 m3_34996_3086# m3_34996_2082# 0.20fF
C1138 col_n[18] rowon_n[1] 0.17fF
C1139 col_n[25] row_n[5] 0.37fF
C1140 col_n[16] rowon_n[0] 0.17fF
C1141 col_n[23] row_n[4] 0.37fF
C1142 col_n[21] row_n[3] 0.37fF
C1143 col_n[19] row_n[2] 0.37fF
C1144 col_n[17] row_n[1] 0.37fF
C1145 vcm col[6] 6.66fF
C1146 col_n[15] row_n[0] 0.37fF
C1147 col_n[22] rowon_n[3] 0.17fF
C1148 col_n[29] row_n[7] 0.37fF
C1149 col_n[20] rowon_n[2] 0.17fF
C1150 col_n[27] row_n[6] 0.37fF
C1151 col_n[31] row_n[8] 0.37fF
C1152 col_n[24] rowon_n[4] 0.17fF
C1153 col_n[26] rowon_n[5] 0.17fF
C1154 col_n[3] col[3] 0.50fF
C1155 col_n[28] rowon_n[6] 0.17fF
C1156 VDD col[9] 11.20fF
C1157 col_n[30] rowon_n[7] 0.17fF
C1158 a_35002_3134# rowoff_n[1] 0.38fF
C1159 a_26970_6146# vcm 0.18fF
C1160 a_24050_6146# m2_24248_6394# 0.19fF
C1161 a_14314_15222# vcm 0.24fF
C1162 a_2475_18218# a_19942_18194# 0.41fF
C1163 a_2275_6170# a_31990_6146# 0.17fF
C1164 a_27062_10162# ctop 4.91fF
C1165 a_16018_17190# row_n[15] 0.43fF
C1166 a_28978_11166# a_29070_11166# 0.45fF
C1167 m2_1732_17010# vcm 1.11fF
C1168 a_26058_7150# row_n[5] 0.43fF
C1169 a_2275_15206# a_9994_15182# 0.71fF
C1170 a_25966_11166# rowon_n[9] 0.14fF
C1171 a_7894_9158# vcm 0.18fF
C1172 a_10998_8154# col_n[8] 0.34fF
C1173 a_2161_16210# rowoff_n[14] 0.14fF
C1174 a_2475_3158# a_24050_3134# 0.68fF
C1175 a_30074_4138# a_30074_3134# 0.84fF
C1176 a_2475_1150# m2_28840_946# 0.62fF
C1177 a_7986_13174# ctop 4.91fF
C1178 a_16930_18194# VDD 0.50fF
C1179 a_2275_13198# col_n[3] 0.17fF
C1180 a_2275_2154# col_n[8] 0.17fF
C1181 a_2275_17214# a_25054_17190# 0.71fF
C1182 a_27062_11166# rowoff_n[9] 1.45fF
C1183 a_2874_15182# rowon_n[13] 0.14fF
C1184 a_15014_4138# m2_15212_4386# 0.19fF
C1185 m2_16792_18014# m2_17220_18442# 0.19fF
C1186 a_22954_13174# vcm 0.18fF
C1187 a_19030_3134# VDD 2.78fF
C1188 a_2275_11190# m2_1732_10986# 0.27fF
C1189 a_20034_5142# a_21038_5142# 0.86fF
C1190 a_31078_7150# col[28] 0.38fF
C1191 a_13006_5142# rowon_n[3] 0.45fF
C1192 a_2275_18218# a_35094_18194# 0.14fF
C1193 a_23046_17190# ctop 4.93fF
C1194 a_9902_14178# a_9994_14178# 0.45fF
C1195 a_2275_14202# a_15318_14218# 0.15fF
C1196 a_2475_14202# a_17934_14178# 0.41fF
C1197 a_1957_3158# row_n[1] 0.29fF
C1198 m2_34864_12994# row_n[11] 0.38fF
C1199 a_2275_2154# a_30074_2130# 0.71fF
C1200 a_2475_9182# col[13] 0.22fF
C1201 a_26362_7190# col_n[23] 0.11fF
C1202 a_34090_7150# VDD 1.23fF
C1203 a_10998_7150# a_10998_6146# 0.84fF
C1204 col_n[16] rowoff_n[13] 0.22fF
C1205 m2_1732_13998# rowoff_n[12] 2.46fF
C1206 a_2275_11190# a_8898_11166# 0.17fF
C1207 a_24050_14178# row_n[12] 0.43fF
C1208 a_5978_1126# vcm 0.15fF
C1209 col[19] rowoff_n[9] 0.22fF
C1210 col[18] rowoff_n[8] 0.23fF
C1211 col[17] rowoff_n[7] 0.23fF
C1212 col[16] rowoff_n[6] 0.24fF
C1213 col[15] rowoff_n[5] 0.25fF
C1214 col[14] rowoff_n[4] 0.25fF
C1215 col[13] rowoff_n[3] 0.26fF
C1216 col[12] rowoff_n[2] 0.27fF
C1217 col[11] rowoff_n[1] 0.27fF
C1218 col[10] rowoff_n[0] 0.28fF
C1219 a_2275_15206# col_n[20] 0.17fF
C1220 a_2475_16210# a_32994_16186# 0.41fF
C1221 a_2275_16210# a_30378_16226# 0.15fF
C1222 a_2275_4162# col_n[25] 0.17fF
C1223 a_34090_4138# row_n[2] 0.43fF
C1224 a_33998_8154# rowon_n[6] 0.14fF
C1225 a_15014_10162# VDD 3.20fF
C1226 a_20034_5142# col[17] 0.38fF
C1227 a_2275_12194# col[10] 0.17fF
C1228 a_2275_13198# a_23958_13174# 0.17fF
C1229 a_2275_1150# col[15] 0.17fF
C1230 a_30074_17190# col[27] 0.38fF
C1231 a_21038_5142# vcm 0.89fF
C1232 a_24962_18194# a_25054_18194# 0.11fF
C1233 a_15014_12170# rowoff_n[10] 2.03fF
C1234 m2_22816_946# vcm 0.71fF
C1235 a_2275_18218# m2_19804_18014# 0.51fF
C1236 a_19942_1126# a_20034_1126# 0.47fF
C1237 a_10998_12170# rowon_n[10] 0.45fF
C1238 a_2475_11190# col[30] 0.22fF
C1239 a_34090_13174# m2_34864_12994# 0.86fF
C1240 vcm rowoff_n[14] 2.43fF
C1241 a_30074_14178# VDD 1.65fF
C1242 a_15318_5182# col_n[12] 0.11fF
C1243 a_26058_11166# a_26058_10162# 0.84fF
C1244 a_2475_10186# a_16018_10162# 0.68fF
C1245 a_21038_2130# rowon_n[0] 0.45fF
C1246 a_25358_17230# col_n[22] 0.11fF
C1247 a_6982_2130# rowoff_n[0] 2.42fF
C1248 col[3] rowoff_n[10] 0.33fF
C1249 a_2475_8178# vcm 1.32fF
C1250 a_31078_16186# rowoff_n[14] 1.25fF
C1251 a_2275_18218# col_n[22] 0.17fF
C1252 a_2275_7174# a_6982_7150# 0.71fF
C1253 a_10998_17190# VDD 3.61fF
C1254 a_16018_12170# a_17022_12170# 0.86fF
C1255 a_2475_12194# a_31078_12170# 0.68fF
C1256 a_2275_14202# col[27] 0.17fF
C1257 a_8990_3134# col[6] 0.38fF
C1258 a_26362_3174# vcm 0.24fF
C1259 a_32082_11166# row_n[9] 0.43fF
C1260 a_31990_15182# rowon_n[13] 0.14fF
C1261 a_19030_15182# col[16] 0.38fF
C1262 a_17022_12170# vcm 0.89fF
C1263 a_13918_2130# VDD 0.29fF
C1264 rowon_n[9] row_n[9] 21.02fF
C1265 vcm col[17] 6.66fF
C1266 col_n[31] rowon_n[2] 0.17fF
C1267 col_n[29] rowon_n[1] 0.17fF
C1268 VDD col[20] 8.48fF
C1269 col_n[27] rowon_n[0] 0.17fF
C1270 col_n[8] col[9] 6.22fF
C1271 col_n[26] row_n[0] 0.37fF
C1272 col_n[28] row_n[1] 0.37fF
C1273 col_n[30] row_n[2] 0.37fF
C1274 a_35002_5142# a_35094_5142# 0.11fF
C1275 a_2275_11190# VDD 3.18fF
C1276 a_34090_11166# col_n[31] 0.34fF
C1277 a_2275_9182# a_22042_9158# 0.71fF
C1278 m2_4744_18014# col_n[2] 0.33fF
C1279 a_4274_3174# col_n[1] 0.11fF
C1280 a_6982_14178# a_6982_13174# 0.84fF
C1281 a_14314_15222# col_n[11] 0.11fF
C1282 a_7286_6186# vcm 0.24fF
C1283 a_2874_13174# rowoff_n[11] 0.74fF
C1284 a_20034_1126# ctop 0.68fF
C1285 a_32082_16186# vcm 0.89fF
C1286 a_28978_6146# VDD 0.29fF
C1287 a_2275_6170# a_12306_6186# 0.15fF
C1288 a_2475_6170# a_14922_6146# 0.41fF
C1289 a_19030_9158# rowon_n[7] 0.45fF
C1290 a_8898_8154# rowoff_n[6] 0.67fF
C1291 a_33390_1166# vcm 0.26fF
C1292 a_31078_16186# a_32082_16186# 0.86fF
C1293 a_2475_7174# col[7] 0.22fF
C1294 a_22346_10202# vcm 0.24fF
C1295 a_19030_17190# rowoff_n[15] 1.84fF
C1296 a_7986_13174# col[5] 0.38fF
C1297 a_2275_3158# a_5886_3134# 0.17fF
C1298 a_17934_6146# rowoff_n[4] 0.57fF
C1299 m3_31984_18146# ctop 0.21fF
C1300 a_9902_9158# VDD 0.29fF
C1301 a_15926_8154# a_16018_8154# 0.45fF
C1302 a_2275_8178# a_27366_8194# 0.15fF
C1303 a_2475_8178# a_29982_8154# 0.41fF
C1304 a_2275_13198# col_n[14] 0.17fF
C1305 a_2275_2154# col_n[19] 0.17fF
C1306 a_23046_9158# col_n[20] 0.34fF
C1307 a_15926_4138# vcm 0.18fF
C1308 a_6890_3134# rowon_n[1] 0.14fF
C1309 a_26970_4138# rowoff_n[2] 0.47fF
C1310 a_2475_17214# a_7986_17190# 0.68fF
C1311 a_3270_13214# vcm 0.24fF
C1312 a_35494_4500# VDD 0.13fF
C1313 a_2275_10186# col[4] 0.17fF
C1314 a_2275_5166# a_20946_5142# 0.17fF
C1315 a_16018_8154# ctop 4.91fF
C1316 a_24962_13174# VDD 0.29fF
C1317 a_2475_9182# col[24] 0.22fF
C1318 a_30986_8154# vcm 0.18fF
C1319 a_2475_2154# a_13006_2130# 0.68fF
C1320 a_6982_2130# a_7986_2130# 0.86fF
C1321 a_18330_17230# vcm 0.24fF
C1322 col_n[27] rowoff_n[13] 0.14fF
C1323 m2_28840_18014# m3_28972_18146# 4.41fF
C1324 a_17022_16186# rowon_n[14] 0.45fF
C1325 a_2275_7174# a_34394_7190# 0.15fF
C1326 a_29070_15182# m2_29268_15430# 0.19fF
C1327 a_31078_12170# ctop 4.91fF
C1328 a_5886_16186# VDD 0.29fF
C1329 col[21] rowoff_n[0] 0.21fF
C1330 col[22] rowoff_n[1] 0.20fF
C1331 col[23] rowoff_n[2] 0.19fF
C1332 col[24] rowoff_n[3] 0.19fF
C1333 col[25] rowoff_n[4] 0.18fF
C1334 col[26] rowoff_n[5] 0.17fF
C1335 col[27] rowoff_n[6] 0.17fF
C1336 col[28] rowoff_n[7] 0.16fF
C1337 col[29] rowoff_n[8] 0.15fF
C1338 col[30] rowoff_n[9] 0.15fF
C1339 a_2275_15206# col_n[31] 0.17fF
C1340 a_30986_12170# a_31078_12170# 0.45fF
C1341 a_27062_6146# rowon_n[4] 0.45fF
C1342 a_2275_16210# a_14010_16186# 0.71fF
C1343 a_12002_7150# col_n[9] 0.34fF
C1344 a_11910_11166# vcm 0.18fF
C1345 a_7986_1126# VDD 0.14fF
C1346 a_32082_5142# a_32082_4138# 0.84fF
C1347 a_2475_4162# a_28066_4138# 0.68fF
C1348 a_2275_12194# col[21] 0.17fF
C1349 a_2275_1150# col[26] 0.17fF
C1350 a_12002_15182# ctop 4.91fF
C1351 a_4974_6146# row_n[4] 0.43fF
C1352 a_2475_13198# a_6890_13174# 0.41fF
C1353 a_2275_13198# a_4274_13214# 0.15fF
C1354 a_4882_10162# rowon_n[8] 0.14fF
C1355 a_28066_10162# rowoff_n[8] 1.40fF
C1356 a_2966_5142# vcm 0.89fF
C1357 a_31990_13174# rowoff_n[11] 0.41fF
C1358 col_n[11] rowoff_n[14] 0.26fF
C1359 a_2275_1150# a_19030_1126# 0.79fF
C1360 a_26970_15182# vcm 0.18fF
C1361 a_23046_5142# VDD 2.37fF
C1362 a_32082_6146# col[29] 0.38fF
C1363 m2_26832_946# VDD 3.70fF
C1364 a_22042_6146# a_23046_6146# 0.86fF
C1365 a_20034_13174# m2_20232_13422# 0.19fF
C1366 col[14] rowoff_n[10] 0.25fF
C1367 a_2475_15206# a_21950_15182# 0.41fF
C1368 a_2275_15206# a_19334_15222# 0.15fF
C1369 a_11910_15182# a_12002_15182# 0.45fF
C1370 a_27366_6186# col_n[24] 0.11fF
C1371 a_2275_3158# a_34090_3134# 0.71fF
C1372 a_7894_18194# vcm 0.18fF
C1373 a_18026_1126# m2_16792_946# 0.86fF
C1374 a_10998_17190# col_n[8] 0.34fF
C1375 a_3970_8154# VDD 4.33fF
C1376 a_13006_8154# a_13006_7150# 0.84fF
C1377 a_2475_5166# col[1] 0.22fF
C1378 a_25054_13174# rowon_n[11] 0.45fF
C1379 a_2275_12194# a_12914_12170# 0.17fF
C1380 a_9994_3134# vcm 0.89fF
C1381 a_2275_17214# a_35398_17230# 0.15fF
C1382 rowon_n[14] ctop 0.37fF
C1383 VDD col[31] 5.75fF
C1384 vcm col[28] 6.66fF
C1385 col_n[14] col[14] 0.50fF
C1386 a_2275_11190# col_n[8] 0.17fF
C1387 a_10998_11166# m2_11196_11414# 0.19fF
C1388 a_19030_12170# VDD 2.78fF
C1389 a_21038_4138# col[18] 0.38fF
C1390 a_2475_9182# a_4974_9158# 0.68fF
C1391 a_31078_16186# col[28] 0.38fF
C1392 a_2275_14202# a_27974_14178# 0.17fF
C1393 a_13006_3134# row_n[1] 0.43fF
C1394 a_12914_7150# rowon_n[5] 0.14fF
C1395 a_25054_7150# vcm 0.89fF
C1396 a_19942_14178# rowoff_n[12] 0.55fF
C1397 a_30074_7150# m2_30272_7398# 0.19fF
C1398 a_21950_2130# a_22042_2130# 0.45fF
C1399 a_16322_4178# col_n[13] 0.11fF
C1400 m2_7756_946# col_n[5] 0.45fF
C1401 a_26362_16226# col_n[23] 0.11fF
C1402 a_34090_16186# VDD 1.23fF
C1403 a_2475_7174# col[18] 0.22fF
C1404 a_2475_11190# a_20034_11166# 0.68fF
C1405 a_28066_12170# a_28066_11166# 0.84fF
C1406 a_15318_1166# vcm 0.25fF
C1407 a_5978_10162# vcm 0.89fF
C1408 a_1957_9182# m2_1732_8978# 0.33fF
C1409 a_2275_13198# col_n[25] 0.17fF
C1410 a_2275_2154# col_n[30] 0.17fF
C1411 a_2275_8178# a_10998_8154# 0.71fF
C1412 a_9994_2130# col[7] 0.38fF
C1413 a_33086_10162# rowon_n[8] 0.45fF
C1414 a_18026_13174# a_19030_13174# 0.86fF
C1415 a_20034_14178# col[17] 0.38fF
C1416 a_30378_5182# vcm 0.24fF
C1417 a_2275_10186# col[15] 0.17fF
C1418 a_21038_5142# m2_21236_5390# 0.19fF
C1419 a_21038_14178# vcm 0.89fF
C1420 a_17934_4138# VDD 0.29fF
C1421 a_2275_10186# a_26058_10162# 0.71fF
C1422 a_10998_10162# row_n[8] 0.43fF
C1423 a_5278_2170# col_n[2] 0.11fF
C1424 a_10906_14178# rowon_n[12] 0.14fF
C1425 a_15318_14218# col_n[12] 0.11fF
C1426 a_8990_15182# a_8990_14178# 0.84fF
C1427 a_11302_8194# vcm 0.24fF
C1428 a_7894_15182# rowoff_n[13] 0.68fF
C1429 a_20946_4138# rowon_n[2] 0.14fF
C1430 a_24050_3134# ctop 4.91fF
C1431 a_2475_17214# vcm 1.32fF
C1432 sample_n rowoff_n[0] 0.55fF
C1433 a_32994_8154# VDD 0.29fF
C1434 a_9902_7150# rowoff_n[5] 0.66fF
C1435 a_2275_7174# a_16322_7190# 0.15fF
C1436 a_2475_7174# a_18938_7150# 0.41fF
C1437 a_4882_2130# vcm 0.18fF
C1438 a_33086_17190# a_34090_17190# 0.86fF
C1439 a_12002_3134# m2_12200_3382# 0.19fF
C1440 a_8990_12170# col[6] 0.38fF
C1441 a_18938_5142# rowoff_n[3] 0.56fF
C1442 a_26362_12210# vcm 0.24fF
C1443 a_2275_4162# a_9902_4138# 0.17fF
C1444 a_4974_6146# ctop 4.91fF
C1445 a_13918_11166# VDD 0.29fF
C1446 a_17934_9158# a_18026_9158# 0.45fF
C1447 a_2475_9182# a_33998_9158# 0.41fF
C1448 a_2275_9182# a_31382_9198# 0.15fF
C1449 a_31078_17190# rowon_n[15] 0.45fF
C1450 a_24050_8154# col_n[21] 0.34fF
C1451 m2_34864_15002# rowon_n[13] 0.42fF
C1452 a_27974_3134# rowoff_n[1] 0.46fF
C1453 a_2275_9182# col_n[2] 0.17fF
C1454 col_n[22] rowoff_n[14] 0.18fF
C1455 m2_1732_4962# m2_2160_5390# 0.19fF
C1456 a_19942_6146# vcm 0.18fF
C1457 a_4274_12210# col_n[1] 0.11fF
C1458 a_1957_2154# sample 0.35fF
C1459 a_19030_2130# a_19030_1126# 0.84fF
C1460 col[25] rowoff_n[10] 0.18fF
C1461 a_7286_15222# vcm 0.24fF
C1462 a_2475_18218# a_12914_18194# 0.41fF
C1463 a_2275_6170# a_24962_6146# 0.17fF
C1464 a_8990_17190# row_n[15] 0.43fF
C1465 a_20034_10162# ctop 4.91fF
C1466 m2_19804_18014# col[17] 0.37fF
C1467 a_28978_15182# VDD 0.29fF
C1468 m2_21812_18014# vcm 0.71fF
C1469 a_19030_7150# row_n[5] 0.43fF
C1470 a_2475_15206# a_3878_15182# 0.41fF
C1471 a_2275_15206# a_2874_15182# 0.17fF
C1472 a_18938_11166# rowon_n[9] 0.14fF
C1473 a_35002_10162# vcm 0.18fF
C1474 a_2475_16210# col[7] 0.22fF
C1475 a_2475_3158# a_17022_3134# 0.68fF
C1476 a_2475_5166# col[12] 0.22fF
C1477 a_8990_3134# a_9994_3134# 0.86fF
C1478 a_2275_1150# m2_11772_946# 0.51fF
C1479 a_29070_2130# m2_28840_946# 0.84fF
C1480 m3_7888_1078# ctop 0.21fF
C1481 a_9902_18194# VDD 0.50fF
C1482 row_n[9] ctop 0.28fF
C1483 col_n[6] rowoff_n[15] 0.29fF
C1484 col_n[19] col[20] 6.22fF
C1485 a_32994_13174# a_33086_13174# 0.45fF
C1486 a_13006_6146# col_n[10] 0.34fF
C1487 a_2275_11190# col_n[19] 0.17fF
C1488 a_20034_11166# rowoff_n[9] 1.79fF
C1489 a_2275_17214# a_18026_17190# 0.71fF
C1490 col[9] rowoff_n[11] 0.29fF
C1491 m2_9764_18014# m2_10192_18442# 0.19fF
C1492 a_15926_13174# vcm 0.18fF
C1493 a_12002_3134# VDD 3.51fF
C1494 a_34090_6146# a_34090_5142# 0.84fF
C1495 a_2475_5166# a_32082_5142# 0.68fF
C1496 a_5978_5142# rowon_n[3] 0.45fF
C1497 a_35494_13536# VDD 0.13fF
C1498 a_2275_18218# a_28066_18194# 0.14fF
C1499 m2_12776_946# m2_13780_946# 0.86fF
C1500 a_16018_17190# ctop 4.93fF
C1501 a_2275_8178# col[9] 0.17fF
C1502 a_29070_9158# rowoff_n[7] 1.35fF
C1503 a_2275_14202# a_8290_14218# 0.15fF
C1504 a_2475_14202# a_10906_14178# 0.41fF
C1505 m2_34864_8978# m2_34864_7974# 0.84fF
C1506 m2_1732_17010# row_n[15] 0.44fF
C1507 a_33086_5142# col[30] 0.38fF
C1508 m2_34864_6970# rowoff_n[5] 1.01fF
C1509 a_2275_2154# a_23046_2130# 0.71fF
C1510 a_30986_17190# vcm 0.18fF
C1511 a_27062_7150# VDD 1.96fF
C1512 a_2475_7174# col[29] 0.22fF
C1513 a_24050_7150# a_25054_7150# 0.86fF
C1514 a_2966_14178# m2_3164_14426# 0.19fF
C1515 a_17022_14178# row_n[12] 0.43fF
C1516 a_33086_2130# vcm 0.89fF
C1517 a_2475_16210# a_25966_16186# 0.41fF
C1518 a_2275_16210# a_23350_16226# 0.15fF
C1519 a_13918_16186# a_14010_16186# 0.45fF
C1520 a_28370_5182# col_n[25] 0.11fF
C1521 a_27062_4138# row_n[2] 0.43fF
C1522 a_12002_16186# col_n[9] 0.34fF
C1523 a_26970_8154# rowon_n[6] 0.14fF
C1524 a_7986_10162# VDD 3.92fF
C1525 a_15014_9158# a_15014_8154# 0.84fF
C1526 a_2275_13198# a_16930_13174# 0.17fF
C1527 a_2275_10186# col[26] 0.17fF
C1528 a_14010_5142# vcm 0.89fF
C1529 a_7986_12170# rowoff_n[10] 2.38fF
C1530 a_2275_18218# m2_5748_18014# 0.51fF
C1531 a_2275_1150# a_28370_1166# 0.15fF
C1532 a_2475_1150# a_30986_1126# 0.41fF
C1533 a_2966_14178# vcm 0.89fF
C1534 a_3970_12170# rowon_n[10] 0.45fF
C1535 m3_26964_18146# VDD 0.11fF
C1536 a_22042_3134# col[19] 0.38fF
C1537 a_23046_14178# VDD 2.37fF
C1538 a_32082_15182# col[29] 0.38fF
C1539 a_4974_10162# a_5978_10162# 0.86fF
C1540 a_2475_10186# a_8990_10162# 0.68fF
C1541 a_14010_2130# rowon_n[0] 0.45fF
C1542 a_2275_15206# a_31990_15182# 0.17fF
C1543 a_29070_9158# vcm 0.89fF
C1544 a_24050_16186# rowoff_n[14] 1.59fF
C1545 a_23958_3134# a_24050_3134# 0.45fF
C1546 a_2275_4162# rowon_n[2] 1.99fF
C1547 a_17326_3174# col_n[14] 0.11fF
C1548 a_27366_15222# col_n[24] 0.11fF
C1549 a_3970_17190# VDD 4.34fF
C1550 a_2475_12194# a_24050_12170# 0.68fF
C1551 a_30074_13174# a_30074_12170# 0.84fF
C1552 a_2475_14202# col[1] 0.22fF
C1553 a_25054_11166# row_n[9] 0.43fF
C1554 a_2475_3158# col[6] 0.22fF
C1555 a_19334_3174# vcm 0.24fF
C1556 a_24962_15182# rowon_n[13] 0.14fF
C1557 a_9994_12170# vcm 0.89fF
C1558 a_6890_2130# VDD 0.29fF
C1559 a_35002_5142# rowon_n[3] 0.14fF
C1560 a_2275_9182# col_n[13] 0.17fF
C1561 a_11910_18194# m2_11772_18014# 0.34fF
C1562 a_2275_9182# a_15014_9158# 0.71fF
C1563 a_21038_13174# col[18] 0.38fF
C1564 a_2475_18218# m2_31852_18014# 0.62fF
C1565 a_20034_14178# a_21038_14178# 0.86fF
C1566 a_35398_7190# vcm 0.24fF
C1567 a_3270_9198# col_n[0] 0.11fF
C1568 a_25054_16186# vcm 0.89fF
C1569 a_2275_6170# col[3] 0.17fF
C1570 a_21950_6146# VDD 0.29fF
C1571 a_4882_6146# a_4974_6146# 0.45fF
C1572 a_26058_14178# m2_26256_14426# 0.19fF
C1573 a_2275_6170# a_5278_6186# 0.15fF
C1574 a_2475_6170# a_7894_6146# 0.41fF
C1575 a_12002_9158# rowon_n[7] 0.45fF
C1576 a_6282_1166# col_n[3] 0.11fF
C1577 a_2275_11190# a_30074_11166# 0.71fF
C1578 a_16322_13214# col_n[13] 0.11fF
C1579 a_27974_1126# vcm 0.18fF
C1580 a_2475_16210# col[18] 0.22fF
C1581 a_10998_16186# a_10998_15182# 0.84fF
C1582 a_2475_5166# col[23] 0.22fF
C1583 a_15318_10202# vcm 0.24fF
C1584 a_12002_17190# rowoff_n[15] 2.18fF
C1585 m2_25828_18014# VDD 2.92fF
C1586 a_10906_6146# rowoff_n[4] 0.65fF
C1587 a_28066_5142# ctop 4.91fF
C1588 a_2161_9182# VDD 0.23fF
C1589 m3_3872_18146# ctop 0.21fF
C1590 col_n[17] rowoff_n[15] 0.21fF
C1591 rowon_n[3] ctop 0.37fF
C1592 col_n[25] col[25] 0.55fF
C1593 a_2475_8178# a_22954_8154# 0.41fF
C1594 a_2275_8178# a_20338_8194# 0.15fF
C1595 a_2275_11190# col_n[30] 0.17fF
C1596 col[20] rowoff_n[11] 0.21fF
C1597 a_8898_4138# vcm 0.18fF
C1598 a_19942_4138# rowoff_n[2] 0.55fF
C1599 a_1957_11190# rowoff_n[9] 0.14fF
C1600 a_9994_11166# col[7] 0.38fF
C1601 a_33086_8154# row_n[6] 0.43fF
C1602 a_30378_14218# vcm 0.24fF
C1603 a_32994_12170# rowon_n[10] 0.14fF
C1604 a_17022_12170# m2_17220_12418# 0.19fF
C1605 a_2275_5166# a_13918_5142# 0.17fF
C1606 a_2275_8178# col[20] 0.17fF
C1607 a_8990_8154# ctop 4.91fF
C1608 a_25054_7150# col_n[22] 0.34fF
C1609 a_17934_13174# VDD 0.29fF
C1610 a_19942_10162# a_20034_10162# 0.45fF
C1611 a_28978_2130# rowoff_n[0] 0.44fF
C1612 a_5278_11206# col_n[2] 0.11fF
C1613 a_23958_8154# vcm 0.18fF
C1614 a_21038_3134# a_21038_2130# 0.84fF
C1615 a_2475_2154# a_5978_2130# 0.68fF
C1616 a_11302_17230# vcm 0.24fF
C1617 a_9994_16186# rowon_n[14] 0.45fF
C1618 a_2275_7174# a_28978_7150# 0.17fF
C1619 a_24050_12170# ctop 4.91fF
C1620 a_32994_17190# VDD 0.29fF
C1621 col[4] rowoff_n[12] 0.32fF
C1622 a_20034_6146# rowon_n[4] 0.45fF
C1623 a_2275_16210# a_6982_16186# 0.71fF
C1624 a_4882_11166# vcm 0.18fF
C1625 a_10998_4138# a_12002_4138# 0.86fF
C1626 a_7986_10162# m2_8184_10410# 0.19fF
C1627 a_2475_4162# a_21038_4138# 0.68fF
C1628 a_30986_18194# m2_30848_18014# 0.34fF
C1629 a_7986_17190# m2_7756_18014# 0.84fF
C1630 a_2475_1150# col[0] 0.20fF
C1631 a_4974_15182# ctop 4.91fF
C1632 a_14010_5142# col_n[11] 0.34fF
C1633 a_35002_14178# a_35094_14178# 0.11fF
C1634 a_24050_17190# col_n[21] 0.34fF
C1635 a_21038_10162# rowoff_n[8] 1.74fF
C1636 a_31078_15182# row_n[13] 0.43fF
C1637 a_24962_13174# rowoff_n[11] 0.49fF
C1638 a_27062_6146# m2_27260_6394# 0.19fF
C1639 a_2275_1150# a_12002_1126# 0.14fF
C1640 a_2275_7174# col_n[7] 0.17fF
C1641 a_19942_15182# vcm 0.18fF
C1642 a_16018_5142# VDD 3.09fF
C1643 a_1957_11190# sample 0.35fF
C1644 a_30074_8154# rowoff_n[6] 1.30fF
C1645 a_2475_15206# a_14922_15182# 0.41fF
C1646 a_2275_15206# a_12306_15222# 0.15fF
C1647 a_34090_4138# col[31] 0.38fF
C1648 a_2275_3158# a_27062_3134# 0.71fF
C1649 a_31078_9158# VDD 1.54fF
C1650 a_2475_14202# col[12] 0.22fF
C1651 a_26058_8154# a_27062_8154# 0.86fF
C1652 a_18026_13174# rowon_n[11] 0.45fF
C1653 a_2475_3158# col[17] 0.22fF
C1654 a_2275_12194# a_5886_12170# 0.17fF
C1655 a_2475_18218# col[3] 0.22fF
C1656 a_29374_4178# col_n[26] 0.11fF
C1657 m2_34864_3958# row_n[2] 0.38fF
C1658 a_2874_3134# vcm 0.18fF
C1659 a_28066_3134# rowon_n[1] 0.45fF
C1660 a_15926_17190# a_16018_17190# 0.45fF
C1661 a_2475_17214# a_29982_17190# 0.41fF
C1662 a_2275_17214# a_27366_17230# 0.15fF
C1663 a_13006_15182# col_n[10] 0.34fF
C1664 a_18026_4138# m2_18224_4386# 0.19fF
C1665 a_2275_9182# col_n[24] 0.17fF
C1666 a_12002_12170# VDD 3.51fF
C1667 a_17022_10162# a_17022_9158# 0.84fF
C1668 a_2275_14202# a_20946_14178# 0.17fF
C1669 a_5978_3134# row_n[1] 0.43fF
C1670 a_2275_17214# col[9] 0.17fF
C1671 a_5886_7150# rowon_n[5] 0.14fF
C1672 a_18026_7150# vcm 0.89fF
C1673 a_2275_6170# col[14] 0.17fF
C1674 a_12914_14178# rowoff_n[12] 0.63fF
C1675 a_2275_2154# a_32386_2170# 0.15fF
C1676 a_2475_2154# a_35002_2130# 0.41fF
C1677 a_23046_2130# col[20] 0.38fF
C1678 a_3878_6146# VDD 0.29fF
C1679 a_33086_14178# col[30] 0.38fF
C1680 a_27062_16186# VDD 1.96fF
C1681 a_2475_16210# col[29] 0.22fF
C1682 a_2475_11190# a_13006_11166# 0.68fF
C1683 a_6982_11166# a_7986_11166# 0.86fF
C1684 a_8290_1166# vcm 0.25fF
C1685 a_2275_16210# a_34394_16226# 0.15fF
C1686 a_33086_11166# vcm 0.89fF
C1687 a_18330_2170# col_n[15] 0.11fF
C1688 a_29982_1126# VDD 0.71fF
C1689 col_n[28] rowoff_n[15] 0.14fF
C1690 col_n[30] col[31] 6.27fF
C1691 a_25966_4138# a_26058_4138# 0.45fF
C1692 a_28370_14218# col_n[25] 0.11fF
C1693 col[31] rowoff_n[11] 0.14fF
C1694 a_27062_17190# m2_26832_18014# 0.84fF
C1695 a_2275_8178# a_3970_8154# 0.71fF
C1696 a_32082_14178# a_32082_13174# 0.84fF
C1697 a_2475_13198# a_28066_13174# 0.68fF
C1698 a_26058_10162# rowon_n[8] 0.45fF
C1699 a_23350_5182# vcm 0.24fF
C1700 a_2275_8178# col[31] 0.17fF
C1701 a_14010_14178# vcm 0.89fF
C1702 a_10906_4138# VDD 0.29fF
C1703 a_2966_12170# m2_1732_11990# 0.86fF
C1704 a_22042_12170# col[19] 0.38fF
C1705 a_2275_10186# a_19030_10162# 0.71fF
C1706 a_3970_10162# row_n[8] 0.43fF
C1707 a_2275_5166# col_n[1] 0.17fF
C1708 a_22042_15182# a_23046_15182# 0.86fF
C1709 a_4274_8194# vcm 0.24fF
C1710 a_13918_4138# rowon_n[2] 0.14fF
C1711 a_29070_18194# vcm 0.15fF
C1712 a_17022_3134# ctop 4.91fF
C1713 col[15] rowoff_n[12] 0.25fF
C1714 a_25966_8154# VDD 0.29fF
C1715 a_2161_7174# rowoff_n[5] 0.14fF
C1716 a_6890_7150# a_6982_7150# 0.45fF
C1717 a_2275_15206# m2_34864_15002# 0.51fF
C1718 a_2475_7174# a_11910_7150# 0.41fF
C1719 a_2275_7174# a_9294_7190# 0.15fF
C1720 a_17326_12210# col_n[14] 0.11fF
C1721 a_2275_2154# row_n[0] 26.41fF
C1722 a_2275_12194# a_34090_12170# 0.71fF
C1723 a_31990_3134# vcm 0.18fF
C1724 a_13006_17190# a_13006_16186# 0.84fF
C1725 a_11910_5142# rowoff_n[3] 0.64fF
C1726 a_19334_12210# vcm 0.24fF
C1727 a_2475_12194# col[6] 0.22fF
C1728 a_2475_1150# col[11] 0.22fF
C1729 a_2475_4162# a_2966_4138# 0.65fF
C1730 a_2161_4162# a_2275_4162# 0.17fF
C1731 a_32082_7150# ctop 4.91fF
C1732 a_6890_11166# VDD 0.29fF
C1733 a_2475_9182# a_26970_9158# 0.41fF
C1734 a_2275_9182# a_24354_9198# 0.15fF
C1735 a_24050_17190# rowon_n[15] 0.45fF
C1736 a_10998_10162# col[8] 0.38fF
C1737 a_20946_3134# rowoff_n[1] 0.54fF
C1738 a_2966_10162# rowoff_n[8] 2.62fF
C1739 a_2275_7174# col_n[18] 0.17fF
C1740 a_34090_7150# rowon_n[5] 0.45fF
C1741 a_12914_6146# vcm 0.18fF
C1742 a_32082_2130# a_33086_2130# 0.86fF
C1743 a_35398_16226# vcm 0.24fF
C1744 a_2475_18218# a_5886_18194# 0.41fF
C1745 a_26058_6146# col_n[23] 0.34fF
C1746 a_3270_18234# col_n[0] 0.11fF
C1747 a_35002_14178# m2_34864_13998# 0.33fF
C1748 a_2275_6170# a_17934_6146# 0.17fF
C1749 a_2475_17214# row_n[15] 0.48fF
C1750 a_13006_10162# ctop 4.91fF
C1751 a_21950_15182# VDD 0.29fF
C1752 a_2275_15206# col[3] 0.17fF
C1753 a_21950_11166# a_22042_11166# 0.45fF
C1754 a_2275_4162# col[8] 0.17fF
C1755 a_6282_10202# col_n[3] 0.11fF
C1756 m2_7756_18014# vcm 0.71fF
C1757 a_12002_7150# row_n[5] 0.43fF
C1758 a_11910_11166# rowon_n[9] 0.14fF
C1759 a_27974_10162# vcm 0.18fF
C1760 a_2475_14202# col[23] 0.22fF
C1761 a_23046_4138# a_23046_3134# 0.84fF
C1762 a_2475_3158# a_9994_3134# 0.68fF
C1763 a_2475_3158# col[28] 0.22fF
C1764 m3_34996_12122# ctop 0.22fF
C1765 a_2275_8178# a_32994_8154# 0.17fF
C1766 a_28066_14178# ctop 4.91fF
C1767 a_2475_18218# col[14] 0.22fF
C1768 a_2275_17214# a_10998_17190# 0.71fF
C1769 a_13006_11166# rowoff_n[9] 2.13fF
C1770 m2_2736_18014# m2_3164_18442# 0.19fF
C1771 a_8898_13174# vcm 0.18fF
C1772 a_4974_3134# VDD 4.23fF
C1773 a_13006_5142# a_14010_5142# 0.86fF
C1774 a_2475_5166# a_25054_5142# 0.68fF
C1775 a_2275_18218# a_21038_18194# 0.14fF
C1776 m2_5748_946# m2_6752_946# 0.86fF
C1777 a_15014_4138# col_n[12] 0.34fF
C1778 a_2275_17214# col[20] 0.17fF
C1779 a_8990_17190# ctop 4.93fF
C1780 a_25054_16186# col_n[22] 0.34fF
C1781 a_22042_9158# rowoff_n[7] 1.69fF
C1782 a_32082_14178# rowon_n[12] 0.45fF
C1783 a_2275_6170# col[25] 0.17fF
C1784 a_2275_18218# col[5] 0.17fF
C1785 a_29070_15182# rowoff_n[13] 1.35fF
C1786 m2_34864_8978# VDD 1.59fF
C1787 a_2275_2154# a_16018_2130# 0.71fF
C1788 a_2966_10162# col_n[0] 0.34fF
C1789 m2_32856_946# col[30] 0.52fF
C1790 a_23958_17190# vcm 0.18fF
C1791 m2_33860_18014# m3_33992_18146# 4.43fF
C1792 a_20034_7150# VDD 2.68fF
C1793 a_31078_7150# rowoff_n[5] 1.25fF
C1794 a_32082_15182# m2_32280_15430# 0.19fF
C1795 a_3970_7150# a_3970_6146# 0.84fF
C1796 a_9994_14178# row_n[12] 0.43fF
C1797 a_26058_2130# vcm 0.89fF
C1798 rowon_n[11] sample_n 0.15fF
C1799 ctop col[6] 0.13fF
C1800 a_2475_16210# a_18938_16186# 0.41fF
C1801 a_2275_16210# a_16322_16226# 0.15fF
C1802 a_20034_4138# row_n[2] 0.43fF
C1803 a_19942_8154# rowon_n[6] 0.14fF
C1804 a_2275_4162# a_31078_4138# 0.71fF
C1805 m3_27968_1078# m3_28972_1078# 0.21fF
C1806 a_28066_9158# a_29070_9158# 0.86fF
C1807 a_3970_17190# m2_4168_17438# 0.19fF
C1808 m2_2736_1950# vcm 0.71fF
C1809 a_3970_2130# col_n[1] 0.33fF
C1810 a_2475_10186# col[0] 0.20fF
C1811 a_30378_3174# col_n[27] 0.11fF
C1812 a_2275_13198# a_9902_13174# 0.17fF
C1813 a_14010_14178# col_n[11] 0.34fF
C1814 a_6982_5142# vcm 0.89fF
C1815 a_17934_18194# a_18026_18194# 0.11fF
C1816 a_2275_1150# a_21342_1166# 0.15fF
C1817 a_12914_1126# a_13006_1126# 0.11fF
C1818 a_2475_1150# a_23958_1126# 0.41fF
C1819 a_23046_13174# m2_23244_13422# 0.19fF
C1820 m2_34864_946# VDD 2.83fF
C1821 a_2275_16210# col_n[7] 0.17fF
C1822 a_16018_14178# VDD 3.09fF
C1823 a_2275_5166# col_n[12] 0.17fF
C1824 a_19030_11166# a_19030_10162# 0.84fF
C1825 a_6982_2130# rowon_n[0] 0.45fF
C1826 a_2275_15206# a_24962_15182# 0.17fF
C1827 a_22042_9158# vcm 0.89fF
C1828 col[26] rowoff_n[12] 0.17fF
C1829 a_17022_16186# rowoff_n[14] 1.94fF
C1830 a_34090_13174# col[31] 0.38fF
C1831 a_2275_2154# col[2] 0.17fF
C1832 a_20946_1126# m2_20808_946# 0.31fF
C1833 a_2475_12194# a_17022_12170# 0.68fF
C1834 a_8990_12170# a_9994_12170# 0.86fF
C1835 a_2475_12194# col[17] 0.22fF
C1836 a_12306_3174# vcm 0.24fF
C1837 a_18026_11166# row_n[9] 0.43fF
C1838 a_2475_1150# col[22] 0.22fF
C1839 a_17934_15182# rowon_n[13] 0.14fF
C1840 a_2874_12170# vcm 0.18fF
C1841 a_29374_13214# col_n[26] 0.11fF
C1842 a_33998_3134# VDD 0.29fF
C1843 a_14010_11166# m2_14208_11414# 0.19fF
C1844 a_27974_5142# a_28066_5142# 0.45fF
C1845 a_27974_5142# rowon_n[3] 0.14fF
C1846 a_2275_9182# a_7986_9158# 0.71fF
C1847 a_2275_7174# col_n[29] 0.17fF
C1848 a_2475_18218# m2_17796_18014# 0.62fF
C1849 a_34090_15182# a_34090_14178# 0.84fF
C1850 a_2475_14202# a_32082_14178# 0.68fF
C1851 a_2275_3158# rowoff_n[1] 0.81fF
C1852 col[10] rowoff_n[13] 0.28fF
C1853 a_27366_7190# vcm 0.24fF
C1854 a_33086_7150# m2_33284_7398# 0.19fF
C1855 a_18026_16186# vcm 0.89fF
C1856 a_2275_15206# col[14] 0.17fF
C1857 a_14922_6146# VDD 0.29fF
C1858 a_2275_4162# col[19] 0.17fF
C1859 a_23046_11166# col[20] 0.38fF
C1860 a_4974_9158# rowon_n[7] 0.45fF
C1861 a_3878_15182# VDD 0.29fF
C1862 a_2275_11190# a_23046_11166# 0.71fF
C1863 a_20946_1126# vcm 0.18fF
C1864 a_24050_16186# a_25054_16186# 0.86fF
C1865 a_8290_10202# vcm 0.24fF
C1866 a_4974_17190# rowoff_n[15] 2.52fF
C1867 m2_11772_18014# VDD 4.37fF
C1868 a_4974_9158# m2_5172_9406# 0.19fF
C1869 a_2475_18218# col[25] 0.22fF
C1870 a_21038_5142# ctop 4.91fF
C1871 a_12002_2130# m2_11772_946# 0.84fF
C1872 a_18330_11206# col_n[15] 0.11fF
C1873 a_29982_10162# VDD 0.29fF
C1874 a_2475_8178# a_15926_8154# 0.41fF
C1875 a_2275_8178# a_13310_8194# 0.15fF
C1876 a_8898_8154# a_8990_8154# 0.45fF
C1877 ctop rowoff_n[14] 0.28fF
C1878 a_34394_5182# vcm 0.24fF
C1879 a_29982_12170# rowoff_n[10] 0.43fF
C1880 a_12914_4138# rowoff_n[2] 0.63fF
C1881 a_24050_5142# m2_24248_5390# 0.19fF
C1882 a_26058_8154# row_n[6] 0.43fF
C1883 a_23350_14218# vcm 0.24fF
C1884 a_25966_12170# rowon_n[10] 0.14fF
C1885 a_2275_17214# col[31] 0.17fF
C1886 a_2275_5166# a_6890_5142# 0.17fF
C1887 a_10906_13174# VDD 0.29fF
C1888 a_2275_18218# col[16] 0.17fF
C1889 a_2475_10186# a_30986_10162# 0.41fF
C1890 a_2275_10186# a_28370_10202# 0.15fF
C1891 a_21950_2130# rowoff_n[0] 0.52fF
C1892 a_12002_9158# col[9] 0.38fF
C1893 m2_1732_15002# sample_n 0.12fF
C1894 a_16930_8154# vcm 0.18fF
C1895 a_2275_14202# col_n[1] 0.17fF
C1896 a_27062_5142# col_n[24] 0.34fF
C1897 a_2275_3158# col_n[6] 0.17fF
C1898 a_4274_17230# vcm 0.24fF
C1899 a_2874_16186# rowon_n[14] 0.14fF
C1900 a_1957_7174# VDD 0.28fF
C1901 a_2275_7174# a_21950_7150# 0.17fF
C1902 m2_34864_5966# rowon_n[4] 0.42fF
C1903 a_17022_12170# ctop 4.91fF
C1904 a_7286_9198# col_n[4] 0.11fF
C1905 a_25966_17190# VDD 0.29fF
C1906 ctop col[17] 0.13fF
C1907 row_n[6] sample_n 0.16fF
C1908 en_bit_n[1] col[15] 0.14fF
C1909 a_2966_7150# col[0] 0.38fF
C1910 a_23958_12170# a_24050_12170# 0.45fF
C1911 a_13006_6146# rowon_n[4] 0.45fF
C1912 a_15014_3134# m2_15212_3382# 0.19fF
C1913 a_31990_12170# vcm 0.18fF
C1914 a_1957_4162# row_n[2] 0.29fF
C1915 a_28066_2130# VDD 1.85fF
C1916 a_2275_10186# m2_1732_9982# 0.27fF
C1917 a_2475_4162# a_14010_4138# 0.68fF
C1918 a_25054_5142# a_25054_4138# 0.84fF
C1919 a_2475_10186# col[11] 0.22fF
C1920 m3_34996_6098# m3_34996_5094# 0.20fF
C1921 a_32082_16186# ctop 4.91fF
C1922 a_14010_10162# rowoff_n[8] 2.08fF
C1923 a_24050_15182# row_n[13] 0.43fF
C1924 a_17934_13174# rowoff_n[11] 0.57fF
C1925 a_2275_1150# a_4974_1126# 0.14fF
C1926 a_2275_16210# col_n[18] 0.17fF
C1927 a_3878_1126# a_3970_1126# 0.47fF
C1928 a_12914_15182# vcm 0.18fF
C1929 a_8990_5142# VDD 3.82fF
C1930 a_2275_5166# col_n[23] 0.17fF
C1931 a_34090_5142# row_n[3] 0.43fF
C1932 a_16018_3134# col_n[13] 0.34fF
C1933 a_2475_6170# a_29070_6146# 0.68fF
C1934 a_15014_6146# a_16018_6146# 0.86fF
C1935 a_33998_9158# rowon_n[7] 0.14fF
C1936 a_23046_8154# rowoff_n[6] 1.64fF
C1937 a_26058_15182# col_n[23] 0.34fF
C1938 a_4882_15182# a_4974_15182# 0.45fF
C1939 a_2475_15206# a_7894_15182# 0.41fF
C1940 a_2275_15206# a_5278_15222# 0.15fF
C1941 a_2275_13198# col[8] 0.17fF
C1942 m2_1732_11990# m2_1732_10986# 0.84fF
C1943 a_2275_2154# col[13] 0.17fF
C1944 a_33998_17190# rowoff_n[15] 0.39fF
C1945 a_32082_6146# rowoff_n[4] 1.20fF
C1946 a_2275_3158# a_20034_3134# 0.71fF
C1947 a_2275_1150# m2_20808_946# 0.51fF
C1948 a_24050_9158# VDD 2.27fF
C1949 m3_22948_1078# ctop 0.21fF
C1950 a_5978_8154# a_5978_7150# 0.84fF
C1951 a_10998_13174# rowon_n[11] 0.45fF
C1952 a_2475_12194# col[28] 0.22fF
C1953 m2_1732_7974# row_n[6] 0.44fF
C1954 a_30074_4138# vcm 0.89fF
C1955 a_21038_3134# rowon_n[1] 0.45fF
C1956 a_2475_17214# a_22954_17190# 0.41fF
C1957 a_2275_17214# a_20338_17230# 0.15fF
C1958 a_2275_5166# a_35094_5142# 0.14fF
C1959 a_34090_12170# m2_34864_11990# 0.86fF
C1960 a_2275_18218# a_30378_18234# 0.15fF
C1961 a_4974_12170# VDD 4.23fF
C1962 m2_16792_946# m2_17220_1374# 0.19fF
C1963 a_30074_10162# a_31078_10162# 0.86fF
C1964 a_31382_2170# col_n[28] 0.11fF
C1965 col[21] rowoff_n[13] 0.21fF
C1966 m2_34864_9982# vcm 0.73fF
C1967 a_15014_13174# col_n[12] 0.34fF
C1968 a_2275_14202# a_13918_14178# 0.17fF
C1969 col_n[4] rowoff_n[9] 0.31fF
C1970 vcm rowoff_n[5] 2.43fF
C1971 VDD rowoff_n[2] 87.22fF
C1972 col_n[3] rowoff_n[8] 0.32fF
C1973 col_n[1] rowoff_n[6] 0.33fF
C1974 col_n[0] rowoff_n[4] 0.34fF
C1975 sample rowoff_n[3] 0.22fF
C1976 col_n[2] rowoff_n[7] 0.32fF
C1977 a_10998_7150# vcm 0.89fF
C1978 a_2275_15206# col[25] 0.17fF
C1979 a_5886_14178# rowoff_n[12] 0.70fF
C1980 a_32082_12170# row_n[10] 0.43fF
C1981 a_2275_4162# col[30] 0.17fF
C1982 a_14922_2130# a_15014_2130# 0.45fF
C1983 a_2475_2154# a_27974_2130# 0.41fF
C1984 a_2275_2154# a_25358_2170# 0.15fF
C1985 a_31990_16186# rowon_n[14] 0.14fF
C1986 a_20034_16186# VDD 2.68fF
C1987 a_2475_11190# a_5978_11166# 0.68fF
C1988 a_21038_12170# a_21038_11166# 0.84fF
C1989 a_2275_1150# vcm 8.49fF
C1990 a_2275_16210# a_28978_16186# 0.17fF
C1991 a_26058_11166# vcm 0.89fF
C1992 a_22954_1126# VDD 0.78fF
C1993 m2_13780_18014# col[11] 0.39fF
C1994 a_2966_5142# ctop 4.82fF
C1995 col[5] rowoff_n[14] 0.31fF
C1996 a_19030_10162# rowon_n[8] 0.45fF
C1997 a_2475_13198# a_21038_13174# 0.68fF
C1998 a_10998_13174# a_12002_13174# 0.86fF
C1999 a_16322_5182# vcm 0.24fF
C2000 a_30378_12210# col_n[27] 0.11fF
C2001 a_3970_11166# col_n[1] 0.34fF
C2002 m2_14784_946# vcm 0.71fF
C2003 a_2475_8178# col[5] 0.22fF
C2004 a_2275_1150# a_35002_1126# 0.17fF
C2005 a_6982_14178# vcm 0.89fF
C2006 a_2275_18218# col[27] 0.17fF
C2007 a_29982_6146# a_30074_6146# 0.45fF
C2008 a_2275_10186# a_12002_10162# 0.71fF
C2009 a_3878_2130# rowoff_n[0] 0.73fF
C2010 a_2275_14202# col_n[12] 0.17fF
C2011 a_2275_3158# col_n[17] 0.17fF
C2012 a_31382_9198# vcm 0.24fF
C2013 m2_1732_11990# VDD 5.46fF
C2014 a_6890_4138# rowon_n[2] 0.14fF
C2015 a_22042_18194# vcm 0.15fF
C2016 a_9994_3134# ctop 4.91fF
C2017 VDD col_n[5] 15.19fF
C2018 vcm col_n[2] 3.22fF
C2019 a_24050_10162# col[21] 0.38fF
C2020 rowon_n[0] sample_n 0.15fF
C2021 ctop col[28] 0.13fF
C2022 a_18938_8154# VDD 0.29fF
C2023 a_2475_7174# a_4882_7150# 0.41fF
C2024 a_2275_7174# a_3878_7150# 0.17fF
C2025 a_2275_11190# col[2] 0.17fF
C2026 m2_29844_18014# col_n[27] 0.34fF
C2027 a_2275_12194# a_27062_12170# 0.71fF
C2028 a_24962_3134# vcm 0.18fF
C2029 a_26058_17190# a_27062_17190# 0.86fF
C2030 a_12306_12210# vcm 0.24fF
C2031 a_4882_5142# rowoff_n[3] 0.72fF
C2032 a_2475_10186# col[22] 0.22fF
C2033 a_19334_10202# col_n[16] 0.11fF
C2034 a_25054_7150# ctop 4.91fF
C2035 a_33998_12170# VDD 0.29fF
C2036 m3_23952_18146# m3_24956_18146# 0.21fF
C2037 a_2475_9182# a_19942_9158# 0.41fF
C2038 a_2275_9182# a_17326_9198# 0.15fF
C2039 a_17022_17190# rowon_n[15] 0.45fF
C2040 a_10906_9158# a_10998_9158# 0.45fF
C2041 a_13918_3134# rowoff_n[1] 0.61fF
C2042 a_2275_16210# col_n[29] 0.17fF
C2043 a_27062_7150# rowon_n[5] 0.45fF
C2044 a_5886_6146# vcm 0.18fF
C2045 a_34090_14178# rowoff_n[12] 1.10fF
C2046 a_27366_16226# vcm 0.24fF
C2047 a_2275_6170# a_10906_6146# 0.17fF
C2048 a_29070_14178# m2_29268_14426# 0.19fF
C2049 a_5978_10162# ctop 4.91fF
C2050 a_13006_8154# col[10] 0.38fF
C2051 a_14922_15182# VDD 0.29fF
C2052 a_2275_13198# col[19] 0.17fF
C2053 a_2475_11190# a_35002_11166# 0.41fF
C2054 a_2275_11190# a_32386_11206# 0.15fF
C2055 a_2275_2154# col[24] 0.17fF
C2056 a_4974_7150# row_n[5] 0.43fF
C2057 a_4882_11166# rowon_n[9] 0.14fF
C2058 a_28066_4138# col_n[25] 0.34fF
C2059 a_20946_10162# vcm 0.18fF
C2060 a_1957_3158# a_2275_3158# 0.19fF
C2061 a_2475_3158# a_2874_3134# 0.41fF
C2062 m3_18932_18146# ctop 0.21fF
C2063 a_8290_8194# col_n[5] 0.11fF
C2064 a_2275_8178# a_25966_8154# 0.17fF
C2065 a_21038_14178# ctop 4.91fF
C2066 a_25966_13174# a_26058_13174# 0.45fF
C2067 a_2966_3134# rowon_n[1] 0.45fF
C2068 a_5978_11166# rowoff_n[9] 2.47fF
C2069 a_2275_17214# a_3970_17190# 0.71fF
C2070 a_34394_14218# vcm 0.24fF
C2071 a_32082_4138# VDD 1.44fF
C2072 a_2475_5166# a_18026_5142# 0.68fF
C2073 a_27062_6146# a_27062_5142# 0.84fF
C2074 a_20034_12170# m2_20232_12418# 0.19fF
C2075 sample_n rowoff_n[13] 0.55fF
C2076 a_2275_18218# a_14010_18194# 0.14fF
C2077 col_n[6] rowoff_n[0] 0.29fF
C2078 col_n[9] rowoff_n[3] 0.27fF
C2079 col_n[12] rowoff_n[6] 0.25fF
C2080 col_n[15] rowoff_n[9] 0.23fF
C2081 col_n[8] rowoff_n[2] 0.28fF
C2082 col_n[13] rowoff_n[7] 0.24fF
C2083 col_n[10] rowoff_n[4] 0.27fF
C2084 col_n[7] rowoff_n[1] 0.29fF
C2085 col_n[14] rowoff_n[8] 0.24fF
C2086 col_n[11] rowoff_n[5] 0.26fF
C2087 a_15014_9158# rowoff_n[7] 2.03fF
C2088 a_25054_14178# rowon_n[12] 0.45fF
C2089 a_22042_15182# rowoff_n[13] 1.69fF
C2090 a_2275_2154# a_8990_2130# 0.71fF
C2091 a_17022_2130# col_n[14] 0.34fF
C2092 a_16930_17190# vcm 0.18fF
C2093 a_13006_7150# VDD 3.40fF
C2094 a_27062_14178# col_n[24] 0.34fF
C2095 a_24050_7150# rowoff_n[5] 1.59fF
C2096 a_2475_7174# a_33086_7150# 0.68fF
C2097 a_17022_7150# a_18026_7150# 0.86fF
C2098 a_2275_12194# col_n[6] 0.17fF
C2099 a_2275_1150# col_n[11] 0.17fF
C2100 a_1957_16210# VDD 0.28fF
C2101 a_7286_18234# col_n[4] 0.11fF
C2102 a_19030_2130# vcm 0.89fF
C2103 a_6890_16186# a_6982_16186# 0.45fF
C2104 a_2475_16210# a_11910_16186# 0.41fF
C2105 a_2275_16210# a_9294_16226# 0.15fF
C2106 a_2966_16186# col[0] 0.38fF
C2107 a_33086_5142# rowoff_n[3] 1.15fF
C2108 a_13006_4138# row_n[2] 0.43fF
C2109 col[16] rowoff_n[14] 0.24fF
C2110 a_12914_8154# rowon_n[6] 0.14fF
C2111 a_2275_4162# a_24050_4138# 0.71fF
C2112 a_10998_10162# m2_11196_10410# 0.19fF
C2113 a_28066_11166# VDD 1.85fF
C2114 m3_13912_1078# m3_14916_1078# 0.21fF
C2115 col_n[0] rowoff_n[10] 0.34fF
C2116 a_7986_9158# a_7986_8154# 0.84fF
C2117 a_2161_13198# a_2275_13198# 0.17fF
C2118 a_2475_13198# a_2966_13174# 0.65fF
C2119 a_2475_8178# col[16] 0.22fF
C2120 a_34090_6146# vcm 0.89fF
C2121 m2_16792_946# col[14] 0.51fF
C2122 a_2275_1150# a_14314_1166# 0.15fF
C2123 a_30074_6146# m2_30272_6394# 0.19fF
C2124 a_2475_1150# a_16930_1126# 0.41fF
C2125 a_32386_1166# col_n[29] 0.11fF
C2126 a_2275_14202# col_n[23] 0.17fF
C2127 a_8990_14178# VDD 3.82fF
C2128 a_32082_11166# a_33086_11166# 0.86fF
C2129 a_16018_12170# col_n[13] 0.34fF
C2130 a_2275_3158# col_n[28] 0.17fF
C2131 a_2275_15206# a_17934_15182# 0.17fF
C2132 a_33086_11166# rowon_n[9] 0.45fF
C2133 a_15014_9158# vcm 0.89fF
C2134 VDD col_n[16] 11.99fF
C2135 vcm col_n[13] 3.22fF
C2136 col[0] rowoff_n[15] 0.34fF
C2137 a_9994_16186# rowoff_n[14] 2.28fF
C2138 a_1957_8178# m2_1732_7974# 0.33fF
C2139 a_2475_3158# a_31990_3134# 0.41fF
C2140 a_2275_3158# a_29374_3174# 0.15fF
C2141 a_16930_3134# a_17022_3134# 0.45fF
C2142 a_2275_11190# col[13] 0.17fF
C2143 a_2475_12194# a_9994_12170# 0.68fF
C2144 a_23046_13174# a_23046_12170# 0.84fF
C2145 a_10998_11166# row_n[9] 0.43fF
C2146 a_5278_3174# vcm 0.24fF
C2147 a_35002_11166# rowoff_n[9] 0.38fF
C2148 a_2275_17214# a_32994_17190# 0.17fF
C2149 a_10906_15182# rowon_n[13] 0.14fF
C2150 a_21038_4138# m2_21236_4386# 0.19fF
C2151 a_30074_13174# vcm 0.89fF
C2152 a_26970_3134# VDD 0.29fF
C2153 a_20946_5142# rowon_n[3] 0.14fF
C2154 m2_28840_946# m2_29844_946# 0.86fF
C2155 a_2475_18218# m2_3740_18014# 0.62fF
C2156 a_2475_14202# a_25054_14178# 0.68fF
C2157 a_13006_14178# a_14010_14178# 0.86fF
C2158 a_4974_10162# col_n[2] 0.34fF
C2159 a_31382_11206# col_n[28] 0.11fF
C2160 a_20338_7190# vcm 0.24fF
C2161 a_33086_2130# ctop 4.93fF
C2162 a_10998_16186# vcm 0.89fF
C2163 a_7894_6146# VDD 0.29fF
C2164 a_2275_13198# col[30] 0.17fF
C2165 a_31990_7150# a_32082_7150# 0.45fF
C2166 a_2275_11190# a_16018_11166# 0.71fF
C2167 a_13918_1126# vcm 0.18fF
C2168 a_3970_16186# a_3970_15182# 0.84fF
C2169 a_2275_10186# vcm 7.71fF
C2170 a_25054_9158# col[22] 0.38fF
C2171 a_33486_1488# VDD 0.12fF
C2172 a_14010_5142# ctop 4.91fF
C2173 a_22954_10162# VDD 0.29fF
C2174 a_2475_8178# a_8898_8154# 0.41fF
C2175 a_2275_8178# a_6282_8194# 0.15fF
C2176 a_2966_14178# ctop 4.82fF
C2177 a_2275_13198# a_31078_13174# 0.71fF
C2178 a_28978_5142# vcm 0.18fF
C2179 a_5886_4138# rowoff_n[2] 0.70fF
C2180 a_22954_12170# rowoff_n[10] 0.51fF
C2181 a_2275_18218# m2_34864_18014# 0.51fF
C2182 a_20338_9198# col_n[17] 0.11fF
C2183 a_19030_8154# row_n[6] 0.43fF
C2184 a_16322_14218# vcm 0.24fF
C2185 a_18938_12170# rowon_n[10] 0.14fF
C2186 a_2475_17214# col[5] 0.22fF
C2187 col_n[21] rowoff_n[4] 0.19fF
C2188 col_n[24] rowoff_n[7] 0.16fF
C2189 col_n[17] rowoff_n[0] 0.21fF
C2190 col_n[20] rowoff_n[3] 0.19fF
C2191 col_n[23] rowoff_n[6] 0.17fF
C2192 col_n[18] rowoff_n[1] 0.21fF
C2193 col_n[25] rowoff_n[8] 0.16fF
C2194 col_n[22] rowoff_n[5] 0.18fF
C2195 col_n[19] rowoff_n[2] 0.20fF
C2196 col_n[26] rowoff_n[9] 0.15fF
C2197 a_29070_9158# ctop 4.91fF
C2198 a_2475_6170# col[10] 0.22fF
C2199 a_2475_10186# a_23958_10162# 0.41fF
C2200 a_2275_10186# a_21342_10202# 0.15fF
C2201 a_12914_10162# a_13006_10162# 0.45fF
C2202 a_14922_2130# rowoff_n[0] 0.60fF
C2203 a_28978_2130# rowon_n[0] 0.14fF
C2204 m2_1732_12994# vcm 1.11fF
C2205 a_9902_8154# vcm 0.18fF
C2206 a_2275_12194# col_n[17] 0.17fF
C2207 a_14010_3134# a_14010_2130# 0.84fF
C2208 a_31382_18234# vcm 0.25fF
C2209 a_2275_1150# col_n[22] 0.17fF
C2210 a_14010_7150# col[11] 0.38fF
C2211 m2_1732_9982# rowon_n[8] 0.43fF
C2212 a_2275_7174# a_14922_7150# 0.17fF
C2213 a_9994_12170# ctop 4.91fF
C2214 a_18938_17190# VDD 0.29fF
C2215 a_2966_12170# a_2966_11166# 0.84fF
C2216 a_5978_6146# rowon_n[4] 0.45fF
C2217 a_29070_3134# col_n[26] 0.34fF
C2218 a_2275_9182# col[7] 0.17fF
C2219 col[27] rowoff_n[14] 0.17fF
C2220 m2_34864_17010# m2_35292_17438# 0.19fF
C2221 a_24962_12170# vcm 0.18fF
C2222 a_21038_2130# VDD 2.58fF
C2223 col_n[10] rowoff_n[10] 0.27fF
C2224 a_9294_7190# col_n[6] 0.11fF
C2225 a_2475_4162# a_6982_4138# 0.68fF
C2226 a_3970_4138# a_4974_4138# 0.86fF
C2227 m3_34996_13126# m3_34996_12122# 0.20fF
C2228 a_2275_9182# a_29982_9158# 0.17fF
C2229 a_2475_8178# col[27] 0.22fF
C2230 a_25054_16186# ctop 4.91fF
C2231 a_27974_14178# a_28066_14178# 0.45fF
C2232 a_6982_10162# rowoff_n[8] 2.42fF
C2233 a_17022_15182# row_n[13] 0.43fF
C2234 a_10906_13174# rowoff_n[11] 0.65fF
C2235 a_5886_15182# vcm 0.18fF
C2236 a_2475_5166# VDD 41.96fF
C2237 a_27062_5142# row_n[3] 0.43fF
C2238 a_2475_6170# a_22042_6146# 0.68fF
C2239 a_29070_7150# a_29070_6146# 0.84fF
C2240 a_2966_13174# m2_3164_13422# 0.19fF
C2241 a_26970_9158# rowon_n[7] 0.14fF
C2242 a_16018_8154# rowoff_n[6] 1.98fF
C2243 vcm col_n[24] 3.22fF
C2244 VDD col_n[27] 9.74fF
C2245 a_13006_17190# col[10] 0.38fF
C2246 col[11] rowoff_n[15] 0.27fF
C2247 a_2275_11190# col[24] 0.17fF
C2248 a_26970_17190# rowoff_n[15] 0.47fF
C2249 a_18026_1126# col_n[15] 0.39fF
C2250 a_25054_6146# rowoff_n[4] 1.54fF
C2251 a_28066_13174# col_n[25] 0.34fF
C2252 a_2275_3158# a_13006_3134# 0.71fF
C2253 a_2475_1150# m2_6752_946# 0.62fF
C2254 m3_1864_4090# ctop 0.22fF
C2255 a_17022_9158# VDD 2.99fF
C2256 a_19030_8154# a_20034_8154# 0.86fF
C2257 a_3970_13174# rowon_n[11] 0.45fF
C2258 a_8290_17230# col_n[5] 0.11fF
C2259 a_23046_4138# vcm 0.89fF
C2260 a_34090_4138# rowoff_n[2] 1.10fF
C2261 a_14010_3134# rowon_n[1] 0.45fF
C2262 a_8898_17190# a_8990_17190# 0.45fF
C2263 a_2275_17214# a_13310_17230# 0.15fF
C2264 a_2475_17214# a_15926_17190# 0.41fF
C2265 a_2275_5166# a_28066_5142# 0.71fF
C2266 a_2275_5166# rowon_n[3] 1.99fF
C2267 a_32082_13174# VDD 1.44fF
C2268 a_2275_18218# a_23350_18234# 0.15fF
C2269 m2_9764_946# m2_10192_1374# 0.19fF
C2270 a_9994_10162# a_9994_9158# 0.84fF
C2271 a_2275_14202# a_6890_14178# 0.17fF
C2272 a_3970_7150# vcm 0.89fF
C2273 a_2475_4162# col[4] 0.22fF
C2274 a_25054_12170# row_n[10] 0.43fF
C2275 a_2475_2154# a_20946_2130# 0.41fF
C2276 a_2275_2154# a_18330_2170# 0.15fF
C2277 a_24962_16186# rowon_n[14] 0.14fF
C2278 a_17022_11166# col_n[14] 0.34fF
C2279 a_13006_16186# VDD 3.40fF
C2280 a_35002_6146# rowon_n[4] 0.14fF
C2281 a_2966_18194# vcm 0.15fF
C2282 a_2275_10186# col_n[11] 0.17fF
C2283 a_28370_2170# vcm 0.24fF
C2284 a_2275_16210# a_21950_16186# 0.17fF
C2285 a_19030_11166# vcm 0.89fF
C2286 a_15926_1126# VDD 0.86fF
C2287 a_2275_4162# a_33390_4178# 0.15fF
C2288 a_18938_4138# a_19030_4138# 0.45fF
C2289 a_6982_17190# m2_7180_17438# 0.19fF
C2290 a_2275_7174# col[1] 0.17fF
C2291 a_12002_10162# rowon_n[8] 0.45fF
C2292 a_25054_14178# a_25054_13174# 0.84fF
C2293 a_2475_13198# a_14010_13174# 0.68fF
C2294 a_9294_5182# vcm 0.24fF
C2295 a_2475_17214# col[16] 0.22fF
C2296 col_n[29] rowoff_n[1] 0.13fF
C2297 col_n[30] rowoff_n[2] 0.12fF
C2298 a_2275_1150# a_26970_1126# 0.17fF
C2299 col_n[31] rowoff_n[3] 0.11fF
C2300 col_n[28] rowoff_n[0] 0.14fF
C2301 a_34090_15182# vcm 0.89fF
C2302 a_2475_6170# col[21] 0.22fF
C2303 a_30986_5142# VDD 0.29fF
C2304 a_26058_13174# m2_26256_13422# 0.19fF
C2305 a_2275_10186# a_4974_10162# 0.71fF
C2306 a_3878_10162# a_3970_10162# 0.45fF
C2307 a_32386_10202# col_n[29] 0.11fF
C2308 a_5978_9158# col_n[3] 0.34fF
C2309 a_2475_15206# a_29070_15182# 0.68fF
C2310 a_15014_15182# a_16018_15182# 0.86fF
C2311 a_2275_12194# col_n[28] 0.17fF
C2312 a_24354_9198# vcm 0.24fF
C2313 a_15014_18194# vcm 0.15fF
C2314 a_33086_9158# row_n[7] 0.43fF
C2315 a_11910_8154# VDD 0.29fF
C2316 a_33998_8154# a_34090_8154# 0.45fF
C2317 a_32994_13174# rowon_n[11] 0.14fF
C2318 a_2275_9182# col[18] 0.17fF
C2319 a_2275_12194# a_20034_12170# 0.71fF
C2320 a_17934_3134# vcm 0.18fF
C2321 m2_26832_946# col[24] 0.51fF
C2322 a_5978_17190# a_5978_16186# 0.84fF
C2323 col_n[21] rowoff_n[10] 0.19fF
C2324 a_26058_8154# col[23] 0.38fF
C2325 a_5278_12210# vcm 0.24fF
C2326 a_17022_11166# m2_17220_11414# 0.19fF
C2327 a_18026_7150# ctop 4.91fF
C2328 a_26970_12170# VDD 0.29fF
C2329 m2_6752_946# m3_6884_1078# 4.41fF
C2330 m3_9896_18146# m3_10900_18146# 0.21fF
C2331 a_2475_9182# a_12914_9158# 0.41fF
C2332 a_2275_9182# a_10298_9198# 0.15fF
C2333 a_9994_17190# rowon_n[15] 0.45fF
C2334 a_2275_14202# a_35094_14178# 0.14fF
C2335 a_6890_3134# rowoff_n[1] 0.69fF
C2336 a_21342_8194# col_n[18] 0.11fF
C2337 a_32994_7150# vcm 0.18fF
C2338 a_20034_7150# rowon_n[5] 0.45fF
C2339 a_27062_14178# rowoff_n[12] 1.45fF
C2340 a_25054_2130# a_26058_2130# 0.86fF
C2341 a_20338_16226# vcm 0.24fF
C2342 a_2874_6146# a_2966_6146# 0.45fF
C2343 a_33086_11166# ctop 4.91fF
C2344 sample row_n[13] 0.92fF
C2345 col_n[2] row_n[15] 0.37fF
C2346 col_n[1] rowon_n[14] 0.17fF
C2347 col_n[0] rowon_n[13] 0.17fF
C2348 vcm row_n[14] 1.08fF
C2349 col_n[3] rowon_n[15] 0.17fF
C2350 VDD rowon_n[12] 4.61fF
C2351 a_7894_15182# VDD 0.29fF
C2352 col[22] rowoff_n[15] 0.20fF
C2353 a_2275_11190# a_25358_11206# 0.15fF
C2354 a_2475_11190# a_27974_11166# 0.41fF
C2355 a_14922_11166# a_15014_11166# 0.45fF
C2356 col_n[5] rowoff_n[11] 0.30fF
C2357 a_13918_10162# vcm 0.18fF
C2358 a_31078_16186# row_n[14] 0.43fF
C2359 a_7986_9158# m2_8184_9406# 0.19fF
C2360 a_15014_6146# col[12] 0.38fF
C2361 a_16018_4138# a_16018_3134# 0.84fF
C2362 a_2275_8178# col_n[5] 0.17fF
C2363 a_2275_8178# a_18938_8154# 0.17fF
C2364 a_14010_14178# ctop 4.91fF
C2365 a_30074_2130# col_n[27] 0.34fF
C2366 a_27062_5142# m2_27260_5390# 0.19fF
C2367 a_28978_14178# vcm 0.18fF
C2368 a_10298_6186# col_n[7] 0.11fF
C2369 a_25054_4138# VDD 2.16fF
C2370 a_20338_18234# col_n[17] 0.11fF
C2371 a_2475_5166# a_10998_5142# 0.68fF
C2372 a_5978_5142# a_6982_5142# 0.86fF
C2373 a_2275_18218# a_6982_18194# 0.14fF
C2374 a_2275_10186# a_33998_10162# 0.17fF
C2375 a_7986_9158# rowoff_n[7] 2.38fF
C2376 a_2475_15206# col[10] 0.22fF
C2377 a_18026_14178# rowon_n[12] 0.45fF
C2378 a_29982_15182# a_30074_15182# 0.45fF
C2379 a_2475_4162# col[15] 0.22fF
C2380 a_15014_15182# rowoff_n[13] 2.03fF
C2381 a_28066_4138# rowon_n[2] 0.45fF
C2382 a_2475_2154# a_2275_2154# 2.96fF
C2383 a_1957_2154# a_2161_2154# 0.11fF
C2384 a_9902_17190# vcm 0.18fF
C2385 a_5978_7150# VDD 4.13fF
C2386 a_17022_7150# rowoff_n[5] 1.94fF
C2387 a_2475_7174# a_26058_7150# 0.68fF
C2388 a_31078_8154# a_31078_7150# 0.84fF
C2389 a_3970_4138# col[1] 0.38fF
C2390 a_2275_10186# col_n[22] 0.17fF
C2391 a_14010_16186# col[11] 0.38fF
C2392 a_12002_2130# vcm 0.89fF
C2393 a_2275_16210# a_3878_16186# 0.17fF
C2394 a_2475_16210# a_4882_16186# 0.41fF
C2395 a_18026_3134# m2_18224_3382# 0.19fF
C2396 a_29070_12170# col_n[26] 0.34fF
C2397 a_5978_4138# row_n[2] 0.43fF
C2398 a_26058_5142# rowoff_n[3] 1.50fF
C2399 a_5886_8154# rowon_n[6] 0.14fF
C2400 a_2275_7174# col[12] 0.17fF
C2401 a_2275_4162# a_17022_4138# 0.71fF
C2402 a_21038_11166# VDD 2.58fF
C2403 m3_1864_2082# m3_1864_1078# 0.20fF
C2404 a_9294_16226# col_n[6] 0.11fF
C2405 a_21038_9158# a_22042_9158# 0.86fF
C2406 a_2475_17214# col[27] 0.22fF
C2407 row_n[8] rowoff_n[8] 0.64fF
C2408 a_27062_6146# vcm 0.89fF
C2409 a_10906_18194# a_10998_18194# 0.11fF
C2410 a_5886_1126# a_5978_1126# 0.11fF
C2411 a_2275_1150# a_7286_1166# 0.15fF
C2412 a_2475_1150# a_9902_1126# 0.41fF
C2413 m2_4744_946# VDD 7.03fF
C2414 a_2275_6170# a_32082_6146# 0.71fF
C2415 a_2475_14202# VDD 41.96fF
C2416 a_12002_11166# a_12002_10162# 0.84fF
C2417 a_2275_15206# a_10906_15182# 0.17fF
C2418 a_26058_11166# rowon_n[9] 0.45fF
C2419 a_7986_9158# vcm 0.89fF
C2420 a_2874_16186# rowoff_n[14] 0.74fF
C2421 a_2475_3158# a_24962_3134# 0.41fF
C2422 a_2275_3158# a_22346_3174# 0.15fF
C2423 a_34090_2130# m2_33860_946# 0.96fF
C2424 a_18026_10162# col_n[15] 0.34fF
C2425 a_2475_1150# m2_29844_946# 0.62fF
C2426 a_2275_9182# col[29] 0.17fF
C2427 a_2475_12194# a_2874_12170# 0.41fF
C2428 a_1957_12194# a_2275_12194# 0.19fF
C2429 a_32386_4178# vcm 0.24fF
C2430 a_3970_11166# row_n[9] 0.43fF
C2431 a_27974_11166# rowoff_n[9] 0.46fF
C2432 a_2275_17214# a_25966_17190# 0.17fF
C2433 a_2275_6170# col_n[0] 0.17fF
C2434 a_23046_13174# vcm 0.89fF
C2435 a_19942_3134# VDD 0.29fF
C2436 a_20946_5142# a_21038_5142# 0.45fF
C2437 a_2966_11166# m2_1732_10986# 0.86fF
C2438 a_13918_5142# rowon_n[3] 0.14fF
C2439 a_2275_18218# a_34394_18234# 0.15fF
C2440 m2_21812_946# m2_22816_946# 0.86fF
C2441 a_2475_14202# a_18026_14178# 0.68fF
C2442 a_27062_15182# a_27062_14178# 0.84fF
C2443 a_2275_3158# row_n[1] 26.41fF
C2444 a_13310_7190# vcm 0.24fF
C2445 a_2275_2154# a_30986_2130# 0.17fF
C2446 col_n[14] rowon_n[15] 0.17fF
C2447 a_26058_2130# ctop 4.93fF
C2448 col_n[3] row_n[10] 0.37fF
C2449 a_3970_16186# vcm 0.89fF
C2450 col_n[12] rowon_n[14] 0.17fF
C2451 col_n[10] rowon_n[13] 0.17fF
C2452 col_n[5] row_n[11] 0.37fF
C2453 VDD row_n[7] 4.64fF
C2454 col_n[13] row_n[15] 0.37fF
C2455 col_n[7] row_n[12] 0.37fF
C2456 col_n[6] rowon_n[11] 0.17fF
C2457 col_n[2] rowon_n[9] 0.17fF
C2458 col_n[4] rowon_n[10] 0.17fF
C2459 sample rowon_n[7] 0.10fF
C2460 vcm rowon_n[8] 0.91fF
C2461 col_n[8] rowon_n[12] 0.17fF
C2462 col_n[0] row_n[8] 0.37fF
C2463 col_n[1] row_n[9] 0.37fF
C2464 col_n[9] row_n[13] 0.37fF
C2465 col_n[11] row_n[14] 0.37fF
C2466 a_35002_7150# VDD 0.36fF
C2467 a_2475_13198# col[4] 0.22fF
C2468 a_2275_14202# m2_34864_13998# 0.51fF
C2469 a_2475_2154# col[9] 0.22fF
C2470 a_33390_9198# col_n[30] 0.11fF
C2471 a_6982_8154# col_n[4] 0.34fF
C2472 col_n[16] rowoff_n[11] 0.22fF
C2473 a_2275_11190# a_8990_11166# 0.71fF
C2474 a_6890_1126# vcm 0.18fF
C2475 a_2475_16210# a_33086_16186# 0.68fF
C2476 a_17022_16186# a_18026_16186# 0.86fF
C2477 m2_2736_1950# ctop 0.12fF
C2478 a_28370_11206# vcm 0.24fF
C2479 a_2275_8178# col_n[16] 0.17fF
C2480 a_26458_1488# VDD 0.13fF
C2481 a_34090_8154# rowon_n[6] 0.45fF
C2482 a_6982_5142# ctop 4.91fF
C2483 a_15926_10162# VDD 0.29fF
C2484 a_2275_13198# a_24050_13174# 0.71fF
C2485 a_2275_16210# col[1] 0.17fF
C2486 m2_1732_2954# m2_2160_3382# 0.19fF
C2487 a_27062_7150# col[24] 0.38fF
C2488 a_21950_5142# vcm 0.18fF
C2489 a_2275_5166# col[6] 0.17fF
C2490 a_15926_12170# rowoff_n[10] 0.59fF
C2491 m2_23820_946# vcm 0.71fF
C2492 a_2275_18218# m2_20808_18014# 0.51fF
C2493 a_12002_8154# row_n[6] 0.43fF
C2494 a_9294_14218# vcm 0.24fF
C2495 a_11910_12170# rowon_n[10] 0.14fF
C2496 a_35002_13174# m2_34864_12994# 0.33fF
C2497 vcm rowoff_n[12] 2.43fF
C2498 a_22042_9158# ctop 4.91fF
C2499 a_2475_15206# col[21] 0.22fF
C2500 a_30986_14178# VDD 0.29fF
C2501 a_2275_10186# a_14314_10202# 0.15fF
C2502 a_2475_10186# a_16930_10162# 0.41fF
C2503 a_2475_4162# col[26] 0.22fF
C2504 a_21950_2130# rowon_n[0] 0.14fF
C2505 a_7894_2130# rowoff_n[0] 0.68fF
C2506 a_22346_7190# col_n[19] 0.11fF
C2507 a_31990_16186# rowoff_n[14] 0.41fF
C2508 a_27062_3134# a_28066_3134# 0.86fF
C2509 a_24354_18234# vcm 0.25fF
C2510 a_2275_7174# a_7894_7150# 0.17fF
C2511 a_11910_17190# VDD 0.29fF
C2512 a_16930_12170# a_17022_12170# 0.45fF
C2513 a_2275_12194# a_29374_12210# 0.15fF
C2514 a_2475_12194# a_31990_12170# 0.41fF
C2515 a_2275_7174# col[23] 0.17fF
C2516 a_32082_15182# rowon_n[13] 0.45fF
C2517 a_16018_5142# col[13] 0.38fF
C2518 a_17934_12170# vcm 0.18fF
C2519 a_14010_2130# VDD 3.30fF
C2520 a_26058_17190# col[23] 0.38fF
C2521 a_18026_5142# a_18026_4138# 0.84fF
C2522 a_2966_11166# VDD 4.45fF
C2523 a_2275_9182# a_22954_9158# 0.17fF
C2524 a_16930_18194# m2_16792_18014# 0.34fF
C2525 a_18026_16186# ctop 4.91fF
C2526 rowon_n[4] rowoff_n[4] 20.66fF
C2527 m2_34864_6970# m2_34864_5966# 0.84fF
C2528 m2_7756_18014# col[5] 0.37fF
C2529 a_9994_15182# row_n[13] 0.43fF
C2530 a_11302_5182# col_n[8] 0.11fF
C2531 a_21342_17230# col_n[18] 0.11fF
C2532 a_32994_16186# vcm 0.18fF
C2533 a_29070_6146# VDD 1.75fF
C2534 a_20034_5142# row_n[3] 0.43fF
C2535 a_2475_6170# a_15014_6146# 0.68fF
C2536 a_32082_14178# m2_32280_14426# 0.19fF
C2537 a_7986_6146# a_8990_6146# 0.86fF
C2538 a_19942_9158# rowon_n[7] 0.14fF
C2539 a_8990_8154# rowoff_n[6] 2.33fF
C2540 a_2161_18218# VDD 0.29fF
C2541 a_31990_16186# a_32082_16186# 0.45fF
C2542 a_19942_17190# rowoff_n[15] 0.55fF
C2543 a_18026_6146# rowoff_n[4] 1.89fF
C2544 a_2275_3158# a_5978_3134# 0.71fF
C2545 a_4974_3134# col[2] 0.38fF
C2546 m3_33992_18146# ctop 0.21fF
C2547 a_9994_9158# VDD 3.71fF
C2548 row_n[10] rowoff_n[10] 0.64fF
C2549 a_3970_16186# m2_4168_16434# 0.19fF
C2550 a_33086_9158# a_33086_8154# 0.84fF
C2551 a_2475_8178# a_30074_8154# 0.68fF
C2552 a_15014_15182# col[12] 0.38fF
C2553 a_2275_17214# col_n[5] 0.17fF
C2554 a_2275_6170# col_n[10] 0.17fF
C2555 a_16018_4138# vcm 0.89fF
C2556 a_6982_3134# rowon_n[1] 0.45fF
C2557 a_27062_4138# rowoff_n[2] 1.45fF
C2558 a_30074_11166# col_n[27] 0.34fF
C2559 a_2475_17214# a_8898_17190# 0.41fF
C2560 a_2275_17214# a_6282_17230# 0.15fF
C2561 a_35398_4178# VDD 0.12fF
C2562 a_23046_12170# m2_23244_12418# 0.19fF
C2563 a_2275_5166# a_21038_5142# 0.71fF
C2564 m2_23820_18014# col_n[21] 0.33fF
C2565 a_10298_15222# col_n[7] 0.11fF
C2566 a_25054_13174# VDD 2.16fF
C2567 a_2275_18218# a_16322_18234# 0.15fF
C2568 a_2275_3158# col[0] 0.16fF
C2569 a_23046_10162# a_24050_10162# 0.86fF
C2570 col_n[15] rowon_n[10] 0.17fF
C2571 col_n[13] rowon_n[9] 0.17fF
C2572 col_n[11] rowon_n[8] 0.17fF
C2573 col_n[18] row_n[12] 0.37fF
C2574 col_n[17] rowon_n[11] 0.17fF
C2575 col_n[9] rowon_n[7] 0.17fF
C2576 col_n[25] rowon_n[15] 0.17fF
C2577 col_n[7] rowon_n[6] 0.17fF
C2578 col_n[14] row_n[10] 0.37fF
C2579 col_n[23] rowon_n[14] 0.17fF
C2580 col_n[5] rowon_n[5] 0.17fF
C2581 col_n[12] row_n[9] 0.37fF
C2582 col_n[19] rowon_n[12] 0.17fF
C2583 col_n[1] rowon_n[3] 0.17fF
C2584 col_n[0] rowon_n[2] 0.17fF
C2585 col_n[2] row_n[4] 0.37fF
C2586 col_n[20] row_n[13] 0.37fF
C2587 VDD rowon_n[1] 4.61fF
C2588 col_n[4] row_n[5] 0.37fF
C2589 sample row_n[2] 0.92fF
C2590 col_n[22] row_n[14] 0.37fF
C2591 col_n[6] row_n[6] 0.37fF
C2592 vcm row_n[3] 1.08fF
C2593 col_n[24] row_n[15] 0.37fF
C2594 col_n[8] row_n[7] 0.37fF
C2595 col_n[16] row_n[11] 0.37fF
C2596 col_n[10] row_n[8] 0.37fF
C2597 col_n[3] rowon_n[4] 0.17fF
C2598 col_n[21] rowon_n[13] 0.17fF
C2599 a_31078_8154# vcm 0.89fF
C2600 a_2475_13198# col[15] 0.22fF
C2601 a_18026_12170# row_n[10] 0.43fF
C2602 a_2475_2154# a_13918_2130# 0.41fF
C2603 a_2275_2154# a_11302_2170# 0.15fF
C2604 a_7894_2130# a_7986_2130# 0.45fF
C2605 a_2475_2154# col[20] 0.22fF
C2606 a_17934_16186# rowon_n[14] 0.14fF
C2607 col_n[27] rowoff_n[11] 0.14fF
C2608 a_5978_16186# VDD 4.13fF
C2609 a_28066_2130# row_n[0] 0.43fF
C2610 a_14010_12170# a_14010_11166# 0.84fF
C2611 a_27974_6146# rowon_n[4] 0.14fF
C2612 a_3970_13174# col[1] 0.38fF
C2613 a_21342_2170# vcm 0.24fF
C2614 a_2275_8178# col_n[27] 0.17fF
C2615 a_2275_16210# a_14922_16186# 0.17fF
C2616 a_12002_11166# vcm 0.89fF
C2617 a_8898_1126# VDD 0.94fF
C2618 a_19030_9158# col_n[16] 0.34fF
C2619 a_14010_10162# m2_14208_10410# 0.19fF
C2620 a_2475_4162# a_28978_4138# 0.41fF
C2621 a_2275_4162# a_26362_4178# 0.15fF
C2622 a_13006_17190# m2_12776_18014# 0.84fF
C2623 a_2275_16210# col[12] 0.17fF
C2624 a_2275_5166# col[17] 0.17fF
C2625 a_4974_10162# rowon_n[8] 0.45fF
C2626 a_2475_13198# a_6982_13174# 0.68fF
C2627 a_3970_13174# a_4974_13174# 0.86fF
C2628 a_28978_10162# rowoff_n[8] 0.44fF
C2629 a_3878_5142# vcm 0.18fF
C2630 a_32082_13174# rowoff_n[11] 1.20fF
C2631 col_n[11] rowoff_n[12] 0.26fF
C2632 a_33086_6146# m2_33284_6394# 0.19fF
C2633 a_2275_1150# a_19942_1126# 0.15fF
C2634 a_27062_15182# vcm 0.89fF
C2635 a_23958_5142# VDD 0.29fF
C2636 m2_27836_946# VDD 3.55fF
C2637 a_22954_6146# a_23046_6146# 0.45fF
C2638 a_3878_2130# rowon_n[0] 0.14fF
C2639 a_29070_16186# a_29070_15182# 0.84fF
C2640 a_2475_15206# a_22042_15182# 0.68fF
C2641 a_17326_9198# vcm 0.24fF
C2642 a_4974_8154# m2_5172_8402# 0.19fF
C2643 a_2275_3158# a_35002_3134# 0.17fF
C2644 a_30074_4138# ctop 4.91fF
C2645 a_7986_18194# vcm 0.15fF
C2646 a_18026_1126# m2_18224_1374# 0.19fF
C2647 a_26058_9158# row_n[7] 0.43fF
C2648 a_4882_8154# VDD 0.29fF
C2649 a_7986_7150# col_n[5] 0.34fF
C2650 a_25966_13174# rowon_n[11] 0.14fF
C2651 a_2275_12194# a_13006_12170# 0.71fF
C2652 a_10906_3134# vcm 0.18fF
C2653 a_19030_17190# a_20034_17190# 0.86fF
C2654 m2_1732_16006# sample 0.31fF
C2655 a_24050_4138# m2_24248_4386# 0.19fF
C2656 m2_27836_18014# m2_28840_18014# 0.86fF
C2657 a_32386_13214# vcm 0.24fF
C2658 ctop rowoff_n[5] 0.28fF
C2659 a_2275_15206# col_n[0] 0.17fF
C2660 a_10998_7150# ctop 4.91fF
C2661 a_19942_12170# VDD 0.29fF
C2662 a_2275_4162# col_n[4] 0.17fF
C2663 m2_32856_946# m2_33284_1374# 0.19fF
C2664 a_2874_17190# rowon_n[15] 0.14fF
C2665 a_2275_9182# a_3270_9198# 0.15fF
C2666 a_2475_9182# a_5886_9158# 0.41fF
C2667 a_28066_6146# col[25] 0.38fF
C2668 a_2275_14202# a_28066_14178# 0.71fF
C2669 a_2475_1150# m2_2736_946# 0.59fF
C2670 a_13006_7150# rowon_n[5] 0.45fF
C2671 a_25966_7150# vcm 0.18fF
C2672 a_20034_14178# rowoff_n[12] 1.79fF
C2673 a_2275_1150# ctop 0.19fF
C2674 a_13310_16226# vcm 0.24fF
C2675 a_1957_5166# row_n[3] 0.29fF
C2676 a_26058_11166# ctop 4.91fF
C2677 a_35002_16186# VDD 0.36fF
C2678 a_23350_6186# col_n[20] 0.11fF
C2679 a_2275_11190# a_18330_11206# 0.15fF
C2680 a_2475_11190# a_20946_11166# 0.41fF
C2681 a_2475_11190# col[9] 0.22fF
C2682 m2_10768_946# col[8] 0.51fF
C2683 a_33390_18234# col_n[30] 0.11fF
C2684 a_6982_17190# col_n[4] 0.34fF
C2685 a_6890_10162# vcm 0.18fF
C2686 a_24050_16186# row_n[14] 0.43fF
C2687 a_2275_9182# m2_1732_8978# 0.27fF
C2688 a_29070_4138# a_30074_4138# 0.86fF
C2689 a_2275_17214# col_n[16] 0.17fF
C2690 a_2275_8178# a_11910_8154# 0.17fF
C2691 a_32082_17190# m2_31852_18014# 0.84fF
C2692 a_2275_6170# col_n[21] 0.17fF
C2693 a_6982_14178# ctop 4.91fF
C2694 a_34090_6146# row_n[4] 0.43fF
C2695 a_2275_18218# col_n[1] 0.17fF
C2696 a_18938_13174# a_19030_13174# 0.45fF
C2697 a_2275_13198# a_33390_13214# 0.15fF
C2698 a_33998_10162# rowon_n[8] 0.14fF
C2699 a_17022_4138# col[14] 0.38fF
C2700 a_27062_16186# col[24] 0.38fF
C2701 a_2275_14202# col[6] 0.17fF
C2702 a_21950_14178# vcm 0.18fF
C2703 a_18026_4138# VDD 2.89fF
C2704 a_2275_3158# col[11] 0.17fF
C2705 a_2275_5166# a_2966_5142# 0.67fF
C2706 a_2475_5166# a_3970_5142# 0.68fF
C2707 a_20034_6146# a_20034_5142# 0.84fF
C2708 a_2275_10186# a_26970_10162# 0.17fF
C2709 col_n[11] row_n[3] 0.37fF
C2710 col_n[30] rowon_n[12] 0.17fF
C2711 col_n[9] row_n[2] 0.37fF
C2712 col_n[7] row_n[1] 0.37fF
C2713 col_n[26] rowon_n[10] 0.17fF
C2714 col_n[5] row_n[0] 0.37fF
C2715 col_n[24] rowon_n[9] 0.17fF
C2716 col_n[22] rowon_n[8] 0.17fF
C2717 col_n[29] row_n[12] 0.37fF
C2718 col_n[8] rowon_n[1] 0.17fF
C2719 col_n[15] row_n[5] 0.37fF
C2720 col_n[13] row_n[4] 0.37fF
C2721 col_n[31] row_n[13] 0.37fF
C2722 col_n[6] rowon_n[0] 0.17fF
C2723 VDD analog_in 0.63fF
C2724 col_n[17] row_n[6] 0.37fF
C2725 col_n[10] rowon_n[2] 0.17fF
C2726 col_n[19] row_n[7] 0.37fF
C2727 col_n[12] rowon_n[3] 0.17fF
C2728 col_n[27] row_n[11] 0.37fF
C2729 col_n[1] en_C0_n 0.19fF
C2730 col_n[21] row_n[8] 0.37fF
C2731 col_n[14] rowon_n[4] 0.17fF
C2732 col_n[23] row_n[9] 0.37fF
C2733 col_n[16] rowon_n[5] 0.17fF
C2734 col_n[25] row_n[10] 0.37fF
C2735 col_n[18] rowon_n[6] 0.17fF
C2736 col_n[20] rowon_n[7] 0.17fF
C2737 col_n[28] rowon_n[11] 0.17fF
C2738 a_10998_14178# rowon_n[12] 0.45fF
C2739 a_2475_13198# col[26] 0.22fF
C2740 a_12306_4178# col_n[9] 0.11fF
C2741 a_2475_2154# col[31] 0.22fF
C2742 a_22346_16226# col_n[19] 0.11fF
C2743 a_7986_15182# rowoff_n[13] 2.38fF
C2744 a_21038_4138# rowon_n[2] 0.45fF
C2745 m2_5748_18014# m3_5880_18146# 4.41fF
C2746 a_33086_8154# VDD 1.34fF
C2747 a_9994_7150# rowoff_n[5] 2.28fF
C2748 a_2475_7174# a_19030_7150# 0.68fF
C2749 a_9994_7150# a_10998_7150# 0.86fF
C2750 a_4974_2130# vcm 0.89fF
C2751 a_33998_17190# a_34090_17190# 0.45fF
C2752 a_19030_5142# rowoff_n[3] 1.84fF
C2753 a_5978_2130# col[3] 0.38fF
C2754 a_2275_16210# col[23] 0.17fF
C2755 a_34090_11166# m2_34864_10986# 0.86fF
C2756 a_2275_4162# a_9994_4138# 0.71fF
C2757 a_16018_14178# col[13] 0.38fF
C2758 a_2275_5166# col[28] 0.17fF
C2759 a_32082_13174# row_n[11] 0.43fF
C2760 a_14010_11166# VDD 3.30fF
C2761 a_31990_17190# rowon_n[15] 0.14fF
C2762 a_2475_9182# a_34090_9158# 0.68fF
C2763 m2_34864_3958# rowoff_n[2] 1.01fF
C2764 a_31078_10162# col_n[28] 0.34fF
C2765 a_28066_3134# rowoff_n[1] 1.40fF
C2766 col_n[22] rowoff_n[12] 0.18fF
C2767 a_20034_6146# vcm 0.89fF
C2768 a_11302_14218# col_n[8] 0.11fF
C2769 a_2275_6170# a_25054_6146# 0.71fF
C2770 a_29070_15182# VDD 1.75fF
C2771 a_25054_11166# a_26058_11166# 0.86fF
C2772 m2_22816_18014# vcm 0.71fF
C2773 a_2874_15182# a_2966_15182# 0.45fF
C2774 a_19030_11166# rowon_n[9] 0.45fF
C2775 a_35094_10162# vcm 0.15fF
C2776 a_2475_3158# a_17934_3134# 0.41fF
C2777 a_2275_3158# a_15318_3174# 0.15fF
C2778 a_9902_3134# a_9994_3134# 0.45fF
C2779 a_2275_1150# m2_12776_946# 0.51fF
C2780 a_2475_9182# col[3] 0.22fF
C2781 m3_9896_1078# ctop 0.21fF
C2782 a_4974_12170# col[2] 0.38fF
C2783 col_n[6] rowoff_n[13] 0.29fF
C2784 a_16018_13174# a_16018_12170# 0.84fF
C2785 a_25358_4178# vcm 0.24fF
C2786 a_2275_17214# a_18938_17190# 0.17fF
C2787 a_20946_11166# rowoff_n[9] 0.54fF
C2788 a_20034_8154# col_n[17] 0.34fF
C2789 col[4] rowoff_n[4] 0.32fF
C2790 col[3] rowoff_n[3] 0.33fF
C2791 col[2] rowoff_n[2] 0.33fF
C2792 col[1] rowoff_n[1] 0.34fF
C2793 col[0] rowoff_n[0] 0.34fF
C2794 col[5] rowoff_n[5] 0.31fF
C2795 col[6] rowoff_n[6] 0.31fF
C2796 col[7] rowoff_n[7] 0.30fF
C2797 col[8] rowoff_n[8] 0.29fF
C2798 col[9] rowoff_n[9] 0.29fF
C2799 a_2275_15206# col_n[10] 0.17fF
C2800 a_16018_13174# vcm 0.89fF
C2801 a_2275_4162# col_n[15] 0.17fF
C2802 a_12914_3134# VDD 0.29fF
C2803 a_2275_5166# a_30378_5182# 0.15fF
C2804 a_2475_5166# a_32994_5142# 0.41fF
C2805 a_6890_5142# rowon_n[3] 0.14fF
C2806 a_2275_18218# a_28978_18194# 0.17fF
C2807 a_35398_13214# VDD 0.12fF
C2808 a_29982_9158# rowoff_n[7] 0.43fF
C2809 a_2275_12194# col[0] 0.16fF
C2810 a_5978_14178# a_6982_14178# 0.86fF
C2811 a_2475_14202# a_10998_14178# 0.68fF
C2812 a_2275_1150# col[5] 0.17fF
C2813 a_6282_7190# vcm 0.24fF
C2814 a_1957_14202# rowoff_n[12] 0.14fF
C2815 a_2275_2154# a_23958_2130# 0.17fF
C2816 a_19030_2130# ctop 4.91fF
C2817 a_31078_17190# vcm 0.89fF
C2818 a_27974_7150# VDD 0.29fF
C2819 a_24962_7150# a_25054_7150# 0.45fF
C2820 a_2475_11190# col[20] 0.22fF
C2821 a_2475_11190# a_2275_11190# 2.96fF
C2822 a_1957_11190# a_2161_11190# 0.11fF
C2823 a_33998_2130# vcm 0.17fF
C2824 a_31078_17190# a_31078_16186# 0.84fF
C2825 a_2475_16210# a_26058_16186# 0.68fF
C2826 a_21342_11206# vcm 0.24fF
C2827 a_2275_17214# col_n[27] 0.17fF
C2828 a_19430_1488# VDD 0.15fF
C2829 a_27062_8154# rowon_n[6] 0.45fF
C2830 a_8990_6146# col_n[6] 0.34fF
C2831 a_34090_6146# ctop 4.80fF
C2832 a_2275_18218# col_n[12] 0.17fF
C2833 a_8898_10162# VDD 0.29fF
C2834 a_9994_17190# m2_10192_17438# 0.19fF
C2835 a_2275_13198# a_17022_13174# 0.71fF
C2836 a_2275_14202# col[17] 0.17fF
C2837 a_14922_5142# vcm 0.18fF
C2838 a_8898_12170# rowoff_n[10] 0.67fF
C2839 a_2275_3158# col[22] 0.17fF
C2840 a_2275_18218# m2_6752_18014# 0.51fF
C2841 a_4974_8154# row_n[6] 0.43fF
C2842 a_3878_14178# vcm 0.18fF
C2843 a_4882_12170# rowon_n[10] 0.14fF
C2844 a_29070_13174# m2_29268_13422# 0.19fF
C2845 col_n[30] row_n[7] 0.37fF
C2846 VDD col[10] 10.96fF
C2847 col_n[21] rowon_n[2] 0.17fF
C2848 col_n[28] row_n[6] 0.37fF
C2849 col_n[3] col[4] 6.22fF
C2850 col_n[19] rowon_n[1] 0.17fF
C2851 col_n[26] row_n[5] 0.37fF
C2852 col_n[17] rowon_n[0] 0.17fF
C2853 col_n[24] row_n[4] 0.37fF
C2854 col_n[22] row_n[3] 0.37fF
C2855 col_n[20] row_n[2] 0.37fF
C2856 col_n[25] rowon_n[4] 0.17fF
C2857 col_n[23] rowon_n[3] 0.17fF
C2858 col_n[27] rowon_n[5] 0.17fF
C2859 vcm col[7] 6.66fF
C2860 col_n[29] rowon_n[6] 0.17fF
C2861 col_n[31] rowon_n[7] 0.17fF
C2862 col_n[16] row_n[0] 0.37fF
C2863 col_n[18] row_n[1] 0.37fF
C2864 a_15014_9158# ctop 4.91fF
C2865 a_23958_14178# VDD 0.29fF
C2866 a_29070_5142# col[26] 0.38fF
C2867 a_5886_10162# a_5978_10162# 0.45fF
C2868 a_2275_10186# a_7286_10202# 0.15fF
C2869 a_2475_10186# a_9902_10162# 0.41fF
C2870 a_14922_2130# rowon_n[0] 0.14fF
C2871 a_2275_15206# a_32082_15182# 0.71fF
C2872 a_29982_9158# vcm 0.18fF
C2873 a_24962_16186# rowoff_n[14] 0.49fF
C2874 a_2966_4138# rowon_n[2] 0.45fF
C2875 a_6982_3134# a_6982_2130# 0.84fF
C2876 a_17326_18234# vcm 0.25fF
C2877 a_25966_1126# m2_25828_946# 0.31fF
C2878 a_24354_5182# col_n[21] 0.11fF
C2879 a_30074_13174# ctop 4.91fF
C2880 a_4882_17190# VDD 0.29fF
C2881 a_7986_16186# col_n[5] 0.34fF
C2882 a_2475_12194# a_24962_12170# 0.41fF
C2883 a_2275_12194# a_22346_12210# 0.15fF
C2884 a_25054_15182# rowon_n[13] 0.45fF
C2885 a_10906_12170# vcm 0.18fF
C2886 m2_2736_946# col[0] 0.51fF
C2887 a_6982_2130# VDD 4.02fF
C2888 a_20034_11166# m2_20232_11414# 0.19fF
C2889 a_31078_5142# a_32082_5142# 0.86fF
C2890 m2_11772_946# m3_11904_1078# 4.41fF
C2891 a_2275_9182# a_15926_9158# 0.17fF
C2892 a_10998_16186# ctop 4.91fF
C2893 a_2275_13198# col_n[4] 0.17fF
C2894 a_2475_18218# m2_32856_18014# 0.62fF
C2895 a_20946_14178# a_21038_14178# 0.45fF
C2896 a_2275_2154# col_n[9] 0.17fF
C2897 a_18026_3134# col[15] 0.38fF
C2898 a_1957_6170# vcm 0.16fF
C2899 a_28066_15182# col[25] 0.38fF
C2900 m2_34864_4962# VDD 1.59fF
C2901 a_25966_16186# vcm 0.18fF
C2902 a_22042_6146# VDD 2.47fF
C2903 a_13006_5142# row_n[3] 0.43fF
C2904 a_22042_7150# a_22042_6146# 0.84fF
C2905 a_2475_6170# a_7986_6146# 0.68fF
C2906 a_2275_10186# ctop 0.14fF
C2907 a_12914_9158# rowon_n[7] 0.14fF
C2908 a_2475_8178# rowoff_n[6] 4.75fF
C2909 a_2275_11190# a_30986_11166# 0.17fF
C2910 a_13310_3174# col_n[10] 0.11fF
C2911 a_28066_1126# vcm 0.15fF
C2912 a_23350_15222# col_n[20] 0.11fF
C2913 a_2475_9182# col[14] 0.22fF
C2914 a_12914_17190# rowoff_n[15] 0.63fF
C2915 m2_26832_18014# VDD 2.85fF
C2916 a_10998_9158# m2_11196_9406# 0.19fF
C2917 a_10998_6146# rowoff_n[4] 2.23fF
C2918 a_17022_2130# m2_16792_946# 0.84fF
C2919 m3_5880_18146# ctop 0.21fF
C2920 a_2874_9158# VDD 0.29fF
C2921 col_n[17] rowoff_n[13] 0.21fF
C2922 a_12002_8154# a_13006_8154# 0.86fF
C2923 a_2475_8178# a_23046_8154# 0.68fF
C2924 a_2275_15206# col_n[21] 0.17fF
C2925 col[11] rowoff_n[0] 0.27fF
C2926 col[12] rowoff_n[1] 0.27fF
C2927 col[13] rowoff_n[2] 0.26fF
C2928 col[14] rowoff_n[3] 0.25fF
C2929 col[15] rowoff_n[4] 0.25fF
C2930 col[16] rowoff_n[5] 0.24fF
C2931 col[17] rowoff_n[6] 0.23fF
C2932 col[18] rowoff_n[7] 0.23fF
C2933 col[19] rowoff_n[8] 0.22fF
C2934 col[20] rowoff_n[9] 0.21fF
C2935 a_2275_4162# col_n[26] 0.17fF
C2936 a_8990_4138# vcm 0.89fF
C2937 a_2275_11190# rowoff_n[9] 0.81fF
C2938 a_20034_4138# rowoff_n[2] 1.79fF
C2939 a_30074_5142# m2_30272_5390# 0.19fF
C2940 a_30986_1126# a_31078_1126# 0.11fF
C2941 a_17022_13174# col[14] 0.38fF
C2942 a_33086_12170# rowon_n[10] 0.45fF
C2943 a_2275_5166# a_14010_5142# 0.71fF
C2944 a_18026_13174# VDD 2.89fF
C2945 a_2275_18218# a_9294_18234# 0.15fF
C2946 a_2275_12194# col[11] 0.17fF
C2947 m2_20808_946# col[18] 0.51fF
C2948 a_2275_1150# col[16] 0.16fF
C2949 a_32082_9158# col_n[29] 0.34fF
C2950 a_29070_2130# rowoff_n[0] 1.35fF
C2951 a_24050_8154# vcm 0.89fF
C2952 a_12306_13214# col_n[9] 0.11fF
C2953 a_10998_12170# row_n[10] 0.43fF
C2954 a_1957_7174# m2_1732_6970# 0.33fF
C2955 a_2475_2154# a_6890_2130# 0.41fF
C2956 a_2275_2154# a_4274_2170# 0.15fF
C2957 a_2475_11190# col[31] 0.22fF
C2958 col_n[1] rowoff_n[14] 0.33fF
C2959 a_10906_16186# rowon_n[14] 0.14fF
C2960 a_2275_7174# a_29070_7150# 0.71fF
C2961 a_21038_2130# row_n[0] 0.43fF
C2962 a_33086_17190# VDD 1.34fF
C2963 col[4] rowoff_n[10] 0.32fF
C2964 a_27062_12170# a_28066_12170# 0.86fF
C2965 a_20946_6146# rowon_n[4] 0.14fF
C2966 a_14314_2170# vcm 0.24fF
C2967 a_2275_16210# a_7894_16186# 0.17fF
C2968 a_21038_3134# m2_21236_3382# 0.19fF
C2969 a_4974_11166# vcm 0.89fF
C2970 a_2275_18218# col_n[23] 0.17fF
C2971 a_2275_4162# a_19334_4178# 0.15fF
C2972 a_2475_4162# a_21950_4138# 0.41fF
C2973 a_11910_4138# a_12002_4138# 0.45fF
C2974 a_5978_11166# col[3] 0.38fF
C2975 a_2275_14202# col[28] 0.17fF
C2976 a_18026_14178# a_18026_13174# 0.84fF
C2977 a_21950_10162# rowoff_n[8] 0.52fF
C2978 a_21038_7150# col_n[18] 0.34fF
C2979 a_29374_6186# vcm 0.24fF
C2980 a_25054_13174# rowoff_n[11] 1.54fF
C2981 col_n[30] rowon_n[1] 0.17fF
C2982 col_n[9] col[9] 0.50fF
C2983 col_n[27] row_n[0] 0.37fF
C2984 a_2275_1150# a_12914_1126# 0.17fF
C2985 VDD col[21] 8.24fF
C2986 col_n[29] row_n[1] 0.37fF
C2987 col_n[31] row_n[2] 0.37fF
C2988 vcm col[18] 6.66fF
C2989 col_n[28] rowon_n[0] 0.17fF
C2990 a_20034_15182# vcm 0.89fF
C2991 a_16930_5142# VDD 0.29fF
C2992 a_2275_6170# a_35398_6186# 0.15fF
C2993 a_30986_8154# rowoff_n[6] 0.42fF
C2994 a_2475_15206# a_15014_15182# 0.68fF
C2995 a_7986_15182# a_8990_15182# 0.86fF
C2996 a_10298_9198# vcm 0.24fF
C2997 a_2275_3158# a_27974_3134# 0.17fF
C2998 a_23046_4138# ctop 4.91fF
C2999 a_19030_9158# row_n[7] 0.43fF
C3000 a_31990_9158# VDD 0.29fF
C3001 a_26970_8154# a_27062_8154# 0.45fF
C3002 a_18938_13174# rowon_n[11] 0.14fF
C3003 a_2275_12194# a_5978_12170# 0.71fF
C3004 a_2475_7174# col[8] 0.22fF
C3005 a_28978_3134# rowon_n[1] 0.14fF
C3006 a_2475_17214# a_30074_17190# 0.68fF
C3007 m2_20808_18014# m2_21812_18014# 0.86fF
C3008 a_9994_5142# col_n[7] 0.34fF
C3009 a_25358_13214# vcm 0.24fF
C3010 a_20034_17190# col_n[17] 0.34fF
C3011 a_3970_7150# ctop 4.91fF
C3012 a_2275_13198# col_n[15] 0.17fF
C3013 a_12914_12170# VDD 0.29fF
C3014 m2_25828_946# m2_26256_1374# 0.19fF
C3015 a_2275_2154# col_n[20] 0.17fF
C3016 m2_1732_10986# sample_n 0.12fF
C3017 a_2275_14202# a_21038_14178# 0.71fF
C3018 a_5978_7150# rowon_n[5] 0.45fF
C3019 a_18938_7150# vcm 0.18fF
C3020 a_13006_14178# rowoff_n[12] 2.13fF
C3021 a_2275_10186# col[5] 0.17fF
C3022 a_18026_2130# a_19030_2130# 0.86fF
C3023 a_6282_16226# vcm 0.24fF
C3024 a_34394_6186# col_n[31] 0.11fF
C3025 a_30074_4138# col[27] 0.38fF
C3026 a_19030_11166# ctop 4.91fF
C3027 a_27974_16186# VDD 0.29fF
C3028 a_7894_11166# a_7986_11166# 0.45fF
C3029 a_2475_11190# a_13918_11166# 0.41fF
C3030 a_2275_11190# a_11302_11206# 0.15fF
C3031 a_2475_9182# col[25] 0.22fF
C3032 a_33998_11166# vcm 0.18fF
C3033 col_n[28] rowoff_n[13] 0.14fF
C3034 a_17022_16186# row_n[14] 0.43fF
C3035 a_8990_4138# a_8990_3134# 0.84fF
C3036 a_25358_4178# col_n[22] 0.11fF
C3037 col[31] rowoff_n[9] 0.14fF
C3038 col[30] rowoff_n[8] 0.15fF
C3039 col[29] rowoff_n[7] 0.15fF
C3040 col[28] rowoff_n[6] 0.16fF
C3041 col[27] rowoff_n[5] 0.17fF
C3042 col[26] rowoff_n[4] 0.17fF
C3043 col[25] rowoff_n[3] 0.18fF
C3044 col[24] rowoff_n[2] 0.19fF
C3045 col[23] rowoff_n[1] 0.19fF
C3046 col[22] rowoff_n[0] 0.20fF
C3047 a_2966_8154# a_3970_8154# 0.86fF
C3048 a_2275_8178# a_4882_8154# 0.17fF
C3049 a_8990_15182# col_n[6] 0.34fF
C3050 a_34090_15182# ctop 4.80fF
C3051 a_27062_6146# row_n[4] 0.43fF
C3052 a_26970_10162# rowon_n[8] 0.14fF
C3053 a_2275_13198# a_26362_13214# 0.15fF
C3054 a_2475_13198# a_28978_13174# 0.41fF
C3055 a_1957_4162# rowoff_n[2] 0.14fF
C3056 a_14922_14178# vcm 0.18fF
C3057 a_10998_4138# VDD 3.61fF
C3058 a_2275_12194# col[22] 0.17fF
C3059 a_33086_6146# a_34090_6146# 0.86fF
C3060 a_2966_12170# m2_3164_12418# 0.19fF
C3061 a_2275_1150# col[27] 0.17fF
C3062 a_2275_10186# a_19942_10162# 0.17fF
C3063 a_19030_2130# col[16] 0.38fF
C3064 a_3970_14178# rowon_n[12] 0.45fF
C3065 a_29070_14178# col[26] 0.38fF
C3066 a_22954_15182# a_23046_15182# 0.45fF
C3067 m2_1732_9982# m2_1732_8978# 0.84fF
C3068 col_n[12] rowoff_n[14] 0.25fF
C3069 a_14010_4138# rowon_n[2] 0.45fF
C3070 a_29982_18194# vcm 0.18fF
C3071 col[15] rowoff_n[10] 0.25fF
C3072 a_26058_8154# VDD 2.06fF
C3073 a_2874_7150# rowoff_n[5] 0.74fF
C3074 a_24050_8154# a_24050_7150# 0.84fF
C3075 a_2475_7174# a_12002_7150# 0.68fF
C3076 a_14314_2170# col_n[11] 0.11fF
C3077 a_2275_12194# a_35002_12170# 0.17fF
C3078 a_2275_6170# rowon_n[4] 1.99fF
C3079 a_24354_14218# col_n[21] 0.11fF
C3080 a_32082_3134# vcm 0.89fF
C3081 a_12002_5142# rowoff_n[3] 2.18fF
C3082 a_2275_4162# a_2874_4138# 0.17fF
C3083 a_2475_4162# a_3878_4138# 0.41fF
C3084 a_25054_13174# row_n[11] 0.43fF
C3085 a_2475_5166# col[2] 0.22fF
C3086 a_6982_11166# VDD 4.02fF
C3087 a_14010_9158# a_15014_9158# 0.86fF
C3088 a_2475_9182# a_27062_9158# 0.68fF
C3089 a_24962_17190# rowon_n[15] 0.14fF
C3090 m2_34864_5966# vcm 0.73fF
C3091 a_3878_10162# rowoff_n[8] 0.73fF
C3092 a_21038_3134# rowoff_n[1] 1.74fF
C3093 vcm col[29] 6.66fF
C3094 row_n[14] ctop 0.28fF
C3095 VDD sample_n 15.71fF
C3096 col_n[14] col[15] 6.22fF
C3097 rowon_n[6] row_n[6] 21.02fF
C3098 a_35002_7150# rowon_n[5] 0.14fF
C3099 a_13006_6146# vcm 0.89fF
C3100 a_2275_11190# col_n[9] 0.17fF
C3101 a_18026_12170# col[15] 0.38fF
C3102 a_32994_2130# a_33086_2130# 0.45fF
C3103 a_1957_15206# vcm 0.16fF
C3104 a_2275_6170# a_18026_6146# 0.71fF
C3105 a_33086_8154# col_n[30] 0.34fF
C3106 a_22042_15182# VDD 2.47fF
C3107 a_4974_11166# a_4974_10162# 0.84fF
C3108 m2_8760_18014# vcm 0.71fF
C3109 a_13310_12210# col_n[10] 0.11fF
C3110 a_12002_11166# rowon_n[9] 0.45fF
C3111 a_28066_10162# vcm 0.89fF
C3112 a_2275_3158# a_8290_3174# 0.15fF
C3113 a_2475_3158# a_10906_3134# 0.41fF
C3114 m3_34996_11118# ctop 0.22fF
C3115 a_2475_7174# col[19] 0.22fF
C3116 a_6982_16186# m2_7180_16434# 0.19fF
C3117 a_2275_8178# a_33086_8154# 0.71fF
C3118 a_29070_13174# a_30074_13174# 0.86fF
C3119 a_18330_4178# vcm 0.24fF
C3120 a_13918_11166# rowoff_n[9] 0.61fF
C3121 a_2275_17214# a_11910_17190# 0.17fF
C3122 a_8990_13174# vcm 0.89fF
C3123 a_2275_13198# col_n[26] 0.17fF
C3124 a_5886_3134# VDD 0.29fF
C3125 a_2275_2154# col_n[31] 0.17fF
C3126 a_6982_10162# col[4] 0.38fF
C3127 a_13918_5142# a_14010_5142# 0.45fF
C3128 a_26058_12170# m2_26256_12418# 0.19fF
C3129 a_2275_5166# a_23350_5182# 0.15fF
C3130 a_2475_5166# a_25966_5142# 0.41fF
C3131 a_2275_18218# a_21950_18194# 0.17fF
C3132 a_33086_10162# row_n[8] 0.43fF
C3133 a_22954_9158# rowoff_n[7] 0.51fF
C3134 a_22042_6146# col_n[19] 0.34fF
C3135 a_32994_14178# rowon_n[12] 0.14fF
C3136 a_20034_15182# a_20034_14178# 0.84fF
C3137 a_2475_14202# a_3970_14178# 0.68fF
C3138 a_2275_14202# a_2966_14178# 0.67fF
C3139 a_2275_10186# col[16] 0.17fF
C3140 a_33390_8194# vcm 0.24fF
C3141 a_29982_15182# rowoff_n[13] 0.43fF
C3142 m2_1732_7974# VDD 5.46fF
C3143 a_2275_2154# a_16930_2130# 0.17fF
C3144 a_12002_2130# ctop 4.93fF
C3145 a_24050_17190# vcm 0.89fF
C3146 a_20946_7150# VDD 0.29fF
C3147 a_31990_7150# rowoff_n[5] 0.41fF
C3148 a_26970_2130# vcm 0.18fF
C3149 a_2475_16210# a_19030_16186# 0.68fF
C3150 a_9994_16186# a_10998_16186# 0.86fF
C3151 a_14314_11206# vcm 0.24fF
C3152 a_12402_1488# VDD 0.16fF
C3153 a_20034_8154# rowon_n[6] 0.45fF
C3154 a_17022_10162# m2_17220_10410# 0.19fF
C3155 a_2275_4162# a_31990_4138# 0.17fF
C3156 a_27062_6146# ctop 4.91fF
C3157 m3_28972_1078# m3_29976_1078# 0.21fF
C3158 a_28978_9158# a_29070_9158# 0.45fF
C3159 a_2275_13198# a_9994_13174# 0.71fF
C3160 a_7894_5142# vcm 0.18fF
C3161 a_10998_4138# col_n[8] 0.34fF
C3162 a_21038_16186# col_n[18] 0.34fF
C3163 a_29374_15222# vcm 0.24fF
C3164 a_2475_18218# a_35002_18194# 0.41fF
C3165 m3_1046_19620# VDD 0.24fF
C3166 a_31078_17190# row_n[15] 0.43fF
C3167 a_7986_9158# ctop 4.91fF
C3168 a_16930_14178# VDD 0.29fF
C3169 m2_34864_15002# row_n[13] 0.38fF
C3170 m2_1732_946# sample_n 0.12fF
C3171 a_2275_9182# col_n[3] 0.17fF
C3172 a_7894_2130# rowon_n[0] 0.14fF
C3173 col_n[23] rowoff_n[14] 0.17fF
C3174 a_2275_15206# a_25054_15182# 0.71fF
C3175 a_22954_9158# vcm 0.18fF
C3176 m2_17796_18014# col_n[15] 0.34fF
C3177 col[26] rowoff_n[10] 0.17fF
C3178 a_17934_16186# rowoff_n[14] 0.57fF
C3179 a_20034_3134# a_21038_3134# 0.86fF
C3180 a_7986_8154# m2_8184_8402# 0.19fF
C3181 a_10298_18234# vcm 0.25fF
C3182 a_31078_3134# col[28] 0.38fF
C3183 a_23046_13174# ctop 4.91fF
C3184 a_31990_18194# VDD 0.50fF
C3185 a_2475_12194# a_17934_12170# 0.41fF
C3186 a_2275_12194# a_15318_12210# 0.15fF
C3187 a_9902_12170# a_9994_12170# 0.45fF
C3188 a_2475_16210# col[8] 0.22fF
C3189 a_18026_15182# rowon_n[13] 0.45fF
C3190 a_27062_4138# m2_27260_4386# 0.19fF
C3191 m2_31852_18014# m2_32280_18442# 0.19fF
C3192 a_2475_5166# col[13] 0.22fF
C3193 a_26362_3174# col_n[23] 0.11fF
C3194 a_34090_3134# VDD 1.23fF
C3195 a_10998_5142# a_10998_4138# 0.84fF
C3196 a_9994_14178# col_n[7] 0.34fF
C3197 a_28066_5142# rowon_n[3] 0.45fF
C3198 a_2275_9182# a_8898_9158# 0.17fF
C3199 rowon_n[8] ctop 0.37fF
C3200 a_3970_16186# ctop 4.91fF
C3201 col_n[7] rowoff_n[15] 0.29fF
C3202 col_n[20] col[20] 0.50fF
C3203 a_2475_18218# m2_18800_18014# 0.62fF
C3204 a_2475_14202# a_32994_14178# 0.41fF
C3205 a_2275_14202# a_30378_14218# 0.15fF
C3206 a_2275_11190# col_n[20] 0.17fF
C3207 a_2966_3134# rowoff_n[1] 2.62fF
C3208 col[10] rowoff_n[11] 0.28fF
C3209 a_18938_16186# vcm 0.18fF
C3210 a_15014_6146# VDD 3.20fF
C3211 a_5978_5142# row_n[3] 0.43fF
C3212 a_5886_9158# rowon_n[7] 0.14fF
C3213 a_20034_1126# col[17] 0.53fF
C3214 a_2275_8178# col[10] 0.17fF
C3215 a_34394_15222# col_n[31] 0.11fF
C3216 a_2275_11190# a_23958_11166# 0.17fF
C3217 a_30074_13174# col[27] 0.38fF
C3218 a_21038_1126# vcm 0.15fF
C3219 a_24962_16186# a_25054_16186# 0.45fF
C3220 a_5886_17190# rowoff_n[15] 0.70fF
C3221 m2_12776_18014# VDD 4.20fF
C3222 a_2475_7174# col[30] 0.22fF
C3223 a_3970_6146# rowoff_n[4] 2.57fF
C3224 a_30074_10162# VDD 1.65fF
C3225 a_15318_1166# col_n[12] 0.11fF
C3226 a_2475_8178# a_16018_8154# 0.68fF
C3227 a_26058_9158# a_26058_8154# 0.84fF
C3228 a_25358_13214# col_n[22] 0.11fF
C3229 ctop rowoff_n[12] 0.28fF
C3230 a_2475_4162# vcm 1.32fF
C3231 a_13006_4138# rowoff_n[2] 2.13fF
C3232 a_30074_12170# rowoff_n[10] 1.30fF
C3233 a_26058_12170# rowon_n[10] 0.45fF
C3234 a_2275_5166# a_6982_5142# 0.71fF
C3235 a_10998_13174# VDD 3.61fF
C3236 a_2275_18218# a_3878_18194# 0.17fF
C3237 a_2475_10186# a_31078_10162# 0.68fF
C3238 a_16018_10162# a_17022_10162# 0.86fF
C3239 a_2275_10186# col[27] 0.17fF
C3240 a_22042_2130# rowoff_n[0] 1.69fF
C3241 a_19030_11166# col[16] 0.38fF
C3242 a_17022_8154# vcm 0.89fF
C3243 a_3970_12170# row_n[10] 0.43fF
C3244 a_35002_3134# a_35094_3134# 0.11fF
C3245 m2_10768_18014# m3_10900_18146# 4.43fF
C3246 a_2275_7174# VDD 3.18fF
C3247 a_34090_7150# col_n[31] 0.34fF
C3248 a_2275_7174# a_22042_7150# 0.71fF
C3249 a_26058_17190# VDD 2.06fF
C3250 a_14010_2130# row_n[0] 0.43fF
C3251 a_6982_12170# a_6982_11166# 0.84fF
C3252 a_13918_6146# rowon_n[4] 0.14fF
C3253 a_14314_11206# col_n[11] 0.11fF
C3254 a_7286_2170# vcm 0.24fF
C3255 a_32082_12170# vcm 0.89fF
C3256 a_2275_4162# row_n[2] 26.41fF
C3257 a_28978_2130# VDD 0.29fF
C3258 a_2966_10162# m2_1732_9982# 0.86fF
C3259 a_2275_4162# a_12306_4178# 0.15fF
C3260 a_2475_4162# a_14922_4138# 0.41fF
C3261 m2_1732_8978# rowoff_n[7] 2.46fF
C3262 m3_1864_5094# m3_1864_4090# 0.20fF
C3263 m2_4744_946# col[2] 0.51fF
C3264 a_2475_14202# col[2] 0.22fF
C3265 a_2475_3158# col[7] 0.22fF
C3266 a_31078_14178# a_32082_14178# 0.86fF
C3267 a_14922_10162# rowoff_n[8] 0.60fF
C3268 a_22346_6186# vcm 0.24fF
C3269 a_18026_13174# rowoff_n[11] 1.89fF
C3270 a_7986_9158# col[5] 0.38fF
C3271 a_2275_1150# a_5886_1126# 0.17fF
C3272 a_13006_15182# vcm 0.89fF
C3273 a_9902_5142# VDD 0.29fF
C3274 a_15926_6146# a_16018_6146# 0.45fF
C3275 a_2275_13198# m2_34864_12994# 0.51fF
C3276 a_2475_6170# a_29982_6146# 0.41fF
C3277 a_2275_6170# a_27366_6186# 0.15fF
C3278 a_2275_9182# col_n[14] 0.17fF
C3279 a_34090_9158# rowon_n[7] 0.45fF
C3280 rowon_n[14] rowoff_n[14] 20.66fF
C3281 a_23958_8154# rowoff_n[6] 0.50fF
C3282 a_23046_5142# col_n[20] 0.34fF
C3283 a_33086_17190# col_n[30] 0.34fF
C3284 a_2475_15206# a_7986_15182# 0.68fF
C3285 a_22042_16186# a_22042_15182# 0.84fF
C3286 a_3270_9198# vcm 0.24fF
C3287 a_34090_17190# rowoff_n[15] 1.10fF
C3288 a_2275_6170# col[4] 0.17fF
C3289 a_2275_3158# a_20946_3134# 0.17fF
C3290 a_32994_6146# rowoff_n[4] 0.40fF
C3291 a_16018_4138# ctop 4.91fF
C3292 a_2275_1150# m2_21812_946# 0.51fF
C3293 a_8898_1126# m2_8760_946# 0.31fF
C3294 m3_24956_1078# ctop 0.21fF
C3295 a_24962_9158# VDD 0.29fF
C3296 a_12002_9158# row_n[7] 0.43fF
C3297 a_11910_13174# rowon_n[11] 0.14fF
C3298 a_2475_16210# col[19] 0.22fF
C3299 a_2475_5166# col[24] 0.22fF
C3300 a_30986_4138# vcm 0.18fF
C3301 a_21950_3134# rowon_n[1] 0.14fF
C3302 a_12002_17190# a_13006_17190# 0.86fF
C3303 a_2475_17214# a_23046_17190# 0.68fF
C3304 m2_13780_18014# m2_14784_18014# 0.86fF
C3305 a_18330_13214# vcm 0.24fF
C3306 col_n[18] rowoff_n[15] 0.21fF
C3307 col_n[25] col[26] 6.11fF
C3308 row_n[3] ctop 0.28fF
C3309 a_2275_5166# a_34394_5182# 0.15fF
C3310 a_35002_12170# m2_34864_11990# 0.33fF
C3311 a_31078_8154# ctop 4.91fF
C3312 a_5886_12170# VDD 0.29fF
C3313 a_2275_11190# col_n[31] 0.17fF
C3314 a_30986_10162# a_31078_10162# 0.45fF
C3315 col[21] rowoff_n[11] 0.21fF
C3316 m2_1732_8978# vcm 1.11fF
C3317 a_2275_14202# a_14010_14178# 0.71fF
C3318 a_12002_3134# col_n[9] 0.34fF
C3319 a_11910_7150# vcm 0.18fF
C3320 a_22042_15182# col_n[19] 0.34fF
C3321 a_5978_14178# rowoff_n[12] 2.47fF
C3322 a_32082_3134# a_32082_2130# 0.84fF
C3323 a_2475_2154# a_28066_2130# 0.68fF
C3324 a_33390_17230# vcm 0.24fF
C3325 a_2275_8178# col[21] 0.17fF
C3326 a_32082_16186# rowon_n[14] 0.45fF
C3327 a_12002_11166# ctop 4.91fF
C3328 a_20946_16186# VDD 0.29fF
C3329 a_2475_11190# a_6890_11166# 0.41fF
C3330 a_2275_11190# a_4274_11206# 0.15fF
C3331 a_2966_1126# vcm 0.15fF
C3332 a_2275_16210# a_29070_16186# 0.71fF
C3333 m2_34864_15002# m2_35292_15430# 0.19fF
C3334 a_3970_2130# m2_2736_1950# 0.86fF
C3335 a_26970_11166# vcm 0.18fF
C3336 a_23046_1126# VDD 0.11fF
C3337 a_9994_16186# row_n[14] 0.43fF
C3338 a_32082_2130# col[29] 0.38fF
C3339 a_22042_4138# a_23046_4138# 0.86fF
C3340 col[5] rowoff_n[12] 0.31fF
C3341 a_13006_17190# m2_13204_17438# 0.19fF
C3342 a_27062_15182# ctop 4.91fF
C3343 a_20034_6146# row_n[4] 0.43fF
C3344 a_2275_13198# a_19334_13214# 0.15fF
C3345 a_2475_13198# a_21950_13174# 0.41fF
C3346 a_11910_13174# a_12002_13174# 0.45fF
C3347 a_19942_10162# rowon_n[8] 0.14fF
C3348 m2_15788_946# vcm 0.71fF
C3349 a_27366_2170# col_n[24] 0.11fF
C3350 a_2275_1150# a_35094_1126# 0.14fF
C3351 a_7894_14178# vcm 0.18fF
C3352 a_10998_13174# col_n[8] 0.34fF
C3353 a_3970_4138# VDD 4.33fF
C3354 a_32082_13174# m2_32280_13422# 0.19fF
C3355 a_13006_6146# a_13006_5142# 0.84fF
C3356 a_2475_1150# col[1] 0.22fF
C3357 a_2275_10186# a_12914_10162# 0.17fF
C3358 a_2275_15206# a_35398_15222# 0.15fF
C3359 a_2275_7174# col_n[8] 0.17fF
C3360 a_6982_4138# rowon_n[2] 0.45fF
C3361 a_22954_18194# vcm 0.18fF
C3362 a_19030_8154# VDD 2.78fF
C3363 a_3970_15182# m2_4168_15430# 0.19fF
C3364 a_2475_7174# a_4974_7150# 0.68fF
C3365 a_31078_12170# col[28] 0.38fF
C3366 a_2275_12194# a_27974_12170# 0.17fF
C3367 a_25054_3134# vcm 0.89fF
C3368 a_26970_17190# a_27062_17190# 0.45fF
C3369 m2_32856_18014# col[30] 0.37fF
C3370 a_4974_5142# rowoff_n[3] 2.52fF
C3371 a_23046_11166# m2_23244_11414# 0.19fF
C3372 a_2475_14202# col[13] 0.22fF
C3373 a_18026_13174# row_n[11] 0.43fF
C3374 a_34090_12170# VDD 1.23fF
C3375 a_26362_12210# col_n[23] 0.11fF
C3376 a_2475_3158# col[18] 0.22fF
C3377 m3_24956_18146# m3_25960_18146# 0.21fF
C3378 m2_16792_946# m3_16924_1078# 4.41fF
C3379 a_2475_9182# a_20034_9158# 0.68fF
C3380 a_28066_10162# a_28066_9158# 0.84fF
C3381 a_17934_17190# rowon_n[15] 0.14fF
C3382 a_2475_18218# col[4] 0.22fF
C3383 a_28066_3134# row_n[1] 0.43fF
C3384 a_14010_3134# rowoff_n[1] 2.08fF
C3385 a_27974_7150# rowon_n[5] 0.14fF
C3386 a_5978_6146# vcm 0.89fF
C3387 a_35002_14178# rowoff_n[12] 0.38fF
C3388 a_2275_9182# col_n[25] 0.17fF
C3389 a_2275_6170# a_10998_6146# 0.71fF
C3390 a_15014_15182# VDD 3.20fF
C3391 a_18026_11166# a_19030_11166# 0.86fF
C3392 a_20034_10162# col[17] 0.38fF
C3393 a_2275_17214# col[10] 0.17fF
C3394 a_30378_1166# vcm 0.25fF
C3395 a_2275_6170# col[15] 0.17fF
C3396 a_4974_11166# rowon_n[9] 0.45fF
C3397 a_21038_10162# vcm 0.89fF
C3398 a_14010_9158# m2_14208_9406# 0.19fF
C3399 m3_20940_18146# ctop 0.21fF
C3400 a_2475_16210# col[30] 0.22fF
C3401 a_2275_8178# a_26058_8154# 0.71fF
C3402 a_15318_10202# col_n[12] 0.11fF
C3403 a_8990_13174# a_8990_12170# 0.84fF
C3404 a_11302_4178# vcm 0.24fF
C3405 a_3878_3134# rowon_n[1] 0.14fF
C3406 a_2966_17190# a_3970_17190# 0.86fF
C3407 a_2275_17214# a_4882_17190# 0.17fF
C3408 a_6890_11166# rowoff_n[9] 0.69fF
C3409 col_n[29] rowoff_n[15] 0.13fF
C3410 col_n[31] col[31] 0.69fF
C3411 m2_34864_17010# rowon_n[15] 0.42fF
C3412 a_33086_5142# m2_33284_5390# 0.19fF
C3413 a_2475_13198# vcm 1.32fF
C3414 a_32994_4138# VDD 0.29fF
C3415 a_2475_5166# a_18938_5142# 0.41fF
C3416 a_2275_5166# a_16322_5182# 0.15fF
C3417 sample_n rowoff_n[11] 0.55fF
C3418 a_2275_18218# a_14922_18194# 0.17fF
C3419 a_26058_10162# row_n[8] 0.43fF
C3420 a_15926_9158# rowoff_n[7] 0.59fF
C3421 a_25966_14178# rowon_n[12] 0.14fF
C3422 a_33086_15182# a_34090_15182# 0.86fF
C3423 a_26362_8194# vcm 0.24fF
C3424 a_8990_8154# col[6] 0.38fF
C3425 a_22954_15182# rowoff_n[13] 0.51fF
C3426 a_2275_2154# a_9902_2130# 0.17fF
C3427 a_4974_7150# m2_5172_7398# 0.19fF
C3428 a_17022_17190# vcm 0.89fF
C3429 a_4974_2130# ctop 4.93fF
C3430 a_13918_7150# VDD 0.29fF
C3431 a_24962_7150# rowoff_n[5] 0.49fF
C3432 a_2475_7174# a_33998_7150# 0.41fF
C3433 a_2275_7174# a_31382_7190# 0.15fF
C3434 a_17934_7150# a_18026_7150# 0.45fF
C3435 a_24050_4138# col_n[21] 0.34fF
C3436 a_2275_16210# VDD 3.18fF
C3437 a_34090_16186# col_n[31] 0.34fF
C3438 a_2275_5166# col_n[2] 0.17fF
C3439 a_19942_2130# vcm 0.18fF
C3440 a_4274_8194# col_n[1] 0.11fF
C3441 a_24050_17190# a_24050_16186# 0.84fF
C3442 a_2475_16210# a_12002_16186# 0.68fF
C3443 a_24050_3134# m2_24248_3382# 0.19fF
C3444 a_33998_5142# rowoff_n[3] 0.39fF
C3445 a_7286_11206# vcm 0.24fF
C3446 a_5374_1488# VDD 0.18fF
C3447 a_13006_8154# rowon_n[6] 0.45fF
C3448 col[16] rowoff_n[12] 0.24fF
C3449 a_2275_4162# a_24962_4138# 0.17fF
C3450 a_20034_6146# ctop 4.91fF
C3451 a_28978_11166# VDD 0.29fF
C3452 m3_14916_1078# m3_15920_1078# 0.21fF
C3453 a_1957_6170# row_n[4] 0.29fF
C3454 a_2475_13198# a_3878_13174# 0.41fF
C3455 a_2275_13198# a_2874_13174# 0.17fF
C3456 a_35002_6146# vcm 0.18fF
C3457 a_2475_12194# col[7] 0.22fF
C3458 a_2475_1150# col[12] 0.22fF
C3459 a_22346_15222# vcm 0.24fF
C3460 a_2475_18218# a_27974_18194# 0.41fF
C3461 a_24050_17190# row_n[15] 0.43fF
C3462 a_9902_14178# VDD 0.29fF
C3463 a_32994_11166# a_33086_11166# 0.45fF
C3464 a_13006_2130# col_n[10] 0.34fF
C3465 a_2275_7174# col_n[19] 0.17fF
C3466 a_23046_14178# col_n[20] 0.34fF
C3467 a_2275_15206# a_18026_15182# 0.71fF
C3468 a_34090_7150# row_n[5] 0.43fF
C3469 a_33998_11166# rowon_n[9] 0.14fF
C3470 a_15926_9158# vcm 0.18fF
C3471 a_10906_16186# rowoff_n[14] 0.65fF
C3472 col[0] rowoff_n[13] 0.34fF
C3473 a_2275_8178# m2_1732_7974# 0.27fF
C3474 a_2475_3158# a_32082_3134# 0.68fF
C3475 a_34090_4138# a_34090_3134# 0.84fF
C3476 a_3270_18234# vcm 0.25fF
C3477 a_35494_9520# VDD 0.13fF
C3478 a_2275_15206# col[4] 0.17fF
C3479 a_16018_13174# ctop 4.91fF
C3480 a_2275_4162# col[9] 0.17fF
C3481 a_24962_18194# VDD 0.50fF
C3482 a_2475_12194# a_10906_12170# 0.41fF
C3483 a_2275_12194# a_8290_12210# 0.15fF
C3484 a_2275_17214# a_33086_17190# 0.71fF
C3485 a_10998_15182# rowon_n[13] 0.45fF
C3486 m2_24824_18014# m2_25252_18442# 0.19fF
C3487 a_2475_14202# col[24] 0.22fF
C3488 a_30986_13174# vcm 0.18fF
C3489 a_27062_3134# VDD 1.96fF
C3490 a_2475_3158# col[29] 0.22fF
C3491 a_24050_5142# a_25054_5142# 0.86fF
C3492 a_2475_18218# col[15] 0.22fF
C3493 a_21038_5142# rowon_n[3] 0.45fF
C3494 a_31078_17190# ctop 4.93fF
C3495 a_2475_18218# m2_4744_18014# 0.62fF
C3496 a_2475_14202# a_25966_14178# 0.41fF
C3497 a_2275_14202# a_23350_14218# 0.15fF
C3498 a_13918_14178# a_14010_14178# 0.45fF
C3499 a_28370_1166# col_n[25] 0.11fF
C3500 a_12002_12170# col_n[9] 0.34fF
C3501 a_11910_16186# vcm 0.18fF
C3502 a_7986_6146# VDD 3.92fF
C3503 a_15014_7150# a_15014_6146# 0.84fF
C3504 a_2275_17214# col[21] 0.17fF
C3505 a_2275_6170# col[26] 0.17fF
C3506 a_32082_14178# row_n[12] 0.43fF
C3507 a_2275_11190# a_16930_11166# 0.17fF
C3508 a_2275_18218# col[6] 0.17fF
C3509 m2_30848_946# col_n[28] 0.48fF
C3510 a_14010_1126# vcm 0.15fF
C3511 a_2966_10162# vcm 0.89fF
C3512 a_34090_10162# m2_34864_9982# 0.86fF
C3513 a_32082_11166# col[29] 0.38fF
C3514 a_23046_10162# VDD 2.37fF
C3515 a_2475_8178# a_8990_8154# 0.68fF
C3516 a_4974_8154# a_5978_8154# 0.86fF
C3517 a_2275_13198# a_31990_13174# 0.17fF
C3518 ctop col[7] 0.13fF
C3519 row_n[11] sample_n 0.16fF
C3520 a_29070_5142# vcm 0.89fF
C3521 a_5978_4138# rowoff_n[2] 2.47fF
C3522 a_23046_12170# rowoff_n[10] 1.64fF
C3523 a_28978_18194# a_29070_18194# 0.11fF
C3524 a_23958_1126# a_24050_1126# 0.11fF
C3525 a_19030_12170# rowon_n[10] 0.45fF
C3526 a_27366_11206# col_n[24] 0.11fF
C3527 a_3970_13174# VDD 4.33fF
C3528 a_2475_10186# a_24050_10162# 0.68fF
C3529 a_30074_11166# a_30074_10162# 0.84fF
C3530 a_2475_10186# col[1] 0.22fF
C3531 a_15014_2130# rowoff_n[0] 2.03fF
C3532 a_29070_2130# rowon_n[0] 0.45fF
C3533 a_9994_8154# vcm 0.89fF
C3534 a_2275_16210# col_n[8] 0.17fF
C3535 a_2275_7174# a_15014_7150# 0.71fF
C3536 a_2275_5166# col_n[13] 0.17fF
C3537 a_6982_2130# row_n[0] 0.43fF
C3538 a_19030_17190# VDD 2.78fF
C3539 a_21038_9158# col[18] 0.38fF
C3540 a_20034_12170# a_21038_12170# 0.86fF
C3541 a_6890_6146# rowon_n[4] 0.14fF
C3542 a_35398_3174# vcm 0.24fF
C3543 col[27] rowoff_n[12] 0.17fF
C3544 a_3270_5182# col_n[0] 0.11fF
C3545 a_25054_12170# vcm 0.89fF
C3546 a_21950_2130# VDD 0.29fF
C3547 a_2275_2154# col[3] 0.17fF
C3548 a_4882_4138# a_4974_4138# 0.45fF
C3549 a_2475_4162# a_7894_4138# 0.41fF
C3550 a_2275_4162# a_5278_4178# 0.15fF
C3551 m3_1864_12122# m3_1864_11118# 0.20fF
C3552 a_16322_9198# col_n[13] 0.11fF
C3553 a_2275_9182# a_30074_9158# 0.71fF
C3554 a_21950_18194# m2_21812_18014# 0.34fF
C3555 a_2475_12194# col[18] 0.22fF
C3556 a_10998_14178# a_10998_13174# 0.84fF
C3557 a_7894_10162# rowoff_n[8] 0.68fF
C3558 a_2475_1150# col[23] 0.22fF
C3559 a_15318_6186# vcm 0.24fF
C3560 a_10998_13174# rowoff_n[11] 2.23fF
C3561 a_5978_15182# vcm 0.89fF
C3562 a_2161_5166# VDD 0.23fF
C3563 a_2475_6170# a_22954_6146# 0.41fF
C3564 a_2275_6170# a_20338_6186# 0.15fF
C3565 a_27062_9158# rowon_n[7] 0.45fF
C3566 a_16930_8154# rowoff_n[6] 0.58fF
C3567 a_2275_7174# col_n[30] 0.17fF
C3568 col[11] rowoff_n[13] 0.27fF
C3569 a_9994_7150# col[7] 0.38fF
C3570 a_30378_10202# vcm 0.24fF
C3571 a_27062_17190# rowoff_n[15] 1.45fF
C3572 a_2275_15206# col[15] 0.17fF
C3573 a_25966_6146# rowoff_n[4] 0.48fF
C3574 a_2275_3158# a_13918_3134# 0.17fF
C3575 a_2275_4162# col[20] 0.17fF
C3576 a_8990_4138# ctop 4.91fF
C3577 a_2475_1150# m2_7756_946# 0.62fF
C3578 a_25054_3134# col_n[22] 0.34fF
C3579 a_17934_9158# VDD 0.29fF
C3580 m3_1864_3086# ctop 0.22fF
C3581 a_4974_9158# row_n[7] 0.43fF
C3582 a_9994_16186# m2_10192_16434# 0.19fF
C3583 a_19942_8154# a_20034_8154# 0.45fF
C3584 a_4882_13174# rowon_n[11] 0.14fF
C3585 a_5278_7190# col_n[2] 0.11fF
C3586 a_23958_4138# vcm 0.18fF
C3587 a_35002_4138# rowoff_n[2] 0.38fF
C3588 a_14922_3134# rowon_n[1] 0.14fF
C3589 a_2475_17214# a_16018_17190# 0.68fF
C3590 m2_6752_18014# m2_7756_18014# 0.86fF
C3591 a_11302_13214# vcm 0.24fF
C3592 a_2475_18218# col[26] 0.22fF
C3593 a_2275_5166# a_28978_5142# 0.17fF
C3594 a_29070_12170# m2_29268_12418# 0.19fF
C3595 a_24050_8154# ctop 4.91fF
C3596 a_2966_5142# rowon_n[3] 0.45fF
C3597 a_32994_13174# VDD 0.29fF
C3598 a_2275_14202# a_6982_14178# 0.71fF
C3599 a_4882_7150# vcm 0.18fF
C3600 a_10998_2130# a_12002_2130# 0.86fF
C3601 a_2475_2154# a_21038_2130# 0.68fF
C3602 a_8990_17190# col[6] 0.38fF
C3603 a_26362_17230# vcm 0.24fF
C3604 a_25054_16186# rowon_n[14] 0.45fF
C3605 a_4974_11166# ctop 4.91fF
C3606 a_2275_18218# col[17] 0.17fF
C3607 a_13918_16186# VDD 0.29fF
C3608 a_35002_12170# a_35094_12170# 0.11fF
C3609 a_24050_13174# col_n[21] 0.34fF
C3610 a_2275_16210# a_22042_16186# 0.71fF
C3611 a_2275_14202# col_n[2] 0.17fF
C3612 a_19942_11166# vcm 0.18fF
C3613 a_2275_3158# col_n[7] 0.17fF
C3614 a_4274_17230# col_n[1] 0.11fF
C3615 a_16018_1126# VDD 0.12fF
C3616 a_1957_7174# sample 0.35fF
C3617 a_20034_10162# m2_20232_10410# 0.19fF
C3618 m2_34864_5966# row_n[4] 0.38fF
C3619 ctop col[18] 0.13fF
C3620 rowon_n[5] sample_n 0.15fF
C3621 a_18026_17190# m2_17796_18014# 0.84fF
C3622 a_20034_15182# ctop 4.91fF
C3623 a_13006_6146# row_n[4] 0.43fF
C3624 a_12914_10162# rowon_n[8] 0.14fF
C3625 a_2475_13198# a_14922_13174# 0.41fF
C3626 a_2275_13198# a_12306_13214# 0.15fF
C3627 m2_34864_4962# m2_34864_3958# 0.84fF
C3628 a_2275_1150# a_27062_1126# 0.14fF
C3629 a_35002_15182# vcm 0.18fF
C3630 a_31078_5142# VDD 1.54fF
C3631 a_2475_10186# col[12] 0.22fF
C3632 a_26058_6146# a_27062_6146# 0.86fF
C3633 m2_2736_946# m2_3164_1374# 0.19fF
C3634 a_2275_10186# a_5886_10162# 0.17fF
C3635 a_15926_15182# a_16018_15182# 0.45fF
C3636 a_2275_15206# a_27366_15222# 0.15fF
C3637 a_2475_15206# a_29982_15182# 0.41fF
C3638 a_13006_11166# col_n[10] 0.34fF
C3639 a_2275_16210# col_n[19] 0.17fF
C3640 a_2275_5166# col_n[24] 0.17fF
C3641 a_10998_8154# m2_11196_8402# 0.19fF
C3642 a_15926_18194# vcm 0.18fF
C3643 a_12002_8154# VDD 3.51fF
C3644 a_17022_8154# a_17022_7150# 0.84fF
C3645 a_33086_13174# rowon_n[11] 0.45fF
C3646 a_35494_18556# VDD 0.13fF
C3647 a_2275_12194# a_20946_12170# 0.17fF
C3648 a_2275_13198# col[9] 0.17fF
C3649 a_18026_3134# vcm 0.89fF
C3650 a_2275_2154# col[14] 0.17fF
C3651 a_30074_4138# m2_30272_4386# 0.19fF
C3652 a_3878_2130# VDD 0.29fF
C3653 a_33086_10162# col[30] 0.38fF
C3654 a_10998_13174# row_n[11] 0.43fF
C3655 a_2475_12194# col[29] 0.22fF
C3656 a_27062_12170# VDD 1.96fF
C3657 m3_10900_18146# m3_11904_18146# 0.21fF
C3658 a_2475_9182# a_13006_9158# 0.68fF
C3659 a_10906_17190# rowon_n[15] 0.14fF
C3660 a_6982_9158# a_7986_9158# 0.86fF
C3661 a_2275_14202# a_34394_14218# 0.15fF
C3662 a_21038_3134# row_n[1] 0.43fF
C3663 a_6982_3134# rowoff_n[1] 2.42fF
C3664 a_33086_7150# vcm 0.89fF
C3665 a_20946_7150# rowon_n[5] 0.14fF
C3666 a_27974_14178# rowoff_n[12] 0.46fF
C3667 a_28370_10202# col_n[25] 0.11fF
C3668 a_1957_6170# m2_1732_5966# 0.33fF
C3669 a_25966_2130# a_26058_2130# 0.45fF
C3670 a_2275_6170# a_3970_6146# 0.71fF
C3671 col[22] rowoff_n[13] 0.20fF
C3672 a_7986_15182# VDD 3.92fF
C3673 a_2475_11190# a_28066_11166# 0.68fF
C3674 a_32082_12170# a_32082_11166# 0.84fF
C3675 col_n[2] rowoff_n[6] 0.32fF
C3676 sample rowoff_n[2] 0.22fF
C3677 a_23350_1166# vcm 0.25fF
C3678 col_n[5] rowoff_n[9] 0.30fF
C3679 col_n[0] rowoff_n[3] 0.34fF
C3680 col_n[1] rowoff_n[5] 0.33fF
C3681 col_n[3] rowoff_n[7] 0.32fF
C3682 VDD rowoff_n[1] 87.22fF
C3683 vcm rowoff_n[4] 2.43fF
C3684 col_n[4] rowoff_n[8] 0.31fF
C3685 a_2275_15206# col[26] 0.17fF
C3686 a_2275_4162# col[31] 0.17fF
C3687 a_14010_10162# vcm 0.89fF
C3688 a_22042_8154# col[19] 0.38fF
C3689 a_2275_8178# a_19030_8154# 0.71fF
C3690 a_22042_13174# a_23046_13174# 0.86fF
C3691 a_2275_1150# col_n[1] 0.14fF
C3692 m2_11772_18014# col_n[9] 0.33fF
C3693 m2_1732_1950# m2_2736_1950# 0.86fF
C3694 a_4274_4178# vcm 0.24fF
C3695 a_29070_14178# vcm 0.89fF
C3696 a_25966_4138# VDD 0.29fF
C3697 a_2475_5166# a_11910_5142# 0.41fF
C3698 a_2275_5166# a_9294_5182# 0.15fF
C3699 a_6890_5142# a_6982_5142# 0.45fF
C3700 col[6] rowoff_n[14] 0.31fF
C3701 a_17326_8194# col_n[14] 0.11fF
C3702 a_2275_18218# a_7894_18194# 0.17fF
C3703 a_2275_10186# a_34090_10162# 0.71fF
C3704 a_19030_10162# row_n[8] 0.43fF
C3705 a_8898_9158# rowoff_n[7] 0.67fF
C3706 a_18938_14178# rowon_n[12] 0.14fF
C3707 a_13006_15182# a_13006_14178# 0.84fF
C3708 a_19334_8194# vcm 0.24fF
C3709 a_2475_8178# col[6] 0.22fF
C3710 a_15926_15182# rowoff_n[13] 0.59fF
C3711 a_2275_18218# col[28] 0.17fF
C3712 a_28978_4138# rowon_n[2] 0.14fF
C3713 a_2161_2154# a_2275_2154# 0.17fF
C3714 a_32082_3134# ctop 4.91fF
C3715 a_9994_17190# vcm 0.89fF
C3716 m2_15788_18014# m3_15920_18146# 4.41fF
C3717 a_6890_7150# VDD 0.29fF
C3718 a_17934_7150# rowoff_n[5] 0.57fF
C3719 a_2475_7174# a_26970_7150# 0.41fF
C3720 a_2275_7174# a_24354_7190# 0.15fF
C3721 a_2275_14202# col_n[13] 0.17fF
C3722 a_10998_6146# col[8] 0.38fF
C3723 a_2275_3158# col_n[18] 0.17fF
C3724 a_12914_2130# vcm 0.18fF
C3725 a_2475_16210# a_4974_16186# 0.68fF
C3726 m2_1732_11990# sample 0.31fF
C3727 a_35398_12210# vcm 0.24fF
C3728 a_26970_5142# rowoff_n[3] 0.47fF
C3729 VDD col_n[6] 14.95fF
C3730 vcm col_n[3] 3.22fF
C3731 a_26058_2130# col_n[23] 0.34fF
C3732 ctop col[29] 0.13fF
C3733 row_n[0] sample_n 0.16fF
C3734 a_5978_8154# rowon_n[6] 0.45fF
C3735 a_3270_14218# col_n[0] 0.11fF
C3736 a_2275_4162# a_17934_4138# 0.17fF
C3737 a_13006_6146# ctop 4.91fF
C3738 a_2275_11190# col[3] 0.17fF
C3739 a_21950_11166# VDD 0.29fF
C3740 m3_2868_2082# m3_2868_1078# 0.20fF
C3741 a_21950_9158# a_22042_9158# 0.45fF
C3742 a_6282_6186# col_n[3] 0.11fF
C3743 a_16322_18234# col_n[13] 0.11fF
C3744 a_19030_1126# en_bit_n[2] 0.28fF
C3745 a_27974_6146# vcm 0.18fF
C3746 a_2475_10186# col[23] 0.22fF
C3747 a_15318_15222# vcm 0.24fF
C3748 a_2475_18218# a_20946_18194# 0.41fF
C3749 m2_5748_946# VDD 6.85fF
C3750 a_2275_6170# a_32994_6146# 0.17fF
C3751 a_28066_10162# ctop 4.91fF
C3752 a_17022_17190# row_n[15] 0.43fF
C3753 a_2161_14202# VDD 0.23fF
C3754 a_2275_16210# col_n[30] 0.17fF
C3755 a_27062_7150# row_n[5] 0.43fF
C3756 a_2275_15206# a_10998_15182# 0.71fF
C3757 a_26970_11166# rowon_n[9] 0.14fF
C3758 a_8898_9158# vcm 0.18fF
C3759 a_9994_16186# col[7] 0.38fF
C3760 a_2475_3158# a_25054_3134# 0.68fF
C3761 a_13006_3134# a_14010_3134# 0.86fF
C3762 a_2475_1150# m2_30848_946# 0.62fF
C3763 a_8990_13174# ctop 4.91fF
C3764 a_2275_13198# col[20] 0.17fF
C3765 a_25054_12170# col_n[22] 0.34fF
C3766 a_17934_18194# VDD 0.50fF
C3767 a_2275_2154# col[25] 0.17fF
C3768 a_28066_11166# rowoff_n[9] 1.40fF
C3769 a_2275_17214# a_26058_17190# 0.71fF
C3770 a_5278_16226# col_n[2] 0.11fF
C3771 a_3970_15182# rowon_n[13] 0.45fF
C3772 m2_17796_18014# m2_18224_18442# 0.19fF
C3773 a_2966_6146# col_n[0] 0.34fF
C3774 a_23958_13174# vcm 0.18fF
C3775 a_20034_3134# VDD 2.68fF
C3776 a_2966_11166# m2_3164_11414# 0.19fF
C3777 a_3970_5142# a_3970_4138# 0.84fF
C3778 a_14010_5142# rowon_n[3] 0.45fF
C3779 a_24050_17190# ctop 4.93fF
C3780 a_2475_14202# a_18938_14178# 0.41fF
C3781 a_2275_14202# a_16322_14218# 0.15fF
C3782 a_2966_3134# row_n[1] 0.41fF
C3783 a_2275_7174# rowon_n[5] 1.99fF
C3784 a_2275_2154# a_31078_2130# 0.71fF
C3785 a_4882_16186# vcm 0.18fF
C3786 a_28066_7150# a_29070_7150# 0.86fF
C3787 col_n[7] rowoff_n[0] 0.29fF
C3788 col_n[10] rowoff_n[3] 0.27fF
C3789 col_n[13] rowoff_n[6] 0.24fF
C3790 col_n[16] rowoff_n[9] 0.22fF
C3791 col_n[11] rowoff_n[4] 0.26fF
C3792 col_n[14] rowoff_n[7] 0.24fF
C3793 col_n[8] rowoff_n[1] 0.28fF
C3794 col_n[15] rowoff_n[8] 0.23fF
C3795 col_n[12] rowoff_n[5] 0.25fF
C3796 col_n[9] rowoff_n[2] 0.27fF
C3797 a_2275_11190# a_9902_11166# 0.17fF
C3798 a_2475_6170# col[0] 0.20fF
C3799 a_25054_14178# row_n[12] 0.43fF
C3800 a_14010_10162# col_n[11] 0.34fF
C3801 a_6982_1126# vcm 0.15fF
C3802 a_2275_16210# a_31382_16226# 0.15fF
C3803 a_2475_16210# a_33998_16186# 0.41fF
C3804 a_17934_16186# a_18026_16186# 0.45fF
C3805 a_35002_8154# rowon_n[6] 0.14fF
C3806 a_2275_12194# col_n[7] 0.17fF
C3807 a_16018_10162# VDD 3.09fF
C3808 a_2275_1150# col_n[12] 0.17fF
C3809 a_1957_16210# sample 0.35fF
C3810 a_16018_17190# m2_16216_17438# 0.19fF
C3811 a_19030_9158# a_19030_8154# 0.84fF
C3812 a_2275_13198# a_24962_13174# 0.17fF
C3813 a_22042_5142# vcm 0.89fF
C3814 a_16018_12170# rowoff_n[10] 1.98fF
C3815 m2_24824_946# vcm 0.71fF
C3816 a_2275_18218# m2_21812_18014# 0.51fF
C3817 col[17] rowoff_n[14] 0.23fF
C3818 a_34090_9158# col[31] 0.38fF
C3819 a_12002_12170# rowon_n[10] 0.45fF
C3820 vcm rowoff_n[10] 2.43fF
C3821 a_31078_14178# VDD 1.54fF
C3822 a_2475_10186# a_17022_10162# 0.68fF
C3823 a_8990_10162# a_9994_10162# 0.86fF
C3824 m2_14784_946# col_n[12] 0.45fF
C3825 a_7986_2130# rowoff_n[0] 2.38fF
C3826 a_22042_2130# rowon_n[0] 0.45fF
C3827 a_2475_8178# col[17] 0.22fF
C3828 a_2874_8154# vcm 0.18fF
C3829 a_29374_9198# col_n[26] 0.11fF
C3830 a_32082_16186# rowoff_n[14] 1.20fF
C3831 a_27974_3134# a_28066_3134# 0.45fF
C3832 a_30986_1126# m2_30848_946# 0.31fF
C3833 a_2275_14202# col_n[24] 0.17fF
C3834 a_6982_15182# m2_7180_15430# 0.19fF
C3835 a_2275_7174# a_7986_7150# 0.71fF
C3836 a_2275_3158# col_n[29] 0.17fF
C3837 a_12002_17190# VDD 3.51fF
C3838 a_34090_13174# a_34090_12170# 0.84fF
C3839 a_2475_12194# a_32082_12170# 0.68fF
C3840 a_27366_3174# vcm 0.24fF
C3841 a_33086_11166# row_n[9] 0.43fF
C3842 vcm col_n[14] 3.22fF
C3843 VDD col_n[17] 11.73fF
C3844 col[1] rowoff_n[15] 0.34fF
C3845 a_32994_15182# rowon_n[13] 0.14fF
C3846 a_18026_12170# vcm 0.89fF
C3847 a_2275_11190# col[14] 0.17fF
C3848 a_14922_2130# VDD 0.29fF
C3849 a_26058_11166# m2_26256_11414# 0.19fF
C3850 a_23046_7150# col[20] 0.38fF
C3851 a_3878_11166# VDD 0.29fF
C3852 m2_22816_946# m3_22948_1078# 4.41fF
C3853 a_2275_9182# a_23046_9158# 0.71fF
C3854 a_24050_14178# a_25054_14178# 0.86fF
C3855 a_8290_6186# vcm 0.24fF
C3856 a_3970_13174# rowoff_n[11] 2.57fF
C3857 a_33086_16186# vcm 0.89fF
C3858 a_18330_7190# col_n[15] 0.11fF
C3859 a_29982_6146# VDD 0.29fF
C3860 a_2475_6170# a_15926_6146# 0.41fF
C3861 a_2275_6170# a_13310_6186# 0.15fF
C3862 a_8898_6146# a_8990_6146# 0.45fF
C3863 m2_34864_946# col_n[31] 0.29fF
C3864 a_20034_9158# rowon_n[7] 0.45fF
C3865 a_9902_8154# rowoff_n[6] 0.66fF
C3866 a_15014_16186# a_15014_15182# 0.84fF
C3867 m2_34864_7974# rowon_n[6] 0.42fF
C3868 a_23350_10202# vcm 0.24fF
C3869 a_20034_17190# rowoff_n[15] 1.79fF
C3870 a_18938_6146# rowoff_n[4] 0.56fF
C3871 a_2275_13198# col[31] 0.17fF
C3872 a_17022_9158# m2_17220_9406# 0.19fF
C3873 a_2275_3158# a_6890_3134# 0.17fF
C3874 m3_1864_17142# ctop 0.22fF
C3875 a_10906_9158# VDD 0.29fF
C3876 a_2475_8178# a_30986_8154# 0.41fF
C3877 a_2275_8178# a_28370_8194# 0.15fF
C3878 a_12002_5142# col[9] 0.38fF
C3879 a_22042_17190# col[19] 0.38fF
C3880 a_16930_4138# vcm 0.18fF
C3881 a_2275_10186# col_n[1] 0.17fF
C3882 a_27974_4138# rowoff_n[2] 0.46fF
C3883 a_7894_3134# rowon_n[1] 0.14fF
C3884 a_2475_17214# a_8990_17190# 0.68fF
C3885 a_4974_17190# a_5978_17190# 0.86fF
C3886 a_4274_13214# vcm 0.24fF
C3887 a_1957_3158# VDD 0.28fF
C3888 a_2275_5166# a_21950_5142# 0.17fF
C3889 a_17022_8154# ctop 4.91fF
C3890 a_7286_5182# col_n[4] 0.11fF
C3891 a_25966_13174# VDD 0.29fF
C3892 a_23958_10162# a_24050_10162# 0.45fF
C3893 a_2966_3134# col[0] 0.38fF
C3894 a_17326_17230# col_n[14] 0.11fF
C3895 m2_26832_18014# col[24] 0.39fF
C3896 a_31990_8154# vcm 0.18fF
C3897 a_7986_7150# m2_8184_7398# 0.19fF
C3898 a_2475_2154# a_14010_2130# 0.68fF
C3899 a_25054_3134# a_25054_2130# 0.84fF
C3900 a_19334_17230# vcm 0.24fF
C3901 a_2475_17214# col[6] 0.22fF
C3902 col_n[19] rowoff_n[1] 0.20fF
C3903 col_n[22] rowoff_n[4] 0.18fF
C3904 col_n[25] rowoff_n[7] 0.16fF
C3905 col_n[18] rowoff_n[0] 0.21fF
C3906 col_n[26] rowoff_n[8] 0.15fF
C3907 col_n[23] rowoff_n[5] 0.17fF
C3908 col_n[20] rowoff_n[2] 0.19fF
C3909 col_n[27] rowoff_n[9] 0.14fF
C3910 col_n[24] rowoff_n[6] 0.16fF
C3911 col_n[21] rowoff_n[3] 0.19fF
C3912 a_18026_16186# rowon_n[14] 0.45fF
C3913 a_2475_6170# col[11] 0.22fF
C3914 a_32082_12170# ctop 4.91fF
C3915 a_6890_16186# VDD 0.29fF
C3916 a_28066_6146# rowon_n[4] 0.45fF
C3917 a_2275_16210# a_15014_16186# 0.71fF
C3918 a_10998_15182# col[8] 0.38fF
C3919 a_27062_3134# m2_27260_3382# 0.19fF
C3920 a_2275_12194# col_n[18] 0.17fF
C3921 a_12914_11166# vcm 0.18fF
C3922 a_8990_1126# VDD 0.14fF
C3923 a_2275_1150# col_n[23] 0.17fF
C3924 a_2475_4162# a_29070_4138# 0.68fF
C3925 a_15014_4138# a_16018_4138# 0.86fF
C3926 m2_1732_9982# row_n[8] 0.44fF
C3927 a_26058_11166# col_n[23] 0.34fF
C3928 a_2475_17214# m2_1732_17010# 0.16fF
C3929 a_13006_15182# ctop 4.91fF
C3930 a_5978_6146# row_n[4] 0.43fF
C3931 a_5886_10162# rowon_n[8] 0.14fF
C3932 a_2475_13198# a_7894_13174# 0.41fF
C3933 a_2275_13198# a_5278_13214# 0.15fF
C3934 a_4882_13174# a_4974_13174# 0.45fF
C3935 a_29070_10162# rowoff_n[8] 1.35fF
C3936 a_2275_9182# col[8] 0.17fF
C3937 col[28] rowoff_n[14] 0.16fF
C3938 a_6282_15222# col_n[3] 0.11fF
C3939 a_32994_13174# rowoff_n[11] 0.40fF
C3940 col_n[11] rowoff_n[10] 0.26fF
C3941 a_2275_1150# a_20034_1126# 0.79fF
C3942 a_27974_15182# vcm 0.18fF
C3943 a_24050_5142# VDD 2.27fF
C3944 m2_28840_946# VDD 3.40fF
C3945 a_5978_6146# a_5978_5142# 0.84fF
C3946 a_2475_8178# col[28] 0.22fF
C3947 a_2475_15206# a_22954_15182# 0.41fF
C3948 a_2275_15206# a_20338_15222# 0.15fF
C3949 a_2275_3158# a_35094_3134# 0.14fF
C3950 a_8898_18194# vcm 0.18fF
C3951 a_4974_8154# VDD 4.23fF
C3952 a_30074_8154# a_31078_8154# 0.86fF
C3953 a_26058_13174# rowon_n[11] 0.45fF
C3954 vcm col_n[25] 3.22fF
C3955 a_15014_9158# col_n[12] 0.34fF
C3956 VDD col_n[28] 9.50fF
C3957 col[12] rowoff_n[15] 0.27fF
C3958 a_2275_12194# a_13918_12170# 0.17fF
C3959 a_10998_3134# vcm 0.89fF
C3960 a_2275_11190# col[25] 0.17fF
C3961 a_19942_17190# a_20034_17190# 0.45fF
C3962 a_2966_15182# col_n[0] 0.34fF
C3963 a_3970_13174# row_n[11] 0.43fF
C3964 a_20034_12170# VDD 2.68fF
C3965 a_2475_9182# a_5978_9158# 0.68fF
C3966 a_21038_10162# a_21038_9158# 0.84fF
C3967 a_2275_14202# a_28978_14178# 0.17fF
C3968 a_14010_3134# row_n[1] 0.43fF
C3969 a_26058_7150# vcm 0.89fF
C3970 a_13918_7150# rowon_n[5] 0.14fF
C3971 a_20946_14178# rowoff_n[12] 0.54fF
C3972 a_2275_5166# row_n[3] 26.41fF
C3973 a_2475_11190# a_21038_11166# 0.68fF
C3974 a_10998_11166# a_12002_11166# 0.86fF
C3975 a_16322_1166# vcm 0.25fF
C3976 a_3970_7150# col_n[1] 0.34fF
C3977 a_30378_8194# col_n[27] 0.11fF
C3978 a_2475_15206# col[0] 0.20fF
C3979 a_2475_4162# col[5] 0.22fF
C3980 a_6982_10162# vcm 0.89fF
C3981 a_1957_17214# rowoff_n[15] 0.14fF
C3982 a_29982_4138# a_30074_4138# 0.45fF
C3983 a_2966_9158# m2_1732_8978# 0.86fF
C3984 a_2275_8178# a_12002_8154# 0.71fF
C3985 a_2275_10186# col_n[12] 0.17fF
C3986 a_34090_10162# rowon_n[8] 0.45fF
C3987 a_31382_5182# vcm 0.24fF
C3988 a_22042_14178# vcm 0.89fF
C3989 a_24050_6146# col[21] 0.38fF
C3990 a_18938_4138# VDD 0.29fF
C3991 a_2275_12194# m2_34864_11990# 0.51fF
C3992 a_2475_5166# a_4882_5142# 0.41fF
C3993 a_2275_5166# a_3878_5142# 0.17fF
C3994 a_2275_7174# col[2] 0.17fF
C3995 a_2275_10186# a_27062_10162# 0.71fF
C3996 a_12002_10162# row_n[8] 0.43fF
C3997 a_11910_14178# rowon_n[12] 0.14fF
C3998 a_26058_15182# a_27062_15182# 0.86fF
C3999 a_2475_17214# col[17] 0.22fF
C4000 a_12306_8194# vcm 0.24fF
C4001 col_n[30] rowoff_n[1] 0.12fF
C4002 col_n[31] rowoff_n[2] 0.11fF
C4003 col_n[29] rowoff_n[0] 0.13fF
C4004 a_8898_15182# rowoff_n[13] 0.67fF
C4005 a_2475_6170# col[22] 0.22fF
C4006 a_19334_6186# col_n[16] 0.11fF
C4007 a_21950_4138# rowon_n[2] 0.14fF
C4008 a_25054_3134# ctop 4.91fF
C4009 a_2874_17190# vcm 0.18fF
C4010 a_29374_18234# col_n[26] 0.11fF
C4011 a_18026_1126# m3_17928_1078# 3.21fF
C4012 a_33998_8154# VDD 0.29fF
C4013 a_10906_7150# rowoff_n[5] 0.65fF
C4014 a_2475_7174# a_19942_7150# 0.41fF
C4015 a_2275_7174# a_17326_7190# 0.15fF
C4016 a_10906_7150# a_10998_7150# 0.45fF
C4017 a_2275_12194# col_n[29] 0.17fF
C4018 a_5886_2130# vcm 0.18fF
C4019 a_17022_17190# a_17022_16186# 0.84fF
C4020 a_19942_5142# rowoff_n[3] 0.55fF
C4021 a_27366_12210# vcm 0.24fF
C4022 a_35002_11166# m2_34864_10986# 0.33fF
C4023 a_2275_4162# a_10906_4138# 0.17fF
C4024 a_5978_6146# ctop 4.91fF
C4025 a_13006_4138# col[10] 0.38fF
C4026 a_14922_11166# VDD 0.29fF
C4027 m2_24824_946# col_n[22] 0.45fF
C4028 a_32082_17190# rowon_n[15] 0.45fF
C4029 a_2275_9182# a_32386_9198# 0.15fF
C4030 a_2475_9182# a_35002_9158# 0.41fF
C4031 a_2275_9182# col[19] 0.17fF
C4032 a_23046_16186# col[20] 0.38fF
C4033 m2_1732_6970# sample_n 0.12fF
C4034 a_28978_3134# rowoff_n[1] 0.44fF
C4035 col_n[22] rowoff_n[10] 0.18fF
C4036 a_20946_6146# vcm 0.18fF
C4037 a_2475_1150# a_2874_1126# 0.41fF
C4038 a_1957_1150# a_2275_1150# 0.19fF
C4039 a_8290_15222# vcm 0.24fF
C4040 a_2475_18218# a_13918_18194# 0.41fF
C4041 a_8290_4178# col_n[5] 0.11fF
C4042 a_2275_6170# a_25966_6146# 0.17fF
C4043 a_21038_10162# ctop 4.91fF
C4044 a_9994_17190# row_n[15] 0.43fF
C4045 a_18330_16226# col_n[15] 0.11fF
C4046 a_29982_15182# VDD 0.29fF
C4047 a_25966_11166# a_26058_11166# 0.45fF
C4048 m2_23820_18014# vcm 0.71fF
C4049 a_20034_7150# row_n[5] 0.43fF
C4050 a_2275_15206# a_3970_15182# 0.71fF
C4051 a_19942_11166# rowon_n[9] 0.14fF
C4052 a_34394_10202# vcm 0.24fF
C4053 a_2475_3158# a_18026_3134# 0.68fF
C4054 a_27062_4138# a_27062_3134# 0.84fF
C4055 a_2275_1150# m2_13780_946# 0.51fF
C4056 col_n[2] rowon_n[14] 0.17fF
C4057 col_n[3] row_n[15] 0.37fF
C4058 sample rowon_n[12] 0.10fF
C4059 VDD row_n[12] 4.64fF
C4060 col_n[4] rowon_n[15] 0.17fF
C4061 vcm rowon_n[13] 0.91fF
C4062 col_n[0] row_n[13] 0.37fF
C4063 col_n[1] row_n[14] 0.37fF
C4064 m3_11904_1078# ctop 0.21fF
C4065 col[23] rowoff_n[15] 0.19fF
C4066 a_13006_16186# m2_13204_16434# 0.19fF
C4067 a_10906_18194# VDD 0.50fF
C4068 col_n[6] rowoff_n[11] 0.29fF
C4069 a_12002_14178# col[9] 0.38fF
C4070 a_21038_11166# rowoff_n[9] 1.74fF
C4071 a_2275_17214# a_19030_17190# 0.71fF
C4072 m2_10768_18014# m2_11196_18442# 0.19fF
C4073 a_16930_13174# vcm 0.18fF
C4074 a_13006_3134# VDD 3.40fF
C4075 a_27062_10162# col_n[24] 0.34fF
C4076 a_32082_12170# m2_32280_12418# 0.19fF
C4077 a_2475_5166# a_33086_5142# 0.68fF
C4078 a_17022_5142# a_18026_5142# 0.86fF
C4079 a_2275_8178# col_n[6] 0.17fF
C4080 a_1957_12194# VDD 0.28fF
C4081 a_6982_5142# rowon_n[3] 0.45fF
C4082 a_2275_18218# a_29070_18194# 0.14fF
C4083 m2_13780_946# m2_14784_946# 0.86fF
C4084 a_17022_17190# ctop 4.93fF
C4085 a_30074_9158# rowoff_n[7] 1.30fF
C4086 a_7286_14218# col_n[4] 0.11fF
C4087 a_2966_12170# col[0] 0.38fF
C4088 a_6890_14178# a_6982_14178# 0.45fF
C4089 a_2275_14202# a_9294_14218# 0.15fF
C4090 a_2475_14202# a_11910_14178# 0.41fF
C4091 m2_1732_7974# m2_1732_6970# 0.84fF
C4092 a_2275_14202# rowoff_n[12] 0.81fF
C4093 a_2275_2154# a_24050_2130# 0.71fF
C4094 a_31990_17190# vcm 0.18fF
C4095 a_28066_7150# VDD 1.85fF
C4096 a_7986_7150# a_7986_6146# 0.84fF
C4097 a_3970_14178# m2_4168_14426# 0.19fF
C4098 a_2475_15206# col[11] 0.22fF
C4099 a_18026_14178# row_n[12] 0.43fF
C4100 a_2475_11190# a_2966_11166# 0.65fF
C4101 a_2161_11190# a_2275_11190# 0.17fF
C4102 a_2475_4162# col[16] 0.22fF
C4103 a_34090_2130# vcm 0.89fF
C4104 a_2275_16210# a_24354_16226# 0.15fF
C4105 a_2475_16210# a_26970_16186# 0.41fF
C4106 a_28066_4138# row_n[2] 0.43fF
C4107 a_27974_8154# rowon_n[6] 0.14fF
C4108 a_23046_10162# m2_23244_10410# 0.19fF
C4109 a_2275_10186# col_n[23] 0.17fF
C4110 a_8990_10162# VDD 3.82fF
C4111 a_16018_8154# col_n[13] 0.34fF
C4112 a_32082_9158# a_33086_9158# 0.86fF
C4113 a_2275_13198# a_17934_13174# 0.17fF
C4114 a_15014_5142# vcm 0.89fF
C4115 a_8990_12170# rowoff_n[10] 2.33fF
C4116 a_21950_18194# a_22042_18194# 0.11fF
C4117 a_2275_18218# m2_7756_18014# 0.51fF
C4118 a_2475_1150# a_31990_1126# 0.41fF
C4119 a_2275_1150# a_29374_1166# 0.15fF
C4120 a_16930_1126# a_17022_1126# 0.11fF
C4121 a_2275_7174# col[13] 0.17fF
C4122 a_4974_12170# rowon_n[10] 0.45fF
C4123 m3_30980_18146# VDD 0.11fF
C4124 a_24050_14178# VDD 2.27fF
C4125 a_23046_11166# a_23046_10162# 0.84fF
C4126 a_2475_10186# a_9994_10162# 0.68fF
C4127 a_2475_17214# col[28] 0.22fF
C4128 a_15014_2130# rowon_n[0] 0.45fF
C4129 a_2275_15206# a_32994_15182# 0.17fF
C4130 a_30074_9158# vcm 0.89fF
C4131 a_25054_16186# rowoff_n[14] 1.54fF
C4132 a_14010_8154# m2_14208_8402# 0.19fF
C4133 a_3878_4138# rowon_n[2] 0.14fF
C4134 a_4974_17190# VDD 4.23fF
C4135 a_13006_12170# a_14010_12170# 0.86fF
C4136 a_2475_12194# a_25054_12170# 0.68fF
C4137 a_31382_7190# col_n[28] 0.11fF
C4138 a_4974_6146# col_n[2] 0.34fF
C4139 a_20338_3174# vcm 0.24fF
C4140 a_26058_11166# row_n[9] 0.43fF
C4141 a_25966_15182# rowon_n[13] 0.14fF
C4142 a_33086_4138# m2_33284_4386# 0.19fF
C4143 a_10998_12170# vcm 0.89fF
C4144 a_7894_2130# VDD 0.29fF
C4145 a_2275_9182# col[30] 0.17fF
C4146 a_31990_5142# a_32082_5142# 0.45fF
C4147 m2_34864_1950# rowoff_n[0] 1.01fF
C4148 m3_1864_18146# m3_1864_17142# 0.20fF
C4149 a_2275_9182# a_16018_9158# 0.71fF
C4150 a_2475_18218# m2_33860_18014# 0.62fF
C4151 a_3970_14178# a_3970_13174# 0.84fF
C4152 a_2275_6170# vcm 7.71fF
C4153 a_25054_5142# col[22] 0.38fF
C4154 m2_1732_3958# VDD 5.46fF
C4155 a_4974_6146# m2_5172_6394# 0.19fF
C4156 a_26058_16186# vcm 0.89fF
C4157 a_22954_6146# VDD 0.29fF
C4158 a_2475_6170# a_8898_6146# 0.41fF
C4159 a_2275_6170# a_6282_6186# 0.15fF
C4160 a_2966_10162# ctop 4.82fF
C4161 a_13006_9158# rowon_n[7] 0.45fF
C4162 a_2161_8178# rowoff_n[6] 0.14fF
C4163 a_2275_11190# a_31078_11166# 0.71fF
C4164 a_28978_1126# vcm 0.18fF
C4165 a_1957_7174# row_n[5] 0.29fF
C4166 a_28066_16186# a_29070_16186# 0.86fF
C4167 m2_1732_11990# rowon_n[10] 0.43fF
C4168 a_20338_5182# col_n[17] 0.11fF
C4169 a_16322_10202# vcm 0.24fF
C4170 col_n[8] row_n[12] 0.37fF
C4171 col_n[7] rowon_n[11] 0.17fF
C4172 vcm row_n[8] 1.08fF
C4173 col_n[15] rowon_n[15] 0.17fF
C4174 sample row_n[7] 0.92fF
C4175 col_n[4] row_n[10] 0.37fF
C4176 VDD rowon_n[6] 4.61fF
C4177 col_n[13] rowon_n[14] 0.17fF
C4178 col_n[2] row_n[9] 0.37fF
C4179 col_n[11] rowon_n[13] 0.17fF
C4180 col_n[6] row_n[11] 0.37fF
C4181 col_n[5] rowon_n[10] 0.17fF
C4182 col_n[3] rowon_n[9] 0.17fF
C4183 col_n[9] rowon_n[12] 0.17fF
C4184 col_n[10] row_n[13] 0.37fF
C4185 col_n[12] row_n[14] 0.37fF
C4186 col_n[0] rowon_n[7] 0.17fF
C4187 col_n[14] row_n[15] 0.37fF
C4188 col_n[1] rowon_n[8] 0.17fF
C4189 a_30378_17230# col_n[27] 0.11fF
C4190 a_3970_16186# col_n[1] 0.34fF
C4191 a_13006_17190# rowoff_n[15] 2.13fF
C4192 m2_27836_18014# VDD 2.73fF
C4193 a_2475_13198# col[5] 0.22fF
C4194 a_11910_6146# rowoff_n[4] 0.64fF
C4195 a_29070_5142# ctop 4.91fF
C4196 a_2475_2154# col[10] 0.22fF
C4197 m3_7888_18146# ctop 0.21fF
C4198 col_n[17] rowoff_n[11] 0.21fF
C4199 a_12914_8154# a_13006_8154# 0.45fF
C4200 a_2275_8178# a_21342_8194# 0.15fF
C4201 a_2475_8178# a_23958_8154# 0.41fF
C4202 a_9902_4138# vcm 0.18fF
C4203 a_20946_4138# rowoff_n[2] 0.54fF
C4204 a_2966_11166# rowoff_n[9] 2.62fF
C4205 a_2275_8178# col_n[17] 0.17fF
C4206 a_34090_8154# row_n[6] 0.43fF
C4207 a_31382_14218# vcm 0.24fF
C4208 a_33998_12170# rowon_n[10] 0.14fF
C4209 a_14010_3134# col[11] 0.38fF
C4210 a_2275_5166# a_14922_5142# 0.17fF
C4211 a_9994_8154# ctop 4.91fF
C4212 a_24050_15182# col[21] 0.38fF
C4213 a_18938_13174# VDD 0.29fF
C4214 a_2966_10162# a_2966_9158# 0.84fF
C4215 a_29982_2130# rowoff_n[0] 0.43fF
C4216 a_2275_16210# col[2] 0.17fF
C4217 a_2275_5166# col[7] 0.17fF
C4218 a_24962_8154# vcm 0.18fF
C4219 a_2275_7174# m2_1732_6970# 0.27fF
C4220 a_2475_2154# a_6982_2130# 0.68fF
C4221 a_3970_2130# a_4974_2130# 0.86fF
C4222 a_9294_3174# col_n[6] 0.11fF
C4223 a_12306_17230# vcm 0.24fF
C4224 a_10998_16186# rowon_n[14] 0.45fF
C4225 col_n[1] rowoff_n[12] 0.33fF
C4226 m2_20808_18014# m3_20940_18146# 4.41fF
C4227 a_19334_15222# col_n[16] 0.11fF
C4228 a_2475_15206# col[22] 0.22fF
C4229 a_2275_7174# a_29982_7150# 0.17fF
C4230 a_2475_4162# col[27] 0.22fF
C4231 a_25054_12170# ctop 4.91fF
C4232 a_33998_17190# VDD 0.29fF
C4233 a_27974_12170# a_28066_12170# 0.45fF
C4234 a_21038_6146# rowon_n[4] 0.45fF
C4235 a_2275_16210# a_7986_16186# 0.71fF
C4236 a_5886_11166# vcm 0.18fF
C4237 a_2475_1150# VDD 47.34fF
C4238 a_2475_4162# a_22042_4138# 0.68fF
C4239 a_29070_5142# a_29070_4138# 0.84fF
C4240 a_5978_15182# ctop 4.91fF
C4241 a_13006_13174# col[10] 0.38fF
C4242 a_22042_10162# rowoff_n[8] 1.69fF
C4243 a_32082_15182# row_n[13] 0.43fF
C4244 a_2275_7174# col[24] 0.17fF
C4245 a_25966_13174# rowoff_n[11] 0.48fF
C4246 a_28066_9158# col_n[25] 0.34fF
C4247 a_2275_1150# a_13006_1126# 0.14fF
C4248 a_20946_15182# vcm 0.18fF
C4249 a_17022_5142# VDD 2.99fF
C4250 a_19030_6146# a_20034_6146# 0.86fF
C4251 m2_5748_18014# col_n[3] 0.34fF
C4252 row_n[4] rowoff_n[4] 0.64fF
C4253 a_31078_8154# rowoff_n[6] 1.25fF
C4254 a_8290_13214# col_n[5] 0.11fF
C4255 a_2475_15206# a_15926_15182# 0.41fF
C4256 a_2275_15206# a_13310_15222# 0.15fF
C4257 a_8898_15182# a_8990_15182# 0.45fF
C4258 a_34090_9158# m2_34864_8978# 0.86fF
C4259 a_2275_3158# a_28066_3134# 0.71fF
C4260 a_13918_1126# m2_13780_946# 0.31fF
C4261 a_32082_9158# VDD 1.44fF
C4262 a_9994_8154# a_9994_7150# 0.84fF
C4263 a_2475_18218# vcm 1.32fF
C4264 a_19030_13174# rowon_n[11] 0.45fF
C4265 a_2275_12194# a_6890_12170# 0.17fF
C4266 a_3970_3134# vcm 0.89fF
C4267 a_29070_3134# rowon_n[1] 0.45fF
C4268 a_2475_17214# a_30986_17190# 0.41fF
C4269 a_2275_17214# a_28370_17230# 0.15fF
C4270 a_17022_7150# col_n[14] 0.34fF
C4271 a_13006_12170# VDD 3.40fF
C4272 a_2275_17214# col_n[6] 0.17fF
C4273 a_2275_6170# col_n[11] 0.17fF
C4274 a_2275_14202# a_21950_14178# 0.17fF
C4275 a_6982_3134# row_n[1] 0.43fF
C4276 a_6890_7150# rowon_n[5] 0.14fF
C4277 a_19030_7150# vcm 0.89fF
C4278 a_13918_14178# rowoff_n[12] 0.61fF
C4279 a_2275_2154# a_33390_2170# 0.15fF
C4280 a_18938_2130# a_19030_2130# 0.45fF
C4281 a_2275_3158# col[1] 0.17fF
C4282 a_28066_16186# VDD 1.85fF
C4283 a_25054_12170# a_25054_11166# 0.84fF
C4284 a_2475_11190# a_14010_11166# 0.68fF
C4285 col_n[16] rowon_n[10] 0.17fF
C4286 VDD row_n[1] 4.64fF
C4287 a_9294_1166# vcm 0.25fF
C4288 col_n[14] rowon_n[9] 0.17fF
C4289 col_n[12] rowon_n[8] 0.17fF
C4290 col_n[19] row_n[12] 0.37fF
C4291 col_n[18] rowon_n[11] 0.17fF
C4292 col_n[10] rowon_n[7] 0.17fF
C4293 col_n[1] row_n[3] 0.37fF
C4294 col_n[0] row_n[2] 0.37fF
C4295 col_n[26] rowon_n[15] 0.17fF
C4296 col_n[8] rowon_n[6] 0.17fF
C4297 col_n[3] row_n[4] 0.37fF
C4298 col_n[20] rowon_n[12] 0.17fF
C4299 col_n[21] row_n[13] 0.37fF
C4300 col_n[5] row_n[5] 0.37fF
C4301 col_n[23] row_n[14] 0.37fF
C4302 col_n[7] row_n[6] 0.37fF
C4303 col_n[25] row_n[15] 0.37fF
C4304 col_n[9] row_n[7] 0.37fF
C4305 col_n[2] rowon_n[3] 0.17fF
C4306 col_n[17] row_n[11] 0.37fF
C4307 col_n[11] row_n[8] 0.37fF
C4308 col_n[4] rowon_n[4] 0.17fF
C4309 sample rowon_n[1] 0.10fF
C4310 col_n[22] rowon_n[13] 0.17fF
C4311 col_n[13] row_n[9] 0.37fF
C4312 col_n[6] rowon_n[5] 0.17fF
C4313 vcm rowon_n[2] 0.91fF
C4314 col_n[24] rowon_n[14] 0.17fF
C4315 col_n[15] row_n[10] 0.37fF
C4316 a_2475_13198# col[16] 0.22fF
C4317 a_34090_11166# vcm 0.89fF
C4318 a_2475_2154# col[21] 0.22fF
C4319 col_n[28] rowoff_n[11] 0.14fF
C4320 a_30986_1126# VDD 0.69fF
C4321 a_3878_8154# a_3970_8154# 0.45fF
C4322 a_2275_8178# a_4974_8154# 0.71fF
C4323 a_19030_17190# m2_19228_17438# 0.19fF
C4324 a_32386_6186# col_n[29] 0.11fF
C4325 a_5978_5142# col_n[3] 0.34fF
C4326 a_15014_13174# a_16018_13174# 0.86fF
C4327 a_16018_17190# col_n[13] 0.34fF
C4328 a_2475_13198# a_29070_13174# 0.68fF
C4329 a_27062_10162# rowon_n[8] 0.45fF
C4330 a_2275_8178# col_n[28] 0.17fF
C4331 a_24354_5182# vcm 0.24fF
C4332 a_2275_4162# rowoff_n[2] 0.81fF
C4333 m2_1732_946# a_2475_1150# 0.16fF
C4334 a_15014_14178# vcm 0.89fF
C4335 a_11910_4138# VDD 0.29fF
C4336 a_33998_6146# a_34090_6146# 0.45fF
C4337 a_2275_16210# col[13] 0.17fF
C4338 a_2275_5166# col[18] 0.17fF
C4339 a_2275_10186# a_20034_10162# 0.71fF
C4340 a_4974_10162# row_n[8] 0.43fF
C4341 a_4882_14178# rowon_n[12] 0.14fF
C4342 a_5978_15182# a_5978_14178# 0.84fF
C4343 a_26058_4138# col[23] 0.38fF
C4344 col_n[12] rowoff_n[12] 0.25fF
C4345 a_5278_8194# vcm 0.24fF
C4346 a_14922_4138# rowon_n[2] 0.14fF
C4347 a_18026_3134# ctop 4.91fF
C4348 a_30074_18194# vcm 0.15fF
C4349 a_26970_8154# VDD 0.29fF
C4350 a_2275_7174# a_10298_7190# 0.15fF
C4351 a_2475_7174# a_12914_7150# 0.41fF
C4352 a_9994_15182# m2_10192_15430# 0.19fF
C4353 a_2275_12194# a_35094_12170# 0.14fF
C4354 a_2966_6146# rowon_n[4] 0.45fF
C4355 a_21342_4178# col_n[18] 0.11fF
C4356 a_32994_3134# vcm 0.18fF
C4357 a_30074_17190# a_31078_17190# 0.86fF
C4358 a_31382_16226# col_n[28] 0.11fF
C4359 a_4974_15182# col_n[2] 0.34fF
C4360 a_12914_5142# rowoff_n[3] 0.63fF
C4361 a_20338_12210# vcm 0.24fF
C4362 a_29070_11166# m2_29268_11414# 0.19fF
C4363 a_2874_4138# a_2966_4138# 0.45fF
C4364 a_33086_7150# ctop 4.91fF
C4365 a_7894_11166# VDD 0.29fF
C4366 m2_27836_946# m3_27968_1078# 4.41fF
C4367 a_14922_9158# a_15014_9158# 0.45fF
C4368 a_25054_17190# rowon_n[15] 0.45fF
C4369 a_2275_9182# a_25358_9198# 0.15fF
C4370 a_2475_9182# a_27974_9158# 0.41fF
C4371 m2_1732_4962# vcm 1.11fF
C4372 a_21950_3134# rowoff_n[1] 0.52fF
C4373 a_13918_6146# vcm 0.18fF
C4374 a_15014_2130# col[12] 0.38fF
C4375 rowon_n[0] rowoff_n[0] 20.66fF
C4376 ctop rowoff_n[4] 0.28fF
C4377 a_2275_15206# vcm 7.71fF
C4378 a_2475_18218# a_6890_18194# 0.41fF
C4379 a_25054_14178# col[22] 0.38fF
C4380 a_2275_4162# col_n[5] 0.17fF
C4381 a_2275_6170# a_18938_6146# 0.17fF
C4382 a_14010_10162# ctop 4.91fF
C4383 a_22954_15182# VDD 0.29fF
C4384 m2_9764_18014# vcm 0.71fF
C4385 a_13006_7150# row_n[5] 0.43fF
C4386 m2_34864_12994# m2_35292_13422# 0.19fF
C4387 a_12914_11166# rowon_n[9] 0.14fF
C4388 a_10298_2170# col_n[7] 0.11fF
C4389 a_28978_10162# vcm 0.18fF
C4390 a_20338_14218# col_n[17] 0.11fF
C4391 a_2475_3158# a_10998_3134# 0.68fF
C4392 a_20034_9158# m2_20232_9406# 0.19fF
C4393 a_5978_3134# a_6982_3134# 0.86fF
C4394 m2_8760_946# col_n[6] 0.45fF
C4395 a_25054_2130# m2_24824_946# 0.84fF
C4396 m3_34996_10114# ctop 0.22fF
C4397 a_2275_8178# a_33998_8154# 0.17fF
C4398 a_29070_14178# ctop 4.91fF
C4399 a_2475_11190# col[10] 0.22fF
C4400 a_29982_13174# a_30074_13174# 0.45fF
C4401 a_2275_17214# a_12002_17190# 0.71fF
C4402 a_14010_11166# rowoff_n[9] 2.08fF
C4403 m2_3740_18014# m2_4168_18442# 0.19fF
C4404 a_9902_13174# vcm 0.18fF
C4405 a_5978_3134# VDD 4.13fF
C4406 a_2275_17214# col_n[17] 0.17fF
C4407 a_31078_6146# a_31078_5142# 0.84fF
C4408 a_2475_5166# a_26058_5142# 0.68fF
C4409 a_2275_6170# col_n[22] 0.17fF
C4410 a_2275_18218# a_22042_18194# 0.14fF
C4411 a_2275_18218# col_n[2] 0.17fF
C4412 m2_6752_946# m2_7756_946# 0.86fF
C4413 a_14010_12170# col[11] 0.38fF
C4414 a_9994_17190# ctop 4.93fF
C4415 a_23046_9158# rowoff_n[7] 1.64fF
C4416 a_33086_14178# rowon_n[12] 0.45fF
C4417 a_2275_14202# a_3878_14178# 0.17fF
C4418 a_2475_14202# a_4882_14178# 0.41fF
C4419 a_29070_8154# col_n[26] 0.34fF
C4420 a_30074_15182# rowoff_n[13] 1.30fF
C4421 a_2275_14202# col[7] 0.17fF
C4422 a_2275_2154# a_17022_2130# 0.71fF
C4423 a_2275_3158# col[12] 0.17fF
C4424 a_10998_7150# m2_11196_7398# 0.19fF
C4425 a_24962_17190# vcm 0.18fF
C4426 a_21038_7150# VDD 2.58fF
C4427 a_32082_7150# rowoff_n[5] 1.20fF
C4428 a_21038_7150# a_22042_7150# 0.86fF
C4429 a_9294_12210# col_n[6] 0.11fF
C4430 col_n[9] rowon_n[1] 0.17fF
C4431 col_n[16] row_n[5] 0.37fF
C4432 col_n[7] rowon_n[0] 0.17fF
C4433 col_n[14] row_n[4] 0.37fF
C4434 col_n[12] row_n[3] 0.37fF
C4435 col_n[31] rowon_n[12] 0.17fF
C4436 col_n[10] row_n[2] 0.37fF
C4437 rowon_n[14] row_n[14] 21.02fF
C4438 col_n[8] row_n[1] 0.37fF
C4439 col_n[27] rowon_n[10] 0.17fF
C4440 col_n[6] row_n[0] 0.37fF
C4441 col_n[28] row_n[11] 0.37fF
C4442 col_n[13] rowon_n[3] 0.17fF
C4443 col_n[20] row_n[7] 0.37fF
C4444 col_n[11] rowon_n[2] 0.17fF
C4445 col_n[18] row_n[6] 0.37fF
C4446 col_n[22] row_n[8] 0.37fF
C4447 VDD col[0] 19.69fF
C4448 col_n[15] rowon_n[4] 0.17fF
C4449 col_n[24] row_n[9] 0.37fF
C4450 col_n[17] rowon_n[5] 0.17fF
C4451 col_n[26] row_n[10] 0.37fF
C4452 col_n[19] rowon_n[6] 0.17fF
C4453 col_n[21] rowon_n[7] 0.17fF
C4454 col_n[29] rowon_n[11] 0.17fF
C4455 col_n[30] row_n[12] 0.37fF
C4456 col_n[23] rowon_n[8] 0.17fF
C4457 col_n[25] rowon_n[9] 0.17fF
C4458 a_10998_14178# row_n[12] 0.43fF
C4459 a_2475_13198# col[27] 0.22fF
C4460 a_27062_2130# vcm 0.89fF
C4461 a_2475_16210# a_19942_16186# 0.41fF
C4462 a_2275_16210# a_17326_16226# 0.15fF
C4463 a_10906_16186# a_10998_16186# 0.45fF
C4464 a_30074_3134# m2_30272_3382# 0.19fF
C4465 a_21038_4138# row_n[2] 0.43fF
C4466 a_20946_8154# rowon_n[6] 0.14fF
C4467 a_2275_4162# a_32082_4138# 0.71fF
C4468 a_2475_10186# VDD 41.96fF
C4469 m3_29976_1078# m3_30980_1078# 0.21fF
C4470 a_12002_9158# a_12002_8154# 0.84fF
C4471 a_2275_13198# a_10906_13174# 0.17fF
C4472 a_7986_5142# vcm 0.89fF
C4473 a_2475_12194# rowoff_n[10] 4.75fF
C4474 m2_22240_2378# a_22042_2130# 0.19fF
C4475 a_1957_5166# m2_1732_4962# 0.33fF
C4476 a_2275_16210# col[24] 0.17fF
C4477 a_2275_1150# a_22346_1166# 0.15fF
C4478 a_2475_1150# a_24962_1126# 0.41fF
C4479 a_18026_6146# col_n[15] 0.34fF
C4480 a_2275_5166# col[29] 0.17fF
C4481 m3_2868_18146# VDD 0.10fF
C4482 a_17022_14178# VDD 2.99fF
C4483 a_2475_10186# a_2874_10162# 0.41fF
C4484 a_1957_10186# a_2275_10186# 0.19fF
C4485 a_7986_2130# rowon_n[0] 0.45fF
C4486 col_n[23] rowoff_n[12] 0.17fF
C4487 a_2275_15206# a_25966_15182# 0.17fF
C4488 a_2275_2154# col_n[0] 0.17fF
C4489 a_23046_9158# vcm 0.89fF
C4490 a_18026_16186# rowoff_n[14] 1.89fF
C4491 a_20946_3134# a_21038_3134# 0.45fF
C4492 m2_20808_18014# col[18] 0.37fF
C4493 a_2475_12194# a_18026_12170# 0.68fF
C4494 a_27062_13174# a_27062_12170# 0.84fF
C4495 a_19030_11166# row_n[9] 0.43fF
C4496 a_13310_3174# vcm 0.24fF
C4497 a_18938_15182# rowon_n[13] 0.14fF
C4498 a_3970_12170# vcm 0.89fF
C4499 a_35002_3134# VDD 0.36fF
C4500 a_2475_9182# col[4] 0.22fF
C4501 a_28978_5142# rowon_n[3] 0.14fF
C4502 a_33390_5182# col_n[30] 0.11fF
C4503 a_6982_4138# col_n[4] 0.34fF
C4504 a_7894_18194# m2_7756_18014# 0.34fF
C4505 a_2275_9182# a_8990_9158# 0.71fF
C4506 col_n[7] rowoff_n[13] 0.29fF
C4507 a_17022_16186# col_n[14] 0.34fF
C4508 a_2475_18218# m2_19804_18014# 0.62fF
C4509 a_17022_14178# a_18026_14178# 0.86fF
C4510 a_2475_14202# a_33086_14178# 0.68fF
C4511 a_3878_3134# rowoff_n[1] 0.73fF
C4512 col[10] rowoff_n[9] 0.28fF
C4513 col[9] rowoff_n[8] 0.29fF
C4514 col[8] rowoff_n[7] 0.29fF
C4515 col[7] rowoff_n[6] 0.30fF
C4516 col[6] rowoff_n[5] 0.31fF
C4517 col[5] rowoff_n[4] 0.31fF
C4518 col[1] rowoff_n[0] 0.34fF
C4519 col[2] rowoff_n[1] 0.33fF
C4520 col[3] rowoff_n[2] 0.33fF
C4521 col[4] rowoff_n[3] 0.32fF
C4522 a_2275_15206# col_n[11] 0.17fF
C4523 a_28370_7190# vcm 0.24fF
C4524 a_2275_4162# col_n[16] 0.17fF
C4525 a_19030_16186# vcm 0.89fF
C4526 a_15926_6146# VDD 0.29fF
C4527 a_5978_9158# rowon_n[7] 0.45fF
C4528 a_2275_11190# a_24050_11166# 0.71fF
C4529 a_2275_12194# col[1] 0.17fF
C4530 a_27062_3134# col[24] 0.38fF
C4531 a_2275_1150# col[6] 0.17fF
C4532 a_21950_1126# vcm 0.18fF
C4533 a_7986_16186# a_7986_15182# 0.84fF
C4534 m2_1732_5966# rowoff_n[4] 2.46fF
C4535 a_9294_10202# vcm 0.24fF
C4536 a_5978_17190# rowoff_n[15] 2.47fF
C4537 m2_13780_18014# VDD 4.14fF
C4538 a_4882_6146# rowoff_n[4] 0.72fF
C4539 a_22042_5142# ctop 4.91fF
C4540 a_2475_11190# col[21] 0.22fF
C4541 a_30986_10162# VDD 0.29fF
C4542 a_2275_8178# a_14314_8194# 0.15fF
C4543 a_2475_8178# a_16930_8154# 0.41fF
C4544 a_22346_3174# col_n[19] 0.11fF
C4545 ctop rowoff_n[10] 0.28fF
C4546 a_5978_14178# col_n[3] 0.34fF
C4547 a_32386_15222# col_n[29] 0.11fF
C4548 a_30986_12170# rowoff_n[10] 0.42fF
C4549 a_13918_4138# rowoff_n[2] 0.61fF
C4550 a_2275_17214# col_n[28] 0.17fF
C4551 a_27062_8154# row_n[6] 0.43fF
C4552 a_24354_14218# vcm 0.24fF
C4553 a_26970_12170# rowon_n[10] 0.14fF
C4554 a_2275_18218# col_n[13] 0.17fF
C4555 a_2275_5166# a_7894_5142# 0.17fF
C4556 a_11910_13174# VDD 0.29fF
C4557 a_16930_10162# a_17022_10162# 0.45fF
C4558 a_2475_10186# a_31990_10162# 0.41fF
C4559 a_2275_10186# a_29374_10202# 0.15fF
C4560 a_22954_2130# rowoff_n[0] 0.51fF
C4561 a_2275_14202# col[18] 0.17fF
C4562 a_2275_3158# col[23] 0.17fF
C4563 a_17934_8154# vcm 0.18fF
C4564 a_26058_13174# col[23] 0.38fF
C4565 a_18026_3134# a_18026_2130# 0.84fF
C4566 a_5278_17230# vcm 0.24fF
C4567 col_n[26] rowon_n[4] 0.17fF
C4568 col_n[24] rowon_n[3] 0.17fF
C4569 col_n[31] row_n[7] 0.37fF
C4570 col_n[22] rowon_n[2] 0.17fF
C4571 col_n[29] row_n[6] 0.37fF
C4572 col_n[4] col[4] 0.50fF
C4573 vcm col[8] 6.66fF
C4574 col_n[20] rowon_n[1] 0.17fF
C4575 col_n[27] row_n[5] 0.37fF
C4576 col_n[18] rowon_n[0] 0.17fF
C4577 col_n[25] row_n[4] 0.37fF
C4578 col_n[23] row_n[3] 0.37fF
C4579 col_n[30] rowon_n[6] 0.17fF
C4580 col_n[28] rowon_n[5] 0.17fF
C4581 col_n[17] row_n[0] 0.37fF
C4582 col_n[19] row_n[1] 0.37fF
C4583 col_n[21] row_n[2] 0.37fF
C4584 VDD col[11] 10.71fF
C4585 a_3970_16186# rowon_n[14] 0.45fF
C4586 a_2966_7150# VDD 4.45fF
C4587 a_2275_7174# a_22954_7150# 0.17fF
C4588 a_18026_12170# ctop 4.91fF
C4589 a_26970_17190# VDD 0.29fF
C4590 a_14010_6146# rowon_n[4] 0.45fF
C4591 a_11302_1166# col_n[8] 0.11fF
C4592 a_21342_13214# col_n[18] 0.11fF
C4593 a_2966_4138# row_n[2] 0.41fF
C4594 a_32994_12170# vcm 0.18fF
C4595 a_29070_2130# VDD 1.75fF
C4596 a_2275_8178# rowon_n[6] 1.99fF
C4597 a_7986_4138# a_8990_4138# 0.86fF
C4598 a_2966_10162# m2_3164_10410# 0.19fF
C4599 a_2475_4162# a_15014_4138# 0.68fF
C4600 m3_34996_5094# m3_34996_4090# 0.20fF
C4601 a_3970_17190# m2_3740_18014# 0.84fF
C4602 a_26970_18194# m2_26832_18014# 0.34fF
C4603 a_33086_16186# ctop 4.91fF
C4604 a_31990_14178# a_32082_14178# 0.45fF
C4605 a_15014_10162# rowoff_n[8] 2.03fF
C4606 a_25054_15182# row_n[13] 0.43fF
C4607 a_18938_13174# rowoff_n[11] 0.56fF
C4608 a_2275_1150# a_5978_1126# 0.14fF
C4609 a_13918_15182# vcm 0.18fF
C4610 a_9994_5142# VDD 3.71fF
C4611 a_15014_11166# col[12] 0.38fF
C4612 a_33086_7150# a_33086_6146# 0.84fF
C4613 a_2475_6170# a_30074_6146# 0.68fF
C4614 a_35002_9158# rowon_n[7] 0.14fF
C4615 a_24050_8154# rowoff_n[6] 1.59fF
C4616 a_2275_13198# col_n[5] 0.17fF
C4617 a_2275_2154# col_n[10] 0.17fF
C4618 a_30074_7150# col_n[27] 0.34fF
C4619 a_2475_15206# a_8898_15182# 0.41fF
C4620 a_2275_15206# a_6282_15222# 0.15fF
C4621 a_35002_17190# rowoff_n[15] 0.38fF
C4622 m2_34864_16006# VDD 1.58fF
C4623 a_2275_3158# a_21038_3134# 0.71fF
C4624 a_33086_6146# rowoff_n[4] 1.15fF
C4625 a_10298_11206# col_n[7] 0.11fF
C4626 a_2275_1150# m2_22816_946# 0.51fF
C4627 m3_26964_1078# ctop 0.21fF
C4628 a_25054_9158# VDD 2.16fF
C4629 a_23046_8154# a_24050_8154# 0.86fF
C4630 a_16018_16186# m2_16216_16434# 0.19fF
C4631 a_12002_13174# rowon_n[11] 0.45fF
C4632 a_31078_4138# vcm 0.89fF
C4633 a_22042_3134# rowon_n[1] 0.45fF
C4634 a_2475_17214# a_23958_17190# 0.41fF
C4635 a_2275_17214# a_21342_17230# 0.15fF
C4636 a_12914_17190# a_13006_17190# 0.45fF
C4637 a_2475_9182# col[15] 0.22fF
C4638 col_n[18] rowoff_n[13] 0.21fF
C4639 a_2275_18218# a_31382_18234# 0.15fF
C4640 a_5978_12170# VDD 4.13fF
C4641 a_14010_10162# a_14010_9158# 0.84fF
C4642 a_3970_9158# col[1] 0.38fF
C4643 col[12] rowoff_n[0] 0.27fF
C4644 col[13] rowoff_n[1] 0.26fF
C4645 col[14] rowoff_n[2] 0.25fF
C4646 col[15] rowoff_n[3] 0.25fF
C4647 col[16] rowoff_n[4] 0.24fF
C4648 col[17] rowoff_n[5] 0.23fF
C4649 col[18] rowoff_n[6] 0.23fF
C4650 col[19] rowoff_n[7] 0.22fF
C4651 col[20] rowoff_n[8] 0.21fF
C4652 col[21] rowoff_n[9] 0.21fF
C4653 a_2275_15206# col_n[22] 0.17fF
C4654 a_2275_4162# col_n[27] 0.17fF
C4655 a_2275_14202# a_14922_14178# 0.17fF
C4656 a_12002_7150# vcm 0.89fF
C4657 a_6890_14178# rowoff_n[12] 0.69fF
C4658 a_19030_5142# col_n[16] 0.34fF
C4659 a_33086_12170# row_n[10] 0.43fF
C4660 a_2275_2154# a_26362_2170# 0.15fF
C4661 a_2475_2154# a_28978_2130# 0.41fF
C4662 a_29070_17190# col_n[26] 0.34fF
C4663 a_32994_16186# rowon_n[14] 0.14fF
C4664 a_2275_12194# col[12] 0.17fF
C4665 a_6982_14178# m2_7180_14426# 0.19fF
C4666 a_21038_16186# VDD 2.58fF
C4667 a_2275_1150# col[17] 0.16fF
C4668 a_3970_11166# a_4974_11166# 0.86fF
C4669 a_2475_11190# a_6982_11166# 0.68fF
C4670 a_3878_1126# vcm 0.18fF
C4671 a_2275_16210# a_29982_16186# 0.17fF
C4672 a_3970_2130# m2_4168_2378# 0.19fF
C4673 a_27062_11166# vcm 0.89fF
C4674 col_n[2] rowoff_n[14] 0.32fF
C4675 a_23958_1126# VDD 0.77fF
C4676 a_22954_4138# a_23046_4138# 0.45fF
C4677 a_26058_10162# m2_26256_10410# 0.19fF
C4678 a_23046_17190# m2_22816_18014# 0.84fF
C4679 col[5] rowoff_n[10] 0.31fF
C4680 a_20034_10162# rowon_n[8] 0.45fF
C4681 a_29070_14178# a_29070_13174# 0.84fF
C4682 a_2475_13198# a_22042_13174# 0.68fF
C4683 a_17326_5182# vcm 0.24fF
C4684 a_2275_18218# col_n[24] 0.17fF
C4685 m2_16792_946# vcm 0.71fF
C4686 a_2275_1150# a_33390_1166# 0.15fF
C4687 a_7986_14178# vcm 0.89fF
C4688 a_4882_4138# VDD 0.29fF
C4689 a_7986_3134# col_n[5] 0.34fF
C4690 a_18026_15182# col_n[15] 0.34fF
C4691 a_2275_14202# col[29] 0.17fF
C4692 a_2275_10186# a_13006_10162# 0.71fF
C4693 a_19030_15182# a_20034_15182# 0.86fF
C4694 VDD col[22] 7.99fF
C4695 col_n[9] col[10] 6.22fF
C4696 col_n[28] row_n[0] 0.37fF
C4697 vcm col[19] 6.66fF
C4698 a_32386_9198# vcm 0.24fF
C4699 col_n[30] row_n[1] 0.37fF
C4700 col_n[29] rowon_n[0] 0.17fF
C4701 col_n[31] rowon_n[1] 0.17fF
C4702 a_7894_4138# rowon_n[2] 0.14fF
C4703 a_17022_8154# m2_17220_8402# 0.19fF
C4704 a_2275_11190# col_n[0] 0.17fF
C4705 a_23046_18194# vcm 0.15fF
C4706 a_10998_3134# ctop 4.91fF
C4707 a_19942_8154# VDD 0.29fF
C4708 a_2275_7174# a_3270_7190# 0.15fF
C4709 a_2475_7174# a_5886_7150# 0.41fF
C4710 a_28066_2130# col[25] 0.38fF
C4711 a_2275_12194# a_28066_12170# 0.71fF
C4712 a_25966_3134# vcm 0.18fF
C4713 a_9994_17190# a_9994_16186# 0.84fF
C4714 a_5886_5142# rowoff_n[3] 0.70fF
C4715 a_13310_12210# vcm 0.24fF
C4716 a_26058_7150# ctop 4.91fF
C4717 a_35002_12170# VDD 0.36fF
C4718 m3_25960_18146# m3_26964_18146# 0.21fF
C4719 a_23350_2170# col_n[20] 0.11fF
C4720 a_2475_9182# a_20946_9158# 0.41fF
C4721 a_2275_9182# a_18330_9198# 0.15fF
C4722 a_18026_17190# rowon_n[15] 0.45fF
C4723 a_2475_7174# col[9] 0.22fF
C4724 a_6982_13174# col_n[4] 0.34fF
C4725 a_33390_14218# col_n[30] 0.11fF
C4726 m2_1732_2954# rowon_n[1] 0.43fF
C4727 a_14922_3134# rowoff_n[1] 0.60fF
C4728 a_28066_7150# rowon_n[5] 0.45fF
C4729 a_6890_6146# vcm 0.18fF
C4730 a_2275_18218# a_2966_18194# 0.14fF
C4731 a_29070_2130# a_30074_2130# 0.86fF
C4732 a_7986_6146# m2_8184_6394# 0.19fF
C4733 a_28370_16226# vcm 0.24fF
C4734 a_2275_13198# col_n[16] 0.17fF
C4735 a_2275_6170# a_11910_6146# 0.17fF
C4736 a_2275_2154# col_n[21] 0.17fF
C4737 a_6982_10162# ctop 4.91fF
C4738 a_15926_15182# VDD 0.29fF
C4739 a_2275_11190# a_33390_11206# 0.15fF
C4740 a_18938_11166# a_19030_11166# 0.45fF
C4741 a_5978_7150# row_n[5] 0.43fF
C4742 a_27062_12170# col[24] 0.38fF
C4743 a_5886_11166# rowon_n[9] 0.14fF
C4744 a_21950_10162# vcm 0.18fF
C4745 a_2275_10186# col[6] 0.17fF
C4746 a_20034_4138# a_20034_3134# 0.84fF
C4747 a_2475_3158# a_3970_3134# 0.68fF
C4748 a_2275_3158# a_2966_3134# 0.67fF
C4749 m3_22948_18146# ctop 0.21fF
C4750 a_2475_16210# m2_1732_16006# 0.16fF
C4751 a_2275_8178# a_26970_8154# 0.17fF
C4752 a_22042_14178# ctop 4.91fF
C4753 a_2475_9182# col[26] 0.22fF
C4754 a_22346_12210# col_n[19] 0.11fF
C4755 a_6982_11166# rowoff_n[9] 2.42fF
C4756 a_2275_17214# a_4974_17190# 0.71fF
C4757 a_3878_17190# a_3970_17190# 0.45fF
C4758 col_n[29] rowoff_n[13] 0.13fF
C4759 a_33086_4138# VDD 1.34fF
C4760 a_9994_5142# a_10998_5142# 0.86fF
C4761 a_2475_5166# a_19030_5142# 0.68fF
C4762 col[23] rowoff_n[0] 0.19fF
C4763 col[24] rowoff_n[1] 0.19fF
C4764 col[25] rowoff_n[2] 0.18fF
C4765 col[26] rowoff_n[3] 0.17fF
C4766 col[27] rowoff_n[4] 0.17fF
C4767 col[28] rowoff_n[5] 0.16fF
C4768 col[29] rowoff_n[6] 0.15fF
C4769 col[30] rowoff_n[7] 0.15fF
C4770 col[31] rowoff_n[8] 0.14fF
C4771 sample_n rowoff_n[9] 0.55fF
C4772 a_2275_18218# a_15014_18194# 0.14fF
C4773 a_16018_9158# rowoff_n[7] 1.98fF
C4774 a_26058_14178# rowon_n[12] 0.45fF
C4775 a_33998_15182# a_34090_15182# 0.45fF
C4776 a_23046_15182# rowoff_n[13] 1.64fF
C4777 a_2275_12194# col[23] 0.17fF
C4778 a_2275_2154# a_9994_2130# 0.71fF
C4779 a_16018_10162# col[13] 0.38fF
C4780 a_17934_17190# vcm 0.18fF
C4781 m2_25828_18014# m3_25960_18146# 4.42fF
C4782 a_2275_1150# col[28] 0.17fF
C4783 a_14010_7150# VDD 3.30fF
C4784 a_25054_7150# rowoff_n[5] 1.54fF
C4785 a_2475_7174# a_34090_7150# 0.68fF
C4786 a_2966_16186# VDD 4.45fF
C4787 a_3970_14178# row_n[12] 0.43fF
C4788 a_31078_6146# col_n[28] 0.34fF
C4789 a_20034_2130# vcm 0.89fF
C4790 col_n[13] rowoff_n[14] 0.24fF
C4791 a_2475_16210# a_12914_16186# 0.41fF
C4792 a_2275_16210# a_10298_16226# 0.15fF
C4793 a_34090_5142# rowoff_n[3] 1.10fF
C4794 a_14010_4138# row_n[2] 0.43fF
C4795 a_11302_10202# col_n[8] 0.11fF
C4796 col[16] rowoff_n[10] 0.24fF
C4797 a_13918_8154# rowon_n[6] 0.14fF
C4798 a_2275_4162# a_25054_4138# 0.71fF
C4799 a_29070_11166# VDD 1.75fF
C4800 m3_15920_1078# m3_16924_1078# 0.21fF
C4801 a_25054_9158# a_26058_9158# 0.86fF
C4802 a_2275_6170# row_n[4] 26.41fF
C4803 a_2874_13174# a_2966_13174# 0.45fF
C4804 a_35094_6146# vcm 0.15fF
C4805 a_14922_18194# a_15014_18194# 0.11fF
C4806 a_2275_1150# a_15318_1166# 0.15fF
C4807 a_9902_1126# a_9994_1126# 0.11fF
C4808 a_2475_1150# a_17934_1126# 0.44fF
C4809 a_2475_5166# col[3] 0.22fF
C4810 a_4974_8154# col[2] 0.38fF
C4811 a_9994_14178# VDD 3.71fF
C4812 a_16018_11166# a_16018_10162# 0.84fF
C4813 col_n[15] col[15] 0.43fF
C4814 rowon_n[13] ctop 0.37fF
C4815 sample sample_n 12.16fF
C4816 VDD rowoff_n[15] 87.23fF
C4817 col_n[31] analog_in 0.22fF
C4818 vcm col[30] 6.66fF
C4819 m2_34864_17010# vcm 0.72fF
C4820 a_2275_15206# a_18938_15182# 0.17fF
C4821 a_20034_4138# col_n[17] 0.34fF
C4822 a_2275_11190# col_n[10] 0.17fF
C4823 a_34090_11166# rowon_n[9] 0.45fF
C4824 a_16018_9158# vcm 0.89fF
C4825 col[0] rowoff_n[11] 0.34fF
C4826 a_30074_16186# col_n[27] 0.34fF
C4827 a_10998_16186# rowoff_n[14] 2.23fF
C4828 a_2966_8154# m2_1732_7974# 0.86fF
C4829 a_2275_3158# a_30378_3174# 0.15fF
C4830 a_2475_3158# a_32994_3134# 0.41fF
C4831 a_35398_9198# VDD 0.12fF
C4832 a_2275_8178# col[0] 0.16fF
C4833 a_2475_12194# a_10998_12170# 0.68fF
C4834 a_5978_12170# a_6982_12170# 0.86fF
C4835 a_12002_11166# row_n[9] 0.43fF
C4836 a_6282_3174# vcm 0.24fF
C4837 a_2275_17214# a_33998_17190# 0.17fF
C4838 a_11910_15182# rowon_n[13] 0.14fF
C4839 a_31078_13174# vcm 0.89fF
C4840 a_27974_3134# VDD 0.29fF
C4841 a_24962_5142# a_25054_5142# 0.45fF
C4842 a_2275_11190# m2_34864_10986# 0.51fF
C4843 a_2475_7174# col[20] 0.22fF
C4844 a_21950_5142# rowon_n[3] 0.14fF
C4845 m2_29844_946# m2_30848_946# 0.86fF
C4846 m2_34864_1950# rowon_n[0] 0.42fF
C4847 a_2475_9182# a_2275_9182# 2.96fF
C4848 a_1957_9182# a_2161_9182# 0.11fF
C4849 a_2475_18218# m2_5748_18014# 0.62fF
C4850 a_31078_15182# a_31078_14178# 0.84fF
C4851 a_2475_14202# a_26058_14178# 0.68fF
C4852 a_21342_7190# vcm 0.24fF
C4853 a_2275_13198# col_n[27] 0.17fF
C4854 a_8990_2130# col_n[6] 0.34fF
C4855 a_12002_16186# vcm 0.89fF
C4856 a_34090_2130# ctop 4.90fF
C4857 a_8898_6146# VDD 0.29fF
C4858 a_19030_14178# col_n[16] 0.34fF
C4859 a_2275_11190# a_17022_11166# 0.71fF
C4860 m2_34864_13998# rowoff_n[12] 1.01fF
C4861 a_2275_10186# col[17] 0.17fF
C4862 a_14922_1126# vcm 0.18fF
C4863 a_21038_16186# a_22042_16186# 0.86fF
C4864 m2_1732_7974# sample 0.31fF
C4865 a_3878_10162# vcm 0.18fF
C4866 m2_33860_946# col[31] 0.33fF
C4867 a_35494_1488# VDD 0.15fF
C4868 a_35002_10162# m2_34864_9982# 0.33fF
C4869 a_15014_5142# ctop 4.91fF
C4870 a_7986_2130# m2_7756_946# 0.84fF
C4871 a_23958_10162# VDD 0.29fF
C4872 a_5886_8154# a_5978_8154# 0.45fF
C4873 a_22042_17190# m2_22240_17438# 0.19fF
C4874 a_2475_8178# a_9902_8154# 0.41fF
C4875 a_2275_8178# a_7286_8194# 0.15fF
C4876 a_2275_13198# a_32082_13174# 0.71fF
C4877 a_29982_5142# vcm 0.18fF
C4878 a_6890_4138# rowoff_n[2] 0.69fF
C4879 a_23958_12170# rowoff_n[10] 0.50fF
C4880 a_20034_8154# row_n[6] 0.43fF
C4881 a_17326_14218# vcm 0.24fF
C4882 a_19942_12170# rowon_n[10] 0.14fF
C4883 a_24354_1166# col_n[21] 0.11fF
C4884 a_30074_9158# ctop 4.91fF
C4885 a_4882_13174# VDD 0.29fF
C4886 a_7986_12170# col_n[5] 0.34fF
C4887 a_2475_10186# a_24962_10162# 0.41fF
C4888 a_2275_10186# a_22346_10202# 0.15fF
C4889 a_15926_2130# rowoff_n[0] 0.59fF
C4890 a_29982_2130# rowon_n[0] 0.14fF
C4891 a_10906_8154# vcm 0.18fF
C4892 a_31078_3134# a_32082_3134# 0.86fF
C4893 a_32386_18234# vcm 0.25fF
C4894 a_13006_15182# m2_13204_15430# 0.19fF
C4895 a_2275_7174# a_15926_7150# 0.17fF
C4896 a_10998_12170# ctop 4.91fF
C4897 a_2275_9182# col_n[4] 0.17fF
C4898 a_19942_17190# VDD 0.29fF
C4899 col_n[24] rowoff_n[14] 0.16fF
C4900 a_20946_12170# a_21038_12170# 0.45fF
C4901 a_6982_6146# rowon_n[4] 0.45fF
C4902 a_1957_2154# vcm 0.16fF
C4903 a_28066_11166# col[25] 0.38fF
C4904 col[27] rowoff_n[10] 0.17fF
C4905 m2_1732_16006# m2_2160_16434# 0.19fF
C4906 a_25966_12170# vcm 0.18fF
C4907 a_22042_2130# VDD 2.47fF
C4908 a_22042_5142# a_22042_4138# 0.84fF
C4909 a_2475_4162# a_7986_4138# 0.68fF
C4910 a_32082_11166# m2_32280_11414# 0.19fF
C4911 a_2275_6170# ctop 0.14fF
C4912 m3_34996_12122# m3_34996_11118# 0.20fF
C4913 m2_32856_946# m3_32988_1078# 4.41fF
C4914 a_2275_9182# a_30986_9158# 0.17fF
C4915 a_26058_16186# ctop 4.91fF
C4916 a_23350_11206# col_n[20] 0.11fF
C4917 a_7986_10162# rowoff_n[8] 2.38fF
C4918 a_2475_16210# col[9] 0.22fF
C4919 a_18026_15182# row_n[13] 0.43fF
C4920 a_2475_5166# col[14] 0.22fF
C4921 a_11910_13174# rowoff_n[11] 0.64fF
C4922 a_6890_15182# vcm 0.18fF
C4923 a_2874_5142# VDD 0.29fF
C4924 a_28066_5142# row_n[3] 0.43fF
C4925 a_3970_13174# m2_4168_13422# 0.19fF
C4926 a_12002_6146# a_13006_6146# 0.86fF
C4927 a_2475_6170# a_23046_6146# 0.68fF
C4928 a_27974_9158# rowon_n[7] 0.14fF
C4929 col_n[20] col[21] 6.22fF
C4930 row_n[8] ctop 0.28fF
C4931 col_n[8] rowoff_n[15] 0.28fF
C4932 rowon_n[3] row_n[3] 21.02fF
C4933 a_17022_8154# rowoff_n[6] 1.94fF
C4934 a_2275_11190# col_n[21] 0.17fF
C4935 col[11] rowoff_n[11] 0.27fF
C4936 a_17022_9158# col[14] 0.38fF
C4937 a_27974_17190# rowoff_n[15] 0.46fF
C4938 a_2275_3158# a_14010_3134# 0.71fF
C4939 a_26058_6146# rowoff_n[4] 1.50fF
C4940 a_23046_9158# m2_23244_9406# 0.19fF
C4941 a_2475_1150# m2_8760_946# 0.62fF
C4942 a_3970_1126# m2_4744_946# 0.86fF
C4943 a_18026_9158# VDD 2.89fF
C4944 a_2275_8178# col[11] 0.17fF
C4945 a_4974_13174# rowon_n[11] 0.45fF
C4946 a_32082_5142# col_n[29] 0.34fF
C4947 a_24050_4138# vcm 0.89fF
C4948 a_15014_3134# rowon_n[1] 0.45fF
C4949 a_2475_17214# a_16930_17190# 0.41fF
C4950 a_2275_17214# a_14314_17230# 0.15fF
C4951 a_12306_9198# col_n[9] 0.11fF
C4952 a_2475_7174# col[31] 0.22fF
C4953 a_2275_5166# a_29070_5142# 0.71fF
C4954 a_3878_5142# rowon_n[3] 0.14fF
C4955 a_33086_13174# VDD 1.34fF
C4956 a_2275_18218# a_24354_18234# 0.15fF
C4957 m2_10768_946# m2_11196_1374# 0.19fF
C4958 a_27062_10162# a_28066_10162# 0.86fF
C4959 a_2275_14202# a_7894_14178# 0.17fF
C4960 a_4974_7150# vcm 0.89fF
C4961 a_26058_12170# row_n[10] 0.43fF
C4962 a_11910_2130# a_12002_2130# 0.45fF
C4963 a_2275_2154# a_19334_2170# 0.15fF
C4964 a_2475_2154# a_21950_2130# 0.41fF
C4965 a_14010_7150# m2_14208_7398# 0.19fF
C4966 a_25966_16186# rowon_n[14] 0.14fF
C4967 a_5978_7150# col[3] 0.38fF
C4968 a_2275_10186# col[28] 0.17fF
C4969 a_14010_16186# VDD 3.30fF
C4970 m2_1732_15002# rowoff_n[13] 2.46fF
C4971 a_18026_12170# a_18026_11166# 0.84fF
C4972 a_21038_3134# col_n[18] 0.34fF
C4973 a_29374_2170# vcm 0.24fF
C4974 a_2275_16210# a_22954_16186# 0.17fF
C4975 a_31078_15182# col_n[28] 0.34fF
C4976 a_33086_3134# m2_33284_3382# 0.19fF
C4977 a_20034_11166# vcm 0.89fF
C4978 a_16930_1126# VDD 0.85fF
C4979 a_2275_4162# a_35398_4178# 0.15fF
C4980 a_7986_13174# a_8990_13174# 0.86fF
C4981 a_2475_13198# a_15014_13174# 0.68fF
C4982 a_13006_10162# rowon_n[8] 0.45fF
C4983 a_10298_5182# vcm 0.24fF
C4984 m2_25252_2378# a_25054_2130# 0.19fF
C4985 a_2275_1150# a_27974_1126# 0.17fF
C4986 a_1957_8178# row_n[6] 0.29fF
C4987 a_4974_5142# m2_5172_5390# 0.19fF
C4988 a_35094_15182# vcm 0.15fF
C4989 a_31990_5142# VDD 0.29fF
C4990 a_26970_6146# a_27062_6146# 0.45fF
C4991 a_2475_14202# col[3] 0.22fF
C4992 a_2275_10186# a_5978_10162# 0.71fF
C4993 a_2475_3158# col[8] 0.22fF
C4994 a_4974_17190# col[2] 0.38fF
C4995 a_2475_15206# a_30074_15182# 0.68fF
C4996 a_33086_16186# a_33086_15182# 0.84fF
C4997 a_25358_9198# vcm 0.24fF
C4998 a_20034_13174# col_n[17] 0.34fF
C4999 a_16018_18194# vcm 0.15fF
C5000 a_3970_3134# ctop 4.93fF
C5001 a_2275_9182# col_n[15] 0.17fF
C5002 a_12914_8154# VDD 0.29fF
C5003 a_34090_9158# row_n[7] 0.43fF
C5004 row_n[14] rowoff_n[14] 0.64fF
C5005 a_33998_13174# rowon_n[11] 0.14fF
C5006 a_35398_18234# VDD 0.14fF
C5007 a_2275_12194# a_21038_12170# 0.71fF
C5008 a_18938_3134# vcm 0.18fF
C5009 a_23046_17190# a_24050_17190# 0.86fF
C5010 a_2275_17214# col[0] 0.16fF
C5011 a_2275_6170# col[5] 0.17fF
C5012 a_6282_12210# vcm 0.24fF
C5013 a_34394_2170# col_n[31] 0.11fF
C5014 a_19030_7150# ctop 4.91fF
C5015 a_27974_12170# VDD 0.29fF
C5016 m3_11904_18146# m3_12908_18146# 0.21fF
C5017 a_2475_9182# a_13918_9158# 0.41fF
C5018 a_2275_9182# a_11302_9198# 0.15fF
C5019 a_10998_17190# rowon_n[15] 0.45fF
C5020 a_7894_9158# a_7986_9158# 0.45fF
C5021 a_2475_16210# col[20] 0.22fF
C5022 a_2475_5166# col[25] 0.22fF
C5023 a_7894_3134# rowoff_n[1] 0.68fF
C5024 a_21038_7150# rowon_n[5] 0.45fF
C5025 a_33998_7150# vcm 0.18fF
C5026 a_28066_14178# rowoff_n[12] 1.40fF
C5027 a_2275_6170# m2_1732_5966# 0.27fF
C5028 col_n[19] rowoff_n[15] 0.20fF
C5029 col_n[26] col[26] 0.55fF
C5030 rowon_n[2] ctop 0.37fF
C5031 a_21342_16226# vcm 0.24fF
C5032 a_8990_11166# col_n[6] 0.34fF
C5033 a_2966_6146# a_3970_6146# 0.86fF
C5034 a_2275_6170# a_4882_6146# 0.17fF
C5035 a_34090_11166# ctop 4.80fF
C5036 a_8898_15182# VDD 0.29fF
C5037 col[22] rowoff_n[11] 0.20fF
C5038 a_2475_11190# a_28978_11166# 0.41fF
C5039 a_2275_11190# a_26362_11206# 0.15fF
C5040 a_14922_10162# vcm 0.18fF
C5041 a_32082_16186# row_n[14] 0.43fF
C5042 a_2275_8178# col[22] 0.17fF
C5043 a_33086_4138# a_34090_4138# 0.86fF
C5044 a_2275_8178# a_19942_8154# 0.17fF
C5045 a_15014_14178# ctop 4.91fF
C5046 a_29070_10162# col[26] 0.38fF
C5047 a_22954_13174# a_23046_13174# 0.45fF
C5048 m2_14784_18014# col[12] 0.39fF
C5049 a_29982_14178# vcm 0.18fF
C5050 a_26058_4138# VDD 2.06fF
C5051 a_2475_5166# a_12002_5142# 0.68fF
C5052 a_24050_6146# a_24050_5142# 0.84fF
C5053 col[6] rowoff_n[12] 0.31fF
C5054 a_2275_18218# a_7986_18194# 0.14fF
C5055 a_2275_10186# a_35002_10162# 0.17fF
C5056 a_24354_10202# col_n[21] 0.11fF
C5057 a_8990_9158# rowoff_n[7] 2.33fF
C5058 a_19030_14178# rowon_n[12] 0.45fF
C5059 a_16018_15182# rowoff_n[13] 1.98fF
C5060 a_2275_2154# a_2874_2130# 0.17fF
C5061 a_2475_2154# a_3878_2130# 0.41fF
C5062 a_34090_8154# m2_34864_7974# 0.86fF
C5063 a_29070_4138# rowon_n[2] 0.45fF
C5064 a_10906_17190# vcm 0.18fF
C5065 a_2475_1150# col[2] 0.21fF
C5066 a_6982_7150# VDD 4.02fF
C5067 a_18026_7150# rowoff_n[5] 1.89fF
C5068 a_2475_7174# a_27062_7150# 0.68fF
C5069 a_14010_7150# a_15014_7150# 0.86fF
C5070 a_13006_2130# vcm 0.89fF
C5071 a_2475_16210# a_5886_16186# 0.41fF
C5072 a_2275_16210# a_3270_16226# 0.15fF
C5073 a_2275_7174# col_n[9] 0.17fF
C5074 a_18026_8154# col[15] 0.38fF
C5075 a_1957_11190# vcm 0.16fF
C5076 a_27062_5142# rowoff_n[3] 1.45fF
C5077 a_6982_4138# row_n[2] 0.43fF
C5078 a_6890_8154# rowon_n[6] 0.14fF
C5079 a_2275_4162# a_18026_4138# 0.71fF
C5080 a_22042_11166# VDD 2.47fF
C5081 a_33086_4138# col_n[30] 0.34fF
C5082 m3_1864_1078# m3_2868_1078# 0.21fF
C5083 a_4974_9158# a_4974_8154# 0.84fF
C5084 m2_30848_18014# col_n[28] 0.32fF
C5085 a_2275_15206# ctop 0.14fF
C5086 a_13310_8194# col_n[10] 0.11fF
C5087 a_28066_6146# vcm 0.89fF
C5088 a_2275_1150# a_8290_1166# 0.15fF
C5089 a_2475_1150# a_10906_1126# 0.41fF
C5090 a_2475_14202# col[14] 0.22fF
C5091 a_2475_3158# col[19] 0.22fF
C5092 a_2275_6170# a_33086_6146# 0.71fF
C5093 m2_6752_946# VDD 6.70fF
C5094 a_2874_14178# VDD 0.29fF
C5095 a_2475_18218# col[5] 0.22fF
C5096 a_29070_11166# a_30074_11166# 0.86fF
C5097 a_2275_15206# a_11910_15182# 0.17fF
C5098 a_27062_11166# rowon_n[9] 0.45fF
C5099 a_8990_9158# vcm 0.89fF
C5100 a_2275_9182# col_n[26] 0.17fF
C5101 a_3970_16186# rowoff_n[14] 2.57fF
C5102 a_6982_6146# col[4] 0.38fF
C5103 a_13918_3134# a_14010_3134# 0.45fF
C5104 a_2475_3158# a_25966_3134# 0.41fF
C5105 a_2275_3158# a_23350_3174# 0.15fF
C5106 a_2475_1150# m2_31852_946# 0.62fF
C5107 a_19030_16186# m2_19228_16434# 0.19fF
C5108 a_22042_2130# col_n[19] 0.34fF
C5109 a_2275_17214# col[11] 0.17fF
C5110 a_2275_12194# a_2966_12170# 0.67fF
C5111 a_2475_12194# a_3970_12170# 0.68fF
C5112 a_20034_13174# a_20034_12170# 0.84fF
C5113 a_32082_14178# col_n[29] 0.34fF
C5114 a_2275_6170# col[16] 0.17fF
C5115 a_4974_11166# row_n[9] 0.43fF
C5116 a_33390_4178# vcm 0.24fF
C5117 a_28978_11166# rowoff_n[9] 0.44fF
C5118 a_2275_17214# a_26970_17190# 0.17fF
C5119 a_4882_15182# rowon_n[13] 0.14fF
C5120 a_24050_13174# vcm 0.89fF
C5121 a_20946_3134# VDD 0.29fF
C5122 a_12306_18234# col_n[9] 0.11fF
C5123 a_2475_16210# col[31] 0.22fF
C5124 a_14922_5142# rowon_n[3] 0.14fF
C5125 m2_22816_946# m2_23820_946# 0.86fF
C5126 a_2475_14202# a_19030_14178# 0.68fF
C5127 a_9994_14178# a_10998_14178# 0.86fF
C5128 sw analog_in 0.80fF
C5129 col_n[30] rowoff_n[15] 0.12fF
C5130 a_2966_7150# rowon_n[5] 0.45fF
C5131 a_14314_7190# vcm 0.24fF
C5132 m2_34864_17010# row_n[15] 0.38fF
C5133 a_2275_2154# a_31990_2130# 0.17fF
C5134 a_4974_16186# vcm 0.89fF
C5135 a_27062_2130# ctop 4.93fF
C5136 a_9994_14178# m2_10192_14426# 0.19fF
C5137 a_28978_7150# a_29070_7150# 0.45fF
C5138 a_5978_16186# col[3] 0.38fF
C5139 a_2275_11190# a_9994_11166# 0.71fF
C5140 a_7894_1126# vcm 0.18fF
C5141 a_2475_16210# a_34090_16186# 0.68fF
C5142 a_21038_12170# col_n[18] 0.34fF
C5143 a_6982_2130# m2_7180_2378# 0.19fF
C5144 a_29374_11206# vcm 0.24fF
C5145 a_27462_1488# VDD 0.13fF
C5146 a_29070_10162# m2_29268_10410# 0.19fF
C5147 a_7986_5142# ctop 4.91fF
C5148 a_16930_10162# VDD 0.29fF
C5149 a_2275_5166# col_n[3] 0.17fF
C5150 m2_1732_2954# sample_n 0.12fF
C5151 a_2275_13198# a_25054_13174# 0.71fF
C5152 a_22954_5142# vcm 0.18fF
C5153 a_16930_12170# rowoff_n[10] 0.58fF
C5154 m2_25828_946# vcm 0.71fF
C5155 a_2275_18218# m2_22816_18014# 0.51fF
C5156 col[17] rowoff_n[12] 0.23fF
C5157 a_13006_8154# row_n[6] 0.43fF
C5158 a_10298_14218# vcm 0.24fF
C5159 a_12914_12170# rowon_n[10] 0.14fF
C5160 a_23046_9158# ctop 4.91fF
C5161 a_31990_14178# VDD 0.29fF
C5162 a_2475_10186# a_17934_10162# 0.41fF
C5163 a_2275_10186# a_15318_10202# 0.15fF
C5164 a_9902_10162# a_9994_10162# 0.45fF
C5165 a_8898_2130# rowoff_n[0] 0.67fF
C5166 a_22954_2130# rowon_n[0] 0.14fF
C5167 a_2475_12194# col[8] 0.22fF
C5168 a_2475_1150# col[13] 0.22fF
C5169 a_32994_16186# rowoff_n[14] 0.40fF
C5170 a_10998_3134# a_10998_2130# 0.84fF
C5171 a_20034_8154# m2_20232_8402# 0.19fF
C5172 a_9994_10162# col_n[7] 0.34fF
C5173 a_25358_18234# vcm 0.25fF
C5174 a_2275_7174# a_8898_7150# 0.17fF
C5175 a_3970_12170# ctop 4.91fF
C5176 a_12914_17190# VDD 0.29fF
C5177 a_2275_7174# col_n[20] 0.17fF
C5178 a_2475_12194# a_32994_12170# 0.41fF
C5179 a_2275_12194# a_30378_12210# 0.15fF
C5180 col[1] rowoff_n[13] 0.34fF
C5181 a_33086_15182# rowon_n[13] 0.45fF
C5182 a_18938_12170# vcm 0.18fF
C5183 a_15014_2130# VDD 3.20fF
C5184 a_2275_15206# col[5] 0.17fF
C5185 a_2275_4162# col[10] 0.17fF
C5186 a_34394_11206# col_n[31] 0.11fF
C5187 a_2275_9182# a_23958_9158# 0.17fF
C5188 a_19030_16186# ctop 4.91fF
C5189 a_30074_9158# col[27] 0.38fF
C5190 a_24962_14178# a_25054_14178# 0.45fF
C5191 a_10998_15182# row_n[13] 0.43fF
C5192 m2_1732_5966# m2_1732_4962# 0.84fF
C5193 a_2475_14202# col[25] 0.22fF
C5194 a_4882_13174# rowoff_n[11] 0.72fF
C5195 a_2475_3158# col[30] 0.22fF
C5196 a_10998_6146# m2_11196_6394# 0.19fF
C5197 a_33998_16186# vcm 0.18fF
C5198 a_30074_6146# VDD 1.65fF
C5199 a_2475_18218# col[16] 0.22fF
C5200 a_21038_5142# row_n[3] 0.43fF
C5201 a_2475_6170# a_16018_6146# 0.68fF
C5202 a_26058_7150# a_26058_6146# 0.84fF
C5203 a_20946_9158# rowon_n[7] 0.14fF
C5204 a_25358_9198# col_n[22] 0.11fF
C5205 a_9994_8154# rowoff_n[6] 2.28fF
C5206 a_20946_17190# rowoff_n[15] 0.54fF
C5207 a_19030_6146# rowoff_n[4] 1.84fF
C5208 a_2275_3158# a_6982_3134# 0.71fF
C5209 a_10998_9158# VDD 3.61fF
C5210 m3_1864_16138# ctop 0.22fF
C5211 a_2275_17214# col[22] 0.17fF
C5212 a_2475_8178# a_31078_8154# 0.68fF
C5213 a_16018_8154# a_17022_8154# 0.86fF
C5214 a_2275_6170# col[27] 0.17fF
C5215 a_2275_18218# col[7] 0.17fF
C5216 a_19030_7150# col[16] 0.38fF
C5217 a_17022_4138# vcm 0.89fF
C5218 a_28066_4138# rowoff_n[2] 1.40fF
C5219 a_7986_3134# rowon_n[1] 0.45fF
C5220 a_5886_17190# a_5978_17190# 0.45fF
C5221 a_2275_17214# a_7286_17230# 0.15fF
C5222 a_2475_17214# a_9902_17190# 0.41fF
C5223 a_1957_4162# m2_1732_3958# 0.33fF
C5224 a_2275_3158# VDD 3.18fF
C5225 a_34090_3134# col_n[31] 0.34fF
C5226 a_2275_5166# a_22042_5142# 0.71fF
C5227 a_2275_18218# a_17326_18234# 0.15fF
C5228 a_26058_13174# VDD 2.06fF
C5229 a_6982_10162# a_6982_9158# 0.84fF
C5230 rowon_n[10] sample_n 0.15fF
C5231 ctop col[8] 0.13fF
C5232 a_14314_7190# col_n[11] 0.11fF
C5233 a_32082_8154# vcm 0.89fF
C5234 a_19030_12170# row_n[10] 0.43fF
C5235 a_2475_2154# a_14922_2130# 0.41fF
C5236 a_2275_2154# a_12306_2170# 0.15fF
C5237 m2_30848_18014# m3_30980_18146# 4.43fF
C5238 a_18938_16186# rowon_n[14] 0.14fF
C5239 a_2475_10186# col[2] 0.22fF
C5240 a_6982_16186# VDD 4.02fF
C5241 a_29070_2130# row_n[0] 0.43fF
C5242 a_31078_12170# a_32082_12170# 0.86fF
C5243 a_28978_6146# rowon_n[4] 0.14fF
C5244 a_22346_2170# vcm 0.24fF
C5245 a_2275_16210# a_15926_16186# 0.17fF
C5246 a_7986_5142# col[5] 0.38fF
C5247 a_13006_11166# vcm 0.89fF
C5248 a_9902_1126# VDD 0.93fF
C5249 a_2275_16210# col_n[9] 0.17fF
C5250 a_18026_17190# col[15] 0.38fF
C5251 a_2475_4162# a_29982_4138# 0.41fF
C5252 a_2275_4162# a_27366_4178# 0.15fF
C5253 a_15926_4138# a_16018_4138# 0.45fF
C5254 a_2275_5166# col_n[14] 0.17fF
C5255 a_33086_13174# col_n[30] 0.34fF
C5256 a_5978_10162# rowon_n[8] 0.45fF
C5257 a_22042_14178# a_22042_13174# 0.84fF
C5258 a_2475_13198# a_7986_13174# 0.68fF
C5259 a_29982_10162# rowoff_n[8] 0.43fF
C5260 col[28] rowoff_n[12] 0.16fF
C5261 a_3270_5182# vcm 0.24fF
C5262 a_33086_13174# rowoff_n[11] 1.15fF
C5263 a_2275_2154# col[4] 0.17fF
C5264 a_13310_17230# col_n[10] 0.11fF
C5265 a_2275_1150# a_20946_1126# 0.17fF
C5266 a_28066_15182# vcm 0.89fF
C5267 a_24962_5142# VDD 0.29fF
C5268 m2_29844_946# VDD 3.25fF
C5269 a_2475_12194# col[19] 0.22fF
C5270 a_2475_1150# col[24] 0.22fF
C5271 a_12002_15182# a_13006_15182# 0.86fF
C5272 a_2475_15206# a_23046_15182# 0.68fF
C5273 a_18330_9198# vcm 0.24fF
C5274 a_2275_3158# a_34394_3174# 0.15fF
C5275 a_8990_18194# vcm 0.15fF
C5276 a_31078_4138# ctop 4.91fF
C5277 a_5886_8154# VDD 0.29fF
C5278 a_27062_9158# row_n[7] 0.43fF
C5279 a_2275_7174# col_n[31] 0.17fF
C5280 a_6982_15182# col[4] 0.38fF
C5281 a_30986_8154# a_31078_8154# 0.45fF
C5282 a_26970_13174# rowon_n[11] 0.14fF
C5283 col[12] rowoff_n[13] 0.27fF
C5284 a_2275_12194# a_14010_12170# 0.71fF
C5285 a_11910_3134# vcm 0.18fF
C5286 a_22042_11166# col_n[19] 0.34fF
C5287 a_2275_15206# col[16] 0.17fF
C5288 m2_28840_18014# m2_29844_18014# 0.86fF
C5289 a_33390_13214# vcm 0.24fF
C5290 a_2275_4162# col[21] 0.17fF
C5291 a_12002_7150# ctop 4.91fF
C5292 a_20946_12170# VDD 0.29fF
C5293 m2_33860_946# m2_34864_946# 0.55fF
C5294 a_2475_9182# a_6890_9158# 0.41fF
C5295 a_2275_9182# a_4274_9198# 0.15fF
C5296 a_3970_17190# rowon_n[15] 0.45fF
C5297 a_2275_14202# a_29070_14178# 0.71fF
C5298 a_2874_1126# m2_2736_946# 0.31fF
C5299 a_26970_7150# vcm 0.18fF
C5300 a_14010_7150# rowon_n[5] 0.45fF
C5301 a_21038_14178# rowoff_n[12] 1.74fF
C5302 a_2475_18218# col[27] 0.22fF
C5303 a_22042_2130# a_23046_2130# 0.86fF
C5304 a_14314_16226# vcm 0.24fF
C5305 a_2966_5142# row_n[3] 0.41fF
C5306 a_27062_11166# ctop 4.91fF
C5307 a_2275_9182# rowon_n[7] 1.99fF
C5308 a_2475_11190# a_21950_11166# 0.41fF
C5309 a_2275_11190# a_19334_11206# 0.15fF
C5310 a_11910_11166# a_12002_11166# 0.45fF
C5311 a_7894_10162# vcm 0.18fF
C5312 a_2275_17214# rowoff_n[15] 0.81fF
C5313 a_10998_9158# col_n[8] 0.34fF
C5314 a_25054_16186# row_n[14] 0.43fF
C5315 a_2966_9158# m2_3164_9406# 0.19fF
C5316 a_13006_4138# a_13006_3134# 0.84fF
C5317 a_2275_18218# col[18] 0.17fF
C5318 a_25054_17190# m2_25252_17438# 0.19fF
C5319 a_2275_8178# a_12914_8154# 0.17fF
C5320 a_7986_14178# ctop 4.91fF
C5321 a_35002_10162# rowon_n[8] 0.14fF
C5322 a_2275_13198# a_35398_13214# 0.15fF
C5323 a_2275_14202# col_n[3] 0.17fF
C5324 a_2275_3158# col_n[8] 0.17fF
C5325 a_22954_14178# vcm 0.18fF
C5326 a_19030_4138# VDD 2.78fF
C5327 a_2475_5166# a_4974_5142# 0.68fF
C5328 en_bit_n[2] col[16] 0.14fF
C5329 row_n[5] sample_n 0.16fF
C5330 ctop col[19] 0.13fF
C5331 a_31078_8154# col[28] 0.38fF
C5332 a_2275_10186# a_27974_10162# 0.17fF
C5333 a_2475_9182# rowoff_n[7] 4.75fF
C5334 a_12002_14178# rowon_n[12] 0.45fF
C5335 a_26970_15182# a_27062_15182# 0.45fF
C5336 a_8990_15182# rowoff_n[13] 2.33fF
C5337 a_22042_4138# rowon_n[2] 0.45fF
C5338 a_2475_10186# col[13] 0.22fF
C5339 a_26362_8194# col_n[23] 0.11fF
C5340 a_34090_8154# VDD 1.23fF
C5341 a_10998_7150# rowoff_n[5] 2.23fF
C5342 a_16018_15182# m2_16216_15430# 0.19fF
C5343 a_2475_7174# a_20034_7150# 0.68fF
C5344 a_28066_8154# a_28066_7150# 0.84fF
C5345 a_5978_2130# vcm 0.89fF
C5346 a_2275_16210# col_n[20] 0.17fF
C5347 a_2275_5166# col_n[25] 0.17fF
C5348 a_20034_5142# rowoff_n[3] 1.79fF
C5349 a_2275_4162# a_10998_4138# 0.71fF
C5350 a_33086_13174# row_n[11] 0.43fF
C5351 a_15014_11166# VDD 3.20fF
C5352 a_32994_17190# rowon_n[15] 0.14fF
C5353 a_18026_9158# a_19030_9158# 0.86fF
C5354 a_20034_6146# col[17] 0.38fF
C5355 a_2275_13198# col[10] 0.17fF
C5356 a_29070_3134# rowoff_n[1] 1.35fF
C5357 m2_27836_946# col[25] 0.51fF
C5358 a_2275_2154# col[15] 0.17fF
C5359 a_21038_6146# vcm 0.89fF
C5360 a_7894_18194# a_7986_18194# 0.11fF
C5361 a_2475_12194# col[30] 0.22fF
C5362 a_2275_6170# a_26058_6146# 0.71fF
C5363 a_6982_13174# m2_7180_13422# 0.19fF
C5364 a_30074_15182# VDD 1.65fF
C5365 a_15318_6186# col_n[12] 0.11fF
C5366 a_8990_11166# a_8990_10162# 0.84fF
C5367 a_25358_18234# col_n[22] 0.11fF
C5368 m2_24824_18014# vcm 0.71fF
C5369 a_2966_15182# a_3970_15182# 0.86fF
C5370 a_2275_15206# a_4882_15182# 0.17fF
C5371 a_20034_11166# rowon_n[9] 0.45fF
C5372 a_2475_9182# vcm 1.32fF
C5373 a_26058_9158# m2_26256_9406# 0.19fF
C5374 a_2475_3158# a_18938_3134# 0.41fF
C5375 a_2275_3158# a_16322_3174# 0.15fF
C5376 a_30074_2130# m2_29844_946# 0.84fF
C5377 a_2275_1150# m2_14784_946# 0.51fF
C5378 m3_13912_1078# ctop 0.21fF
C5379 col[23] rowoff_n[13] 0.19fF
C5380 VDD rowoff_n[0] 87.22fF
C5381 col_n[3] rowoff_n[6] 0.32fF
C5382 col_n[1] rowoff_n[4] 0.33fF
C5383 col_n[6] rowoff_n[9] 0.29fF
C5384 vcm rowoff_n[3] 2.43fF
C5385 col_n[4] rowoff_n[7] 0.31fF
C5386 col_n[0] rowoff_n[2] 0.34fF
C5387 col_n[5] rowoff_n[8] 0.30fF
C5388 sample rowoff_n[1] 0.22fF
C5389 col_n[2] rowoff_n[5] 0.32fF
C5390 a_33086_13174# a_34090_13174# 0.86fF
C5391 a_2275_15206# col[27] 0.17fF
C5392 a_26362_4178# vcm 0.24fF
C5393 a_8990_4138# col[6] 0.38fF
C5394 a_21950_11166# rowoff_n[9] 0.52fF
C5395 a_2275_17214# a_19942_17190# 0.17fF
C5396 a_19030_16186# col[16] 0.38fF
C5397 a_17022_13174# vcm 0.89fF
C5398 a_13918_3134# VDD 0.29fF
C5399 a_2475_5166# a_33998_5142# 0.41fF
C5400 a_2275_5166# a_31382_5182# 0.15fF
C5401 a_17934_5142# a_18026_5142# 0.45fF
C5402 a_7894_5142# rowon_n[3] 0.14fF
C5403 a_2275_12194# VDD 3.18fF
C5404 a_2275_18218# a_29982_18194# 0.17fF
C5405 a_34090_12170# col_n[31] 0.34fF
C5406 a_2275_1150# col_n[2] 0.17fF
C5407 a_30986_9158# rowoff_n[7] 0.42fF
C5408 a_4274_4178# col_n[1] 0.11fF
C5409 a_2475_14202# a_12002_14178# 0.68fF
C5410 a_24050_15182# a_24050_14178# 0.84fF
C5411 a_14314_16226# col_n[11] 0.11fF
C5412 a_7286_7190# vcm 0.24fF
C5413 a_2966_14178# rowoff_n[12] 2.62fF
C5414 a_17022_7150# m2_17220_7398# 0.19fF
C5415 a_2275_2154# a_24962_2130# 0.17fF
C5416 a_32082_17190# vcm 0.89fF
C5417 a_20034_2130# ctop 4.93fF
C5418 col[7] rowoff_n[14] 0.30fF
C5419 a_28978_7150# VDD 0.29fF
C5420 a_2275_11190# a_2874_11166# 0.17fF
C5421 a_2475_11190# a_3878_11166# 0.41fF
C5422 a_35002_2130# vcm 0.18fF
C5423 a_2475_8178# col[7] 0.22fF
C5424 a_2475_16210# a_27062_16186# 0.68fF
C5425 a_14010_16186# a_15014_16186# 0.86fF
C5426 a_22346_11206# vcm 0.24fF
C5427 a_2275_18218# col[29] 0.17fF
C5428 a_20434_1488# VDD 0.14fF
C5429 a_28066_8154# rowon_n[6] 0.45fF
C5430 a_7986_14178# col[5] 0.38fF
C5431 a_9902_10162# VDD 0.29fF
C5432 a_32994_9158# a_33086_9158# 0.45fF
C5433 a_2275_14202# col_n[14] 0.17fF
C5434 a_2275_3158# col_n[19] 0.17fF
C5435 a_23046_10162# col_n[20] 0.34fF
C5436 a_2275_13198# a_18026_13174# 0.71fF
C5437 a_15926_5142# vcm 0.18fF
C5438 m2_28264_2378# a_28066_2130# 0.19fF
C5439 a_9902_12170# rowoff_n[10] 0.66fF
C5440 a_2275_18218# m2_8760_18014# 0.51fF
C5441 VDD col_n[7] 14.72fF
C5442 vcm col_n[4] 3.22fF
C5443 ctop col[30] 0.13fF
C5444 a_7986_5142# m2_8184_5390# 0.19fF
C5445 a_5978_8154# row_n[6] 0.43fF
C5446 a_3270_14218# vcm 0.24fF
C5447 a_5886_12170# rowon_n[10] 0.14fF
C5448 a_35494_5504# VDD 0.13fF
C5449 a_2275_11190# col[4] 0.17fF
C5450 a_16018_9158# ctop 4.91fF
C5451 a_24962_14178# VDD 0.29fF
C5452 a_2275_10186# a_8290_10202# 0.15fF
C5453 a_2475_10186# a_10906_10162# 0.41fF
C5454 a_15926_2130# rowon_n[0] 0.14fF
C5455 a_2275_15206# a_33086_15182# 0.71fF
C5456 a_2475_10186# col[24] 0.22fF
C5457 m2_34864_10986# m2_35292_11414# 0.19fF
C5458 a_30986_9158# vcm 0.18fF
C5459 a_25966_16186# rowoff_n[14] 0.48fF
C5460 a_24050_3134# a_25054_3134# 0.86fF
C5461 a_18330_18234# vcm 0.25fF
C5462 a_2475_15206# m2_1732_15002# 0.16fF
C5463 a_31078_13174# ctop 4.91fF
C5464 a_5886_17190# VDD 0.29fF
C5465 a_2275_16210# col_n[31] 0.17fF
C5466 a_13918_12170# a_14010_12170# 0.45fF
C5467 a_2275_12194# a_23350_12210# 0.15fF
C5468 a_2475_12194# a_25966_12170# 0.41fF
C5469 m2_2736_946# VDD 7.29fF
C5470 a_12002_8154# col_n[9] 0.34fF
C5471 a_26058_15182# rowon_n[13] 0.45fF
C5472 a_11910_12170# vcm 0.18fF
C5473 a_1957_5166# rowoff_n[3] 0.14fF
C5474 a_7986_2130# VDD 3.92fF
C5475 a_15014_5142# a_15014_4138# 0.84fF
C5476 a_2275_13198# col[21] 0.17fF
C5477 a_2275_9182# a_16930_9158# 0.17fF
C5478 a_12914_18194# m2_12776_18014# 0.35fF
C5479 a_2275_2154# col[26] 0.17fF
C5480 a_12002_16186# ctop 4.91fF
C5481 a_2475_18218# m2_34864_18014# 0.55fF
C5482 a_3970_15182# row_n[13] 0.43fF
C5483 a_2966_6146# vcm 0.89fF
C5484 a_26970_16186# vcm 0.18fF
C5485 a_32082_7150# col[29] 0.38fF
C5486 a_23046_6146# VDD 2.37fF
C5487 a_14010_5142# row_n[3] 0.43fF
C5488 a_2475_6170# a_8990_6146# 0.68fF
C5489 a_4974_6146# a_5978_6146# 0.86fF
C5490 a_13918_9158# rowon_n[7] 0.14fF
C5491 a_2874_8154# rowoff_n[6] 0.74fF
C5492 a_2275_11190# a_31990_11166# 0.17fF
C5493 a_29070_1126# vcm 0.15fF
C5494 a_2275_7174# row_n[5] 26.41fF
C5495 a_28978_16186# a_29070_16186# 0.45fF
C5496 a_13918_17190# rowoff_n[15] 0.61fF
C5497 m2_28840_18014# VDD 2.54fF
C5498 a_27366_7190# col_n[24] 0.11fF
C5499 a_12002_6146# rowoff_n[4] 2.18fF
C5500 m3_9896_18146# ctop 0.21fF
C5501 a_3970_9158# VDD 4.33fF
C5502 col_n[12] rowoff_n[4] 0.25fF
C5503 col_n[15] rowoff_n[7] 0.23fF
C5504 col_n[8] rowoff_n[0] 0.28fF
C5505 col_n[11] rowoff_n[3] 0.26fF
C5506 col_n[14] rowoff_n[6] 0.24fF
C5507 col_n[9] rowoff_n[1] 0.27fF
C5508 col_n[16] rowoff_n[8] 0.22fF
C5509 col_n[13] rowoff_n[5] 0.24fF
C5510 col_n[10] rowoff_n[2] 0.27fF
C5511 col_n[17] rowoff_n[9] 0.21fF
C5512 a_30074_9158# a_30074_8154# 0.84fF
C5513 a_2475_8178# a_24050_8154# 0.68fF
C5514 a_2475_6170# col[1] 0.22fF
C5515 a_9994_4138# vcm 0.89fF
C5516 a_21038_4138# rowoff_n[2] 1.74fF
C5517 a_3878_11166# rowoff_n[9] 0.73fF
C5518 a_2275_12194# col_n[8] 0.17fF
C5519 a_34090_12170# rowon_n[10] 0.45fF
C5520 a_2275_5166# a_15014_5142# 0.71fF
C5521 a_2275_1150# col_n[13] 0.17fF
C5522 a_19030_13174# VDD 2.78fF
C5523 a_2275_18218# a_10298_18234# 0.15fF
C5524 a_21038_5142# col[18] 0.38fF
C5525 a_20034_10162# a_21038_10162# 0.86fF
C5526 a_31078_17190# col[28] 0.38fF
C5527 a_30074_2130# rowoff_n[0] 1.30fF
C5528 a_3270_1166# col_n[0] 0.11fF
C5529 a_25054_8154# vcm 0.89fF
C5530 col[18] rowoff_n[14] 0.23fF
C5531 a_12002_12170# row_n[10] 0.43fF
C5532 a_2966_7150# m2_1732_6970# 0.86fF
C5533 a_2475_2154# a_7894_2130# 0.41fF
C5534 a_2275_2154# a_5278_2170# 0.15fF
C5535 a_4882_2130# a_4974_2130# 0.45fF
C5536 col_n[1] rowoff_n[10] 0.33fF
C5537 a_11910_16186# rowon_n[14] 0.14fF
C5538 a_2275_7174# a_30074_7150# 0.71fF
C5539 a_16322_5182# col_n[13] 0.11fF
C5540 a_22042_2130# row_n[0] 0.43fF
C5541 a_26362_17230# col_n[23] 0.11fF
C5542 a_34090_17190# VDD 1.24fF
C5543 a_2475_8178# col[18] 0.22fF
C5544 a_10998_12170# a_10998_11166# 0.84fF
C5545 a_21950_6146# rowon_n[4] 0.14fF
C5546 a_15318_2170# vcm 0.24fF
C5547 a_2275_16210# a_8898_16186# 0.17fF
C5548 a_5978_11166# vcm 0.89fF
C5549 a_2161_1150# VDD 0.40fF
C5550 a_2275_14202# col_n[25] 0.17fF
C5551 a_2275_10186# m2_34864_9982# 0.51fF
C5552 a_2475_4162# a_22954_4138# 0.41fF
C5553 a_2275_4162# a_20338_4178# 0.15fF
C5554 a_2275_3158# col_n[30] 0.17fF
C5555 a_31990_18194# m2_31852_18014# 0.34fF
C5556 a_8990_17190# m2_8760_18014# 0.84fF
C5557 m2_1732_946# m2_2736_946# 0.86fF
C5558 a_9994_3134# col[7] 0.38fF
C5559 a_22954_10162# rowoff_n[8] 0.51fF
C5560 vcm col_n[15] 3.19fF
C5561 VDD col_n[18] 11.97fF
C5562 col[2] rowoff_n[15] 0.33fF
C5563 a_20034_15182# col[17] 0.38fF
C5564 a_30378_6186# vcm 0.24fF
C5565 a_26058_13174# rowoff_n[11] 1.50fF
C5566 a_2275_11190# col[15] 0.17fF
C5567 a_2275_1150# a_13918_1126# 0.17fF
C5568 a_21038_15182# vcm 0.89fF
C5569 a_17934_5142# VDD 0.29fF
C5570 a_19942_6146# a_20034_6146# 0.45fF
C5571 a_31990_8154# rowoff_n[6] 0.41fF
C5572 a_5278_3174# col_n[2] 0.11fF
C5573 m2_8760_18014# col[6] 0.37fF
C5574 a_15318_15222# col_n[12] 0.11fF
C5575 a_2475_15206# a_16018_15182# 0.68fF
C5576 a_26058_16186# a_26058_15182# 0.84fF
C5577 a_11302_9198# vcm 0.24fF
C5578 a_35002_9158# m2_34864_8978# 0.33fF
C5579 a_2275_3158# a_28978_3134# 0.17fF
C5580 a_24050_4138# ctop 4.91fF
C5581 a_20034_9158# row_n[7] 0.43fF
C5582 a_32994_9158# VDD 0.29fF
C5583 a_22042_16186# m2_22240_16434# 0.19fF
C5584 a_19942_13174# rowon_n[11] 0.14fF
C5585 a_2275_12194# a_6982_12170# 0.71fF
C5586 m2_34864_7974# row_n[6] 0.38fF
C5587 a_4882_3134# vcm 0.18fF
C5588 a_29982_3134# rowon_n[1] 0.14fF
C5589 a_2475_17214# a_31078_17190# 0.68fF
C5590 a_16018_17190# a_17022_17190# 0.86fF
C5591 m2_21812_18014# m2_22816_18014# 0.86fF
C5592 a_8990_13174# col[6] 0.38fF
C5593 a_26362_13214# vcm 0.24fF
C5594 a_4974_7150# ctop 4.91fF
C5595 a_13918_12170# VDD 0.29fF
C5596 m2_26832_946# m2_27260_1374# 0.19fF
C5597 a_35002_10162# a_35094_10162# 0.11fF
C5598 a_24050_9158# col_n[21] 0.34fF
C5599 a_2275_14202# a_22042_14178# 0.71fF
C5600 a_2275_10186# col_n[2] 0.17fF
C5601 a_19942_7150# vcm 0.18fF
C5602 a_6982_7150# rowon_n[5] 0.45fF
C5603 a_14010_14178# rowoff_n[12] 2.08fF
C5604 a_4274_13214# col_n[1] 0.11fF
C5605 a_1957_3158# sample 0.35fF
C5606 a_7286_16226# vcm 0.24fF
C5607 m2_24824_18014# col_n[22] 0.33fF
C5608 a_13006_14178# m2_13204_14426# 0.19fF
C5609 a_20034_11166# ctop 4.91fF
C5610 a_28978_16186# VDD 0.29fF
C5611 a_2275_11190# a_12306_11206# 0.15fF
C5612 a_2475_11190# a_14922_11166# 0.41fF
C5613 a_9994_2130# m2_10192_2378# 0.19fF
C5614 a_35002_11166# vcm 0.18fF
C5615 a_2475_17214# col[7] 0.22fF
C5616 col_n[27] rowoff_n[8] 0.14fF
C5617 col_n[20] rowoff_n[1] 0.19fF
C5618 col_n[23] rowoff_n[4] 0.17fF
C5619 col_n[26] rowoff_n[7] 0.15fF
C5620 col_n[21] rowoff_n[2] 0.19fF
C5621 col_n[24] rowoff_n[5] 0.16fF
C5622 col_n[28] rowoff_n[9] 0.14fF
C5623 col_n[25] rowoff_n[6] 0.16fF
C5624 col_n[22] rowoff_n[3] 0.18fF
C5625 a_18026_16186# row_n[14] 0.43fF
C5626 col_n[19] rowoff_n[0] 0.20fF
C5627 a_2475_6170# col[12] 0.22fF
C5628 a_32082_10162# m2_32280_10410# 0.19fF
C5629 a_26058_4138# a_27062_4138# 0.86fF
C5630 a_2275_8178# a_5886_8154# 0.17fF
C5631 a_28066_17190# m2_27836_18014# 0.84fF
C5632 a_28066_6146# row_n[4] 0.43fF
C5633 a_27974_10162# rowon_n[8] 0.14fF
C5634 a_15926_13174# a_16018_13174# 0.45fF
C5635 a_2475_13198# a_29982_13174# 0.41fF
C5636 a_2275_13198# a_27366_13214# 0.15fF
C5637 a_13006_7150# col_n[10] 0.34fF
C5638 a_2275_12194# col_n[19] 0.17fF
C5639 a_2966_4138# rowoff_n[2] 2.62fF
C5640 a_2275_1150# col_n[24] 0.17fF
C5641 a_15926_14178# vcm 0.18fF
C5642 a_12002_4138# VDD 3.51fF
C5643 a_17022_6146# a_17022_5142# 0.84fF
C5644 a_3970_12170# m2_4168_12418# 0.19fF
C5645 a_35494_14540# VDD 0.13fF
C5646 a_2275_10186# a_20946_10162# 0.17fF
C5647 a_2275_9182# col[9] 0.17fF
C5648 col[29] rowoff_n[14] 0.15fF
C5649 a_4974_14178# rowon_n[12] 0.45fF
C5650 col_n[12] rowoff_n[10] 0.25fF
C5651 a_2475_15206# rowoff_n[13] 4.75fF
C5652 m2_34864_11990# VDD 1.58fF
C5653 a_33086_6146# col[30] 0.38fF
C5654 a_15014_4138# rowon_n[2] 0.45fF
C5655 a_23046_8154# m2_23244_8402# 0.19fF
C5656 a_30986_18194# vcm 0.18fF
C5657 a_27062_8154# VDD 1.96fF
C5658 a_2475_8178# col[29] 0.22fF
C5659 a_3970_7150# rowoff_n[5] 2.57fF
C5660 a_2475_7174# a_13006_7150# 0.68fF
C5661 a_6982_7150# a_7986_7150# 0.86fF
C5662 a_2275_12194# a_34394_12210# 0.15fF
C5663 a_3878_6146# rowon_n[4] 0.14fF
C5664 a_33086_3134# vcm 0.89fF
C5665 a_30986_17190# a_31078_17190# 0.45fF
C5666 a_28370_6186# col_n[25] 0.11fF
C5667 a_13006_5142# rowoff_n[3] 2.13fF
C5668 a_12002_17190# col_n[9] 0.34fF
C5669 a_2275_4162# a_3970_4138# 0.71fF
C5670 a_26058_13174# row_n[11] 0.43fF
C5671 a_7986_11166# VDD 3.92fF
C5672 a_25966_17190# rowon_n[15] 0.14fF
C5673 a_32082_10162# a_32082_9158# 0.84fF
C5674 a_2475_9182# a_28066_9158# 0.68fF
C5675 vcm col_n[26] 3.22fF
C5676 VDD col_n[29] 9.25fF
C5677 col[13] rowoff_n[15] 0.26fF
C5678 a_2275_11190# col[26] 0.17fF
C5679 a_22042_3134# rowoff_n[1] 1.69fF
C5680 a_14010_6146# vcm 0.89fF
C5681 a_14010_6146# m2_14208_6394# 0.19fF
C5682 a_2966_15182# vcm 0.89fF
C5683 a_2275_6170# a_19030_6146# 0.71fF
C5684 a_22042_4138# col[19] 0.38fF
C5685 a_32082_16186# col[29] 0.38fF
C5686 a_23046_15182# VDD 2.37fF
C5687 a_22042_11166# a_23046_11166# 0.86fF
C5688 m2_10768_18014# vcm 0.71fF
C5689 a_13006_11166# rowon_n[9] 0.45fF
C5690 a_29070_10162# vcm 0.89fF
C5691 a_2475_3158# a_11910_3134# 0.41fF
C5692 a_2275_3158# a_9294_3174# 0.15fF
C5693 a_6890_3134# a_6982_3134# 0.45fF
C5694 a_17326_4178# col_n[14] 0.11fF
C5695 m3_34996_9110# ctop 0.22fF
C5696 a_1957_9182# row_n[7] 0.29fF
C5697 a_27366_16226# col_n[24] 0.11fF
C5698 a_2275_8178# a_34090_8154# 0.71fF
C5699 m2_11772_946# col[9] 0.51fF
C5700 a_13006_13174# a_13006_12170# 0.84fF
C5701 a_2475_15206# col[1] 0.22fF
C5702 a_19334_4178# vcm 0.24fF
C5703 a_2475_4162# col[6] 0.22fF
C5704 a_14922_11166# rowoff_n[9] 0.60fF
C5705 a_2275_17214# a_12914_17190# 0.17fF
C5706 a_4974_4138# m2_5172_4386# 0.19fF
C5707 a_9994_13174# vcm 0.89fF
C5708 a_6890_3134# VDD 0.29fF
C5709 a_2275_5166# a_24354_5182# 0.15fF
C5710 a_2475_5166# a_26970_5142# 0.41fF
C5711 a_2275_18218# a_22954_18194# 0.17fF
C5712 a_2275_10186# col_n[13] 0.17fF
C5713 a_34090_10162# row_n[8] 0.43fF
C5714 a_10998_2130# col[8] 0.38fF
C5715 a_23958_9158# rowoff_n[7] 0.50fF
C5716 a_21038_14178# col[18] 0.38fF
C5717 a_33998_14178# rowon_n[12] 0.14fF
C5718 a_2475_14202# a_4974_14178# 0.68fF
C5719 a_35398_8194# vcm 0.24fF
C5720 a_30986_15182# rowoff_n[13] 0.42fF
C5721 a_3270_10202# col_n[0] 0.11fF
C5722 a_2275_2154# a_17934_2130# 0.17fF
C5723 a_13006_2130# ctop 4.93fF
C5724 a_25054_17190# vcm 0.89fF
C5725 m2_1732_17010# m3_1864_17142# 4.42fF
C5726 a_2275_7174# col[3] 0.17fF
C5727 a_21950_7150# VDD 0.29fF
C5728 a_32994_7150# rowoff_n[5] 0.40fF
C5729 a_21950_7150# a_22042_7150# 0.45fF
C5730 a_6282_2170# col_n[3] 0.11fF
C5731 a_16322_14218# col_n[13] 0.11fF
C5732 a_27974_2130# vcm 0.18fF
C5733 a_2475_17214# col[18] 0.22fF
C5734 col_n[31] rowoff_n[1] 0.11fF
C5735 col_n[30] rowoff_n[0] 0.12fF
C5736 a_2475_16210# a_20034_16186# 0.68fF
C5737 a_28066_17190# a_28066_16186# 0.84fF
C5738 a_2475_6170# col[23] 0.22fF
C5739 a_15318_11206# vcm 0.24fF
C5740 a_13406_1488# VDD 0.16fF
C5741 a_21038_8154# rowon_n[6] 0.45fF
C5742 a_2275_4162# a_32994_4138# 0.17fF
C5743 a_28066_6146# ctop 4.91fF
C5744 a_2161_10186# VDD 0.23fF
C5745 m3_30980_1078# m3_31984_1078# 0.21fF
C5746 a_2275_12194# col_n[30] 0.17fF
C5747 a_2275_13198# a_10998_13174# 0.71fF
C5748 a_8898_5142# vcm 0.18fF
C5749 a_9994_12170# col[7] 0.38fF
C5750 a_2161_12194# rowoff_n[10] 0.14fF
C5751 a_2275_5166# m2_1732_4962# 0.27fF
C5752 a_30378_15222# vcm 0.24fF
C5753 a_8990_9158# ctop 4.91fF
C5754 a_2275_9182# col[20] 0.17fF
C5755 a_32082_17190# row_n[15] 0.43fF
C5756 a_25054_8154# col_n[22] 0.34fF
C5757 a_17934_14178# VDD 0.29fF
C5758 m2_1732_2954# rowoff_n[1] 2.46fF
C5759 a_8898_2130# rowon_n[0] 0.14fF
C5760 col_n[23] rowoff_n[10] 0.17fF
C5761 a_2275_15206# a_26058_15182# 0.71fF
C5762 a_5278_12210# col_n[2] 0.11fF
C5763 a_23958_9158# vcm 0.18fF
C5764 a_18938_16186# rowoff_n[14] 0.56fF
C5765 a_3970_3134# a_3970_2130# 0.84fF
C5766 a_11302_18234# vcm 0.25fF
C5767 a_21950_1126# m2_21812_946# 0.31fF
C5768 a_24050_13174# ctop 4.91fF
C5769 a_32994_18194# VDD 0.50fF
C5770 a_2275_12194# a_16322_12210# 0.15fF
C5771 a_2475_12194# a_18938_12170# 0.41fF
C5772 a_19030_15182# rowon_n[13] 0.45fF
C5773 m2_32856_18014# m2_33284_18442# 0.19fF
C5774 a_4882_12170# vcm 0.18fF
C5775 col_n[0] rowon_n[12] 0.17fF
C5776 VDD rowon_n[11] 4.61fF
C5777 col_n[5] rowon_n[15] 0.17fF
C5778 col_n[3] rowon_n[14] 0.17fF
C5779 vcm row_n[13] 1.08fF
C5780 col_n[4] row_n[15] 0.37fF
C5781 sample row_n[12] 0.92fF
C5782 col_n[1] rowon_n[13] 0.17fF
C5783 col_n[2] row_n[14] 0.37fF
C5784 a_28066_5142# a_29070_5142# 0.86fF
C5785 col[24] rowoff_n[15] 0.19fF
C5786 a_29070_5142# rowon_n[3] 0.45fF
C5787 a_2475_2154# col[0] 0.20fF
C5788 a_2275_9182# a_9902_9158# 0.17fF
C5789 a_4974_16186# ctop 4.91fF
C5790 col_n[7] rowoff_n[11] 0.29fF
C5791 a_14010_6146# col_n[11] 0.34fF
C5792 a_2475_18218# m2_20808_18014# 0.62fF
C5793 a_17934_14178# a_18026_14178# 0.45fF
C5794 a_2275_14202# a_31382_14218# 0.15fF
C5795 a_2475_14202# a_33998_14178# 0.41fF
C5796 a_34090_7150# m2_34864_6970# 0.86fF
C5797 a_19942_16186# vcm 0.18fF
C5798 a_2275_8178# col_n[7] 0.17fF
C5799 m2_1732_13998# m3_1864_14130# 4.42fF
C5800 a_16018_6146# VDD 3.09fF
C5801 a_6982_5142# row_n[3] 0.43fF
C5802 a_1957_12194# sample 0.35fF
C5803 a_19030_7150# a_19030_6146# 0.84fF
C5804 a_6890_9158# rowon_n[7] 0.14fF
C5805 a_2275_11190# a_24962_11166# 0.17fF
C5806 a_22042_1126# vcm 0.15fF
C5807 a_34090_5142# col[31] 0.38fF
C5808 m2_34864_1950# VDD 1.58fF
C5809 a_6890_17190# rowoff_n[15] 0.69fF
C5810 m2_14784_18014# VDD 4.08fF
C5811 a_4974_6146# rowoff_n[4] 2.52fF
C5812 a_13006_2130# m2_12776_946# 0.84fF
C5813 a_31078_10162# VDD 1.54fF
C5814 a_8990_8154# a_9994_8154# 0.86fF
C5815 a_2475_8178# a_17022_8154# 0.68fF
C5816 a_28066_17190# m2_28264_17438# 0.19fF
C5817 a_2475_15206# col[12] 0.22fF
C5818 a_2475_4162# col[17] 0.22fF
C5819 a_29374_5182# col_n[26] 0.11fF
C5820 a_2874_4138# vcm 0.18fF
C5821 a_14010_4138# rowoff_n[2] 2.08fF
C5822 a_32994_18194# a_33086_18194# 0.11fF
C5823 a_31078_12170# rowoff_n[10] 1.25fF
C5824 a_13006_16186# col_n[10] 0.34fF
C5825 a_27974_1126# a_28066_1126# 0.11fF
C5826 a_27062_12170# rowon_n[10] 0.45fF
C5827 a_2275_10186# col_n[24] 0.17fF
C5828 a_2275_5166# a_7986_5142# 0.71fF
C5829 a_12002_13174# VDD 3.51fF
C5830 a_2275_18218# a_3270_18234# 0.15fF
C5831 a_34090_11166# a_34090_10162# 0.84fF
C5832 a_2475_10186# a_32082_10162# 0.68fF
C5833 a_23046_2130# rowoff_n[0] 1.64fF
C5834 m2_34864_12994# vcm 0.72fF
C5835 a_18026_8154# vcm 0.89fF
C5836 a_2275_7174# col[14] 0.17fF
C5837 a_4974_12170# row_n[10] 0.43fF
C5838 a_23046_3134# col[20] 0.38fF
C5839 a_4882_16186# rowon_n[14] 0.14fF
C5840 a_3878_7150# VDD 0.29fF
C5841 a_33086_15182# col[30] 0.38fF
C5842 m2_34864_9982# rowon_n[8] 0.42fF
C5843 a_2275_7174# a_23046_7150# 0.71fF
C5844 a_19030_15182# m2_19228_15430# 0.19fF
C5845 a_27062_17190# VDD 1.96fF
C5846 a_15014_2130# row_n[0] 0.43fF
C5847 a_2475_17214# col[29] 0.22fF
C5848 rowon_n[7] rowoff_n[7] 20.66fF
C5849 a_24050_12170# a_25054_12170# 0.86fF
C5850 a_14922_6146# rowon_n[4] 0.14fF
C5851 a_8290_2170# vcm 0.24fF
C5852 a_2874_18194# VDD 0.50fF
C5853 a_33086_12170# vcm 0.89fF
C5854 a_18330_3174# col_n[15] 0.11fF
C5855 a_29982_2130# VDD 0.29fF
C5856 a_2966_8154# rowon_n[6] 0.45fF
C5857 a_2275_4162# a_13310_4178# 0.15fF
C5858 a_2475_4162# a_15926_4138# 0.41fF
C5859 a_28370_15222# col_n[25] 0.11fF
C5860 a_8898_4138# a_8990_4138# 0.45fF
C5861 m3_1864_4090# m3_1864_3086# 0.20fF
C5862 a_15014_14178# a_15014_13174# 0.84fF
C5863 a_15926_10162# rowoff_n[8] 0.59fF
C5864 a_23350_6186# vcm 0.24fF
C5865 a_19030_13174# rowoff_n[11] 1.84fF
C5866 a_2275_9182# col[31] 0.17fF
C5867 a_2275_1150# a_6890_1126# 0.17fF
C5868 a_14010_15182# vcm 0.89fF
C5869 m2_1732_10986# m3_1864_11118# 4.42fF
C5870 a_10906_5142# VDD 0.29fF
C5871 a_2275_6170# a_28370_6186# 0.15fF
C5872 a_2475_6170# a_30986_6146# 0.41fF
C5873 a_9994_13174# m2_10192_13422# 0.19fF
C5874 a_24962_8154# rowoff_n[6] 0.49fF
C5875 a_22042_13174# col[19] 0.38fF
C5876 a_2275_6170# col_n[1] 0.17fF
C5877 a_2475_15206# a_8990_15182# 0.68fF
C5878 a_4974_15182# a_5978_15182# 0.86fF
C5879 m2_1732_3958# sample 0.31fF
C5880 a_4274_9198# vcm 0.24fF
C5881 m2_1732_15002# VDD 5.46fF
C5882 a_2275_3158# a_21950_3134# 0.17fF
C5883 a_29070_9158# m2_29268_9406# 0.19fF
C5884 a_33998_6146# rowoff_n[4] 0.39fF
C5885 a_17022_4138# ctop 4.91fF
C5886 a_2275_1150# m2_23820_946# 0.51fF
C5887 m3_28972_1078# ctop 0.21fF
C5888 a_13006_9158# row_n[7] 0.43fF
C5889 a_25966_9158# VDD 0.29fF
C5890 a_7286_1166# col_n[4] 0.11fF
C5891 a_23958_8154# a_24050_8154# 0.45fF
C5892 a_17326_13214# col_n[14] 0.11fF
C5893 a_12914_13174# rowon_n[11] 0.14fF
C5894 m2_1732_11990# row_n[10] 0.44fF
C5895 a_31990_4138# vcm 0.18fF
C5896 a_22954_3134# rowon_n[1] 0.14fF
C5897 a_2475_17214# a_24050_17190# 0.68fF
C5898 col_n[6] rowon_n[10] 0.17fF
C5899 sample rowon_n[6] 0.10fF
C5900 col_n[4] rowon_n[9] 0.17fF
C5901 col_n[2] rowon_n[8] 0.17fF
C5902 col_n[9] row_n[12] 0.37fF
C5903 col_n[8] rowon_n[11] 0.17fF
C5904 col_n[16] rowon_n[15] 0.17fF
C5905 col_n[5] row_n[10] 0.37fF
C5906 col_n[14] rowon_n[14] 0.17fF
C5907 col_n[3] row_n[9] 0.37fF
C5908 col_n[12] rowon_n[13] 0.17fF
C5909 col_n[10] rowon_n[12] 0.17fF
C5910 col_n[1] row_n[8] 0.37fF
C5911 col_n[0] row_n[7] 0.37fF
C5912 vcm rowon_n[7] 0.91fF
C5913 col_n[11] row_n[13] 0.37fF
C5914 col_n[13] row_n[14] 0.37fF
C5915 VDD row_n[6] 4.64fF
C5916 col_n[15] row_n[15] 0.37fF
C5917 col_n[7] row_n[11] 0.37fF
C5918 m2_14784_18014# m2_15788_18014# 0.86fF
C5919 a_19334_13214# vcm 0.24fF
C5920 a_2475_13198# col[6] 0.22fF
C5921 a_2475_2154# col[11] 0.22fF
C5922 col_n[18] rowoff_n[11] 0.21fF
C5923 a_32082_8154# ctop 4.91fF
C5924 a_6890_12170# VDD 0.29fF
C5925 a_2275_14202# a_15014_14178# 0.71fF
C5926 a_10998_11166# col[8] 0.38fF
C5927 a_2275_8178# col_n[18] 0.17fF
C5928 a_12914_7150# vcm 0.18fF
C5929 a_6982_14178# rowoff_n[12] 2.42fF
C5930 a_2475_2154# a_29070_2130# 0.68fF
C5931 a_20034_7150# m2_20232_7398# 0.19fF
C5932 a_15014_2130# a_16018_2130# 0.86fF
C5933 a_35398_17230# vcm 0.24fF
C5934 a_33086_16186# rowon_n[14] 0.45fF
C5935 a_26058_7150# col_n[23] 0.34fF
C5936 a_13006_11166# ctop 4.91fF
C5937 m2_21812_946# col[19] 0.51fF
C5938 a_2275_16210# col[3] 0.17fF
C5939 a_21950_16186# VDD 0.29fF
C5940 a_4882_11166# a_4974_11166# 0.45fF
C5941 a_2275_11190# a_5278_11206# 0.15fF
C5942 a_2475_11190# a_7894_11166# 0.41fF
C5943 a_2275_5166# col[8] 0.17fF
C5944 a_6282_11206# col_n[3] 0.11fF
C5945 a_2275_16210# a_30074_16186# 0.71fF
C5946 m2_1732_13998# m2_2160_14426# 0.19fF
C5947 a_27974_11166# vcm 0.18fF
C5948 a_24050_1126# VDD 0.10fF
C5949 col_n[2] rowoff_n[12] 0.32fF
C5950 a_10998_16186# row_n[14] 0.43fF
C5951 a_2475_15206# col[23] 0.22fF
C5952 a_5978_4138# a_5978_3134# 0.84fF
C5953 a_2475_4162# col[28] 0.22fF
C5954 a_28066_15182# ctop 4.91fF
C5955 a_21038_6146# row_n[4] 0.43fF
C5956 a_2475_13198# a_22954_13174# 0.41fF
C5957 a_2275_13198# a_20338_13214# 0.15fF
C5958 a_20946_10162# rowon_n[8] 0.14fF
C5959 m2_31276_2378# a_31078_2130# 0.19fF
C5960 a_10998_5142# m2_11196_5390# 0.19fF
C5961 a_18026_1126# a_18330_1166# 0.10fF
C5962 a_8898_14178# vcm 0.18fF
C5963 m2_1732_7974# m3_1864_8106# 4.42fF
C5964 a_4974_4138# VDD 4.23fF
C5965 a_30074_6146# a_31078_6146# 0.86fF
C5966 a_15014_5142# col_n[12] 0.34fF
C5967 a_2275_10186# a_13918_10162# 0.17fF
C5968 a_25054_17190# col_n[22] 0.34fF
C5969 a_2275_7174# col[25] 0.17fF
C5970 a_19942_15182# a_20034_15182# 0.45fF
C5971 a_7986_4138# rowon_n[2] 0.45fF
C5972 a_2966_11166# col_n[0] 0.34fF
C5973 a_23958_18194# vcm 0.18fF
C5974 a_20034_8154# VDD 2.68fF
C5975 a_21038_8154# a_21038_7150# 0.84fF
C5976 a_2475_7174# a_5978_7150# 0.68fF
C5977 a_2275_12194# a_28978_12170# 0.17fF
C5978 a_26058_3134# vcm 0.89fF
C5979 a_1957_3158# m2_1732_2954# 0.33fF
C5980 m2_34864_18014# m2_34864_17010# 0.84fF
C5981 a_5978_5142# rowoff_n[3] 2.47fF
C5982 a_19030_13174# row_n[11] 0.43fF
C5983 m3_26964_18146# m3_27968_18146# 0.21fF
C5984 a_10998_9158# a_12002_9158# 0.86fF
C5985 a_18938_17190# rowon_n[15] 0.14fF
C5986 a_2475_9182# a_21038_9158# 0.68fF
C5987 a_3970_3134# col_n[1] 0.34fF
C5988 a_30378_4178# col_n[27] 0.11fF
C5989 a_2475_11190# col[0] 0.20fF
C5990 a_15014_3134# rowoff_n[1] 2.03fF
C5991 a_29070_3134# row_n[1] 0.43fF
C5992 a_14010_15182# col_n[11] 0.34fF
C5993 a_28978_7150# rowon_n[5] 0.14fF
C5994 a_6982_6146# vcm 0.89fF
C5995 a_29982_2130# a_30074_2130# 0.45fF
C5996 a_2275_6170# a_12002_6146# 0.71fF
C5997 a_2275_17214# col_n[7] 0.17fF
C5998 a_16018_15182# VDD 3.09fF
C5999 a_2275_6170# col_n[12] 0.17fF
C6000 a_31382_1166# vcm 0.25fF
C6001 a_5978_11166# rowon_n[9] 0.45fF
C6002 a_22042_10162# vcm 0.89fF
C6003 a_24050_2130# col[21] 0.38fF
C6004 a_2275_3158# a_3878_3134# 0.17fF
C6005 a_2475_3158# a_4882_3134# 0.41fF
C6006 a_34090_14178# col[31] 0.38fF
C6007 a_2275_3158# col[2] 0.17fF
C6008 m3_24956_18146# ctop 0.21fF
C6009 a_2275_8178# a_27062_8154# 0.71fF
C6010 VDD rowon_n[0] 4.61fF
C6011 col_n[2] row_n[3] 0.37fF
C6012 col_n[21] rowon_n[12] 0.17fF
C6013 col_n[17] rowon_n[10] 0.17fF
C6014 col_n[1] rowon_n[2] 0.17fF
C6015 col_n[0] rowon_n[1] 0.17fF
C6016 col_n[15] rowon_n[9] 0.17fF
C6017 col_n[13] rowon_n[8] 0.17fF
C6018 col_n[20] row_n[12] 0.37fF
C6019 col_n[24] row_n[14] 0.37fF
C6020 vcm row_n[2] 1.08fF
C6021 col_n[6] row_n[5] 0.37fF
C6022 col_n[4] row_n[4] 0.37fF
C6023 sample row_n[1] 0.92fF
C6024 col_n[22] row_n[13] 0.37fF
C6025 col_n[8] row_n[6] 0.37fF
C6026 col_n[26] row_n[15] 0.37fF
C6027 col_n[10] row_n[7] 0.37fF
C6028 col_n[3] rowon_n[3] 0.17fF
C6029 col_n[18] row_n[11] 0.37fF
C6030 col_n[12] row_n[8] 0.37fF
C6031 col_n[5] rowon_n[4] 0.17fF
C6032 col_n[23] rowon_n[13] 0.17fF
C6033 col_n[14] row_n[9] 0.37fF
C6034 col_n[7] rowon_n[5] 0.17fF
C6035 col_n[25] rowon_n[14] 0.17fF
C6036 col_n[16] row_n[10] 0.37fF
C6037 col_n[9] rowon_n[6] 0.17fF
C6038 col_n[27] rowon_n[15] 0.17fF
C6039 col_n[11] rowon_n[7] 0.17fF
C6040 col_n[19] rowon_n[11] 0.17fF
C6041 a_26058_13174# a_27062_13174# 0.86fF
C6042 a_2475_13198# col[17] 0.22fF
C6043 a_12306_4178# vcm 0.24fF
C6044 a_2275_17214# a_5886_17190# 0.17fF
C6045 a_7894_11166# rowoff_n[9] 0.68fF
C6046 a_2475_2154# col[22] 0.22fF
C6047 a_19334_2170# col_n[16] 0.11fF
C6048 col_n[29] rowoff_n[11] 0.13fF
C6049 a_2874_13174# vcm 0.18fF
C6050 a_29374_14218# col_n[26] 0.11fF
C6051 m2_1732_4962# m3_1864_5094# 4.42fF
C6052 a_33998_4138# VDD 0.29fF
C6053 a_10906_5142# a_10998_5142# 0.45fF
C6054 a_2275_5166# a_17326_5182# 0.15fF
C6055 a_2475_5166# a_19942_5142# 0.41fF
C6056 a_2275_18218# a_15926_18194# 0.17fF
C6057 a_27062_10162# row_n[8] 0.43fF
C6058 a_2275_8178# col_n[29] 0.17fF
C6059 a_16930_9158# rowoff_n[7] 0.58fF
C6060 a_26970_14178# rowon_n[12] 0.14fF
C6061 a_17022_15182# a_17022_14178# 0.84fF
C6062 a_27366_8194# vcm 0.24fF
C6063 a_23958_15182# rowoff_n[13] 0.50fF
C6064 a_2275_2154# a_10906_2130# 0.17fF
C6065 a_5978_2130# ctop 4.93fF
C6066 a_18026_17190# vcm 0.89fF
C6067 a_2275_16210# col[14] 0.17fF
C6068 a_14922_7150# VDD 0.29fF
C6069 a_25966_7150# rowoff_n[5] 0.48fF
C6070 a_2275_7174# a_32386_7190# 0.15fF
C6071 a_2475_7174# a_35002_7150# 0.41fF
C6072 a_2275_5166# col[19] 0.17fF
C6073 a_23046_12170# col[20] 0.38fF
C6074 a_3878_16186# VDD 0.29fF
C6075 a_20946_2130# vcm 0.18fF
C6076 col_n[13] rowoff_n[12] 0.24fF
C6077 a_2475_16210# a_13006_16186# 0.68fF
C6078 a_6982_16186# a_7986_16186# 0.86fF
C6079 a_35002_5142# rowoff_n[3] 0.38fF
C6080 a_8290_11206# vcm 0.24fF
C6081 a_6378_1488# VDD 0.18fF
C6082 a_14010_8154# rowon_n[6] 0.45fF
C6083 a_2275_4162# a_25966_4138# 0.17fF
C6084 a_21038_6146# ctop 4.91fF
C6085 a_18330_12210# col_n[15] 0.11fF
C6086 a_29982_11166# VDD 0.29fF
C6087 m3_16924_1078# m3_17928_1078# 0.21fF
C6088 a_25966_9158# a_26058_9158# 0.45fF
C6089 a_2966_6146# row_n[4] 0.41fF
C6090 a_2275_10186# rowon_n[8] 1.99fF
C6091 a_2275_13198# a_3970_13174# 0.71fF
C6092 a_34394_6186# vcm 0.24fF
C6093 a_2475_1150# a_18026_1126# 0.66fF
C6094 a_23350_15222# vcm 0.24fF
C6095 a_2475_18218# a_28978_18194# 0.41fF
C6096 a_25054_17190# row_n[15] 0.43fF
C6097 a_10906_14178# VDD 0.29fF
C6098 a_12002_10162# col[9] 0.38fF
C6099 VDD rowoff_n[13] 87.22fF
C6100 m2_1732_16006# vcm 1.11fF
C6101 a_2275_15206# a_19030_15182# 0.71fF
C6102 a_35002_11166# rowon_n[9] 0.14fF
C6103 a_16930_9158# vcm 0.18fF
C6104 ctop rowoff_n[3] 0.28fF
C6105 a_2275_15206# col_n[1] 0.17fF
C6106 row_n[0] rowoff_n[0] 0.64fF
C6107 col[0] rowoff_n[9] 0.34fF
C6108 a_11910_16186# rowoff_n[14] 0.64fF
C6109 a_27062_6146# col_n[24] 0.34fF
C6110 a_17022_3134# a_18026_3134# 0.86fF
C6111 a_2966_8154# m2_3164_8402# 0.19fF
C6112 a_2475_3158# a_33086_3134# 0.68fF
C6113 a_2275_4162# col_n[6] 0.17fF
C6114 a_4274_18234# vcm 0.25fF
C6115 a_1957_8178# VDD 0.28fF
C6116 a_25054_16186# m2_25252_16434# 0.19fF
C6117 a_17022_13174# ctop 4.91fF
C6118 a_25966_18194# VDD 0.50fF
C6119 a_7286_10202# col_n[4] 0.11fF
C6120 a_2966_8154# col[0] 0.38fF
C6121 a_6890_12170# a_6982_12170# 0.45fF
C6122 a_2475_12194# a_11910_12170# 0.41fF
C6123 a_2275_12194# a_9294_12210# 0.15fF
C6124 a_2275_17214# a_34090_17190# 0.71fF
C6125 a_12002_15182# rowon_n[13] 0.45fF
C6126 m2_25828_18014# m2_26256_18442# 0.19fF
C6127 a_31990_13174# vcm 0.18fF
C6128 m2_1732_1950# m3_1864_2082# 4.42fF
C6129 a_28066_3134# VDD 1.85fF
C6130 a_7986_5142# a_7986_4138# 0.84fF
C6131 a_22042_5142# rowon_n[3] 0.45fF
C6132 a_2475_11190# col[11] 0.22fF
C6133 a_2475_9182# a_2966_9158# 0.65fF
C6134 a_2161_9182# a_2275_9182# 0.17fF
C6135 a_32082_17190# ctop 4.93fF
C6136 a_2475_18218# m2_6752_18014# 0.62fF
C6137 a_2475_14202# a_26970_14178# 0.41fF
C6138 a_2275_14202# a_24354_14218# 0.15fF
C6139 a_2275_17214# col_n[18] 0.17fF
C6140 a_12914_16186# vcm 0.18fF
C6141 a_2275_6170# col_n[23] 0.17fF
C6142 a_8990_6146# VDD 3.82fF
C6143 a_16018_14178# m2_16216_14426# 0.19fF
C6144 a_32082_7150# a_33086_7150# 0.86fF
C6145 a_2275_18218# col_n[3] 0.17fF
C6146 a_16018_4138# col_n[13] 0.34fF
C6147 a_26058_16186# col_n[23] 0.34fF
C6148 a_33086_14178# row_n[12] 0.43fF
C6149 a_2275_11190# a_17934_11166# 0.17fF
C6150 a_15014_1126# vcm 0.15fF
C6151 a_21950_16186# a_22042_16186# 0.45fF
C6152 a_2275_14202# col[8] 0.17fF
C6153 a_13006_2130# m2_13204_2378# 0.19fF
C6154 a_2275_3158# col[13] 0.17fF
C6155 a_35398_1166# VDD 0.13fF
C6156 a_24050_10162# VDD 2.27fF
C6157 col_n[12] rowon_n[2] 0.17fF
C6158 col_n[19] row_n[6] 0.37fF
C6159 col_n[10] rowon_n[1] 0.17fF
C6160 col_n[17] row_n[5] 0.37fF
C6161 col_n[8] rowon_n[0] 0.17fF
C6162 col_n[15] row_n[4] 0.37fF
C6163 VDD col[1] 13.18fF
C6164 col_n[13] row_n[3] 0.37fF
C6165 col_n[11] row_n[2] 0.37fF
C6166 col_n[16] rowon_n[4] 0.17fF
C6167 col_n[23] row_n[8] 0.37fF
C6168 col_n[21] row_n[7] 0.37fF
C6169 col_n[14] rowon_n[3] 0.17fF
C6170 col_n[29] row_n[11] 0.37fF
C6171 col_n[25] row_n[9] 0.37fF
C6172 col_n[18] rowon_n[5] 0.17fF
C6173 col_n[27] row_n[10] 0.37fF
C6174 col_n[20] rowon_n[6] 0.17fF
C6175 col_n[22] rowon_n[7] 0.17fF
C6176 col_n[30] rowon_n[11] 0.17fF
C6177 col_n[31] row_n[12] 0.37fF
C6178 col_n[24] rowon_n[8] 0.17fF
C6179 col_n[26] rowon_n[9] 0.17fF
C6180 col_n[7] row_n[0] 0.37fF
C6181 col_n[28] rowon_n[10] 0.17fF
C6182 col_n[9] row_n[1] 0.37fF
C6183 m2_2736_18014# col[0] 0.39fF
C6184 a_23046_9158# a_23046_8154# 0.84fF
C6185 a_2475_8178# a_9994_8154# 0.68fF
C6186 a_2475_13198# col[28] 0.22fF
C6187 a_2275_13198# a_32994_13174# 0.17fF
C6188 rowon_n[11] rowoff_n[11] 20.66fF
C6189 a_30074_5142# vcm 0.89fF
C6190 a_24050_12170# rowoff_n[10] 1.59fF
C6191 a_6982_4138# rowoff_n[2] 2.42fF
C6192 a_20034_12170# rowon_n[10] 0.45fF
C6193 a_6982_12170# m2_7180_12418# 0.19fF
C6194 a_4974_13174# VDD 4.23fF
C6195 a_13006_10162# a_14010_10162# 0.86fF
C6196 a_2475_10186# a_25054_10162# 0.68fF
C6197 a_31382_3174# col_n[28] 0.11fF
C6198 a_4974_2130# col_n[2] 0.34fF
C6199 a_30074_2130# rowon_n[0] 0.45fF
C6200 a_16018_2130# rowoff_n[0] 1.98fF
C6201 a_15014_14178# col_n[12] 0.34fF
C6202 a_2275_16210# col[25] 0.17fF
C6203 a_10998_8154# vcm 0.89fF
C6204 a_2275_5166# col[30] 0.17fF
C6205 a_31990_3134# a_32082_3134# 0.45fF
C6206 a_26058_8154# m2_26256_8402# 0.19fF
C6207 m2_2736_18014# m3_2868_18146# 4.43fF
C6208 m2_1732_13998# rowon_n[12] 0.43fF
C6209 a_2275_7174# a_16018_7150# 0.71fF
C6210 a_7986_2130# row_n[0] 0.43fF
C6211 a_20034_17190# VDD 2.68fF
C6212 col_n[24] rowoff_n[12] 0.16fF
C6213 a_3970_12170# a_3970_11166# 0.84fF
C6214 a_7894_6146# rowon_n[4] 0.14fF
C6215 a_2275_2154# vcm 7.73fF
C6216 m2_18800_18014# col_n[16] 0.32fF
C6217 a_26058_12170# vcm 0.89fF
C6218 a_22954_2130# VDD 0.29fF
C6219 a_2275_4162# a_6282_4178# 0.15fF
C6220 a_2475_4162# a_8898_4138# 0.41fF
C6221 a_2966_6146# ctop 4.82fF
C6222 m3_1864_11118# m3_1864_10114# 0.20fF
C6223 a_2275_9182# a_31078_9158# 0.71fF
C6224 a_28066_14178# a_29070_14178# 0.86fF
C6225 a_8898_10162# rowoff_n[8] 0.67fF
C6226 m2_33860_946# analog_in 1.05fF
C6227 a_16322_6186# vcm 0.24fF
C6228 a_12002_13174# rowoff_n[11] 2.18fF
C6229 a_3970_12170# col_n[1] 0.34fF
C6230 a_30378_13214# col_n[27] 0.11fF
C6231 a_2475_9182# col[5] 0.22fF
C6232 a_17022_6146# m2_17220_6394# 0.19fF
C6233 a_6982_15182# vcm 0.89fF
C6234 a_12914_6146# a_13006_6146# 0.45fF
C6235 a_2275_6170# a_21342_6186# 0.15fF
C6236 a_2475_6170# a_23958_6146# 0.41fF
C6237 col_n[8] rowoff_n[13] 0.28fF
C6238 a_28066_9158# rowon_n[7] 0.45fF
C6239 a_17934_8154# rowoff_n[6] 0.57fF
C6240 col[4] rowoff_n[2] 0.32fF
C6241 col[3] rowoff_n[1] 0.33fF
C6242 col[2] rowoff_n[0] 0.33fF
C6243 col[5] rowoff_n[3] 0.31fF
C6244 col[6] rowoff_n[4] 0.31fF
C6245 col[7] rowoff_n[5] 0.30fF
C6246 col[8] rowoff_n[6] 0.29fF
C6247 col[9] rowoff_n[7] 0.29fF
C6248 col[10] rowoff_n[8] 0.28fF
C6249 col[11] rowoff_n[9] 0.27fF
C6250 a_2275_15206# col_n[12] 0.17fF
C6251 a_19030_16186# a_19030_15182# 0.84fF
C6252 a_2275_4162# col_n[17] 0.17fF
C6253 a_31382_10202# vcm 0.24fF
C6254 a_28066_17190# rowoff_n[15] 1.40fF
C6255 a_2275_3158# a_14922_3134# 0.17fF
C6256 a_26970_6146# rowoff_n[4] 0.47fF
C6257 a_9994_4138# ctop 4.91fF
C6258 a_24050_11166# col[21] 0.38fF
C6259 a_4882_1126# m2_4744_946# 0.31fF
C6260 a_2475_1150# m2_9764_946# 0.62fF
C6261 m3_34996_2082# ctop 0.22fF
C6262 a_5978_9158# row_n[7] 0.43fF
C6263 a_18938_9158# VDD 0.29fF
C6264 a_2966_8154# a_2966_7150# 0.84fF
C6265 a_5886_13174# rowon_n[11] 0.14fF
C6266 a_2275_12194# col[2] 0.17fF
C6267 a_2275_1150# col[7] 0.17fF
C6268 a_24962_4138# vcm 0.18fF
C6269 a_15926_3134# rowon_n[1] 0.14fF
C6270 a_2475_17214# a_17022_17190# 0.68fF
C6271 a_8990_17190# a_9994_17190# 0.86fF
C6272 a_7986_4138# m2_8184_4386# 0.19fF
C6273 m2_7756_18014# m2_8760_18014# 0.86fF
C6274 a_12306_13214# vcm 0.24fF
C6275 a_19334_11206# col_n[16] 0.11fF
C6276 a_2475_11190# col[22] 0.22fF
C6277 a_2275_5166# a_29982_5142# 0.17fF
C6278 a_25054_8154# ctop 4.91fF
C6279 a_33998_13174# VDD 0.29fF
C6280 a_27974_10162# a_28066_10162# 0.45fF
C6281 a_2275_14202# a_7986_14178# 0.71fF
C6282 a_2275_17214# col_n[29] 0.17fF
C6283 a_5886_7150# vcm 0.18fF
C6284 a_2275_18218# col_n[14] 0.17fF
C6285 a_29070_3134# a_29070_2130# 0.84fF
C6286 a_2475_2154# a_22042_2130# 0.68fF
C6287 a_27366_17230# vcm 0.24fF
C6288 a_26058_16186# rowon_n[14] 0.45fF
C6289 a_2475_14202# m2_1732_13998# 0.16fF
C6290 a_5978_11166# ctop 4.91fF
C6291 a_14922_16186# VDD 0.29fF
C6292 a_13006_9158# col[10] 0.38fF
C6293 a_2275_14202# col[19] 0.17fF
C6294 a_2275_3158# col[24] 0.17fF
C6295 a_2275_16210# a_23046_16186# 0.71fF
C6296 a_28066_5142# col_n[25] 0.34fF
C6297 a_20946_11166# vcm 0.18fF
C6298 col_n[29] rowon_n[5] 0.17fF
C6299 col_n[27] rowon_n[4] 0.17fF
C6300 col_n[25] rowon_n[3] 0.17fF
C6301 col_n[23] rowon_n[2] 0.17fF
C6302 col_n[30] row_n[6] 0.37fF
C6303 rowon_n[11] row_n[11] 21.02fF
C6304 col_n[21] rowon_n[1] 0.17fF
C6305 col_n[28] row_n[5] 0.37fF
C6306 VDD col[12] 10.46fF
C6307 col_n[31] rowon_n[6] 0.17fF
C6308 a_3970_16186# row_n[14] 0.43fF
C6309 col_n[18] row_n[0] 0.37fF
C6310 a_17022_1126# VDD 0.12fF
C6311 col_n[20] row_n[1] 0.37fF
C6312 vcm col[9] 6.66fF
C6313 col_n[4] col[5] 6.22fF
C6314 col_n[22] row_n[2] 0.37fF
C6315 col_n[24] row_n[3] 0.37fF
C6316 col_n[26] row_n[4] 0.37fF
C6317 col_n[19] rowon_n[0] 0.17fF
C6318 a_19030_4138# a_20034_4138# 0.86fF
C6319 a_8290_9198# col_n[5] 0.11fF
C6320 a_21038_15182# ctop 4.91fF
C6321 a_14010_6146# row_n[4] 0.43fF
C6322 a_13918_10162# rowon_n[8] 0.14fF
C6323 a_8898_13174# a_8990_13174# 0.45fF
C6324 a_2275_13198# a_13310_13214# 0.15fF
C6325 a_2475_13198# a_15926_13174# 0.41fF
C6326 m2_1732_3958# m2_1732_2954# 0.84fF
C6327 a_2275_1150# a_28066_1126# 0.14fF
C6328 a_2275_8178# row_n[6] 26.41fF
C6329 a_34394_15222# vcm 0.24fF
C6330 a_32082_5142# VDD 1.44fF
C6331 a_9994_6146# a_9994_5142# 0.84fF
C6332 m2_5748_946# col[3] 0.51fF
C6333 a_2275_10186# a_6890_10162# 0.17fF
C6334 a_2275_15206# a_28370_15222# 0.15fF
C6335 a_2475_15206# a_30986_15182# 0.41fF
C6336 a_17022_3134# col_n[14] 0.34fF
C6337 a_16930_18194# vcm 0.18fF
C6338 a_13006_8154# VDD 3.40fF
C6339 a_27062_15182# col_n[24] 0.34fF
C6340 a_2275_13198# col_n[6] 0.17fF
C6341 a_34090_13174# rowon_n[11] 0.45fF
C6342 a_2275_2154# col_n[11] 0.17fF
C6343 a_1957_17214# VDD 0.28fF
C6344 a_2275_12194# a_21950_12170# 0.17fF
C6345 a_19030_3134# vcm 0.89fF
C6346 a_2966_17190# col[0] 0.38fF
C6347 a_23958_17190# a_24050_17190# 0.45fF
C6348 a_2475_1150# col_n[31] 0.21fF
C6349 a_12002_13174# row_n[11] 0.43fF
C6350 a_28066_12170# VDD 1.85fF
C6351 m3_12908_18146# m3_13912_18146# 0.21fF
C6352 m2_8760_946# m3_8892_1078# 4.41fF
C6353 a_2475_9182# a_14010_9158# 0.68fF
C6354 a_25054_10162# a_25054_9158# 0.84fF
C6355 a_11910_17190# rowon_n[15] 0.14fF
C6356 a_22042_3134# row_n[1] 0.43fF
C6357 a_7986_3134# rowoff_n[1] 2.38fF
C6358 a_2475_9182# col[16] 0.22fF
C6359 a_21950_7150# rowon_n[5] 0.14fF
C6360 a_34090_7150# vcm 0.89fF
C6361 a_28978_14178# rowoff_n[12] 0.44fF
C6362 a_2966_6146# m2_1732_5966# 0.86fF
C6363 col_n[19] rowoff_n[13] 0.20fF
C6364 a_3878_6146# a_3970_6146# 0.45fF
C6365 a_2275_6170# a_4974_6146# 0.71fF
C6366 a_32386_2170# col_n[29] 0.11fF
C6367 col[22] rowoff_n[9] 0.20fF
C6368 col[21] rowoff_n[8] 0.21fF
C6369 col[20] rowoff_n[7] 0.21fF
C6370 col[19] rowoff_n[6] 0.22fF
C6371 col[18] rowoff_n[5] 0.23fF
C6372 col[17] rowoff_n[4] 0.23fF
C6373 col[16] rowoff_n[3] 0.24fF
C6374 col[15] rowoff_n[2] 0.25fF
C6375 col[14] rowoff_n[1] 0.25fF
C6376 col[13] rowoff_n[0] 0.26fF
C6377 a_2275_15206# col_n[23] 0.17fF
C6378 a_8990_15182# VDD 3.82fF
C6379 a_2475_11190# a_29070_11166# 0.68fF
C6380 a_16018_13174# col_n[13] 0.34fF
C6381 a_15014_11166# a_16018_11166# 0.86fF
C6382 a_2275_4162# col_n[28] 0.17fF
C6383 a_24354_1166# vcm 0.25fF
C6384 a_15014_10162# vcm 0.89fF
C6385 a_33998_4138# a_34090_4138# 0.45fF
C6386 a_2275_9182# m2_34864_8978# 0.51fF
C6387 a_2275_12194# col[13] 0.17fF
C6388 a_2275_1150# col[18] 0.16fF
C6389 a_31078_17190# m2_31276_17438# 0.19fF
C6390 a_2275_8178# a_20034_8154# 0.71fF
C6391 a_5978_13174# a_5978_12170# 0.84fF
C6392 a_5278_4178# vcm 0.24fF
C6393 col_n[3] rowoff_n[14] 0.32fF
C6394 a_30074_14178# vcm 0.89fF
C6395 a_26970_4138# VDD 0.29fF
C6396 a_2275_5166# a_10298_5182# 0.15fF
C6397 a_2475_5166# a_12914_5142# 0.41fF
C6398 col[6] rowoff_n[10] 0.31fF
C6399 a_2275_18218# a_8898_18194# 0.17fF
C6400 a_2275_10186# a_35094_10162# 0.14fF
C6401 a_20034_10162# row_n[8] 0.43fF
C6402 a_9902_9158# rowoff_n[7] 0.66fF
C6403 a_19942_14178# rowon_n[12] 0.14fF
C6404 a_30074_15182# a_31078_15182# 0.86fF
C6405 a_4974_11166# col_n[2] 0.34fF
C6406 a_2275_18218# col_n[25] 0.17fF
C6407 a_31382_12210# col_n[28] 0.11fF
C6408 a_20338_8194# vcm 0.24fF
C6409 a_16930_15182# rowoff_n[13] 0.58fF
C6410 a_2874_2130# a_2966_2130# 0.11fF
C6411 a_29982_4138# rowon_n[2] 0.14fF
C6412 a_35002_8154# m2_34864_7974# 0.33fF
C6413 a_33086_3134# ctop 4.91fF
C6414 a_10998_17190# vcm 0.89fF
C6415 a_7894_7150# VDD 0.29fF
C6416 a_2275_14202# col[30] 0.17fF
C6417 a_18938_7150# rowoff_n[5] 0.56fF
C6418 a_14922_7150# a_15014_7150# 0.45fF
C6419 a_22042_15182# m2_22240_15430# 0.19fF
C6420 a_2475_7174# a_27974_7150# 0.41fF
C6421 a_2275_7174# a_25358_7190# 0.15fF
C6422 a_13918_2130# vcm 0.18fF
C6423 vcm col[20] 6.66fF
C6424 col_n[31] row_n[1] 0.37fF
C6425 col_n[29] row_n[0] 0.37fF
C6426 col_n[30] rowon_n[0] 0.17fF
C6427 VDD col[23] 7.74fF
C6428 col_n[10] col[10] 0.50fF
C6429 a_21038_17190# a_21038_16186# 0.84fF
C6430 a_2475_16210# a_5978_16186# 0.68fF
C6431 a_27974_5142# rowoff_n[3] 0.46fF
C6432 a_2275_11190# vcm 7.71fF
C6433 a_25054_10162# col[22] 0.38fF
C6434 a_6982_8154# rowon_n[6] 0.45fF
C6435 a_2275_4162# a_18938_4138# 0.17fF
C6436 a_14010_6146# ctop 4.91fF
C6437 a_22954_11166# VDD 0.29fF
C6438 m3_2868_1078# m3_3872_1078# 0.13fF
C6439 a_2966_15182# ctop 4.82fF
C6440 m2_33860_18014# col[31] 0.39fF
C6441 a_28978_6146# vcm 0.18fF
C6442 a_20338_10202# col_n[17] 0.11fF
C6443 a_16322_15222# vcm 0.24fF
C6444 a_2475_18218# a_21950_18194# 0.41fF
C6445 m2_7756_946# VDD 6.55fF
C6446 a_13006_13174# m2_13204_13422# 0.19fF
C6447 a_2275_6170# a_33998_6146# 0.17fF
C6448 a_18026_17190# row_n[15] 0.43fF
C6449 a_29070_10162# ctop 4.91fF
C6450 a_2475_7174# col[10] 0.22fF
C6451 a_29982_11166# a_30074_11166# 0.45fF
C6452 m2_1732_2954# row_n[1] 0.44fF
C6453 a_28066_7150# row_n[5] 0.43fF
C6454 a_2275_15206# a_12002_15182# 0.71fF
C6455 a_27974_11166# rowon_n[9] 0.14fF
C6456 a_9902_9158# vcm 0.18fF
C6457 a_4882_16186# rowoff_n[14] 0.72fF
C6458 a_2275_13198# col_n[17] 0.17fF
C6459 a_31078_4138# a_31078_3134# 0.84fF
C6460 a_2475_3158# a_26058_3134# 0.68fF
C6461 a_32082_9158# m2_32280_9406# 0.19fF
C6462 a_2475_1150# m2_32856_946# 0.65fF
C6463 a_2275_2154# col_n[22] 0.17fF
C6464 a_14010_8154# col[11] 0.38fF
C6465 a_9994_13174# ctop 4.91fF
C6466 a_18938_18194# VDD 0.50fF
C6467 a_2475_12194# a_4882_12170# 0.41fF
C6468 a_2275_12194# a_3878_12170# 0.17fF
C6469 a_29070_4138# col_n[26] 0.34fF
C6470 a_2275_17214# a_27062_17190# 0.71fF
C6471 a_29070_11166# rowoff_n[9] 1.35fF
C6472 a_2275_10186# col[7] 0.17fF
C6473 a_4974_15182# rowon_n[13] 0.45fF
C6474 m2_18800_18014# m2_19228_18442# 0.19fF
C6475 a_24962_13174# vcm 0.18fF
C6476 a_21038_3134# VDD 2.58fF
C6477 a_9294_8194# col_n[6] 0.11fF
C6478 a_3970_11166# m2_4168_11414# 0.19fF
C6479 a_21038_5142# a_22042_5142# 0.86fF
C6480 a_15014_5142# rowon_n[3] 0.45fF
C6481 a_2475_9182# col[27] 0.22fF
C6482 a_25054_17190# ctop 4.93fF
C6483 a_2475_14202# a_19942_14178# 0.41fF
C6484 a_2275_14202# a_17326_14218# 0.15fF
C6485 a_10906_14178# a_10998_14178# 0.45fF
C6486 col_n[30] rowoff_n[13] 0.12fF
C6487 a_3878_7150# rowon_n[5] 0.14fF
C6488 a_2275_2154# a_32082_2130# 0.71fF
C6489 a_23046_7150# m2_23244_7398# 0.19fF
C6490 a_5886_16186# vcm 0.18fF
C6491 sample_n rowoff_n[8] 0.55fF
C6492 col[31] rowoff_n[7] 0.14fF
C6493 col[30] rowoff_n[6] 0.15fF
C6494 col[29] rowoff_n[5] 0.15fF
C6495 col[28] rowoff_n[4] 0.16fF
C6496 col[27] rowoff_n[3] 0.17fF
C6497 col[26] rowoff_n[2] 0.17fF
C6498 col[25] rowoff_n[1] 0.18fF
C6499 col[24] rowoff_n[0] 0.19fF
C6500 a_2475_6170# VDD 41.96fF
C6501 a_12002_7150# a_12002_6146# 0.84fF
C6502 a_26058_14178# row_n[12] 0.43fF
C6503 a_2275_11190# a_10906_11166# 0.17fF
C6504 a_7986_1126# vcm 0.15fF
C6505 a_2475_16210# a_35002_16186# 0.41fF
C6506 a_2275_16210# a_32386_16226# 0.15fF
C6507 a_2275_12194# col[24] 0.17fF
C6508 a_18026_2130# col_n[15] 0.33fF
C6509 a_2275_1150# col[29] 0.17fF
C6510 a_28066_14178# col_n[25] 0.34fF
C6511 a_17022_10162# VDD 2.99fF
C6512 a_1957_8178# a_2275_8178# 0.19fF
C6513 a_2475_8178# a_2874_8154# 0.41fF
C6514 a_8290_18234# col_n[5] 0.11fF
C6515 a_2275_13198# a_25966_13174# 0.17fF
C6516 col_n[14] rowoff_n[14] 0.24fF
C6517 a_23046_5142# vcm 0.89fF
C6518 a_17022_12170# rowoff_n[10] 1.94fF
C6519 m2_34288_2378# a_34090_2130# 0.19fF
C6520 a_25966_18194# a_26058_18194# 0.11fF
C6521 a_2275_18218# m2_23820_18014# 0.51fF
C6522 m2_26832_946# vcm 0.71fF
C6523 col[17] rowoff_n[10] 0.23fF
C6524 a_20946_1126# a_21038_1126# 0.11fF
C6525 a_14010_5142# m2_14208_5390# 0.19fF
C6526 a_13006_12170# rowon_n[10] 0.45fF
C6527 a_32082_14178# VDD 1.44fF
C6528 a_2475_10186# a_18026_10162# 0.68fF
C6529 a_27062_11166# a_27062_10162# 0.84fF
C6530 a_1957_10186# row_n[8] 0.29fF
C6531 a_8990_2130# rowoff_n[0] 2.33fF
C6532 a_23046_2130# rowon_n[0] 0.45fF
C6533 a_3970_8154# vcm 0.89fF
C6534 a_33086_16186# rowoff_n[14] 1.15fF
C6535 a_2475_5166# col[4] 0.22fF
C6536 a_2275_7174# a_8990_7150# 0.71fF
C6537 a_17022_12170# col_n[14] 0.34fF
C6538 a_13006_17190# VDD 3.41fF
C6539 vcm col[31] 6.41fF
C6540 sample rowoff_n[15] 0.23fF
C6541 row_n[13] ctop 0.28fF
C6542 col_n[15] col[16] 6.27fF
C6543 a_2475_12194# a_33086_12170# 0.68fF
C6544 a_17022_12170# a_18026_12170# 0.86fF
C6545 a_2275_11190# col_n[11] 0.17fF
C6546 a_34090_11166# row_n[9] 0.43fF
C6547 a_28370_3174# vcm 0.24fF
C6548 col[1] rowoff_n[11] 0.34fF
C6549 a_33998_15182# rowon_n[13] 0.14fF
C6550 a_4974_3134# m2_5172_3382# 0.19fF
C6551 a_19030_12170# vcm 0.89fF
C6552 a_15926_2130# VDD 0.29fF
C6553 a_17934_18194# m2_17796_18014# 0.34fF
C6554 a_2275_9182# a_24050_9158# 0.71fF
C6555 a_2275_8178# col[1] 0.17fF
C6556 a_7986_14178# a_7986_13174# 0.84fF
C6557 a_9294_6186# vcm 0.24fF
C6558 a_4974_13174# rowoff_n[11] 2.52fF
C6559 a_34090_16186# vcm 0.89fF
C6560 a_2475_18218# a_3878_18194# 0.41fF
C6561 a_2475_7174# col[21] 0.22fF
C6562 a_30986_6146# VDD 0.29fF
C6563 m2_34864_1950# row_n[0] 0.38fF
C6564 a_2475_6170# a_16930_6146# 0.41fF
C6565 a_2275_6170# a_14314_6186# 0.15fF
C6566 a_21038_9158# rowon_n[7] 0.45fF
C6567 a_10906_8154# rowoff_n[6] 0.65fF
C6568 a_5978_10162# col_n[3] 0.34fF
C6569 a_32386_11206# col_n[29] 0.11fF
C6570 a_32082_16186# a_33086_16186# 0.86fF
C6571 a_2275_13198# col_n[28] 0.17fF
C6572 a_24354_10202# vcm 0.24fF
C6573 a_21038_17190# rowoff_n[15] 1.74fF
C6574 a_2275_3158# a_7894_3134# 0.17fF
C6575 a_19942_6146# rowoff_n[4] 0.55fF
C6576 m3_1864_15134# ctop 0.22fF
C6577 a_11910_9158# VDD 0.29fF
C6578 a_2475_8178# a_31990_8154# 0.41fF
C6579 a_2275_8178# a_29374_8194# 0.15fF
C6580 a_16930_8154# a_17022_8154# 0.45fF
C6581 m2_31852_946# col_n[29] 0.49fF
C6582 a_2275_10186# col[18] 0.17fF
C6583 a_17934_4138# vcm 0.18fF
C6584 a_28978_4138# rowoff_n[2] 0.44fF
C6585 a_8898_3134# rowon_n[1] 0.14fF
C6586 a_2475_17214# a_9994_17190# 0.68fF
C6587 a_26058_9158# col[23] 0.38fF
C6588 a_2275_4162# m2_1732_3958# 0.27fF
C6589 a_5278_13214# vcm 0.24fF
C6590 a_2966_3134# VDD 4.45fF
C6591 a_2275_5166# a_22954_5142# 0.17fF
C6592 a_18026_8154# ctop 4.91fF
C6593 a_26970_13174# VDD 0.29fF
C6594 m2_34864_8978# m2_35292_9406# 0.19fF
C6595 a_21342_9198# col_n[18] 0.11fF
C6596 a_32994_8154# vcm 0.18fF
C6597 a_7986_2130# a_8990_2130# 0.86fF
C6598 a_2475_2154# a_15014_2130# 0.68fF
C6599 a_20338_17230# vcm 0.24fF
C6600 a_19030_16186# rowon_n[14] 0.45fF
C6601 a_33086_12170# ctop 4.91fF
C6602 a_7894_16186# VDD 0.29fF
C6603 a_31990_12170# a_32082_12170# 0.45fF
C6604 a_29070_6146# rowon_n[4] 0.45fF
C6605 a_2275_16210# a_16018_16186# 0.71fF
C6606 a_13918_11166# vcm 0.18fF
C6607 a_9994_1126# VDD 0.14fF
C6608 a_15014_7150# col[12] 0.38fF
C6609 a_2475_4162# a_30074_4138# 0.68fF
C6610 a_33086_5142# a_33086_4138# 0.84fF
C6611 a_2275_9182# col_n[5] 0.17fF
C6612 col_n[25] rowoff_n[14] 0.16fF
C6613 a_14010_17190# m2_13780_18014# 0.84fF
C6614 a_14010_15182# ctop 4.91fF
C6615 a_6982_6146# row_n[4] 0.43fF
C6616 a_2275_13198# a_6282_13214# 0.15fF
C6617 a_2475_13198# a_8898_13174# 0.41fF
C6618 a_6890_10162# rowon_n[8] 0.14fF
C6619 a_30074_3134# col_n[27] 0.34fF
C6620 a_30074_10162# rowoff_n[8] 1.30fF
C6621 col[28] rowoff_n[10] 0.16fF
C6622 a_33998_13174# rowoff_n[11] 0.39fF
C6623 a_2275_1150# a_21038_1126# 0.14fF
C6624 a_34090_6146# m2_34864_5966# 0.86fF
C6625 a_28978_15182# vcm 0.18fF
C6626 a_10298_7190# col_n[7] 0.11fF
C6627 a_25054_5142# VDD 2.16fF
C6628 m2_30848_946# VDD 3.10fF
C6629 a_23046_6146# a_24050_6146# 0.86fF
C6630 a_2475_16210# col[10] 0.22fF
C6631 a_12914_15182# a_13006_15182# 0.45fF
C6632 a_2275_15206# a_21342_15222# 0.15fF
C6633 a_2475_15206# a_23958_15182# 0.41fF
C6634 a_2475_5166# col[15] 0.22fF
C6635 a_9902_18194# vcm 0.18fF
C6636 col_n[9] rowoff_n[15] 0.27fF
C6637 a_5978_8154# VDD 4.13fF
C6638 rowon_n[7] ctop 0.37fF
C6639 col_n[21] col[21] 0.50fF
C6640 a_28066_16186# m2_28264_16434# 0.19fF
C6641 a_14010_8154# a_14010_7150# 0.84fF
C6642 a_3970_5142# col[1] 0.38fF
C6643 a_27062_13174# rowon_n[11] 0.45fF
C6644 a_2275_11190# col_n[22] 0.17fF
C6645 a_14010_17190# col[11] 0.38fF
C6646 col[12] rowoff_n[11] 0.27fF
C6647 a_2275_12194# a_14922_12170# 0.17fF
C6648 a_12002_3134# vcm 0.89fF
C6649 a_2966_17190# a_2966_16186# 0.84fF
C6650 a_19030_1126# col_n[16] 0.39fF
C6651 a_29070_13174# col_n[26] 0.34fF
C6652 a_2275_8178# col[12] 0.17fF
C6653 a_4974_13174# row_n[11] 0.43fF
C6654 a_21038_12170# VDD 2.58fF
C6655 m2_34864_946# m2_35292_1374# 0.19fF
C6656 a_9294_17230# col_n[6] 0.11fF
C6657 a_2475_9182# a_6982_9158# 0.68fF
C6658 a_4882_17190# rowon_n[15] 0.14fF
C6659 a_3970_9158# a_4974_9158# 0.86fF
C6660 a_2275_14202# a_29982_14178# 0.17fF
C6661 a_15014_3134# row_n[1] 0.43fF
C6662 a_14922_7150# rowon_n[5] 0.14fF
C6663 a_27062_7150# vcm 0.89fF
C6664 a_21950_14178# rowoff_n[12] 0.52fF
C6665 a_22954_2130# a_23046_2130# 0.45fF
C6666 a_19030_14178# m2_19228_14426# 0.19fF
C6667 a_2966_9158# rowon_n[7] 0.45fF
C6668 a_2475_15206# VDD 41.96fF
C6669 a_2475_11190# a_22042_11166# 0.68fF
C6670 a_29070_12170# a_29070_11166# 0.84fF
C6671 a_17326_1166# vcm 0.25fF
C6672 a_16018_2130# m2_16216_2378# 0.19fF
C6673 a_7986_10162# vcm 0.89fF
C6674 a_2966_17190# rowoff_n[15] 2.62fF
C6675 a_18026_11166# col_n[15] 0.34fF
C6676 a_2275_10186# col[29] 0.17fF
C6677 a_33086_17190# m2_32856_18014# 0.84fF
C6678 a_2275_8178# a_13006_8154# 0.71fF
C6679 a_19030_13174# a_20034_13174# 0.86fF
C6680 a_32386_5182# vcm 0.24fF
C6681 a_2275_7174# col_n[0] 0.17fF
C6682 a_23046_14178# vcm 0.89fF
C6683 a_19942_4138# VDD 0.29fF
C6684 m2_1732_4962# rowon_n[3] 0.43fF
C6685 a_2475_5166# a_5886_5142# 0.41fF
C6686 a_2275_5166# a_3270_5182# 0.15fF
C6687 a_9994_12170# m2_10192_12418# 0.19fF
C6688 a_2275_10186# a_28066_10162# 0.71fF
C6689 a_13006_10162# row_n[8] 0.43fF
C6690 a_2161_9182# rowoff_n[7] 0.14fF
C6691 a_2475_18218# a_2275_18218# 2.94fF
C6692 a_12914_14178# rowon_n[12] 0.14fF
C6693 a_9994_15182# a_9994_14178# 0.84fF
C6694 a_13310_8194# vcm 0.24fF
C6695 a_9902_15182# rowoff_n[13] 0.66fF
C6696 a_29070_8154# m2_29268_8402# 0.19fF
C6697 a_22954_4138# rowon_n[2] 0.14fF
C6698 a_3970_17190# vcm 0.89fF
C6699 a_26058_3134# ctop 4.91fF
C6700 m2_7756_18014# m3_7888_18146# 4.41fF
C6701 a_35002_8154# VDD 0.36fF
C6702 a_2475_14202# col[4] 0.22fF
C6703 a_11910_7150# rowoff_n[5] 0.64fF
C6704 a_2475_7174# a_20946_7150# 0.41fF
C6705 a_2275_7174# a_18330_7190# 0.15fF
C6706 a_2475_3158# col[9] 0.22fF
C6707 a_6982_9158# col_n[4] 0.34fF
C6708 a_33390_10202# col_n[30] 0.11fF
C6709 a_6890_2130# vcm 0.18fF
C6710 a_28370_12210# vcm 0.24fF
C6711 a_20946_5142# rowoff_n[3] 0.54fF
C6712 a_2275_9182# col_n[16] 0.17fF
C6713 a_2275_4162# a_11910_4138# 0.17fF
C6714 a_6982_6146# ctop 4.91fF
C6715 a_15926_11166# VDD 0.29fF
C6716 a_2275_9182# a_33390_9198# 0.15fF
C6717 a_33086_17190# rowon_n[15] 0.45fF
C6718 a_18938_9158# a_19030_9158# 0.45fF
C6719 a_29982_3134# rowoff_n[1] 0.43fF
C6720 a_2275_17214# col[1] 0.17fF
C6721 a_27062_8154# col[24] 0.38fF
C6722 a_21950_6146# vcm 0.18fF
C6723 a_2275_6170# col[6] 0.17fF
C6724 a_2275_1150# a_2966_1126# 0.14fF
C6725 a_20034_6146# m2_20232_6394# 0.19fF
C6726 a_2475_1150# a_3970_1126# 0.66fF
C6727 a_20034_2130# a_20034_1126# 0.84fF
C6728 a_9294_15222# vcm 0.24fF
C6729 a_2475_18218# a_14922_18194# 0.41fF
C6730 a_2275_6170# a_26970_6146# 0.17fF
C6731 a_10998_17190# row_n[15] 0.43fF
C6732 a_22042_10162# ctop 4.91fF
C6733 a_2475_16210# col[21] 0.22fF
C6734 a_30986_15182# VDD 0.29fF
C6735 a_2475_5166# col[26] 0.22fF
C6736 m2_25828_18014# vcm 0.71fF
C6737 a_22346_8194# col_n[19] 0.11fF
C6738 a_3878_15182# a_3970_15182# 0.45fF
C6739 a_2275_15206# a_4974_15182# 0.71fF
C6740 a_21038_7150# row_n[5] 0.43fF
C6741 a_20946_11166# rowon_n[9] 0.14fF
C6742 row_n[2] ctop 0.28fF
C6743 col_n[20] rowoff_n[15] 0.19fF
C6744 rowon_n[0] row_n[0] 21.02fF
C6745 col_n[26] col[27] 6.14fF
C6746 a_9994_3134# a_10998_3134# 0.86fF
C6747 a_2475_3158# a_19030_3134# 0.68fF
C6748 a_2275_1150# m2_15788_946# 0.51fF
C6749 m3_15920_1078# ctop 0.21fF
C6750 col[23] rowoff_n[11] 0.19fF
C6751 a_11910_18194# VDD 0.50fF
C6752 a_33998_13174# a_34090_13174# 0.45fF
C6753 a_22042_11166# rowoff_n[9] 1.69fF
C6754 a_2275_17214# a_20034_17190# 0.71fF
C6755 a_2275_8178# col[23] 0.17fF
C6756 m2_11772_18014# m2_12200_18442# 0.19fF
C6757 a_10998_4138# m2_11196_4386# 0.19fF
C6758 a_17934_13174# vcm 0.18fF
C6759 a_16018_6146# col[13] 0.38fF
C6760 a_14010_3134# VDD 3.30fF
C6761 a_2475_5166# a_34090_5142# 0.68fF
C6762 a_2966_12170# VDD 4.45fF
C6763 a_7986_5142# rowon_n[3] 0.45fF
C6764 a_2275_18218# a_30074_18194# 0.14fF
C6765 m2_14784_946# m2_15788_946# 0.86fF
C6766 a_31078_2130# col_n[28] 0.34fF
C6767 a_18026_17190# ctop 4.93fF
C6768 a_31078_9158# rowoff_n[7] 1.25fF
C6769 m2_12776_18014# col_n[10] 0.33fF
C6770 a_2475_14202# a_12914_14178# 0.41fF
C6771 a_2275_14202# a_10298_14218# 0.15fF
C6772 a_11302_6186# col_n[8] 0.11fF
C6773 a_3878_14178# rowoff_n[12] 0.73fF
C6774 m2_34864_7974# VDD 1.58fF
C6775 a_21342_18234# col_n[18] 0.11fF
C6776 a_2275_2154# a_25054_2130# 0.71fF
C6777 a_32994_17190# vcm 0.18fF
C6778 col[7] rowoff_n[12] 0.30fF
C6779 a_29070_7150# VDD 1.75fF
C6780 a_25054_7150# a_26058_7150# 0.86fF
C6781 a_19030_14178# row_n[12] 0.43fF
C6782 a_2874_11166# a_2966_11166# 0.45fF
C6783 a_35094_2130# vcm 0.15fF
C6784 a_14922_16186# a_15014_16186# 0.45fF
C6785 a_2275_16210# a_25358_16226# 0.15fF
C6786 a_2475_16210# a_27974_16186# 0.41fF
C6787 a_1957_2154# m2_1732_1950# 0.33fF
C6788 a_29070_4138# row_n[2] 0.43fF
C6789 a_2475_1150# col[3] 0.22fF
C6790 a_28978_8154# rowon_n[6] 0.14fF
C6791 a_4974_4138# col[2] 0.38fF
C6792 a_9994_10162# VDD 3.71fF
C6793 a_15014_16186# col[12] 0.38fF
C6794 a_16018_9158# a_16018_8154# 0.84fF
C6795 a_2275_13198# a_18938_13174# 0.17fF
C6796 a_2275_7174# col_n[10] 0.17fF
C6797 a_16018_5142# vcm 0.89fF
C6798 a_30074_12170# col_n[27] 0.34fF
C6799 a_9994_12170# rowoff_n[10] 2.28fF
C6800 a_2275_18218# m2_9764_18014# 0.51fF
C6801 a_2475_1150# a_32994_1126# 0.41fF
C6802 a_2275_1150# a_30378_1166# 0.15fF
C6803 a_35398_5182# VDD 0.12fF
C6804 a_5978_12170# rowon_n[10] 0.45fF
C6805 m3_34996_18146# VDD 0.12fF
C6806 a_10298_16226# col_n[7] 0.11fF
C6807 a_25054_14178# VDD 2.16fF
C6808 a_2475_10186# a_10998_10162# 0.68fF
C6809 a_2275_4162# col[0] 0.16fF
C6810 a_5978_10162# a_6982_10162# 0.86fF
C6811 a_2475_2154# rowoff_n[0] 4.75fF
C6812 a_16018_2130# rowon_n[0] 0.45fF
C6813 a_2275_15206# a_33998_15182# 0.17fF
C6814 a_1957_18218# a_2161_18218# 0.11fF
C6815 a_31078_9158# vcm 0.89fF
C6816 a_26058_16186# rowoff_n[14] 1.50fF
C6817 a_2475_14202# col[15] 0.22fF
C6818 a_24962_3134# a_25054_3134# 0.45fF
C6819 a_2475_3158# col[20] 0.22fF
C6820 a_26970_1126# m2_26832_946# 0.31fF
C6821 a_2475_7174# a_2275_7174# 2.96fF
C6822 a_1957_7174# a_2161_7174# 0.11fF
C6823 a_2475_18218# col[6] 0.22fF
C6824 a_5978_17190# VDD 4.13fF
C6825 a_31078_13174# a_31078_12170# 0.84fF
C6826 a_2475_12194# a_26058_12170# 0.68fF
C6827 a_3970_14178# col[1] 0.38fF
C6828 a_27062_11166# row_n[9] 0.43fF
C6829 a_21342_3174# vcm 0.24fF
C6830 a_2275_9182# col_n[27] 0.17fF
C6831 a_26970_15182# rowon_n[13] 0.14fF
C6832 a_2275_5166# rowoff_n[3] 0.81fF
C6833 a_12002_12170# vcm 0.89fF
C6834 a_8898_2130# VDD 0.29fF
C6835 a_19030_10162# col_n[16] 0.34fF
C6836 m2_13780_946# m3_13912_1078# 4.41fF
C6837 a_2275_9182# a_17022_9158# 0.71fF
C6838 a_2275_17214# col[12] 0.17fF
C6839 a_2275_6170# col[17] 0.17fF
C6840 a_21038_14178# a_22042_14178# 0.86fF
C6841 a_3878_6146# vcm 0.18fF
C6842 a_27062_16186# vcm 0.89fF
C6843 a_23958_6146# VDD 0.29fF
C6844 a_2475_6170# a_9902_6146# 0.41fF
C6845 a_2275_6170# a_7286_6186# 0.15fF
C6846 a_5886_6146# a_5978_6146# 0.45fF
C6847 a_14010_9158# rowon_n[7] 0.45fF
C6848 a_2275_11190# a_32082_11166# 0.71fF
C6849 rowon_n[15] sample_n 0.14fF
C6850 col_n[31] rowoff_n[15] 0.11fF
C6851 a_29982_1126# vcm 0.18fF
C6852 a_2966_7150# row_n[5] 0.41fF
C6853 a_12002_16186# a_12002_15182# 0.84fF
C6854 a_2275_11190# rowon_n[9] 1.99fF
C6855 a_17326_10202# vcm 0.24fF
C6856 a_14010_17190# rowoff_n[15] 2.08fF
C6857 m2_29844_18014# VDD 2.50fF
C6858 a_12914_6146# rowoff_n[4] 0.63fF
C6859 a_30074_5142# ctop 4.91fF
C6860 a_4882_9158# VDD 0.29fF
C6861 m3_11904_18146# ctop 0.21fF
C6862 a_7986_8154# col_n[5] 0.34fF
C6863 a_34090_17190# m2_34288_17438# 0.19fF
C6864 a_2475_8178# a_24962_8154# 0.41fF
C6865 a_2275_8178# a_22346_8194# 0.15fF
C6866 a_10906_4138# vcm 0.18fF
C6867 a_21950_4138# rowoff_n[2] 0.52fF
C6868 a_1957_17214# a_2275_17214# 0.19fF
C6869 a_2475_17214# a_2874_17190# 0.41fF
C6870 a_32386_14218# vcm 0.24fF
C6871 a_35002_12170# rowon_n[10] 0.14fF
C6872 a_2275_5166# a_15926_5142# 0.17fF
C6873 a_2275_16210# col_n[0] 0.17fF
C6874 a_10998_8154# ctop 4.91fF
C6875 a_19942_13174# VDD 0.29fF
C6876 a_2275_5166# col_n[4] 0.17fF
C6877 a_20946_10162# a_21038_10162# 0.45fF
C6878 a_30986_2130# rowoff_n[0] 0.42fF
C6879 a_28066_7150# col[25] 0.38fF
C6880 m2_1732_13998# sample_n 0.12fF
C6881 col[18] rowoff_n[12] 0.23fF
C6882 a_25966_8154# vcm 0.18fF
C6883 a_2966_7150# m2_3164_7398# 0.19fF
C6884 a_2475_2154# a_7986_2130# 0.68fF
C6885 a_22042_3134# a_22042_2130# 0.84fF
C6886 a_2275_2154# ctop 0.13fF
C6887 a_13310_17230# vcm 0.24fF
C6888 a_12002_16186# rowon_n[14] 0.45fF
C6889 a_25054_15182# m2_25252_15430# 0.19fF
C6890 a_2275_7174# a_30986_7150# 0.17fF
C6891 a_26058_12170# ctop 4.91fF
C6892 m2_15788_946# col_n[13] 0.45fF
C6893 a_35002_17190# VDD 0.36fF
C6894 a_23350_7190# col_n[20] 0.11fF
C6895 a_22042_6146# rowon_n[4] 0.45fF
C6896 a_2475_12194# col[9] 0.22fF
C6897 a_2475_1150# col[14] 0.22fF
C6898 a_2275_16210# a_8990_16186# 0.71fF
C6899 a_6890_11166# vcm 0.18fF
C6900 a_2874_1126# VDD 1.01fF
C6901 a_2475_4162# a_23046_4138# 0.68fF
C6902 a_12002_4138# a_13006_4138# 0.86fF
C6903 m2_34864_8978# rowoff_n[7] 1.01fF
C6904 a_2275_7174# col_n[21] 0.17fF
C6905 a_6982_15182# ctop 4.91fF
C6906 a_23046_10162# rowoff_n[8] 1.64fF
C6907 col[2] rowoff_n[13] 0.33fF
C6908 a_33086_15182# row_n[13] 0.43fF
C6909 a_17022_5142# col[14] 0.38fF
C6910 a_26970_13174# rowoff_n[11] 0.47fF
C6911 a_2275_1150# a_14010_1126# 0.14fF
C6912 a_27062_17190# col[24] 0.38fF
C6913 a_21950_15182# vcm 0.18fF
C6914 a_2275_15206# col[6] 0.17fF
C6915 a_18026_5142# VDD 2.89fF
C6916 a_2275_4162# col[11] 0.17fF
C6917 a_16018_13174# m2_16216_13422# 0.19fF
C6918 a_32082_8154# rowoff_n[6] 1.20fF
C6919 a_2275_15206# a_14314_15222# 0.15fF
C6920 a_2475_15206# a_16930_15182# 0.41fF
C6921 a_2475_14202# col[26] 0.22fF
C6922 a_12306_5182# col_n[9] 0.11fF
C6923 a_2475_3158# col[31] 0.22fF
C6924 a_22346_17230# col_n[19] 0.11fF
C6925 a_2475_18218# col[17] 0.22fF
C6926 a_2275_3158# a_29070_3134# 0.71fF
C6927 a_33086_9158# VDD 1.34fF
C6928 a_27062_8154# a_28066_8154# 0.86fF
C6929 a_20034_13174# rowon_n[11] 0.45fF
C6930 a_2275_12194# a_7894_12170# 0.17fF
C6931 a_4974_3134# vcm 0.89fF
C6932 a_30074_3134# rowon_n[1] 0.45fF
C6933 a_2275_17214# a_29374_17230# 0.15fF
C6934 a_2475_17214# a_31990_17190# 0.41fF
C6935 a_16930_17190# a_17022_17190# 0.45fF
C6936 a_5978_3134# col[3] 0.38fF
C6937 a_2275_17214# col[23] 0.17fF
C6938 a_6982_11166# m2_7180_11414# 0.19fF
C6939 a_16018_15182# col[13] 0.38fF
C6940 a_2275_6170# col[28] 0.17fF
C6941 a_14010_12170# VDD 3.30fF
C6942 a_2275_18218# col[8] 0.17fF
C6943 a_18026_10162# a_18026_9158# 0.84fF
C6944 m2_34864_8978# vcm 0.72fF
C6945 a_2275_14202# a_22954_14178# 0.17fF
C6946 a_7986_3134# row_n[1] 0.43fF
C6947 a_31078_11166# col_n[28] 0.34fF
C6948 a_20034_7150# vcm 0.89fF
C6949 a_7894_7150# rowon_n[5] 0.14fF
C6950 a_14922_14178# rowoff_n[12] 0.60fF
C6951 a_26058_7150# m2_26256_7398# 0.19fF
C6952 a_2275_2154# a_35398_2170# 0.15fF
C6953 a_11302_15222# col_n[8] 0.11fF
C6954 m2_34864_16006# m3_34996_16138# 4.48fF
C6955 ctop col[9] 0.13fF
C6956 row_n[10] sample_n 0.16fF
C6957 a_29070_16186# VDD 1.75fF
C6958 m2_27836_18014# col[25] 0.37fF
C6959 a_2475_11190# a_15014_11166# 0.68fF
C6960 a_7986_11166# a_8990_11166# 0.86fF
C6961 a_10298_1166# vcm 0.25fF
C6962 a_35094_11166# vcm 0.15fF
C6963 a_31990_1126# VDD 0.68fF
C6964 a_26970_4138# a_27062_4138# 0.45fF
C6965 a_2475_10186# col[3] 0.22fF
C6966 a_2275_8178# a_5978_8154# 0.71fF
C6967 a_4974_13174# col[2] 0.38fF
C6968 a_28066_10162# rowon_n[8] 0.45fF
C6969 a_2475_13198# a_30074_13174# 0.68fF
C6970 a_33086_14178# a_33086_13174# 0.84fF
C6971 a_25358_5182# vcm 0.24fF
C6972 a_3878_4138# rowoff_n[2] 0.73fF
C6973 m2_34864_946# vcm 0.72fF
C6974 a_20034_9158# col_n[17] 0.34fF
C6975 a_2275_16210# col_n[10] 0.17fF
C6976 a_17022_5142# m2_17220_5390# 0.19fF
C6977 a_16018_14178# vcm 0.89fF
C6978 a_2275_5166# col_n[15] 0.17fF
C6979 a_12914_4138# VDD 0.29fF
C6980 a_35398_14218# VDD 0.12fF
C6981 a_2275_10186# a_21038_10162# 0.71fF
C6982 a_5978_10162# row_n[8] 0.43fF
C6983 col[29] rowoff_n[12] 0.15fF
C6984 a_5886_14178# rowon_n[12] 0.14fF
C6985 a_2275_13198# col[0] 0.16fF
C6986 a_23046_15182# a_24050_15182# 0.86fF
C6987 a_2275_2154# col[5] 0.17fF
C6988 a_6282_8194# vcm 0.24fF
C6989 a_2161_15206# rowoff_n[13] 0.14fF
C6990 m2_1732_10986# VDD 5.46fF
C6991 a_15926_4138# rowon_n[2] 0.14fF
C6992 a_19030_3134# ctop 4.91fF
C6993 a_31078_18194# vcm 0.15fF
C6994 a_35002_1126# m2_34864_946# 0.30fF
C6995 a_27974_8154# VDD 0.29fF
C6996 a_4882_7150# rowoff_n[5] 0.72fF
C6997 a_2475_7174# a_13918_7150# 0.41fF
C6998 a_2275_7174# a_11302_7190# 0.15fF
C6999 a_7894_7150# a_7986_7150# 0.45fF
C7000 a_2475_12194# col[20] 0.22fF
C7001 a_2475_1150# col[25] 0.22fF
C7002 a_33998_3134# vcm 0.18fF
C7003 a_14010_17190# a_14010_16186# 0.84fF
C7004 a_7986_3134# m2_8184_3382# 0.19fF
C7005 a_13918_5142# rowoff_n[3] 0.61fF
C7006 a_21342_12210# vcm 0.24fF
C7007 a_2275_4162# a_4882_4138# 0.17fF
C7008 a_2966_4138# a_3970_4138# 0.86fF
C7009 a_8990_7150# col_n[6] 0.34fF
C7010 a_34090_7150# ctop 4.80fF
C7011 a_8898_11166# VDD 0.29fF
C7012 a_26058_17190# rowon_n[15] 0.45fF
C7013 a_2275_9182# a_26362_9198# 0.15fF
C7014 a_2475_9182# a_28978_9158# 0.41fF
C7015 col[13] rowoff_n[13] 0.26fF
C7016 a_22954_3134# rowoff_n[1] 0.51fF
C7017 a_2275_15206# col[17] 0.17fF
C7018 a_14922_6146# vcm 0.18fF
C7019 a_2275_4162# col[22] 0.17fF
C7020 a_33086_2130# a_34090_2130# 0.86fF
C7021 a_3878_15182# vcm 0.18fF
C7022 a_2475_18218# a_7894_18194# 0.41fF
C7023 m2_34864_12994# m3_34996_13126# 4.42fF
C7024 a_2275_6170# a_19942_6146# 0.17fF
C7025 a_2475_13198# m2_1732_12994# 0.16fF
C7026 a_15014_10162# ctop 4.91fF
C7027 a_3970_17190# row_n[15] 0.43fF
C7028 a_23958_15182# VDD 0.29fF
C7029 a_22954_11166# a_23046_11166# 0.45fF
C7030 a_29070_6146# col[26] 0.38fF
C7031 m2_11772_18014# vcm 0.71fF
C7032 a_14010_7150# row_n[5] 0.43fF
C7033 a_2475_18218# col[28] 0.22fF
C7034 m2_1732_11990# m2_2160_12418# 0.19fF
C7035 a_13918_11166# rowon_n[9] 0.14fF
C7036 a_29982_10162# vcm 0.18fF
C7037 a_2475_3158# a_12002_3134# 0.68fF
C7038 a_24050_4138# a_24050_3134# 0.84fF
C7039 a_2275_9182# row_n[7] 26.41fF
C7040 m3_34996_8106# ctop 0.22fF
C7041 a_2275_8178# a_35002_8154# 0.17fF
C7042 a_24354_6186# col_n[21] 0.11fF
C7043 a_30074_14178# ctop 4.91fF
C7044 a_4882_18194# VDD 0.50fF
C7045 a_7986_17190# col_n[5] 0.34fF
C7046 a_15014_11166# rowoff_n[9] 2.03fF
C7047 a_2275_17214# a_13006_17190# 0.71fF
C7048 m2_4744_18014# m2_5172_18442# 0.19fF
C7049 a_10906_13174# vcm 0.18fF
C7050 a_6982_3134# VDD 4.02fF
C7051 a_2275_18218# col[19] 0.17fF
C7052 a_2475_5166# a_27062_5142# 0.68fF
C7053 a_14010_5142# a_15014_5142# 0.86fF
C7054 a_2275_18218# a_23046_18194# 0.14fF
C7055 m2_7756_946# m2_8760_946# 0.86fF
C7056 a_10998_17190# ctop 4.93fF
C7057 a_24050_9158# rowoff_n[7] 1.59fF
C7058 a_2275_14202# col_n[4] 0.17fF
C7059 a_34090_14178# rowon_n[12] 0.45fF
C7060 a_2475_14202# a_5886_14178# 0.41fF
C7061 a_2275_14202# a_3270_14218# 0.15fF
C7062 a_18026_4138# col[15] 0.38fF
C7063 a_2275_3158# col_n[9] 0.17fF
C7064 a_1957_7174# vcm 0.16fF
C7065 a_28066_16186# col[25] 0.38fF
C7066 a_31078_15182# rowoff_n[13] 1.25fF
C7067 a_2275_2154# a_18026_2130# 0.71fF
C7068 a_25966_17190# vcm 0.18fF
C7069 rowon_n[4] sample_n 0.15fF
C7070 ctop col[20] 0.13fF
C7071 a_22042_7150# VDD 2.47fF
C7072 a_33086_7150# rowoff_n[5] 1.15fF
C7073 a_4974_7150# a_4974_6146# 0.84fF
C7074 a_2275_11190# ctop 0.14fF
C7075 a_12002_14178# row_n[12] 0.43fF
C7076 a_13310_4178# col_n[10] 0.11fF
C7077 a_28066_2130# vcm 0.89fF
C7078 a_23350_16226# col_n[20] 0.11fF
C7079 a_2275_16210# a_18330_16226# 0.15fF
C7080 a_2475_16210# a_20946_16186# 0.41fF
C7081 m2_34864_16006# m2_34864_15002# 0.84fF
C7082 a_22042_4138# row_n[2] 0.43fF
C7083 a_2475_10186# col[14] 0.22fF
C7084 a_21950_8154# rowon_n[6] 0.14fF
C7085 a_2275_4162# a_33086_4138# 0.71fF
C7086 a_2874_10162# VDD 0.29fF
C7087 m3_31984_1078# m3_32988_1078# 0.21fF
C7088 a_29070_9158# a_30074_9158# 0.86fF
C7089 a_2275_13198# a_11910_13174# 0.17fF
C7090 a_2275_16210# col_n[21] 0.17fF
C7091 a_8990_5142# vcm 0.89fF
C7092 a_2275_5166# col_n[26] 0.17fF
C7093 a_18938_18194# a_19030_18194# 0.11fF
C7094 a_2874_12170# rowoff_n[10] 0.74fF
C7095 a_6982_2130# col[4] 0.38fF
C7096 a_2475_1150# a_25966_1126# 0.41fF
C7097 a_13918_1126# a_14010_1126# 0.11fF
C7098 a_2966_5142# m2_1732_4962# 0.86fF
C7099 a_2275_1150# a_23350_1166# 0.15fF
C7100 m2_34864_9982# m3_34996_10114# 4.42fF
C7101 a_17022_14178# col[14] 0.38fF
C7102 m2_25828_946# col_n[23] 0.45fF
C7103 m3_6884_18146# VDD 0.10fF
C7104 a_18026_14178# VDD 2.89fF
C7105 a_2275_13198# col[11] 0.17fF
C7106 a_20034_11166# a_20034_10162# 0.84fF
C7107 a_2475_10186# a_3970_10162# 0.68fF
C7108 a_2275_10186# a_2966_10162# 0.67fF
C7109 a_32082_10162# col_n[29] 0.34fF
C7110 a_2275_2154# col[16] 0.17fF
C7111 a_8990_2130# rowon_n[0] 0.45fF
C7112 a_2275_15206# a_26970_15182# 0.17fF
C7113 a_24050_9158# vcm 0.89fF
C7114 a_19030_16186# rowoff_n[14] 1.84fF
C7115 a_12306_14218# col_n[9] 0.11fF
C7116 a_2475_12194# col[31] 0.22fF
C7117 a_2275_8178# m2_34864_7974# 0.51fF
C7118 a_31078_16186# m2_31276_16434# 0.19fF
C7119 a_9994_12170# a_10998_12170# 0.86fF
C7120 a_2475_12194# a_19030_12170# 0.68fF
C7121 a_14314_3174# vcm 0.24fF
C7122 a_20034_11166# row_n[9] 0.43fF
C7123 a_19942_15182# rowon_n[13] 0.14fF
C7124 a_4974_12170# vcm 0.89fF
C7125 col[24] rowoff_n[13] 0.19fF
C7126 a_28978_5142# a_29070_5142# 0.45fF
C7127 a_5978_12170# col[3] 0.38fF
C7128 a_29982_5142# rowon_n[3] 0.14fF
C7129 a_2275_9182# a_9994_9158# 0.71fF
C7130 col_n[0] rowoff_n[1] 0.34fF
C7131 col_n[4] rowoff_n[6] 0.31fF
C7132 vcm rowoff_n[2] 2.43fF
C7133 col_n[7] rowoff_n[9] 0.29fF
C7134 col_n[2] rowoff_n[4] 0.32fF
C7135 sample rowoff_n[0] 0.22fF
C7136 col_n[5] rowoff_n[7] 0.30fF
C7137 col_n[6] rowoff_n[8] 0.29fF
C7138 col_n[1] rowoff_n[3] 0.33fF
C7139 col_n[3] rowoff_n[5] 0.32fF
C7140 a_2275_15206# col[28] 0.17fF
C7141 a_2475_18218# m2_21812_18014# 0.62fF
C7142 a_2475_14202# a_34090_14178# 0.68fF
C7143 a_21038_8154# col_n[18] 0.34fF
C7144 a_29374_7190# vcm 0.24fF
C7145 a_35002_7150# m2_34864_6970# 0.33fF
C7146 a_20034_16186# vcm 0.89fF
C7147 a_16930_6146# VDD 0.29fF
C7148 a_22042_14178# m2_22240_14426# 0.19fF
C7149 a_2275_1150# col_n[3] 0.17fF
C7150 a_6982_9158# rowon_n[7] 0.45fF
C7151 a_2275_11190# a_25054_11166# 0.71fF
C7152 a_22954_1126# vcm 0.18fF
C7153 a_25054_16186# a_26058_16186# 0.86fF
C7154 a_19030_2130# m2_19228_2378# 0.19fF
C7155 m2_1732_946# VDD 8.31fF
C7156 a_10298_10202# vcm 0.24fF
C7157 a_6982_17190# rowoff_n[15] 2.42fF
C7158 col[8] rowoff_n[14] 0.29fF
C7159 m2_15788_18014# VDD 3.98fF
C7160 a_5886_6146# rowoff_n[4] 0.70fF
C7161 a_23046_5142# ctop 4.91fF
C7162 a_31990_10162# VDD 0.29fF
C7163 a_2275_8178# a_15318_8194# 0.15fF
C7164 a_2475_8178# a_17934_8154# 0.41fF
C7165 a_9902_8154# a_9994_8154# 0.45fF
C7166 a_2475_8178# col[8] 0.22fF
C7167 a_2275_18218# col[30] 0.17fF
C7168 a_14922_4138# rowoff_n[2] 0.60fF
C7169 a_31990_12170# rowoff_n[10] 0.41fF
C7170 a_28066_8154# row_n[6] 0.43fF
C7171 a_25358_14218# vcm 0.24fF
C7172 a_9994_6146# col_n[7] 0.34fF
C7173 m2_34864_6970# m3_34996_7102# 4.42fF
C7174 a_27974_12170# rowon_n[10] 0.14fF
C7175 a_2275_5166# a_8898_5142# 0.17fF
C7176 a_13006_12170# m2_13204_12418# 0.19fF
C7177 a_3970_8154# ctop 4.91fF
C7178 a_2275_14202# col_n[15] 0.17fF
C7179 a_12914_13174# VDD 0.29fF
C7180 a_2275_10186# a_30378_10202# 0.15fF
C7181 a_2475_10186# a_32994_10162# 0.41fF
C7182 a_2275_3158# col_n[20] 0.17fF
C7183 a_23958_2130# rowoff_n[0] 0.50fF
C7184 m2_1732_11990# vcm 1.11fF
C7185 vcm col_n[5] 3.22fF
C7186 VDD col_n[8] 14.45fF
C7187 ctop col[31] 0.40fF
C7188 a_18938_8154# vcm 0.18fF
C7189 a_32082_8154# m2_32280_8402# 0.19fF
C7190 a_2275_11190# col[5] 0.17fF
C7191 a_6282_17230# vcm 0.24fF
C7192 a_4974_16186# rowon_n[14] 0.45fF
C7193 m2_12776_18014# m3_12908_18146# 4.41fF
C7194 a_34394_7190# col_n[31] 0.11fF
C7195 a_2275_7174# a_23958_7150# 0.17fF
C7196 a_30074_5142# col[27] 0.38fF
C7197 a_19030_12170# ctop 4.91fF
C7198 a_27974_17190# VDD 0.29fF
C7199 a_24962_12170# a_25054_12170# 0.45fF
C7200 a_15014_6146# rowon_n[4] 0.45fF
C7201 a_2475_10186# col[25] 0.22fF
C7202 a_1957_16210# a_2161_16210# 0.11fF
C7203 a_2475_16210# a_2275_16210# 2.96fF
C7204 a_33998_12170# vcm 0.18fF
C7205 a_30074_2130# VDD 1.65fF
C7206 a_3878_8154# rowon_n[6] 0.14fF
C7207 a_26058_5142# a_26058_4138# 0.84fF
C7208 a_2475_4162# a_16018_4138# 0.68fF
C7209 a_3970_10162# m2_4168_10410# 0.19fF
C7210 a_25358_5182# col_n[22] 0.11fF
C7211 m3_34996_4090# m3_34996_3086# 0.20fF
C7212 a_8990_16186# col_n[6] 0.34fF
C7213 a_34090_16186# ctop 4.80fF
C7214 a_16018_10162# rowoff_n[8] 1.98fF
C7215 a_26058_15182# row_n[13] 0.43fF
C7216 a_19942_13174# rowoff_n[11] 0.55fF
C7217 m2_34864_1950# a_2475_2154# 0.56fF
C7218 a_3970_1126# a_4274_1166# 0.10fF
C7219 a_2275_1150# a_6982_1126# 0.14fF
C7220 a_23046_6146# m2_23244_6394# 0.19fF
C7221 a_14922_15182# vcm 0.18fF
C7222 a_2275_13198# col[22] 0.17fF
C7223 a_10998_5142# VDD 3.61fF
C7224 a_2475_6170# a_31078_6146# 0.68fF
C7225 a_16018_6146# a_17022_6146# 0.86fF
C7226 a_2275_2154# col[27] 0.17fF
C7227 a_25054_8154# rowoff_n[6] 1.54fF
C7228 a_19030_3134# col[16] 0.38fF
C7229 a_29070_15182# col[26] 0.38fF
C7230 a_2275_15206# a_7286_15222# 0.15fF
C7231 a_2475_15206# a_9902_15182# 0.41fF
C7232 a_5886_15182# a_5978_15182# 0.45fF
C7233 a_34090_6146# rowoff_n[4] 1.10fF
C7234 a_2275_3158# a_22042_3134# 0.71fF
C7235 a_9902_1126# m2_9764_946# 0.31fF
C7236 a_2275_1150# m2_24824_946# 0.51fF
C7237 m3_30980_1078# ctop 0.21fF
C7238 a_26058_9158# VDD 2.06fF
C7239 a_6982_8154# a_6982_7150# 0.84fF
C7240 a_13006_13174# rowon_n[11] 0.45fF
C7241 a_14314_3174# col_n[11] 0.11fF
C7242 a_24354_15222# col_n[21] 0.11fF
C7243 a_32082_4138# vcm 0.89fF
C7244 a_1957_11190# row_n[9] 0.29fF
C7245 a_23046_3134# rowon_n[1] 0.45fF
C7246 a_2275_17214# a_22346_17230# 0.15fF
C7247 a_2475_17214# a_24962_17190# 0.41fF
C7248 a_14010_4138# m2_14208_4386# 0.19fF
C7249 m2_34864_3958# m3_34996_4090# 4.42fF
C7250 col_n[10] rowoff_n[1] 0.27fF
C7251 col_n[13] rowoff_n[4] 0.24fF
C7252 col_n[16] rowoff_n[7] 0.22fF
C7253 col_n[9] rowoff_n[0] 0.27fF
C7254 col_n[17] rowoff_n[8] 0.21fF
C7255 col_n[14] rowoff_n[5] 0.24fF
C7256 col_n[11] rowoff_n[2] 0.26fF
C7257 col_n[18] rowoff_n[9] 0.21fF
C7258 col_n[15] rowoff_n[6] 0.23fF
C7259 col_n[12] rowoff_n[3] 0.25fF
C7260 a_2475_6170# col[2] 0.22fF
C7261 a_2275_18218# a_32386_18234# 0.15fF
C7262 a_6982_12170# VDD 4.02fF
C7263 a_31078_10162# a_32082_10162# 0.86fF
C7264 a_2275_14202# a_15926_14178# 0.17fF
C7265 a_13006_7150# vcm 0.89fF
C7266 a_7894_14178# rowoff_n[12] 0.68fF
C7267 a_18026_13174# col[15] 0.38fF
C7268 a_2275_12194# col_n[9] 0.17fF
C7269 a_34090_12170# row_n[10] 0.43fF
C7270 a_2475_2154# a_29982_2130# 0.41fF
C7271 a_2275_2154# a_27366_2170# 0.15fF
C7272 a_15926_2130# a_16018_2130# 0.45fF
C7273 a_1957_16210# vcm 0.16fF
C7274 a_2275_1150# col_n[14] 0.17fF
C7275 a_33998_16186# rowon_n[14] 0.14fF
C7276 a_33086_9158# col_n[30] 0.34fF
C7277 a_22042_16186# VDD 2.47fF
C7278 a_22042_12170# a_22042_11166# 0.84fF
C7279 a_2475_11190# a_7986_11166# 0.68fF
C7280 a_3270_1166# vcm 0.25fF
C7281 col[19] rowoff_n[14] 0.22fF
C7282 a_2275_16210# a_30986_16186# 0.17fF
C7283 a_13310_13214# col_n[10] 0.11fF
C7284 a_28066_11166# vcm 0.89fF
C7285 col_n[2] rowoff_n[10] 0.32fF
C7286 a_24962_1126# VDD 0.76fF
C7287 a_2475_8178# col[19] 0.22fF
C7288 a_21038_10162# rowon_n[8] 0.45fF
C7289 a_12002_13174# a_13006_13174# 0.86fF
C7290 a_2475_13198# a_23046_13174# 0.68fF
C7291 a_18330_5182# vcm 0.24fF
C7292 a_2275_14202# col_n[26] 0.17fF
C7293 a_8990_14178# vcm 0.89fF
C7294 a_5886_4138# VDD 0.29fF
C7295 a_2275_3158# col_n[31] 0.17fF
C7296 a_6982_11166# col[4] 0.38fF
C7297 a_30986_6146# a_31078_6146# 0.45fF
C7298 a_2275_10186# a_14010_10162# 0.71fF
C7299 vcm col_n[16] 3.19fF
C7300 VDD col_n[19] 11.72fF
C7301 col[3] rowoff_n[15] 0.33fF
C7302 a_22042_7150# col_n[19] 0.34fF
C7303 a_2275_11190# col[16] 0.17fF
C7304 a_33390_9198# vcm 0.24fF
C7305 a_8898_4138# rowon_n[2] 0.14fF
C7306 a_24050_18194# vcm 0.15fF
C7307 a_12002_3134# ctop 4.91fF
C7308 m2_6752_18014# col_n[4] 0.32fF
C7309 a_20946_8154# VDD 0.29fF
C7310 a_2275_7174# a_4274_7190# 0.15fF
C7311 a_2475_7174# a_6890_7150# 0.41fF
C7312 a_2275_12194# a_29070_12170# 0.71fF
C7313 a_26970_3134# vcm 0.18fF
C7314 a_27062_17190# a_28066_17190# 0.86fF
C7315 a_2275_3158# m2_1732_2954# 0.27fF
C7316 a_6890_5142# rowoff_n[3] 0.69fF
C7317 a_14314_12210# vcm 0.24fF
C7318 a_27062_7150# ctop 4.91fF
C7319 m3_27968_18146# m3_28972_18146# 0.21fF
C7320 a_11910_9158# a_12002_9158# 0.45fF
C7321 a_19030_17190# rowon_n[15] 0.45fF
C7322 a_2275_9182# a_19334_9198# 0.15fF
C7323 a_2475_9182# a_21950_9158# 0.41fF
C7324 a_15926_3134# rowoff_n[1] 0.59fF
C7325 a_7894_6146# vcm 0.18fF
C7326 a_29070_7150# rowon_n[5] 0.45fF
C7327 a_10998_5142# col_n[8] 0.34fF
C7328 a_21038_17190# col_n[18] 0.34fF
C7329 a_29374_16226# vcm 0.24fF
C7330 a_2275_6170# a_12914_6146# 0.17fF
C7331 a_7986_10162# ctop 4.91fF
C7332 a_16930_15182# VDD 0.29fF
C7333 a_2275_11190# a_35398_11206# 0.15fF
C7334 a_2275_10186# col_n[3] 0.17fF
C7335 a_6982_7150# row_n[5] 0.43fF
C7336 a_6890_11166# rowon_n[9] 0.14fF
C7337 a_22954_10162# vcm 0.18fF
C7338 a_2475_3158# a_4974_3134# 0.68fF
C7339 a_31078_4138# col[28] 0.38fF
C7340 a_21038_2130# m2_20808_946# 0.84fF
C7341 m3_26964_18146# ctop 0.21fF
C7342 a_2275_8178# a_27974_8154# 0.17fF
C7343 a_23046_14178# ctop 4.91fF
C7344 a_26970_13174# a_27062_13174# 0.45fF
C7345 a_7986_11166# rowoff_n[9] 2.38fF
C7346 a_2275_17214# a_5978_17190# 0.71fF
C7347 a_2475_17214# col[8] 0.22fF
C7348 col_n[25] rowoff_n[5] 0.16fF
C7349 col_n[28] rowoff_n[8] 0.14fF
C7350 col_n[21] rowoff_n[1] 0.19fF
C7351 col_n[24] rowoff_n[4] 0.16fF
C7352 col_n[22] rowoff_n[2] 0.18fF
C7353 col_n[29] rowoff_n[9] 0.13fF
C7354 col_n[26] rowoff_n[6] 0.15fF
C7355 col_n[23] rowoff_n[3] 0.17fF
C7356 col_n[20] rowoff_n[0] 0.19fF
C7357 col_n[27] rowoff_n[7] 0.14fF
C7358 a_34090_5142# m2_34864_4962# 0.86fF
C7359 a_2475_6170# col[13] 0.22fF
C7360 a_26362_4178# col_n[23] 0.11fF
C7361 a_34090_4138# VDD 1.23fF
C7362 a_28066_6146# a_28066_5142# 0.84fF
C7363 a_2475_5166# a_20034_5142# 0.68fF
C7364 a_9994_15182# col_n[7] 0.34fF
C7365 a_2275_18218# a_16018_18194# 0.14fF
C7366 a_3970_17190# ctop 4.93fF
C7367 a_17022_9158# rowoff_n[7] 1.94fF
C7368 a_27062_14178# rowon_n[12] 0.45fF
C7369 a_2275_12194# col_n[20] 0.17fF
C7370 a_2275_1150# col_n[25] 0.17fF
C7371 a_24050_15182# rowoff_n[13] 1.59fF
C7372 a_2275_2154# a_10998_2130# 0.71fF
C7373 a_18938_17190# vcm 0.18fF
C7374 a_15014_7150# VDD 3.20fF
C7375 a_26058_7150# rowoff_n[5] 1.50fF
C7376 a_18026_7150# a_19030_7150# 0.86fF
C7377 a_28066_15182# m2_28264_15430# 0.19fF
C7378 a_20034_2130# col[17] 0.38fF
C7379 a_2275_9182# col[10] 0.17fF
C7380 a_34394_16226# col_n[31] 0.11fF
C7381 col[30] rowoff_n[14] 0.15fF
C7382 a_4974_14178# row_n[12] 0.43fF
C7383 a_30074_14178# col[27] 0.38fF
C7384 a_21038_2130# vcm 0.89fF
C7385 col_n[13] rowoff_n[10] 0.24fF
C7386 a_2275_16210# a_11302_16226# 0.15fF
C7387 a_2475_16210# a_13918_16186# 0.41fF
C7388 a_7894_16186# a_7986_16186# 0.45fF
C7389 a_15014_4138# row_n[2] 0.43fF
C7390 a_2475_8178# col[30] 0.22fF
C7391 a_14922_8154# rowon_n[6] 0.14fF
C7392 a_2275_4162# a_26058_4138# 0.71fF
C7393 a_30074_11166# VDD 1.65fF
C7394 m3_34996_2082# m3_34996_1078# 0.20fF
C7395 a_15318_2170# col_n[12] 0.11fF
C7396 a_8990_9158# a_8990_8154# 0.84fF
C7397 a_25358_14218# col_n[22] 0.11fF
C7398 a_2275_13198# a_4882_13174# 0.17fF
C7399 a_2966_13174# a_3970_13174# 0.86fF
C7400 a_2966_10162# rowon_n[8] 0.45fF
C7401 a_2475_5166# vcm 1.32fF
C7402 a_2475_1150# a_18938_1126# 0.44fF
C7403 a_2275_1150# a_16322_1166# 0.15fF
C7404 a_19030_13174# m2_19228_13422# 0.19fF
C7405 VDD col_n[30] 8.98fF
C7406 vcm col_n[27] 3.22fF
C7407 col[14] rowoff_n[15] 0.25fF
C7408 a_10998_14178# VDD 3.61fF
C7409 a_33086_11166# a_34090_11166# 0.86fF
C7410 a_2275_11190# col[27] 0.17fF
C7411 a_2475_2154# rowon_n[0] 0.40fF
C7412 VDD rowoff_n[11] 87.22fF
C7413 a_2275_15206# a_19942_15182# 0.17fF
C7414 a_19030_12170# col[16] 0.38fF
C7415 a_17022_9158# vcm 0.89fF
C7416 a_12002_16186# rowoff_n[14] 2.18fF
C7417 a_2275_3158# a_31382_3174# 0.15fF
C7418 a_2475_3158# a_33998_3134# 0.41fF
C7419 a_17934_3134# a_18026_3134# 0.45fF
C7420 a_2275_8178# VDD 3.18fF
C7421 a_34090_8154# col_n[31] 0.34fF
C7422 a_24050_13174# a_24050_12170# 0.84fF
C7423 a_2475_12194# a_12002_12170# 0.68fF
C7424 a_14314_12210# col_n[11] 0.11fF
C7425 a_7286_3174# vcm 0.24fF
C7426 a_13006_11166# row_n[9] 0.43fF
C7427 a_2275_17214# a_35002_17190# 0.17fF
C7428 a_12914_15182# rowon_n[13] 0.14fF
C7429 a_32082_13174# vcm 0.89fF
C7430 m2_9764_946# col_n[7] 0.45fF
C7431 a_28978_3134# VDD 0.29fF
C7432 a_9994_11166# m2_10192_11414# 0.19fF
C7433 a_22954_5142# rowon_n[3] 0.14fF
C7434 m2_30848_946# m2_31852_946# 0.86fF
C7435 a_2275_9182# a_2874_9158# 0.17fF
C7436 a_2475_9182# a_3878_9158# 0.41fF
C7437 a_2475_15206# col[2] 0.22fF
C7438 a_2475_18218# m2_7756_18014# 0.62fF
C7439 a_2475_4162# col[7] 0.22fF
C7440 a_14010_14178# a_15014_14178# 0.86fF
C7441 a_2475_14202# a_27062_14178# 0.68fF
C7442 a_22346_7190# vcm 0.24fF
C7443 a_29070_7150# m2_29268_7398# 0.19fF
C7444 a_7986_10162# col[5] 0.38fF
C7445 a_13006_16186# vcm 0.89fF
C7446 a_9902_6146# VDD 0.29fF
C7447 a_32994_7150# a_33086_7150# 0.45fF
C7448 a_2275_10186# col_n[14] 0.17fF
C7449 a_2275_11190# a_18026_11166# 0.71fF
C7450 a_23046_6146# col_n[20] 0.34fF
C7451 a_15926_1126# vcm 0.18fF
C7452 a_4974_16186# a_4974_15182# 0.84fF
C7453 a_3270_10202# vcm 0.24fF
C7454 m2_1732_18014# VDD 5.99fF
C7455 a_2275_7174# col[4] 0.17fF
C7456 a_16018_5142# ctop 4.91fF
C7457 a_24962_10162# VDD 0.29fF
C7458 a_2275_8178# a_8290_8194# 0.15fF
C7459 a_2475_8178# a_10906_8154# 0.41fF
C7460 a_2475_17214# col[19] 0.22fF
C7461 a_2275_13198# a_33086_13174# 0.71fF
C7462 col_n[31] rowoff_n[0] 0.11fF
C7463 a_2475_6170# col[24] 0.22fF
C7464 a_30986_5142# vcm 0.18fF
C7465 a_7894_4138# rowoff_n[2] 0.68fF
C7466 a_24962_12170# rowoff_n[10] 0.49fF
C7467 a_21038_8154# row_n[6] 0.43fF
C7468 a_20034_5142# m2_20232_5390# 0.19fF
C7469 a_18330_14218# vcm 0.24fF
C7470 a_20946_12170# rowon_n[10] 0.14fF
C7471 a_31078_9158# ctop 4.91fF
C7472 a_5886_13174# VDD 0.29fF
C7473 a_2275_12194# col_n[31] 0.17fF
C7474 a_13918_10162# a_14010_10162# 0.45fF
C7475 a_2275_10186# a_23350_10202# 0.15fF
C7476 a_2475_10186# a_25966_10162# 0.41fF
C7477 a_30986_2130# rowon_n[0] 0.14fF
C7478 a_16930_2130# rowoff_n[0] 0.58fF
C7479 a_12002_4138# col_n[9] 0.34fF
C7480 a_22042_16186# col_n[19] 0.34fF
C7481 a_11910_8154# vcm 0.18fF
C7482 a_15014_3134# a_15014_2130# 0.84fF
C7483 a_33390_18234# vcm 0.25fF
C7484 a_2275_9182# col[21] 0.17fF
C7485 a_2275_7174# a_16930_7150# 0.17fF
C7486 a_12002_12170# ctop 4.91fF
C7487 a_20946_17190# VDD 0.29fF
C7488 col_n[24] rowoff_n[10] 0.16fF
C7489 a_7986_6146# rowon_n[4] 0.45fF
C7490 a_2966_2130# vcm 0.15fF
C7491 a_10998_3134# m2_11196_3382# 0.19fF
C7492 a_26970_12170# vcm 0.18fF
C7493 a_23046_2130# VDD 2.37fF
C7494 a_32082_3134# col[29] 0.38fF
C7495 a_2475_4162# a_8990_4138# 0.68fF
C7496 a_4974_4138# a_5978_4138# 0.86fF
C7497 m2_21812_18014# col[19] 0.39fF
C7498 m3_34996_11118# m3_34996_10114# 0.20fF
C7499 m2_33860_946# m3_34568_1078# 1.25fF
C7500 a_2275_9182# a_31990_9158# 0.17fF
C7501 a_22954_18194# m2_22816_18014# 0.34fF
C7502 a_27062_16186# ctop 4.91fF
C7503 a_28978_14178# a_29070_14178# 0.45fF
C7504 a_8990_10162# rowoff_n[8] 2.33fF
C7505 a_19030_15182# row_n[13] 0.43fF
C7506 a_12914_13174# rowoff_n[11] 0.63fF
C7507 a_27366_3174# col_n[24] 0.11fF
C7508 col_n[1] row_n[13] 0.37fF
C7509 col_n[6] rowon_n[15] 0.17fF
C7510 col_n[4] rowon_n[14] 0.17fF
C7511 col_n[2] rowon_n[13] 0.17fF
C7512 sample rowon_n[11] 0.10fF
C7513 col_n[3] row_n[14] 0.37fF
C7514 vcm rowon_n[12] 0.91fF
C7515 col_n[5] row_n[15] 0.37fF
C7516 VDD row_n[11] 4.64fF
C7517 col_n[0] row_n[12] 0.37fF
C7518 col[25] rowoff_n[15] 0.18fF
C7519 a_7894_15182# vcm 0.18fF
C7520 a_10998_14178# col_n[8] 0.34fF
C7521 a_3970_5142# VDD 4.33fF
C7522 a_29070_5142# row_n[3] 0.43fF
C7523 a_30074_7150# a_30074_6146# 0.84fF
C7524 a_2475_6170# a_24050_6146# 0.68fF
C7525 a_2475_2154# col[1] 0.22fF
C7526 a_28978_9158# rowon_n[7] 0.14fF
C7527 col_n[8] rowoff_n[11] 0.28fF
C7528 a_18026_8154# rowoff_n[6] 1.89fF
C7529 a_2275_8178# col_n[8] 0.17fF
C7530 a_28978_17190# rowoff_n[15] 0.44fF
C7531 a_2275_3158# a_15014_3134# 0.71fF
C7532 a_27062_6146# rowoff_n[4] 1.45fF
C7533 a_2475_1150# m2_10768_946# 0.62fF
C7534 a_19030_9158# VDD 2.78fF
C7535 a_20034_8154# a_21038_8154# 0.86fF
C7536 a_5978_13174# rowon_n[11] 0.45fF
C7537 a_31078_13174# col[28] 0.38fF
C7538 a_25054_4138# vcm 0.89fF
C7539 a_16018_3134# rowon_n[1] 0.45fF
C7540 a_2475_17214# a_17934_17190# 0.41fF
C7541 a_2275_17214# a_15318_17230# 0.15fF
C7542 a_9902_17190# a_9994_17190# 0.45fF
C7543 a_16322_1166# col_n[13] 0.11fF
C7544 a_2275_5166# a_30074_5142# 0.71fF
C7545 a_2475_15206# col[13] 0.22fF
C7546 a_26362_13214# col_n[23] 0.11fF
C7547 a_34090_13174# VDD 1.23fF
C7548 a_2275_18218# a_25358_18234# 0.15fF
C7549 a_2475_4162# col[18] 0.22fF
C7550 m2_11772_946# m2_12200_1374# 0.19fF
C7551 a_10998_10162# a_10998_9158# 0.84fF
C7552 a_2275_14202# a_8898_14178# 0.17fF
C7553 a_5978_7150# vcm 0.89fF
C7554 a_27062_12170# row_n[10] 0.43fF
C7555 a_2275_2154# a_20338_2170# 0.15fF
C7556 a_2475_2154# a_22954_2130# 0.41fF
C7557 a_2275_10186# col_n[25] 0.17fF
C7558 a_26970_16186# rowon_n[14] 0.14fF
C7559 a_15014_16186# VDD 3.20fF
C7560 a_20034_11166# col[17] 0.38fF
C7561 a_30378_2170# vcm 0.24fF
C7562 a_2275_16210# a_23958_16186# 0.17fF
C7563 a_2275_7174# col[15] 0.17fF
C7564 a_21038_11166# vcm 0.89fF
C7565 a_17934_1126# VDD 0.73fF
C7566 a_19942_4138# a_20034_4138# 0.45fF
C7567 m2_34864_9982# row_n[8] 0.38fF
C7568 a_2475_17214# col[30] 0.22fF
C7569 row_n[7] rowoff_n[7] 0.64fF
C7570 a_19030_17190# m2_18800_18014# 0.84fF
C7571 a_2475_17214# m2_34864_17010# 0.56fF
C7572 a_15318_11206# col_n[12] 0.11fF
C7573 a_2475_13198# a_16018_13174# 0.68fF
C7574 a_26058_14178# a_26058_13174# 0.84fF
C7575 a_14010_10162# rowon_n[8] 0.45fF
C7576 a_11302_5182# vcm 0.24fF
C7577 m2_4744_946# vcm 0.71fF
C7578 a_2874_18194# m2_2736_18014# 0.34fF
C7579 a_2966_8154# row_n[6] 0.41fF
C7580 a_2275_1150# a_28978_1126# 0.17fF
C7581 a_2475_14202# vcm 1.32fF
C7582 a_32994_5142# VDD 0.29fF
C7583 a_2275_12194# rowon_n[10] 1.99fF
C7584 a_2275_10186# a_6982_10162# 0.71fF
C7585 a_2475_15206# a_31078_15182# 0.68fF
C7586 a_16018_15182# a_17022_15182# 0.86fF
C7587 a_8990_9158# col[6] 0.38fF
C7588 a_26362_9198# vcm 0.24fF
C7589 a_4974_3134# ctop 4.91fF
C7590 a_17022_18194# vcm 0.15fF
C7591 a_13918_8154# VDD 0.29fF
C7592 a_35002_8154# a_35094_8154# 0.11fF
C7593 a_34090_16186# m2_34288_16434# 0.19fF
C7594 a_24050_5142# col_n[21] 0.34fF
C7595 a_35002_13174# rowon_n[11] 0.14fF
C7596 a_2275_17214# VDD 3.18fF
C7597 a_34090_17190# col_n[31] 0.34fF
C7598 a_2275_12194# a_22042_12170# 0.71fF
C7599 a_2275_6170# col_n[2] 0.17fF
C7600 a_19942_3134# vcm 0.18fF
C7601 a_4274_9198# col_n[1] 0.11fF
C7602 a_6982_17190# a_6982_16186# 0.84fF
C7603 m2_1732_15002# sample 0.31fF
C7604 a_7286_12210# vcm 0.24fF
C7605 a_20034_7150# ctop 4.91fF
C7606 a_28978_12170# VDD 0.29fF
C7607 m3_13912_18146# m3_14916_18146# 0.21fF
C7608 a_12002_17190# rowon_n[15] 0.45fF
C7609 a_2275_9182# a_12306_9198# 0.15fF
C7610 a_2475_9182# a_14922_9158# 0.41fF
C7611 a_8898_3134# rowoff_n[1] 0.67fF
C7612 col_n[7] rowon_n[10] 0.17fF
C7613 col_n[5] rowon_n[9] 0.17fF
C7614 col_n[3] rowon_n[8] 0.17fF
C7615 col_n[10] row_n[12] 0.37fF
C7616 col_n[9] rowon_n[11] 0.17fF
C7617 col_n[17] rowon_n[15] 0.17fF
C7618 vcm row_n[7] 1.08fF
C7619 col_n[6] row_n[10] 0.37fF
C7620 col_n[11] rowon_n[12] 0.17fF
C7621 col_n[12] row_n[13] 0.37fF
C7622 col_n[0] rowon_n[6] 0.17fF
C7623 col_n[14] row_n[14] 0.37fF
C7624 col_n[1] rowon_n[7] 0.17fF
C7625 col_n[16] row_n[15] 0.37fF
C7626 col_n[8] row_n[11] 0.37fF
C7627 col_n[2] row_n[8] 0.37fF
C7628 col_n[13] rowon_n[13] 0.17fF
C7629 VDD rowon_n[5] 4.61fF
C7630 col_n[4] row_n[9] 0.37fF
C7631 sample row_n[6] 0.92fF
C7632 col_n[15] rowon_n[14] 0.17fF
C7633 m2_34864_6970# m2_35292_7398# 0.19fF
C7634 a_22042_7150# rowon_n[5] 0.45fF
C7635 a_35002_7150# vcm 0.18fF
C7636 a_29070_14178# rowoff_n[12] 1.35fF
C7637 a_2475_13198# col[7] 0.22fF
C7638 a_26058_2130# a_27062_2130# 0.86fF
C7639 a_2475_2154# col[12] 0.22fF
C7640 a_2966_6146# m2_3164_6394# 0.19fF
C7641 col_n[19] rowoff_n[11] 0.20fF
C7642 a_22346_16226# vcm 0.24fF
C7643 a_25054_14178# m2_25252_14426# 0.19fF
C7644 a_2275_6170# a_5886_6146# 0.17fF
C7645 a_9902_15182# VDD 0.29fF
C7646 a_15926_11166# a_16018_11166# 0.45fF
C7647 a_2475_11190# a_29982_11166# 0.41fF
C7648 a_2275_11190# a_27366_11206# 0.15fF
C7649 a_13006_3134# col_n[10] 0.34fF
C7650 a_2275_8178# col_n[19] 0.17fF
C7651 a_23046_15182# col_n[20] 0.34fF
C7652 a_15926_10162# vcm 0.18fF
C7653 a_33086_16186# row_n[14] 0.43fF
C7654 a_17022_4138# a_17022_3134# 0.84fF
C7655 a_35494_10524# VDD 0.13fF
C7656 a_2275_16210# col[4] 0.17fF
C7657 a_2275_8178# a_20946_8154# 0.17fF
C7658 a_16018_14178# ctop 4.91fF
C7659 a_2275_5166# col[9] 0.17fF
C7660 a_33086_2130# col[30] 0.38fF
C7661 col_n[3] rowoff_n[12] 0.32fF
C7662 a_2475_15206# col[24] 0.22fF
C7663 a_30986_14178# vcm 0.18fF
C7664 a_27062_4138# VDD 1.96fF
C7665 a_2475_4162# col[29] 0.22fF
C7666 a_6982_5142# a_7986_5142# 0.86fF
C7667 a_16018_12170# m2_16216_12418# 0.19fF
C7668 a_2475_5166# a_13006_5142# 0.68fF
C7669 a_2275_18218# a_8990_18194# 0.14fF
C7670 a_2275_10186# a_34394_10202# 0.15fF
C7671 a_9994_9158# rowoff_n[7] 2.28fF
C7672 a_20034_14178# rowon_n[12] 0.45fF
C7673 a_30986_15182# a_31078_15182# 0.45fF
C7674 a_28370_2170# col_n[25] 0.11fF
C7675 a_17022_15182# rowoff_n[13] 1.94fF
C7676 a_12002_13174# col_n[9] 0.34fF
C7677 a_2275_2154# a_3970_2130# 0.71fF
C7678 a_30074_4138# rowon_n[2] 0.45fF
C7679 a_11910_17190# vcm 0.18fF
C7680 m2_17796_18014# m3_17928_18146# 4.41fF
C7681 a_7986_7150# VDD 3.92fF
C7682 a_19030_7150# rowoff_n[5] 1.84fF
C7683 a_32082_8154# a_32082_7150# 0.84fF
C7684 a_2475_7174# a_28066_7150# 0.68fF
C7685 a_2275_7174# col[26] 0.17fF
C7686 a_14010_2130# vcm 0.89fF
C7687 a_2475_16210# a_6890_16186# 0.41fF
C7688 a_2275_16210# a_4274_16226# 0.15fF
C7689 a_28066_5142# rowoff_n[3] 1.40fF
C7690 a_2966_11166# vcm 0.89fF
C7691 a_7986_4138# row_n[2] 0.43fF
C7692 rowon_n[3] rowoff_n[3] 20.66fF
C7693 a_7894_8154# rowon_n[6] 0.14fF
C7694 a_6982_10162# m2_7180_10410# 0.19fF
C7695 a_2275_4162# a_19030_4138# 0.71fF
C7696 a_23046_11166# VDD 2.37fF
C7697 a_32082_12170# col[29] 0.38fF
C7698 m3_3872_1078# m3_4876_1078# 0.21fF
C7699 a_22042_9158# a_23046_9158# 0.86fF
C7700 a_29070_6146# vcm 0.89fF
C7701 a_11910_18194# a_12002_18194# 0.11fF
C7702 a_2475_1150# a_11910_1126# 0.41fF
C7703 a_26058_6146# m2_26256_6394# 0.19fF
C7704 a_2275_1150# a_9294_1166# 0.15fF
C7705 a_6890_1126# a_6982_1126# 0.11fF
C7706 a_27366_12210# col_n[24] 0.11fF
C7707 m2_8760_946# VDD 6.40fF
C7708 a_2275_6170# a_34090_6146# 0.71fF
C7709 a_3970_14178# VDD 4.33fF
C7710 a_13006_11166# a_13006_10162# 0.84fF
C7711 a_2475_11190# col[1] 0.22fF
C7712 a_2275_15206# a_12914_15182# 0.17fF
C7713 a_28066_11166# rowon_n[9] 0.45fF
C7714 a_9994_9158# vcm 0.89fF
C7715 a_4974_16186# rowoff_n[14] 2.52fF
C7716 a_2275_3158# a_24354_3174# 0.15fF
C7717 a_2475_3158# a_26970_3134# 0.41fF
C7718 a_2475_1150# m2_33860_946# 0.42fF
C7719 a_2275_17214# col_n[8] 0.17fF
C7720 a_2275_6170# col_n[13] 0.17fF
C7721 a_21038_10162# col[18] 0.38fF
C7722 a_2475_12194# a_4974_12170# 0.68fF
C7723 a_5978_11166# row_n[9] 0.43fF
C7724 a_35398_4178# vcm 0.24fF
C7725 a_29982_11166# rowoff_n[9] 0.43fF
C7726 a_2275_17214# a_27974_17190# 0.17fF
C7727 a_5886_15182# rowon_n[13] 0.14fF
C7728 a_3270_6186# col_n[0] 0.11fF
C7729 a_17022_4138# m2_17220_4386# 0.19fF
C7730 a_25054_13174# vcm 0.89fF
C7731 a_2275_3158# col[3] 0.17fF
C7732 a_21950_3134# VDD 0.29fF
C7733 a_21950_5142# a_22042_5142# 0.45fF
C7734 a_15926_5142# rowon_n[3] 0.14fF
C7735 m2_23820_946# m2_24824_946# 0.86fF
C7736 a_16322_10202# col_n[13] 0.11fF
C7737 col_n[25] row_n[14] 0.37fF
C7738 col_n[7] row_n[5] 0.37fF
C7739 col_n[23] row_n[13] 0.37fF
C7740 col_n[5] row_n[4] 0.37fF
C7741 col_n[3] row_n[3] 0.37fF
C7742 col_n[22] rowon_n[12] 0.17fF
C7743 col_n[18] rowon_n[10] 0.17fF
C7744 col_n[16] rowon_n[9] 0.17fF
C7745 col_n[11] row_n[7] 0.37fF
C7746 col_n[2] rowon_n[2] 0.17fF
C7747 col_n[27] row_n[15] 0.37fF
C7748 col_n[9] row_n[6] 0.37fF
C7749 col_n[4] rowon_n[3] 0.17fF
C7750 col_n[19] row_n[11] 0.37fF
C7751 sample rowon_n[0] 0.10fF
C7752 col_n[13] row_n[8] 0.37fF
C7753 col_n[6] rowon_n[4] 0.17fF
C7754 vcm rowon_n[1] 0.91fF
C7755 col_n[24] rowon_n[13] 0.17fF
C7756 col_n[15] row_n[9] 0.37fF
C7757 col_n[8] rowon_n[5] 0.17fF
C7758 col_n[26] rowon_n[14] 0.17fF
C7759 col_n[0] row_n[1] 0.37fF
C7760 col_n[1] row_n[2] 0.37fF
C7761 col_n[17] row_n[10] 0.37fF
C7762 col_n[10] rowon_n[6] 0.17fF
C7763 col_n[28] rowon_n[15] 0.17fF
C7764 col_n[12] rowon_n[7] 0.17fF
C7765 col_n[20] rowon_n[11] 0.17fF
C7766 col_n[21] row_n[12] 0.37fF
C7767 col_n[14] rowon_n[8] 0.17fF
C7768 VDD row_n[0] 4.64fF
C7769 a_2475_13198# col[18] 0.22fF
C7770 a_28066_15182# a_28066_14178# 0.84fF
C7771 a_2475_14202# a_20034_14178# 0.68fF
C7772 a_2475_2154# col[23] 0.22fF
C7773 col_n[30] rowoff_n[11] 0.12fF
C7774 a_15318_7190# vcm 0.24fF
C7775 a_2275_2154# a_32994_2130# 0.17fF
C7776 a_28066_2130# ctop 4.93fF
C7777 a_5978_16186# vcm 0.89fF
C7778 a_2161_6170# VDD 0.23fF
C7779 a_2275_8178# col_n[30] 0.17fF
C7780 a_2275_11190# a_10998_11166# 0.71fF
C7781 a_8898_1126# vcm 0.18fF
C7782 a_18026_16186# a_19030_16186# 0.86fF
C7783 a_9994_8154# col[7] 0.38fF
C7784 a_30378_11206# vcm 0.24fF
C7785 a_28466_1488# VDD 0.13fF
C7786 a_2275_16210# col[15] 0.17fF
C7787 a_2275_5166# col[20] 0.17fF
C7788 a_8990_5142# ctop 4.91fF
C7789 a_25054_4138# col_n[22] 0.34fF
C7790 a_17934_10162# VDD 0.29fF
C7791 a_2275_13198# a_26058_13174# 0.71fF
C7792 col_n[14] rowoff_n[12] 0.24fF
C7793 a_5278_8194# col_n[2] 0.11fF
C7794 a_23958_5142# vcm 0.18fF
C7795 a_17934_12170# rowoff_n[10] 0.57fF
C7796 m2_27836_946# vcm 0.71fF
C7797 a_2275_18218# m2_24824_18014# 0.51fF
C7798 a_14010_8154# row_n[6] 0.43fF
C7799 a_11302_14218# vcm 0.24fF
C7800 a_13918_12170# rowon_n[10] 0.14fF
C7801 a_2475_12194# m2_1732_11990# 0.16fF
C7802 a_24050_9158# ctop 4.91fF
C7803 a_32994_14178# VDD 0.29fF
C7804 a_2475_10186# a_18938_10162# 0.41fF
C7805 a_2275_10186# a_16322_10202# 0.15fF
C7806 a_2275_10186# row_n[8] 26.41fF
C7807 a_23958_2130# rowon_n[0] 0.14fF
C7808 a_9902_2130# rowoff_n[0] 0.66fF
C7809 a_4882_8154# vcm 0.18fF
C7810 a_33998_16186# rowoff_n[14] 0.39fF
C7811 a_28066_3134# a_29070_3134# 0.86fF
C7812 a_26362_18234# vcm 0.25fF
C7813 a_31990_1126# m2_31852_946# 0.31fF
C7814 a_2275_7174# a_9902_7150# 0.17fF
C7815 a_4974_12170# ctop 4.91fF
C7816 a_14010_2130# col_n[11] 0.34fF
C7817 a_13918_17190# VDD 0.29fF
C7818 sample rowoff_n[13] 0.22fF
C7819 a_2475_12194# a_33998_12170# 0.41fF
C7820 a_2275_12194# a_31382_12210# 0.15fF
C7821 a_17934_12170# a_18026_12170# 0.45fF
C7822 a_24050_14178# col_n[21] 0.34fF
C7823 col[0] rowoff_n[8] 0.34fF
C7824 col[1] rowoff_n[9] 0.34fF
C7825 a_2275_15206# col_n[2] 0.17fF
C7826 ctop rowoff_n[2] 0.28fF
C7827 a_34090_15182# rowon_n[13] 0.45fF
C7828 a_2275_4162# col_n[7] 0.17fF
C7829 a_19942_12170# vcm 0.18fF
C7830 a_4274_18234# col_n[1] 0.11fF
C7831 a_16018_2130# VDD 3.09fF
C7832 a_1957_8178# sample 0.35fF
C7833 a_19030_5142# a_19030_4138# 0.84fF
C7834 m3_34996_18146# m3_34996_17142# 0.20fF
C7835 m2_24824_946# m3_24956_1078# 4.41fF
C7836 a_2275_9182# a_24962_9158# 0.17fF
C7837 a_20034_16186# ctop 4.91fF
C7838 a_2475_10186# rowoff_n[8] 4.75fF
C7839 a_12002_15182# row_n[13] 0.43fF
C7840 a_5886_13174# rowoff_n[11] 0.70fF
C7841 m2_34864_3958# VDD 1.59fF
C7842 a_35002_16186# vcm 0.18fF
C7843 a_31078_6146# VDD 1.54fF
C7844 a_22042_5142# row_n[3] 0.43fF
C7845 a_8990_6146# a_9994_6146# 0.86fF
C7846 a_2475_6170# a_17022_6146# 0.68fF
C7847 a_2475_11190# col[12] 0.22fF
C7848 a_21950_9158# rowon_n[7] 0.14fF
C7849 a_10998_8154# rowoff_n[6] 2.23fF
C7850 a_29374_1166# col_n[26] 0.11fF
C7851 a_32994_16186# a_33086_16186# 0.45fF
C7852 m2_34864_11990# rowon_n[10] 0.42fF
C7853 a_13006_12170# col_n[10] 0.34fF
C7854 a_2275_17214# col_n[19] 0.17fF
C7855 a_21950_17190# rowoff_n[15] 0.52fF
C7856 a_2275_6170# col_n[24] 0.17fF
C7857 a_2275_3158# a_7986_3134# 0.71fF
C7858 a_20034_6146# rowoff_n[4] 1.79fF
C7859 a_2275_18218# col_n[4] 0.17fF
C7860 m3_1864_14130# ctop 0.22fF
C7861 a_12002_9158# VDD 3.51fF
C7862 a_2475_8178# a_32082_8154# 0.68fF
C7863 a_34090_9158# a_34090_8154# 0.84fF
C7864 a_2275_14202# col[9] 0.17fF
C7865 a_18026_4138# vcm 0.89fF
C7866 a_2475_17214# a_10906_17190# 0.41fF
C7867 a_2275_17214# a_8290_17230# 0.15fF
C7868 a_8990_3134# rowon_n[1] 0.45fF
C7869 a_29070_4138# rowoff_n[2] 1.35fF
C7870 a_2275_3158# col[14] 0.17fF
C7871 a_2966_4138# m2_1732_3958# 0.86fF
C7872 a_3878_3134# VDD 0.29fF
C7873 a_33086_11166# col[30] 0.38fF
C7874 col_n[17] rowon_n[4] 0.17fF
C7875 col_n[24] row_n[8] 0.37fF
C7876 col_n[30] row_n[11] 0.37fF
C7877 col_n[15] rowon_n[3] 0.17fF
C7878 col_n[22] row_n[7] 0.37fF
C7879 col_n[13] rowon_n[2] 0.17fF
C7880 col_n[20] row_n[6] 0.37fF
C7881 col_n[11] rowon_n[1] 0.17fF
C7882 col_n[18] row_n[5] 0.37fF
C7883 col_n[9] rowon_n[0] 0.17fF
C7884 col_n[16] row_n[4] 0.37fF
C7885 col_n[0] col[0] 0.50fF
C7886 a_2275_5166# a_23046_5142# 0.71fF
C7887 col_n[14] row_n[3] 0.37fF
C7888 col_n[21] rowon_n[6] 0.17fF
C7889 col_n[28] row_n[10] 0.37fF
C7890 vcm analog_in 0.13fF
C7891 col_n[19] rowon_n[5] 0.17fF
C7892 col_n[26] row_n[9] 0.37fF
C7893 col_n[23] rowon_n[7] 0.17fF
C7894 col_n[31] rowon_n[11] 0.17fF
C7895 col_n[25] rowon_n[8] 0.17fF
C7896 col_n[27] rowon_n[9] 0.17fF
C7897 VDD col[2] 12.90fF
C7898 col_n[8] row_n[0] 0.37fF
C7899 col_n[29] rowon_n[10] 0.17fF
C7900 col_n[10] row_n[1] 0.37fF
C7901 col_n[12] row_n[2] 0.37fF
C7902 a_27062_13174# VDD 1.96fF
C7903 a_2475_13198# col[29] 0.22fF
C7904 a_2275_18218# a_18330_18234# 0.15fF
C7905 m2_4744_946# m2_5172_1374# 0.19fF
C7906 a_24050_10162# a_25054_10162# 0.86fF
C7907 row_n[11] rowoff_n[11] 0.64fF
C7908 a_33086_8154# vcm 0.89fF
C7909 a_20034_12170# row_n[10] 0.43fF
C7910 a_8898_2130# a_8990_2130# 0.45fF
C7911 a_2275_2154# a_13310_2170# 0.15fF
C7912 a_2475_2154# a_15926_2130# 0.41fF
C7913 a_28370_11206# col_n[25] 0.11fF
C7914 a_2275_7174# m2_34864_6970# 0.51fF
C7915 a_19942_16186# rowon_n[14] 0.14fF
C7916 a_31078_15182# m2_31276_15430# 0.19fF
C7917 a_30074_2130# row_n[0] 0.43fF
C7918 a_7986_16186# VDD 3.92fF
C7919 a_15014_12170# a_15014_11166# 0.84fF
C7920 a_29982_6146# rowon_n[4] 0.14fF
C7921 a_23350_2170# vcm 0.24fF
C7922 a_2275_16210# col[26] 0.17fF
C7923 a_2275_16210# a_16930_16186# 0.17fF
C7924 a_2275_5166# col[31] 0.17fF
C7925 a_14010_11166# vcm 0.89fF
C7926 a_10906_1126# VDD 0.92fF
C7927 m2_1732_13998# row_n[12] 0.44fF
C7928 a_2275_4162# a_28370_4178# 0.15fF
C7929 a_2475_4162# a_30986_4138# 0.41fF
C7930 col_n[25] rowoff_n[12] 0.16fF
C7931 a_22042_9158# col[19] 0.38fF
C7932 a_2275_2154# col_n[1] 0.17fF
C7933 a_6982_10162# rowon_n[8] 0.45fF
C7934 a_4974_13174# a_5978_13174# 0.86fF
C7935 a_2475_13198# a_8990_13174# 0.68fF
C7936 a_30986_10162# rowoff_n[8] 0.42fF
C7937 a_4274_5182# vcm 0.24fF
C7938 a_34090_13174# rowoff_n[11] 1.10fF
C7939 a_2275_1150# a_21950_1126# 0.17fF
C7940 a_35002_6146# m2_34864_5966# 0.33fF
C7941 a_29070_15182# vcm 0.89fF
C7942 a_25966_5142# VDD 0.29fF
C7943 a_23958_6146# a_24050_6146# 0.45fF
C7944 m2_31852_946# VDD 2.95fF
C7945 a_22042_13174# m2_22240_13422# 0.19fF
C7946 a_17326_9198# col_n[14] 0.11fF
C7947 a_2475_15206# a_24050_15182# 0.68fF
C7948 a_30074_16186# a_30074_15182# 0.84fF
C7949 a_19334_9198# vcm 0.24fF
C7950 a_2475_9182# col[6] 0.22fF
C7951 a_32082_4138# ctop 4.91fF
C7952 a_9994_18194# vcm 0.15fF
C7953 col_n[9] rowoff_n[13] 0.27fF
C7954 a_28066_9158# row_n[7] 0.43fF
C7955 a_6890_8154# VDD 0.29fF
C7956 a_27974_13174# rowon_n[11] 0.14fF
C7957 col[12] rowoff_n[9] 0.27fF
C7958 col[11] rowoff_n[8] 0.27fF
C7959 col[10] rowoff_n[7] 0.28fF
C7960 col[9] rowoff_n[6] 0.29fF
C7961 col[8] rowoff_n[5] 0.29fF
C7962 col[7] rowoff_n[4] 0.30fF
C7963 col[6] rowoff_n[3] 0.31fF
C7964 col[5] rowoff_n[2] 0.31fF
C7965 col[3] rowoff_n[0] 0.33fF
C7966 col[4] rowoff_n[1] 0.32fF
C7967 a_2275_15206# col_n[13] 0.17fF
C7968 a_2275_12194# a_15014_12170# 0.71fF
C7969 a_10998_7150# col[8] 0.38fF
C7970 a_2275_4162# col_n[18] 0.17fF
C7971 a_12914_3134# vcm 0.18fF
C7972 a_20034_17190# a_21038_17190# 0.86fF
C7973 m2_29844_18014# m2_30848_18014# 0.86fF
C7974 a_35398_13214# vcm 0.24fF
C7975 a_26058_3134# col_n[23] 0.34fF
C7976 a_3270_15222# col_n[0] 0.11fF
C7977 a_13006_11166# m2_13204_11414# 0.19fF
C7978 a_13006_7150# ctop 4.91fF
C7979 a_21950_12170# VDD 0.29fF
C7980 a_2275_12194# col[3] 0.17fF
C7981 a_4882_9158# a_4974_9158# 0.45fF
C7982 a_2475_9182# a_7894_9158# 0.41fF
C7983 a_2275_9182# a_5278_9198# 0.15fF
C7984 a_4974_17190# rowon_n[15] 0.45fF
C7985 a_2275_1150# col[8] 0.17fF
C7986 a_6282_7190# col_n[3] 0.11fF
C7987 m2_1732_9982# sample_n 0.12fF
C7988 a_2275_14202# a_30074_14178# 0.71fF
C7989 a_3970_1126# m2_2736_946# 0.86fF
C7990 a_15014_7150# rowon_n[5] 0.45fF
C7991 a_27974_7150# vcm 0.18fF
C7992 a_22042_14178# rowoff_n[12] 1.69fF
C7993 a_2475_11190# col[23] 0.22fF
C7994 a_32082_7150# m2_32280_7398# 0.19fF
C7995 a_15318_16226# vcm 0.24fF
C7996 a_28066_11166# ctop 4.91fF
C7997 a_3878_9158# rowon_n[7] 0.14fF
C7998 a_2161_15206# VDD 0.23fF
C7999 a_2475_11190# a_22954_11166# 0.41fF
C8000 a_2275_11190# a_20338_11206# 0.15fF
C8001 a_2275_17214# col_n[30] 0.17fF
C8002 a_2275_18218# col_n[15] 0.17fF
C8003 a_8898_10162# vcm 0.18fF
C8004 a_3878_17190# rowoff_n[15] 0.73fF
C8005 a_9994_17190# col[7] 0.38fF
C8006 a_26058_16186# row_n[14] 0.43fF
C8007 a_3970_9158# m2_4168_9406# 0.19fF
C8008 a_30074_4138# a_31078_4138# 0.86fF
C8009 a_1957_6170# rowoff_n[4] 0.14fF
C8010 a_2275_8178# a_13918_8154# 0.17fF
C8011 a_2275_14202# col[20] 0.17fF
C8012 a_8990_14178# ctop 4.91fF
C8013 a_25054_13174# col_n[22] 0.34fF
C8014 a_2275_3158# col[25] 0.17fF
C8015 a_19942_13174# a_20034_13174# 0.45fF
C8016 a_5278_17230# col_n[2] 0.11fF
C8017 vcm col[10] 6.66fF
C8018 col_n[30] rowon_n[5] 0.17fF
C8019 col_n[28] rowon_n[4] 0.17fF
C8020 VDD col[13] 10.21fF
C8021 col_n[26] rowon_n[3] 0.17fF
C8022 col_n[24] rowon_n[2] 0.17fF
C8023 col_n[31] row_n[6] 0.37fF
C8024 col_n[19] row_n[0] 0.37fF
C8025 col_n[21] row_n[1] 0.37fF
C8026 col_n[5] col[5] 0.50fF
C8027 col_n[23] row_n[2] 0.37fF
C8028 col_n[25] row_n[3] 0.37fF
C8029 col_n[27] row_n[4] 0.37fF
C8030 col_n[20] rowon_n[0] 0.17fF
C8031 col_n[29] row_n[5] 0.37fF
C8032 col_n[22] rowon_n[1] 0.17fF
C8033 a_2966_7150# col_n[0] 0.34fF
C8034 a_23046_5142# m2_23244_5390# 0.19fF
C8035 a_23958_14178# vcm 0.18fF
C8036 a_20034_4138# VDD 2.68fF
C8037 a_21038_6146# a_21038_5142# 0.84fF
C8038 a_2475_5166# a_5978_5142# 0.68fF
C8039 a_2275_10186# a_28978_10162# 0.17fF
C8040 a_2874_9158# rowoff_n[7] 0.74fF
C8041 a_13006_14178# rowon_n[12] 0.45fF
C8042 a_9994_15182# rowoff_n[13] 2.28fF
C8043 a_1957_12194# row_n[10] 0.29fF
C8044 a_23046_4138# rowon_n[2] 0.45fF
C8045 a_4882_17190# vcm 0.18fF
C8046 a_12002_7150# rowoff_n[5] 2.18fF
C8047 a_10998_7150# a_12002_7150# 0.86fF
C8048 a_2475_7174# a_21038_7150# 0.68fF
C8049 a_2475_7174# col[0] 0.20fF
C8050 a_14010_11166# col_n[11] 0.34fF
C8051 a_6982_2130# vcm 0.89fF
C8052 a_35002_17190# a_35094_17190# 0.11fF
C8053 a_14010_3134# m2_14208_3382# 0.19fF
C8054 a_21038_5142# rowoff_n[3] 1.74fF
C8055 a_2275_4162# a_12002_4138# 0.71fF
C8056 a_2275_13198# col_n[7] 0.17fF
C8057 a_34090_13174# row_n[11] 0.43fF
C8058 a_16018_11166# VDD 3.09fF
C8059 a_2275_2154# col_n[12] 0.17fF
C8060 a_1957_17214# sample 0.35fF
C8061 a_33998_17190# rowon_n[15] 0.14fF
C8062 m2_34864_4962# vcm 0.72fF
C8063 a_30074_3134# rowoff_n[1] 1.30fF
C8064 a_22042_6146# vcm 0.89fF
C8065 a_2475_1150# a_4882_1126# 0.41fF
C8066 a_2275_1150# a_3878_1126# 0.15fF
C8067 a_34090_10162# col[31] 0.38fF
C8068 a_2275_6170# a_27062_6146# 0.71fF
C8069 a_31078_15182# VDD 1.54fF
C8070 a_26058_11166# a_27062_11166# 0.86fF
C8071 a_2475_9182# col[17] 0.22fF
C8072 m2_26832_18014# vcm 0.71fF
C8073 a_2275_15206# a_5886_15182# 0.17fF
C8074 a_21038_11166# rowon_n[9] 0.45fF
C8075 a_2874_9158# vcm 0.18fF
C8076 a_29374_10202# col_n[26] 0.11fF
C8077 col_n[20] rowoff_n[13] 0.19fF
C8078 a_10906_3134# a_10998_3134# 0.45fF
C8079 a_2275_3158# a_17326_3174# 0.15fF
C8080 a_2475_3158# a_19942_3134# 0.41fF
C8081 a_2275_1150# m2_16792_946# 0.51fF
C8082 m3_17928_1078# ctop 0.37fF
C8083 col[14] rowoff_n[0] 0.25fF
C8084 col[15] rowoff_n[1] 0.25fF
C8085 col[16] rowoff_n[2] 0.24fF
C8086 col[17] rowoff_n[3] 0.23fF
C8087 col[18] rowoff_n[4] 0.23fF
C8088 col[19] rowoff_n[5] 0.22fF
C8089 col[20] rowoff_n[6] 0.21fF
C8090 col[21] rowoff_n[7] 0.21fF
C8091 col[22] rowoff_n[8] 0.20fF
C8092 col[23] rowoff_n[9] 0.19fF
C8093 a_2275_15206# col_n[24] 0.17fF
C8094 a_2275_4162# col_n[29] 0.17fF
C8095 a_17022_13174# a_17022_12170# 0.84fF
C8096 a_27366_4178# vcm 0.24fF
C8097 a_2275_17214# a_20946_17190# 0.17fF
C8098 a_22954_11166# rowoff_n[9] 0.51fF
C8099 a_18026_13174# vcm 0.89fF
C8100 a_2275_12194# col[14] 0.17fF
C8101 a_14922_3134# VDD 0.29fF
C8102 a_2275_1150# col[19] 0.17fF
C8103 a_2475_5166# a_35002_5142# 0.41fF
C8104 a_2275_5166# a_32386_5182# 0.15fF
C8105 a_23046_8154# col[20] 0.38fF
C8106 a_3878_12170# VDD 0.29fF
C8107 a_8898_5142# rowon_n[3] 0.14fF
C8108 a_2275_18218# a_30986_18194# 0.17fF
C8109 a_31990_9158# rowoff_n[7] 0.41fF
C8110 a_2475_14202# a_13006_14178# 0.68fF
C8111 a_6982_14178# a_7986_14178# 0.86fF
C8112 col_n[4] rowoff_n[14] 0.31fF
C8113 m2_15788_18014# col[13] 0.39fF
C8114 a_8290_7190# vcm 0.24fF
C8115 m2_1732_6970# VDD 5.46fF
C8116 a_2275_2154# a_25966_2130# 0.17fF
C8117 a_33086_17190# vcm 0.89fF
C8118 a_21038_2130# ctop 4.93fF
C8119 a_18330_8194# col_n[15] 0.11fF
C8120 col[7] rowoff_n[10] 0.30fF
C8121 a_29982_7150# VDD 0.29fF
C8122 a_25966_7150# a_26058_7150# 0.45fF
C8123 a_2275_11190# a_3970_11166# 0.71fF
C8124 a_2275_18218# col_n[26] 0.17fF
C8125 a_34394_2170# vcm 0.24fF
C8126 a_32082_17190# a_32082_16186# 0.84fF
C8127 a_2475_16210# a_28066_16186# 0.68fF
C8128 a_2275_2154# m2_1732_1950# 0.27fF
C8129 a_23350_11206# vcm 0.24fF
C8130 a_21438_1488# VDD 0.14fF
C8131 a_29070_8154# rowon_n[6] 0.45fF
C8132 a_2275_14202# col[31] 0.17fF
C8133 a_10906_10162# VDD 0.29fF
C8134 a_12002_6146# col[9] 0.38fF
C8135 a_2275_13198# a_19030_13174# 0.71fF
C8136 col_n[30] row_n[0] 0.37fF
C8137 VDD col[24] 7.50fF
C8138 col_n[10] col[11] 6.22fF
C8139 col_n[31] rowon_n[0] 0.17fF
C8140 vcm col[21] 6.66fF
C8141 rowon_n[8] row_n[8] 21.02fF
C8142 a_16930_5142# vcm 0.18fF
C8143 a_10906_12170# rowoff_n[10] 0.65fF
C8144 a_2275_11190# col_n[1] 0.17fF
C8145 a_2275_18218# m2_10768_18014# 0.51fF
C8146 a_27062_2130# col_n[24] 0.34fF
C8147 a_6982_8154# row_n[6] 0.43fF
C8148 a_4274_14218# vcm 0.24fF
C8149 a_1957_4162# VDD 0.28fF
C8150 a_6890_12170# rowon_n[10] 0.14fF
C8151 a_17022_9158# ctop 4.91fF
C8152 m2_31852_18014# col_n[29] 0.32fF
C8153 a_7286_6186# col_n[4] 0.11fF
C8154 a_25966_14178# VDD 0.29fF
C8155 a_2966_4138# col[0] 0.38fF
C8156 a_2475_10186# a_11910_10162# 0.41fF
C8157 a_2275_10186# a_9294_10202# 0.15fF
C8158 a_6890_10162# a_6982_10162# 0.45fF
C8159 a_17326_18234# col_n[14] 0.11fF
C8160 a_2161_2154# rowoff_n[0] 0.14fF
C8161 a_16930_2130# rowon_n[0] 0.14fF
C8162 a_20034_1126# en_bit_n[0] 0.28fF
C8163 a_2275_15206# a_34090_15182# 0.71fF
C8164 m2_1732_9982# m2_2160_10410# 0.19fF
C8165 a_31990_9158# vcm 0.18fF
C8166 a_26970_16186# rowoff_n[14] 0.47fF
C8167 a_7986_3134# a_7986_2130# 0.84fF
C8168 a_19334_18234# vcm 0.25fF
C8169 a_2475_7174# col[11] 0.22fF
C8170 a_2161_7174# a_2275_7174# 0.17fF
C8171 a_2475_7174# a_2966_7150# 0.65fF
C8172 a_32082_13174# ctop 4.91fF
C8173 a_6890_17190# VDD 0.29fF
C8174 a_2475_12194# a_26970_12170# 0.41fF
C8175 a_2275_12194# a_24354_12210# 0.15fF
C8176 a_10998_16186# col[8] 0.38fF
C8177 a_27062_15182# rowon_n[13] 0.45fF
C8178 a_34090_4138# m2_34864_3958# 0.86fF
C8179 a_2275_13198# col_n[18] 0.17fF
C8180 a_12914_12170# vcm 0.18fF
C8181 a_2966_5142# rowoff_n[3] 2.62fF
C8182 a_8990_2130# VDD 3.82fF
C8183 a_2275_2154# col_n[23] 0.17fF
C8184 a_32082_5142# a_33086_5142# 0.86fF
C8185 a_26058_12170# col_n[23] 0.34fF
C8186 a_2275_9182# a_17934_9158# 0.17fF
C8187 a_13006_16186# ctop 4.91fF
C8188 a_21950_14178# a_22042_14178# 0.45fF
C8189 a_2275_10186# col[8] 0.17fF
C8190 a_6282_16226# col_n[3] 0.11fF
C8191 a_4974_15182# row_n[13] 0.43fF
C8192 a_27974_16186# vcm 0.18fF
C8193 a_24050_6146# VDD 2.27fF
C8194 a_15014_5142# row_n[3] 0.43fF
C8195 a_28066_14178# m2_28264_14426# 0.19fF
C8196 a_2475_6170# a_9994_6146# 0.68fF
C8197 a_23046_7150# a_23046_6146# 0.84fF
C8198 a_14922_9158# rowon_n[7] 0.14fF
C8199 m3_34568_1078# sw_n 0.10fF
C8200 a_2475_9182# col[28] 0.22fF
C8201 a_3970_8154# rowoff_n[6] 2.57fF
C8202 a_2275_11190# a_32994_11166# 0.17fF
C8203 col_n[31] rowoff_n[13] 0.11fF
C8204 a_30074_1126# vcm 0.15fF
C8205 m2_1732_16006# rowon_n[14] 0.43fF
C8206 m2_34864_13998# m2_34864_12994# 0.84fF
C8207 m2_34864_5966# rowoff_n[4] 1.01fF
C8208 a_2966_11166# rowon_n[9] 0.45fF
C8209 a_14922_17190# rowoff_n[15] 0.60fF
C8210 sample_n rowoff_n[7] 0.55fF
C8211 col[31] rowoff_n[6] 0.14fF
C8212 col[30] rowoff_n[5] 0.15fF
C8213 col[29] rowoff_n[4] 0.15fF
C8214 col[28] rowoff_n[3] 0.16fF
C8215 col[27] rowoff_n[2] 0.17fF
C8216 col[26] rowoff_n[1] 0.17fF
C8217 col[25] rowoff_n[0] 0.18fF
C8218 m2_30848_18014# VDD 2.44fF
C8219 a_13006_6146# rowoff_n[4] 2.13fF
C8220 m3_13912_18146# ctop 0.21fF
C8221 a_4974_9158# VDD 4.23fF
C8222 a_2475_8178# a_25054_8154# 0.68fF
C8223 a_13006_8154# a_14010_8154# 0.86fF
C8224 a_15014_10162# col_n[12] 0.34fF
C8225 a_2275_12194# col[25] 0.17fF
C8226 a_10998_4138# vcm 0.89fF
C8227 a_2475_3158# rowon_n[1] 0.40fF
C8228 a_22042_4138# rowoff_n[2] 1.69fF
C8229 a_2275_1150# col[30] 0.17fF
C8230 a_31990_1126# a_32082_1126# 0.11fF
C8231 a_2966_16186# col_n[0] 0.34fF
C8232 a_2275_5166# a_16018_5142# 0.71fF
C8233 a_19030_12170# m2_19228_12418# 0.19fF
C8234 a_20034_13174# VDD 2.68fF
C8235 a_2275_18218# a_11302_18234# 0.15fF
C8236 a_3970_10162# a_3970_9158# 0.84fF
C8237 col_n[15] rowoff_n[14] 0.23fF
C8238 a_31078_2130# rowoff_n[0] 1.25fF
C8239 col[18] rowoff_n[10] 0.23fF
C8240 a_26058_8154# vcm 0.89fF
C8241 a_13006_12170# row_n[10] 0.43fF
C8242 a_2275_2154# a_6282_2170# 0.15fF
C8243 a_2475_2154# a_8898_2130# 0.41fF
C8244 m2_22816_18014# m3_22948_18146# 4.43fF
C8245 a_12914_16186# rowon_n[14] 0.14fF
C8246 a_2275_7174# a_31078_7150# 0.71fF
C8247 a_23046_2130# row_n[0] 0.43fF
C8248 a_28066_12170# a_29070_12170# 0.86fF
C8249 a_22954_6146# rowon_n[4] 0.14fF
C8250 a_16322_2170# vcm 0.24fF
C8251 a_2275_16210# a_9902_16186# 0.17fF
C8252 a_30378_9198# col_n[27] 0.11fF
C8253 a_3970_8154# col_n[1] 0.34fF
C8254 a_2475_16210# col[0] 0.20fF
C8255 a_2475_5166# col[5] 0.22fF
C8256 a_6982_11166# vcm 0.89fF
C8257 a_3366_1488# VDD 0.19fF
C8258 a_12914_4138# a_13006_4138# 0.45fF
C8259 a_2475_4162# a_23958_4138# 0.41fF
C8260 a_2275_4162# a_21342_4178# 0.15fF
C8261 a_9994_10162# m2_10192_10410# 0.19fF
C8262 col_n[0] rowoff_n[15] 0.34fF
C8263 vcm sample_n 5.83fF
C8264 rowon_n[12] ctop 0.37fF
C8265 col_n[16] col[16] 0.43fF
C8266 a_2275_11190# col_n[12] 0.17fF
C8267 a_19030_14178# a_19030_13174# 0.84fF
C8268 a_23958_10162# rowoff_n[8] 0.50fF
C8269 col[2] rowoff_n[11] 0.33fF
C8270 a_31382_6186# vcm 0.24fF
C8271 a_27062_13174# rowoff_n[11] 1.45fF
C8272 a_2275_1150# a_14922_1126# 0.17fF
C8273 a_29070_6146# m2_29268_6394# 0.19fF
C8274 a_22042_15182# vcm 0.89fF
C8275 a_24050_7150# col[21] 0.38fF
C8276 a_18938_5142# VDD 0.29fF
C8277 a_2966_6146# a_2966_5142# 0.84fF
C8278 a_2275_8178# col[2] 0.17fF
C8279 a_32994_8154# rowoff_n[6] 0.40fF
C8280 a_8990_15182# a_9994_15182# 0.86fF
C8281 a_2475_15206# a_17022_15182# 0.68fF
C8282 a_12306_9198# vcm 0.24fF
C8283 a_2475_7174# col[22] 0.22fF
C8284 a_19334_7190# col_n[16] 0.11fF
C8285 a_2275_3158# a_29982_3134# 0.17fF
C8286 a_25054_4138# ctop 4.91fF
C8287 a_14922_1126# m2_14784_946# 0.31fF
C8288 a_33998_9158# VDD 0.29fF
C8289 a_21038_9158# row_n[7] 0.43fF
C8290 a_27974_8154# a_28066_8154# 0.45fF
C8291 a_20946_13174# rowon_n[11] 0.14fF
C8292 a_2275_12194# a_7986_12170# 0.71fF
C8293 a_2275_13198# col_n[29] 0.17fF
C8294 a_5886_3134# vcm 0.18fF
C8295 a_30986_3134# rowon_n[1] 0.14fF
C8296 a_2475_17214# a_32082_17190# 0.68fF
C8297 m2_22816_18014# m2_23820_18014# 0.86fF
C8298 a_20034_4138# m2_20232_4386# 0.19fF
C8299 a_27366_13214# vcm 0.24fF
C8300 a_5978_7150# ctop 4.91fF
C8301 a_14922_12170# VDD 0.29fF
C8302 a_13006_5142# col[10] 0.38fF
C8303 m2_27836_946# m2_28264_1374# 0.19fF
C8304 a_2275_10186# col[19] 0.17fF
C8305 a_23046_17190# col[20] 0.38fF
C8306 m2_1732_7974# vcm 1.11fF
C8307 a_2275_14202# a_23046_14178# 0.71fF
C8308 a_20946_7150# vcm 0.18fF
C8309 a_7986_7150# rowon_n[5] 0.45fF
C8310 a_15014_14178# rowoff_n[12] 2.03fF
C8311 a_19030_2130# a_20034_2130# 0.86fF
C8312 a_8290_16226# vcm 0.24fF
C8313 a_8290_5182# col_n[5] 0.11fF
C8314 a_21038_11166# ctop 4.91fF
C8315 a_18330_17230# col_n[15] 0.11fF
C8316 a_29982_16186# VDD 0.29fF
C8317 a_2275_11190# a_13310_11206# 0.15fF
C8318 a_2475_11190# a_15926_11166# 0.41fF
C8319 a_8898_11166# a_8990_11166# 0.45fF
C8320 a_34394_11206# vcm 0.24fF
C8321 a_19030_16186# row_n[14] 0.43fF
C8322 a_9994_4138# a_9994_3134# 0.84fF
C8323 a_2275_8178# a_6890_8154# 0.17fF
C8324 a_29070_6146# row_n[4] 0.43fF
C8325 a_28978_10162# rowon_n[8] 0.14fF
C8326 a_2275_13198# a_28370_13214# 0.15fF
C8327 a_2475_13198# a_30986_13174# 0.41fF
C8328 a_12002_15182# col[9] 0.38fF
C8329 a_16930_14178# vcm 0.18fF
C8330 a_13006_4138# VDD 3.40fF
C8331 a_27062_11166# col_n[24] 0.34fF
C8332 a_2275_9182# col_n[6] 0.17fF
C8333 col_n[26] rowoff_n[14] 0.15fF
C8334 a_1957_13198# VDD 0.28fF
C8335 a_2275_10186# a_21950_10162# 0.17fF
C8336 a_7286_15222# col_n[4] 0.11fF
C8337 col[29] rowoff_n[10] 0.15fF
C8338 a_5978_14178# rowon_n[12] 0.45fF
C8339 a_23958_15182# a_24050_15182# 0.45fF
C8340 a_2966_13174# col[0] 0.38fF
C8341 a_2874_15182# rowoff_n[13] 0.74fF
C8342 a_16018_4138# rowon_n[2] 0.45fF
C8343 a_31990_18194# vcm 0.18fF
C8344 a_28066_8154# VDD 1.85fF
C8345 a_4974_7150# rowoff_n[5] 2.52fF
C8346 a_2475_7174# a_14010_7150# 0.68fF
C8347 a_25054_8154# a_25054_7150# 0.84fF
C8348 a_2475_16210# col[11] 0.22fF
C8349 a_2475_5166# col[16] 0.22fF
C8350 a_34090_3134# vcm 0.89fF
C8351 a_14010_5142# rowoff_n[3] 2.08fF
C8352 col_n[10] rowoff_n[15] 0.27fF
C8353 col_n[21] col[22] 6.22fF
C8354 row_n[7] ctop 0.28fF
C8355 a_3878_4138# a_3970_4138# 0.45fF
C8356 a_2275_4162# a_4974_4138# 0.71fF
C8357 a_27062_13174# row_n[11] 0.43fF
C8358 a_8990_11166# VDD 3.82fF
C8359 a_2275_11190# col_n[23] 0.17fF
C8360 m2_29844_946# m3_29976_1078# 4.41fF
C8361 a_2475_9182# a_29070_9158# 0.68fF
C8362 a_26970_17190# rowon_n[15] 0.14fF
C8363 a_15014_9158# a_16018_9158# 0.86fF
C8364 a_16018_9158# col_n[13] 0.34fF
C8365 col[13] rowoff_n[11] 0.26fF
C8366 m2_34864_2954# rowon_n[1] 0.42fF
C8367 a_23046_3134# rowoff_n[1] 1.64fF
C8368 a_15014_6146# vcm 0.89fF
C8369 a_4882_18194# a_4974_18194# 0.11fF
C8370 a_33998_2130# a_34090_2130# 0.48fF
C8371 a_2275_8178# col[13] 0.17fF
C8372 a_2275_6170# a_20034_6146# 0.71fF
C8373 a_24050_15182# VDD 2.27fF
C8374 a_5978_11166# a_5978_10162# 0.84fF
C8375 m2_12776_18014# vcm 0.71fF
C8376 a_14010_11166# rowon_n[9] 0.45fF
C8377 a_30074_10162# vcm 0.89fF
C8378 a_2475_3158# a_12914_3134# 0.41fF
C8379 a_2275_3158# a_10298_3174# 0.15fF
C8380 a_26058_2130# m2_25828_946# 0.84fF
C8381 m3_34996_7102# ctop 0.22fF
C8382 a_2966_9158# row_n[7] 0.41fF
C8383 a_2275_8178# a_35094_8154# 0.14fF
C8384 a_2475_16210# m2_34864_16006# 0.56fF
C8385 a_2275_13198# rowon_n[11] 1.99fF
C8386 a_30074_13174# a_31078_13174# 0.86fF
C8387 a_4974_7150# col_n[2] 0.34fF
C8388 a_31382_8194# col_n[28] 0.11fF
C8389 a_20338_4178# vcm 0.24fF
C8390 a_15926_11166# rowoff_n[9] 0.59fF
C8391 a_2275_17214# a_13918_17190# 0.17fF
C8392 a_10998_13174# vcm 0.89fF
C8393 a_7894_3134# VDD 0.29fF
C8394 a_2275_10186# col[30] 0.17fF
C8395 a_2475_5166# a_27974_5142# 0.41fF
C8396 a_2275_5166# a_25358_5182# 0.15fF
C8397 a_14922_5142# a_15014_5142# 0.45fF
C8398 a_2275_18218# a_23958_18194# 0.17fF
C8399 a_24962_9158# rowoff_n[7] 0.49fF
C8400 a_35002_14178# rowon_n[12] 0.14fF
C8401 a_2475_14202# a_5978_14178# 0.68fF
C8402 a_21038_15182# a_21038_14178# 0.84fF
C8403 a_2275_7174# vcm 7.71fF
C8404 a_31990_15182# rowoff_n[13] 0.41fF
C8405 a_25054_6146# col[22] 0.38fF
C8406 m2_1732_4962# row_n[3] 0.44fF
C8407 a_2275_2154# a_18938_2130# 0.17fF
C8408 a_14010_2130# ctop 4.93fF
C8409 a_26058_17190# vcm 0.89fF
C8410 a_22954_7150# VDD 0.29fF
C8411 a_33998_7150# rowoff_n[5] 0.39fF
C8412 a_34090_15182# m2_34288_15430# 0.19fF
C8413 a_2966_11166# ctop 4.82fF
C8414 a_28978_2130# vcm 0.18fF
C8415 a_10998_16186# a_12002_16186# 0.86fF
C8416 a_2475_16210# a_21038_16186# 0.68fF
C8417 a_20338_6186# col_n[17] 0.11fF
C8418 a_16322_11206# vcm 0.24fF
C8419 a_30378_18234# col_n[27] 0.11fF
C8420 a_3970_17190# col_n[1] 0.34fF
C8421 a_14410_1488# VDD 0.16fF
C8422 a_22042_8154# rowon_n[6] 0.45fF
C8423 a_2275_4162# a_33998_4138# 0.17fF
C8424 a_2475_14202# col[5] 0.22fF
C8425 a_29070_6146# ctop 4.91fF
C8426 a_2475_3158# col[10] 0.22fF
C8427 m3_32988_1078# m3_33992_1078# 0.21fF
C8428 a_29982_9158# a_30074_9158# 0.45fF
C8429 a_5978_17190# m2_6176_17438# 0.19fF
C8430 a_2275_13198# a_12002_13174# 0.71fF
C8431 a_9902_5142# vcm 0.18fF
C8432 a_2275_9182# col_n[17] 0.17fF
C8433 a_2966_5142# m2_3164_5390# 0.19fF
C8434 a_31382_15222# vcm 0.24fF
C8435 a_14010_4138# col[11] 0.38fF
C8436 a_25054_13174# m2_25252_13422# 0.19fF
C8437 a_33086_17190# row_n[15] 0.43fF
C8438 a_9994_9158# ctop 4.91fF
C8439 a_24050_16186# col[21] 0.38fF
C8440 a_18938_14178# VDD 0.29fF
C8441 a_2275_10186# a_3878_10162# 0.17fF
C8442 a_2475_10186# a_4882_10162# 0.41fF
C8443 a_2275_17214# col[2] 0.17fF
C8444 a_9902_2130# rowon_n[0] 0.14fF
C8445 m2_28840_946# col[26] 0.52fF
C8446 a_2275_6170# col[7] 0.17fF
C8447 a_2275_15206# a_27062_15182# 0.71fF
C8448 a_24962_9158# vcm 0.18fF
C8449 a_19942_16186# rowoff_n[14] 0.55fF
C8450 a_9294_4178# col_n[6] 0.11fF
C8451 a_21038_3134# a_22042_3134# 0.86fF
C8452 a_12306_18234# vcm 0.25fF
C8453 a_19334_16226# col_n[16] 0.11fF
C8454 a_2475_16210# col[22] 0.22fF
C8455 a_25054_13174# ctop 4.91fF
C8456 a_2475_5166# col[27] 0.22fF
C8457 a_33998_18194# VDD 0.50fF
C8458 a_2275_12194# a_17326_12210# 0.15fF
C8459 a_2475_12194# a_19942_12170# 0.41fF
C8460 a_10906_12170# a_10998_12170# 0.45fF
C8461 rowon_n[1] ctop 0.37fF
C8462 col_n[21] rowoff_n[15] 0.19fF
C8463 col_n[27] col[27] 0.55fF
C8464 a_20034_15182# rowon_n[13] 0.45fF
C8465 m2_33860_18014# m2_34288_18442# 0.19fF
C8466 a_5886_12170# vcm 0.18fF
C8467 a_2475_2154# VDD 41.97fF
C8468 col[24] rowoff_n[11] 0.19fF
C8469 a_16018_11166# m2_16216_11414# 0.19fF
C8470 a_12002_5142# a_12002_4138# 0.84fF
C8471 a_30074_5142# rowon_n[3] 0.45fF
C8472 a_8898_18194# m2_8760_18014# 0.34fF
C8473 a_2275_9182# a_10906_9158# 0.17fF
C8474 a_5978_16186# ctop 4.91fF
C8475 a_13006_14178# col[10] 0.38fF
C8476 a_2475_18218# m2_22816_18014# 0.62fF
C8477 a_2275_14202# a_32386_14218# 0.15fF
C8478 a_2475_14202# a_35002_14178# 0.41fF
C8479 a_2275_8178# col[24] 0.17fF
C8480 a_28066_10162# col_n[25] 0.34fF
C8481 a_20946_16186# vcm 0.18fF
C8482 a_17022_6146# VDD 2.99fF
C8483 a_7986_5142# row_n[3] 0.43fF
C8484 a_1957_6170# a_2275_6170# 0.19fF
C8485 a_2475_6170# a_2874_6146# 0.41fF
C8486 a_7894_9158# rowon_n[7] 0.14fF
C8487 a_8290_14218# col_n[5] 0.11fF
C8488 a_2275_11190# a_25966_11166# 0.17fF
C8489 a_23046_1126# vcm 0.15fF
C8490 a_25966_16186# a_26058_16186# 0.45fF
C8491 a_7894_17190# rowoff_n[15] 0.68fF
C8492 col[8] rowoff_n[12] 0.29fF
C8493 m2_16792_18014# VDD 3.78fF
C8494 a_5978_6146# rowoff_n[4] 2.47fF
C8495 a_6982_9158# m2_7180_9406# 0.19fF
C8496 a_32082_10162# VDD 1.44fF
C8497 a_27062_9158# a_27062_8154# 0.84fF
C8498 a_2475_8178# a_18026_8154# 0.68fF
C8499 a_3970_4138# vcm 0.89fF
C8500 a_15014_4138# rowoff_n[2] 2.03fF
C8501 a_32082_12170# rowoff_n[10] 1.20fF
C8502 a_2475_1150# col[4] 0.22fF
C8503 a_26058_5142# m2_26256_5390# 0.19fF
C8504 a_28066_12170# rowon_n[10] 0.45fF
C8505 a_2275_5166# a_8990_5142# 0.71fF
C8506 a_17022_8154# col_n[14] 0.34fF
C8507 a_2275_18218# a_4274_18234# 0.15fF
C8508 a_13006_13174# VDD 3.40fF
C8509 a_2475_10186# a_33086_10162# 0.68fF
C8510 a_17022_10162# a_18026_10162# 0.86fF
C8511 a_24050_2130# rowoff_n[0] 1.59fF
C8512 a_2275_7174# col_n[11] 0.17fF
C8513 a_19030_8154# vcm 0.89fF
C8514 a_5978_12170# row_n[10] 0.43fF
C8515 a_5886_16186# rowon_n[14] 0.14fF
C8516 a_2275_7174# a_24050_7150# 0.71fF
C8517 a_2275_4162# col[1] 0.17fF
C8518 a_16018_2130# row_n[0] 0.43fF
C8519 a_28066_17190# VDD 1.85fF
C8520 a_7986_12170# a_7986_11166# 0.84fF
C8521 a_15926_6146# rowon_n[4] 0.14fF
C8522 a_9294_2170# vcm 0.24fF
C8523 a_2161_16210# a_2275_16210# 0.17fF
C8524 a_2475_16210# a_2966_16186# 0.65fF
C8525 a_2475_14202# col[16] 0.22fF
C8526 a_17022_3134# m2_17220_3382# 0.19fF
C8527 a_34090_12170# vcm 0.89fF
C8528 a_2475_3158# col[21] 0.22fF
C8529 a_30986_2130# VDD 0.29fF
C8530 a_2475_4162# a_16930_4138# 0.41fF
C8531 a_2275_4162# a_14314_4178# 0.15fF
C8532 a_2475_18218# col[7] 0.22fF
C8533 m3_1864_3086# m3_1864_2082# 0.20fF
C8534 a_27974_18194# m2_27836_18014# 0.34fF
C8535 a_4974_17190# m2_4744_18014# 0.84fF
C8536 a_5978_6146# col_n[3] 0.34fF
C8537 a_32386_7190# col_n[29] 0.11fF
C8538 a_32082_14178# a_33086_14178# 0.86fF
C8539 a_16930_10162# rowoff_n[8] 0.58fF
C8540 a_2275_9182# col_n[28] 0.17fF
C8541 a_24354_6186# vcm 0.24fF
C8542 a_20034_13174# rowoff_n[11] 1.79fF
C8543 a_2275_1150# a_7894_1126# 0.17fF
C8544 a_15014_15182# vcm 0.89fF
C8545 a_11910_5142# VDD 0.29fF
C8546 a_2275_6170# a_29374_6186# 0.15fF
C8547 a_2475_6170# a_31990_6146# 0.41fF
C8548 a_16930_6146# a_17022_6146# 0.45fF
C8549 a_2275_17214# col[13] 0.17fF
C8550 a_25966_8154# rowoff_n[6] 0.48fF
C8551 a_2275_6170# col[18] 0.17fF
C8552 a_23046_16186# a_23046_15182# 0.84fF
C8553 a_2475_15206# a_9994_15182# 0.68fF
C8554 a_26058_5142# col[23] 0.38fF
C8555 a_5278_9198# vcm 0.24fF
C8556 a_35002_6146# rowoff_n[4] 0.38fF
C8557 a_2275_3158# a_22954_3134# 0.17fF
C8558 a_18026_4138# ctop 4.91fF
C8559 a_2275_1150# m2_25828_946# 0.51fF
C8560 m3_32988_1078# ctop 0.21fF
C8561 a_14010_9158# row_n[7] 0.43fF
C8562 a_26970_9158# VDD 0.29fF
C8563 a_13918_13174# rowon_n[11] 0.14fF
C8564 ctop analog_in 0.79fF
C8565 rowon_n[15] rowoff_n[15] 20.65fF
C8566 row_n[15] sample_n 0.16fF
C8567 a_21342_5182# col_n[18] 0.11fF
C8568 a_32994_4138# vcm 0.18fF
C8569 a_2275_11190# row_n[9] 26.41fF
C8570 a_23958_3134# rowon_n[1] 0.14fF
C8571 a_2475_17214# a_25054_17190# 0.68fF
C8572 a_13006_17190# a_14010_17190# 0.86fF
C8573 a_4974_16186# col_n[2] 0.34fF
C8574 a_31382_17230# col_n[28] 0.11fF
C8575 m2_15788_18014# m2_16792_18014# 0.86fF
C8576 a_20338_13214# vcm 0.24fF
C8577 a_2475_11190# m2_1732_10986# 0.16fF
C8578 a_33086_8154# ctop 4.91fF
C8579 a_7894_12170# VDD 0.29fF
C8580 m2_20808_946# m2_21236_1374# 0.19fF
C8581 a_31990_10162# a_32082_10162# 0.45fF
C8582 a_2275_14202# a_16018_14178# 0.71fF
C8583 a_13918_7150# vcm 0.18fF
C8584 a_7986_14178# rowoff_n[12] 2.38fF
C8585 a_2475_2154# a_30074_2130# 0.68fF
C8586 a_33086_3134# a_33086_2130# 0.84fF
C8587 a_15014_3134# col[12] 0.38fF
C8588 a_2275_16210# vcm 7.71fF
C8589 a_34090_16186# rowon_n[14] 0.45fF
C8590 a_25054_15182# col[22] 0.38fF
C8591 a_2275_5166# col_n[5] 0.17fF
C8592 a_14010_11166# ctop 4.91fF
C8593 a_22954_16186# VDD 0.29fF
C8594 m2_34864_15002# rowoff_n[13] 1.01fF
C8595 a_2275_11190# a_6282_11206# 0.15fF
C8596 a_2475_11190# a_8898_11166# 0.41fF
C8597 col[19] rowoff_n[12] 0.22fF
C8598 a_2275_16210# a_31078_16186# 0.71fF
C8599 a_10298_3174# col_n[7] 0.11fF
C8600 a_28978_11166# vcm 0.18fF
C8601 a_25054_1126# VDD 0.10fF
C8602 a_12002_16186# row_n[14] 0.43fF
C8603 a_20338_15222# col_n[17] 0.11fF
C8604 a_23046_4138# a_24050_4138# 0.86fF
C8605 a_24050_17190# m2_23820_18014# 0.84fF
C8606 a_29070_15182# ctop 4.91fF
C8607 a_22042_6146# row_n[4] 0.43fF
C8608 a_2475_12194# col[10] 0.22fF
C8609 a_21950_10162# rowon_n[8] 0.14fF
C8610 a_12914_13174# a_13006_13174# 0.45fF
C8611 a_2475_13198# a_23958_13174# 0.41fF
C8612 a_2275_13198# a_21342_13214# 0.15fF
C8613 a_2475_1150# col[15] 0.22fF
C8614 a_9902_14178# vcm 0.18fF
C8615 a_5978_4138# VDD 4.13fF
C8616 a_14010_6146# a_14010_5142# 0.84fF
C8617 a_3970_1126# col[1] 0.53fF
C8618 a_2275_7174# col_n[22] 0.17fF
C8619 a_14010_13174# col[11] 0.38fF
C8620 a_2275_10186# a_14922_10162# 0.17fF
C8621 col[3] rowoff_n[13] 0.33fF
C8622 a_2966_15182# a_2966_14178# 0.84fF
C8623 a_29070_9158# col_n[26] 0.34fF
C8624 a_2275_15206# col[7] 0.17fF
C8625 a_2275_4162# col[12] 0.17fF
C8626 a_8990_4138# rowon_n[2] 0.45fF
C8627 a_24962_18194# vcm 0.18fF
C8628 a_21038_8154# VDD 2.58fF
C8629 a_2475_7174# a_6982_7150# 0.68fF
C8630 a_9294_13214# col_n[6] 0.11fF
C8631 a_3970_7150# a_4974_7150# 0.86fF
C8632 m2_9764_18014# col[7] 0.39fF
C8633 a_2275_12194# a_29982_12170# 0.17fF
C8634 a_2475_14202# col[27] 0.22fF
C8635 a_27062_3134# vcm 0.89fF
C8636 a_27974_17190# a_28066_17190# 0.45fF
C8637 m2_1732_17010# m2_1732_16006# 0.84fF
C8638 a_2966_3134# m2_1732_2954# 0.86fF
C8639 a_2475_18218# col[18] 0.22fF
C8640 a_6982_5142# rowoff_n[3] 2.42fF
C8641 a_20034_13174# row_n[11] 0.43fF
C8642 a_2475_11190# VDD 41.96fF
C8643 m3_28972_18146# m3_29976_18146# 0.21fF
C8644 a_19942_17190# rowon_n[15] 0.14fF
C8645 a_29070_10162# a_29070_9158# 0.84fF
C8646 a_2475_9182# a_22042_9158# 0.68fF
C8647 m2_1732_6970# rowon_n[5] 0.43fF
C8648 a_16018_3134# rowoff_n[1] 1.98fF
C8649 a_30074_3134# row_n[1] 0.43fF
C8650 a_7986_6146# vcm 0.89fF
C8651 a_29982_7150# rowon_n[5] 0.14fF
C8652 a_1957_13198# rowoff_n[11] 0.14fF
C8653 a_2275_6170# m2_34864_5966# 0.51fF
C8654 a_2275_17214# col[24] 0.17fF
C8655 a_18026_7150# col_n[15] 0.34fF
C8656 a_2275_6170# col[29] 0.17fF
C8657 a_2275_18218# col[9] 0.17fF
C8658 a_2275_6170# a_13006_6146# 0.71fF
C8659 a_31078_14178# m2_31276_14426# 0.19fF
C8660 a_17022_15182# VDD 2.99fF
C8661 a_19030_11166# a_20034_11166# 0.86fF
C8662 m2_1732_10986# rowoff_n[9] 2.46fF
C8663 a_32386_1166# vcm 0.25fF
C8664 a_6982_11166# rowon_n[9] 0.45fF
C8665 a_2275_3158# col_n[0] 0.17fF
C8666 a_23046_10162# vcm 0.89fF
C8667 m2_25828_18014# col_n[23] 0.34fF
C8668 a_2475_3158# a_5886_3134# 0.41fF
C8669 a_2275_3158# a_3270_3174# 0.15fF
C8670 m3_28972_18146# ctop 0.21fF
C8671 ctop col[10] 0.13fF
C8672 rowon_n[9] sample_n 0.15fF
C8673 a_2275_8178# a_28066_8154# 0.71fF
C8674 a_9994_13174# a_9994_12170# 0.84fF
C8675 a_13310_4178# vcm 0.24fF
C8676 a_8898_11166# rowoff_n[9] 0.67fF
C8677 a_2275_17214# a_6890_17190# 0.17fF
C8678 a_35002_5142# m2_34864_4962# 0.33fF
C8679 a_3970_13174# vcm 0.89fF
C8680 a_35002_4138# VDD 0.36fF
C8681 a_2475_10186# col[4] 0.22fF
C8682 a_2275_5166# a_18330_5182# 0.15fF
C8683 a_2475_5166# a_20946_5142# 0.41fF
C8684 a_22042_12170# m2_22240_12418# 0.19fF
C8685 a_2275_18218# a_16930_18194# 0.17fF
C8686 a_33390_6186# col_n[30] 0.11fF
C8687 a_6982_5142# col_n[4] 0.34fF
C8688 a_28066_10162# row_n[8] 0.43fF
C8689 a_17022_17190# col_n[14] 0.34fF
C8690 a_17934_9158# rowoff_n[7] 0.57fF
C8691 a_27974_14178# rowon_n[12] 0.14fF
C8692 a_2275_16210# col_n[11] 0.17fF
C8693 a_28370_8194# vcm 0.24fF
C8694 a_24962_15182# rowoff_n[13] 0.49fF
C8695 a_2275_5166# col_n[16] 0.17fF
C8696 a_2275_2154# a_11910_2130# 0.17fF
C8697 a_19030_17190# vcm 0.89fF
C8698 a_6982_2130# ctop 4.93fF
C8699 m2_27836_18014# m3_27968_18146# 4.43fF
C8700 a_15926_7150# VDD 0.29fF
C8701 a_26970_7150# rowoff_n[5] 0.47fF
C8702 a_2275_7174# a_33390_7190# 0.15fF
C8703 a_18938_7150# a_19030_7150# 0.45fF
C8704 col[30] rowoff_n[12] 0.15fF
C8705 m2_1732_16006# rowoff_n[14] 2.46fF
C8706 a_2275_13198# col[1] 0.17fF
C8707 a_27062_4138# col[24] 0.38fF
C8708 a_21950_2130# vcm 0.18fF
C8709 a_2275_2154# col[6] 0.17fF
C8710 a_2475_16210# a_14010_16186# 0.68fF
C8711 a_25054_17190# a_25054_16186# 0.84fF
C8712 m2_1732_10986# sample 0.31fF
C8713 a_9294_11206# vcm 0.24fF
C8714 a_7382_1488# VDD 0.18fF
C8715 a_15014_8154# rowon_n[6] 0.45fF
C8716 a_2275_4162# a_26970_4138# 0.17fF
C8717 a_13006_10162# m2_13204_10410# 0.19fF
C8718 a_22042_6146# ctop 4.91fF
C8719 a_2475_12194# col[21] 0.22fF
C8720 a_30986_11166# VDD 0.29fF
C8721 m3_18932_1078# m3_19936_1078# 0.12fF
C8722 a_2475_1150# col[26] 0.22fF
C8723 a_22346_4178# col_n[19] 0.11fF
C8724 a_3878_10162# rowon_n[8] 0.14fF
C8725 a_2275_13198# a_4974_13174# 0.71fF
C8726 a_3878_13174# a_3970_13174# 0.45fF
C8727 a_5978_15182# col_n[3] 0.34fF
C8728 a_32386_16226# col_n[29] 0.11fF
C8729 m2_34864_4962# m2_35292_5390# 0.19fF
C8730 a_32082_6146# m2_32280_6394# 0.19fF
C8731 a_2475_1150# a_19030_1126# 0.66fF
C8732 a_24354_15222# vcm 0.24fF
C8733 a_2475_18218# a_29982_18194# 0.41fF
C8734 a_26058_17190# row_n[15] 0.43fF
C8735 col[14] rowoff_n[13] 0.25fF
C8736 a_11910_14178# VDD 0.29fF
C8737 a_33998_11166# a_34090_11166# 0.45fF
C8738 VDD rowoff_n[9] 87.22fF
C8739 a_2275_15206# col[18] 0.17fF
C8740 a_2275_15206# a_20034_15182# 0.71fF
C8741 a_2275_4162# col[23] 0.17fF
C8742 a_16018_2130# col[13] 0.38fF
C8743 a_17934_9158# vcm 0.18fF
C8744 a_12914_16186# rowoff_n[14] 0.63fF
C8745 a_26058_14178# col[23] 0.38fF
C8746 a_2475_3158# a_34090_3134# 0.68fF
C8747 a_3970_8154# m2_4168_8402# 0.19fF
C8748 a_5278_18234# vcm 0.25fF
C8749 a_2966_8154# VDD 4.45fF
C8750 a_18026_13174# ctop 4.91fF
C8751 a_26970_18194# VDD 0.50fF
C8752 a_2275_12194# a_10298_12210# 0.15fF
C8753 a_2475_12194# a_12914_12170# 0.41fF
C8754 a_2475_18218# col[29] 0.22fF
C8755 a_11302_2170# col_n[8] 0.11fF
C8756 a_2275_17214# a_35094_17190# 0.14fF
C8757 a_13006_15182# rowon_n[13] 0.45fF
C8758 m2_26832_18014# m2_27260_18442# 0.19fF
C8759 a_23046_4138# m2_23244_4386# 0.19fF
C8760 a_21342_14218# col_n[18] 0.11fF
C8761 a_32994_13174# vcm 0.18fF
C8762 a_29070_3134# VDD 1.75fF
C8763 a_25054_5142# a_26058_5142# 0.86fF
C8764 a_1957_13198# row_n[11] 0.29fF
C8765 a_23046_5142# rowon_n[3] 0.45fF
C8766 a_2874_9158# a_2966_9158# 0.45fF
C8767 m2_12776_946# col[10] 0.51fF
C8768 a_33086_17190# ctop 4.93fF
C8769 a_2475_18218# m2_8760_18014# 0.62fF
C8770 a_14922_14178# a_15014_14178# 0.45fF
C8771 a_2275_14202# a_25358_14218# 0.15fF
C8772 a_2475_14202# a_27974_14178# 0.41fF
C8773 a_2275_18218# col[20] 0.17fF
C8774 a_13918_16186# vcm 0.18fF
C8775 a_9994_6146# VDD 3.71fF
C8776 a_16018_7150# a_16018_6146# 0.84fF
C8777 a_15014_12170# col[12] 0.38fF
C8778 a_2275_14202# col_n[5] 0.17fF
C8779 a_2275_11190# a_18938_11166# 0.17fF
C8780 a_34090_14178# row_n[12] 0.43fF
C8781 a_2275_3158# col_n[10] 0.17fF
C8782 a_16018_1126# vcm 0.15fF
C8783 a_30074_8154# col_n[27] 0.34fF
C8784 VDD sample 6.38fF
C8785 ctop col[21] 0.13fF
C8786 m2_2736_18014# VDD 5.31fF
C8787 en_bit_n[0] col[17] 0.14fF
C8788 row_n[4] sample_n 0.16fF
C8789 a_10298_12210# col_n[7] 0.11fF
C8790 a_8990_2130# m2_8760_946# 0.84fF
C8791 a_25054_10162# VDD 2.16fF
C8792 a_2475_8178# a_10998_8154# 0.68fF
C8793 a_5978_8154# a_6982_8154# 0.86fF
C8794 a_2275_13198# a_33998_13174# 0.17fF
C8795 a_31078_5142# vcm 0.89fF
C8796 a_7986_4138# rowoff_n[2] 2.38fF
C8797 a_25054_12170# rowoff_n[10] 1.54fF
C8798 a_29982_18194# a_30074_18194# 0.11fF
C8799 a_2475_10186# col[15] 0.22fF
C8800 a_24962_1126# a_25054_1126# 0.11fF
C8801 a_21038_12170# rowon_n[10] 0.45fF
C8802 a_1957_5166# a_2161_5166# 0.11fF
C8803 a_2475_5166# a_2275_5166# 2.96fF
C8804 a_5978_13174# VDD 4.13fF
C8805 a_31078_11166# a_31078_10162# 0.84fF
C8806 a_2475_10186# a_26058_10162# 0.68fF
C8807 a_3970_10162# col[1] 0.38fF
C8808 a_31078_2130# rowon_n[0] 0.45fF
C8809 a_2275_16210# col_n[22] 0.17fF
C8810 a_17022_2130# rowoff_n[0] 1.94fF
C8811 a_2275_5166# col_n[27] 0.17fF
C8812 a_12002_8154# vcm 0.89fF
C8813 a_19030_6146# col_n[16] 0.34fF
C8814 a_2275_7174# a_17022_7150# 0.71fF
C8815 a_2275_13198# col[12] 0.17fF
C8816 a_8990_2130# row_n[0] 0.43fF
C8817 a_2275_2154# col[17] 0.17fF
C8818 a_21038_17190# VDD 2.58fF
C8819 a_21038_12170# a_22042_12170# 0.86fF
C8820 a_8898_6146# rowon_n[4] 0.14fF
C8821 a_3878_2130# vcm 0.18fF
C8822 a_27062_12170# vcm 0.89fF
C8823 a_23958_2130# VDD 0.29fF
C8824 a_2275_4162# a_7286_4178# 0.15fF
C8825 a_2475_4162# a_9902_4138# 0.41fF
C8826 a_5886_4138# a_5978_4138# 0.45fF
C8827 m3_1864_10114# m3_1864_9110# 0.20fF
C8828 m2_34864_946# m3_34996_1078# 4.42fF
C8829 a_2275_9182# a_32082_9158# 0.71fF
C8830 a_12002_14178# a_12002_13174# 0.84fF
C8831 a_9902_10162# rowoff_n[8] 0.66fF
C8832 a_17326_6186# vcm 0.24fF
C8833 a_13006_13174# rowoff_n[11] 2.13fF
C8834 a_7986_15182# vcm 0.89fF
C8835 col[25] rowoff_n[13] 0.18fF
C8836 a_4882_5142# VDD 0.29fF
C8837 a_7986_4138# col_n[5] 0.34fF
C8838 a_2275_6170# a_22346_6186# 0.15fF
C8839 a_2475_6170# a_24962_6146# 0.41fF
C8840 col_n[3] rowoff_n[4] 0.32fF
C8841 col_n[1] rowoff_n[2] 0.33fF
C8842 col_n[6] rowoff_n[7] 0.29fF
C8843 col_n[2] rowoff_n[3] 0.32fF
C8844 col_n[5] rowoff_n[6] 0.30fF
C8845 col_n[7] rowoff_n[8] 0.29fF
C8846 vcm rowoff_n[1] 2.43fF
C8847 col_n[4] rowoff_n[5] 0.31fF
C8848 col_n[0] rowoff_n[0] 0.34fF
C8849 col_n[8] rowoff_n[9] 0.28fF
C8850 a_18026_16186# col_n[15] 0.34fF
C8851 a_29070_9158# rowon_n[7] 0.45fF
C8852 a_2275_15206# col[29] 0.17fF
C8853 a_18938_8154# rowoff_n[6] 0.56fF
C8854 a_1957_15206# a_2275_15206# 0.19fF
C8855 a_2475_15206# a_2874_15182# 0.41fF
C8856 a_32386_10202# vcm 0.24fF
C8857 a_29070_17190# rowoff_n[15] 1.35fF
C8858 a_2275_12194# col_n[0] 0.17fF
C8859 a_27974_6146# rowoff_n[4] 0.46fF
C8860 a_2275_3158# a_15926_3134# 0.17fF
C8861 a_10998_4138# ctop 4.91fF
C8862 a_2475_1150# m2_11772_946# 0.62fF
C8863 a_6982_9158# row_n[7] 0.43fF
C8864 m3_4876_1078# ctop 0.21fF
C8865 a_19942_9158# VDD 0.29fF
C8866 a_2275_1150# col_n[4] 0.17fF
C8867 a_20946_8154# a_21038_8154# 0.45fF
C8868 a_6890_13174# rowon_n[11] 0.14fF
C8869 a_28066_3134# col[25] 0.38fF
C8870 a_25966_4138# vcm 0.18fF
C8871 m2_1732_946# sample 0.31fF
C8872 a_16930_3134# rowon_n[1] 0.14fF
C8873 a_2475_17214# a_18026_17190# 0.68fF
C8874 col[9] rowoff_n[14] 0.29fF
C8875 m2_8760_18014# m2_9764_18014# 0.86fF
C8876 a_13310_13214# vcm 0.24fF
C8877 a_2275_5166# a_30986_5142# 0.17fF
C8878 a_26058_8154# ctop 4.91fF
C8879 a_35002_13174# VDD 0.36fF
C8880 a_23350_3174# col_n[20] 0.11fF
C8881 a_2475_8178# col[9] 0.22fF
C8882 a_33390_15222# col_n[30] 0.11fF
C8883 a_6982_14178# col_n[4] 0.34fF
C8884 a_2275_14202# a_8990_14178# 0.71fF
C8885 a_2275_18218# col[31] 0.17fF
C8886 a_6890_7150# vcm 0.18fF
C8887 a_2475_2154# a_23046_2130# 0.68fF
C8888 a_12002_2130# a_13006_2130# 0.86fF
C8889 a_28370_17230# vcm 0.24fF
C8890 a_27062_16186# rowon_n[14] 0.45fF
C8891 a_2275_14202# col_n[16] 0.17fF
C8892 a_6982_11166# ctop 4.91fF
C8893 a_2275_3158# col_n[21] 0.17fF
C8894 a_15926_16186# VDD 0.29fF
C8895 vcm col_n[6] 3.22fF
C8896 VDD col_n[9] 14.20fF
C8897 a_2275_16210# a_24050_16186# 0.71fF
C8898 a_34090_3134# m2_34864_2954# 0.86fF
C8899 a_27062_13174# col[24] 0.38fF
C8900 a_2275_11190# col[6] 0.17fF
C8901 a_21950_11166# vcm 0.18fF
C8902 a_18026_1126# VDD 5.11fF
C8903 a_4974_16186# row_n[14] 0.43fF
C8904 a_8990_17190# m2_9188_17438# 0.19fF
C8905 a_22042_15182# ctop 4.91fF
C8906 a_15014_6146# row_n[4] 0.43fF
C8907 a_2475_10186# col[26] 0.22fF
C8908 a_14922_10162# rowon_n[8] 0.14fF
C8909 a_2275_13198# a_14314_13214# 0.15fF
C8910 a_2475_13198# a_16930_13174# 0.41fF
C8911 a_12306_1166# col_n[9] 0.11fF
C8912 a_22346_13214# col_n[19] 0.11fF
C8913 m2_5748_946# vcm 0.71fF
C8914 a_2275_1150# a_29070_1126# 0.14fF
C8915 a_2966_12170# rowon_n[10] 0.45fF
C8916 a_33086_5142# VDD 1.34fF
C8917 a_27062_6146# a_28066_6146# 0.86fF
C8918 a_28066_13174# m2_28264_13422# 0.19fF
C8919 a_2275_10186# a_7894_10162# 0.17fF
C8920 m2_2736_946# col_n[0] 0.45fF
C8921 a_2475_15206# a_31990_15182# 0.41fF
C8922 a_2275_15206# a_29374_15222# 0.15fF
C8923 a_16930_15182# a_17022_15182# 0.45fF
C8924 a_2275_13198# col[23] 0.17fF
C8925 a_2475_4162# rowon_n[2] 0.40fF
C8926 a_16018_11166# col[13] 0.38fF
C8927 a_17934_18194# vcm 0.18fF
C8928 a_2275_2154# col[28] 0.17fF
C8929 a_14010_8154# VDD 3.30fF
C8930 a_18026_8154# a_18026_7150# 0.84fF
C8931 a_2966_17190# VDD 4.45fF
C8932 a_2275_12194# a_22954_12170# 0.17fF
C8933 a_31078_7150# col_n[28] 0.34fF
C8934 a_20034_3134# vcm 0.89fF
C8935 a_11302_11206# col_n[8] 0.11fF
C8936 a_19030_11166# m2_19228_11414# 0.19fF
C8937 a_13006_13174# row_n[11] 0.43fF
C8938 a_29070_12170# VDD 1.75fF
C8939 m3_14916_18146# m3_15920_18146# 0.21fF
C8940 a_7986_9158# a_8990_9158# 0.86fF
C8941 a_12914_17190# rowon_n[15] 0.14fF
C8942 a_2475_9182# a_15014_9158# 0.68fF
C8943 a_8990_3134# rowoff_n[1] 2.33fF
C8944 a_23046_3134# row_n[1] 0.43fF
C8945 a_22954_7150# rowon_n[5] 0.14fF
C8946 a_35094_7150# vcm 0.15fF
C8947 a_29982_14178# rowoff_n[12] 0.43fF
C8948 a_26970_2130# a_27062_2130# 0.45fF
C8949 col_n[18] rowoff_n[8] 0.21fF
C8950 col_n[11] rowoff_n[1] 0.26fF
C8951 col_n[14] rowoff_n[4] 0.24fF
C8952 col_n[17] rowoff_n[7] 0.21fF
C8953 col_n[12] rowoff_n[2] 0.25fF
C8954 col_n[15] rowoff_n[5] 0.23fF
C8955 col_n[19] rowoff_n[9] 0.20fF
C8956 col_n[16] rowoff_n[6] 0.22fF
C8957 col_n[13] rowoff_n[3] 0.24fF
C8958 col_n[10] rowoff_n[0] 0.27fF
C8959 a_2475_6170# col[3] 0.22fF
C8960 a_2275_6170# a_5978_6146# 0.71fF
C8961 a_4974_9158# col[2] 0.38fF
C8962 a_9994_15182# VDD 3.71fF
C8963 a_33086_12170# a_33086_11166# 0.84fF
C8964 a_2475_11190# a_30074_11166# 0.68fF
C8965 a_25358_1166# vcm 0.25fF
C8966 a_2275_12194# col_n[10] 0.17fF
C8967 a_20034_5142# col_n[17] 0.34fF
C8968 a_16018_10162# vcm 0.89fF
C8969 a_30074_17190# col_n[27] 0.34fF
C8970 a_2275_1150# col_n[15] 0.14fF
C8971 a_9994_9158# m2_10192_9406# 0.19fF
C8972 m2_22816_946# col[20] 0.51fF
C8973 a_35398_10202# VDD 0.12fF
C8974 a_2275_8178# a_21038_8154# 0.71fF
C8975 a_2275_9182# col[0] 0.16fF
C8976 a_23046_13174# a_24050_13174# 0.86fF
C8977 col[20] rowoff_n[14] 0.21fF
C8978 a_6282_4178# vcm 0.24fF
C8979 col_n[3] rowoff_n[10] 0.32fF
C8980 a_29070_5142# m2_29268_5390# 0.19fF
C8981 a_31078_14178# vcm 0.89fF
C8982 a_27974_4138# VDD 0.29fF
C8983 a_2275_5166# a_11302_5182# 0.15fF
C8984 a_2475_5166# a_13918_5142# 0.41fF
C8985 a_7894_5142# a_7986_5142# 0.45fF
C8986 a_2475_8178# col[20] 0.22fF
C8987 a_2275_18218# a_9902_18194# 0.17fF
C8988 a_21038_10162# row_n[8] 0.43fF
C8989 a_10906_9158# rowoff_n[7] 0.65fF
C8990 a_20946_14178# rowon_n[12] 0.14fF
C8991 a_14010_15182# a_14010_14178# 0.84fF
C8992 a_21342_8194# vcm 0.24fF
C8993 a_2275_14202# col_n[27] 0.17fF
C8994 a_17934_15182# rowoff_n[13] 0.57fF
C8995 a_30986_4138# rowon_n[2] 0.14fF
C8996 a_2275_2154# a_4882_2130# 0.17fF
C8997 a_8990_3134# col_n[6] 0.34fF
C8998 a_34090_3134# ctop 4.80fF
C8999 a_12002_17190# vcm 0.89fF
C9000 a_19030_15182# col_n[16] 0.34fF
C9001 a_8898_7150# VDD 0.29fF
C9002 a_19942_7150# rowoff_n[5] 0.55fF
C9003 a_2275_7174# a_26362_7190# 0.15fF
C9004 a_2475_7174# a_28978_7150# 0.41fF
C9005 vcm col_n[17] 3.19fF
C9006 VDD col_n[20] 11.48fF
C9007 col[4] rowoff_n[15] 0.32fF
C9008 a_2275_11190# col[17] 0.17fF
C9009 a_14922_2130# vcm 0.18fF
C9010 a_2475_16210# a_6982_16186# 0.68fF
C9011 a_3970_16186# a_4974_16186# 0.86fF
C9012 a_20034_3134# m2_20232_3382# 0.19fF
C9013 a_28978_5142# rowoff_n[3] 0.44fF
C9014 a_3878_11166# vcm 0.18fF
C9015 a_7986_8154# rowon_n[6] 0.45fF
C9016 a_2275_4162# a_19942_4138# 0.17fF
C9017 a_15014_6146# ctop 4.91fF
C9018 a_23958_11166# VDD 0.29fF
C9019 m3_4876_1078# m3_5880_1078# 0.21fF
C9020 a_29070_2130# col[26] 0.38fF
C9021 a_22954_9158# a_23046_9158# 0.45fF
C9022 m2_1732_5966# sample_n 0.12fF
C9023 a_29982_6146# vcm 0.18fF
C9024 a_17326_15222# vcm 0.24fF
C9025 a_2475_18218# a_22954_18194# 0.41fF
C9026 m2_9764_946# VDD 6.25fF
C9027 a_2275_6170# a_35002_6146# 0.17fF
C9028 a_24354_2170# col_n[21] 0.11fF
C9029 a_19030_17190# row_n[15] 0.43fF
C9030 a_30074_10162# ctop 4.91fF
C9031 a_4882_14178# VDD 0.29fF
C9032 a_7986_13174# col_n[5] 0.34fF
C9033 a_29070_7150# row_n[5] 0.43fF
C9034 a_2275_15206# a_13006_15182# 0.71fF
C9035 a_28978_11166# rowon_n[9] 0.14fF
C9036 a_10906_9158# vcm 0.18fF
C9037 a_5886_16186# rowoff_n[14] 0.70fF
C9038 a_2475_3158# a_27062_3134# 0.68fF
C9039 a_14010_3134# a_15014_3134# 0.86fF
C9040 a_10998_13174# ctop 4.91fF
C9041 a_2275_10186# col_n[4] 0.17fF
C9042 a_19942_18194# VDD 0.50fF
C9043 a_2275_12194# a_3270_12210# 0.15fF
C9044 a_2475_12194# a_5886_12170# 0.41fF
C9045 a_28066_12170# col[25] 0.38fF
C9046 a_1957_3158# vcm 0.16fF
C9047 a_30074_11166# rowoff_n[9] 1.30fF
C9048 a_2275_17214# a_28066_17190# 0.71fF
C9049 a_5978_15182# rowon_n[13] 0.45fF
C9050 m2_19804_18014# m2_20232_18442# 0.19fF
C9051 a_25966_13174# vcm 0.18fF
C9052 a_22042_3134# VDD 2.47fF
C9053 a_4974_5142# a_4974_4138# 0.84fF
C9054 a_2275_7174# ctop 0.14fF
C9055 a_16018_5142# rowon_n[3] 0.45fF
C9056 a_26058_17190# ctop 4.93fF
C9057 a_23350_12210# col_n[20] 0.11fF
C9058 a_2275_14202# a_18330_14218# 0.15fF
C9059 a_2475_14202# a_20946_14178# 0.41fF
C9060 a_2475_17214# col[9] 0.22fF
C9061 col_n[23] rowoff_n[2] 0.17fF
C9062 col_n[26] rowoff_n[5] 0.15fF
C9063 col_n[29] rowoff_n[8] 0.13fF
C9064 col_n[22] rowoff_n[1] 0.18fF
C9065 col_n[27] rowoff_n[6] 0.14fF
C9066 col_n[30] rowoff_n[9] 0.12fF
C9067 col_n[24] rowoff_n[3] 0.16fF
C9068 col_n[21] rowoff_n[0] 0.19fF
C9069 col_n[28] rowoff_n[7] 0.14fF
C9070 col_n[25] rowoff_n[4] 0.16fF
C9071 a_2475_6170# col[14] 0.22fF
C9072 a_2275_2154# a_33086_2130# 0.71fF
C9073 a_6890_16186# vcm 0.18fF
C9074 a_2874_6146# VDD 0.29fF
C9075 a_29070_7150# a_30074_7150# 0.86fF
C9076 a_2275_11190# a_11910_11166# 0.17fF
C9077 a_27062_14178# row_n[12] 0.43fF
C9078 a_2275_12194# col_n[21] 0.17fF
C9079 a_8990_1126# vcm 0.15fF
C9080 a_2275_1150# col_n[26] 0.17fF
C9081 a_2275_16210# a_33390_16226# 0.15fF
C9082 a_18938_16186# a_19030_16186# 0.45fF
C9083 a_17022_10162# col[14] 0.38fF
C9084 a_18026_10162# VDD 2.89fF
C9085 a_2275_9182# col[11] 0.17fF
C9086 a_20034_9158# a_20034_8154# 0.84fF
C9087 a_2475_8178# a_3970_8154# 0.68fF
C9088 a_2275_8178# a_2966_8154# 0.67fF
C9089 col[31] rowoff_n[14] 0.14fF
C9090 a_32082_6146# col_n[29] 0.34fF
C9091 a_2275_13198# a_26970_13174# 0.17fF
C9092 col_n[14] rowoff_n[10] 0.24fF
C9093 a_24050_5142# vcm 0.89fF
C9094 a_18026_12170# rowoff_n[10] 1.89fF
C9095 m2_28840_946# vcm 0.71fF
C9096 a_12306_10202# col_n[9] 0.11fF
C9097 a_2275_18218# m2_25828_18014# 0.51fF
C9098 a_2475_8178# col[31] 0.22fF
C9099 a_14010_12170# rowon_n[10] 0.45fF
C9100 a_33086_14178# VDD 1.34fF
C9101 a_9994_10162# a_10998_10162# 0.86fF
C9102 a_2475_10186# a_19030_10162# 0.68fF
C9103 a_2966_10162# row_n[8] 0.41fF
C9104 a_24050_2130# rowon_n[0] 0.45fF
C9105 a_9994_2130# rowoff_n[0] 2.28fF
C9106 a_2275_14202# rowon_n[12] 1.99fF
C9107 a_4974_8154# vcm 0.89fF
C9108 a_34090_16186# rowoff_n[14] 1.10fF
C9109 a_28978_3134# a_29070_3134# 0.45fF
C9110 VDD col_n[31] 8.61fF
C9111 vcm col_n[28] 3.22fF
C9112 col[15] rowoff_n[15] 0.25fF
C9113 a_5978_8154# col[3] 0.38fF
C9114 a_2275_7174# a_9994_7150# 0.71fF
C9115 a_2475_15206# m2_34864_15002# 0.56fF
C9116 a_2275_11190# col[28] 0.17fF
C9117 a_2475_2154# row_n[0] 0.48fF
C9118 a_14010_17190# VDD 3.30fF
C9119 sample rowoff_n[11] 0.22fF
C9120 a_2475_12194# a_34090_12170# 0.68fF
C9121 a_21038_4138# col_n[18] 0.34fF
C9122 a_29374_3174# vcm 0.24fF
C9123 a_31078_16186# col_n[28] 0.34fF
C9124 a_35002_15182# rowon_n[13] 0.14fF
C9125 a_20034_12170# vcm 0.89fF
C9126 a_16930_2130# VDD 0.29fF
C9127 m3_1864_17142# m3_1864_16138# 0.20fF
C9128 a_2275_9182# a_25054_9158# 0.71fF
C9129 a_25054_14178# a_26058_14178# 0.86fF
C9130 a_2161_10186# rowoff_n[8] 0.14fF
C9131 a_10298_6186# vcm 0.24fF
C9132 a_5978_13174# rowoff_n[11] 2.47fF
C9133 m2_1732_2954# VDD 5.46fF
C9134 a_35094_16186# vcm 0.15fF
C9135 a_31990_6146# VDD 0.29fF
C9136 a_9902_6146# a_9994_6146# 0.45fF
C9137 a_34090_14178# m2_34288_14426# 0.19fF
C9138 a_2275_6170# a_15318_6186# 0.15fF
C9139 a_2475_6170# a_17934_6146# 0.41fF
C9140 a_22042_9158# rowon_n[7] 0.45fF
C9141 a_2475_15206# col[3] 0.22fF
C9142 a_11910_8154# rowoff_n[6] 0.64fF
C9143 a_2475_4162# col[8] 0.22fF
C9144 a_16018_16186# a_16018_15182# 0.84fF
C9145 a_9994_2130# col_n[7] 0.34fF
C9146 a_25358_10202# vcm 0.24fF
C9147 a_22042_17190# rowoff_n[15] 1.69fF
C9148 a_20034_14178# col_n[17] 0.34fF
C9149 a_2275_3158# a_8898_3134# 0.17fF
C9150 a_20946_6146# rowoff_n[4] 0.54fF
C9151 a_3970_4138# ctop 4.91fF
C9152 a_2275_10186# col_n[15] 0.17fF
C9153 m3_1864_13126# ctop 0.22fF
C9154 a_12914_9158# VDD 0.29fF
C9155 a_5978_16186# m2_6176_16434# 0.19fF
C9156 a_2275_8178# a_30378_8194# 0.15fF
C9157 a_2475_8178# a_32994_8154# 0.41fF
C9158 a_18938_4138# vcm 0.18fF
C9159 a_9902_3134# rowon_n[1] 0.14fF
C9160 a_29982_4138# rowoff_n[2] 0.43fF
C9161 a_2475_17214# a_10998_17190# 0.68fF
C9162 a_5978_17190# a_6982_17190# 0.86fF
C9163 m2_1732_18014# sample 0.32fF
C9164 a_2966_4138# m2_3164_4386# 0.19fF
C9165 a_2275_7174# col[5] 0.17fF
C9166 m2_1732_18014# m2_2736_18014# 0.86fF
C9167 a_6282_13214# vcm 0.24fF
C9168 a_34394_3174# col_n[31] 0.11fF
C9169 a_25054_12170# m2_25252_12418# 0.19fF
C9170 a_2275_5166# a_23958_5142# 0.17fF
C9171 m2_3740_18014# col[1] 0.37fF
C9172 a_19030_8154# ctop 4.91fF
C9173 a_27974_13174# VDD 0.29fF
C9174 a_24962_10162# a_25054_10162# 0.45fF
C9175 a_2475_17214# col[20] 0.22fF
C9176 a_2475_6170# col[25] 0.22fF
C9177 a_1957_14202# a_2161_14202# 0.11fF
C9178 a_2475_14202# a_2275_14202# 2.96fF
C9179 m2_1732_7974# m2_2160_8402# 0.19fF
C9180 a_33998_8154# vcm 0.18fF
C9181 a_26058_3134# a_26058_2130# 0.84fF
C9182 a_2475_2154# a_16018_2130# 0.68fF
C9183 a_21342_17230# vcm 0.24fF
C9184 a_25358_1166# col_n[22] 0.11fF
C9185 m2_32856_18014# m3_32988_18146# 4.41fF
C9186 a_20034_16186# rowon_n[14] 0.45fF
C9187 a_8990_12170# col_n[6] 0.34fF
C9188 a_34090_12170# ctop 4.80fF
C9189 a_8898_16186# VDD 0.29fF
C9190 a_30074_6146# rowon_n[4] 0.45fF
C9191 a_2275_16210# a_17022_16186# 0.71fF
C9192 a_14922_11166# vcm 0.18fF
C9193 a_10998_1126# VDD 0.13fF
C9194 a_2275_9182# col[22] 0.17fF
C9195 a_16018_4138# a_17022_4138# 0.86fF
C9196 a_16018_10162# m2_16216_10410# 0.19fF
C9197 a_2475_4162# a_31078_4138# 0.68fF
C9198 col_n[25] rowoff_n[10] 0.16fF
C9199 a_15014_15182# ctop 4.91fF
C9200 a_7986_6146# row_n[4] 0.43fF
C9201 a_2275_13198# a_7286_13214# 0.15fF
C9202 a_2475_13198# a_9902_13174# 0.41fF
C9203 a_5886_13174# a_5978_13174# 0.45fF
C9204 a_29070_11166# col[26] 0.38fF
C9205 a_7894_10162# rowon_n[8] 0.14fF
C9206 a_31078_10162# rowoff_n[8] 1.25fF
C9207 m2_19804_18014# col_n[17] 0.33fF
C9208 a_35002_13174# rowoff_n[11] 0.38fF
C9209 a_2275_1150# a_22042_1126# 0.14fF
C9210 a_29982_15182# vcm 0.18fF
C9211 a_26058_5142# VDD 2.06fF
C9212 m2_32856_946# VDD 2.81fF
C9213 a_6982_6146# a_6982_5142# 0.84fF
C9214 a_24354_11206# col_n[21] 0.11fF
C9215 a_2475_15206# a_24962_15182# 0.41fF
C9216 a_2275_15206# a_22346_15222# 0.15fF
C9217 m2_34864_11990# m2_34864_10986# 0.84fF
C9218 VDD rowon_n[10] 4.61fF
C9219 sample row_n[11] 0.92fF
C9220 col_n[7] rowon_n[15] 0.17fF
C9221 col_n[1] rowon_n[12] 0.17fF
C9222 col_n[5] rowon_n[14] 0.17fF
C9223 col_n[3] rowon_n[13] 0.17fF
C9224 vcm row_n[12] 1.08fF
C9225 col_n[2] row_n[13] 0.37fF
C9226 col_n[4] row_n[14] 0.37fF
C9227 col_n[6] row_n[15] 0.37fF
C9228 col_n[0] rowon_n[11] 0.17fF
C9229 col[26] rowoff_n[15] 0.17fF
C9230 a_6982_8154# m2_7180_8402# 0.19fF
C9231 a_10906_18194# vcm 0.18fF
C9232 a_2475_2154# col[2] 0.22fF
C9233 a_20034_1126# m2_20232_1374# 0.19fF
C9234 a_6982_8154# VDD 4.02fF
C9235 col_n[9] rowoff_n[11] 0.27fF
C9236 a_31078_8154# a_32082_8154# 0.86fF
C9237 a_28066_13174# rowon_n[11] 0.45fF
C9238 a_2275_12194# a_15926_12170# 0.17fF
C9239 a_13006_3134# vcm 0.89fF
C9240 a_20946_17190# a_21038_17190# 0.45fF
C9241 a_2275_8178# col_n[9] 0.17fF
C9242 a_18026_9158# col[15] 0.38fF
C9243 a_26058_4138# m2_26256_4386# 0.19fF
C9244 a_1957_12194# vcm 0.16fF
C9245 a_5978_13174# row_n[11] 0.43fF
C9246 a_22042_12170# VDD 2.47fF
C9247 a_33086_5142# col_n[30] 0.34fF
C9248 a_5886_17190# rowon_n[15] 0.14fF
C9249 a_22042_10162# a_22042_9158# 0.84fF
C9250 a_2475_9182# a_7986_9158# 0.68fF
C9251 a_2275_16210# ctop 0.14fF
C9252 a_2275_14202# a_30986_14178# 0.17fF
C9253 a_2475_3158# rowoff_n[1] 4.75fF
C9254 a_16018_3134# row_n[1] 0.43fF
C9255 a_13310_9198# col_n[10] 0.11fF
C9256 a_15926_7150# rowon_n[5] 0.14fF
C9257 a_28066_7150# vcm 0.89fF
C9258 a_22954_14178# rowoff_n[12] 0.51fF
C9259 a_2475_15206# col[14] 0.22fF
C9260 a_2475_4162# col[19] 0.22fF
C9261 a_2874_15182# VDD 0.29fF
C9262 a_12002_11166# a_13006_11166# 0.86fF
C9263 a_2475_11190# a_23046_11166# 0.68fF
C9264 a_18330_1166# vcm 0.24fF
C9265 a_2275_10186# col_n[26] 0.17fF
C9266 a_8990_10162# vcm 0.89fF
C9267 a_6982_7150# col[4] 0.38fF
C9268 a_30986_4138# a_31078_4138# 0.45fF
C9269 a_2275_6170# rowoff_n[4] 0.81fF
C9270 a_2275_8178# a_14010_8154# 0.71fF
C9271 a_22042_3134# col_n[19] 0.34fF
C9272 a_2275_7174# col[16] 0.17fF
C9273 a_32082_15182# col_n[29] 0.34fF
C9274 a_33390_5182# vcm 0.24fF
C9275 a_24050_14178# vcm 0.89fF
C9276 a_20946_4138# VDD 0.29fF
C9277 a_2275_5166# a_4274_5182# 0.15fF
C9278 a_2475_5166# a_6890_5142# 0.41fF
C9279 a_2475_17214# col[31] 0.22fF
C9280 a_2275_10186# a_29070_10162# 0.71fF
C9281 a_14010_10162# row_n[8] 0.43fF
C9282 a_13918_14178# rowon_n[12] 0.14fF
C9283 a_27062_15182# a_28066_15182# 0.86fF
C9284 a_14314_8194# vcm 0.24fF
C9285 a_10906_15182# rowoff_n[13] 0.65fF
C9286 a_2275_12194# row_n[10] 26.41fF
C9287 a_23958_4138# rowon_n[2] 0.14fF
C9288 m2_6752_946# col[4] 0.51fF
C9289 a_4974_17190# vcm 0.89fF
C9290 a_27062_3134# ctop 4.91fF
C9291 a_12914_7150# rowoff_n[5] 0.63fF
C9292 a_11910_7150# a_12002_7150# 0.45fF
C9293 a_2275_7174# a_19334_7190# 0.15fF
C9294 a_2475_7174# a_21950_7150# 0.41fF
C9295 a_5978_17190# col[3] 0.38fF
C9296 a_7894_2130# vcm 0.18fF
C9297 a_18026_17190# a_18026_16186# 0.84fF
C9298 a_21038_13174# col_n[18] 0.34fF
C9299 a_21950_5142# rowoff_n[3] 0.52fF
C9300 a_29374_12210# vcm 0.24fF
C9301 a_2275_4162# a_12914_4138# 0.17fF
C9302 a_2475_10186# m2_1732_9982# 0.16fF
C9303 a_7986_6146# ctop 4.91fF
C9304 a_16930_11166# VDD 0.29fF
C9305 a_2275_9182# a_35398_9198# 0.15fF
C9306 a_34090_17190# rowon_n[15] 0.45fF
C9307 a_2275_6170# col_n[3] 0.17fF
C9308 m2_1732_3958# vcm 1.11fF
C9309 a_30986_3134# rowoff_n[1] 0.42fF
C9310 a_22954_6146# vcm 0.18fF
C9311 a_10298_15222# vcm 0.24fF
C9312 a_2475_18218# a_15926_18194# 0.41fF
C9313 a_2275_6170# a_27974_6146# 0.17fF
C9314 a_12002_17190# row_n[15] 0.43fF
C9315 a_23046_10162# ctop 4.91fF
C9316 a_31990_15182# VDD 0.29fF
C9317 a_26970_11166# a_27062_11166# 0.45fF
C9318 col_n[12] rowon_n[12] 0.17fF
C9319 col_n[1] row_n[7] 0.37fF
C9320 col_n[0] row_n[6] 0.37fF
C9321 col_n[8] rowon_n[10] 0.17fF
C9322 vcm rowon_n[6] 0.91fF
C9323 col_n[6] rowon_n[9] 0.17fF
C9324 sample rowon_n[5] 0.10fF
C9325 col_n[4] rowon_n[8] 0.17fF
C9326 col_n[11] row_n[12] 0.37fF
C9327 col_n[10] rowon_n[11] 0.17fF
C9328 col_n[15] row_n[14] 0.37fF
C9329 VDD row_n[5] 4.64fF
C9330 col_n[13] row_n[13] 0.37fF
C9331 col_n[17] row_n[15] 0.37fF
C9332 col_n[9] row_n[11] 0.37fF
C9333 col_n[3] row_n[8] 0.37fF
C9334 col_n[14] rowon_n[13] 0.17fF
C9335 col_n[5] row_n[9] 0.37fF
C9336 col_n[16] rowon_n[14] 0.17fF
C9337 col_n[7] row_n[10] 0.37fF
C9338 col_n[18] rowon_n[15] 0.17fF
C9339 col_n[2] rowon_n[7] 0.17fF
C9340 m2_27836_18014# vcm 0.71fF
C9341 a_22042_7150# row_n[5] 0.43fF
C9342 a_2275_15206# a_5978_15182# 0.71fF
C9343 a_2475_13198# col[8] 0.22fF
C9344 a_21950_11166# rowon_n[9] 0.14fF
C9345 a_2475_2154# col[13] 0.22fF
C9346 col_n[20] rowoff_n[11] 0.19fF
C9347 a_28066_4138# a_28066_3134# 0.84fF
C9348 a_2475_3158# a_20034_3134# 0.68fF
C9349 a_9994_11166# col_n[7] 0.34fF
C9350 a_2475_1150# m2_20808_946# 0.62fF
C9351 a_31078_2130# m2_30848_946# 0.84fF
C9352 m3_19936_1078# ctop 0.34fF
C9353 a_3970_13174# ctop 4.91fF
C9354 a_12914_18194# VDD 0.50fF
C9355 a_2275_8178# col_n[20] 0.17fF
C9356 a_23046_11166# rowoff_n[9] 1.64fF
C9357 a_2275_17214# a_21038_17190# 0.71fF
C9358 m2_12776_18014# m2_13204_18442# 0.19fF
C9359 a_18938_13174# vcm 0.18fF
C9360 a_15014_3134# VDD 3.20fF
C9361 a_18026_5142# a_19030_5142# 0.86fF
C9362 a_2275_16210# col[5] 0.17fF
C9363 a_8990_5142# rowon_n[3] 0.45fF
C9364 a_2275_5166# col[10] 0.17fF
C9365 a_2275_18218# a_31078_18194# 0.14fF
C9366 m2_15788_946# m2_16792_946# 0.86fF
C9367 a_34394_12210# col_n[31] 0.11fF
C9368 a_30074_10162# col[27] 0.38fF
C9369 a_19030_17190# ctop 4.93fF
C9370 a_32082_9158# rowoff_n[7] 1.20fF
C9371 a_2275_14202# a_11302_14218# 0.15fF
C9372 a_2475_14202# a_13918_14178# 0.41fF
C9373 a_7894_14178# a_7986_14178# 0.45fF
C9374 col_n[4] rowoff_n[12] 0.31fF
C9375 a_2475_15206# col[25] 0.22fF
C9376 a_2475_4162# col[30] 0.22fF
C9377 a_2275_2154# a_26058_2130# 0.71fF
C9378 a_33998_17190# vcm 0.18fF
C9379 a_30074_7150# VDD 1.65fF
C9380 a_8990_7150# a_8990_6146# 0.84fF
C9381 a_25358_10202# col_n[22] 0.11fF
C9382 a_20034_14178# row_n[12] 0.43fF
C9383 a_2966_11166# a_3970_11166# 0.86fF
C9384 a_2275_11190# a_4882_11166# 0.17fF
C9385 a_2475_1150# vcm 1.28fF
C9386 a_2475_16210# a_28978_16186# 0.41fF
C9387 a_2275_16210# a_26362_16226# 0.15fF
C9388 a_2275_2154# m2_2736_1950# 0.48fF
C9389 a_30074_4138# row_n[2] 0.43fF
C9390 a_29982_8154# rowon_n[6] 0.14fF
C9391 a_10998_10162# VDD 3.61fF
C9392 a_33086_9158# a_34090_9158# 0.86fF
C9393 a_12002_17190# m2_12200_17438# 0.19fF
C9394 a_2275_7174# col[27] 0.17fF
C9395 a_2275_13198# a_19942_13174# 0.17fF
C9396 a_19030_8154# col[16] 0.38fF
C9397 a_17022_5142# vcm 0.89fF
C9398 a_10998_12170# rowoff_n[10] 2.23fF
C9399 a_22954_18194# a_23046_18194# 0.11fF
C9400 a_2275_18218# m2_11772_18014# 0.51fF
C9401 row_n[3] rowoff_n[3] 0.64fF
C9402 a_2475_1150# a_35002_1126# 0.41fF
C9403 a_2275_1150# a_31382_1166# 0.15fF
C9404 a_17934_1126# a_18026_1126# 0.48fF
C9405 a_2275_5166# m2_34864_4962# 0.51fF
C9406 a_2275_4162# VDD 3.18fF
C9407 a_6982_12170# rowon_n[10] 0.45fF
C9408 a_34090_4138# col_n[31] 0.34fF
C9409 a_31078_13174# m2_31276_13422# 0.19fF
C9410 a_26058_14178# VDD 2.06fF
C9411 a_2475_10186# a_12002_10162# 0.68fF
C9412 a_24050_11166# a_24050_10162# 0.84fF
C9413 m2_34864_2954# rowoff_n[1] 1.02fF
C9414 a_17022_2130# rowon_n[0] 0.45fF
C9415 a_2874_2130# rowoff_n[0] 0.74fF
C9416 a_14314_8194# col_n[11] 0.11fF
C9417 a_2275_15206# a_35002_15182# 0.17fF
C9418 a_32082_9158# vcm 0.89fF
C9419 a_27062_16186# rowoff_n[14] 1.45fF
C9420 a_2275_7174# a_2874_7150# 0.17fF
C9421 a_2475_7174# a_3878_7150# 0.41fF
C9422 a_2475_11190# col[2] 0.22fF
C9423 a_6982_17190# VDD 4.03fF
C9424 a_2475_12194# a_27062_12170# 0.68fF
C9425 a_14010_12170# a_15014_12170# 0.86fF
C9426 a_28066_11166# row_n[9] 0.43fF
C9427 a_22346_3174# vcm 0.24fF
C9428 a_27974_15182# rowon_n[13] 0.14fF
C9429 a_7986_6146# col[5] 0.38fF
C9430 a_35002_4138# m2_34864_3958# 0.33fF
C9431 a_3878_5142# rowoff_n[3] 0.73fF
C9432 a_13006_12170# vcm 0.89fF
C9433 a_9902_2130# VDD 0.29fF
C9434 a_2275_17214# col_n[9] 0.17fF
C9435 a_22042_11166# m2_22240_11414# 0.19fF
C9436 a_32994_5142# a_33086_5142# 0.45fF
C9437 a_2275_6170# col_n[14] 0.17fF
C9438 a_23046_2130# col_n[20] 0.34fF
C9439 a_13918_18194# m2_13780_18014# 0.34fF
C9440 a_2275_9182# a_18026_9158# 0.71fF
C9441 a_33086_14178# col_n[30] 0.34fF
C9442 a_4974_14178# a_4974_13174# 0.84fF
C9443 a_3270_6186# vcm 0.24fF
C9444 a_13310_18234# col_n[10] 0.11fF
C9445 a_2275_3158# col[4] 0.17fF
C9446 a_28066_16186# vcm 0.89fF
C9447 a_24962_6146# VDD 0.29fF
C9448 a_2275_6170# a_8290_6186# 0.15fF
C9449 a_2475_6170# a_10906_6146# 0.41fF
C9450 col_n[3] rowon_n[2] 0.17fF
C9451 col_n[28] row_n[15] 0.37fF
C9452 col_n[10] row_n[6] 0.37fF
C9453 col_n[26] row_n[14] 0.37fF
C9454 col_n[8] row_n[5] 0.37fF
C9455 col_n[24] row_n[13] 0.37fF
C9456 vcm row_n[1] 1.08fF
C9457 col_n[6] row_n[4] 0.37fF
C9458 sample row_n[0] 0.89fF
C9459 col_n[4] row_n[3] 0.37fF
C9460 col_n[23] rowon_n[12] 0.17fF
C9461 col_n[2] row_n[2] 0.37fF
C9462 col_n[25] rowon_n[13] 0.17fF
C9463 col_n[7] rowon_n[4] 0.17fF
C9464 col_n[14] row_n[8] 0.37fF
C9465 col_n[20] row_n[11] 0.37fF
C9466 col_n[12] row_n[7] 0.37fF
C9467 col_n[5] rowon_n[3] 0.17fF
C9468 col_n[16] row_n[9] 0.37fF
C9469 col_n[9] rowon_n[5] 0.17fF
C9470 col_n[27] rowon_n[14] 0.17fF
C9471 col_n[18] row_n[10] 0.37fF
C9472 col_n[11] rowon_n[6] 0.17fF
C9473 col_n[29] rowon_n[15] 0.17fF
C9474 col_n[13] rowon_n[7] 0.17fF
C9475 col_n[21] rowon_n[11] 0.17fF
C9476 col_n[22] row_n[12] 0.37fF
C9477 VDD sw 0.56fF
C9478 col_n[15] rowon_n[8] 0.17fF
C9479 col_n[0] rowon_n[0] 0.17fF
C9480 col_n[1] rowon_n[1] 0.17fF
C9481 col_n[17] rowon_n[9] 0.17fF
C9482 col_n[19] rowon_n[10] 0.17fF
C9483 a_15014_9158# rowon_n[7] 0.45fF
C9484 a_4882_8154# rowoff_n[6] 0.72fF
C9485 a_2475_13198# col[19] 0.22fF
C9486 a_2275_11190# a_33086_11166# 0.71fF
C9487 a_2475_2154# col[24] 0.22fF
C9488 col_n[31] rowoff_n[11] 0.11fF
C9489 a_30986_1126# vcm 0.18fF
C9490 a_29070_16186# a_30074_16186# 0.86fF
C9491 a_3878_11166# rowon_n[9] 0.14fF
C9492 a_18330_10202# vcm 0.24fF
C9493 a_15014_17190# rowoff_n[15] 2.03fF
C9494 m2_31852_18014# VDD 2.32fF
C9495 a_13006_9158# m2_13204_9406# 0.19fF
C9496 a_13918_6146# rowoff_n[4] 0.61fF
C9497 a_31078_5142# ctop 4.91fF
C9498 a_5886_9158# VDD 0.29fF
C9499 m3_15920_18146# ctop 0.21fF
C9500 a_2275_8178# col_n[31] 0.17fF
C9501 a_6982_16186# col[4] 0.38fF
C9502 a_13918_8154# a_14010_8154# 0.45fF
C9503 a_2475_8178# a_25966_8154# 0.41fF
C9504 a_2275_8178# a_23350_8194# 0.15fF
C9505 a_22042_12170# col_n[19] 0.34fF
C9506 a_11910_4138# vcm 0.18fF
C9507 a_2475_17214# a_3970_17190# 0.68fF
C9508 a_2275_17214# a_2966_17190# 0.67fF
C9509 a_22954_4138# rowoff_n[2] 0.51fF
C9510 a_2275_16210# col[16] 0.17fF
C9511 a_32082_5142# m2_32280_5390# 0.19fF
C9512 a_33390_14218# vcm 0.24fF
C9513 a_2275_5166# col[21] 0.17fF
C9514 a_2275_5166# a_16930_5142# 0.17fF
C9515 a_12002_8154# ctop 4.91fF
C9516 a_20946_13174# VDD 0.29fF
C9517 a_31990_2130# rowoff_n[0] 0.41fF
C9518 col_n[15] rowoff_n[12] 0.23fF
C9519 a_26970_8154# vcm 0.18fF
C9520 a_4974_2130# a_5978_2130# 0.86fF
C9521 a_2475_2154# a_8990_2130# 0.68fF
C9522 a_3970_7150# m2_4168_7398# 0.19fF
C9523 a_14314_17230# vcm 0.24fF
C9524 a_13006_16186# rowon_n[14] 0.45fF
C9525 a_2275_7174# a_31990_7150# 0.17fF
C9526 a_27062_12170# ctop 4.91fF
C9527 a_1957_14202# row_n[12] 0.29fF
C9528 a_28978_12170# a_29070_12170# 0.45fF
C9529 a_23046_6146# rowon_n[4] 0.45fF
C9530 a_2275_16210# a_9994_16186# 0.71fF
C9531 a_23046_3134# m2_23244_3382# 0.19fF
C9532 a_7894_11166# vcm 0.18fF
C9533 a_10998_10162# col_n[8] 0.34fF
C9534 a_3970_1126# VDD 7.24fF
C9535 a_30074_5142# a_30074_4138# 0.84fF
C9536 a_2475_4162# a_24050_4138# 0.68fF
C9537 col_n[0] rowoff_n[13] 0.34fF
C9538 a_32994_18194# m2_32856_18014# 0.34fF
C9539 a_9994_17190# m2_9764_18014# 0.84fF
C9540 a_7986_15182# ctop 4.91fF
C9541 a_24050_10162# rowoff_n[8] 1.59fF
C9542 ctop rowoff_n[1] 0.28fF
C9543 a_2275_15206# col_n[3] 0.17fF
C9544 col[2] rowoff_n[9] 0.33fF
C9545 col[1] rowoff_n[8] 0.34fF
C9546 col[0] rowoff_n[7] 0.34fF
C9547 a_34090_15182# row_n[13] 0.43fF
C9548 a_2275_4162# col_n[8] 0.17fF
C9549 a_27974_13174# rowoff_n[11] 0.46fF
C9550 a_2275_1150# a_15014_1126# 0.14fF
C9551 a_22954_15182# vcm 0.18fF
C9552 a_19030_5142# VDD 2.78fF
C9553 a_20034_6146# a_21038_6146# 0.86fF
C9554 a_31078_9158# col[28] 0.38fF
C9555 a_33086_8154# rowoff_n[6] 1.15fF
C9556 a_9902_15182# a_9994_15182# 0.45fF
C9557 a_2275_15206# a_15318_15222# 0.15fF
C9558 a_2475_15206# a_17934_15182# 0.41fF
C9559 m2_34864_15002# VDD 1.59fF
C9560 a_2275_3158# a_30074_3134# 0.71fF
C9561 a_2475_11190# col[13] 0.22fF
C9562 a_34090_9158# VDD 1.23fF
C9563 a_26362_9198# col_n[23] 0.11fF
C9564 a_10998_8154# a_10998_7150# 0.84fF
C9565 a_21038_13174# rowon_n[11] 0.45fF
C9566 a_2275_12194# a_8898_12170# 0.17fF
C9567 m2_34864_11990# row_n[10] 0.38fF
C9568 a_5978_3134# vcm 0.89fF
C9569 a_2275_17214# col_n[20] 0.17fF
C9570 a_31078_3134# rowon_n[1] 0.45fF
C9571 a_2475_17214# a_32994_17190# 0.41fF
C9572 a_2275_17214# a_30378_17230# 0.15fF
C9573 a_2275_6170# col_n[25] 0.17fF
C9574 a_2275_18218# col_n[5] 0.17fF
C9575 a_15014_12170# VDD 3.20fF
C9576 m2_32856_946# col_n[30] 0.54fF
C9577 a_20034_7150# col[17] 0.38fF
C9578 a_2275_14202# col[10] 0.17fF
C9579 a_2275_14202# a_23958_14178# 0.17fF
C9580 a_2275_3158# col[15] 0.17fF
C9581 a_8990_3134# row_n[1] 0.43fF
C9582 a_8898_7150# rowon_n[5] 0.14fF
C9583 a_21038_7150# vcm 0.89fF
C9584 a_15926_14178# rowoff_n[12] 0.59fF
C9585 a_19942_2130# a_20034_2130# 0.45fF
C9586 col_n[29] row_n[10] 0.37fF
C9587 col_n[20] rowon_n[5] 0.17fF
C9588 VDD col[3] 12.69fF
C9589 col_n[27] row_n[9] 0.37fF
C9590 col_n[18] rowon_n[4] 0.17fF
C9591 col_n[25] row_n[8] 0.37fF
C9592 col_n[31] row_n[11] 0.37fF
C9593 col_n[16] rowon_n[3] 0.17fF
C9594 col_n[23] row_n[7] 0.37fF
C9595 col_n[14] rowon_n[2] 0.17fF
C9596 col_n[21] row_n[6] 0.37fF
C9597 col_n[12] rowon_n[1] 0.17fF
C9598 col_n[19] row_n[5] 0.37fF
C9599 col_n[10] rowon_n[0] 0.17fF
C9600 vcm col[0] 6.58fF
C9601 col_n[24] rowon_n[7] 0.17fF
C9602 col_n[22] rowon_n[6] 0.17fF
C9603 col_n[26] rowon_n[8] 0.17fF
C9604 col_n[0] col[1] 6.24fF
C9605 col_n[28] rowon_n[9] 0.17fF
C9606 col_n[9] row_n[0] 0.37fF
C9607 col_n[30] rowon_n[10] 0.17fF
C9608 col_n[11] row_n[1] 0.37fF
C9609 col_n[13] row_n[2] 0.37fF
C9610 col_n[15] row_n[3] 0.37fF
C9611 col_n[17] row_n[4] 0.37fF
C9612 a_2475_13198# col[30] 0.22fF
C9613 a_30074_16186# VDD 1.65fF
C9614 a_15318_7190# col_n[12] 0.11fF
C9615 a_2475_11190# a_16018_11166# 0.68fF
C9616 a_26058_12170# a_26058_11166# 0.84fF
C9617 a_11302_1166# vcm 0.25fF
C9618 a_2475_10186# vcm 1.32fF
C9619 a_32994_1126# VDD 0.68fF
C9620 a_29070_17190# m2_28840_18014# 0.84fF
C9621 a_2275_8178# a_6982_8154# 0.71fF
C9622 a_2475_13198# a_31078_13174# 0.68fF
C9623 a_16018_13174# a_17022_13174# 0.86fF
C9624 a_29070_10162# rowon_n[8] 0.45fF
C9625 a_2275_16210# col[27] 0.17fF
C9626 a_8990_5142# col[6] 0.38fF
C9627 a_26362_5182# vcm 0.24fF
C9628 a_19030_17190# col[16] 0.38fF
C9629 a_17022_14178# vcm 0.89fF
C9630 a_13918_4138# VDD 0.29fF
C9631 a_35002_6146# a_35094_6146# 0.11fF
C9632 col_n[26] rowoff_n[12] 0.15fF
C9633 a_2275_13198# VDD 3.18fF
C9634 a_34090_13174# col_n[31] 0.34fF
C9635 a_2275_10186# a_22042_10162# 0.71fF
C9636 a_2275_2154# col_n[2] 0.17fF
C9637 a_6982_10162# row_n[8] 0.43fF
C9638 a_6890_14178# rowon_n[12] 0.14fF
C9639 a_4274_5182# col_n[1] 0.11fF
C9640 a_6982_15182# a_6982_14178# 0.84fF
C9641 a_14314_17230# col_n[11] 0.11fF
C9642 a_7286_8194# vcm 0.24fF
C9643 a_16930_4138# rowon_n[2] 0.14fF
C9644 a_20034_3134# ctop 4.91fF
C9645 a_32082_18194# vcm 0.15fF
C9646 a_28978_8154# VDD 0.29fF
C9647 a_5886_7150# rowoff_n[5] 0.70fF
C9648 a_2475_7174# a_14922_7150# 0.41fF
C9649 a_2275_7174# a_12306_7190# 0.15fF
C9650 a_35002_3134# vcm 0.18fF
C9651 a_31078_17190# a_32082_17190# 0.86fF
C9652 a_2475_9182# col[7] 0.22fF
C9653 a_14922_5142# rowoff_n[3] 0.60fF
C9654 a_22346_12210# vcm 0.24fF
C9655 col_n[10] rowoff_n[13] 0.27fF
C9656 a_2275_4162# a_5886_4138# 0.17fF
C9657 a_7986_15182# col[5] 0.38fF
C9658 a_9902_11166# VDD 0.29fF
C9659 a_2475_9182# a_29982_9158# 0.41fF
C9660 a_2275_9182# a_27366_9198# 0.15fF
C9661 a_27062_17190# rowon_n[15] 0.45fF
C9662 a_15926_9158# a_16018_9158# 0.45fF
C9663 a_2275_15206# col_n[14] 0.17fF
C9664 col[4] rowoff_n[0] 0.32fF
C9665 col[5] rowoff_n[1] 0.31fF
C9666 col[6] rowoff_n[2] 0.31fF
C9667 col[7] rowoff_n[3] 0.30fF
C9668 col[8] rowoff_n[4] 0.29fF
C9669 col[9] rowoff_n[5] 0.29fF
C9670 col[10] rowoff_n[6] 0.28fF
C9671 col[11] rowoff_n[7] 0.27fF
C9672 col[12] rowoff_n[8] 0.27fF
C9673 col[13] rowoff_n[9] 0.26fF
C9674 a_2275_4162# col_n[19] 0.17fF
C9675 a_23046_11166# col_n[20] 0.34fF
C9676 a_23958_3134# rowoff_n[1] 0.50fF
C9677 a_15926_6146# vcm 0.18fF
C9678 a_3270_15222# vcm 0.24fF
C9679 a_2475_18218# a_8898_18194# 0.41fF
C9680 a_35494_6508# VDD 0.13fF
C9681 a_2275_12194# col[4] 0.17fF
C9682 a_2275_6170# a_20946_6146# 0.17fF
C9683 a_4974_17190# row_n[15] 0.43fF
C9684 a_16018_10162# ctop 4.91fF
C9685 a_2275_1150# col[9] 0.17fF
C9686 a_24962_15182# VDD 0.29fF
C9687 m2_13780_18014# vcm 0.71fF
C9688 a_15014_7150# row_n[5] 0.43fF
C9689 a_14922_11166# rowon_n[9] 0.14fF
C9690 a_2475_11190# col[24] 0.22fF
C9691 a_30986_10162# vcm 0.18fF
C9692 a_6982_3134# a_7986_3134# 0.86fF
C9693 a_2475_3158# a_13006_3134# 0.68fF
C9694 m3_34996_6098# ctop 0.22fF
C9695 a_2275_8178# a_34394_8194# 0.15fF
C9696 a_8990_16186# m2_9188_16434# 0.19fF
C9697 a_2966_13174# rowon_n[11] 0.45fF
C9698 a_31078_14178# ctop 4.91fF
C9699 a_5886_18194# VDD 0.50fF
C9700 a_2275_17214# col_n[31] 0.17fF
C9701 a_30986_13174# a_31078_13174# 0.45fF
C9702 a_2275_18218# col_n[16] 0.17fF
C9703 a_2275_17214# a_14010_17190# 0.71fF
C9704 a_16018_11166# rowoff_n[9] 1.98fF
C9705 a_12002_9158# col_n[9] 0.34fF
C9706 m2_5748_18014# m2_6176_18442# 0.19fF
C9707 a_11910_13174# vcm 0.18fF
C9708 a_7986_3134# VDD 3.92fF
C9709 a_2475_5166# a_28066_5142# 0.68fF
C9710 a_32082_6146# a_32082_5142# 0.84fF
C9711 a_28066_12170# m2_28264_12418# 0.19fF
C9712 a_2275_14202# col[21] 0.17fF
C9713 a_2275_18218# a_24050_18194# 0.14fF
C9714 a_2475_5166# rowon_n[3] 0.40fF
C9715 m2_8760_946# m2_9764_946# 0.86fF
C9716 a_2275_3158# col[26] 0.17fF
C9717 a_12002_17190# ctop 4.93fF
C9718 a_25054_9158# rowoff_n[7] 1.54fF
C9719 a_2475_14202# a_6890_14178# 0.41fF
C9720 a_2275_14202# a_4274_14218# 0.15fF
C9721 col_n[5] col[6] 6.22fF
C9722 col_n[31] rowon_n[5] 0.17fF
C9723 col_n[29] rowon_n[4] 0.17fF
C9724 col_n[22] row_n[1] 0.37fF
C9725 col_n[20] row_n[0] 0.37fF
C9726 col_n[24] row_n[2] 0.37fF
C9727 col_n[26] row_n[3] 0.37fF
C9728 VDD col[14] 9.97fF
C9729 col_n[28] row_n[4] 0.37fF
C9730 col_n[21] rowon_n[0] 0.17fF
C9731 col_n[30] row_n[5] 0.37fF
C9732 col_n[23] rowon_n[1] 0.17fF
C9733 col_n[15] en_bit_n[1] 0.19fF
C9734 vcm col[11] 6.66fF
C9735 col_n[25] rowon_n[2] 0.17fF
C9736 col_n[27] rowon_n[3] 0.17fF
C9737 a_2966_7150# vcm 0.89fF
C9738 a_32082_15182# rowoff_n[13] 1.20fF
C9739 a_2275_2154# a_19030_2130# 0.71fF
C9740 a_26970_17190# vcm 0.18fF
C9741 a_32082_8154# col[29] 0.38fF
C9742 a_23046_7150# VDD 2.37fF
C9743 a_34090_7150# rowoff_n[5] 1.10fF
C9744 a_22042_7150# a_23046_7150# 0.86fF
C9745 a_13006_14178# row_n[12] 0.43fF
C9746 a_29070_2130# vcm 0.89fF
C9747 a_11910_16186# a_12002_16186# 0.45fF
C9748 a_2475_16210# a_21950_16186# 0.41fF
C9749 a_2275_16210# a_19334_16226# 0.15fF
C9750 m2_1732_15002# m2_1732_13998# 0.84fF
C9751 a_23046_4138# row_n[2] 0.43fF
C9752 a_22954_8154# rowon_n[6] 0.14fF
C9753 a_27366_8194# col_n[24] 0.11fF
C9754 a_2275_4162# a_34090_4138# 0.71fF
C9755 a_19030_10162# m2_19228_10410# 0.19fF
C9756 a_3970_10162# VDD 4.33fF
C9757 a_13006_9158# a_13006_8154# 0.84fF
C9758 a_2475_7174# col[1] 0.22fF
C9759 a_2275_13198# a_12914_13174# 0.17fF
C9760 a_9994_5142# vcm 0.89fF
C9761 a_3970_12170# rowoff_n[10] 2.57fF
C9762 a_2275_1150# a_24354_1166# 0.15fF
C9763 a_2475_1150# a_26970_1126# 0.41fF
C9764 a_2275_13198# col_n[8] 0.17fF
C9765 a_2275_2154# col_n[13] 0.17fF
C9766 m3_10900_18146# VDD 0.10fF
C9767 a_19030_14178# VDD 2.78fF
C9768 a_21038_6146# col[18] 0.38fF
C9769 a_2475_10186# a_4974_10162# 0.68fF
C9770 a_9994_2130# rowon_n[0] 0.45fF
C9771 m2_34864_16006# vcm 0.72fF
C9772 a_2275_15206# a_27974_15182# 0.17fF
C9773 a_3270_2170# col_n[0] 0.11fF
C9774 a_25054_9158# vcm 0.89fF
C9775 a_20034_16186# rowoff_n[14] 1.79fF
C9776 a_21950_3134# a_22042_3134# 0.45fF
C9777 a_9994_8154# m2_10192_8402# 0.19fF
C9778 a_22954_1126# m2_22816_946# 0.31fF
C9779 a_16322_6186# col_n[13] 0.11fF
C9780 a_26362_18234# col_n[23] 0.11fF
C9781 a_2475_9182# col[18] 0.22fF
C9782 a_28066_13174# a_28066_12170# 0.84fF
C9783 a_2475_12194# a_20034_12170# 0.68fF
C9784 a_21038_11166# row_n[9] 0.43fF
C9785 a_15318_3174# vcm 0.24fF
C9786 col_n[21] rowoff_n[13] 0.19fF
C9787 a_20946_15182# rowon_n[13] 0.14fF
C9788 a_29070_4138# m2_29268_4386# 0.19fF
C9789 a_5978_12170# vcm 0.89fF
C9790 a_2161_2154# VDD 0.23fF
C9791 col[24] rowoff_n[9] 0.19fF
C9792 col[23] rowoff_n[8] 0.19fF
C9793 col[22] rowoff_n[7] 0.20fF
C9794 col[21] rowoff_n[6] 0.21fF
C9795 col[20] rowoff_n[5] 0.21fF
C9796 col[19] rowoff_n[4] 0.22fF
C9797 col[18] rowoff_n[3] 0.23fF
C9798 col[17] rowoff_n[2] 0.23fF
C9799 col[16] rowoff_n[1] 0.24fF
C9800 col[15] rowoff_n[0] 0.25fF
C9801 a_2275_15206# col_n[25] 0.17fF
C9802 a_2275_4162# col_n[30] 0.17fF
C9803 a_30986_5142# rowon_n[3] 0.14fF
C9804 m2_5748_946# m3_5880_1078# 4.41fF
C9805 a_2275_9182# a_10998_9158# 0.71fF
C9806 a_9994_4138# col[7] 0.38fF
C9807 a_2475_18218# m2_23820_18014# 0.62fF
C9808 a_18026_14178# a_19030_14178# 0.86fF
C9809 a_20034_16186# col[17] 0.38fF
C9810 a_30378_7190# vcm 0.24fF
C9811 a_2275_12194# col[15] 0.17fF
C9812 a_2275_1150# col[20] 0.17fF
C9813 a_21038_16186# vcm 0.89fF
C9814 a_17934_6146# VDD 0.29fF
C9815 a_7986_9158# rowon_n[7] 0.45fF
C9816 m2_13780_18014# col_n[11] 0.34fF
C9817 a_2275_11190# a_26058_11166# 0.71fF
C9818 a_5278_4178# col_n[2] 0.11fF
C9819 a_23958_1126# vcm 0.18fF
C9820 col_n[5] rowoff_n[14] 0.30fF
C9821 a_15318_16226# col_n[12] 0.11fF
C9822 a_8990_16186# a_8990_15182# 0.84fF
C9823 m2_1732_6970# sample 0.31fF
C9824 a_11302_10202# vcm 0.24fF
C9825 a_7986_17190# rowoff_n[15] 2.38fF
C9826 col[8] rowoff_n[10] 0.29fF
C9827 m2_17796_18014# VDD 3.73fF
C9828 a_6890_6146# rowoff_n[4] 0.69fF
C9829 a_24050_5142# ctop 4.91fF
C9830 a_14010_2130# m2_13780_946# 0.84fF
C9831 a_32994_10162# VDD 0.29fF
C9832 a_2475_8178# a_18938_8154# 0.41fF
C9833 a_2275_8178# a_16322_8194# 0.15fF
C9834 a_2275_18218# col_n[27] 0.17fF
C9835 m2_34864_2954# m2_35292_3382# 0.19fF
C9836 a_4882_4138# vcm 0.18fF
C9837 a_15926_4138# rowoff_n[2] 0.59fF
C9838 a_32994_12170# rowoff_n[10] 0.40fF
C9839 a_29070_8154# row_n[6] 0.43fF
C9840 a_8990_14178# col[6] 0.38fF
C9841 a_26362_14218# vcm 0.24fF
C9842 a_28978_12170# rowon_n[10] 0.14fF
C9843 a_2275_5166# a_9902_5142# 0.17fF
C9844 a_4974_8154# ctop 4.91fF
C9845 a_13918_13174# VDD 0.29fF
C9846 a_2275_10186# a_31382_10202# 0.15fF
C9847 a_2475_10186# a_33998_10162# 0.41fF
C9848 a_17934_10162# a_18026_10162# 0.45fF
C9849 a_24050_10162# col_n[21] 0.34fF
C9850 vcm col[22] 6.66fF
C9851 a_24962_2130# rowoff_n[0] 0.49fF
C9852 col_n[31] row_n[0] 0.37fF
C9853 VDD col[25] 7.25fF
C9854 col_n[11] col[11] 0.50fF
C9855 a_2275_11190# col_n[2] 0.17fF
C9856 a_19942_8154# vcm 0.18fF
C9857 a_4274_14218# col_n[1] 0.11fF
C9858 a_1957_4162# sample 0.35fF
C9859 a_19030_3134# a_19030_2130# 0.84fF
C9860 a_7286_17230# vcm 0.24fF
C9861 a_5978_16186# rowon_n[14] 0.45fF
C9862 m2_34864_13998# rowon_n[12] 0.42fF
C9863 a_2275_7174# a_24962_7150# 0.17fF
C9864 a_20034_12170# ctop 4.91fF
C9865 a_28978_17190# VDD 0.29fF
C9866 a_16018_6146# rowon_n[4] 0.45fF
C9867 a_2475_16210# a_3878_16186# 0.41fF
C9868 a_2275_16210# a_2874_16186# 0.17fF
C9869 a_35002_12170# vcm 0.18fF
C9870 a_31078_2130# VDD 1.54fF
C9871 a_2475_7174# col[12] 0.22fF
C9872 a_8990_4138# a_9994_4138# 0.86fF
C9873 a_2475_4162# a_17022_4138# 0.68fF
C9874 a_32994_14178# a_33086_14178# 0.45fF
C9875 a_17022_10162# rowoff_n[8] 1.94fF
C9876 a_13006_8154# col_n[10] 0.34fF
C9877 a_27062_15182# row_n[13] 0.43fF
C9878 a_2275_13198# col_n[19] 0.17fF
C9879 a_20946_13174# rowoff_n[11] 0.54fF
C9880 a_2275_2154# col_n[24] 0.17fF
C9881 a_2275_1150# a_7986_1126# 0.14fF
C9882 a_15926_15182# vcm 0.18fF
C9883 a_12002_5142# VDD 3.51fF
C9884 a_2475_6170# a_32082_6146# 0.68fF
C9885 a_34090_7150# a_34090_6146# 0.84fF
C9886 a_26058_8154# rowoff_n[6] 1.50fF
C9887 a_35494_15544# VDD 0.13fF
C9888 a_2275_10186# col[9] 0.17fF
C9889 a_2475_15206# a_10906_15182# 0.41fF
C9890 a_2275_15206# a_8290_15222# 0.15fF
C9891 a_1957_16210# rowoff_n[14] 0.14fF
C9892 a_33086_7150# col[30] 0.38fF
C9893 a_2275_3158# a_23046_3134# 0.71fF
C9894 a_2275_1150# m2_26832_946# 0.51fF
C9895 a_2475_9182# col[29] 0.22fF
C9896 a_27062_9158# VDD 1.96fF
C9897 m3_34568_1078# ctop 0.35fF
C9898 a_24050_8154# a_25054_8154# 0.86fF
C9899 a_14010_13174# rowon_n[11] 0.45fF
C9900 m2_1732_16006# row_n[14] 0.44fF
C9901 a_33086_4138# vcm 0.89fF
C9902 a_2966_11166# row_n[9] 0.41fF
C9903 a_13918_17190# a_14010_17190# 0.45fF
C9904 a_24050_3134# rowon_n[1] 0.45fF
C9905 a_2275_17214# a_23350_17230# 0.15fF
C9906 a_2475_17214# a_25966_17190# 0.41fF
C9907 col[26] rowoff_n[0] 0.17fF
C9908 col[27] rowoff_n[1] 0.17fF
C9909 col[28] rowoff_n[2] 0.16fF
C9910 col[29] rowoff_n[3] 0.15fF
C9911 col[30] rowoff_n[4] 0.15fF
C9912 col[31] rowoff_n[5] 0.14fF
C9913 sample_n rowoff_n[6] 0.55fF
C9914 a_2275_15206# rowon_n[13] 1.99fF
C9915 a_28370_7190# col_n[25] 0.11fF
C9916 a_2275_18218# a_33390_18234# 0.15fF
C9917 a_7986_12170# VDD 3.92fF
C9918 a_15014_10162# a_15014_9158# 0.84fF
C9919 a_2275_12194# col[26] 0.17fF
C9920 a_2275_14202# a_16930_14178# 0.17fF
C9921 a_2475_3158# row_n[1] 0.48fF
C9922 a_14010_7150# vcm 0.89fF
C9923 a_8898_14178# rowoff_n[12] 0.67fF
C9924 a_2475_2154# a_30986_2130# 0.41fF
C9925 a_2275_2154# a_28370_2170# 0.15fF
C9926 a_2966_16186# vcm 0.89fF
C9927 a_35002_16186# rowon_n[14] 0.14fF
C9928 a_2475_14202# m2_34864_13998# 0.56fF
C9929 a_22042_5142# col[19] 0.38fF
C9930 a_23046_16186# VDD 2.37fF
C9931 col_n[16] rowoff_n[14] 0.22fF
C9932 a_32082_17190# col[29] 0.38fF
C9933 a_2475_11190# a_8990_11166# 0.68fF
C9934 a_4974_11166# a_5978_11166# 0.86fF
C9935 a_4274_1166# vcm 0.24fF
C9936 col[19] rowoff_n[10] 0.22fF
C9937 a_2275_16210# a_31990_16186# 0.17fF
C9938 a_29070_11166# vcm 0.89fF
C9939 a_25966_1126# VDD 0.75fF
C9940 a_23958_4138# a_24050_4138# 0.45fF
C9941 a_17326_5182# col_n[14] 0.11fF
C9942 m2_16792_946# col_n[14] 0.45fF
C9943 a_27366_17230# col_n[24] 0.11fF
C9944 a_15014_17190# m2_15212_17438# 0.19fF
C9945 a_22042_10162# rowon_n[8] 0.45fF
C9946 a_30074_14178# a_30074_13174# 0.84fF
C9947 a_2475_13198# a_24050_13174# 0.68fF
C9948 a_2475_16210# col[1] 0.22fF
C9949 a_19334_5182# vcm 0.24fF
C9950 a_2475_5166# col[6] 0.22fF
C9951 a_9994_14178# vcm 0.89fF
C9952 a_6890_4138# VDD 0.29fF
C9953 m2_1732_7974# rowoff_n[6] 2.46fF
C9954 a_34090_13174# m2_34288_13422# 0.19fF
C9955 col_n[16] col[17] 6.27fF
C9956 row_n[12] ctop 0.28fF
C9957 rowon_n[5] row_n[5] 21.02fF
C9958 vcm rowoff_n[15] 2.43fF
C9959 a_2275_10186# a_15014_10162# 0.71fF
C9960 a_2275_11190# col_n[13] 0.17fF
C9961 a_10998_3134# col[8] 0.38fF
C9962 col[3] rowoff_n[11] 0.33fF
C9963 a_21038_15182# col[18] 0.38fF
C9964 a_20034_15182# a_21038_15182# 0.86fF
C9965 a_35398_9198# vcm 0.24fF
C9966 a_9902_4138# rowon_n[2] 0.14fF
C9967 a_3270_11206# col_n[0] 0.11fF
C9968 a_25054_18194# vcm 0.15fF
C9969 a_13006_3134# ctop 4.91fF
C9970 a_21950_8154# VDD 0.29fF
C9971 a_2275_8178# col[3] 0.17fF
C9972 a_5978_15182# m2_6176_15430# 0.19fF
C9973 a_2475_7174# a_7894_7150# 0.41fF
C9974 a_2275_7174# a_5278_7190# 0.15fF
C9975 a_4882_7150# a_4974_7150# 0.45fF
C9976 a_6282_3174# col_n[3] 0.11fF
C9977 a_2275_12194# a_30074_12170# 0.71fF
C9978 a_16322_15222# col_n[13] 0.11fF
C9979 a_27974_3134# vcm 0.18fF
C9980 a_10998_17190# a_10998_16186# 0.84fF
C9981 a_2475_7174# col[23] 0.22fF
C9982 a_2966_3134# m2_3164_3382# 0.19fF
C9983 a_15318_12210# vcm 0.24fF
C9984 a_7894_5142# rowoff_n[3] 0.68fF
C9985 a_25054_11166# m2_25252_11414# 0.19fF
C9986 a_28066_7150# ctop 4.91fF
C9987 a_2161_11190# VDD 0.23fF
C9988 m3_29976_18146# m3_30980_18146# 0.21fF
C9989 a_20034_17190# rowon_n[15] 0.45fF
C9990 a_2275_9182# a_20338_9198# 0.15fF
C9991 a_2475_9182# a_22954_9158# 0.41fF
C9992 a_2275_13198# col_n[30] 0.17fF
C9993 a_16930_3134# rowoff_n[1] 0.58fF
C9994 a_8898_6146# vcm 0.18fF
C9995 a_30074_7150# rowon_n[5] 0.45fF
C9996 a_9994_13174# col[7] 0.38fF
C9997 a_2275_13198# rowoff_n[11] 0.81fF
C9998 a_30074_2130# a_31078_2130# 0.86fF
C9999 a_30378_16226# vcm 0.24fF
C10000 a_2275_6170# a_13918_6146# 0.17fF
C10001 a_2275_10186# col[20] 0.17fF
C10002 a_8990_10162# ctop 4.91fF
C10003 a_25054_9158# col_n[22] 0.34fF
C10004 a_17934_15182# VDD 0.29fF
C10005 a_19942_11166# a_20034_11166# 0.45fF
C10006 a_7986_7150# row_n[5] 0.43fF
C10007 a_5278_13214# col_n[2] 0.11fF
C10008 a_7894_11166# rowon_n[9] 0.14fF
C10009 a_2966_3134# col_n[0] 0.34fF
C10010 a_23958_10162# vcm 0.18fF
C10011 a_16018_9158# m2_16216_9406# 0.19fF
C10012 a_2475_3158# a_5978_3134# 0.68fF
C10013 a_21038_4138# a_21038_3134# 0.84fF
C10014 m3_30980_18146# ctop 0.21fF
C10015 m2_28840_18014# col[26] 0.37fF
C10016 a_2275_8178# a_28978_8154# 0.17fF
C10017 a_24050_14178# ctop 4.91fF
C10018 a_8990_11166# rowoff_n[9] 2.33fF
C10019 a_2275_17214# a_6982_17190# 0.71fF
C10020 a_4882_13174# vcm 0.18fF
C10021 a_2475_5166# a_21038_5142# 0.68fF
C10022 a_10998_5142# a_12002_5142# 0.86fF
C10023 a_2275_18218# a_17022_18194# 0.14fF
C10024 a_2475_3158# col[0] 0.20fF
C10025 a_4974_17190# ctop 4.93fF
C10026 a_18026_9158# rowoff_n[7] 1.89fF
C10027 a_14010_7150# col_n[11] 0.34fF
C10028 a_28066_14178# rowon_n[12] 0.45fF
C10029 a_35002_15182# a_35094_15182# 0.11fF
C10030 a_25054_15182# rowoff_n[13] 1.54fF
C10031 a_6982_7150# m2_7180_7398# 0.19fF
C10032 a_2275_2154# a_12002_2130# 0.71fF
C10033 a_2275_9182# col_n[7] 0.17fF
C10034 a_19942_17190# vcm 0.18fF
C10035 col_n[27] rowoff_n[14] 0.14fF
C10036 a_16018_7150# VDD 3.09fF
C10037 a_27062_7150# rowoff_n[5] 1.45fF
C10038 a_1957_13198# sample 0.35fF
C10039 col[30] rowoff_n[10] 0.15fF
C10040 a_5978_14178# row_n[12] 0.43fF
C10041 a_22042_2130# vcm 0.89fF
C10042 a_2275_16210# a_12306_16226# 0.15fF
C10043 a_2475_16210# a_14922_16186# 0.41fF
C10044 a_34090_6146# col[31] 0.38fF
C10045 a_26058_3134# m2_26256_3382# 0.19fF
C10046 a_16018_4138# row_n[2] 0.43fF
C10047 a_15926_8154# rowon_n[6] 0.14fF
C10048 a_2275_4162# a_27062_4138# 0.71fF
C10049 a_31078_11166# VDD 1.54fF
C10050 m3_19936_1078# m3_20940_1078# 0.21fF
C10051 a_26058_9158# a_27062_9158# 0.86fF
C10052 a_2475_16210# col[12] 0.22fF
C10053 a_2475_5166# col[17] 0.22fF
C10054 a_2275_13198# a_5886_13174# 0.17fF
C10055 a_2874_5142# vcm 0.18fF
C10056 a_29374_6186# col_n[26] 0.11fF
C10057 a_15926_18194# a_16018_18194# 0.11fF
C10058 a_13006_17190# col_n[10] 0.34fF
C10059 col_n[11] rowoff_n[15] 0.26fF
C10060 col_n[22] col[22] 0.50fF
C10061 rowon_n[6] ctop 0.37fF
C10062 a_2275_1150# a_17326_1166# 0.15fF
C10063 a_10906_1126# a_10998_1126# 0.11fF
C10064 a_2475_1150# a_19942_1126# 0.44fF
C10065 a_2275_11190# col_n[24] 0.17fF
C10066 col[14] rowoff_n[11] 0.25fF
C10067 a_12002_14178# VDD 3.51fF
C10068 a_17022_11166# a_17022_10162# 0.84fF
C10069 m2_34864_2954# row_n[1] 0.38fF
C10070 a_2874_2130# rowon_n[0] 0.14fF
C10071 a_2275_15206# a_20946_15182# 0.17fF
C10072 a_18026_9158# vcm 0.89fF
C10073 a_13006_16186# rowoff_n[14] 2.13fF
C10074 a_2275_8178# col[14] 0.17fF
C10075 a_2475_3158# a_35002_3134# 0.41fF
C10076 a_2275_3158# a_32386_3174# 0.15fF
C10077 a_23046_4138# col[20] 0.38fF
C10078 a_3878_8154# VDD 0.29fF
C10079 a_33086_16186# col[30] 0.38fF
C10080 a_2475_12194# a_13006_12170# 0.68fF
C10081 a_6982_12170# a_7986_12170# 0.86fF
C10082 a_8290_3174# vcm 0.24fF
C10083 a_14010_11166# row_n[9] 0.43fF
C10084 a_2275_17214# a_34394_17230# 0.15fF
C10085 a_13918_15182# rowon_n[13] 0.14fF
C10086 a_33086_13174# vcm 0.89fF
C10087 a_18330_4178# col_n[15] 0.11fF
C10088 a_29982_3134# VDD 0.29fF
C10089 a_25966_5142# a_26058_5142# 0.45fF
C10090 a_28370_16226# col_n[25] 0.11fF
C10091 a_2275_13198# row_n[11] 26.41fF
C10092 a_23958_5142# rowon_n[3] 0.14fF
C10093 m2_31852_946# m2_32856_946# 0.86fF
C10094 a_2275_9182# a_3970_9158# 0.71fF
C10095 a_2475_18218# m2_9764_18014# 0.62fF
C10096 a_2475_14202# a_28066_14178# 0.68fF
C10097 a_32082_15182# a_32082_14178# 0.84fF
C10098 a_23350_7190# vcm 0.24fF
C10099 a_2275_10186# col[31] 0.17fF
C10100 a_2475_1150# ctop 0.16fF
C10101 a_14010_16186# vcm 0.89fF
C10102 a_10906_6146# VDD 0.29fF
C10103 a_12002_2130# col[9] 0.38fF
C10104 a_2275_11190# a_19030_11166# 0.71fF
C10105 a_22042_14178# col[19] 0.38fF
C10106 a_16930_1126# vcm 0.18fF
C10107 a_2275_7174# col_n[1] 0.17fF
C10108 a_22042_16186# a_23046_16186# 0.86fF
C10109 a_4274_10202# vcm 0.24fF
C10110 m2_3740_18014# VDD 5.20fF
C10111 a_2475_9182# m2_1732_8978# 0.16fF
C10112 a_17022_5142# ctop 4.91fF
C10113 a_7286_2170# col_n[4] 0.11fF
C10114 a_25966_10162# VDD 0.29fF
C10115 a_2161_18218# a_2275_18218# 0.17fF
C10116 a_2275_8178# a_9294_8194# 0.15fF
C10117 a_2475_8178# a_11910_8154# 0.41fF
C10118 a_6890_8154# a_6982_8154# 0.45fF
C10119 a_17326_14218# col_n[14] 0.11fF
C10120 m2_1732_1950# sample_n 0.12fF
C10121 a_2275_13198# a_34090_13174# 0.71fF
C10122 a_31990_5142# vcm 0.18fF
C10123 a_8898_4138# rowoff_n[2] 0.67fF
C10124 a_25966_12170# rowoff_n[10] 0.48fF
C10125 a_22042_8154# row_n[6] 0.43fF
C10126 a_2475_14202# col[6] 0.22fF
C10127 a_19334_14218# vcm 0.24fF
C10128 a_21950_12170# rowon_n[10] 0.14fF
C10129 a_2475_3158# col[11] 0.22fF
C10130 a_2161_5166# a_2275_5166# 0.17fF
C10131 a_2475_5166# a_2966_5142# 0.65fF
C10132 a_32082_9158# ctop 4.91fF
C10133 a_6890_13174# VDD 0.29fF
C10134 a_2275_10186# a_24354_10202# 0.15fF
C10135 a_2475_10186# a_26970_10162# 0.41fF
C10136 a_17934_2130# rowoff_n[0] 0.57fF
C10137 a_31990_2130# rowon_n[0] 0.14fF
C10138 a_10998_12170# col[8] 0.38fF
C10139 a_2275_9182# col_n[18] 0.17fF
C10140 a_12914_8154# vcm 0.18fF
C10141 a_32082_3134# a_33086_3134# 0.86fF
C10142 a_35398_18234# vcm 0.24fF
C10143 m2_26832_946# col_n[24] 0.45fF
C10144 m2_4744_18014# m3_4876_18146# 4.41fF
C10145 a_26058_8154# col_n[23] 0.34fF
C10146 a_2275_7174# a_17934_7150# 0.17fF
C10147 a_13006_12170# ctop 4.91fF
C10148 a_21950_17190# VDD 0.29fF
C10149 a_2275_17214# col[3] 0.17fF
C10150 a_21950_12170# a_22042_12170# 0.45fF
C10151 a_8990_6146# rowon_n[4] 0.45fF
C10152 a_2275_6170# col[8] 0.17fF
C10153 a_6282_12210# col_n[3] 0.11fF
C10154 a_27974_12170# vcm 0.18fF
C10155 a_24050_2130# VDD 2.27fF
C10156 a_2475_16210# col[23] 0.22fF
C10157 a_2475_4162# a_9994_4138# 0.68fF
C10158 a_23046_5142# a_23046_4138# 0.84fF
C10159 a_2475_5166# col[28] 0.22fF
C10160 m3_34996_10114# m3_34996_9110# 0.20fF
C10161 a_2275_9182# a_32994_9158# 0.17fF
C10162 a_28066_16186# ctop 4.91fF
C10163 a_9994_10162# rowoff_n[8] 2.28fF
C10164 col_n[27] col[28] 6.14fF
C10165 row_n[1] ctop 0.28fF
C10166 col_n[22] rowoff_n[15] 0.18fF
C10167 a_20034_15182# row_n[13] 0.43fF
C10168 a_13918_13174# rowoff_n[11] 0.61fF
C10169 col[25] rowoff_n[11] 0.18fF
C10170 a_8898_15182# vcm 0.18fF
C10171 a_4974_5142# VDD 4.23fF
C10172 a_30074_5142# row_n[3] 0.43fF
C10173 a_2475_6170# a_25054_6146# 0.68fF
C10174 a_13006_6146# a_14010_6146# 0.86fF
C10175 a_29982_9158# rowon_n[7] 0.14fF
C10176 a_19030_8154# rowoff_n[6] 1.84fF
C10177 a_15014_6146# col_n[12] 0.34fF
C10178 a_2275_8178# col[25] 0.17fF
C10179 a_29982_17190# rowoff_n[15] 0.43fF
C10180 a_28066_6146# rowoff_n[4] 1.40fF
C10181 a_2966_12170# col_n[0] 0.34fF
C10182 a_2275_3158# a_16018_3134# 0.71fF
C10183 a_5886_1126# m2_5748_946# 0.31fF
C10184 a_2475_1150# m2_12776_946# 0.62fF
C10185 m3_6884_1078# ctop 0.21fF
C10186 a_20034_9158# VDD 2.68fF
C10187 a_12002_16186# m2_12200_16434# 0.19fF
C10188 a_3970_8154# a_3970_7150# 0.84fF
C10189 a_6982_13174# rowon_n[11] 0.45fF
C10190 a_26058_4138# vcm 0.89fF
C10191 a_17022_3134# rowon_n[1] 0.45fF
C10192 a_2275_17214# a_16322_17230# 0.15fF
C10193 a_2475_17214# a_18938_17190# 0.41fF
C10194 col[9] rowoff_n[12] 0.29fF
C10195 a_2275_4162# m2_34864_3958# 0.51fF
C10196 a_2275_5166# a_31078_5142# 0.71fF
C10197 a_31078_12170# m2_31276_12418# 0.19fF
C10198 a_2275_18218# a_26362_18234# 0.15fF
C10199 m2_12776_946# m2_13204_1374# 0.19fF
C10200 a_28066_10162# a_29070_10162# 0.86fF
C10201 a_2475_12194# col[0] 0.20fF
C10202 a_30378_5182# col_n[27] 0.11fF
C10203 a_3970_4138# col_n[1] 0.34fF
C10204 a_2275_14202# a_9902_14178# 0.17fF
C10205 a_2475_1150# col[5] 0.22fF
C10206 a_14010_16186# col_n[11] 0.34fF
C10207 a_6982_7150# vcm 0.89fF
C10208 a_28066_12170# row_n[10] 0.43fF
C10209 a_2475_2154# a_23958_2130# 0.41fF
C10210 a_2275_2154# a_21342_2170# 0.15fF
C10211 a_12914_2130# a_13006_2130# 0.45fF
C10212 a_27974_16186# rowon_n[14] 0.14fF
C10213 a_16018_16186# VDD 3.09fF
C10214 a_2275_7174# col_n[12] 0.17fF
C10215 a_19030_12170# a_19030_11166# 0.84fF
C10216 a_31382_2170# vcm 0.24fF
C10217 a_2275_16210# a_24962_16186# 0.17fF
C10218 a_35002_3134# m2_34864_2954# 0.33fF
C10219 a_22042_11166# vcm 0.89fF
C10220 a_24050_3134# col[21] 0.38fF
C10221 a_18938_1126# VDD 0.72fF
C10222 a_34090_15182# col[31] 0.38fF
C10223 a_22042_10162# m2_22240_10410# 0.19fF
C10224 a_2966_4138# a_2966_3134# 0.84fF
C10225 a_2275_4162# col[2] 0.17fF
C10226 a_15014_10162# rowon_n[8] 0.45fF
C10227 a_2475_13198# a_17022_13174# 0.68fF
C10228 a_8990_13174# a_9994_13174# 0.86fF
C10229 a_2475_14202# col[17] 0.22fF
C10230 a_12306_5182# vcm 0.24fF
C10231 m2_6752_946# vcm 0.71fF
C10232 a_2475_3158# col[22] 0.22fF
C10233 a_19334_3174# col_n[16] 0.11fF
C10234 a_2275_1150# a_29982_1126# 0.17fF
C10235 a_29374_15222# col_n[26] 0.11fF
C10236 a_2874_14178# vcm 0.18fF
C10237 a_2475_18218# col[8] 0.22fF
C10238 a_3878_12170# rowon_n[10] 0.14fF
C10239 a_33998_5142# VDD 0.29fF
C10240 a_27974_6146# a_28066_6146# 0.45fF
C10241 a_2275_10186# a_7986_10162# 0.71fF
C10242 a_2275_9182# col_n[29] 0.17fF
C10243 a_34090_16186# a_34090_15182# 0.84fF
C10244 a_2475_15206# a_32082_15182# 0.68fF
C10245 a_27366_9198# vcm 0.24fF
C10246 a_13006_8154# m2_13204_8402# 0.19fF
C10247 a_5978_3134# ctop 4.91fF
C10248 a_18026_18194# vcm 0.15fF
C10249 a_2275_17214# col[14] 0.17fF
C10250 a_14922_8154# VDD 0.29fF
C10251 a_2275_6170# col[19] 0.17fF
C10252 a_23046_13174# col[20] 0.38fF
C10253 a_3878_17190# VDD 0.29fF
C10254 a_2275_12194# a_23046_12170# 0.71fF
C10255 a_20946_3134# vcm 0.18fF
C10256 a_24050_17190# a_25054_17190# 0.86fF
C10257 a_32082_4138# m2_32280_4386# 0.19fF
C10258 a_8290_12210# vcm 0.24fF
C10259 a_8290_1166# col_n[5] 0.11fF
C10260 a_21038_7150# ctop 4.91fF
C10261 a_18330_13214# col_n[15] 0.11fF
C10262 a_29982_12170# VDD 0.29fF
C10263 m2_10768_946# m3_10900_1078# 4.41fF
C10264 m3_15920_18146# m3_16924_18146# 0.21fF
C10265 a_13006_17190# rowon_n[15] 0.45fF
C10266 a_2275_9182# a_13310_9198# 0.15fF
C10267 a_2475_9182# a_15926_9158# 0.41fF
C10268 a_8898_9158# a_8990_9158# 0.45fF
C10269 row_n[15] rowoff_n[15] 0.64fF
C10270 rowon_n[14] sample_n 0.15fF
C10271 a_9902_3134# rowoff_n[1] 0.66fF
C10272 m2_1732_5966# m2_2160_6394# 0.19fF
C10273 a_1957_15206# row_n[13] 0.29fF
C10274 a_34394_7190# vcm 0.24fF
C10275 a_23046_7150# rowon_n[5] 0.45fF
C10276 a_30074_14178# rowoff_n[12] 1.30fF
C10277 a_3970_6146# m2_4168_6394# 0.19fF
C10278 a_23350_16226# vcm 0.24fF
C10279 a_2275_6170# a_6890_6146# 0.17fF
C10280 a_10906_15182# VDD 0.29fF
C10281 a_2275_11190# a_28370_11206# 0.15fF
C10282 a_2475_11190# a_30986_11166# 0.41fF
C10283 a_12002_11166# col[9] 0.38fF
C10284 a_16930_10162# vcm 0.18fF
C10285 a_2275_16210# col_n[1] 0.17fF
C10286 a_34090_16186# row_n[14] 0.43fF
C10287 a_27062_7150# col_n[24] 0.34fF
C10288 a_2275_5166# col_n[6] 0.17fF
C10289 a_1957_9182# VDD 0.28fF
C10290 m3_2868_18146# ctop 0.21fF
C10291 a_2275_8178# a_21950_8154# 0.17fF
C10292 a_17022_14178# ctop 4.91fF
C10293 a_7286_11206# col_n[4] 0.11fF
C10294 a_2966_9158# col[0] 0.38fF
C10295 a_23958_13174# a_24050_13174# 0.45fF
C10296 col[20] rowoff_n[12] 0.21fF
C10297 a_2475_11190# rowoff_n[9] 4.75fF
C10298 a_31990_14178# vcm 0.18fF
C10299 m2_34864_4962# rowon_n[3] 0.42fF
C10300 a_28066_4138# VDD 1.85fF
C10301 a_25054_6146# a_25054_5142# 0.84fF
C10302 a_2475_5166# a_14010_5142# 0.68fF
C10303 a_2275_18218# a_9994_18194# 0.14fF
C10304 a_2475_12194# col[11] 0.22fF
C10305 a_10998_9158# rowoff_n[7] 2.23fF
C10306 a_2475_1150# col[16] 0.21fF
C10307 a_21038_14178# rowon_n[12] 0.45fF
C10308 m2_34864_9982# m2_34864_8978# 0.84fF
C10309 a_18026_15182# rowoff_n[13] 1.89fF
C10310 a_31078_4138# rowon_n[2] 0.45fF
C10311 a_2275_2154# a_4974_2130# 0.71fF
C10312 a_3878_2130# a_3970_2130# 0.45fF
C10313 a_12914_17190# vcm 0.18fF
C10314 a_2275_7174# col_n[23] 0.17fF
C10315 a_8990_7150# VDD 3.82fF
C10316 a_20034_7150# rowoff_n[5] 1.79fF
C10317 a_2475_7174# a_29070_7150# 0.68fF
C10318 a_15014_7150# a_16018_7150# 0.86fF
C10319 a_16018_5142# col_n[13] 0.34fF
C10320 a_26058_17190# col_n[23] 0.34fF
C10321 col[4] rowoff_n[13] 0.32fF
C10322 a_15014_2130# vcm 0.89fF
C10323 a_2275_16210# a_5278_16226# 0.15fF
C10324 a_2475_16210# a_7894_16186# 0.41fF
C10325 a_4882_16186# a_4974_16186# 0.45fF
C10326 a_2275_15206# col[8] 0.17fF
C10327 a_8990_4138# row_n[2] 0.43fF
C10328 a_2275_4162# col[13] 0.17fF
C10329 a_29070_5142# rowoff_n[3] 1.35fF
C10330 m2_7756_18014# col_n[5] 0.33fF
C10331 a_8898_8154# rowon_n[6] 0.14fF
C10332 a_2275_4162# a_20034_4138# 0.71fF
C10333 a_24050_11166# VDD 2.27fF
C10334 m3_5880_1078# m3_6884_1078# 0.21fF
C10335 a_5978_9158# a_5978_8154# 0.84fF
C10336 a_2475_14202# col[28] 0.22fF
C10337 a_30074_6146# vcm 0.89fF
C10338 a_2475_18218# col[19] 0.22fF
C10339 a_2275_1150# a_10298_1166# 0.15fF
C10340 a_2475_1150# a_12914_1126# 0.41fF
C10341 m2_10768_946# VDD 6.10fF
C10342 a_2275_6170# a_35094_6146# 0.14fF
C10343 a_4974_14178# VDD 4.23fF
C10344 m2_1732_6970# row_n[5] 0.44fF
C10345 a_30074_11166# a_31078_11166# 0.86fF
C10346 a_31382_4178# col_n[28] 0.11fF
C10347 a_4974_3134# col_n[2] 0.34fF
C10348 a_15014_15182# col_n[12] 0.34fF
C10349 a_2275_15206# a_13918_15182# 0.17fF
C10350 a_29070_11166# rowon_n[9] 0.45fF
C10351 a_2275_17214# col[25] 0.17fF
C10352 a_10998_9158# vcm 0.89fF
C10353 a_5978_16186# rowoff_n[14] 2.47fF
C10354 a_2275_6170# col[30] 0.17fF
C10355 a_2275_3158# a_25358_3174# 0.15fF
C10356 a_2475_3158# a_27974_3134# 0.41fF
C10357 a_14922_3134# a_15014_3134# 0.45fF
C10358 a_2275_18218# col[10] 0.17fF
C10359 a_2275_1150# m2_34864_946# 0.48fF
C10360 a_21038_13174# a_21038_12170# 0.84fF
C10361 a_2475_12194# a_5978_12170# 0.68fF
C10362 a_2275_3158# vcm 7.71fF
C10363 a_6982_11166# row_n[9] 0.43fF
C10364 a_30986_11166# rowoff_n[9] 0.42fF
C10365 a_2275_17214# a_28978_17190# 0.17fF
C10366 a_25054_2130# col[22] 0.38fF
C10367 a_6890_15182# rowon_n[13] 0.14fF
C10368 a_26058_13174# vcm 0.89fF
C10369 a_22954_3134# VDD 0.29fF
C10370 row_n[9] sample_n 0.16fF
C10371 ctop col[11] 0.13fF
C10372 a_2966_7150# ctop 4.82fF
C10373 a_16930_5142# rowon_n[3] 0.14fF
C10374 m2_24824_946# m2_25828_946# 0.86fF
C10375 a_2475_14202# a_21038_14178# 0.68fF
C10376 a_10998_14178# a_12002_14178# 0.86fF
C10377 a_20338_2170# col_n[17] 0.11fF
C10378 a_16322_7190# vcm 0.24fF
C10379 a_3970_13174# col_n[1] 0.34fF
C10380 a_30378_14218# col_n[27] 0.11fF
C10381 a_2275_2154# a_33998_2130# 0.17fF
C10382 a_2475_10186# col[5] 0.22fF
C10383 a_29070_2130# ctop 4.93fF
C10384 a_6982_16186# vcm 0.89fF
C10385 a_29982_7150# a_30074_7150# 0.45fF
C10386 a_2275_11190# a_12002_11166# 0.71fF
C10387 a_9902_1126# vcm 0.18fF
C10388 a_2275_16210# col_n[12] 0.17fF
C10389 a_2275_5166# col_n[17] 0.17fF
C10390 a_31382_11206# vcm 0.24fF
C10391 a_29470_1488# VDD 0.12fF
C10392 a_9994_5142# ctop 4.91fF
C10393 a_24050_12170# col[21] 0.38fF
C10394 a_18938_10162# VDD 0.29fF
C10395 col[31] rowoff_n[12] 0.14fF
C10396 a_2275_8178# a_3878_8154# 0.17fF
C10397 a_2475_8178# a_4882_8154# 0.41fF
C10398 a_18026_17190# m2_18224_17438# 0.19fF
C10399 a_2275_13198# col[2] 0.17fF
C10400 a_2275_2154# col[7] 0.17fF
C10401 a_2275_13198# a_27062_13174# 0.71fF
C10402 a_24962_5142# vcm 0.18fF
C10403 a_18938_12170# rowoff_n[10] 0.56fF
C10404 m2_29844_946# vcm 0.71fF
C10405 a_2275_18218# m2_26832_18014# 0.51fF
C10406 a_15014_8154# row_n[6] 0.43fF
C10407 a_12306_14218# vcm 0.24fF
C10408 a_14922_12170# rowon_n[10] 0.14fF
C10409 a_2475_12194# col[22] 0.22fF
C10410 a_19334_12210# col_n[16] 0.11fF
C10411 a_2475_1150# col[27] 0.22fF
C10412 a_25054_9158# ctop 4.91fF
C10413 a_33998_14178# VDD 0.29fF
C10414 a_10906_10162# a_10998_10162# 0.45fF
C10415 a_2275_10186# a_17326_10202# 0.15fF
C10416 a_2475_10186# a_19942_10162# 0.41fF
C10417 a_24962_2130# rowon_n[0] 0.14fF
C10418 a_10906_2130# rowoff_n[0] 0.65fF
C10419 a_2966_14178# rowon_n[12] 0.45fF
C10420 a_5886_8154# vcm 0.18fF
C10421 a_35002_16186# rowoff_n[14] 0.38fF
C10422 a_12002_3134# a_12002_2130# 0.84fF
C10423 a_27366_18234# vcm 0.25fF
C10424 col[15] rowoff_n[13] 0.25fF
C10425 a_1957_7174# rowoff_n[5] 0.14fF
C10426 a_2275_7174# a_10906_7150# 0.17fF
C10427 a_8990_15182# m2_9188_15430# 0.19fF
C10428 a_5978_12170# ctop 4.91fF
C10429 a_13006_10162# col[10] 0.38fF
C10430 a_14922_17190# VDD 0.29fF
C10431 sample rowoff_n[9] 0.22fF
C10432 VDD rowoff_n[8] 87.22fF
C10433 a_2275_15206# col[19] 0.17fF
C10434 a_2275_12194# a_32386_12210# 0.15fF
C10435 a_2475_12194# a_35002_12170# 0.41fF
C10436 a_2475_6170# rowon_n[4] 0.40fF
C10437 a_2275_4162# col[24] 0.17fF
C10438 a_28066_6146# col_n[25] 0.34fF
C10439 a_20946_12170# vcm 0.18fF
C10440 a_17022_2130# VDD 2.99fF
C10441 a_1957_4162# a_2275_4162# 0.19fF
C10442 a_2475_4162# a_2874_4138# 0.41fF
C10443 a_28066_11166# m2_28264_11414# 0.19fF
C10444 m3_34996_17142# m3_34996_16138# 0.20fF
C10445 a_8290_10202# col_n[5] 0.11fF
C10446 a_2275_9182# a_25966_9158# 0.17fF
C10447 a_18938_18194# m2_18800_18014# 0.34fF
C10448 a_21038_16186# ctop 4.91fF
C10449 a_2475_18218# col[30] 0.22fF
C10450 a_25966_14178# a_26058_14178# 0.45fF
C10451 a_2874_10162# rowoff_n[8] 0.74fF
C10452 a_13006_15182# row_n[13] 0.43fF
C10453 a_6890_13174# rowoff_n[11] 0.69fF
C10454 m2_10768_946# col_n[8] 0.45fF
C10455 a_34394_16226# vcm 0.24fF
C10456 a_32082_6146# VDD 1.44fF
C10457 a_23046_5142# row_n[3] 0.43fF
C10458 a_27062_7150# a_27062_6146# 0.84fF
C10459 a_2475_6170# a_18026_6146# 0.68fF
C10460 a_22954_9158# rowon_n[7] 0.14fF
C10461 a_12002_8154# rowoff_n[6] 2.18fF
C10462 a_2275_18218# col[21] 0.17fF
C10463 a_22954_17190# rowoff_n[15] 0.51fF
C10464 a_21038_6146# rowoff_n[4] 1.74fF
C10465 a_2275_3158# a_8990_3134# 0.71fF
C10466 a_19030_9158# m2_19228_9406# 0.19fF
C10467 a_17022_4138# col_n[14] 0.34fF
C10468 m3_1864_12122# ctop 0.22fF
C10469 a_13006_9158# VDD 3.40fF
C10470 a_27062_16186# col_n[24] 0.34fF
C10471 a_2275_14202# col_n[6] 0.17fF
C10472 a_17022_8154# a_18026_8154# 0.86fF
C10473 a_2475_8178# a_33086_8154# 0.68fF
C10474 a_2275_3158# col_n[11] 0.17fF
C10475 a_19030_4138# vcm 0.89fF
C10476 a_9994_3134# rowon_n[1] 0.45fF
C10477 a_30074_4138# rowoff_n[2] 1.30fF
C10478 a_2275_17214# a_9294_17230# 0.15fF
C10479 a_2475_17214# a_11910_17190# 0.41fF
C10480 a_6890_17190# a_6982_17190# 0.45fF
C10481 VDD col_n[0] 16.44fF
C10482 rowon_n[3] sample_n 0.15fF
C10483 ctop col[22] 0.13fF
C10484 a_2275_5166# a_24050_5142# 0.71fF
C10485 a_2275_18218# a_19334_18234# 0.15fF
C10486 a_28066_13174# VDD 1.85fF
C10487 m2_5748_946# m2_6176_1374# 0.19fF
C10488 a_7986_10162# a_7986_9158# 0.84fF
C10489 a_2475_14202# a_2966_14178# 0.65fF
C10490 a_2161_14202# a_2275_14202# 0.17fF
C10491 a_2475_10186# col[16] 0.22fF
C10492 a_34090_8154# vcm 0.89fF
C10493 m2_1732_946# m3_1864_1078# 4.44fF
C10494 a_21038_12170# row_n[10] 0.43fF
C10495 a_2275_2154# a_14314_2170# 0.15fF
C10496 a_2475_2154# a_16930_2130# 0.41fF
C10497 a_9994_7150# m2_10192_7398# 0.19fF
C10498 a_20946_16186# rowon_n[14] 0.14fF
C10499 a_32386_3174# col_n[29] 0.11fF
C10500 a_5978_2130# col_n[3] 0.34fF
C10501 a_2275_16210# col_n[23] 0.17fF
C10502 a_31078_2130# row_n[0] 0.43fF
C10503 a_8990_16186# VDD 3.82fF
C10504 a_16018_14178# col_n[13] 0.34fF
C10505 a_32082_12170# a_33086_12170# 0.86fF
C10506 a_2275_5166# col_n[28] 0.17fF
C10507 a_30986_6146# rowon_n[4] 0.14fF
C10508 a_24354_2170# vcm 0.24fF
C10509 a_2275_16210# a_17934_16186# 0.17fF
C10510 a_29070_3134# m2_29268_3382# 0.19fF
C10511 a_15014_11166# vcm 0.89fF
C10512 a_11910_1126# VDD 0.91fF
C10513 a_2275_4162# a_29374_4178# 0.15fF
C10514 a_2475_4162# a_31990_4138# 0.41fF
C10515 a_16930_4138# a_17022_4138# 0.45fF
C10516 a_2275_13198# col[13] 0.17fF
C10517 a_2275_2154# col[18] 0.17fF
C10518 a_15014_17190# m2_14784_18014# 0.84fF
C10519 a_7986_10162# rowon_n[8] 0.45fF
C10520 a_2475_13198# a_9994_13174# 0.68fF
C10521 a_23046_14178# a_23046_13174# 0.84fF
C10522 a_31990_10162# rowoff_n[8] 0.41fF
C10523 a_5278_5182# vcm 0.24fF
C10524 m2_21236_2378# a_21038_2130# 0.19fF
C10525 a_2275_1150# a_22954_1126# 0.17fF
C10526 m2_22816_18014# col[20] 0.39fF
C10527 a_30074_15182# vcm 0.89fF
C10528 a_26970_5142# VDD 0.29fF
C10529 m2_33860_946# VDD 1.49fF
C10530 a_21342_1166# col_n[18] 0.11fF
C10531 a_2475_15206# a_25054_15182# 0.68fF
C10532 a_13006_15182# a_14010_15182# 0.86fF
C10533 a_31382_13214# col_n[28] 0.11fF
C10534 a_4974_12170# col_n[2] 0.34fF
C10535 a_20338_9198# vcm 0.24fF
C10536 col[26] rowoff_n[13] 0.17fF
C10537 a_33086_4138# ctop 4.91fF
C10538 a_10998_18194# vcm 0.15fF
C10539 col_n[4] rowoff_n[4] 0.31fF
C10540 vcm rowoff_n[0] 2.43fF
C10541 col_n[7] rowoff_n[7] 0.29fF
C10542 col_n[8] rowoff_n[8] 0.28fF
C10543 col_n[5] rowoff_n[5] 0.30fF
C10544 col_n[2] rowoff_n[2] 0.32fF
C10545 col_n[9] rowoff_n[9] 0.27fF
C10546 col_n[6] rowoff_n[6] 0.29fF
C10547 col_n[1] rowoff_n[1] 0.33fF
C10548 col_n[3] rowoff_n[3] 0.32fF
C10549 a_29070_9158# row_n[7] 0.43fF
C10550 a_7894_8154# VDD 0.29fF
C10551 a_2275_15206# col[30] 0.17fF
C10552 a_31990_8154# a_32082_8154# 0.45fF
C10553 a_28978_13174# rowon_n[11] 0.14fF
C10554 a_2275_12194# a_16018_12170# 0.71fF
C10555 a_13918_3134# vcm 0.18fF
C10556 a_3970_17190# a_3970_16186# 0.84fF
C10557 m2_30848_18014# m2_31852_18014# 0.86fF
C10558 a_2275_12194# vcm 7.71fF
C10559 a_25054_11166# col[22] 0.38fF
C10560 a_2275_1150# col_n[5] 0.17fF
C10561 a_14010_7150# ctop 4.91fF
C10562 a_22954_12170# VDD 0.29fF
C10563 m3_1864_18146# m3_2868_18146# 0.21fF
C10564 a_5978_17190# rowon_n[15] 0.45fF
C10565 a_2275_9182# a_6282_9198# 0.15fF
C10566 a_2475_9182# a_8898_9158# 0.41fF
C10567 a_2966_16186# ctop 4.82fF
C10568 a_2275_14202# a_31078_14178# 0.71fF
C10569 a_2161_3158# rowoff_n[1] 0.14fF
C10570 col[10] rowoff_n[14] 0.28fF
C10571 a_16018_7150# rowon_n[5] 0.45fF
C10572 a_28978_7150# vcm 0.18fF
C10573 a_23046_14178# rowoff_n[12] 1.64fF
C10574 a_20338_11206# col_n[17] 0.11fF
C10575 a_23046_2130# a_24050_2130# 0.86fF
C10576 a_16322_16226# vcm 0.24fF
C10577 a_29070_11166# ctop 4.91fF
C10578 a_2475_8178# col[10] 0.22fF
C10579 a_12914_11166# a_13006_11166# 0.45fF
C10580 a_2275_11190# a_21342_11206# 0.15fF
C10581 a_2475_11190# a_23958_11166# 0.41fF
C10582 a_9902_10162# vcm 0.18fF
C10583 a_27062_16186# row_n[14] 0.43fF
C10584 a_2275_14202# col_n[17] 0.17fF
C10585 a_2966_6146# rowoff_n[4] 2.62fF
C10586 a_14010_4138# a_14010_3134# 0.84fF
C10587 a_2275_3158# col_n[22] 0.17fF
C10588 a_14010_9158# col[11] 0.38fF
C10589 a_2275_8178# a_14922_8154# 0.17fF
C10590 a_34090_17190# m2_33860_18014# 0.84fF
C10591 a_9994_14178# ctop 4.91fF
C10592 vcm col_n[7] 3.22fF
C10593 VDD col_n[10] 13.96fF
C10594 a_2966_13174# a_2966_12170# 0.84fF
C10595 ctop rowoff_n[15] 0.28fF
C10596 a_29070_5142# col_n[26] 0.34fF
C10597 a_2275_11190# col[7] 0.17fF
C10598 a_24962_14178# vcm 0.18fF
C10599 m2_1732_8978# rowon_n[7] 0.43fF
C10600 a_21038_4138# VDD 2.58fF
C10601 a_2475_5166# a_6982_5142# 0.68fF
C10602 a_3970_5142# a_4974_5142# 0.86fF
C10603 a_9294_9198# col_n[6] 0.11fF
C10604 a_2275_10186# a_29982_10162# 0.17fF
C10605 a_2475_10186# col[27] 0.22fF
C10606 a_3970_9158# rowoff_n[7] 2.57fF
C10607 a_14010_14178# rowon_n[12] 0.45fF
C10608 a_27974_15182# a_28066_15182# 0.45fF
C10609 a_10998_15182# rowoff_n[13] 2.23fF
C10610 m2_34864_10986# VDD 1.59fF
C10611 a_2966_12170# row_n[10] 0.41fF
C10612 a_24050_4138# rowon_n[2] 0.45fF
C10613 a_5886_17190# vcm 0.18fF
C10614 m2_9764_18014# m3_9896_18146# 4.41fF
C10615 a_20034_1126# m3_19936_1078# 3.79fF
C10616 a_2275_16210# rowon_n[14] 1.99fF
C10617 a_2475_7174# VDD 41.96fF
C10618 a_13006_7150# rowoff_n[5] 2.13fF
C10619 a_29070_8154# a_29070_7150# 0.84fF
C10620 a_2475_7174# a_22042_7150# 0.68fF
C10621 m2_2736_946# vcm 0.71fF
C10622 a_7986_2130# vcm 0.89fF
C10623 a_2275_13198# col[24] 0.17fF
C10624 a_22042_5142# rowoff_n[3] 1.69fF
C10625 a_2475_4162# row_n[2] 0.48fF
C10626 a_18026_3134# col_n[15] 0.34fF
C10627 a_2275_2154# col[29] 0.17fF
C10628 a_2275_4162# a_13006_4138# 0.71fF
C10629 a_28066_15182# col_n[25] 0.34fF
C10630 a_17022_11166# VDD 2.99fF
C10631 a_2966_17190# m2_2736_18014# 0.84fF
C10632 a_19030_9158# a_20034_9158# 0.86fF
C10633 a_35002_17190# rowon_n[15] 0.14fF
C10634 a_31078_3134# rowoff_n[1] 1.25fF
C10635 a_23046_6146# vcm 0.89fF
C10636 a_8898_18194# a_8990_18194# 0.11fF
C10637 a_2475_1150# a_5886_1126# 0.41fF
C10638 a_2275_1150# a_3270_1166# 0.15fF
C10639 a_2475_13198# m2_34864_12994# 0.56fF
C10640 a_2275_6170# a_28066_6146# 0.71fF
C10641 a_32082_15182# VDD 1.44fF
C10642 a_9994_11166# a_9994_10162# 0.84fF
C10643 m2_28840_18014# vcm 0.71fF
C10644 a_2275_15206# a_6890_15182# 0.17fF
C10645 a_22042_11166# rowon_n[9] 0.45fF
C10646 a_3970_9158# vcm 0.89fF
C10647 col_n[16] rowoff_n[5] 0.22fF
C10648 col_n[19] rowoff_n[8] 0.20fF
C10649 col_n[12] rowoff_n[1] 0.25fF
C10650 col_n[15] rowoff_n[4] 0.23fF
C10651 col_n[18] rowoff_n[7] 0.21fF
C10652 col_n[13] rowoff_n[2] 0.24fF
C10653 col_n[20] rowoff_n[9] 0.19fF
C10654 col_n[17] rowoff_n[6] 0.21fF
C10655 col_n[14] rowoff_n[3] 0.24fF
C10656 col_n[11] rowoff_n[0] 0.26fF
C10657 a_2475_6170# col[4] 0.22fF
C10658 a_2275_3158# a_18330_3174# 0.15fF
C10659 a_2475_3158# a_20946_3134# 0.41fF
C10660 a_2475_1150# m2_21812_946# 0.62fF
C10661 a_33390_2170# col_n[30] 0.11fF
C10662 m3_21944_1078# ctop 0.21fF
C10663 a_15014_16186# m2_15212_16434# 0.19fF
C10664 a_17022_13174# col_n[14] 0.34fF
C10665 a_2275_12194# col_n[11] 0.17fF
C10666 a_28370_4178# vcm 0.24fF
C10667 m2_20808_946# col_n[18] 0.45fF
C10668 a_23958_11166# rowoff_n[9] 0.50fF
C10669 a_2275_17214# a_21950_17190# 0.17fF
C10670 a_2275_1150# col_n[16] 0.14fF
C10671 a_19030_13174# vcm 0.89fF
C10672 a_15926_3134# VDD 0.29fF
C10673 a_18938_5142# a_19030_5142# 0.45fF
C10674 a_34090_12170# m2_34288_12418# 0.19fF
C10675 a_2275_5166# a_33390_5182# 0.15fF
C10676 a_9902_5142# rowon_n[3] 0.14fF
C10677 a_2275_18218# a_31990_18194# 0.17fF
C10678 a_2275_9182# col[1] 0.17fF
C10679 col[21] rowoff_n[14] 0.21fF
C10680 a_32994_9158# rowoff_n[7] 0.40fF
C10681 a_2475_14202# a_14010_14178# 0.68fF
C10682 a_25054_15182# a_25054_14178# 0.84fF
C10683 col_n[4] rowoff_n[10] 0.31fF
C10684 a_9294_7190# vcm 0.24fF
C10685 a_2275_2154# a_26970_2130# 0.17fF
C10686 a_22042_2130# ctop 4.93fF
C10687 a_34090_17190# vcm 0.89fF
C10688 a_2475_8178# col[21] 0.22fF
C10689 a_30986_7150# VDD 0.29fF
C10690 a_5978_14178# m2_6176_14426# 0.19fF
C10691 a_3878_11166# a_3970_11166# 0.45fF
C10692 a_2275_11190# a_4974_11166# 0.71fF
C10693 a_32386_12210# col_n[29] 0.11fF
C10694 a_5978_11166# col_n[3] 0.34fF
C10695 a_2475_16210# a_29070_16186# 0.68fF
C10696 a_15014_16186# a_16018_16186# 0.86fF
C10697 a_2275_14202# col_n[28] 0.17fF
C10698 a_24354_11206# vcm 0.24fF
C10699 a_22442_1488# VDD 0.14fF
C10700 a_30074_8154# rowon_n[6] 0.45fF
C10701 a_25054_10162# m2_25252_10410# 0.19fF
C10702 a_11910_10162# VDD 0.29fF
C10703 VDD col_n[21] 11.23fF
C10704 vcm col_n[18] 3.22fF
C10705 col[5] rowoff_n[15] 0.31fF
C10706 a_33998_9158# a_34090_9158# 0.45fF
C10707 a_2275_11190# col[18] 0.17fF
C10708 a_2275_13198# a_20034_13174# 0.71fF
C10709 a_17934_5142# vcm 0.18fF
C10710 a_11910_12170# rowoff_n[10] 0.64fF
C10711 a_2275_18218# m2_12776_18014# 0.51fF
C10712 a_26058_10162# col[23] 0.38fF
C10713 a_7986_8154# row_n[6] 0.43fF
C10714 a_5278_14218# vcm 0.24fF
C10715 a_2966_4138# VDD 4.45fF
C10716 a_7894_12170# rowon_n[10] 0.14fF
C10717 a_18026_9158# ctop 4.91fF
C10718 a_26970_14178# VDD 0.29fF
C10719 a_2275_10186# a_10298_10202# 0.15fF
C10720 a_2475_10186# a_12914_10162# 0.41fF
C10721 a_17934_2130# rowon_n[0] 0.14fF
C10722 m2_1732_17010# sample_n 0.12fF
C10723 a_2275_15206# a_35094_15182# 0.14fF
C10724 a_21342_10202# col_n[18] 0.11fF
C10725 a_32994_9158# vcm 0.18fF
C10726 a_27974_16186# rowoff_n[14] 0.46fF
C10727 a_25054_3134# a_26058_3134# 0.86fF
C10728 a_16018_8154# m2_16216_8402# 0.19fF
C10729 a_20338_18234# vcm 0.25fF
C10730 a_27974_1126# m2_27836_946# 0.31fF
C10731 a_2874_7150# a_2966_7150# 0.45fF
C10732 a_33086_13174# ctop 4.91fF
C10733 a_7894_17190# VDD 0.29fF
C10734 a_14922_12170# a_15014_12170# 0.45fF
C10735 a_2475_12194# a_27974_12170# 0.41fF
C10736 a_2275_12194# a_25358_12210# 0.15fF
C10737 a_28066_15182# rowon_n[13] 0.45fF
C10738 a_13918_12170# vcm 0.18fF
C10739 a_9994_2130# VDD 3.71fF
C10740 a_16018_5142# a_16018_4138# 0.84fF
C10741 a_15014_8154# col[12] 0.38fF
C10742 m2_15788_946# m3_15920_1078# 4.41fF
C10743 a_2275_10186# col_n[5] 0.17fF
C10744 a_2275_9182# a_18938_9158# 0.17fF
C10745 a_14010_16186# ctop 4.91fF
C10746 a_30074_4138# col_n[27] 0.34fF
C10747 a_5978_15182# row_n[13] 0.43fF
C10748 a_6982_6146# m2_7180_6394# 0.19fF
C10749 a_10298_8194# col_n[7] 0.11fF
C10750 a_28978_16186# vcm 0.18fF
C10751 a_25054_6146# VDD 2.16fF
C10752 a_16018_5142# row_n[3] 0.43fF
C10753 a_5978_6146# a_6982_6146# 0.86fF
C10754 a_2475_6170# a_10998_6146# 0.68fF
C10755 a_15926_9158# rowon_n[7] 0.14fF
C10756 a_4974_8154# rowoff_n[6] 2.52fF
C10757 a_2275_11190# a_33998_11166# 0.17fF
C10758 a_2475_17214# col[10] 0.22fF
C10759 col_n[31] rowoff_n[9] 0.11fF
C10760 col_n[24] rowoff_n[2] 0.16fF
C10761 col_n[27] rowoff_n[5] 0.14fF
C10762 col_n[30] rowoff_n[8] 0.12fF
C10763 col_n[25] rowoff_n[3] 0.16fF
C10764 col_n[28] rowoff_n[6] 0.14fF
C10765 col_n[22] rowoff_n[0] 0.18fF
C10766 a_31078_1126# vcm 0.15fF
C10767 col_n[29] rowoff_n[7] 0.13fF
C10768 col_n[26] rowoff_n[4] 0.15fF
C10769 col_n[23] rowoff_n[1] 0.17fF
C10770 a_29982_16186# a_30074_16186# 0.45fF
C10771 a_2475_6170# col[15] 0.22fF
C10772 m2_1732_12994# m2_1732_11990# 0.84fF
C10773 a_15926_17190# rowoff_n[15] 0.59fF
C10774 m2_32856_18014# VDD 2.13fF
C10775 a_14010_6146# rowoff_n[4] 2.08fF
C10776 a_1957_3158# a_2161_3158# 0.11fF
C10777 a_2475_3158# a_2275_3158# 2.96fF
C10778 m3_17928_18146# ctop 0.21fF
C10779 a_5978_9158# VDD 4.13fF
C10780 a_31078_9158# a_31078_8154# 0.84fF
C10781 a_2475_8178# a_26058_8154# 0.68fF
C10782 a_3970_6146# col[1] 0.38fF
C10783 a_2275_12194# col_n[22] 0.17fF
C10784 a_2275_1150# col_n[27] 0.17fF
C10785 a_12002_4138# vcm 0.89fF
C10786 a_2874_3134# rowon_n[1] 0.14fF
C10787 a_23046_4138# rowoff_n[2] 1.64fF
C10788 a_2475_17214# a_4882_17190# 0.41fF
C10789 a_2275_17214# a_3878_17190# 0.17fF
C10790 a_19030_2130# col_n[16] 0.33fF
C10791 a_29070_14178# col_n[26] 0.34fF
C10792 a_2275_5166# a_17022_5142# 0.71fF
C10793 a_2275_9182# col[12] 0.17fF
C10794 sample_n rowoff_n[14] 0.55fF
C10795 a_21038_13174# VDD 2.58fF
C10796 a_2275_18218# a_12306_18234# 0.15fF
C10797 a_9294_18234# col_n[6] 0.11fF
C10798 a_21038_10162# a_22042_10162# 0.86fF
C10799 a_32082_2130# rowoff_n[0] 1.20fF
C10800 col_n[15] rowoff_n[10] 0.23fF
C10801 m2_34864_11990# vcm 0.72fF
C10802 a_27062_8154# vcm 0.89fF
C10803 a_14010_12170# row_n[10] 0.43fF
C10804 a_2275_2154# a_7286_2170# 0.15fF
C10805 a_2475_2154# a_9902_2130# 0.41fF
C10806 a_5886_2130# a_5978_2130# 0.45fF
C10807 a_13918_16186# rowon_n[14] 0.14fF
C10808 a_2275_7174# a_32082_7150# 0.71fF
C10809 a_24050_2130# row_n[0] 0.43fF
C10810 a_2475_16210# VDD 41.96fF
C10811 a_12002_12170# a_12002_11166# 0.84fF
C10812 a_2275_14202# row_n[12] 26.41fF
C10813 a_23958_6146# rowon_n[4] 0.14fF
C10814 a_17326_2170# vcm 0.24fF
C10815 a_2275_16210# a_10906_16186# 0.17fF
C10816 a_7986_11166# vcm 0.89fF
C10817 VDD rowon_n[15] 4.68fF
C10818 vcm col_n[29] 3.22fF
C10819 a_4882_1126# VDD 0.99fF
C10820 col[16] rowoff_n[15] 0.24fF
C10821 a_2275_4162# a_22346_4178# 0.15fF
C10822 a_2475_4162# a_24962_4138# 0.41fF
C10823 a_18026_12170# col_n[15] 0.34fF
C10824 a_2275_11190# col[29] 0.17fF
C10825 col_n[0] rowoff_n[11] 0.34fF
C10826 a_2475_13198# a_2874_13174# 0.41fF
C10827 a_1957_13198# a_2275_13198# 0.19fF
C10828 a_24962_10162# rowoff_n[8] 0.49fF
C10829 a_32386_6186# vcm 0.24fF
C10830 a_28066_13174# rowoff_n[11] 1.40fF
C10831 a_2275_8178# col_n[0] 0.17fF
C10832 a_2275_1150# a_15926_1126# 0.17fF
C10833 a_23046_15182# vcm 0.89fF
C10834 a_19942_5142# VDD 0.29fF
C10835 a_20946_6146# a_21038_6146# 0.45fF
C10836 a_33998_8154# rowoff_n[6] 0.39fF
C10837 a_27062_16186# a_27062_15182# 0.84fF
C10838 a_2475_15206# a_18026_15182# 0.68fF
C10839 m2_1732_2954# sample 0.31fF
C10840 a_13310_9198# vcm 0.24fF
C10841 m2_1732_13998# VDD 5.46fF
C10842 a_2275_3158# a_30986_3134# 0.17fF
C10843 a_2475_8178# m2_1732_7974# 0.16fF
C10844 a_26058_4138# ctop 4.91fF
C10845 a_3970_18194# vcm 0.15fF
C10846 a_35002_9158# VDD 0.36fF
C10847 a_22042_9158# row_n[7] 0.43fF
C10848 a_2475_15206# col[4] 0.22fF
C10849 a_21950_13174# rowon_n[11] 0.14fF
C10850 a_2475_4162# col[9] 0.22fF
C10851 a_6982_10162# col_n[4] 0.34fF
C10852 a_33390_11206# col_n[30] 0.11fF
C10853 a_2275_12194# a_8990_12170# 0.71fF
C10854 a_6890_3134# vcm 0.18fF
C10855 a_2475_17214# a_33086_17190# 0.68fF
C10856 a_31990_3134# rowon_n[1] 0.14fF
C10857 a_17022_17190# a_18026_17190# 0.86fF
C10858 m2_23820_18014# m2_24824_18014# 0.86fF
C10859 a_28370_13214# vcm 0.24fF
C10860 a_2275_10186# col_n[16] 0.17fF
C10861 a_6982_7150# ctop 4.91fF
C10862 a_15926_12170# VDD 0.29fF
C10863 m2_28840_946# m2_29268_1374# 0.19fF
C10864 a_2275_14202# a_24050_14178# 0.71fF
C10865 a_27062_9158# col[24] 0.38fF
C10866 a_2275_7174# col[6] 0.17fF
C10867 a_8990_7150# rowon_n[5] 0.45fF
C10868 a_21950_7150# vcm 0.18fF
C10869 a_16018_14178# rowoff_n[12] 1.98fF
C10870 a_9294_16226# vcm 0.24fF
C10871 a_22042_11166# ctop 4.91fF
C10872 a_2475_17214# col[21] 0.22fF
C10873 a_30986_16186# VDD 0.29fF
C10874 a_2475_6170# col[26] 0.22fF
C10875 a_2475_11190# a_16930_11166# 0.41fF
C10876 a_2275_11190# a_14314_11206# 0.15fF
C10877 a_22346_9198# col_n[19] 0.11fF
C10878 a_20034_16186# row_n[14] 0.43fF
C10879 a_27062_4138# a_28066_4138# 0.86fF
C10880 a_2275_8178# a_7894_8154# 0.17fF
C10881 a_21038_17190# m2_21236_17438# 0.19fF
C10882 a_30074_6146# row_n[4] 0.43fF
C10883 a_29982_10162# rowon_n[8] 0.14fF
C10884 a_16930_13174# a_17022_13174# 0.45fF
C10885 a_2475_13198# a_31990_13174# 0.41fF
C10886 a_2275_13198# a_29374_13214# 0.15fF
C10887 a_2275_9182# col[23] 0.17fF
C10888 a_16018_7150# col[13] 0.38fF
C10889 a_17934_14178# vcm 0.18fF
C10890 a_14010_4138# VDD 3.30fF
C10891 a_18026_6146# a_18026_5142# 0.84fF
C10892 col_n[26] rowoff_n[10] 0.15fF
C10893 a_2966_13174# VDD 4.45fF
C10894 a_2275_10186# a_22954_10162# 0.17fF
C10895 a_31078_3134# col_n[28] 0.34fF
C10896 a_6982_14178# rowon_n[12] 0.45fF
C10897 a_11302_7190# col_n[8] 0.11fF
C10898 a_3970_15182# rowoff_n[13] 2.57fF
C10899 a_17022_4138# rowon_n[2] 0.45fF
C10900 a_32994_18194# vcm 0.18fF
C10901 a_29070_8154# VDD 1.75fF
C10902 a_5978_7150# rowoff_n[5] 2.47fF
C10903 a_7986_7150# a_8990_7150# 0.86fF
C10904 a_2475_7174# a_15014_7150# 0.68fF
C10905 a_12002_15182# m2_12200_15430# 0.19fF
C10906 a_35094_3134# vcm 0.15fF
C10907 vcm rowon_n[11] 0.91fF
C10908 col_n[8] rowon_n[15] 0.17fF
C10909 sample rowon_n[10] 0.10fF
C10910 col_n[0] row_n[11] 0.37fF
C10911 col_n[2] rowon_n[12] 0.17fF
C10912 col_n[3] row_n[13] 0.37fF
C10913 col_n[5] row_n[14] 0.37fF
C10914 col_n[1] row_n[12] 0.37fF
C10915 col_n[7] row_n[15] 0.37fF
C10916 col_n[4] rowon_n[13] 0.17fF
C10917 VDD row_n[10] 4.64fF
C10918 col_n[6] rowon_n[14] 0.17fF
C10919 a_31990_17190# a_32082_17190# 0.45fF
C10920 col[27] rowoff_n[15] 0.17fF
C10921 a_2275_3158# m2_34864_2954# 0.51fF
C10922 a_15014_5142# rowoff_n[3] 2.03fF
C10923 a_2475_2154# col[3] 0.22fF
C10924 col_n[10] rowoff_n[11] 0.27fF
C10925 a_2275_4162# a_5978_4138# 0.71fF
C10926 a_31078_11166# m2_31276_11414# 0.19fF
C10927 a_28066_13174# row_n[11] 0.43fF
C10928 a_4974_5142# col[2] 0.38fF
C10929 a_9994_11166# VDD 3.71fF
C10930 a_15014_17190# col[12] 0.38fF
C10931 a_27974_17190# rowon_n[15] 0.14fF
C10932 a_2475_9182# a_30074_9158# 0.68fF
C10933 a_33086_10162# a_33086_9158# 0.84fF
C10934 a_24050_3134# rowoff_n[1] 1.59fF
C10935 a_2275_8178# col_n[10] 0.17fF
C10936 a_20034_1126# col_n[17] 0.39fF
C10937 a_16018_6146# vcm 0.89fF
C10938 a_30074_13174# col_n[27] 0.34fF
C10939 a_35398_6186# VDD 0.12fF
C10940 a_2275_6170# a_21038_6146# 0.71fF
C10941 a_10298_17230# col_n[7] 0.11fF
C10942 a_25054_15182# VDD 2.16fF
C10943 a_2275_5166# col[0] 0.16fF
C10944 a_23046_11166# a_24050_11166# 0.86fF
C10945 m2_34864_1950# vcm 0.73fF
C10946 m2_14784_18014# vcm 0.71fF
C10947 a_15014_11166# rowon_n[9] 0.45fF
C10948 a_31078_10162# vcm 0.89fF
C10949 a_2475_15206# col[15] 0.22fF
C10950 a_7894_3134# a_7986_3134# 0.45fF
C10951 a_2275_3158# a_11302_3174# 0.15fF
C10952 a_2475_3158# a_13918_3134# 0.41fF
C10953 a_22042_9158# m2_22240_9406# 0.19fF
C10954 a_2475_4162# col[20] 0.22fF
C10955 a_2275_1150# m2_4744_946# 0.51fF
C10956 m3_34996_5094# ctop 0.22fF
C10957 a_3878_13174# rowon_n[11] 0.14fF
C10958 a_14010_13174# a_14010_12170# 0.84fF
C10959 a_3970_15182# col[1] 0.38fF
C10960 a_21342_4178# vcm 0.24fF
C10961 a_16930_11166# rowoff_n[9] 0.58fF
C10962 a_2275_10186# col_n[27] 0.17fF
C10963 a_2275_17214# a_14922_17190# 0.17fF
C10964 a_12002_13174# vcm 0.89fF
C10965 a_19030_11166# col_n[16] 0.34fF
C10966 a_8898_3134# VDD 0.29fF
C10967 a_2275_5166# a_26362_5182# 0.15fF
C10968 a_2475_5166# a_28978_5142# 0.41fF
C10969 a_2275_18218# a_24962_18194# 0.17fF
C10970 a_25966_9158# rowoff_n[7] 0.48fF
C10971 a_2275_7174# col[17] 0.17fF
C10972 a_2475_14202# a_6982_14178# 0.68fF
C10973 a_3970_14178# a_4974_14178# 0.86fF
C10974 a_3878_7150# vcm 0.18fF
C10975 a_32994_15182# rowoff_n[13] 0.40fF
C10976 a_2275_2154# a_19942_2130# 0.17fF
C10977 a_13006_7150# m2_13204_7398# 0.19fF
C10978 a_15014_2130# ctop 4.93fF
C10979 a_27062_17190# vcm 0.89fF
C10980 rowon_n[6] rowoff_n[6] 20.66fF
C10981 a_23958_7150# VDD 0.29fF
C10982 a_35002_7150# rowoff_n[5] 0.38fF
C10983 a_22954_7150# a_23046_7150# 0.45fF
C10984 a_2874_18194# vcm 0.18fF
C10985 m2_4744_946# col_n[2] 0.45fF
C10986 a_29982_2130# vcm 0.18fF
C10987 a_29070_17190# a_29070_16186# 0.84fF
C10988 a_2475_16210# a_22042_16186# 0.68fF
C10989 a_32082_3134# m2_32280_3382# 0.19fF
C10990 a_17326_11206# vcm 0.24fF
C10991 a_15414_1488# VDD 0.16fF
C10992 a_1957_16210# row_n[14] 0.29fF
C10993 a_23046_8154# rowon_n[6] 0.45fF
C10994 a_2275_4162# a_35002_4138# 0.17fF
C10995 a_30074_6146# ctop 4.91fF
C10996 a_4882_10162# VDD 0.29fF
C10997 a_7986_9158# col_n[5] 0.34fF
C10998 m3_34568_1078# m3_34996_1078# 0.21fF
C10999 a_2275_13198# a_13006_13174# 0.71fF
C11000 a_10906_5142# vcm 0.18fF
C11001 a_4882_12170# rowoff_n[10] 0.72fF
C11002 m2_24248_2378# a_24050_2130# 0.19fF
C11003 a_3970_5142# m2_4168_5390# 0.19fF
C11004 a_32386_15222# vcm 0.24fF
C11005 a_2275_17214# col_n[0] 0.17fF
C11006 a_34090_17190# row_n[15] 0.43fF
C11007 a_10998_9158# ctop 4.91fF
C11008 a_2275_6170# col_n[4] 0.17fF
C11009 a_19942_14178# VDD 0.29fF
C11010 a_2475_10186# a_5886_10162# 0.41fF
C11011 a_2275_10186# a_3270_10202# 0.15fF
C11012 a_10906_2130# rowon_n[0] 0.14fF
C11013 m2_1732_15002# vcm 1.11fF
C11014 a_28066_8154# col[25] 0.38fF
C11015 a_2275_15206# a_28066_15182# 0.71fF
C11016 a_25966_9158# vcm 0.18fF
C11017 a_20946_16186# rowoff_n[14] 0.54fF
C11018 a_4974_3134# a_4974_2130# 0.84fF
C11019 a_2275_3158# ctop 0.14fF
C11020 a_13310_18234# vcm 0.25fF
C11021 a_26058_13174# ctop 4.91fF
C11022 a_35002_18194# VDD 0.56fF
C11023 col_n[1] rowon_n[6] 0.17fF
C11024 col_n[14] row_n[13] 0.37fF
C11025 col_n[0] rowon_n[5] 0.17fF
C11026 col_n[13] rowon_n[12] 0.17fF
C11027 col_n[9] rowon_n[10] 0.17fF
C11028 col_n[7] rowon_n[9] 0.17fF
C11029 col_n[2] row_n[7] 0.37fF
C11030 col_n[18] row_n[15] 0.37fF
C11031 col_n[16] row_n[14] 0.37fF
C11032 col_n[10] row_n[11] 0.37fF
C11033 VDD rowon_n[4] 4.61fF
C11034 col_n[4] row_n[8] 0.37fF
C11035 sample row_n[5] 0.92fF
C11036 col_n[15] rowon_n[13] 0.17fF
C11037 col_n[6] row_n[9] 0.37fF
C11038 vcm row_n[6] 1.08fF
C11039 col_n[17] rowon_n[14] 0.17fF
C11040 col_n[8] row_n[10] 0.37fF
C11041 col_n[19] rowon_n[15] 0.17fF
C11042 col_n[3] rowon_n[7] 0.17fF
C11043 col_n[11] rowon_n[11] 0.17fF
C11044 col_n[12] row_n[12] 0.37fF
C11045 col_n[5] rowon_n[8] 0.17fF
C11046 a_23350_8194# col_n[20] 0.11fF
C11047 a_2475_12194# a_20946_12170# 0.41fF
C11048 a_2275_12194# a_18330_12210# 0.15fF
C11049 a_2475_13198# col[9] 0.22fF
C11050 a_2475_2154# col[14] 0.22fF
C11051 col_n[21] rowoff_n[11] 0.19fF
C11052 a_21038_15182# rowon_n[13] 0.45fF
C11053 m2_34864_18014# m2_35292_18442# 0.19fF
C11054 a_6890_12170# vcm 0.18fF
C11055 a_2874_2130# VDD 0.29fF
C11056 a_29070_5142# a_30074_5142# 0.86fF
C11057 a_31078_5142# rowon_n[3] 0.45fF
C11058 a_2275_9182# a_11910_9158# 0.17fF
C11059 a_6982_16186# ctop 4.91fF
C11060 a_2275_8178# col_n[21] 0.17fF
C11061 a_2475_18218# m2_24824_18014# 0.62fF
C11062 a_2275_14202# a_33390_14218# 0.15fF
C11063 a_18938_14178# a_19030_14178# 0.45fF
C11064 a_17022_6146# col[14] 0.38fF
C11065 a_2275_16210# col[6] 0.17fF
C11066 a_21950_16186# vcm 0.18fF
C11067 a_18026_6146# VDD 2.89fF
C11068 a_2275_5166# col[11] 0.17fF
C11069 a_8990_5142# row_n[3] 0.43fF
C11070 a_20034_7150# a_20034_6146# 0.84fF
C11071 a_2475_6170# a_3970_6146# 0.68fF
C11072 a_2275_6170# a_2966_6146# 0.67fF
C11073 a_32082_2130# col_n[29] 0.34fF
C11074 a_8898_9158# rowon_n[7] 0.14fF
C11075 a_2275_11190# a_26970_11166# 0.17fF
C11076 col_n[5] rowoff_n[12] 0.30fF
C11077 a_24050_1126# vcm 0.15fF
C11078 m2_16792_18014# col[14] 0.37fF
C11079 a_2475_15206# col[26] 0.22fF
C11080 a_12306_6186# col_n[9] 0.11fF
C11081 a_2475_4162# col[31] 0.22fF
C11082 a_22346_18234# col_n[19] 0.11fF
C11083 a_8898_17190# rowoff_n[15] 0.67fF
C11084 m2_18800_18014# VDD 3.67fF
C11085 a_6982_6146# rowoff_n[4] 2.42fF
C11086 a_33086_10162# VDD 1.34fF
C11087 a_9994_8154# a_10998_8154# 0.86fF
C11088 a_2475_8178# a_19030_8154# 0.68fF
C11089 a_4974_4138# vcm 0.89fF
C11090 a_33998_18194# a_34090_18194# 0.11fF
C11091 a_33086_12170# rowoff_n[10] 1.15fF
C11092 a_16018_4138# rowoff_n[2] 1.98fF
C11093 a_28978_1126# a_29070_1126# 0.11fF
C11094 a_5978_4138# col[3] 0.38fF
C11095 a_29070_12170# rowon_n[10] 0.45fF
C11096 a_2275_5166# a_9994_5142# 0.71fF
C11097 a_16018_16186# col[13] 0.38fF
C11098 a_2275_7174# col[28] 0.17fF
C11099 a_14010_13174# VDD 3.30fF
C11100 a_2275_18218# a_5278_18234# 0.15fF
C11101 a_2475_10186# a_34090_10162# 0.68fF
C11102 a_25054_2130# rowoff_n[0] 1.54fF
C11103 a_31078_12170# col_n[28] 0.34fF
C11104 a_20034_8154# vcm 0.89fF
C11105 a_6982_12170# row_n[10] 0.43fF
C11106 m2_14784_18014# m3_14916_18146# 4.43fF
C11107 a_11302_16226# col_n[8] 0.11fF
C11108 a_6890_16186# rowon_n[14] 0.14fF
C11109 m2_32856_18014# col_n[30] 0.33fF
C11110 a_2275_7174# a_25054_7150# 0.71fF
C11111 a_29070_17190# VDD 1.75fF
C11112 a_17022_2130# row_n[0] 0.43fF
C11113 a_25054_12170# a_26058_12170# 0.86fF
C11114 a_16930_6146# rowon_n[4] 0.14fF
C11115 a_10298_2170# vcm 0.24fF
C11116 a_2874_16186# a_2966_16186# 0.45fF
C11117 a_35094_12170# vcm 0.15fF
C11118 a_31990_2130# VDD 0.29fF
C11119 a_9902_4138# a_9994_4138# 0.45fF
C11120 a_2275_4162# a_15318_4178# 0.15fF
C11121 a_2475_4162# a_17934_4138# 0.41fF
C11122 a_2475_11190# col[3] 0.22fF
C11123 a_4974_14178# col[2] 0.38fF
C11124 a_16018_14178# a_16018_13174# 0.84fF
C11125 a_17934_10162# rowoff_n[8] 0.57fF
C11126 a_25358_6186# vcm 0.24fF
C11127 a_21038_13174# rowoff_n[11] 1.74fF
C11128 a_2275_17214# col_n[10] 0.17fF
C11129 a_20034_10162# col_n[17] 0.34fF
C11130 a_2275_1150# a_8898_1126# 0.17fF
C11131 a_16018_15182# vcm 0.89fF
C11132 a_2275_6170# col_n[15] 0.17fF
C11133 a_12914_5142# VDD 0.29fF
C11134 a_2475_6170# a_32994_6146# 0.41fF
C11135 a_2275_6170# a_30378_6186# 0.15fF
C11136 a_26970_8154# rowoff_n[6] 0.47fF
C11137 a_35398_15222# VDD 0.12fF
C11138 a_5978_15182# a_6982_15182# 0.86fF
C11139 a_2475_15206# a_10998_15182# 0.68fF
C11140 a_2275_14202# col[0] 0.16fF
C11141 a_2275_3158# col[5] 0.17fF
C11142 a_6282_9198# vcm 0.24fF
C11143 a_2275_16210# rowoff_n[14] 0.81fF
C11144 a_2275_3158# a_23958_3134# 0.17fF
C11145 a_19030_4138# ctop 4.91fF
C11146 a_2275_1150# m2_27836_946# 0.51fF
C11147 a_10906_1126# m2_10768_946# 0.31fF
C11148 col_n[8] rowon_n[4] 0.17fF
C11149 col_n[15] row_n[8] 0.37fF
C11150 VDD sw_n 0.58fF
C11151 vcm rowon_n[0] 0.91fF
C11152 col_n[21] row_n[11] 0.37fF
C11153 col_n[6] rowon_n[3] 0.17fF
C11154 col_n[13] row_n[7] 0.37fF
C11155 col_n[4] rowon_n[2] 0.17fF
C11156 col_n[29] row_n[15] 0.37fF
C11157 col_n[11] row_n[6] 0.37fF
C11158 col_n[2] rowon_n[1] 0.17fF
C11159 col_n[27] row_n[14] 0.37fF
C11160 col_n[9] row_n[5] 0.37fF
C11161 col_n[25] row_n[13] 0.37fF
C11162 col_n[7] row_n[4] 0.37fF
C11163 col_n[5] row_n[3] 0.37fF
C11164 col_n[12] rowon_n[6] 0.17fF
C11165 col_n[19] row_n[10] 0.37fF
C11166 col_n[28] rowon_n[14] 0.17fF
C11167 col_n[10] rowon_n[5] 0.17fF
C11168 col_n[17] row_n[9] 0.37fF
C11169 col_n[1] row_n[1] 0.37fF
C11170 col_n[26] rowon_n[13] 0.17fF
C11171 col_n[0] row_n[0] 0.37fF
C11172 col_n[30] rowon_n[15] 0.17fF
C11173 col_n[14] rowon_n[7] 0.17fF
C11174 col_n[22] rowon_n[11] 0.17fF
C11175 col_n[23] row_n[12] 0.37fF
C11176 col_n[16] rowon_n[8] 0.17fF
C11177 col_n[18] rowon_n[9] 0.17fF
C11178 col_n[20] rowon_n[10] 0.17fF
C11179 col_n[3] row_n[2] 0.37fF
C11180 col_n[24] rowon_n[12] 0.17fF
C11181 a_27974_9158# VDD 0.29fF
C11182 a_15014_9158# row_n[7] 0.43fF
C11183 a_18026_16186# m2_18224_16434# 0.19fF
C11184 a_24962_8154# a_25054_8154# 0.45fF
C11185 a_14922_13174# rowon_n[11] 0.14fF
C11186 a_2475_13198# col[20] 0.22fF
C11187 a_2475_2154# col[25] 0.22fF
C11188 a_1957_12194# a_2161_12194# 0.11fF
C11189 a_2475_12194# a_2275_12194# 2.96fF
C11190 m2_1732_4962# rowoff_n[3] 2.46fF
C11191 a_33998_4138# vcm 0.18fF
C11192 a_24962_3134# rowon_n[1] 0.14fF
C11193 a_2475_17214# a_26058_17190# 0.68fF
C11194 a_2966_15182# rowon_n[13] 0.45fF
C11195 m2_16792_18014# m2_17796_18014# 0.86fF
C11196 a_21342_13214# vcm 0.24fF
C11197 a_8990_8154# col_n[6] 0.34fF
C11198 a_34090_8154# ctop 4.80fF
C11199 a_8898_12170# VDD 0.29fF
C11200 m2_21812_946# m2_22240_1374# 0.19fF
C11201 a_2275_14202# a_17022_14178# 0.71fF
C11202 a_2275_16210# col[17] 0.17fF
C11203 a_2475_7174# rowon_n[5] 0.40fF
C11204 a_14922_7150# vcm 0.18fF
C11205 a_8990_14178# rowoff_n[12] 2.33fF
C11206 a_2275_5166# col[22] 0.17fF
C11207 a_16018_2130# a_17022_2130# 0.86fF
C11208 a_2475_2154# a_31078_2130# 0.68fF
C11209 a_3878_16186# vcm 0.18fF
C11210 a_8990_14178# m2_9188_14426# 0.19fF
C11211 a_15014_11166# ctop 4.91fF
C11212 col_n[16] rowoff_n[12] 0.22fF
C11213 a_23958_16186# VDD 0.29fF
C11214 a_29070_7150# col[26] 0.38fF
C11215 a_2475_11190# a_9902_11166# 0.41fF
C11216 a_2275_11190# a_7286_11206# 0.15fF
C11217 a_5886_11166# a_5978_11166# 0.45fF
C11218 a_2275_16210# a_32082_16186# 0.71fF
C11219 a_5978_2130# m2_6176_2378# 0.19fF
C11220 a_29982_11166# vcm 0.18fF
C11221 a_13006_16186# row_n[14] 0.43fF
C11222 a_6982_4138# a_6982_3134# 0.84fF
C11223 a_28066_10162# m2_28264_10410# 0.19fF
C11224 a_30074_15182# ctop 4.91fF
C11225 a_24354_7190# col_n[21] 0.11fF
C11226 a_23046_6146# row_n[4] 0.43fF
C11227 a_22954_10162# rowon_n[8] 0.14fF
C11228 a_2275_13198# a_22346_13214# 0.15fF
C11229 a_2475_13198# a_24962_13174# 0.41fF
C11230 a_19030_1126# a_19334_1166# 0.10fF
C11231 a_10906_14178# vcm 0.18fF
C11232 a_6982_4138# VDD 4.02fF
C11233 a_31078_6146# a_32082_6146# 0.86fF
C11234 vcm rowoff_n[13] 2.43fF
C11235 a_2275_10186# a_15926_10162# 0.17fF
C11236 col[0] rowoff_n[6] 0.34fF
C11237 col[1] rowoff_n[7] 0.34fF
C11238 col[2] rowoff_n[8] 0.33fF
C11239 col[3] rowoff_n[9] 0.33fF
C11240 ctop rowoff_n[0] 0.27fF
C11241 a_2275_15206# col_n[4] 0.17fF
C11242 a_20946_15182# a_21038_15182# 0.45fF
C11243 a_2275_4162# col_n[9] 0.17fF
C11244 a_18026_5142# col[15] 0.38fF
C11245 a_1957_8178# vcm 0.16fF
C11246 a_28066_17190# col[25] 0.38fF
C11247 a_9994_4138# rowon_n[2] 0.45fF
C11248 a_19030_8154# m2_19228_8402# 0.19fF
C11249 a_25966_18194# vcm 0.18fF
C11250 a_22042_8154# VDD 2.47fF
C11251 a_2475_7174# a_7986_7150# 0.68fF
C11252 a_22042_8154# a_22042_7150# 0.84fF
C11253 a_2275_12194# ctop 0.14fF
C11254 a_2275_12194# a_30986_12170# 0.17fF
C11255 a_13310_5182# col_n[10] 0.11fF
C11256 a_28066_3134# vcm 0.89fF
C11257 a_23350_17230# col_n[20] 0.11fF
C11258 a_7986_5142# rowoff_n[3] 2.38fF
C11259 a_2475_11190# col[14] 0.22fF
C11260 a_21038_13174# row_n[11] 0.43fF
C11261 a_2874_11166# VDD 0.29fF
C11262 m3_30980_18146# m3_31984_18146# 0.21fF
C11263 m2_21812_946# m3_21944_1078# 4.41fF
C11264 a_2475_9182# a_23046_9158# 0.68fF
C11265 a_20946_17190# rowon_n[15] 0.14fF
C11266 a_12002_9158# a_13006_9158# 0.86fF
C11267 a_31078_3134# row_n[1] 0.43fF
C11268 a_17022_3134# rowoff_n[1] 1.94fF
C11269 a_2275_17214# col_n[21] 0.17fF
C11270 a_30986_7150# rowon_n[5] 0.14fF
C11271 a_8990_6146# vcm 0.89fF
C11272 a_2275_6170# col_n[26] 0.17fF
C11273 a_2966_13174# rowoff_n[11] 2.62fF
C11274 a_2275_18218# col_n[6] 0.17fF
C11275 a_6982_3134# col[4] 0.38fF
C11276 a_30986_2130# a_31078_2130# 0.45fF
C11277 a_9994_6146# m2_10192_6394# 0.19fF
C11278 a_17022_15182# col[14] 0.38fF
C11279 a_2275_6170# a_14010_6146# 0.71fF
C11280 a_18026_15182# VDD 2.89fF
C11281 a_2275_14202# col[11] 0.17fF
C11282 a_1957_18218# VDD 0.59fF
C11283 a_2275_3158# col[16] 0.17fF
C11284 a_32082_11166# col_n[29] 0.34fF
C11285 a_35398_1166# vcm 0.24fF
C11286 a_7986_11166# rowon_n[9] 0.45fF
C11287 a_24050_10162# vcm 0.89fF
C11288 col_n[25] rowon_n[7] 0.17fF
C11289 col_n[23] rowon_n[6] 0.17fF
C11290 col_n[30] row_n[10] 0.37fF
C11291 col_n[21] rowon_n[5] 0.17fF
C11292 col_n[28] row_n[9] 0.37fF
C11293 col_n[19] rowon_n[4] 0.17fF
C11294 col_n[26] row_n[8] 0.37fF
C11295 vcm col[1] 6.67fF
C11296 col_n[17] rowon_n[3] 0.17fF
C11297 col_n[24] row_n[7] 0.37fF
C11298 col_n[15] rowon_n[2] 0.17fF
C11299 col_n[22] row_n[6] 0.37fF
C11300 col_n[29] rowon_n[9] 0.17fF
C11301 rowon_n[13] row_n[13] 21.02fF
C11302 col_n[27] rowon_n[8] 0.17fF
C11303 col_n[10] row_n[0] 0.37fF
C11304 col_n[31] rowon_n[10] 0.17fF
C11305 col_n[12] row_n[1] 0.37fF
C11306 col_n[14] row_n[2] 0.37fF
C11307 col_n[16] row_n[3] 0.37fF
C11308 col_n[18] row_n[4] 0.37fF
C11309 col_n[11] rowon_n[0] 0.17fF
C11310 VDD col[4] 12.44fF
C11311 col_n[20] row_n[5] 0.37fF
C11312 col_n[13] rowon_n[1] 0.17fF
C11313 a_12306_15222# col_n[9] 0.11fF
C11314 a_2475_13198# col[31] 0.22fF
C11315 a_2275_3158# a_4274_3174# 0.15fF
C11316 a_2475_3158# a_6890_3134# 0.41fF
C11317 a_22042_2130# m2_21812_946# 0.84fF
C11318 m3_32988_18146# ctop 0.21fF
C11319 a_2275_8178# a_29070_8154# 0.71fF
C11320 a_27062_13174# a_28066_13174# 0.86fF
C11321 a_14314_4178# vcm 0.24fF
C11322 a_2275_17214# a_7894_17190# 0.17fF
C11323 a_9902_11166# rowoff_n[9] 0.66fF
C11324 a_4974_13174# vcm 0.89fF
C11325 a_11910_5142# a_12002_5142# 0.45fF
C11326 a_2475_5166# a_21950_5142# 0.41fF
C11327 a_2275_5166# a_19334_5182# 0.15fF
C11328 a_5978_13174# col[3] 0.38fF
C11329 a_2275_18218# a_17934_18194# 0.17fF
C11330 a_29070_10162# row_n[8] 0.43fF
C11331 a_18938_9158# rowoff_n[7] 0.56fF
C11332 a_2275_16210# col[28] 0.17fF
C11333 a_28978_14178# rowon_n[12] 0.14fF
C11334 a_18026_15182# a_18026_14178# 0.84fF
C11335 a_21038_9158# col_n[18] 0.34fF
C11336 a_29374_8194# vcm 0.24fF
C11337 a_25966_15182# rowoff_n[13] 0.48fF
C11338 a_2275_2154# a_12914_2130# 0.17fF
C11339 a_20034_17190# vcm 0.89fF
C11340 a_7986_2130# ctop 4.93fF
C11341 col_n[27] rowoff_n[12] 0.14fF
C11342 a_16930_7150# VDD 0.29fF
C11343 a_27974_7150# rowoff_n[5] 0.46fF
C11344 a_2275_7174# a_35398_7190# 0.15fF
C11345 a_2275_2154# col_n[3] 0.17fF
C11346 a_22954_2130# vcm 0.18fF
C11347 a_7986_16186# a_8990_16186# 0.86fF
C11348 a_2475_16210# a_15014_16186# 0.68fF
C11349 a_10298_11206# vcm 0.24fF
C11350 a_8386_1488# VDD 0.17fF
C11351 a_16018_8154# rowon_n[6] 0.45fF
C11352 a_2275_4162# a_27974_4138# 0.17fF
C11353 a_23046_6146# ctop 4.91fF
C11354 a_31990_11166# VDD 0.29fF
C11355 m3_20940_1078# m3_21944_1078# 0.21fF
C11356 a_26970_9158# a_27062_9158# 0.45fF
C11357 a_2275_13198# a_5978_13174# 0.71fF
C11358 a_2475_9182# col[8] 0.22fF
C11359 m2_1732_3958# m2_2160_4386# 0.19fF
C11360 col_n[11] rowoff_n[13] 0.26fF
C11361 a_2475_1150# a_20034_1126# 0.66fF
C11362 a_9994_7150# col_n[7] 0.34fF
C11363 a_25358_15222# vcm 0.24fF
C11364 a_2475_18218# a_30986_18194# 0.41fF
C11365 a_27062_17190# row_n[15] 0.43fF
C11366 a_3970_9158# ctop 4.91fF
C11367 a_2275_15206# col_n[15] 0.17fF
C11368 col[14] rowoff_n[9] 0.25fF
C11369 col[13] rowoff_n[8] 0.26fF
C11370 col[12] rowoff_n[7] 0.27fF
C11371 col[11] rowoff_n[6] 0.27fF
C11372 col[10] rowoff_n[5] 0.28fF
C11373 col[9] rowoff_n[4] 0.29fF
C11374 col[8] rowoff_n[3] 0.29fF
C11375 col[7] rowoff_n[2] 0.30fF
C11376 col[6] rowoff_n[1] 0.31fF
C11377 col[5] rowoff_n[0] 0.31fF
C11378 a_12914_14178# VDD 0.29fF
C11379 a_2275_4162# col_n[20] 0.17fF
C11380 a_2275_15206# a_21038_15182# 0.71fF
C11381 a_18938_9158# vcm 0.18fF
C11382 a_13918_16186# rowoff_n[14] 0.61fF
C11383 a_18026_3134# a_19030_3134# 0.86fF
C11384 a_2275_12194# col[5] 0.17fF
C11385 a_6282_18234# vcm 0.25fF
C11386 a_2275_1150# col[10] 0.17fF
C11387 a_34394_8194# col_n[31] 0.11fF
C11388 a_19030_13174# ctop 4.91fF
C11389 a_30074_6146# col[27] 0.38fF
C11390 a_27974_18194# VDD 0.50fF
C11391 a_2275_12194# a_11302_12210# 0.15fF
C11392 a_2475_12194# a_13918_12170# 0.41fF
C11393 a_7894_12170# a_7986_12170# 0.45fF
C11394 a_2475_11190# col[25] 0.22fF
C11395 a_14010_15182# rowon_n[13] 0.45fF
C11396 m2_27836_18014# m2_28264_18442# 0.19fF
C11397 a_33998_13174# vcm 0.18fF
C11398 a_30074_3134# VDD 1.65fF
C11399 a_8990_5142# a_8990_4138# 0.84fF
C11400 a_2966_13174# row_n[11] 0.41fF
C11401 a_25358_6186# col_n[22] 0.11fF
C11402 a_24050_5142# rowon_n[3] 0.45fF
C11403 a_8990_17190# col_n[6] 0.34fF
C11404 a_2275_17214# rowon_n[15] 1.99fF
C11405 a_4882_18194# m2_4744_18014# 0.34fF
C11406 a_2275_9182# a_4882_9158# 0.17fF
C11407 a_2966_9158# a_3970_9158# 0.86fF
C11408 a_34090_17190# ctop 4.80fF
C11409 a_2475_18218# m2_10768_18014# 0.62fF
C11410 a_2475_14202# a_28978_14178# 0.41fF
C11411 a_2275_14202# a_26362_14218# 0.15fF
C11412 a_2275_18218# col_n[17] 0.17fF
C11413 m2_34864_7974# m2_34864_6970# 0.84fF
C11414 a_14922_16186# vcm 0.18fF
C11415 a_10998_6146# VDD 3.61fF
C11416 a_2275_14202# col[22] 0.17fF
C11417 a_2475_5166# row_n[3] 0.48fF
C11418 a_33086_7150# a_34090_7150# 0.86fF
C11419 a_2275_3158# col[27] 0.17fF
C11420 a_2275_11190# a_19942_11166# 0.17fF
C11421 a_19030_4138# col[16] 0.38fF
C11422 col_n[23] row_n[1] 0.37fF
C11423 col_n[21] row_n[0] 0.37fF
C11424 VDD col[15] 9.72fF
C11425 col_n[6] col[6] 0.50fF
C11426 col_n[27] row_n[3] 0.37fF
C11427 col_n[25] row_n[2] 0.37fF
C11428 vcm col[12] 6.66fF
C11429 col_n[29] row_n[4] 0.37fF
C11430 col_n[22] rowon_n[0] 0.17fF
C11431 a_17022_1126# vcm 0.15fF
C11432 col_n[31] row_n[5] 0.37fF
C11433 col_n[24] rowon_n[1] 0.17fF
C11434 col_n[26] rowon_n[2] 0.17fF
C11435 col_n[28] rowon_n[3] 0.17fF
C11436 col_n[30] rowon_n[4] 0.17fF
C11437 a_22954_16186# a_23046_16186# 0.45fF
C11438 a_29070_16186# col[26] 0.38fF
C11439 m2_4744_18014# VDD 5.01fF
C11440 a_26058_10162# VDD 2.06fF
C11441 a_24050_17190# m2_24248_17438# 0.19fF
C11442 a_2475_8178# a_12002_8154# 0.68fF
C11443 a_24050_9158# a_24050_8154# 0.84fF
C11444 a_14314_4178# col_n[11] 0.11fF
C11445 a_2275_13198# a_35002_13174# 0.17fF
C11446 a_24354_16226# col_n[21] 0.11fF
C11447 a_32082_5142# vcm 0.89fF
C11448 a_8990_4138# rowoff_n[2] 2.33fF
C11449 a_26058_12170# rowoff_n[10] 1.50fF
C11450 a_22042_12170# rowon_n[10] 0.45fF
C11451 a_2475_12194# m2_34864_11990# 0.56fF
C11452 a_2475_5166# a_3878_5142# 0.41fF
C11453 a_2275_5166# a_2874_5142# 0.17fF
C11454 a_2475_7174# col[2] 0.22fF
C11455 a_6982_13174# VDD 4.02fF
C11456 a_2475_10186# a_27062_10162# 0.68fF
C11457 a_14010_10162# a_15014_10162# 0.86fF
C11458 a_18026_2130# rowoff_n[0] 1.89fF
C11459 a_32082_2130# rowon_n[0] 0.45fF
C11460 a_7986_2130# col[5] 0.38fF
C11461 a_13006_8154# vcm 0.89fF
C11462 rowon_n[12] rowoff_n[12] 20.66fF
C11463 a_2275_13198# col_n[9] 0.17fF
C11464 a_18026_14178# col[15] 0.38fF
C11465 a_32994_3134# a_33086_3134# 0.45fF
C11466 a_2275_2154# col_n[14] 0.17fF
C11467 a_1957_17214# vcm 0.16fF
C11468 a_15014_15182# m2_15212_15430# 0.19fF
C11469 a_2275_7174# a_18026_7150# 0.71fF
C11470 a_9994_2130# row_n[0] 0.43fF
C11471 m2_29844_946# col[27] 0.52fF
C11472 a_22042_17190# VDD 2.47fF
C11473 a_33086_10162# col_n[30] 0.34fF
C11474 a_4974_12170# a_4974_11166# 0.84fF
C11475 a_9902_6146# rowon_n[4] 0.14fF
C11476 a_3270_2170# vcm 0.25fF
C11477 a_13310_14218# col_n[10] 0.11fF
C11478 a_28066_12170# vcm 0.89fF
C11479 a_24962_2130# VDD 0.29fF
C11480 a_34090_11166# m2_34288_11414# 0.19fF
C11481 a_2475_4162# a_10906_4138# 0.41fF
C11482 a_2275_4162# a_8290_4178# 0.15fF
C11483 m3_1864_9110# m3_1864_8106# 0.20fF
C11484 a_2275_9182# a_33086_9158# 0.71fF
C11485 a_2475_9182# col[19] 0.22fF
C11486 a_23958_18194# m2_23820_18014# 0.34fF
C11487 a_29070_14178# a_30074_14178# 0.86fF
C11488 a_10906_10162# rowoff_n[8] 0.65fF
C11489 col_n[22] rowoff_n[13] 0.18fF
C11490 a_18330_6186# vcm 0.24fF
C11491 a_14010_13174# rowoff_n[11] 2.08fF
C11492 a_8990_15182# vcm 0.89fF
C11493 a_2275_15206# col_n[26] 0.17fF
C11494 col[16] rowoff_n[0] 0.24fF
C11495 col[17] rowoff_n[1] 0.23fF
C11496 col[18] rowoff_n[2] 0.23fF
C11497 col[19] rowoff_n[3] 0.22fF
C11498 col[20] rowoff_n[4] 0.21fF
C11499 col[21] rowoff_n[5] 0.21fF
C11500 col[22] rowoff_n[6] 0.20fF
C11501 col[23] rowoff_n[7] 0.19fF
C11502 col[24] rowoff_n[8] 0.19fF
C11503 col[25] rowoff_n[9] 0.18fF
C11504 a_5886_5142# VDD 0.29fF
C11505 a_6982_12170# col[4] 0.38fF
C11506 a_2275_4162# col_n[31] 0.17fF
C11507 a_5978_13174# m2_6176_13422# 0.19fF
C11508 a_2475_6170# a_25966_6146# 0.41fF
C11509 a_2275_6170# a_23350_6186# 0.15fF
C11510 a_13918_6146# a_14010_6146# 0.45fF
C11511 a_30074_9158# rowon_n[7] 0.45fF
C11512 a_19942_8154# rowoff_n[6] 0.55fF
C11513 a_22042_8154# col_n[19] 0.34fF
C11514 a_2275_15206# a_2966_15182# 0.67fF
C11515 a_2475_15206# a_3970_15182# 0.68fF
C11516 a_20034_16186# a_20034_15182# 0.84fF
C11517 a_2275_12194# col[16] 0.17fF
C11518 a_33390_10202# vcm 0.24fF
C11519 a_2275_1150# col[21] 0.17fF
C11520 a_30074_17190# rowoff_n[15] 1.30fF
C11521 a_28978_6146# rowoff_n[4] 0.44fF
C11522 a_25054_9158# m2_25252_9406# 0.19fF
C11523 a_2275_3158# a_16930_3134# 0.17fF
C11524 a_12002_4138# ctop 4.91fF
C11525 a_2475_1150# m2_13780_946# 0.62fF
C11526 a_20946_9158# VDD 0.29fF
C11527 m3_8892_1078# ctop 0.21fF
C11528 a_7986_9158# row_n[7] 0.43fF
C11529 a_7894_13174# rowon_n[11] 0.14fF
C11530 col_n[6] rowoff_n[14] 0.29fF
C11531 a_26970_4138# vcm 0.18fF
C11532 a_9994_17190# a_10998_17190# 0.86fF
C11533 a_17934_3134# rowon_n[1] 0.14fF
C11534 a_2475_17214# a_19030_17190# 0.68fF
C11535 col[9] rowoff_n[10] 0.29fF
C11536 m2_9764_18014# m2_10768_18014# 0.86fF
C11537 a_14314_13214# vcm 0.24fF
C11538 a_2275_5166# a_31990_5142# 0.17fF
C11539 a_27062_8154# ctop 4.91fF
C11540 a_2275_18218# col_n[28] 0.17fF
C11541 a_28978_10162# a_29070_10162# 0.45fF
C11542 a_2275_14202# a_9994_14178# 0.71fF
C11543 a_7894_7150# vcm 0.18fF
C11544 a_10998_6146# col_n[8] 0.34fF
C11545 a_2475_14202# rowoff_n[12] 4.75fF
C11546 a_16018_7150# m2_16216_7398# 0.19fF
C11547 a_2475_2154# a_24050_2130# 0.68fF
C11548 a_30074_3134# a_30074_2130# 0.84fF
C11549 a_29374_17230# vcm 0.24fF
C11550 a_28066_16186# rowon_n[14] 0.45fF
C11551 a_7986_11166# ctop 4.91fF
C11552 a_16930_16186# VDD 0.29fF
C11553 col_n[11] col[12] 6.22fF
C11554 VDD col[26] 7.00fF
C11555 vcm col[23] 6.66fF
C11556 a_2275_11190# col_n[3] 0.17fF
C11557 a_2275_16210# a_25054_16186# 0.71fF
C11558 a_22954_11166# vcm 0.18fF
C11559 a_5978_16186# row_n[14] 0.43fF
C11560 a_19030_1126# VDD 4.98fF
C11561 m2_34864_13998# row_n[12] 0.38fF
C11562 a_20034_4138# a_21038_4138# 0.86fF
C11563 a_31078_5142# col[28] 0.38fF
C11564 a_20034_17190# m2_19804_18014# 0.84fF
C11565 a_23046_15182# ctop 4.91fF
C11566 a_16018_6146# row_n[4] 0.43fF
C11567 a_15926_10162# rowon_n[8] 0.14fF
C11568 a_9902_13174# a_9994_13174# 0.45fF
C11569 a_2475_13198# a_17934_13174# 0.41fF
C11570 a_2275_13198# a_15318_13214# 0.15fF
C11571 m2_27260_2378# a_27062_2130# 0.19fF
C11572 m2_7756_946# vcm 0.71fF
C11573 a_6982_5142# m2_7180_5390# 0.19fF
C11574 a_2275_1150# a_30074_1126# 0.14fF
C11575 a_2475_7174# col[13] 0.22fF
C11576 a_34090_5142# VDD 1.23fF
C11577 a_26362_5182# col_n[23] 0.11fF
C11578 a_10998_6146# a_10998_5142# 0.84fF
C11579 a_9994_16186# col_n[7] 0.34fF
C11580 a_2275_10186# a_8898_10162# 0.17fF
C11581 m2_34864_1950# m2_34864_2954# 0.84fF
C11582 a_2275_13198# col_n[20] 0.17fF
C11583 a_2475_15206# a_32994_15182# 0.41fF
C11584 a_2275_15206# a_30378_15222# 0.15fF
C11585 a_2275_2154# col_n[25] 0.17fF
C11586 a_2874_4138# rowon_n[2] 0.14fF
C11587 a_18938_18194# vcm 0.18fF
C11588 a_15014_8154# VDD 3.20fF
C11589 a_2275_10186# col[10] 0.17fF
C11590 a_20034_3134# col[17] 0.38fF
C11591 a_34394_17230# col_n[31] 0.11fF
C11592 a_2275_12194# a_23958_12170# 0.17fF
C11593 a_30074_15182# col[27] 0.38fF
C11594 a_21038_3134# vcm 0.89fF
C11595 a_24962_17190# a_25054_17190# 0.45fF
C11596 a_2475_9182# col[30] 0.22fF
C11597 a_14010_13174# row_n[11] 0.43fF
C11598 a_30074_12170# VDD 1.65fF
C11599 m3_16924_18146# m3_17928_18146# 0.21fF
C11600 a_15318_3174# col_n[12] 0.11fF
C11601 a_13918_17190# rowon_n[15] 0.14fF
C11602 a_26058_10162# a_26058_9158# 0.84fF
C11603 a_2475_9182# a_16018_9158# 0.68fF
C11604 a_25358_15222# col_n[22] 0.11fF
C11605 a_24050_3134# row_n[1] 0.43fF
C11606 a_9994_3134# rowoff_n[1] 2.28fF
C11607 sample_n rowoff_n[5] 0.55fF
C11608 col[31] rowoff_n[4] 0.14fF
C11609 col[30] rowoff_n[3] 0.15fF
C11610 col[29] rowoff_n[2] 0.15fF
C11611 col[28] rowoff_n[1] 0.16fF
C11612 col[27] rowoff_n[0] 0.17fF
C11613 a_2275_15206# row_n[13] 26.41fF
C11614 a_2475_6170# vcm 1.32fF
C11615 a_23958_7150# rowon_n[5] 0.14fF
C11616 a_30986_14178# rowoff_n[12] 0.42fF
C11617 a_2275_6170# a_6982_6146# 0.71fF
C11618 a_10998_15182# VDD 3.61fF
C11619 a_2475_11190# a_31078_11166# 0.68fF
C11620 a_16018_11166# a_17022_11166# 0.86fF
C11621 a_2275_12194# col[27] 0.17fF
C11622 a_26362_1166# vcm 0.25fF
C11623 a_19030_13174# col[16] 0.38fF
C11624 a_17022_10162# vcm 0.89fF
C11625 a_35002_4138# a_35094_4138# 0.11fF
C11626 m3_4876_18146# ctop 0.21fF
C11627 a_2275_9182# VDD 3.18fF
C11628 col_n[17] rowoff_n[14] 0.21fF
C11629 a_34090_9158# col_n[31] 0.34fF
C11630 a_2275_8178# a_22042_8154# 0.71fF
C11631 a_6982_13174# a_6982_12170# 0.84fF
C11632 col[20] rowoff_n[10] 0.21fF
C11633 a_14314_13214# col_n[11] 0.11fF
C11634 a_7286_4178# vcm 0.24fF
C11635 a_2161_11190# rowoff_n[9] 0.14fF
C11636 a_32082_14178# vcm 0.89fF
C11637 a_28978_4138# VDD 0.29fF
C11638 a_2475_5166# a_14922_5142# 0.41fF
C11639 a_2275_5166# a_12306_5182# 0.15fF
C11640 a_2275_18218# a_10906_18194# 0.17fF
C11641 a_22042_10162# row_n[8] 0.43fF
C11642 a_11910_9158# rowoff_n[7] 0.64fF
C11643 a_2475_16210# col[2] 0.22fF
C11644 a_21950_14178# rowon_n[12] 0.14fF
C11645 a_2475_5166# col[7] 0.22fF
C11646 a_31078_15182# a_32082_15182# 0.86fF
C11647 a_22346_8194# vcm 0.24fF
C11648 a_18938_15182# rowoff_n[13] 0.56fF
C11649 a_2475_7174# m2_1732_6970# 0.16fF
C11650 a_31990_4138# rowon_n[2] 0.14fF
C11651 a_2275_2154# a_5886_2130# 0.17fF
C11652 a_7986_11166# col[5] 0.38fF
C11653 a_13006_17190# vcm 0.89fF
C11654 col_n[17] col[17] 0.43fF
C11655 rowon_n[11] ctop 0.37fF
C11656 col_n[1] rowoff_n[15] 0.33fF
C11657 m2_19804_18014# m3_19936_18146# 4.41fF
C11658 a_9902_7150# VDD 0.29fF
C11659 a_20946_7150# rowoff_n[5] 0.54fF
C11660 a_2275_7174# a_27366_7190# 0.15fF
C11661 a_2475_7174# a_29982_7150# 0.41fF
C11662 a_15926_7150# a_16018_7150# 0.45fF
C11663 a_2275_11190# col_n[14] 0.17fF
C11664 col[4] rowoff_n[11] 0.32fF
C11665 a_23046_7150# col_n[20] 0.34fF
C11666 a_15926_2130# vcm 0.18fF
C11667 a_2475_16210# a_7986_16186# 0.68fF
C11668 a_22042_17190# a_22042_16186# 0.84fF
C11669 a_3270_11206# vcm 0.24fF
C11670 a_29982_5142# rowoff_n[3] 0.43fF
C11671 a_35494_2492# VDD 0.13fF
C11672 a_2275_8178# col[4] 0.17fF
C11673 a_8990_8154# rowon_n[6] 0.45fF
C11674 a_2275_4162# a_20946_4138# 0.17fF
C11675 a_16018_6146# ctop 4.91fF
C11676 a_24962_11166# VDD 0.29fF
C11677 m3_6884_1078# m3_7888_1078# 0.21fF
C11678 m2_10768_18014# col[8] 0.39fF
C11679 a_2475_7174# col[24] 0.22fF
C11680 a_30986_6146# vcm 0.18fF
C11681 a_18330_15222# vcm 0.24fF
C11682 a_2475_18218# a_23958_18194# 0.41fF
C11683 a_2275_6170# a_34394_6186# 0.15fF
C11684 m2_11772_946# VDD 5.95fF
C11685 a_31078_10162# ctop 4.91fF
C11686 a_20034_17190# row_n[15] 0.43fF
C11687 a_5886_14178# VDD 0.29fF
C11688 a_2275_13198# col_n[31] 0.17fF
C11689 a_30986_11166# a_31078_11166# 0.45fF
C11690 a_30074_7150# row_n[5] 0.43fF
C11691 a_2275_15206# a_14010_15182# 0.71fF
C11692 a_12002_5142# col_n[9] 0.34fF
C11693 a_29982_11166# rowon_n[9] 0.14fF
C11694 a_11910_9158# vcm 0.18fF
C11695 a_22042_17190# col_n[19] 0.34fF
C11696 a_6890_16186# rowoff_n[14] 0.69fF
C11697 a_2475_3158# a_28066_3134# 0.68fF
C11698 a_32082_4138# a_32082_3134# 0.84fF
C11699 a_2275_10186# col[21] 0.17fF
C11700 a_21038_16186# m2_21236_16434# 0.19fF
C11701 a_12002_13174# ctop 4.91fF
C11702 a_1957_18218# m2_1732_18014# 0.33fF
C11703 a_20946_18194# VDD 0.50fF
C11704 a_2275_12194# a_4274_12210# 0.15fF
C11705 a_2475_12194# a_6890_12170# 0.41fF
C11706 a_2966_3134# vcm 0.89fF
C11707 a_31078_11166# rowoff_n[9] 1.25fF
C11708 a_2275_17214# a_29070_17190# 0.71fF
C11709 m2_26832_18014# col_n[24] 0.32fF
C11710 a_6982_15182# rowon_n[13] 0.45fF
C11711 m2_20808_18014# m2_21236_18442# 0.19fF
C11712 a_26970_13174# vcm 0.18fF
C11713 a_32082_4138# col[29] 0.38fF
C11714 a_23046_3134# VDD 2.37fF
C11715 a_22042_5142# a_23046_5142# 0.86fF
C11716 a_17022_5142# rowon_n[3] 0.45fF
C11717 a_27062_17190# ctop 4.93fF
C11718 a_11910_14178# a_12002_14178# 0.45fF
C11719 a_2275_14202# a_19334_14218# 0.15fF
C11720 a_2475_14202# a_21950_14178# 0.41fF
C11721 m2_34864_6970# VDD 1.58fF
C11722 a_27366_4178# col_n[24] 0.11fF
C11723 a_2275_2154# a_34090_2130# 0.71fF
C11724 a_7894_16186# vcm 0.18fF
C11725 a_10998_15182# col_n[8] 0.34fF
C11726 a_3970_6146# VDD 4.33fF
C11727 a_13006_7150# a_13006_6146# 0.84fF
C11728 a_12002_14178# m2_12200_14426# 0.19fF
C11729 a_2475_3158# col[1] 0.22fF
C11730 a_28066_14178# row_n[12] 0.43fF
C11731 a_2275_11190# a_12914_11166# 0.17fF
C11732 a_9994_1126# vcm 0.15fF
C11733 a_2275_16210# a_35398_16226# 0.15fF
C11734 a_8990_2130# m2_9188_2378# 0.19fF
C11735 a_2275_9182# col_n[8] 0.17fF
C11736 col_n[28] rowoff_n[14] 0.14fF
C11737 a_31078_10162# m2_31276_10410# 0.19fF
C11738 a_4974_2130# m2_4744_946# 0.84fF
C11739 a_19030_10162# VDD 2.78fF
C11740 a_21038_2130# col[18] 0.38fF
C11741 col[31] rowoff_n[10] 0.14fF
C11742 a_2475_8178# a_4974_8154# 0.68fF
C11743 a_31078_14178# col[28] 0.38fF
C11744 a_2275_13198# a_27974_13174# 0.17fF
C11745 a_25054_5142# vcm 0.89fF
C11746 a_2475_4162# rowoff_n[2] 4.75fF
C11747 a_26970_18194# a_27062_18194# 0.11fF
C11748 a_19030_12170# rowoff_n[10] 1.84fF
C11749 m2_30848_946# vcm 0.71fF
C11750 a_2275_18218# m2_27836_18014# 0.51fF
C11751 a_21950_1126# a_22042_1126# 0.11fF
C11752 a_15014_12170# rowon_n[10] 0.45fF
C11753 a_16322_2170# col_n[13] 0.11fF
C11754 a_2475_16210# col[13] 0.22fF
C11755 a_26362_14218# col_n[23] 0.11fF
C11756 a_34090_14178# VDD 1.23fF
C11757 a_2475_5166# col[18] 0.22fF
C11758 a_28066_11166# a_28066_10162# 0.84fF
C11759 a_2475_10186# a_20034_10162# 0.68fF
C11760 a_10998_2130# rowoff_n[0] 2.23fF
C11761 a_25054_2130# rowon_n[0] 0.45fF
C11762 a_3878_14178# rowon_n[12] 0.14fF
C11763 row_n[6] ctop 0.28fF
C11764 rowon_n[2] row_n[2] 21.02fF
C11765 col_n[22] col[23] 6.22fF
C11766 col_n[12] rowoff_n[15] 0.25fF
C11767 a_5978_8154# vcm 0.89fF
C11768 a_2275_11190# col_n[25] 0.17fF
C11769 a_22042_8154# m2_22240_8402# 0.19fF
C11770 a_32994_1126# m2_32856_946# 0.30fF
C11771 col[15] rowoff_n[11] 0.25fF
C11772 a_2275_7174# rowoff_n[5] 0.81fF
C11773 a_2275_7174# a_10998_7150# 0.71fF
C11774 a_15014_17190# VDD 3.20fF
C11775 a_18026_12170# a_19030_12170# 0.86fF
C11776 a_20034_12170# col[17] 0.38fF
C11777 a_30378_3174# vcm 0.24fF
C11778 a_2275_8178# col[15] 0.17fF
C11779 a_21038_12170# vcm 0.89fF
C11780 a_17934_2130# VDD 0.29fF
C11781 m2_26832_946# m3_26964_1078# 4.41fF
C11782 m3_1864_16138# m3_1864_15134# 0.20fF
C11783 a_2275_9182# a_26058_9158# 0.71fF
C11784 a_15318_12210# col_n[12] 0.11fF
C11785 a_8990_14178# a_8990_13174# 0.84fF
C11786 a_11302_6186# vcm 0.24fF
C11787 a_6982_13174# rowoff_n[11] 2.42fF
C11788 a_13006_6146# m2_13204_6394# 0.19fF
C11789 a_2475_15206# vcm 1.32fF
C11790 a_32994_6146# VDD 0.29fF
C11791 a_2275_6170# a_16322_6186# 0.15fF
C11792 a_2475_6170# a_18938_6146# 0.41fF
C11793 m2_13780_946# col[11] 0.51fF
C11794 a_1957_17214# row_n[15] 0.29fF
C11795 a_23046_9158# rowon_n[7] 0.45fF
C11796 a_12914_8154# rowoff_n[6] 0.63fF
C11797 m2_34864_16006# rowon_n[14] 0.42fF
C11798 a_33086_16186# a_34090_16186# 0.86fF
C11799 a_26362_10202# vcm 0.24fF
C11800 a_8990_10162# col[6] 0.38fF
C11801 a_23046_17190# rowoff_n[15] 1.64fF
C11802 a_21950_6146# rowoff_n[4] 0.52fF
C11803 a_2275_3158# a_9902_3134# 0.17fF
C11804 a_4974_4138# ctop 4.91fF
C11805 m3_1864_11118# ctop 0.22fF
C11806 a_13918_9158# VDD 0.29fF
C11807 a_2275_8178# a_31382_8194# 0.15fF
C11808 a_2475_8178# a_33998_8154# 0.41fF
C11809 a_17934_8154# a_18026_8154# 0.45fF
C11810 a_24050_6146# col_n[21] 0.34fF
C11811 a_2275_7174# col_n[2] 0.17fF
C11812 a_19942_4138# vcm 0.18fF
C11813 a_30986_4138# rowoff_n[2] 0.42fF
C11814 a_4274_10202# col_n[1] 0.11fF
C11815 a_10906_3134# rowon_n[1] 0.14fF
C11816 a_2475_17214# a_12002_17190# 0.68fF
C11817 m2_2736_18014# m2_3740_18014# 0.86fF
C11818 a_3970_4138# m2_4168_4386# 0.19fF
C11819 a_7286_13214# vcm 0.24fF
C11820 a_2275_5166# a_24962_5142# 0.17fF
C11821 a_20034_8154# ctop 4.91fF
C11822 a_28978_13174# VDD 0.29fF
C11823 m2_1732_12994# sample_n 0.12fF
C11824 a_2475_14202# a_3878_14178# 0.41fF
C11825 a_2275_14202# a_2874_14178# 0.17fF
C11826 a_35002_8154# vcm 0.18fF
C11827 a_2475_14202# col[7] 0.22fF
C11828 a_2475_3158# col[12] 0.22fF
C11829 a_2475_2154# a_17022_2130# 0.68fF
C11830 a_8990_2130# a_9994_2130# 0.86fF
C11831 a_22346_17230# vcm 0.24fF
C11832 a_21038_16186# rowon_n[14] 0.45fF
C11833 a_9902_16186# VDD 0.29fF
C11834 a_32994_12170# a_33086_12170# 0.45fF
C11835 a_31078_6146# rowon_n[4] 0.45fF
C11836 a_13006_4138# col_n[10] 0.34fF
C11837 a_2275_9182# col_n[19] 0.17fF
C11838 a_23046_16186# col_n[20] 0.34fF
C11839 a_2275_16210# a_18026_16186# 0.71fF
C11840 a_15926_11166# vcm 0.18fF
C11841 a_12002_1126# VDD 0.13fF
C11842 a_34090_5142# a_34090_4138# 0.84fF
C11843 a_2475_4162# a_32082_4138# 0.68fF
C11844 a_35494_11528# VDD 0.13fF
C11845 a_2275_17214# col[4] 0.17fF
C11846 a_16018_15182# ctop 4.91fF
C11847 a_2275_6170# col[9] 0.17fF
C11848 a_8990_6146# row_n[4] 0.43fF
C11849 a_8898_10162# rowon_n[8] 0.14fF
C11850 a_2475_13198# a_10906_13174# 0.41fF
C11851 a_2275_13198# a_8290_13214# 0.15fF
C11852 a_32082_10162# rowoff_n[8] 1.20fF
C11853 a_33086_3134# col[30] 0.38fF
C11854 a_2275_1150# a_23046_1126# 0.14fF
C11855 a_2475_16210# col[24] 0.22fF
C11856 a_30986_15182# vcm 0.18fF
C11857 a_2475_5166# col[29] 0.22fF
C11858 a_27062_5142# VDD 1.96fF
C11859 a_24050_6146# a_25054_6146# 0.86fF
C11860 col_n[28] col[28] 0.54fF
C11861 rowon_n[0] ctop 0.36fF
C11862 col_n[23] rowoff_n[15] 0.17fF
C11863 a_2475_15206# a_25966_15182# 0.41fF
C11864 a_2275_15206# a_23350_15222# 0.15fF
C11865 a_13918_15182# a_14010_15182# 0.45fF
C11866 a_28370_3174# col_n[25] 0.11fF
C11867 m2_1732_10986# m2_1732_9982# 0.84fF
C11868 col[26] rowoff_n[11] 0.17fF
C11869 a_12002_14178# col_n[9] 0.34fF
C11870 a_11910_18194# vcm 0.18fF
C11871 a_7986_8154# VDD 3.92fF
C11872 a_15014_8154# a_15014_7150# 0.84fF
C11873 a_29070_13174# rowon_n[11] 0.45fF
C11874 a_2275_12194# a_16930_12170# 0.17fF
C11875 a_2275_8178# col[26] 0.17fF
C11876 a_14010_3134# vcm 0.89fF
C11877 a_2966_12170# vcm 0.89fF
C11878 a_6982_13174# row_n[11] 0.43fF
C11879 a_23046_12170# VDD 2.37fF
C11880 a_32082_13174# col[29] 0.38fF
C11881 m3_2868_18146# m3_3872_18146# 0.21fF
C11882 a_6890_17190# rowon_n[15] 0.14fF
C11883 a_2475_9182# a_8990_9158# 0.68fF
C11884 a_4974_9158# a_5978_9158# 0.86fF
C11885 m2_34864_7974# vcm 0.72fF
C11886 a_2275_14202# a_31990_14178# 0.17fF
C11887 a_2874_3134# rowoff_n[1] 0.74fF
C11888 a_17022_3134# row_n[1] 0.43fF
C11889 col[10] rowoff_n[12] 0.28fF
C11890 a_29070_7150# vcm 0.89fF
C11891 a_16930_7150# rowon_n[5] 0.14fF
C11892 a_23958_14178# rowoff_n[12] 0.50fF
C11893 a_23958_2130# a_24050_2130# 0.45fF
C11894 a_17326_1166# col_n[14] 0.11fF
C11895 a_27366_13214# col_n[24] 0.11fF
C11896 a_3970_15182# VDD 4.33fF
C11897 a_30074_12170# a_30074_11166# 0.84fF
C11898 a_2475_11190# a_24050_11166# 0.68fF
C11899 a_2475_12194# col[1] 0.22fF
C11900 a_2475_1150# col[6] 0.22fF
C11901 a_19334_1166# vcm 0.24fF
C11902 a_9994_10162# vcm 0.89fF
C11903 a_3878_6146# rowoff_n[4] 0.73fF
C11904 a_2275_7174# col_n[13] 0.17fF
C11905 a_2275_8178# a_15014_8154# 0.71fF
C11906 a_27062_17190# m2_27260_17438# 0.19fF
C11907 a_21038_11166# col[18] 0.38fF
C11908 a_20034_13174# a_21038_13174# 0.86fF
C11909 ctop rowoff_n[13] 0.28fF
C11910 a_35398_5182# vcm 0.24fF
C11911 a_3270_7190# col_n[0] 0.11fF
C11912 a_25054_14178# vcm 0.89fF
C11913 a_2275_4162# col[3] 0.17fF
C11914 a_21950_4138# VDD 0.29fF
C11915 a_2275_5166# a_5278_5182# 0.15fF
C11916 a_2475_5166# a_7894_5142# 0.41fF
C11917 a_4882_5142# a_4974_5142# 0.45fF
C11918 a_2275_10186# a_30074_10162# 0.71fF
C11919 a_16322_11206# col_n[13] 0.11fF
C11920 a_15014_10162# row_n[8] 0.43fF
C11921 a_4882_9158# rowoff_n[7] 0.72fF
C11922 a_2475_14202# col[18] 0.22fF
C11923 a_14922_14178# rowon_n[12] 0.14fF
C11924 a_10998_15182# a_10998_14178# 0.84fF
C11925 a_2475_3158# col[23] 0.22fF
C11926 a_15318_8194# vcm 0.24fF
C11927 a_11910_15182# rowoff_n[13] 0.64fF
C11928 m2_1732_9982# VDD 5.46fF
C11929 a_2475_18218# col[9] 0.22fF
C11930 a_24962_4138# rowon_n[2] 0.14fF
C11931 a_28066_3134# ctop 4.91fF
C11932 a_5978_17190# vcm 0.89fF
C11933 a_2966_16186# rowon_n[14] 0.45fF
C11934 a_2161_7174# VDD 0.23fF
C11935 a_13918_7150# rowoff_n[5] 0.61fF
C11936 a_2275_7174# a_20338_7190# 0.15fF
C11937 a_2475_7174# a_22954_7150# 0.41fF
C11938 a_18026_15182# m2_18224_15430# 0.19fF
C11939 a_2275_9182# col_n[30] 0.17fF
C11940 a_8898_2130# vcm 0.18fF
C11941 a_9994_9158# col[7] 0.38fF
C11942 a_22954_5142# rowoff_n[3] 0.51fF
C11943 a_30378_12210# vcm 0.24fF
C11944 a_2275_17214# col[15] 0.17fF
C11945 a_2475_8178# rowon_n[6] 0.40fF
C11946 a_2275_4162# a_13918_4138# 0.17fF
C11947 a_8990_6146# ctop 4.91fF
C11948 a_2275_6170# col[20] 0.17fF
C11949 a_25054_5142# col_n[22] 0.34fF
C11950 a_17934_11166# VDD 0.29fF
C11951 a_2275_18218# col[0] 0.16fF
C11952 a_19942_9158# a_20034_9158# 0.45fF
C11953 a_31990_3134# rowoff_n[1] 0.41fF
C11954 a_5278_9198# col_n[2] 0.11fF
C11955 a_23958_6146# vcm 0.18fF
C11956 a_11302_15222# vcm 0.24fF
C11957 a_2475_18218# a_16930_18194# 0.41fF
C11958 a_2275_6170# a_28978_6146# 0.17fF
C11959 a_8990_13174# m2_9188_13422# 0.19fF
C11960 a_24050_10162# ctop 4.91fF
C11961 a_13006_17190# row_n[15] 0.43fF
C11962 row_n[14] sample_n 0.16fF
C11963 ctop col[1] 0.13fF
C11964 a_32994_15182# VDD 0.29fF
C11965 m2_29844_18014# vcm 0.71fF
C11966 a_23046_7150# row_n[5] 0.43fF
C11967 a_2275_15206# a_6982_15182# 0.71fF
C11968 a_22954_11166# rowon_n[9] 0.14fF
C11969 a_4882_9158# vcm 0.18fF
C11970 a_2475_3158# a_21038_3134# 0.68fF
C11971 a_28066_9158# m2_28264_9406# 0.19fF
C11972 a_10998_3134# a_12002_3134# 0.86fF
C11973 a_2475_1150# m2_22816_946# 0.62fF
C11974 m3_23952_1078# ctop 0.21fF
C11975 a_4974_13174# ctop 4.91fF
C11976 a_13918_18194# VDD 0.50fF
C11977 a_14010_3134# col_n[11] 0.34fF
C11978 a_35002_13174# a_35094_13174# 0.11fF
C11979 a_24050_15182# col_n[21] 0.34fF
C11980 a_24050_11166# rowoff_n[9] 1.59fF
C11981 a_2275_17214# a_22042_17190# 0.71fF
C11982 a_2275_16210# col_n[2] 0.17fF
C11983 m2_13780_18014# m2_14208_18442# 0.19fF
C11984 a_2275_5166# col_n[7] 0.17fF
C11985 a_19942_13174# vcm 0.18fF
C11986 a_16018_3134# VDD 3.09fF
C11987 m2_23820_946# col[21] 0.51fF
C11988 a_1957_9182# sample 0.35fF
C11989 a_9994_5142# rowon_n[3] 0.45fF
C11990 a_2275_18218# a_32082_18194# 0.14fF
C11991 a_20034_17190# ctop 4.93fF
C11992 col[21] rowoff_n[12] 0.21fF
C11993 a_33086_9158# rowoff_n[7] 1.15fF
C11994 a_2275_14202# a_12306_14218# 0.15fF
C11995 a_2475_14202# a_14922_14178# 0.41fF
C11996 a_34090_2130# col[31] 0.38fF
C11997 m2_34864_4962# row_n[3] 0.38fF
C11998 a_2275_2154# a_27062_2130# 0.71fF
C11999 a_19030_7150# m2_19228_7398# 0.19fF
C12000 a_35002_17190# vcm 0.18fF
C12001 m2_1732_16006# m3_1864_16138# 4.42fF
C12002 a_31078_7150# VDD 1.54fF
C12003 a_2475_12194# col[12] 0.22fF
C12004 a_26058_7150# a_27062_7150# 0.86fF
C12005 a_2475_1150# col[17] 0.21fF
C12006 a_2275_11190# a_5886_11166# 0.17fF
C12007 a_21038_14178# row_n[12] 0.43fF
C12008 a_2874_1126# vcm 0.18fF
C12009 a_29374_2170# col_n[26] 0.11fF
C12010 a_2275_16210# a_27366_16226# 0.15fF
C12011 a_2475_16210# a_29982_16186# 0.41fF
C12012 a_15926_16186# a_16018_16186# 0.45fF
C12013 a_13006_13174# col_n[10] 0.34fF
C12014 a_31078_4138# row_n[2] 0.43fF
C12015 a_2275_7174# col_n[24] 0.17fF
C12016 a_30986_8154# rowon_n[6] 0.14fF
C12017 a_12002_10162# VDD 3.51fF
C12018 col[5] rowoff_n[13] 0.31fF
C12019 a_17022_9158# a_17022_8154# 0.84fF
C12020 a_2275_13198# a_20946_13174# 0.17fF
C12021 a_2275_15206# col[9] 0.17fF
C12022 a_18026_5142# vcm 0.89fF
C12023 a_12002_12170# rowoff_n[10] 2.18fF
C12024 a_2275_4162# col[14] 0.17fF
C12025 m2_30272_2378# a_30074_2130# 0.19fF
C12026 a_2275_18218# m2_13780_18014# 0.51fF
C12027 a_2275_1150# a_32386_1166# 0.15fF
C12028 a_9994_5142# m2_10192_5390# 0.19fF
C12029 a_7986_12170# rowon_n[10] 0.45fF
C12030 a_3878_4138# VDD 0.29fF
C12031 a_33086_12170# col[30] 0.38fF
C12032 a_27062_14178# VDD 1.96fF
C12033 a_2475_14202# col[29] 0.22fF
C12034 a_6982_10162# a_7986_10162# 0.86fF
C12035 a_2475_10186# a_13006_10162# 0.68fF
C12036 a_18026_2130# rowon_n[0] 0.45fF
C12037 a_3970_2130# rowoff_n[0] 2.57fF
C12038 a_2275_15206# a_34394_15222# 0.15fF
C12039 a_2475_18218# col[20] 0.22fF
C12040 a_33086_9158# vcm 0.89fF
C12041 a_28066_16186# rowoff_n[14] 1.40fF
C12042 a_28370_12210# col_n[25] 0.11fF
C12043 a_25966_3134# a_26058_3134# 0.45fF
C12044 a_2275_7174# a_3970_7150# 0.71fF
C12045 a_7986_17190# VDD 3.92fF
C12046 a_32082_13174# a_32082_12170# 0.84fF
C12047 a_2475_12194# a_28066_12170# 0.68fF
C12048 a_23350_3174# vcm 0.24fF
C12049 a_29070_11166# row_n[9] 0.43fF
C12050 a_2275_17214# col[26] 0.17fF
C12051 a_28978_15182# rowon_n[13] 0.14fF
C12052 a_2275_6170# col[31] 0.17fF
C12053 a_14010_12170# vcm 0.89fF
C12054 a_2275_18218# col[11] 0.17fF
C12055 a_10906_2130# VDD 0.29fF
C12056 a_2275_9182# a_19030_9158# 0.71fF
C12057 a_22042_10162# col[19] 0.38fF
C12058 a_2275_3158# col_n[1] 0.17fF
C12059 a_22042_14178# a_23046_14178# 0.86fF
C12060 a_4274_6186# vcm 0.24fF
C12061 ctop col[12] 0.13fF
C12062 a_29070_16186# vcm 0.89fF
C12063 rowon_n[8] sample_n 0.15fF
C12064 m2_1732_12994# m3_1864_13126# 4.42fF
C12065 a_25966_6146# VDD 0.29fF
C12066 a_2275_6170# a_9294_6186# 0.15fF
C12067 a_2475_6170# a_11910_6146# 0.41fF
C12068 a_6890_6146# a_6982_6146# 0.45fF
C12069 a_17326_10202# col_n[14] 0.11fF
C12070 a_16018_9158# rowon_n[7] 0.45fF
C12071 a_5886_8154# rowoff_n[6] 0.70fF
C12072 a_2275_11190# a_34090_11166# 0.71fF
C12073 a_31990_1126# vcm 0.18fF
C12074 a_13006_16186# a_13006_15182# 0.84fF
C12075 a_2475_10186# col[6] 0.22fF
C12076 a_19334_10202# vcm 0.24fF
C12077 a_16018_17190# rowoff_n[15] 1.98fF
C12078 m2_33860_18014# VDD 2.09fF
C12079 a_2161_3158# a_2275_3158# 0.17fF
C12080 a_14922_6146# rowoff_n[4] 0.60fF
C12081 a_2475_3158# a_2966_3134# 0.65fF
C12082 a_32082_5142# ctop 4.91fF
C12083 m3_19936_18146# ctop 0.21fF
C12084 a_6890_9158# VDD 0.29fF
C12085 a_2275_8178# a_24354_8194# 0.15fF
C12086 a_2475_8178# a_26970_8154# 0.41fF
C12087 a_2275_16210# col_n[13] 0.17fF
C12088 a_10998_8154# col[8] 0.38fF
C12089 a_2275_5166# col_n[18] 0.17fF
C12090 a_12914_4138# vcm 0.18fF
C12091 a_23958_4138# rowoff_n[2] 0.50fF
C12092 a_2475_17214# a_4974_17190# 0.68fF
C12093 a_35398_14218# vcm 0.24fF
C12094 a_26058_4138# col_n[23] 0.34fF
C12095 a_2275_5166# a_17934_5142# 0.17fF
C12096 a_3270_16226# col_n[0] 0.11fF
C12097 sample_n rowoff_n[12] 0.55fF
C12098 a_13006_8154# ctop 4.91fF
C12099 a_21950_13174# VDD 0.29fF
C12100 a_2275_13198# col[3] 0.17fF
C12101 a_21950_10162# a_22042_10162# 0.45fF
C12102 a_2275_2154# col[8] 0.17fF
C12103 a_32994_2130# rowoff_n[0] 0.40fF
C12104 a_6282_8194# col_n[3] 0.11fF
C12105 m2_1732_10986# vcm 1.11fF
C12106 a_27974_8154# vcm 0.18fF
C12107 a_2475_12194# col[23] 0.22fF
C12108 a_23046_3134# a_23046_2130# 0.84fF
C12109 a_2475_2154# a_9994_2130# 0.68fF
C12110 a_15318_17230# vcm 0.24fF
C12111 m2_24824_18014# m3_24956_18146# 4.41fF
C12112 a_2475_1150# col[28] 0.22fF
C12113 a_14010_16186# rowon_n[14] 0.45fF
C12114 a_2275_7174# a_32994_7150# 0.17fF
C12115 a_28066_12170# ctop 4.91fF
C12116 a_2161_16210# VDD 0.23fF
C12117 a_2966_14178# row_n[12] 0.41fF
C12118 a_24050_6146# rowon_n[4] 0.45fF
C12119 a_2275_16210# a_10998_16186# 0.71fF
C12120 m2_34864_16006# m2_35292_16434# 0.19fF
C12121 a_8898_11166# vcm 0.18fF
C12122 a_4974_1126# VDD 0.15fF
C12123 col[16] rowoff_n[13] 0.24fF
C12124 a_2475_4162# a_25054_4138# 0.68fF
C12125 a_13006_4138# a_14010_4138# 0.86fF
C12126 a_15014_2130# col_n[12] 0.34fF
C12127 VDD rowoff_n[7] 87.22fF
C12128 col_n[0] rowoff_n[9] 0.34fF
C12129 sample rowoff_n[8] 0.22fF
C12130 a_8990_15182# ctop 4.91fF
C12131 a_2275_15206# col[20] 0.17fF
C12132 a_2475_6170# row_n[4] 0.48fF
C12133 a_25054_14178# col_n[22] 0.34fF
C12134 a_2275_4162# col[25] 0.17fF
C12135 a_25054_10162# rowoff_n[8] 1.54fF
C12136 a_28978_13174# rowoff_n[11] 0.44fF
C12137 a_5278_18234# col_n[2] 0.11fF
C12138 a_2966_8154# col_n[0] 0.34fF
C12139 a_2275_1150# a_16018_1126# 0.14fF
C12140 a_23958_15182# vcm 0.18fF
C12141 m2_1732_9982# m3_1864_10114# 4.42fF
C12142 a_20034_5142# VDD 2.68fF
C12143 m2_20808_946# VDD 4.63fF
C12144 a_3970_6146# a_3970_5142# 0.84fF
C12145 a_34090_8154# rowoff_n[6] 1.10fF
C12146 a_2475_18218# col[31] 0.22fF
C12147 a_2475_15206# a_18938_15182# 0.41fF
C12148 a_2275_15206# a_16322_15222# 0.15fF
C12149 col[0] rowoff_n[14] 0.34fF
C12150 a_2275_3158# a_31078_3134# 0.71fF
C12151 a_4882_18194# vcm 0.18fF
C12152 a_15926_1126# m2_15788_946# 0.31fF
C12153 a_28066_8154# a_29070_8154# 0.86fF
C12154 a_24050_16186# m2_24248_16434# 0.19fF
C12155 a_22042_13174# rowon_n[11] 0.45fF
C12156 a_30378_1166# col_n[27] 0.11fF
C12157 a_2475_8178# col[0] 0.20fF
C12158 a_2275_12194# a_9902_12170# 0.17fF
C12159 a_14010_12170# col_n[11] 0.34fF
C12160 a_6982_3134# vcm 0.89fF
C12161 a_2275_18218# col[22] 0.17fF
C12162 a_32082_3134# rowon_n[1] 0.45fF
C12163 a_2275_17214# a_31382_17230# 0.15fF
C12164 a_2475_17214# a_33998_17190# 0.41fF
C12165 a_17934_17190# a_18026_17190# 0.45fF
C12166 a_2475_11190# m2_34864_10986# 0.56fF
C12167 a_2275_14202# col_n[7] 0.17fF
C12168 a_16018_12170# VDD 3.09fF
C12169 a_2275_3158# col_n[12] 0.17fF
C12170 a_19030_10162# a_19030_9158# 0.84fF
C12171 a_2275_14202# a_24962_14178# 0.17fF
C12172 a_9994_3134# row_n[1] 0.43fF
C12173 VDD vcm 39.10fF
C12174 ctop col[23] 0.13fF
C12175 row_n[3] sample_n 0.16fF
C12176 m2_2736_18014# col_n[0] 0.32fF
C12177 a_9902_7150# rowon_n[5] 0.14fF
C12178 a_22042_7150# vcm 0.89fF
C12179 a_16930_14178# rowoff_n[12] 0.58fF
C12180 a_34090_11166# col[31] 0.38fF
C12181 m2_4744_18014# col[2] 0.37fF
C12182 a_15014_14178# m2_15212_14426# 0.19fF
C12183 a_31078_16186# VDD 1.54fF
C12184 a_8990_11166# a_9994_11166# 0.86fF
C12185 a_2475_11190# a_17022_11166# 0.68fF
C12186 a_2475_10186# col[17] 0.22fF
C12187 a_12306_1166# vcm 0.25fF
C12188 a_12002_2130# m2_12200_2378# 0.19fF
C12189 a_29374_11206# col_n[26] 0.11fF
C12190 a_2874_10162# vcm 0.18fF
C12191 a_35002_1126# VDD 0.74fF
C12192 a_27974_4138# a_28066_4138# 0.45fF
C12193 a_34090_10162# m2_34288_10410# 0.19fF
C12194 a_2275_16210# col_n[24] 0.17fF
C12195 a_2275_8178# a_7986_8154# 0.71fF
C12196 a_2275_5166# col_n[29] 0.17fF
C12197 a_30074_10162# rowon_n[8] 0.45fF
C12198 a_2475_13198# a_32082_13174# 0.68fF
C12199 a_34090_14178# a_34090_13174# 0.84fF
C12200 a_27366_5182# vcm 0.24fF
C12201 a_18026_14178# vcm 0.89fF
C12202 m2_1732_6970# m3_1864_7102# 4.42fF
C12203 a_2275_13198# col[14] 0.17fF
C12204 a_14922_4138# VDD 0.29fF
C12205 a_5978_12170# m2_6176_12418# 0.19fF
C12206 a_2275_2154# col[19] 0.17fF
C12207 a_23046_9158# col[20] 0.38fF
C12208 a_3878_13174# VDD 0.29fF
C12209 a_2275_10186# a_23046_10162# 0.71fF
C12210 a_7986_10162# row_n[8] 0.43fF
C12211 m2_20808_18014# col_n[18] 0.33fF
C12212 a_7894_14178# rowon_n[12] 0.14fF
C12213 a_24050_15182# a_25054_15182# 0.86fF
C12214 a_8290_8194# vcm 0.24fF
C12215 a_4882_15182# rowoff_n[13] 0.72fF
C12216 a_17934_4138# rowon_n[2] 0.14fF
C12217 a_25054_8154# m2_25252_8402# 0.19fF
C12218 a_21038_3134# ctop 4.91fF
C12219 a_33086_18194# vcm 0.15fF
C12220 a_18330_9198# col_n[15] 0.11fF
C12221 m2_1046_19620# m3_1046_19620# 0.25fF
C12222 a_29982_8154# VDD 0.29fF
C12223 a_6890_7150# rowoff_n[5] 0.69fF
C12224 a_8898_7150# a_8990_7150# 0.45fF
C12225 a_2275_7174# a_13310_7190# 0.15fF
C12226 a_2475_7174# a_15926_7150# 0.41fF
C12227 a_34394_3174# vcm 0.24fF
C12228 a_15014_17190# a_15014_16186# 0.84fF
C12229 col[27] rowoff_n[13] 0.17fF
C12230 a_15926_5142# rowoff_n[3] 0.59fF
C12231 a_23350_12210# vcm 0.24fF
C12232 col_n[2] rowoff_n[1] 0.32fF
C12233 col_n[5] rowoff_n[4] 0.30fF
C12234 col_n[8] rowoff_n[7] 0.28fF
C12235 col_n[1] rowoff_n[0] 0.33fF
C12236 col_n[6] rowoff_n[5] 0.29fF
C12237 col_n[9] rowoff_n[8] 0.27fF
C12238 col_n[3] rowoff_n[2] 0.32fF
C12239 col_n[10] rowoff_n[9] 0.27fF
C12240 col_n[7] rowoff_n[6] 0.29fF
C12241 col_n[4] rowoff_n[3] 0.31fF
C12242 a_2275_4162# a_6890_4138# 0.17fF
C12243 a_2275_15206# col[31] 0.17fF
C12244 a_10906_11166# VDD 0.29fF
C12245 m2_31852_946# m3_31984_1078# 4.41fF
C12246 a_28066_17190# rowon_n[15] 0.45fF
C12247 a_2275_9182# a_28370_9198# 0.15fF
C12248 a_2475_9182# a_30986_9158# 0.41fF
C12249 a_12002_7150# col[9] 0.38fF
C12250 m2_34864_6970# rowon_n[5] 0.42fF
C12251 a_24962_3134# rowoff_n[1] 0.49fF
C12252 a_16930_6146# vcm 0.18fF
C12253 a_2275_12194# col_n[1] 0.17fF
C12254 a_27062_3134# col_n[24] 0.34fF
C12255 a_2275_1150# col_n[6] 0.17fF
C12256 a_16018_6146# m2_16216_6394# 0.19fF
C12257 a_4274_15222# vcm 0.24fF
C12258 a_2475_18218# a_9902_18194# 0.41fF
C12259 a_1957_5166# VDD 0.28fF
C12260 a_2275_6170# a_21950_6146# 0.17fF
C12261 a_5978_17190# row_n[15] 0.43fF
C12262 a_17022_10162# ctop 4.91fF
C12263 a_25966_15182# VDD 0.29fF
C12264 a_7286_7190# col_n[4] 0.11fF
C12265 a_2966_5142# col[0] 0.38fF
C12266 m2_34864_10986# rowoff_n[9] 1.01fF
C12267 a_23958_11166# a_24050_11166# 0.45fF
C12268 m2_1732_946# vcm 1.11fF
C12269 m2_15788_18014# vcm 0.71fF
C12270 col[11] rowoff_n[14] 0.27fF
C12271 a_16018_7150# row_n[5] 0.43fF
C12272 a_15926_11166# rowon_n[9] 0.14fF
C12273 a_31990_10162# vcm 0.18fF
C12274 a_25054_4138# a_25054_3134# 0.84fF
C12275 a_2475_3158# a_14010_3134# 0.68fF
C12276 a_2275_1150# m2_5748_946# 0.51fF
C12277 a_27062_2130# m2_26832_946# 0.84fF
C12278 m3_34996_4090# ctop 0.22fF
C12279 a_2475_8178# col[11] 0.22fF
C12280 a_32082_14178# ctop 4.91fF
C12281 a_6890_18194# VDD 0.50fF
C12282 a_17022_11166# rowoff_n[9] 1.94fF
C12283 a_2275_17214# a_15014_17190# 0.71fF
C12284 a_10998_17190# col[8] 0.38fF
C12285 a_6982_4138# m2_7180_4386# 0.19fF
C12286 a_2275_14202# col_n[18] 0.17fF
C12287 m2_6752_18014# m2_7180_18442# 0.19fF
C12288 a_12914_13174# vcm 0.18fF
C12289 m2_1732_3958# m3_1864_4090# 4.42fF
C12290 a_2275_3158# col_n[23] 0.17fF
C12291 a_8990_3134# VDD 3.82fF
C12292 a_15014_5142# a_16018_5142# 0.86fF
C12293 a_2475_5166# a_29070_5142# 0.68fF
C12294 a_26058_13174# col_n[23] 0.34fF
C12295 a_2874_5142# rowon_n[3] 0.14fF
C12296 a_2275_18218# a_25054_18194# 0.14fF
C12297 m2_9764_946# m2_10768_946# 0.86fF
C12298 a_13006_17190# ctop 4.93fF
C12299 vcm col_n[8] 3.22fF
C12300 VDD col_n[11] 13.72fF
C12301 a_26058_9158# rowoff_n[7] 1.50fF
C12302 a_4882_14178# a_4974_14178# 0.45fF
C12303 a_2275_14202# a_5278_14218# 0.15fF
C12304 a_2475_14202# a_7894_14178# 0.41fF
C12305 a_2275_11190# col[8] 0.17fF
C12306 a_6282_17230# col_n[3] 0.11fF
C12307 a_33086_15182# rowoff_n[13] 1.15fF
C12308 m2_1732_8978# row_n[7] 0.44fF
C12309 a_2275_2154# a_20034_2130# 0.71fF
C12310 a_27974_17190# vcm 0.18fF
C12311 a_24050_7150# VDD 2.27fF
C12312 a_5978_7150# a_5978_6146# 0.84fF
C12313 a_2475_10186# col[28] 0.22fF
C12314 m2_34864_16006# rowoff_n[14] 1.02fF
C12315 a_14010_14178# row_n[12] 0.43fF
C12316 a_30074_2130# vcm 0.89fF
C12317 a_2275_16210# a_20338_16226# 0.15fF
C12318 a_2475_16210# a_22954_16186# 0.41fF
C12319 a_24050_4138# row_n[2] 0.43fF
C12320 m2_7756_946# col[5] 0.51fF
C12321 a_2275_16210# row_n[14] 26.41fF
C12322 a_23958_8154# rowon_n[6] 0.14fF
C12323 a_2275_4162# a_35094_4138# 0.14fF
C12324 a_4974_10162# VDD 4.23fF
C12325 a_30074_9158# a_31078_9158# 0.86fF
C12326 a_15014_11166# col_n[12] 0.34fF
C12327 a_2275_13198# a_13918_13174# 0.17fF
C12328 a_2275_13198# col[25] 0.17fF
C12329 a_10998_5142# vcm 0.89fF
C12330 a_4974_12170# rowoff_n[10] 2.52fF
C12331 a_19942_18194# a_20034_18194# 0.11fF
C12332 a_2275_2154# col[30] 0.17fF
C12333 a_2275_1150# a_25358_1166# 0.15fF
C12334 a_14922_1126# a_15014_1126# 0.11fF
C12335 a_2475_1150# a_27974_1126# 0.41fF
C12336 m3_14916_18146# VDD 0.10fF
C12337 a_2966_17190# col_n[0] 0.34fF
C12338 a_20034_14178# VDD 2.68fF
C12339 a_21038_11166# a_21038_10162# 0.84fF
C12340 a_2475_10186# a_5978_10162# 0.68fF
C12341 a_10998_2130# rowon_n[0] 0.45fF
C12342 a_2275_15206# a_28978_15182# 0.17fF
C12343 a_26058_9158# vcm 0.89fF
C12344 a_21038_16186# rowoff_n[14] 1.74fF
C12345 a_2966_3134# ctop 4.82fF
C12346 a_10998_12170# a_12002_12170# 0.86fF
C12347 a_2475_12194# a_21038_12170# 0.68fF
C12348 a_22042_11166# row_n[9] 0.43fF
C12349 a_16322_3174# vcm 0.24fF
C12350 a_2475_17214# col[0] 0.20fF
C12351 a_3970_9158# col_n[1] 0.34fF
C12352 a_30378_10202# col_n[27] 0.11fF
C12353 col_n[14] rowoff_n[2] 0.24fF
C12354 col_n[17] rowoff_n[5] 0.21fF
C12355 col_n[20] rowoff_n[8] 0.19fF
C12356 col_n[13] rowoff_n[1] 0.24fF
C12357 col_n[21] rowoff_n[9] 0.19fF
C12358 col_n[18] rowoff_n[6] 0.21fF
C12359 col_n[15] rowoff_n[3] 0.23fF
C12360 col_n[12] rowoff_n[0] 0.25fF
C12361 col_n[19] rowoff_n[7] 0.20fF
C12362 col_n[16] rowoff_n[4] 0.22fF
C12363 a_21950_15182# rowon_n[13] 0.14fF
C12364 a_2475_6170# col[5] 0.22fF
C12365 a_6982_12170# vcm 0.89fF
C12366 a_29982_5142# a_30074_5142# 0.45fF
C12367 a_31990_5142# rowon_n[3] 0.14fF
C12368 a_9902_18194# m2_9764_18014# 0.34fF
C12369 a_2275_9182# a_12002_9158# 0.71fF
C12370 a_2275_12194# col_n[12] 0.17fF
C12371 a_2475_18218# m2_25828_18014# 0.62fF
C12372 a_2275_1150# col_n[17] 0.14fF
C12373 a_31382_7190# vcm 0.24fF
C12374 a_2475_6170# m2_1732_5966# 0.16fF
C12375 a_22042_16186# vcm 0.89fF
C12376 a_24050_8154# col[21] 0.38fF
C12377 a_18938_6146# VDD 0.29fF
C12378 a_2275_6170# a_3878_6146# 0.17fF
C12379 a_2475_6170# a_4882_6146# 0.41fF
C12380 a_2275_9182# col[2] 0.17fF
C12381 a_8990_9158# rowon_n[7] 0.45fF
C12382 col[22] rowoff_n[14] 0.20fF
C12383 m2_1732_11990# rowoff_n[10] 2.46fF
C12384 a_2275_11190# a_27062_11166# 0.71fF
C12385 col_n[5] rowoff_n[10] 0.30fF
C12386 a_24962_1126# vcm 0.18fF
C12387 a_26058_16186# a_27062_16186# 0.86fF
C12388 a_12306_10202# vcm 0.24fF
C12389 a_8990_17190# rowoff_n[15] 2.33fF
C12390 m2_19804_18014# VDD 3.56fF
C12391 a_19334_8194# col_n[16] 0.11fF
C12392 a_2475_8178# col[22] 0.22fF
C12393 a_7894_6146# rowoff_n[4] 0.68fF
C12394 a_25054_5142# ctop 4.91fF
C12395 a_33998_10162# VDD 0.29fF
C12396 a_10906_8154# a_10998_8154# 0.45fF
C12397 a_2275_8178# a_17326_8194# 0.15fF
C12398 a_2475_8178# a_19942_8154# 0.41fF
C12399 a_30074_17190# m2_30272_17438# 0.19fF
C12400 a_2275_14202# col_n[29] 0.17fF
C12401 m2_1732_1950# m2_2160_2378# 0.19fF
C12402 a_5886_4138# vcm 0.18fF
C12403 a_33998_12170# rowoff_n[10] 0.39fF
C12404 a_16930_4138# rowoff_n[2] 0.58fF
C12405 a_30074_8154# row_n[6] 0.43fF
C12406 a_27366_14218# vcm 0.24fF
C12407 a_29982_12170# rowon_n[10] 0.14fF
C12408 a_2275_5166# a_10906_5142# 0.17fF
C12409 VDD col_n[22] 10.98fF
C12410 vcm col_n[19] 3.22fF
C12411 col[6] rowoff_n[15] 0.31fF
C12412 a_5978_8154# ctop 4.91fF
C12413 a_14922_13174# VDD 0.29fF
C12414 a_13006_6146# col[10] 0.38fF
C12415 a_2275_11190# col[19] 0.17fF
C12416 a_2475_10186# a_35002_10162# 0.41fF
C12417 a_2275_10186# a_32386_10202# 0.15fF
C12418 a_25966_2130# rowoff_n[0] 0.48fF
C12419 a_28066_2130# col_n[25] 0.34fF
C12420 a_20946_8154# vcm 0.18fF
C12421 a_2475_2154# a_2874_2130# 0.41fF
C12422 a_1957_2154# a_2275_2154# 0.19fF
C12423 a_8290_17230# vcm 0.24fF
C12424 a_6982_16186# rowon_n[14] 0.45fF
C12425 a_8290_6186# col_n[5] 0.11fF
C12426 a_2275_7174# a_25966_7150# 0.17fF
C12427 a_21038_15182# m2_21236_15430# 0.19fF
C12428 a_21038_12170# ctop 4.91fF
C12429 a_18330_18234# col_n[15] 0.11fF
C12430 m2_1732_1950# rowoff_n[0] 2.46fF
C12431 a_29982_17190# VDD 0.29fF
C12432 m2_1732_17010# rowoff_n[15] 2.46fF
C12433 a_25966_12170# a_26058_12170# 0.45fF
C12434 a_17022_6146# rowon_n[4] 0.45fF
C12435 a_2275_16210# a_3970_16186# 0.71fF
C12436 a_34394_12210# vcm 0.24fF
C12437 a_32082_2130# VDD 1.44fF
C12438 a_27062_5142# a_27062_4138# 0.84fF
C12439 a_2475_4162# a_18026_4138# 0.68fF
C12440 a_5978_17190# m2_5748_18014# 0.84fF
C12441 a_28978_18194# m2_28840_18014# 0.34fF
C12442 a_18026_10162# rowoff_n[8] 1.89fF
C12443 a_12002_16186# col[9] 0.38fF
C12444 a_28066_15182# row_n[13] 0.43fF
C12445 m2_34864_5966# m2_34864_4962# 0.84fF
C12446 a_21950_13174# rowoff_n[11] 0.52fF
C12447 a_2275_1150# a_8990_1126# 0.14fF
C12448 a_16930_15182# vcm 0.18fF
C12449 a_13006_5142# VDD 3.40fF
C12450 a_27062_12170# col_n[24] 0.34fF
C12451 a_12002_13174# m2_12200_13422# 0.19fF
C12452 a_2275_10186# col_n[6] 0.17fF
C12453 a_17022_6146# a_18026_6146# 0.86fF
C12454 a_2475_6170# a_33086_6146# 0.68fF
C12455 a_27062_8154# rowoff_n[6] 1.45fF
C12456 a_1957_14202# VDD 0.28fF
C12457 a_7286_16226# col_n[4] 0.11fF
C12458 a_2475_15206# a_11910_15182# 0.41fF
C12459 a_2275_15206# a_9294_15222# 0.15fF
C12460 a_6890_15182# a_6982_15182# 0.45fF
C12461 a_2966_14178# col[0] 0.38fF
C12462 a_2966_16186# rowoff_n[14] 2.62fF
C12463 a_2275_3158# a_24050_3134# 0.71fF
C12464 a_31078_9158# m2_31276_9406# 0.19fF
C12465 a_2275_1150# m2_28840_946# 0.51fF
C12466 a_28066_9158# VDD 1.85fF
C12467 a_7986_8154# a_7986_7150# 0.84fF
C12468 a_15014_13174# rowon_n[11] 0.45fF
C12469 a_2475_17214# col[11] 0.22fF
C12470 col_n[26] rowoff_n[3] 0.15fF
C12471 col_n[29] rowoff_n[6] 0.13fF
C12472 col_n[25] rowoff_n[2] 0.16fF
C12473 col_n[28] rowoff_n[5] 0.14fF
C12474 col_n[23] rowoff_n[0] 0.17fF
C12475 col_n[30] rowoff_n[7] 0.12fF
C12476 col_n[27] rowoff_n[4] 0.14fF
C12477 col_n[24] rowoff_n[1] 0.16fF
C12478 col_n[31] rowoff_n[8] 0.11fF
C12479 a_2161_12194# a_2275_12194# 0.17fF
C12480 a_2475_12194# a_2966_12170# 0.65fF
C12481 a_2475_6170# col[16] 0.22fF
C12482 a_34090_4138# vcm 0.89fF
C12483 a_25054_3134# rowon_n[1] 0.45fF
C12484 a_2475_17214# a_26970_17190# 0.41fF
C12485 a_2275_17214# a_24354_17230# 0.15fF
C12486 a_3878_15182# rowon_n[13] 0.14fF
C12487 a_8990_12170# VDD 3.82fF
C12488 a_2275_12194# col_n[23] 0.17fF
C12489 a_2275_18218# a_35398_18234# 0.15fF
C12490 a_16018_10162# col_n[13] 0.34fF
C12491 a_32082_10162# a_33086_10162# 0.86fF
C12492 a_2275_1150# col_n[28] 0.17fF
C12493 a_2275_14202# a_17934_14178# 0.17fF
C12494 a_15014_7150# vcm 0.89fF
C12495 a_9902_14178# rowoff_n[12] 0.66fF
C12496 a_16930_2130# a_17022_2130# 0.45fF
C12497 a_2275_2154# a_29374_2170# 0.15fF
C12498 a_2475_2154# a_31990_2130# 0.41fF
C12499 a_22042_7150# m2_22240_7398# 0.19fF
C12500 a_2275_9182# col[13] 0.17fF
C12501 col_n[16] rowoff_n[10] 0.22fF
C12502 a_24050_16186# VDD 2.27fF
C12503 a_2475_11190# a_9994_11166# 0.68fF
C12504 a_23046_12170# a_23046_11166# 0.84fF
C12505 a_5278_1166# vcm 0.25fF
C12506 a_2275_16210# a_32994_16186# 0.17fF
C12507 a_30074_11166# vcm 0.89fF
C12508 a_26970_1126# VDD 0.74fF
C12509 a_25054_17190# m2_24824_18014# 0.84fF
C12510 a_13006_13174# a_14010_13174# 0.86fF
C12511 a_2475_13198# a_25054_13174# 0.68fF
C12512 a_23046_10162# rowon_n[8] 0.45fF
C12513 a_4974_8154# col_n[2] 0.34fF
C12514 a_31382_9198# col_n[28] 0.11fF
C12515 a_20338_5182# vcm 0.24fF
C12516 m2_33284_2378# a_33086_2130# 0.19fF
C12517 sample rowon_n[15] 0.10fF
C12518 vcm col_n[30] 3.24fF
C12519 VDD row_n[15] 4.64fF
C12520 a_13006_5142# m2_13204_5390# 0.19fF
C12521 col[17] rowoff_n[15] 0.23fF
C12522 a_10998_14178# vcm 0.89fF
C12523 a_7894_4138# VDD 0.29fF
C12524 a_2275_11190# col[30] 0.17fF
C12525 a_31990_6146# a_32082_6146# 0.45fF
C12526 vcm rowoff_n[11] 2.43fF
C12527 a_2275_10186# a_16018_10162# 0.71fF
C12528 a_3970_15182# a_3970_14178# 0.84fF
C12529 a_2275_8178# vcm 7.71fF
C12530 a_25054_7150# col[22] 0.38fF
C12531 a_10906_4138# rowon_n[2] 0.14fF
C12532 a_26058_18194# vcm 0.15fF
C12533 a_14010_3134# ctop 4.91fF
C12534 a_22954_8154# VDD 0.29fF
C12535 a_2275_7174# a_6282_7190# 0.15fF
C12536 a_2475_7174# a_8898_7150# 0.41fF
C12537 a_2966_12170# ctop 4.82fF
C12538 a_2275_12194# a_31078_12170# 0.71fF
C12539 a_28978_3134# vcm 0.18fF
C12540 a_28066_17190# a_29070_17190# 0.86fF
C12541 m2_1732_13998# sample 0.31fF
C12542 a_20338_7190# col_n[17] 0.11fF
C12543 a_3970_3134# m2_4168_3382# 0.19fF
C12544 a_16322_12210# vcm 0.24fF
C12545 a_8898_5142# rowoff_n[3] 0.67fF
C12546 a_2475_15206# col[5] 0.22fF
C12547 a_29070_7150# ctop 4.91fF
C12548 a_2475_4162# col[10] 0.22fF
C12549 m3_31984_18146# m3_32988_18146# 0.21fF
C12550 a_21038_17190# rowon_n[15] 0.45fF
C12551 a_12914_9158# a_13006_9158# 0.45fF
C12552 a_2475_9182# a_23958_9158# 0.41fF
C12553 a_2275_9182# a_21342_9198# 0.15fF
C12554 m2_1732_10986# rowon_n[9] 0.43fF
C12555 a_17934_3134# rowoff_n[1] 0.57fF
C12556 a_31078_7150# rowon_n[5] 0.45fF
C12557 a_9902_6146# vcm 0.18fF
C12558 a_3878_13174# rowoff_n[11] 0.73fF
C12559 a_2275_10186# col_n[17] 0.17fF
C12560 a_31382_16226# vcm 0.24fF
C12561 a_14010_5142# col[11] 0.38fF
C12562 a_2275_6170# a_14922_6146# 0.17fF
C12563 m2_33860_946# col_n[31] 0.74fF
C12564 a_9994_10162# ctop 4.91fF
C12565 a_24050_17190# col[21] 0.38fF
C12566 a_18938_15182# VDD 0.29fF
C12567 a_2966_11166# a_2966_10162# 0.84fF
C12568 m2_1732_18014# vcm 1.11fF
C12569 a_8990_7150# row_n[5] 0.43fF
C12570 a_2275_7174# col[7] 0.17fF
C12571 a_8898_11166# rowon_n[9] 0.14fF
C12572 a_24962_10162# vcm 0.18fF
C12573 a_9294_5182# col_n[6] 0.11fF
C12574 a_3970_3134# a_4974_3134# 0.86fF
C12575 a_2475_3158# a_6982_3134# 0.68fF
C12576 a_19334_17230# col_n[16] 0.11fF
C12577 a_2475_17214# col[22] 0.22fF
C12578 a_2275_8178# a_29982_8154# 0.17fF
C12579 a_25054_14178# ctop 4.91fF
C12580 a_2475_6170# col[27] 0.22fF
C12581 a_27974_13174# a_28066_13174# 0.45fF
C12582 a_9994_11166# rowoff_n[9] 2.28fF
C12583 a_2275_17214# a_7986_17190# 0.71fF
C12584 a_5886_13174# vcm 0.18fF
C12585 a_2475_3158# VDD 41.96fF
C12586 a_29070_6146# a_29070_5142# 0.84fF
C12587 a_2475_5166# a_22042_5142# 0.68fF
C12588 a_2275_18218# a_18026_18194# 0.14fF
C12589 a_5978_17190# ctop 4.93fF
C12590 a_19030_9158# rowoff_n[7] 1.84fF
C12591 a_13006_15182# col[10] 0.38fF
C12592 a_29070_14178# rowon_n[12] 0.45fF
C12593 a_2275_9182# col[24] 0.17fF
C12594 a_26058_15182# rowoff_n[13] 1.50fF
C12595 a_2275_2154# a_13006_2130# 0.71fF
C12596 a_28066_11166# col_n[25] 0.34fF
C12597 a_20946_17190# vcm 0.18fF
C12598 m2_29844_18014# m3_29976_18146# 4.43fF
C12599 col_n[27] rowoff_n[10] 0.14fF
C12600 a_17022_7150# VDD 2.99fF
C12601 a_28066_7150# rowoff_n[5] 1.40fF
C12602 a_19030_7150# a_20034_7150# 0.86fF
C12603 a_8290_15222# col_n[5] 0.11fF
C12604 a_6982_14178# row_n[12] 0.43fF
C12605 a_23046_2130# vcm 0.89fF
C12606 a_8898_16186# a_8990_16186# 0.45fF
C12607 a_2475_16210# a_15926_16186# 0.41fF
C12608 a_2275_16210# a_13310_16226# 0.15fF
C12609 a_17022_4138# row_n[2] 0.43fF
C12610 a_16930_8154# rowon_n[6] 0.14fF
C12611 a_2275_4162# a_28066_4138# 0.71fF
C12612 a_32082_11166# VDD 1.44fF
C12613 m3_21944_1078# m3_22948_1078# 0.21fF
C12614 a_9994_9158# a_9994_8154# 0.84fF
C12615 a_2275_13198# a_6890_13174# 0.17fF
C12616 col_n[3] rowon_n[12] 0.17fF
C12617 sample row_n[10] 0.92fF
C12618 VDD rowon_n[9] 4.61fF
C12619 col_n[2] row_n[12] 0.37fF
C12620 col_n[6] row_n[14] 0.37fF
C12621 col_n[4] row_n[13] 0.37fF
C12622 col_n[1] rowon_n[11] 0.17fF
C12623 col_n[8] row_n[15] 0.37fF
C12624 col_n[5] rowon_n[13] 0.17fF
C12625 col_n[0] rowon_n[10] 0.17fF
C12626 col_n[7] rowon_n[14] 0.17fF
C12627 col_n[9] rowon_n[15] 0.17fF
C12628 vcm row_n[11] 1.08fF
C12629 col[28] rowoff_n[15] 0.16fF
C12630 a_3970_5142# vcm 0.89fF
C12631 a_2475_2154# col[4] 0.22fF
C12632 col_n[11] rowoff_n[11] 0.26fF
C12633 a_2275_1150# a_18330_1166# 0.19fF
C12634 a_2475_1150# a_20946_1126# 0.41fF
C12635 a_17022_9158# col_n[14] 0.34fF
C12636 a_13006_14178# VDD 3.40fF
C12637 a_3970_2130# rowon_n[0] 0.45fF
C12638 a_2275_8178# col_n[11] 0.17fF
C12639 a_2275_15206# a_21950_15182# 0.17fF
C12640 a_19030_9158# vcm 0.89fF
C12641 a_14010_16186# rowoff_n[14] 2.08fF
C12642 a_18938_3134# a_19030_3134# 0.45fF
C12643 a_2275_3158# a_33390_3174# 0.15fF
C12644 a_27062_16186# m2_27260_16434# 0.19fF
C12645 a_2275_5166# col[1] 0.17fF
C12646 a_2475_12194# a_14010_12170# 0.68fF
C12647 a_25054_13174# a_25054_12170# 0.84fF
C12648 a_15014_11166# row_n[9] 0.43fF
C12649 a_9294_3174# vcm 0.24fF
C12650 a_14922_15182# rowon_n[13] 0.14fF
C12651 a_2475_15206# col[16] 0.22fF
C12652 a_34090_13174# vcm 0.89fF
C12653 a_2475_4162# col[21] 0.22fF
C12654 a_30986_3134# VDD 0.29fF
C12655 a_24962_5142# rowon_n[3] 0.14fF
C12656 m2_32856_946# m2_33860_946# 0.86fF
C12657 a_3878_9158# a_3970_9158# 0.45fF
C12658 a_2275_9182# a_4974_9158# 0.71fF
C12659 a_2966_17190# rowon_n[15] 0.45fF
C12660 a_5978_7150# col_n[3] 0.34fF
C12661 a_32386_8194# col_n[29] 0.11fF
C12662 a_2475_18218# m2_11772_18014# 0.62fF
C12663 a_2475_14202# a_29070_14178# 0.68fF
C12664 a_15014_14178# a_16018_14178# 0.86fF
C12665 a_2275_10186# col_n[28] 0.17fF
C12666 a_24354_7190# vcm 0.24fF
C12667 a_15014_16186# vcm 0.89fF
C12668 a_11910_6146# VDD 0.29fF
C12669 a_18026_14178# m2_18224_14426# 0.19fF
C12670 a_33998_7150# a_34090_7150# 0.45fF
C12671 a_2475_9182# rowon_n[7] 0.40fF
C12672 a_2275_7174# col[18] 0.17fF
C12673 a_2275_11190# a_20034_11166# 0.71fF
C12674 a_17934_1126# vcm 0.18fF
C12675 a_5978_16186# a_5978_15182# 0.84fF
C12676 a_26058_6146# col[23] 0.38fF
C12677 a_15014_2130# m2_15212_2378# 0.19fF
C12678 a_5278_10202# vcm 0.24fF
C12679 a_2475_17214# rowoff_n[15] 4.75fF
C12680 row_n[6] rowoff_n[6] 0.64fF
C12681 m2_5748_18014# VDD 4.97fF
C12682 a_18026_5142# ctop 4.91fF
C12683 a_9994_2130# m2_9764_946# 0.84fF
C12684 a_26970_10162# VDD 0.29fF
C12685 a_2475_8178# a_12914_8154# 0.41fF
C12686 a_2275_8178# a_10298_8194# 0.15fF
C12687 a_2275_13198# a_35094_13174# 0.14fF
C12688 a_21342_6186# col_n[18] 0.11fF
C12689 a_32994_5142# vcm 0.18fF
C12690 a_26970_12170# rowoff_n[10] 0.47fF
C12691 a_9902_4138# rowoff_n[2] 0.66fF
C12692 a_31382_18234# col_n[28] 0.11fF
C12693 a_4974_17190# col_n[2] 0.34fF
C12694 a_23046_8154# row_n[6] 0.43fF
C12695 a_20338_14218# vcm 0.24fF
C12696 a_22954_12170# rowon_n[10] 0.14fF
C12697 a_2874_5142# a_2966_5142# 0.45fF
C12698 a_8990_12170# m2_9188_12418# 0.19fF
C12699 a_33086_9158# ctop 4.91fF
C12700 a_7894_13174# VDD 0.29fF
C12701 a_2475_10186# a_27974_10162# 0.41fF
C12702 a_2275_10186# a_25358_10202# 0.15fF
C12703 a_14922_10162# a_15014_10162# 0.45fF
C12704 a_18938_2130# rowoff_n[0] 0.56fF
C12705 a_32994_2130# rowon_n[0] 0.14fF
C12706 a_13918_8154# vcm 0.18fF
C12707 a_15014_4138# col[12] 0.38fF
C12708 a_16018_3134# a_16018_2130# 0.84fF
C12709 a_28066_8154# m2_28264_8402# 0.19fF
C12710 a_2275_17214# vcm 7.71fF
C12711 a_25054_16186# col[22] 0.38fF
C12712 a_2275_6170# col_n[5] 0.17fF
C12713 a_2275_7174# a_18938_7150# 0.17fF
C12714 a_14010_12170# ctop 4.91fF
C12715 a_22954_17190# VDD 0.29fF
C12716 a_9994_6146# rowon_n[4] 0.45fF
C12717 a_28978_12170# vcm 0.18fF
C12718 a_10298_4178# col_n[7] 0.11fF
C12719 a_25054_2130# VDD 2.16fF
C12720 a_20338_16226# col_n[17] 0.11fF
C12721 a_5978_4138# a_6982_4138# 0.86fF
C12722 a_2475_4162# a_10998_4138# 0.68fF
C12723 m3_34996_9110# m3_34996_8106# 0.20fF
C12724 col_n[19] row_n[15] 0.37fF
C12725 col_n[17] row_n[14] 0.37fF
C12726 col_n[15] row_n[13] 0.37fF
C12727 VDD row_n[4] 4.64fF
C12728 col_n[14] rowon_n[12] 0.17fF
C12729 col_n[16] rowon_n[13] 0.17fF
C12730 col_n[5] row_n[8] 0.37fF
C12731 col_n[11] row_n[11] 0.37fF
C12732 col_n[3] row_n[7] 0.37fF
C12733 col_n[7] row_n[9] 0.37fF
C12734 col_n[18] rowon_n[14] 0.17fF
C12735 col_n[9] row_n[10] 0.37fF
C12736 col_n[2] rowon_n[6] 0.17fF
C12737 col_n[20] rowon_n[15] 0.17fF
C12738 col_n[4] rowon_n[7] 0.17fF
C12739 sample rowon_n[4] 0.10fF
C12740 col_n[12] rowon_n[11] 0.17fF
C12741 col_n[13] row_n[12] 0.37fF
C12742 col_n[6] rowon_n[8] 0.17fF
C12743 vcm rowon_n[5] 0.91fF
C12744 col_n[8] rowon_n[9] 0.17fF
C12745 col_n[0] row_n[5] 0.37fF
C12746 col_n[1] row_n[6] 0.37fF
C12747 col_n[10] rowon_n[10] 0.17fF
C12748 a_2275_9182# a_33998_9158# 0.17fF
C12749 a_29070_16186# ctop 4.91fF
C12750 a_2475_13198# col[10] 0.22fF
C12751 a_29982_14178# a_30074_14178# 0.45fF
C12752 a_2475_2154# col[15] 0.22fF
C12753 a_10998_10162# rowoff_n[8] 2.23fF
C12754 col_n[22] rowoff_n[11] 0.18fF
C12755 a_21038_15182# row_n[13] 0.43fF
C12756 a_14922_13174# rowoff_n[11] 0.60fF
C12757 m2_34864_2954# VDD 1.58fF
C12758 a_1957_1150# a_2161_1150# 0.11fF
C12759 a_2475_1150# a_2275_1150# 2.86fF
C12760 a_19030_6146# m2_19228_6394# 0.19fF
C12761 a_9902_15182# vcm 0.18fF
C12762 a_5978_5142# VDD 4.13fF
C12763 a_31078_5142# row_n[3] 0.43fF
C12764 m2_2736_1950# col[0] 0.37fF
C12765 a_2475_6170# a_26058_6146# 0.68fF
C12766 a_31078_7150# a_31078_6146# 0.84fF
C12767 a_3970_2130# col[1] 0.38fF
C12768 a_30986_9158# rowon_n[7] 0.14fF
C12769 a_2275_8178# col_n[22] 0.17fF
C12770 a_20034_8154# rowoff_n[6] 1.79fF
C12771 a_14010_14178# col[11] 0.38fF
C12772 a_2475_15206# a_4882_15182# 0.41fF
C12773 a_2275_15206# a_3878_15182# 0.17fF
C12774 a_29070_10162# col_n[26] 0.34fF
C12775 a_30986_17190# rowoff_n[15] 0.42fF
C12776 a_2275_16210# col[7] 0.17fF
C12777 a_29070_6146# rowoff_n[4] 1.35fF
C12778 a_2275_5166# col[12] 0.17fF
C12779 a_2275_3158# a_17022_3134# 0.71fF
C12780 a_2475_1150# m2_14784_946# 0.62fF
C12781 a_21038_9158# VDD 2.58fF
C12782 m3_10900_1078# ctop 0.21fF
C12783 m2_14784_18014# col_n[12] 0.32fF
C12784 a_9294_14218# col_n[6] 0.11fF
C12785 a_21038_8154# a_22042_8154# 0.86fF
C12786 a_7986_13174# rowon_n[11] 0.45fF
C12787 col_n[6] rowoff_n[12] 0.29fF
C12788 a_2475_15206# col[27] 0.22fF
C12789 a_27062_4138# vcm 0.89fF
C12790 a_18026_3134# rowon_n[1] 0.45fF
C12791 a_10906_17190# a_10998_17190# 0.45fF
C12792 a_2475_17214# a_19942_17190# 0.41fF
C12793 a_2275_17214# a_17326_17230# 0.15fF
C12794 a_9994_4138# m2_10192_4386# 0.19fF
C12795 a_2275_5166# a_32082_5142# 0.71fF
C12796 a_2475_12194# VDD 41.96fF
C12797 a_2275_18218# a_27366_18234# 0.15fF
C12798 m2_13780_946# m2_14208_1374# 0.19fF
C12799 a_12002_10162# a_12002_9158# 0.84fF
C12800 a_2275_14202# a_10906_14178# 0.17fF
C12801 a_7986_7150# vcm 0.89fF
C12802 a_2161_14202# rowoff_n[12] 0.14fF
C12803 a_29070_12170# row_n[10] 0.43fF
C12804 a_2275_2154# a_22346_2170# 0.15fF
C12805 a_2475_2154# a_24962_2130# 0.41fF
C12806 a_18026_8154# col_n[15] 0.34fF
C12807 a_28978_16186# rowon_n[14] 0.14fF
C12808 a_2275_7174# col[29] 0.17fF
C12809 a_17022_16186# VDD 2.99fF
C12810 a_1957_11190# a_2275_11190# 0.19fF
C12811 a_2475_11190# a_2874_11166# 0.41fF
C12812 a_32386_2170# vcm 0.24fF
C12813 rowon_n[2] rowoff_n[2] 20.66fF
C12814 a_2275_16210# a_25966_16186# 0.17fF
C12815 a_2275_4162# col_n[0] 0.17fF
C12816 a_23046_11166# vcm 0.89fF
C12817 a_19942_1126# VDD 0.71fF
C12818 a_20946_4138# a_21038_4138# 0.45fF
C12819 a_16018_10162# rowon_n[8] 0.45fF
C12820 a_27062_14178# a_27062_13174# 0.84fF
C12821 a_2475_13198# a_18026_13174# 0.68fF
C12822 a_13310_5182# vcm 0.24fF
C12823 m2_8760_946# vcm 0.71fF
C12824 a_2275_1150# a_30986_1126# 0.17fF
C12825 a_3970_14178# vcm 0.89fF
C12826 a_35002_5142# VDD 0.36fF
C12827 a_2475_11190# col[4] 0.22fF
C12828 a_6982_6146# col_n[4] 0.34fF
C12829 a_33390_7190# col_n[30] 0.11fF
C12830 a_2275_10186# a_8990_10162# 0.71fF
C12831 a_17022_15182# a_18026_15182# 0.86fF
C12832 a_2475_15206# a_33086_15182# 0.68fF
C12833 a_2275_17214# col_n[11] 0.17fF
C12834 a_28370_9198# vcm 0.24fF
C12835 a_2275_6170# col_n[16] 0.17fF
C12836 a_6982_3134# ctop 4.91fF
C12837 a_19030_18194# vcm 0.15fF
C12838 a_15926_8154# VDD 0.29fF
C12839 a_2275_12194# a_24050_12170# 0.71fF
C12840 a_2275_14202# col[1] 0.17fF
C12841 a_27062_5142# col[24] 0.38fF
C12842 a_21950_3134# vcm 0.18fF
C12843 a_2275_3158# col[6] 0.17fF
C12844 a_7986_17190# a_7986_16186# 0.84fF
C12845 a_9294_12210# vcm 0.24fF
C12846 col_n[29] rowon_n[14] 0.17fF
C12847 col_n[11] rowon_n[5] 0.17fF
C12848 col_n[18] row_n[9] 0.37fF
C12849 col_n[27] rowon_n[13] 0.17fF
C12850 col_n[9] rowon_n[4] 0.17fF
C12851 col_n[16] row_n[8] 0.37fF
C12852 col_n[22] row_n[11] 0.37fF
C12853 col_n[7] rowon_n[3] 0.17fF
C12854 col_n[14] row_n[7] 0.37fF
C12855 col_n[5] rowon_n[2] 0.17fF
C12856 col_n[30] row_n[15] 0.37fF
C12857 col_n[12] row_n[6] 0.37fF
C12858 col_n[3] rowon_n[1] 0.17fF
C12859 col_n[28] row_n[14] 0.37fF
C12860 col_n[10] row_n[5] 0.37fF
C12861 col_n[26] row_n[13] 0.37fF
C12862 col_n[24] row_n[12] 0.37fF
C12863 col_n[23] rowon_n[11] 0.17fF
C12864 col_n[15] rowon_n[7] 0.17fF
C12865 col_n[31] rowon_n[15] 0.17fF
C12866 col_n[20] row_n[10] 0.37fF
C12867 col_n[13] rowon_n[6] 0.17fF
C12868 col_n[1] rowon_n[0] 0.17fF
C12869 col_n[17] rowon_n[8] 0.17fF
C12870 col_n[19] rowon_n[9] 0.17fF
C12871 col_n[21] rowon_n[10] 0.17fF
C12872 col_n[2] row_n[1] 0.37fF
C12873 col_n[4] row_n[2] 0.37fF
C12874 col_n[25] rowon_n[12] 0.17fF
C12875 col_n[6] row_n[3] 0.37fF
C12876 vcm row_n[0] 1.06fF
C12877 VDD ctop 10.52fF
C12878 col_n[8] row_n[4] 0.37fF
C12879 a_22042_7150# ctop 4.91fF
C12880 a_2475_13198# col[21] 0.22fF
C12881 a_30986_12170# VDD 0.29fF
C12882 m3_17928_18146# m3_18932_18146# 0.21fF
C12883 a_2475_2154# col[26] 0.22fF
C12884 a_2475_9182# a_16930_9158# 0.41fF
C12885 a_2275_9182# a_14314_9198# 0.15fF
C12886 a_14010_17190# rowon_n[15] 0.45fF
C12887 m2_1732_8978# sample_n 0.12fF
C12888 a_22346_5182# col_n[19] 0.11fF
C12889 a_10906_3134# rowoff_n[1] 0.65fF
C12890 a_5978_16186# col_n[3] 0.34fF
C12891 a_32386_17230# col_n[29] 0.11fF
C12892 a_2966_15182# row_n[13] 0.41fF
C12893 a_24050_7150# rowon_n[5] 0.45fF
C12894 a_31078_14178# rowoff_n[12] 1.25fF
C12895 a_27062_2130# a_28066_2130# 0.86fF
C12896 a_24354_16226# vcm 0.24fF
C12897 a_2275_6170# a_7894_6146# 0.17fF
C12898 a_11910_15182# VDD 0.29fF
C12899 a_1957_8178# rowoff_n[6] 0.14fF
C12900 a_2275_11190# a_29374_11206# 0.15fF
C12901 a_2475_11190# a_31990_11166# 0.41fF
C12902 a_16930_11166# a_17022_11166# 0.45fF
C12903 a_2275_16210# col[18] 0.17fF
C12904 a_2475_7174# row_n[5] 0.48fF
C12905 a_2275_5166# col[23] 0.17fF
C12906 a_17934_10162# vcm 0.18fF
C12907 a_16018_3134# col[13] 0.38fF
C12908 a_26058_15182# col[23] 0.38fF
C12909 a_18026_4138# a_18026_3134# 0.84fF
C12910 a_2966_9158# VDD 4.45fF
C12911 m3_6884_18146# ctop 0.21fF
C12912 col_n[17] rowoff_n[12] 0.21fF
C12913 a_33086_17190# m2_33284_17438# 0.19fF
C12914 a_2275_8178# a_22954_8154# 0.17fF
C12915 a_18026_14178# ctop 4.91fF
C12916 a_11302_3174# col_n[8] 0.11fF
C12917 a_2874_11166# rowoff_n[9] 0.74fF
C12918 a_21342_15222# col_n[18] 0.11fF
C12919 a_32994_14178# vcm 0.18fF
C12920 a_29070_4138# VDD 1.75fF
C12921 a_7986_5142# a_8990_5142# 0.86fF
C12922 a_2475_5166# a_15014_5142# 0.68fF
C12923 a_2275_18218# a_10998_18194# 0.14fF
C12924 m2_33860_946# sw 0.38fF
C12925 a_12002_9158# rowoff_n[7] 2.18fF
C12926 a_22042_14178# rowon_n[12] 0.45fF
C12927 a_31990_15182# a_32082_15182# 0.45fF
C12928 m2_1732_8978# m2_1732_7974# 0.84fF
C12929 a_19030_15182# rowoff_n[13] 1.84fF
C12930 a_32082_4138# rowon_n[2] 0.45fF
C12931 a_2275_2154# a_5978_2130# 0.71fF
C12932 a_13918_17190# vcm 0.18fF
C12933 col_n[1] rowoff_n[13] 0.33fF
C12934 a_9994_7150# VDD 3.71fF
C12935 a_21038_7150# rowoff_n[5] 1.74fF
C12936 a_24050_15182# m2_24248_15430# 0.19fF
C12937 a_15014_13174# col[12] 0.38fF
C12938 a_2475_7174# a_30074_7150# 0.68fF
C12939 a_33086_8154# a_33086_7150# 0.84fF
C12940 col[4] rowoff_n[9] 0.32fF
C12941 col[3] rowoff_n[8] 0.33fF
C12942 col[2] rowoff_n[7] 0.33fF
C12943 col[1] rowoff_n[6] 0.34fF
C12944 col[0] rowoff_n[5] 0.34fF
C12945 a_2275_15206# col_n[5] 0.17fF
C12946 a_2275_4162# col_n[10] 0.17fF
C12947 a_16018_2130# vcm 0.89fF
C12948 a_30074_9158# col_n[27] 0.34fF
C12949 a_2475_16210# a_8898_16186# 0.41fF
C12950 a_2275_16210# a_6282_16226# 0.15fF
C12951 a_30074_5142# rowoff_n[3] 1.30fF
C12952 a_9994_4138# row_n[2] 0.43fF
C12953 a_35398_2170# VDD 0.12fF
C12954 a_9902_8154# rowon_n[6] 0.14fF
C12955 a_2475_10186# m2_34864_9982# 0.56fF
C12956 a_2275_4162# a_21038_4138# 0.71fF
C12957 a_10298_13214# col_n[7] 0.11fF
C12958 a_25054_11166# VDD 2.16fF
C12959 m3_7888_1078# m3_8892_1078# 0.21fF
C12960 a_2275_1150# col[0] 0.16fF
C12961 a_23046_9158# a_24050_9158# 0.86fF
C12962 m2_34864_3958# vcm 0.72fF
C12963 a_31078_6146# vcm 0.89fF
C12964 a_12914_18194# a_13006_18194# 0.11fF
C12965 a_2475_11190# col[15] 0.22fF
C12966 a_7894_1126# a_7986_1126# 0.11fF
C12967 a_2275_1150# a_11302_1166# 0.15fF
C12968 a_2475_1150# a_13918_1126# 0.41fF
C12969 m2_12776_946# VDD 5.80fF
C12970 a_15014_13174# m2_15212_13422# 0.19fF
C12971 a_5978_14178# VDD 4.13fF
C12972 a_14010_11166# a_14010_10162# 0.84fF
C12973 a_3970_11166# col[1] 0.38fF
C12974 a_2275_17214# col_n[22] 0.17fF
C12975 a_2275_6170# col_n[27] 0.17fF
C12976 a_2275_15206# a_14922_15182# 0.17fF
C12977 a_2275_18218# col_n[7] 0.17fF
C12978 a_30074_11166# rowon_n[9] 0.45fF
C12979 a_12002_9158# vcm 0.89fF
C12980 a_6982_16186# rowoff_n[14] 2.42fF
C12981 a_19030_7150# col_n[16] 0.34fF
C12982 a_34090_9158# m2_34288_9406# 0.19fF
C12983 a_2475_3158# a_28978_3134# 0.41fF
C12984 a_2275_3158# a_26362_3174# 0.15fF
C12985 a_2275_14202# col[12] 0.17fF
C12986 a_1957_18218# sample 0.35fF
C12987 a_2275_3158# col[17] 0.17fF
C12988 a_2475_12194# a_6982_12170# 0.68fF
C12989 a_3970_12170# a_4974_12170# 0.86fF
C12990 a_7986_11166# row_n[9] 0.43fF
C12991 a_3878_3134# vcm 0.18fF
C12992 a_31990_11166# rowoff_n[9] 0.41fF
C12993 a_2275_17214# a_29982_17190# 0.17fF
C12994 col_n[1] col[1] 0.43fF
C12995 col_n[28] rowon_n[8] 0.17fF
C12996 col_n[26] rowon_n[7] 0.17fF
C12997 col_n[24] rowon_n[6] 0.17fF
C12998 col_n[31] row_n[10] 0.37fF
C12999 col_n[22] rowon_n[5] 0.17fF
C13000 col_n[29] row_n[9] 0.37fF
C13001 col_n[20] rowon_n[4] 0.17fF
C13002 col_n[27] row_n[8] 0.37fF
C13003 col_n[18] rowon_n[3] 0.17fF
C13004 col_n[13] row_n[1] 0.37fF
C13005 VDD col[5] 12.19fF
C13006 col_n[11] row_n[0] 0.37fF
C13007 col_n[30] rowon_n[9] 0.17fF
C13008 col_n[15] row_n[2] 0.37fF
C13009 col_n[17] row_n[3] 0.37fF
C13010 vcm col[2] 6.66fF
C13011 col_n[19] row_n[4] 0.37fF
C13012 col_n[12] rowon_n[0] 0.17fF
C13013 col_n[21] row_n[5] 0.37fF
C13014 col_n[14] rowon_n[1] 0.17fF
C13015 col_n[23] row_n[6] 0.37fF
C13016 col_n[16] rowon_n[2] 0.17fF
C13017 col_n[25] row_n[7] 0.37fF
C13018 a_7894_15182# rowon_n[13] 0.14fF
C13019 a_27062_13174# vcm 0.89fF
C13020 a_23958_3134# VDD 0.29fF
C13021 a_22954_5142# a_23046_5142# 0.45fF
C13022 a_5978_11166# m2_6176_11414# 0.19fF
C13023 m2_29844_18014# col[27] 0.39fF
C13024 a_17934_5142# rowon_n[3] 0.14fF
C13025 m2_25828_946# m2_26832_946# 0.86fF
C13026 a_29070_15182# a_29070_14178# 0.84fF
C13027 a_2475_14202# a_22042_14178# 0.68fF
C13028 a_17326_7190# vcm 0.24fF
C13029 m2_1732_5966# VDD 5.46fF
C13030 a_25054_7150# m2_25252_7398# 0.19fF
C13031 a_2275_2154# a_35002_2130# 0.17fF
C13032 a_30074_2130# ctop 4.93fF
C13033 a_7986_16186# vcm 0.89fF
C13034 a_4882_6146# VDD 0.29fF
C13035 a_7986_5142# col_n[5] 0.34fF
C13036 a_18026_17190# col_n[15] 0.34fF
C13037 a_2275_16210# col[29] 0.17fF
C13038 a_2275_11190# a_13006_11166# 0.71fF
C13039 a_10906_1126# vcm 0.18fF
C13040 a_19030_16186# a_20034_16186# 0.86fF
C13041 a_32386_11206# vcm 0.24fF
C13042 a_30474_1488# VDD 0.12fF
C13043 col_n[28] rowoff_n[12] 0.14fF
C13044 a_2275_13198# col_n[0] 0.17fF
C13045 a_10998_5142# ctop 4.91fF
C13046 a_2275_2154# col_n[4] 0.17fF
C13047 a_19942_10162# VDD 0.29fF
C13048 a_2475_8178# a_5886_8154# 0.41fF
C13049 a_2275_8178# a_3270_8194# 0.15fF
C13050 a_28066_4138# col[25] 0.38fF
C13051 a_2275_13198# a_28066_13174# 0.71fF
C13052 a_25966_5142# vcm 0.18fF
C13053 a_2161_4162# rowoff_n[2] 0.14fF
C13054 a_19942_12170# rowoff_n[10] 0.55fF
C13055 m2_31852_946# vcm 0.71fF
C13056 a_2275_18218# m2_28840_18014# 0.51fF
C13057 a_16018_5142# m2_16216_5390# 0.19fF
C13058 a_16018_8154# row_n[6] 0.43fF
C13059 a_13310_14218# vcm 0.24fF
C13060 a_15926_12170# rowon_n[10] 0.14fF
C13061 a_26058_9158# ctop 4.91fF
C13062 a_35002_14178# VDD 0.36fF
C13063 a_23350_4178# col_n[20] 0.11fF
C13064 a_2275_10186# a_18330_10202# 0.15fF
C13065 a_2475_10186# a_20946_10162# 0.41fF
C13066 a_11910_2130# rowoff_n[0] 0.64fF
C13067 a_25966_2130# rowon_n[0] 0.14fF
C13068 a_2475_9182# col[9] 0.22fF
C13069 a_6982_15182# col_n[4] 0.34fF
C13070 a_33390_16226# col_n[30] 0.11fF
C13071 a_6890_8154# vcm 0.18fF
C13072 col_n[12] rowoff_n[13] 0.25fF
C13073 a_29070_3134# a_30074_3134# 0.86fF
C13074 a_28370_18234# vcm 0.25fF
C13075 col[15] rowoff_n[9] 0.25fF
C13076 col[14] rowoff_n[8] 0.25fF
C13077 col[13] rowoff_n[7] 0.26fF
C13078 col[12] rowoff_n[6] 0.27fF
C13079 col[11] rowoff_n[5] 0.27fF
C13080 col[10] rowoff_n[4] 0.28fF
C13081 col[9] rowoff_n[3] 0.29fF
C13082 col[8] rowoff_n[2] 0.29fF
C13083 col[7] rowoff_n[1] 0.30fF
C13084 col[6] rowoff_n[0] 0.31fF
C13085 a_2275_15206# col_n[16] 0.17fF
C13086 a_2966_7150# rowoff_n[5] 2.62fF
C13087 a_2275_7174# a_11910_7150# 0.17fF
C13088 a_6982_12170# ctop 4.91fF
C13089 a_2275_4162# col_n[21] 0.17fF
C13090 m2_1732_1950# rowon_n[0] 0.43fF
C13091 a_15926_17190# VDD 0.29fF
C13092 a_2275_12194# a_33390_12210# 0.15fF
C13093 a_18938_12170# a_19030_12170# 0.45fF
C13094 a_2874_6146# rowon_n[4] 0.14fF
C13095 a_17022_2130# col[14] 0.38fF
C13096 a_27062_14178# col[24] 0.38fF
C13097 a_6982_3134# m2_7180_3382# 0.19fF
C13098 a_21950_12170# vcm 0.18fF
C13099 a_2275_12194# col[6] 0.17fF
C13100 a_18026_2130# VDD 2.89fF
C13101 a_2275_1150# col[11] 0.17fF
C13102 a_2275_4162# a_2966_4138# 0.67fF
C13103 a_2475_4162# a_3970_4138# 0.68fF
C13104 a_20034_5142# a_20034_4138# 0.84fF
C13105 m3_34996_16138# m3_34996_15134# 0.20fF
C13106 a_2275_9182# a_26970_9158# 0.17fF
C13107 a_22042_16186# ctop 4.91fF
C13108 a_2475_11190# col[26] 0.22fF
C13109 a_12306_2170# col_n[9] 0.11fF
C13110 a_3970_10162# rowoff_n[8] 2.57fF
C13111 a_14010_15182# row_n[13] 0.43fF
C13112 a_22346_14218# col_n[19] 0.11fF
C13113 a_7894_13174# rowoff_n[11] 0.68fF
C13114 a_3878_18194# a_3970_18194# 0.11fF
C13115 a_33086_6146# VDD 1.34fF
C13116 a_24050_5142# row_n[3] 0.43fF
C13117 a_2475_6170# a_19030_6146# 0.68fF
C13118 a_9994_6146# a_10998_6146# 0.86fF
C13119 a_2275_17214# row_n[15] 26.41fF
C13120 a_23958_9158# rowon_n[7] 0.14fF
C13121 a_13006_8154# rowoff_n[6] 2.13fF
C13122 a_2275_18218# col_n[18] 0.17fF
C13123 a_33998_16186# a_34090_16186# 0.45fF
C13124 a_23958_17190# rowoff_n[15] 0.50fF
C13125 a_2275_14202# col[23] 0.17fF
C13126 a_22042_6146# rowoff_n[4] 1.69fF
C13127 a_2275_3158# a_9994_3134# 0.71fF
C13128 a_16018_12170# col[13] 0.38fF
C13129 a_2275_3158# col[28] 0.17fF
C13130 a_14010_9158# VDD 3.30fF
C13131 m3_1864_10114# ctop 0.22fF
C13132 a_2475_8178# a_34090_8154# 0.68fF
C13133 col_n[26] row_n[2] 0.37fF
C13134 col_n[24] row_n[1] 0.37fF
C13135 col_n[22] row_n[0] 0.37fF
C13136 vcm col[13] 6.66fF
C13137 rowon_n[10] row_n[10] 21.02fF
C13138 col_n[23] rowon_n[0] 0.17fF
C13139 col_n[30] row_n[4] 0.37fF
C13140 col_n[28] row_n[3] 0.37fF
C13141 col_n[25] rowon_n[1] 0.17fF
C13142 col_n[16] en_bit_n[2] 0.19fF
C13143 col_n[27] rowon_n[2] 0.17fF
C13144 col_n[6] col[7] 6.22fF
C13145 col_n[29] rowon_n[3] 0.17fF
C13146 col_n[31] rowon_n[4] 0.17fF
C13147 VDD col[16] 9.44fF
C13148 a_31078_8154# col_n[28] 0.34fF
C13149 a_20034_4138# vcm 0.89fF
C13150 a_31078_4138# rowoff_n[2] 1.25fF
C13151 a_10998_3134# rowon_n[1] 0.45fF
C13152 a_2275_17214# a_10298_17230# 0.15fF
C13153 a_2475_17214# a_12914_17190# 0.41fF
C13154 a_11302_12210# col_n[8] 0.11fF
C13155 a_2275_5166# a_25054_5142# 0.71fF
C13156 a_29070_13174# VDD 1.75fF
C13157 a_2275_18218# a_20338_18234# 0.15fF
C13158 m2_6752_946# m2_7180_1374# 0.19fF
C13159 a_25054_10162# a_26058_10162# 0.86fF
C13160 a_2874_14178# a_2966_14178# 0.45fF
C13161 a_35094_8154# vcm 0.15fF
C13162 a_22042_12170# row_n[10] 0.43fF
C13163 a_9902_2130# a_9994_2130# 0.45fF
C13164 a_2475_2154# a_17934_2130# 0.41fF
C13165 a_2275_2154# a_15318_2170# 0.15fF
C13166 m2_34864_18014# m3_34996_18146# 4.48fF
C13167 a_21950_16186# rowon_n[14] 0.14fF
C13168 a_2475_7174# col[3] 0.22fF
C13169 a_4974_10162# col[2] 0.38fF
C13170 a_9994_16186# VDD 3.71fF
C13171 a_32082_2130# row_n[0] 0.43fF
C13172 a_16018_12170# a_16018_11166# 0.84fF
C13173 a_31990_6146# rowon_n[4] 0.14fF
C13174 a_25358_2170# vcm 0.24fF
C13175 row_n[12] rowoff_n[12] 0.64fF
C13176 a_2275_16210# a_18938_16186# 0.17fF
C13177 a_2275_13198# col_n[10] 0.17fF
C13178 a_20034_6146# col_n[17] 0.34fF
C13179 a_16018_11166# vcm 0.89fF
C13180 m2_27836_946# col_n[25] 0.51fF
C13181 a_2275_2154# col_n[15] 0.17fF
C13182 a_12914_1126# VDD 0.90fF
C13183 a_2475_4162# a_32994_4138# 0.41fF
C13184 a_2275_4162# a_30378_4178# 0.15fF
C13185 a_35398_11206# VDD 0.12fF
C13186 a_8990_10162# rowon_n[8] 0.45fF
C13187 a_2275_10186# col[0] 0.16fF
C13188 a_2475_13198# a_10998_13174# 0.68fF
C13189 a_5978_13174# a_6982_13174# 0.86fF
C13190 a_32994_10162# rowoff_n[8] 0.40fF
C13191 a_6282_5182# vcm 0.24fF
C13192 a_2475_5166# m2_1732_4962# 0.16fF
C13193 a_2275_1150# a_23958_1126# 0.17fF
C13194 a_31078_15182# vcm 0.89fF
C13195 a_27974_5142# VDD 0.29fF
C13196 a_24962_6146# a_25054_6146# 0.45fF
C13197 a_2475_9182# col[20] 0.22fF
C13198 a_1957_10186# a_2161_10186# 0.11fF
C13199 a_2475_10186# a_2275_10186# 2.96fF
C13200 col_n[23] rowoff_n[13] 0.17fF
C13201 a_31078_16186# a_31078_15182# 0.84fF
C13202 a_2475_15206# a_26058_15182# 0.68fF
C13203 a_21342_9198# vcm 0.24fF
C13204 col[26] rowoff_n[9] 0.17fF
C13205 col[25] rowoff_n[8] 0.18fF
C13206 col[24] rowoff_n[7] 0.19fF
C13207 col[23] rowoff_n[6] 0.19fF
C13208 col[22] rowoff_n[5] 0.20fF
C13209 col[21] rowoff_n[4] 0.21fF
C13210 col[20] rowoff_n[3] 0.21fF
C13211 col[19] rowoff_n[2] 0.22fF
C13212 col[18] rowoff_n[1] 0.23fF
C13213 col[17] rowoff_n[0] 0.23fF
C13214 a_2275_15206# col_n[27] 0.17fF
C13215 a_8990_4138# col_n[6] 0.34fF
C13216 a_34090_4138# ctop 4.80fF
C13217 a_12002_18194# vcm 0.15fF
C13218 a_8898_8154# VDD 0.29fF
C13219 a_30074_9158# row_n[7] 0.43fF
C13220 a_19030_16186# col_n[16] 0.34fF
C13221 a_30074_16186# m2_30272_16434# 0.19fF
C13222 a_29982_13174# rowon_n[11] 0.14fF
C13223 a_2275_12194# a_17022_12170# 0.71fF
C13224 a_2275_12194# col[17] 0.17fF
C13225 a_14922_3134# vcm 0.18fF
C13226 a_21038_17190# a_22042_17190# 0.86fF
C13227 a_2275_1150# col[22] 0.17fF
C13228 m2_31852_18014# m2_32856_18014# 0.86fF
C13229 a_3878_12170# vcm 0.18fF
C13230 a_15014_7150# ctop 4.91fF
C13231 a_23958_12170# VDD 0.29fF
C13232 m3_3872_18146# m3_4876_18146# 0.21fF
C13233 a_29070_3134# col[26] 0.38fF
C13234 a_6982_17190# rowon_n[15] 0.45fF
C13235 a_2275_9182# a_7286_9198# 0.15fF
C13236 a_2475_9182# a_9902_9158# 0.41fF
C13237 a_5886_9158# a_5978_9158# 0.45fF
C13238 col_n[7] rowoff_n[14] 0.29fF
C13239 m2_1732_6970# vcm 1.11fF
C13240 a_2275_14202# a_32082_14178# 0.71fF
C13241 col[10] rowoff_n[10] 0.28fF
C13242 a_29982_7150# vcm 0.18fF
C13243 a_17022_7150# rowon_n[5] 0.45fF
C13244 a_24050_14178# rowoff_n[12] 1.59fF
C13245 a_17326_16226# vcm 0.24fF
C13246 m2_34864_15002# m3_34996_15134# 4.42fF
C13247 a_2275_18218# col_n[29] 0.17fF
C13248 a_21038_14178# m2_21236_14426# 0.19fF
C13249 a_30074_11166# ctop 4.91fF
C13250 a_24354_3174# col_n[21] 0.11fF
C13251 a_4882_15182# VDD 0.29fF
C13252 a_7986_14178# col_n[5] 0.34fF
C13253 a_2275_11190# a_22346_11206# 0.15fF
C13254 a_2475_11190# a_24962_11166# 0.41fF
C13255 a_18026_2130# m2_18224_2378# 0.19fF
C13256 m2_34864_13998# m2_35292_14426# 0.19fF
C13257 a_10906_10162# vcm 0.18fF
C13258 a_28066_16186# row_n[14] 0.43fF
C13259 a_31078_4138# a_32082_4138# 0.86fF
C13260 VDD col[27] 6.75fF
C13261 vcm col[24] 6.66fF
C13262 col_n[31] sw_n 0.53fF
C13263 col_n[12] col[12] 0.50fF
C13264 a_2275_8178# a_15926_8154# 0.17fF
C13265 a_10998_14178# ctop 4.91fF
C13266 a_2275_11190# col_n[4] 0.17fF
C13267 a_20946_13174# a_21038_13174# 0.45fF
C13268 a_18026_1126# col[15] 0.53fF
C13269 ctop rowoff_n[11] 0.28fF
C13270 a_28066_13174# col[25] 0.38fF
C13271 a_1957_4162# vcm 0.16fF
C13272 a_25966_14178# vcm 0.18fF
C13273 a_22042_4138# VDD 2.47fF
C13274 a_2475_5166# a_7986_5142# 0.68fF
C13275 a_22042_6146# a_22042_5142# 0.84fF
C13276 a_12002_12170# m2_12200_12418# 0.19fF
C13277 a_2275_8178# ctop 0.14fF
C13278 a_2275_18218# a_3970_18194# 0.14fF
C13279 a_2275_10186# a_30986_10162# 0.17fF
C13280 a_4974_9158# rowoff_n[7] 2.52fF
C13281 a_13310_1166# col_n[10] 0.11fF
C13282 a_15014_14178# rowon_n[12] 0.45fF
C13283 a_23350_13214# col_n[20] 0.11fF
C13284 a_12002_15182# rowoff_n[13] 2.18fF
C13285 a_2475_7174# col[14] 0.22fF
C13286 a_31078_8154# m2_31276_8402# 0.19fF
C13287 a_25054_4138# rowon_n[2] 0.45fF
C13288 a_6890_17190# vcm 0.18fF
C13289 a_3878_16186# rowon_n[14] 0.14fF
C13290 a_2874_7150# VDD 0.29fF
C13291 a_14010_7150# rowoff_n[5] 2.08fF
C13292 a_2475_7174# a_23046_7150# 0.68fF
C13293 a_12002_7150# a_13006_7150# 0.86fF
C13294 a_2275_13198# col_n[21] 0.17fF
C13295 a_8990_2130# vcm 0.89fF
C13296 a_2275_2154# col_n[26] 0.17fF
C13297 a_23046_5142# rowoff_n[3] 1.64fF
C13298 a_17022_11166# col[14] 0.38fF
C13299 a_2275_4162# a_14010_4138# 0.71fF
C13300 a_18026_11166# VDD 2.89fF
C13301 a_2275_10186# col[11] 0.17fF
C13302 a_32082_7150# col_n[29] 0.34fF
C13303 a_32082_3134# rowoff_n[1] 1.20fF
C13304 a_24050_6146# vcm 0.89fF
C13305 a_12306_11206# col_n[9] 0.11fF
C13306 a_2475_9182# col[31] 0.22fF
C13307 a_2275_1150# a_4274_1166# 0.19fF
C13308 a_22042_6146# m2_22240_6394# 0.19fF
C13309 a_2475_1150# a_6890_1126# 0.41fF
C13310 m2_34864_11990# m3_34996_12122# 4.46fF
C13311 a_2275_6170# a_29070_6146# 0.71fF
C13312 a_33086_15182# VDD 1.34fF
C13313 a_27062_11166# a_28066_11166# 0.86fF
C13314 col[28] rowoff_n[0] 0.16fF
C13315 col[29] rowoff_n[1] 0.15fF
C13316 col[30] rowoff_n[2] 0.15fF
C13317 col[31] rowoff_n[3] 0.14fF
C13318 sample_n rowoff_n[4] 0.55fF
C13319 m2_30848_18014# vcm 0.71fF
C13320 a_2275_15206# a_7894_15182# 0.17fF
C13321 a_23046_11166# rowon_n[9] 0.45fF
C13322 a_4974_9158# vcm 0.89fF
C13323 a_2475_3158# a_21950_3134# 0.41fF
C13324 a_2275_3158# a_19334_3174# 0.15fF
C13325 a_11910_3134# a_12002_3134# 0.45fF
C13326 a_32082_2130# m2_31852_946# 0.84fF
C13327 a_2475_1150# m2_23820_946# 0.62fF
C13328 a_5978_9158# col[3] 0.38fF
C13329 m3_25960_1078# ctop 0.21fF
C13330 a_2275_12194# col[28] 0.17fF
C13331 a_18026_13174# a_18026_12170# 0.84fF
C13332 a_21038_5142# col_n[18] 0.34fF
C13333 a_29374_4178# vcm 0.24fF
C13334 a_24962_11166# rowoff_n[9] 0.49fF
C13335 a_2275_17214# a_22954_17190# 0.17fF
C13336 a_31078_17190# col_n[28] 0.34fF
C13337 a_13006_4138# m2_13204_4386# 0.19fF
C13338 a_20034_13174# vcm 0.89fF
C13339 a_16930_3134# VDD 0.29fF
C13340 col_n[18] rowoff_n[14] 0.21fF
C13341 a_2275_5166# a_35398_5182# 0.15fF
C13342 a_10906_5142# rowon_n[3] 0.14fF
C13343 a_2275_18218# a_32994_18194# 0.17fF
C13344 col[21] rowoff_n[10] 0.21fF
C13345 a_33998_9158# rowoff_n[7] 0.39fF
C13346 a_7986_14178# a_8990_14178# 0.86fF
C13347 a_2475_14202# a_15014_14178# 0.68fF
C13348 a_10298_7190# vcm 0.24fF
C13349 a_2275_2154# a_27974_2130# 0.17fF
C13350 a_23046_2130# ctop 4.93fF
C13351 a_35094_17190# vcm 0.15fF
C13352 a_31990_7150# VDD 0.29fF
C13353 a_26970_7150# a_27062_7150# 0.45fF
C13354 a_2475_16210# col[3] 0.22fF
C13355 a_2275_11190# a_5978_11166# 0.71fF
C13356 a_2475_5166# col[8] 0.22fF
C13357 a_2475_16210# a_30074_16186# 0.68fF
C13358 a_33086_17190# a_33086_16186# 0.84fF
C13359 a_25358_11206# vcm 0.24fF
C13360 a_9994_3134# col_n[7] 0.34fF
C13361 col_n[2] rowoff_n[15] 0.32fF
C13362 row_n[11] ctop 0.28fF
C13363 col_n[17] col[18] 6.24fF
C13364 a_23446_1488# VDD 0.14fF
C13365 a_20034_15182# col_n[17] 0.34fF
C13366 a_31078_8154# rowon_n[6] 0.45fF
C13367 a_3970_5142# ctop 4.91fF
C13368 a_2275_11190# col_n[15] 0.17fF
C13369 a_12914_10162# VDD 0.29fF
C13370 col[5] rowoff_n[11] 0.31fF
C13371 a_2275_13198# a_21038_13174# 0.71fF
C13372 a_18938_5142# vcm 0.18fF
C13373 a_12914_12170# rowoff_n[10] 0.63fF
C13374 a_2275_18218# m2_14784_18014# 0.51fF
C13375 m2_8760_18014# col_n[6] 0.33fF
C13376 a_8990_8154# row_n[6] 0.43fF
C13377 a_18026_1126# a_19030_1126# 0.86fF
C13378 a_2275_8178# col[5] 0.17fF
C13379 a_6282_14218# vcm 0.24fF
C13380 m2_34864_8978# m3_34996_9110# 4.42fF
C13381 a_8898_12170# rowon_n[10] 0.14fF
C13382 a_34394_4178# col_n[31] 0.11fF
C13383 a_19030_9158# ctop 4.91fF
C13384 a_30074_2130# col[27] 0.38fF
C13385 a_27974_14178# VDD 0.29fF
C13386 a_2275_10186# a_11302_10202# 0.15fF
C13387 a_2475_10186# a_13918_10162# 0.41fF
C13388 a_7894_10162# a_7986_10162# 0.45fF
C13389 a_4882_2130# rowoff_n[0] 0.72fF
C13390 a_18938_2130# rowon_n[0] 0.14fF
C13391 a_2475_7174# col[25] 0.22fF
C13392 a_33998_9158# vcm 0.18fF
C13393 a_28978_16186# rowoff_n[14] 0.44fF
C13394 a_8990_3134# a_8990_2130# 0.84fF
C13395 a_21342_18234# vcm 0.25fF
C13396 a_25358_2170# col_n[22] 0.11fF
C13397 a_2275_7174# a_4882_7150# 0.17fF
C13398 a_8990_13174# col_n[6] 0.34fF
C13399 a_2966_7150# a_3970_7150# 0.86fF
C13400 a_34090_13174# ctop 4.80fF
C13401 a_8898_17190# VDD 0.29fF
C13402 a_2275_12194# a_26362_12210# 0.15fF
C13403 a_2475_12194# a_28978_12170# 0.41fF
C13404 a_29070_15182# rowon_n[13] 0.45fF
C13405 a_14922_12170# vcm 0.18fF
C13406 a_2275_10186# col[22] 0.17fF
C13407 a_10998_2130# VDD 3.61fF
C13408 a_33086_5142# a_34090_5142# 0.86fF
C13409 a_2275_9182# a_19942_9158# 0.17fF
C13410 a_14922_18194# m2_14784_18014# 0.34fF
C13411 a_15014_16186# ctop 4.91fF
C13412 a_22954_14178# a_23046_14178# 0.45fF
C13413 a_29070_12170# col[26] 0.38fF
C13414 a_6982_15182# row_n[13] 0.43fF
C13415 a_2275_18218# a_2874_18194# 0.17fF
C13416 a_29982_16186# vcm 0.18fF
C13417 a_26058_6146# VDD 2.06fF
C13418 a_17022_5142# row_n[3] 0.43fF
C13419 a_24050_7150# a_24050_6146# 0.84fF
C13420 a_2475_6170# a_12002_6146# 0.68fF
C13421 a_16930_9158# rowon_n[7] 0.14fF
C13422 a_5978_8154# rowoff_n[6] 2.47fF
C13423 a_2275_11190# a_35002_11166# 0.17fF
C13424 a_24354_12210# col_n[21] 0.11fF
C13425 a_32082_1126# vcm 0.15fF
C13426 a_16930_17190# rowoff_n[15] 0.58fF
C13427 m2_34864_18014# VDD 2.39fF
C13428 a_15014_6146# rowoff_n[4] 2.03fF
C13429 a_2475_3158# a_3878_3134# 0.41fF
C13430 a_2275_3158# a_2874_3134# 0.17fF
C13431 a_2475_3158# col[2] 0.22fF
C13432 m3_21944_18146# ctop 0.21fF
C13433 a_6982_9158# VDD 4.02fF
C13434 a_2475_8178# a_27062_8154# 0.68fF
C13435 a_14010_8154# a_15014_8154# 0.86fF
C13436 a_13006_4138# vcm 0.89fF
C13437 a_3970_3134# rowon_n[1] 0.45fF
C13438 a_24050_4138# rowoff_n[2] 1.59fF
C13439 a_2475_17214# a_5886_17190# 0.41fF
C13440 a_2275_17214# a_3270_17230# 0.15fF
C13441 a_18026_10162# col[15] 0.38fF
C13442 a_2275_9182# col_n[9] 0.17fF
C13443 col_n[29] rowoff_n[14] 0.13fF
C13444 a_32994_1126# a_33086_1126# 0.11fF
C13445 a_1957_13198# vcm 0.16fF
C13446 m2_34864_5966# m3_34996_6098# 4.45fF
C13447 a_2275_5166# a_18026_5142# 0.71fF
C13448 sample_n rowoff_n[10] 0.55fF
C13449 a_33086_6146# col_n[30] 0.34fF
C13450 a_22042_13174# VDD 2.47fF
C13451 a_2275_18218# a_13310_18234# 0.15fF
C13452 a_4974_10162# a_4974_9158# 0.84fF
C13453 a_2275_17214# ctop 0.14fF
C13454 a_33086_2130# rowoff_n[0] 1.15fF
C13455 a_13310_10202# col_n[10] 0.11fF
C13456 a_28066_8154# vcm 0.89fF
C13457 a_15014_12170# row_n[10] 0.43fF
C13458 a_2475_2154# a_10906_2130# 0.41fF
C13459 a_2275_2154# a_8290_2170# 0.15fF
C13460 a_14922_16186# rowon_n[14] 0.14fF
C13461 a_2475_16210# col[14] 0.22fF
C13462 a_2475_5166# col[19] 0.22fF
C13463 a_2275_7174# a_33086_7150# 0.71fF
C13464 a_27062_15182# m2_27260_15430# 0.19fF
C13465 a_2874_16186# VDD 0.29fF
C13466 a_25054_2130# row_n[0] 0.43fF
C13467 a_29070_12170# a_30074_12170# 0.86fF
C13468 a_24962_6146# rowon_n[4] 0.14fF
C13469 a_18330_2170# vcm 0.24fF
C13470 col_n[23] col[23] 0.50fF
C13471 rowon_n[5] ctop 0.37fF
C13472 col_n[13] rowoff_n[15] 0.24fF
C13473 a_2275_16210# a_11910_16186# 0.17fF
C13474 a_2275_11190# col_n[26] 0.17fF
C13475 a_8990_11166# vcm 0.89fF
C13476 a_5886_1126# VDD 0.98fF
C13477 a_6982_8154# col[4] 0.38fF
C13478 col[16] rowoff_n[11] 0.24fF
C13479 a_2275_4162# a_23350_4178# 0.15fF
C13480 a_2475_4162# a_25966_4138# 0.41fF
C13481 a_13918_4138# a_14010_4138# 0.45fF
C13482 a_33998_18194# m2_33860_18014# 0.34fF
C13483 a_10998_17190# m2_10768_18014# 0.84fF
C13484 a_22042_4138# col_n[19] 0.34fF
C13485 a_2475_10186# rowon_n[8] 0.40fF
C13486 a_2475_13198# a_3970_13174# 0.68fF
C13487 a_2275_13198# a_2966_13174# 0.67fF
C13488 a_20034_14178# a_20034_13174# 0.84fF
C13489 a_25966_10162# rowoff_n[8] 0.48fF
C13490 a_2275_8178# col[16] 0.17fF
C13491 a_32082_16186# col_n[29] 0.34fF
C13492 a_33390_6186# vcm 0.24fF
C13493 a_29070_13174# rowoff_n[11] 1.35fF
C13494 a_2275_1150# a_16930_1126# 0.17fF
C13495 a_24050_15182# vcm 0.89fF
C13496 a_20946_5142# VDD 0.29fF
C13497 m2_21812_946# VDD 4.45fF
C13498 a_18026_13174# m2_18224_13422# 0.19fF
C13499 a_35002_8154# rowoff_n[6] 0.38fF
C13500 a_2475_15206# a_19030_15182# 0.68fF
C13501 a_9994_15182# a_10998_15182# 0.86fF
C13502 m2_11772_946# col_n[9] 0.45fF
C13503 a_14314_9198# vcm 0.24fF
C13504 col[0] rowoff_n[12] 0.34fF
C13505 a_2275_3158# a_31990_3134# 0.17fF
C13506 a_27062_4138# ctop 4.91fF
C13507 a_4974_18194# vcm 0.15fF
C13508 a_23046_9158# row_n[7] 0.43fF
C13509 a_28978_8154# a_29070_8154# 0.45fF
C13510 a_22954_13174# rowon_n[11] 0.14fF
C13511 a_2275_12194# a_9994_12170# 0.71fF
C13512 m2_34864_16006# row_n[14] 0.38fF
C13513 a_7894_3134# vcm 0.18fF
C13514 a_32994_3134# rowon_n[1] 0.14fF
C13515 a_10998_2130# col_n[8] 0.34fF
C13516 a_2475_17214# a_34090_17190# 0.68fF
C13517 a_21038_14178# col_n[18] 0.34fF
C13518 m2_24824_18014# m2_25828_18014# 0.86fF
C13519 a_29374_13214# vcm 0.24fF
C13520 m2_34864_2954# m3_34996_3086# 4.47fF
C13521 a_8990_11166# m2_9188_11414# 0.19fF
C13522 a_7986_7150# ctop 4.91fF
C13523 a_16930_12170# VDD 0.29fF
C13524 m2_29844_946# m2_30272_1374# 0.19fF
C13525 a_2275_7174# col_n[3] 0.17fF
C13526 a_2275_14202# a_25054_14178# 0.71fF
C13527 a_22954_7150# vcm 0.18fF
C13528 a_9994_7150# rowon_n[5] 0.45fF
C13529 a_17022_14178# rowoff_n[12] 1.94fF
C13530 a_28066_7150# m2_28264_7398# 0.19fF
C13531 a_20034_2130# a_21038_2130# 0.86fF
C13532 a_10298_16226# vcm 0.24fF
C13533 a_23046_11166# ctop 4.91fF
C13534 a_31990_16186# VDD 0.29fF
C13535 a_9902_11166# a_9994_11166# 0.45fF
C13536 a_2275_11190# a_15318_11206# 0.15fF
C13537 a_2475_11190# a_17934_11166# 0.41fF
C13538 a_2475_14202# col[8] 0.22fF
C13539 a_2475_3158# col[13] 0.22fF
C13540 a_26362_1166# col_n[23] 0.11fF
C13541 a_21038_16186# row_n[14] 0.43fF
C13542 a_10998_4138# a_10998_3134# 0.84fF
C13543 a_9994_12170# col_n[7] 0.34fF
C13544 a_2275_8178# a_8898_8154# 0.17fF
C13545 a_30074_17190# m2_29844_18014# 0.84fF
C13546 a_3970_14178# ctop 4.91fF
C13547 a_31078_6146# row_n[4] 0.43fF
C13548 a_2275_9182# col_n[20] 0.17fF
C13549 a_2475_13198# a_32994_13174# 0.41fF
C13550 a_2275_13198# a_30378_13214# 0.15fF
C13551 a_30986_10162# rowon_n[8] 0.14fF
C13552 m2_34864_3958# m2_34864_2954# 0.84fF
C13553 a_19030_5142# m2_19228_5390# 0.19fF
C13554 a_18938_14178# vcm 0.18fF
C13555 m2_34864_7974# rowoff_n[6] 1.01fF
C13556 a_15014_4138# VDD 3.20fF
C13557 a_2275_17214# col[5] 0.17fF
C13558 a_2275_6170# col[10] 0.17fF
C13559 a_34394_13214# col_n[31] 0.11fF
C13560 a_2275_10186# a_23958_10162# 0.17fF
C13561 a_30074_11166# col[27] 0.38fF
C13562 a_7986_14178# rowon_n[12] 0.45fF
C13563 a_24962_15182# a_25054_15182# 0.45fF
C13564 a_2475_16210# col[25] 0.22fF
C13565 m2_23820_18014# col[21] 0.37fF
C13566 a_4974_15182# rowoff_n[13] 2.52fF
C13567 a_2475_5166# col[30] 0.22fF
C13568 a_18026_4138# rowon_n[2] 0.45fF
C13569 a_33998_18194# vcm 0.18fF
C13570 m2_1732_18014# m3_1864_18146# 4.44fF
C13571 a_30074_8154# VDD 1.65fF
C13572 a_6982_7150# rowoff_n[5] 2.42fF
C13573 a_26058_8154# a_26058_7150# 0.84fF
C13574 a_2475_7174# a_16018_7150# 0.68fF
C13575 a_25358_11206# col_n[22] 0.11fF
C13576 row_n[0] ctop 0.27fF
C13577 col_n[24] rowoff_n[15] 0.16fF
C13578 sw sw_n 0.22fF
C13579 col_n[28] col[29] 6.15fF
C13580 a_2475_2154# vcm 1.32fF
C13581 col[27] rowoff_n[11] 0.17fF
C13582 a_9994_3134# m2_10192_3382# 0.19fF
C13583 a_16018_5142# rowoff_n[3] 1.98fF
C13584 a_2275_4162# a_6982_4138# 0.71fF
C13585 a_29070_13174# row_n[11] 0.43fF
C13586 a_10998_11166# VDD 3.61fF
C13587 a_28978_17190# rowon_n[15] 0.14fF
C13588 a_16018_9158# a_17022_9158# 0.86fF
C13589 a_2475_9182# a_31078_9158# 0.68fF
C13590 a_2275_8178# col[27] 0.17fF
C13591 a_25054_3134# rowoff_n[1] 1.54fF
C13592 a_19030_9158# col[16] 0.38fF
C13593 a_17022_6146# vcm 0.89fF
C13594 a_5886_18194# a_5978_18194# 0.11fF
C13595 a_35002_2130# a_35094_2130# 0.11fF
C13596 a_2275_5166# VDD 3.18fF
C13597 a_34090_5142# col_n[31] 0.34fF
C13598 a_2275_6170# a_22042_6146# 0.71fF
C13599 a_26058_15182# VDD 2.06fF
C13600 a_6982_11166# a_6982_10162# 0.84fF
C13601 a_14314_9198# col_n[11] 0.11fF
C13602 col[11] rowoff_n[12] 0.27fF
C13603 m2_16792_18014# vcm 0.71fF
C13604 a_16018_11166# rowon_n[9] 0.45fF
C13605 a_32082_10162# vcm 0.89fF
C13606 a_2275_3158# a_12306_3174# 0.15fF
C13607 a_2475_3158# a_14922_3134# 0.41fF
C13608 a_3970_1126# m2_4168_1374# 0.19fF
C13609 a_2275_1150# m2_6752_946# 0.51fF
C13610 m3_34996_3086# ctop 0.22fF
C13611 a_2475_12194# col[2] 0.22fF
C13612 a_2475_1150# col[7] 0.22fF
C13613 a_31078_13174# a_32082_13174# 0.86fF
C13614 a_22346_4178# vcm 0.24fF
C13615 a_17934_11166# rowoff_n[9] 0.57fF
C13616 a_2275_17214# a_15926_17190# 0.17fF
C13617 a_7986_7150# col[5] 0.38fF
C13618 a_13006_13174# vcm 0.89fF
C13619 a_9902_3134# VDD 0.29fF
C13620 a_2275_5166# a_27366_5182# 0.15fF
C13621 a_2475_5166# a_29982_5142# 0.41fF
C13622 a_15926_5142# a_16018_5142# 0.45fF
C13623 a_2275_7174# col_n[14] 0.17fF
C13624 a_2275_18218# a_25966_18194# 0.17fF
C13625 a_23046_3134# col_n[20] 0.34fF
C13626 a_26970_9158# rowoff_n[7] 0.47fF
C13627 a_33086_15182# col_n[30] 0.34fF
C13628 a_2475_14202# a_7986_14178# 0.68fF
C13629 a_22042_15182# a_22042_14178# 0.84fF
C13630 a_3270_7190# vcm 0.24fF
C13631 a_33998_15182# rowoff_n[13] 0.39fF
C13632 a_2275_4162# col[4] 0.17fF
C13633 a_2275_2154# a_20946_2130# 0.17fF
C13634 a_16018_2130# ctop 4.93fF
C13635 a_28066_17190# vcm 0.89fF
C13636 a_24962_7150# VDD 0.29fF
C13637 a_2475_14202# col[19] 0.22fF
C13638 a_2475_3158# col[24] 0.22fF
C13639 a_30986_2130# vcm 0.18fF
C13640 a_2475_16210# a_23046_16186# 0.68fF
C13641 a_12002_16186# a_13006_16186# 0.86fF
C13642 m2_1732_9982# sample 0.31fF
C13643 a_2475_18218# col[10] 0.22fF
C13644 a_18330_11206# vcm 0.24fF
C13645 a_16418_1488# VDD 0.15fF
C13646 a_2966_16186# row_n[14] 0.41fF
C13647 a_24050_8154# rowon_n[6] 0.45fF
C13648 a_2275_4162# a_34394_4178# 0.15fF
C13649 a_31078_6146# ctop 4.91fF
C13650 a_5886_10162# VDD 0.29fF
C13651 a_6982_17190# col[4] 0.38fF
C13652 a_2275_9182# col_n[31] 0.17fF
C13653 a_30986_9158# a_31078_9158# 0.45fF
C13654 a_2275_13198# a_14010_13174# 0.71fF
C13655 a_22042_13174# col_n[19] 0.34fF
C13656 a_11910_5142# vcm 0.18fF
C13657 a_5886_12170# rowoff_n[10] 0.70fF
C13658 a_2275_17214# col[16] 0.17fF
C13659 a_2475_8178# row_n[6] 0.48fF
C13660 a_33390_15222# vcm 0.24fF
C13661 a_2275_6170# col[21] 0.17fF
C13662 a_2275_18218# col[1] 0.17fF
C13663 a_12002_9158# ctop 4.91fF
C13664 a_20946_14178# VDD 0.29fF
C13665 a_2275_10186# a_4274_10202# 0.15fF
C13666 a_2475_10186# a_6890_10162# 0.41fF
C13667 a_11910_2130# rowon_n[0] 0.14fF
C13668 a_2275_15206# a_29070_15182# 0.71fF
C13669 a_26970_9158# vcm 0.18fF
C13670 a_21950_16186# rowoff_n[14] 0.52fF
C13671 a_22042_3134# a_23046_3134# 0.86fF
C13672 a_14314_18234# vcm 0.25fF
C13673 a_23958_1126# m2_23820_946# 0.31fF
C13674 en_C0_n col[1] 0.14fF
C13675 ctop col[2] 0.13fF
C13676 rowon_n[13] sample_n 0.15fF
C13677 a_33086_16186# m2_33284_16434# 0.19fF
C13678 a_27062_13174# ctop 4.91fF
C13679 a_11910_12170# a_12002_12170# 0.45fF
C13680 a_2275_12194# a_19334_12210# 0.15fF
C13681 a_2475_12194# a_21950_12170# 0.41fF
C13682 a_22042_15182# rowon_n[13] 0.45fF
C13683 m2_1732_17010# m2_2160_17438# 0.19fF
C13684 a_7894_12170# vcm 0.18fF
C13685 a_10998_11166# col_n[8] 0.34fF
C13686 a_3970_2130# VDD 4.33fF
C13687 a_13006_5142# a_13006_4138# 0.84fF
C13688 a_32082_5142# rowon_n[3] 0.45fF
C13689 m2_7756_946# m3_7888_1078# 4.41fF
C13690 a_2275_9182# a_12914_9158# 0.17fF
C13691 a_7986_16186# ctop 4.91fF
C13692 a_2475_18218# m2_26832_18014# 0.62fF
C13693 a_2275_14202# a_35398_14218# 0.15fF
C13694 m2_21812_946# col_n[19] 0.45fF
C13695 a_2275_16210# col_n[3] 0.17fF
C13696 a_2275_5166# col_n[8] 0.17fF
C13697 a_22954_16186# vcm 0.18fF
C13698 a_19030_6146# VDD 2.78fF
C13699 a_9994_5142# row_n[3] 0.43fF
C13700 a_2475_6170# a_4974_6146# 0.68fF
C13701 a_24050_14178# m2_24248_14426# 0.19fF
C13702 a_31078_10162# col[28] 0.38fF
C13703 a_9902_9158# rowon_n[7] 0.14fF
C13704 col[22] rowoff_n[12] 0.20fF
C13705 a_2275_11190# a_27974_11166# 0.17fF
C13706 a_25054_1126# vcm 0.15fF
C13707 a_26970_16186# a_27062_16186# 0.45fF
C13708 a_9902_17190# rowoff_n[15] 0.66fF
C13709 m2_20808_18014# VDD 3.37fF
C13710 a_2475_9182# m2_34864_8978# 0.56fF
C13711 a_7986_6146# rowoff_n[4] 2.38fF
C13712 a_2475_12194# col[13] 0.22fF
C13713 a_15014_2130# m2_14784_946# 0.84fF
C13714 a_26362_10202# col_n[23] 0.11fF
C13715 a_34090_10162# VDD 1.23fF
C13716 a_2475_1150# col[18] 0.21fF
C13717 a_28066_9158# a_28066_8154# 0.84fF
C13718 a_2475_8178# a_20034_8154# 0.68fF
C13719 a_5978_4138# vcm 0.89fF
C13720 a_34090_12170# rowoff_n[10] 1.10fF
C13721 a_17022_4138# rowoff_n[2] 1.94fF
C13722 a_2275_7174# col_n[25] 0.17fF
C13723 a_30074_12170# rowon_n[10] 0.45fF
C13724 a_15014_12170# m2_15212_12418# 0.19fF
C13725 a_2275_5166# a_10998_5142# 0.71fF
C13726 col[6] rowoff_n[13] 0.31fF
C13727 a_15014_13174# VDD 3.20fF
C13728 a_2275_18218# a_6282_18234# 0.15fF
C13729 a_18026_10162# a_19030_10162# 0.86fF
C13730 a_26058_2130# rowoff_n[0] 1.50fF
C13731 a_2275_15206# col[10] 0.17fF
C13732 a_20034_8154# col[17] 0.38fF
C13733 a_2275_4162# col[15] 0.17fF
C13734 a_21038_8154# vcm 0.89fF
C13735 a_7986_12170# row_n[10] 0.43fF
C13736 a_34090_8154# m2_34288_8402# 0.19fF
C13737 a_7894_16186# rowon_n[14] 0.14fF
C13738 a_2475_14202# col[30] 0.22fF
C13739 a_2275_7174# a_26058_7150# 0.71fF
C13740 m2_2736_1950# rowoff_n[0] 2.51fF
C13741 a_30074_17190# VDD 1.65fF
C13742 a_18026_2130# row_n[0] 0.43fF
C13743 a_15318_8194# col_n[12] 0.11fF
C13744 a_8990_12170# a_8990_11166# 0.84fF
C13745 a_17934_6146# rowon_n[4] 0.14fF
C13746 a_2475_18218# col[21] 0.22fF
C13747 a_11302_2170# vcm 0.24fF
C13748 a_2275_16210# a_4882_16186# 0.17fF
C13749 a_2966_16186# a_3970_16186# 0.86fF
C13750 a_2475_11190# vcm 1.32fF
C13751 a_32994_2130# VDD 0.29fF
C13752 a_5978_10162# m2_6176_10410# 0.19fF
C13753 a_2275_4162# a_16322_4178# 0.15fF
C13754 a_2475_4162# a_18938_4138# 0.41fF
C13755 a_33086_14178# a_34090_14178# 0.86fF
C13756 a_18938_10162# rowoff_n[8] 0.56fF
C13757 a_2275_17214# col[27] 0.17fF
C13758 a_8990_6146# col[6] 0.38fF
C13759 a_26362_6186# vcm 0.24fF
C13760 a_22042_13174# rowoff_n[11] 1.69fF
C13761 a_2275_18218# col[12] 0.17fF
C13762 a_25054_6146# m2_25252_6394# 0.19fF
C13763 a_2275_1150# a_9902_1126# 0.17fF
C13764 a_17022_15182# vcm 0.89fF
C13765 a_13918_5142# VDD 0.29fF
C13766 a_17934_6146# a_18026_6146# 0.45fF
C13767 a_2275_6170# a_31382_6186# 0.15fF
C13768 a_2475_6170# a_33998_6146# 0.41fF
C13769 a_24050_2130# col_n[21] 0.34fF
C13770 a_2275_14202# VDD 3.18fF
C13771 a_27974_8154# rowoff_n[6] 0.46fF
C13772 a_34090_14178# col_n[31] 0.34fF
C13773 a_2275_3158# col_n[2] 0.17fF
C13774 a_4274_6186# col_n[1] 0.11fF
C13775 a_24050_16186# a_24050_15182# 0.84fF
C13776 a_2475_15206# a_12002_15182# 0.68fF
C13777 a_14314_18234# col_n[11] 0.11fF
C13778 a_7286_9198# vcm 0.24fF
C13779 row_n[8] sample_n 0.16fF
C13780 a_3878_16186# rowoff_n[14] 0.73fF
C13781 ctop col[13] 0.13fF
C13782 a_2275_3158# a_24962_3134# 0.17fF
C13783 a_20034_4138# ctop 4.91fF
C13784 a_2275_1150# m2_29844_946# 0.51fF
C13785 a_16018_9158# row_n[7] 0.43fF
C13786 a_28978_9158# VDD 0.29fF
C13787 a_15926_13174# rowon_n[11] 0.14fF
C13788 a_2275_12194# a_2874_12170# 0.17fF
C13789 a_2475_12194# a_3878_12170# 0.41fF
C13790 a_35002_4138# vcm 0.18fF
C13791 a_25966_3134# rowon_n[1] 0.14fF
C13792 a_2475_10186# col[7] 0.22fF
C13793 a_2475_17214# a_27062_17190# 0.68fF
C13794 a_14010_17190# a_15014_17190# 0.86fF
C13795 a_16018_4138# m2_16216_4386# 0.19fF
C13796 m2_17796_18014# m2_18800_18014# 0.86fF
C13797 a_22346_13214# vcm 0.24fF
C13798 a_7986_16186# col[5] 0.38fF
C13799 a_9902_12170# VDD 0.29fF
C13800 m2_22816_946# m2_23244_1374# 0.19fF
C13801 a_32994_10162# a_33086_10162# 0.45fF
C13802 a_2275_16210# col_n[14] 0.17fF
C13803 a_2275_5166# col_n[19] 0.17fF
C13804 a_23046_12170# col_n[20] 0.34fF
C13805 a_2275_14202# a_18026_14178# 0.71fF
C13806 a_2874_7150# rowon_n[5] 0.14fF
C13807 a_15926_7150# vcm 0.18fF
C13808 a_9994_14178# rowoff_n[12] 2.28fF
C13809 a_34090_3134# a_34090_2130# 0.84fF
C13810 a_2475_2154# a_32082_2130# 0.68fF
C13811 a_3270_16226# vcm 0.24fF
C13812 a_35494_7512# VDD 0.13fF
C13813 a_2275_13198# col[4] 0.17fF
C13814 a_16018_11166# ctop 4.91fF
C13815 a_2275_2154# col[9] 0.17fF
C13816 a_24962_16186# VDD 0.29fF
C13817 a_2275_11190# a_8290_11206# 0.15fF
C13818 a_2475_11190# a_10906_11166# 0.41fF
C13819 m2_2736_1950# m2_2736_946# 0.84fF
C13820 a_2275_16210# a_33086_16186# 0.71fF
C13821 a_2475_12194# col[24] 0.22fF
C13822 a_30986_11166# vcm 0.18fF
C13823 a_2475_1150# col[29] 0.22fF
C13824 a_14010_16186# row_n[14] 0.43fF
C13825 a_24050_4138# a_25054_4138# 0.86fF
C13826 a_31078_15182# ctop 4.91fF
C13827 a_24050_6146# row_n[4] 0.43fF
C13828 a_23958_10162# rowon_n[8] 0.14fF
C13829 a_13918_13174# a_14010_13174# 0.45fF
C13830 a_2475_13198# a_25966_13174# 0.41fF
C13831 a_2275_13198# a_23350_13214# 0.15fF
C13832 a_12002_10162# col_n[9] 0.34fF
C13833 col[17] rowoff_n[13] 0.23fF
C13834 a_11910_14178# vcm 0.18fF
C13835 a_7986_4138# VDD 3.92fF
C13836 a_15014_6146# a_15014_5142# 0.84fF
C13837 col_n[0] rowoff_n[8] 0.34fF
C13838 vcm rowoff_n[9] 2.43fF
C13839 sample rowoff_n[7] 0.22fF
C13840 VDD rowoff_n[6] 87.22fF
C13841 a_2275_15206# col[21] 0.17fF
C13842 a_2275_4162# col[26] 0.17fF
C13843 a_2275_10186# a_16930_10162# 0.17fF
C13844 a_2966_8154# vcm 0.89fF
C13845 a_10998_4138# rowon_n[2] 0.45fF
C13846 a_26970_18194# vcm 0.18fF
C13847 a_23046_8154# VDD 2.37fF
C13848 a_32082_9158# col[29] 0.38fF
C13849 a_4974_7150# a_5978_7150# 0.86fF
C13850 a_2475_7174# a_8990_7150# 0.68fF
C13851 a_2275_12194# a_31990_12170# 0.17fF
C13852 a_29070_3134# vcm 0.89fF
C13853 a_28978_17190# a_29070_17190# 0.45fF
C13854 col[1] rowoff_n[14] 0.34fF
C13855 a_8990_5142# rowoff_n[3] 2.33fF
C13856 a_27366_9198# col_n[24] 0.11fF
C13857 a_22042_13174# row_n[11] 0.43fF
C13858 a_3970_11166# VDD 4.33fF
C13859 m3_32988_18146# m3_33992_18146# 0.21fF
C13860 a_21950_17190# rowon_n[15] 0.14fF
C13861 a_30074_10162# a_30074_9158# 0.84fF
C13862 a_2475_9182# a_24050_9158# 0.68fF
C13863 a_2475_8178# col[1] 0.22fF
C13864 a_2275_18218# col[23] 0.17fF
C13865 a_32082_3134# row_n[1] 0.43fF
C13866 a_18026_3134# rowoff_n[1] 1.89fF
C13867 a_31990_7150# rowon_n[5] 0.14fF
C13868 a_9994_6146# vcm 0.89fF
C13869 a_2275_14202# col_n[8] 0.17fF
C13870 a_2275_3158# col_n[13] 0.17fF
C13871 a_2275_6170# a_15014_6146# 0.71fF
C13872 a_19030_15182# VDD 2.78fF
C13873 a_21038_7150# col[18] 0.38fF
C13874 a_20034_11166# a_21038_11166# 0.86fF
C13875 VDD col_n[1] 15.69fF
C13876 sample vcm 17.23fF
C13877 ctop col[24] 0.13fF
C13878 m2_2736_18014# vcm 0.71fF
C13879 rowon_n[2] sample_n 0.15fF
C13880 a_3270_3174# col_n[0] 0.11fF
C13881 a_8990_11166# rowon_n[9] 0.45fF
C13882 a_25054_10162# vcm 0.89fF
C13883 a_2275_3158# a_5278_3174# 0.15fF
C13884 a_2475_3158# a_7894_3134# 0.41fF
C13885 a_4882_3134# a_4974_3134# 0.45fF
C13886 m3_34996_17142# ctop 0.22fF
C13887 a_16322_7190# col_n[13] 0.11fF
C13888 a_2275_8178# a_30074_8154# 0.71fF
C13889 a_2475_10186# col[18] 0.22fF
C13890 a_10998_13174# a_10998_12170# 0.84fF
C13891 a_15318_4178# vcm 0.24fF
C13892 a_10906_11166# rowoff_n[9] 0.65fF
C13893 a_2275_17214# a_8898_17190# 0.17fF
C13894 a_2475_4162# m2_1732_3958# 0.16fF
C13895 a_5978_13174# vcm 0.89fF
C13896 a_2161_3158# VDD 0.23fF
C13897 a_2275_16210# col_n[25] 0.17fF
C13898 a_2275_5166# a_20338_5182# 0.15fF
C13899 a_2475_5166# a_22954_5142# 0.41fF
C13900 a_2275_5166# col_n[30] 0.17fF
C13901 a_2275_18218# a_18938_18194# 0.17fF
C13902 a_30074_10162# row_n[8] 0.43fF
C13903 a_19942_9158# rowoff_n[7] 0.55fF
C13904 a_29982_14178# rowon_n[12] 0.14fF
C13905 a_9994_5142# col[7] 0.38fF
C13906 a_20034_17190# col[17] 0.38fF
C13907 a_30378_8194# vcm 0.24fF
C13908 a_26970_15182# rowoff_n[13] 0.47fF
C13909 a_2275_13198# col[15] 0.17fF
C13910 a_2275_2154# a_13918_2130# 0.17fF
C13911 a_8990_2130# ctop 4.93fF
C13912 a_2275_2154# col[20] 0.17fF
C13913 a_21038_17190# vcm 0.89fF
C13914 a_17934_7150# VDD 0.29fF
C13915 a_28978_7150# rowoff_n[5] 0.44fF
C13916 a_19942_7150# a_20034_7150# 0.45fF
C13917 a_30074_15182# m2_30272_15430# 0.19fF
C13918 a_5278_5182# col_n[2] 0.11fF
C13919 a_15318_17230# col_n[12] 0.11fF
C13920 a_23958_2130# vcm 0.18fF
C13921 a_26058_17190# a_26058_16186# 0.84fF
C13922 a_2475_16210# a_16018_16186# 0.68fF
C13923 a_11302_11206# vcm 0.24fF
C13924 a_9390_1488# VDD 0.17fF
C13925 a_17022_8154# rowon_n[6] 0.45fF
C13926 a_2275_4162# a_28978_4138# 0.17fF
C13927 a_24050_6146# ctop 4.91fF
C13928 a_32994_11166# VDD 0.29fF
C13929 m3_22948_1078# m3_23952_1078# 0.21fF
C13930 a_1957_17214# m2_1732_17010# 0.33fF
C13931 m2_1732_4962# sample_n 0.12fF
C13932 a_2275_13198# a_6982_13174# 0.71fF
C13933 col[28] rowoff_n[13] 0.16fF
C13934 a_4882_5142# vcm 0.18fF
C13935 col_n[7] rowoff_n[5] 0.29fF
C13936 col_n[10] rowoff_n[8] 0.27fF
C13937 col_n[3] rowoff_n[1] 0.32fF
C13938 col_n[6] rowoff_n[4] 0.29fF
C13939 col_n[9] rowoff_n[7] 0.27fF
C13940 col_n[4] rowoff_n[2] 0.31fF
C13941 col_n[11] rowoff_n[9] 0.26fF
C13942 col_n[8] rowoff_n[6] 0.28fF
C13943 col_n[5] rowoff_n[3] 0.30fF
C13944 col_n[2] rowoff_n[0] 0.32fF
C13945 a_8990_15182# col[6] 0.38fF
C13946 a_26362_15222# vcm 0.24fF
C13947 a_2475_18218# a_31990_18194# 0.41fF
C13948 a_21038_13174# m2_21236_13422# 0.19fF
C13949 a_28066_17190# row_n[15] 0.43fF
C13950 a_4974_9158# ctop 4.91fF
C13951 a_13918_14178# VDD 0.29fF
C13952 m2_34864_6970# row_n[5] 0.38fF
C13953 a_35002_11166# a_35094_11166# 0.11fF
C13954 a_24050_11166# col_n[21] 0.34fF
C13955 a_4882_2130# rowon_n[0] 0.14fF
C13956 a_2275_15206# a_22042_15182# 0.71fF
C13957 a_2275_12194# col_n[2] 0.17fF
C13958 a_2275_1150# col_n[7] 0.17fF
C13959 a_19942_9158# vcm 0.18fF
C13960 a_4274_15222# col_n[1] 0.11fF
C13961 a_14922_16186# rowoff_n[14] 0.60fF
C13962 a_1957_5166# sample 0.35fF
C13963 a_7286_18234# vcm 0.25fF
C13964 a_20034_13174# ctop 4.91fF
C13965 a_28978_18194# VDD 0.50fF
C13966 col[12] rowoff_n[14] 0.27fF
C13967 a_2475_12194# a_14922_12170# 0.41fF
C13968 a_2275_12194# a_12306_12210# 0.15fF
C13969 a_15014_15182# rowon_n[13] 0.45fF
C13970 m2_28840_18014# m2_29268_18442# 0.19fF
C13971 a_35002_13174# vcm 0.18fF
C13972 a_31078_3134# VDD 1.54fF
C13973 a_12002_11166# m2_12200_11414# 0.19fF
C13974 a_26058_5142# a_27062_5142# 0.86fF
C13975 a_2475_8178# col[12] 0.22fF
C13976 a_25054_5142# rowon_n[3] 0.45fF
C13977 a_3878_17190# rowon_n[15] 0.14fF
C13978 a_2275_9182# a_5886_9158# 0.17fF
C13979 a_2475_18218# m2_12776_18014# 0.62fF
C13980 a_2475_14202# a_29982_14178# 0.41fF
C13981 a_2275_14202# a_27366_14218# 0.15fF
C13982 a_15926_14178# a_16018_14178# 0.45fF
C13983 a_2275_1150# m2_2736_946# 0.48fF
C13984 a_13006_9158# col_n[10] 0.34fF
C13985 m2_1732_6970# m2_1732_5966# 0.84fF
C13986 a_2275_14202# col_n[19] 0.17fF
C13987 a_2275_3158# col_n[24] 0.17fF
C13988 a_31078_7150# m2_31276_7398# 0.19fF
C13989 a_15926_16186# vcm 0.18fF
C13990 a_12002_6146# VDD 3.51fF
C13991 a_17022_7150# a_17022_6146# 0.84fF
C13992 VDD col_n[12] 13.46fF
C13993 vcm col_n[9] 3.22fF
C13994 a_35494_16548# VDD 0.13fF
C13995 a_2275_11190# a_20946_11166# 0.17fF
C13996 a_2275_11190# col[9] 0.17fF
C13997 a_18026_1126# vcm 0.89fF
C13998 a_2161_17214# rowoff_n[15] 0.14fF
C13999 m2_6752_18014# VDD 4.90fF
C14000 a_33086_8154# col[30] 0.38fF
C14001 a_27062_10162# VDD 1.96fF
C14002 a_2475_10186# col[29] 0.22fF
C14003 a_6982_8154# a_7986_8154# 0.86fF
C14004 a_2475_8178# a_13006_8154# 0.68fF
C14005 m2_5748_946# col_n[3] 0.45fF
C14006 a_2275_13198# a_34394_13214# 0.15fF
C14007 a_33086_5142# vcm 0.89fF
C14008 a_27062_12170# rowoff_n[10] 1.45fF
C14009 a_9994_4138# rowoff_n[2] 2.28fF
C14010 a_30986_18194# a_31078_18194# 0.11fF
C14011 a_22042_5142# m2_22240_5390# 0.19fF
C14012 a_28370_8194# col_n[25] 0.11fF
C14013 a_25966_1126# a_26058_1126# 0.11fF
C14014 a_23046_12170# rowon_n[10] 0.45fF
C14015 a_2275_5166# a_3970_5142# 0.71fF
C14016 a_7986_13174# VDD 3.92fF
C14017 a_2475_10186# a_28066_10162# 0.68fF
C14018 a_32082_11166# a_32082_10162# 0.84fF
C14019 a_19030_2130# rowoff_n[0] 1.84fF
C14020 a_33086_2130# rowon_n[0] 0.45fF
C14021 a_2275_13198# col[26] 0.17fF
C14022 a_2275_2154# col[31] 0.17fF
C14023 a_14010_8154# vcm 0.89fF
C14024 a_2966_17190# vcm 0.89fF
C14025 m2_6752_18014# m3_6884_18146# 4.43fF
C14026 a_22042_6146# col[19] 0.38fF
C14027 a_2275_7174# a_19030_7150# 0.71fF
C14028 a_23046_17190# VDD 2.37fF
C14029 a_10998_2130# row_n[0] 0.43fF
C14030 a_22042_12170# a_23046_12170# 0.86fF
C14031 a_10906_6146# rowon_n[4] 0.14fF
C14032 a_4274_2170# vcm 0.24fF
C14033 a_13006_3134# m2_13204_3382# 0.19fF
C14034 a_29070_12170# vcm 0.89fF
C14035 a_25966_2130# VDD 0.29fF
C14036 a_6890_4138# a_6982_4138# 0.45fF
C14037 a_2275_4162# a_9294_4178# 0.15fF
C14038 a_2475_4162# a_11910_4138# 0.41fF
C14039 a_17326_6186# col_n[14] 0.11fF
C14040 a_27366_18234# col_n[24] 0.11fF
C14041 m3_1864_8106# m3_1864_7102# 0.20fF
C14042 a_2275_9182# a_34090_9158# 0.71fF
C14043 a_13006_14178# a_13006_13174# 0.84fF
C14044 a_11910_10162# rowoff_n[8] 0.64fF
C14045 a_2475_17214# col[1] 0.22fF
C14046 col_n[22] rowoff_n[9] 0.18fF
C14047 col_n[15] rowoff_n[2] 0.23fF
C14048 col_n[18] rowoff_n[5] 0.21fF
C14049 col_n[21] rowoff_n[8] 0.19fF
C14050 col_n[16] rowoff_n[3] 0.22fF
C14051 col_n[19] rowoff_n[6] 0.20fF
C14052 col_n[13] rowoff_n[0] 0.24fF
C14053 col_n[20] rowoff_n[7] 0.19fF
C14054 col_n[17] rowoff_n[4] 0.21fF
C14055 col_n[14] rowoff_n[1] 0.24fF
C14056 a_2475_6170# col[6] 0.22fF
C14057 a_19334_6186# vcm 0.24fF
C14058 a_15014_13174# rowoff_n[11] 2.03fF
C14059 m2_1732_1950# VDD 5.46fF
C14060 a_2161_1150# a_2275_1150# 0.17fF
C14061 a_9994_15182# vcm 0.89fF
C14062 a_6890_5142# VDD 0.29fF
C14063 a_2275_6170# a_24354_6186# 0.15fF
C14064 a_2475_6170# a_26970_6146# 0.41fF
C14065 a_31078_9158# rowon_n[7] 0.45fF
C14066 a_20946_8154# rowoff_n[6] 0.54fF
C14067 a_2275_12194# col_n[13] 0.17fF
C14068 a_10998_4138# col[8] 0.38fF
C14069 a_2275_1150# col_n[18] 0.17fF
C14070 a_21038_16186# col[18] 0.38fF
C14071 a_2475_15206# a_4974_15182# 0.68fF
C14072 a_35398_10202# vcm 0.24fF
C14073 a_31078_17190# rowoff_n[15] 1.25fF
C14074 a_2275_3158# a_17934_3134# 0.17fF
C14075 a_3270_12210# col_n[0] 0.11fF
C14076 a_29982_6146# rowoff_n[4] 0.43fF
C14077 a_13006_4138# ctop 4.91fF
C14078 a_6890_1126# m2_6752_946# 0.31fF
C14079 a_2475_1150# m2_15788_946# 0.62fF
C14080 a_21950_9158# VDD 0.29fF
C14081 m3_12908_1078# ctop 0.21fF
C14082 a_8990_9158# row_n[7] 0.43fF
C14083 a_2275_9182# col[3] 0.17fF
C14084 col[23] rowoff_n[14] 0.19fF
C14085 a_21950_8154# a_22042_8154# 0.45fF
C14086 a_8898_13174# rowon_n[11] 0.14fF
C14087 a_6282_4178# col_n[3] 0.11fF
C14088 col_n[6] rowoff_n[10] 0.29fF
C14089 a_16322_16226# col_n[13] 0.11fF
C14090 m2_17796_18014# col[15] 0.39fF
C14091 a_27974_4138# vcm 0.18fF
C14092 a_18938_3134# rowon_n[1] 0.14fF
C14093 a_2475_17214# a_20034_17190# 0.68fF
C14094 a_2475_8178# col[23] 0.22fF
C14095 m2_10768_18014# m2_11772_18014# 0.86fF
C14096 a_15318_13214# vcm 0.24fF
C14097 a_2275_5166# a_32994_5142# 0.17fF
C14098 a_28066_8154# ctop 4.91fF
C14099 a_2161_12194# VDD 0.23fF
C14100 a_2275_14202# col_n[30] 0.17fF
C14101 a_2275_14202# a_10998_14178# 0.71fF
C14102 a_8898_7150# vcm 0.18fF
C14103 a_2874_14178# rowoff_n[12] 0.74fF
C14104 a_9994_14178# col[7] 0.38fF
C14105 a_13006_2130# a_14010_2130# 0.86fF
C14106 a_2475_2154# a_25054_2130# 0.68fF
C14107 VDD col_n[23] 10.73fF
C14108 vcm col_n[20] 3.22fF
C14109 a_30378_17230# vcm 0.24fF
C14110 col[7] rowoff_n[15] 0.30fF
C14111 a_29070_16186# rowon_n[14] 0.45fF
C14112 a_2275_11190# col[20] 0.17fF
C14113 a_8990_11166# ctop 4.91fF
C14114 a_25054_10162# col_n[22] 0.34fF
C14115 a_17934_16186# VDD 0.29fF
C14116 a_2275_16210# a_26058_16186# 0.71fF
C14117 a_5278_14218# col_n[2] 0.11fF
C14118 a_2966_4138# col_n[0] 0.34fF
C14119 a_23958_11166# vcm 0.18fF
C14120 a_20034_1126# VDD 4.83fF
C14121 a_6982_16186# row_n[14] 0.43fF
C14122 m2_33860_18014# col_n[31] 0.34fF
C14123 a_3970_4138# a_3970_3134# 0.84fF
C14124 a_24050_15182# ctop 4.91fF
C14125 a_17022_6146# row_n[4] 0.43fF
C14126 a_2275_13198# a_16322_13214# 0.15fF
C14127 a_2475_13198# a_18938_13174# 0.41fF
C14128 a_16930_10162# rowon_n[8] 0.14fF
C14129 m2_9764_946# vcm 0.71fF
C14130 a_2275_1150# a_31078_1126# 0.14fF
C14131 a_4882_14178# vcm 0.18fF
C14132 a_28066_6146# a_29070_6146# 0.86fF
C14133 a_2275_10186# a_9902_10162# 0.17fF
C14134 a_2475_4162# col[0] 0.20fF
C14135 a_14010_8154# col_n[11] 0.34fF
C14136 m2_1732_946# m2_1732_1950# 0.84fF
C14137 a_17934_15182# a_18026_15182# 0.45fF
C14138 a_2275_15206# a_31382_15222# 0.15fF
C14139 a_2475_15206# a_33998_15182# 0.41fF
C14140 a_3970_4138# rowon_n[2] 0.45fF
C14141 a_2275_10186# col_n[7] 0.17fF
C14142 a_19942_18194# vcm 0.18fF
C14143 a_3970_1126# m3_3872_1078# 3.79fF
C14144 a_16018_8154# VDD 3.09fF
C14145 a_1957_14202# sample 0.35fF
C14146 a_19030_8154# a_19030_7150# 0.84fF
C14147 a_2275_12194# a_24962_12170# 0.17fF
C14148 a_22042_3134# vcm 0.89fF
C14149 a_34090_7150# col[31] 0.38fF
C14150 a_2475_5166# rowoff_n[3] 4.75fF
C14151 a_15014_13174# row_n[11] 0.43fF
C14152 a_31078_12170# VDD 1.54fF
C14153 m3_18932_18146# m3_19936_18146# 0.21fF
C14154 m2_12776_946# m3_12908_1078# 4.41fF
C14155 a_2475_17214# col[12] 0.22fF
C14156 a_14922_17190# rowon_n[15] 0.14fF
C14157 a_8990_9158# a_9994_9158# 0.86fF
C14158 a_2475_9182# a_17022_9158# 0.68fF
C14159 col_n[24] rowoff_n[0] 0.16fF
C14160 col_n[27] rowoff_n[3] 0.14fF
C14161 col_n[30] rowoff_n[6] 0.12fF
C14162 col_n[31] rowoff_n[7] 0.11fF
C14163 col_n[28] rowoff_n[4] 0.14fF
C14164 col_n[25] rowoff_n[1] 0.16fF
C14165 col_n[29] rowoff_n[5] 0.13fF
C14166 col_n[26] rowoff_n[2] 0.15fF
C14167 a_2475_6170# col[17] 0.22fF
C14168 a_25054_3134# row_n[1] 0.43fF
C14169 a_10998_3134# rowoff_n[1] 2.23fF
C14170 a_24962_7150# rowon_n[5] 0.14fF
C14171 a_2874_6146# vcm 0.18fF
C14172 a_29374_7190# col_n[26] 0.11fF
C14173 a_31990_14178# rowoff_n[12] 0.41fF
C14174 a_27974_2130# a_28066_2130# 0.45fF
C14175 a_2275_12194# col_n[24] 0.17fF
C14176 a_27062_14178# m2_27260_14426# 0.19fF
C14177 a_2275_6170# a_7986_6146# 0.71fF
C14178 a_2275_1150# col_n[29] 0.17fF
C14179 a_2275_8178# rowoff_n[6] 0.81fF
C14180 a_12002_15182# VDD 3.51fF
C14181 a_2475_11190# a_32082_11166# 0.68fF
C14182 a_34090_12170# a_34090_11166# 0.84fF
C14183 a_27366_1166# vcm 0.25fF
C14184 a_2475_11190# rowon_n[9] 0.40fF
C14185 a_18026_10162# vcm 0.89fF
C14186 a_2275_9182# col[14] 0.17fF
C14187 a_23046_5142# col[20] 0.38fF
C14188 a_3878_9158# VDD 0.29fF
C14189 m3_8892_18146# ctop 0.21fF
C14190 col_n[17] rowoff_n[10] 0.21fF
C14191 a_33086_17190# col[30] 0.38fF
C14192 a_2275_8178# a_23046_8154# 0.71fF
C14193 a_24050_13174# a_25054_13174# 0.86fF
C14194 a_8290_4178# vcm 0.24fF
C14195 a_33086_14178# vcm 0.89fF
C14196 a_18330_5182# col_n[15] 0.11fF
C14197 m2_34864_8978# rowon_n[7] 0.42fF
C14198 a_29982_4138# VDD 0.29fF
C14199 a_8898_5142# a_8990_5142# 0.45fF
C14200 a_28370_17230# col_n[25] 0.11fF
C14201 a_18026_12170# m2_18224_12418# 0.19fF
C14202 a_2275_5166# a_13310_5182# 0.15fF
C14203 a_2475_5166# a_15926_5142# 0.41fF
C14204 a_2275_18218# a_11910_18194# 0.17fF
C14205 a_23046_10162# row_n[8] 0.43fF
C14206 a_12914_9158# rowoff_n[7] 0.63fF
C14207 a_22954_14178# rowon_n[12] 0.14fF
C14208 a_15014_15182# a_15014_14178# 0.84fF
C14209 vcm col_n[31] 3.32fF
C14210 col_n[0] rowon_n[15] 0.17fF
C14211 VDD rowon_n[14] 4.61fF
C14212 sample row_n[15] 0.92fF
C14213 col[18] rowoff_n[15] 0.23fF
C14214 a_23350_8194# vcm 0.24fF
C14215 a_19942_15182# rowoff_n[13] 0.55fF
C14216 a_2275_2154# a_6890_2130# 0.17fF
C14217 a_2275_11190# col[31] 0.17fF
C14218 a_32994_4138# rowon_n[2] 0.14fF
C14219 a_14010_17190# vcm 0.89fF
C14220 col_n[1] rowoff_n[11] 0.33fF
C14221 a_10906_7150# VDD 0.29fF
C14222 a_21950_7150# rowoff_n[5] 0.52fF
C14223 a_2475_7174# a_30986_7150# 0.41fF
C14224 a_2275_7174# a_28370_7190# 0.15fF
C14225 a_12002_3134# col[9] 0.38fF
C14226 a_22042_15182# col[19] 0.38fF
C14227 a_16930_2130# vcm 0.18fF
C14228 a_2275_8178# col_n[1] 0.17fF
C14229 a_4974_16186# a_5978_16186# 0.86fF
C14230 a_2475_16210# a_8990_16186# 0.68fF
C14231 a_30986_5142# rowoff_n[3] 0.42fF
C14232 a_4274_11206# vcm 0.24fF
C14233 a_1957_1150# VDD 0.70fF
C14234 a_9994_8154# rowon_n[6] 0.45fF
C14235 a_8990_10162# m2_9188_10410# 0.19fF
C14236 a_2275_4162# a_21950_4138# 0.17fF
C14237 a_17022_6146# ctop 4.91fF
C14238 a_7286_3174# col_n[4] 0.11fF
C14239 a_25966_11166# VDD 0.29fF
C14240 m3_8892_1078# m3_9896_1078# 0.21fF
C14241 a_23958_9158# a_24050_9158# 0.45fF
C14242 a_17326_15222# col_n[14] 0.11fF
C14243 m2_1732_2954# vcm 1.11fF
C14244 a_31990_6146# vcm 0.18fF
C14245 a_28066_6146# m2_28264_6394# 0.19fF
C14246 a_19334_15222# vcm 0.24fF
C14247 a_2475_15206# col[6] 0.22fF
C14248 a_2475_18218# a_24962_18194# 0.41fF
C14249 a_2475_4162# col[11] 0.22fF
C14250 m2_13780_946# VDD 5.65fF
C14251 a_32082_10162# ctop 4.91fF
C14252 a_21038_17190# row_n[15] 0.43fF
C14253 a_6890_14178# VDD 0.29fF
C14254 m2_1732_10986# row_n[9] 0.44fF
C14255 a_31078_7150# row_n[5] 0.43fF
C14256 a_2275_15206# a_15014_15182# 0.71fF
C14257 a_10998_13174# col[8] 0.38fF
C14258 m2_34864_11990# m2_35292_12418# 0.19fF
C14259 a_30986_11166# rowon_n[9] 0.14fF
C14260 a_2275_10186# col_n[18] 0.17fF
C14261 a_12914_9158# vcm 0.18fF
C14262 a_7894_16186# rowoff_n[14] 0.68fF
C14263 a_15014_3134# a_16018_3134# 0.86fF
C14264 a_2475_3158# a_29070_3134# 0.68fF
C14265 a_26058_9158# col_n[23] 0.34fF
C14266 a_13006_13174# ctop 4.91fF
C14267 a_21950_18194# VDD 0.50fF
C14268 a_2475_12194# a_7894_12170# 0.41fF
C14269 a_2275_12194# a_5278_12210# 0.15fF
C14270 a_4882_12170# a_4974_12170# 0.45fF
C14271 a_2275_7174# col[8] 0.17fF
C14272 a_6282_13214# col_n[3] 0.11fF
C14273 a_32082_11166# rowoff_n[9] 1.20fF
C14274 a_2275_17214# a_30074_17190# 0.71fF
C14275 a_7986_15182# rowon_n[13] 0.45fF
C14276 m2_21812_18014# m2_22240_18442# 0.19fF
C14277 a_19030_4138# m2_19228_4386# 0.19fF
C14278 a_27974_13174# vcm 0.18fF
C14279 a_24050_3134# VDD 2.27fF
C14280 a_2475_17214# col[23] 0.22fF
C14281 rowon_n[9] rowoff_n[9] 20.66fF
C14282 a_5978_5142# a_5978_4138# 0.84fF
C14283 a_2475_6170# col[28] 0.22fF
C14284 a_18026_5142# rowon_n[3] 0.45fF
C14285 a_28066_17190# ctop 4.93fF
C14286 a_2475_14202# a_22954_14178# 0.41fF
C14287 a_2275_14202# a_20338_14218# 0.15fF
C14288 a_2275_2154# a_35094_2130# 0.14fF
C14289 a_8898_16186# vcm 0.18fF
C14290 a_4974_6146# VDD 4.23fF
C14291 a_30074_7150# a_31078_7150# 0.86fF
C14292 a_15014_7150# col_n[12] 0.34fF
C14293 a_29070_14178# row_n[12] 0.43fF
C14294 a_2275_11190# a_13918_11166# 0.17fF
C14295 a_2275_9182# col[25] 0.17fF
C14296 a_10998_1126# vcm 0.15fF
C14297 a_19942_16186# a_20034_16186# 0.45fF
C14298 col_n[28] rowoff_n[10] 0.14fF
C14299 a_2966_13174# col_n[0] 0.34fF
C14300 a_20034_10162# VDD 2.68fF
C14301 a_2475_8178# a_5978_8154# 0.68fF
C14302 a_21038_9158# a_21038_8154# 0.84fF
C14303 a_2275_13198# a_28978_13174# 0.17fF
C14304 a_26058_5142# vcm 0.89fF
C14305 a_20034_12170# rowoff_n[10] 1.79fF
C14306 a_2874_4138# rowoff_n[2] 0.74fF
C14307 m2_1732_946# a_1957_1150# 0.33fF
C14308 m2_32856_946# vcm 0.82fF
C14309 a_2275_18218# m2_29844_18014# 0.51fF
C14310 a_16018_12170# rowon_n[10] 0.45fF
C14311 a_2475_10186# a_21038_10162# 0.68fF
C14312 a_10998_10162# a_12002_10162# 0.86fF
C14313 col_n[0] row_n[10] 0.37fF
C14314 a_12002_2130# rowoff_n[0] 2.18fF
C14315 col_n[5] row_n[13] 0.37fF
C14316 vcm rowon_n[10] 0.91fF
C14317 sample rowon_n[9] 0.10fF
C14318 col_n[4] rowon_n[12] 0.17fF
C14319 col_n[1] row_n[11] 0.37fF
C14320 col_n[9] row_n[15] 0.37fF
C14321 col_n[7] row_n[14] 0.37fF
C14322 VDD row_n[9] 4.64fF
C14323 col_n[6] rowon_n[13] 0.17fF
C14324 col_n[8] rowon_n[14] 0.17fF
C14325 a_26058_2130# rowon_n[0] 0.45fF
C14326 col_n[10] rowon_n[15] 0.17fF
C14327 col_n[2] rowon_n[11] 0.17fF
C14328 col_n[3] row_n[12] 0.37fF
C14329 col[29] rowoff_n[15] 0.15fF
C14330 a_2475_13198# col[0] 0.20fF
C14331 a_30378_6186# col_n[27] 0.11fF
C14332 a_3970_5142# col_n[1] 0.34fF
C14333 a_2475_2154# col[5] 0.22fF
C14334 a_14010_17190# col_n[11] 0.34fF
C14335 col_n[12] rowoff_n[11] 0.25fF
C14336 a_6982_8154# vcm 0.89fF
C14337 a_29982_3134# a_30074_3134# 0.45fF
C14338 a_3878_7150# rowoff_n[5] 0.73fF
C14339 a_2275_7174# a_12002_7150# 0.71fF
C14340 m2_2736_1950# rowon_n[0] 0.42fF
C14341 a_16018_17190# VDD 3.10fF
C14342 a_3970_2130# row_n[0] 0.43fF
C14343 a_2275_8178# col_n[12] 0.17fF
C14344 a_31382_3174# vcm 0.24fF
C14345 a_22042_12170# vcm 0.89fF
C14346 a_24050_4138# col[21] 0.38fF
C14347 a_18938_2130# VDD 0.29fF
C14348 a_2275_4162# a_3878_4138# 0.17fF
C14349 a_2475_4162# a_4882_4138# 0.41fF
C14350 a_34090_16186# col[31] 0.38fF
C14351 a_2275_5166# col[2] 0.17fF
C14352 m3_1864_15134# m3_1864_14130# 0.20fF
C14353 a_19942_18194# m2_19804_18014# 0.34fF
C14354 a_2275_9182# a_27062_9158# 0.71fF
C14355 a_26058_14178# a_27062_14178# 0.86fF
C14356 a_4882_10162# rowoff_n[8] 0.72fF
C14357 a_2475_15206# col[17] 0.22fF
C14358 a_12306_6186# vcm 0.24fF
C14359 a_7986_13174# rowoff_n[11] 2.38fF
C14360 a_19334_4178# col_n[16] 0.11fF
C14361 a_2475_4162# col[22] 0.22fF
C14362 a_2874_15182# vcm 0.18fF
C14363 a_29374_16226# col_n[26] 0.11fF
C14364 a_33998_6146# VDD 0.29fF
C14365 a_2475_6170# a_19942_6146# 0.41fF
C14366 a_2275_6170# a_17326_6186# 0.15fF
C14367 a_10906_6146# a_10998_6146# 0.45fF
C14368 a_2966_17190# row_n[15] 0.41fF
C14369 a_24050_9158# rowon_n[7] 0.45fF
C14370 a_13918_8154# rowoff_n[6] 0.61fF
C14371 a_2275_10186# col_n[29] 0.17fF
C14372 a_17022_16186# a_17022_15182# 0.84fF
C14373 a_27366_10202# vcm 0.24fF
C14374 a_24050_17190# rowoff_n[15] 1.59fF
C14375 a_22954_6146# rowoff_n[4] 0.51fF
C14376 a_2275_3158# a_10906_3134# 0.17fF
C14377 a_5978_4138# ctop 4.91fF
C14378 a_14922_9158# VDD 0.29fF
C14379 m3_1864_9110# ctop 0.22fF
C14380 a_13006_2130# col[10] 0.38fF
C14381 a_2475_9182# row_n[7] 0.48fF
C14382 a_2275_7174# col[19] 0.17fF
C14383 a_2475_8178# a_35002_8154# 0.41fF
C14384 a_2275_8178# a_32386_8194# 0.15fF
C14385 a_23046_14178# col[20] 0.38fF
C14386 a_3878_18194# VDD 0.50fF
C14387 a_20946_4138# vcm 0.18fF
C14388 a_31990_4138# rowoff_n[2] 0.41fF
C14389 a_11910_3134# rowon_n[1] 0.14fF
C14390 a_6982_17190# a_7986_17190# 0.86fF
C14391 a_2475_17214# a_13006_17190# 0.68fF
C14392 m2_3740_18014# m2_4744_18014# 0.86fF
C14393 a_8290_13214# vcm 0.24fF
C14394 a_8290_2170# col_n[5] 0.11fF
C14395 a_2275_5166# a_25966_5142# 0.17fF
C14396 a_21038_8154# ctop 4.91fF
C14397 a_18330_14218# col_n[15] 0.11fF
C14398 a_29982_13174# VDD 0.29fF
C14399 a_25966_10162# a_26058_10162# 0.45fF
C14400 a_2275_14202# a_3970_14178# 0.71fF
C14401 a_34394_8194# vcm 0.24fF
C14402 a_27062_3134# a_27062_2130# 0.84fF
C14403 a_2475_2154# a_18026_2130# 0.68fF
C14404 a_23350_17230# vcm 0.24fF
C14405 a_22042_16186# rowon_n[14] 0.45fF
C14406 a_33086_15182# m2_33284_15430# 0.19fF
C14407 a_10906_16186# VDD 0.29fF
C14408 a_32082_6146# rowon_n[4] 0.45fF
C14409 a_12002_12170# col[9] 0.38fF
C14410 a_2275_16210# a_19030_16186# 0.71fF
C14411 a_16930_11166# vcm 0.18fF
C14412 a_2275_17214# col_n[1] 0.17fF
C14413 a_13006_1126# VDD 0.13fF
C14414 a_27062_8154# col_n[24] 0.34fF
C14415 a_2275_6170# col_n[6] 0.17fF
C14416 a_2475_4162# a_33086_4138# 0.68fF
C14417 a_17022_4138# a_18026_4138# 0.86fF
C14418 a_1957_10186# VDD 0.28fF
C14419 m2_30848_946# col[28] 0.52fF
C14420 a_16018_17190# m2_15788_18014# 0.84fF
C14421 a_4974_17190# m2_5172_17438# 0.19fF
C14422 a_17022_15182# ctop 4.91fF
C14423 a_9994_6146# row_n[4] 0.43fF
C14424 a_7286_12210# col_n[4] 0.11fF
C14425 a_9902_10162# rowon_n[8] 0.14fF
C14426 a_2966_10162# col[0] 0.38fF
C14427 a_6890_13174# a_6982_13174# 0.45fF
C14428 a_2475_13198# a_11910_13174# 0.41fF
C14429 a_2275_13198# a_9294_13214# 0.15fF
C14430 a_33086_10162# rowoff_n[8] 1.15fF
C14431 a_1957_12194# rowoff_n[10] 0.14fF
C14432 a_2275_1150# a_24050_1126# 0.14fF
C14433 a_31990_15182# vcm 0.18fF
C14434 a_28066_5142# VDD 1.85fF
C14435 a_24050_13174# m2_24248_13422# 0.19fF
C14436 a_7986_6146# a_7986_5142# 0.84fF
C14437 vcm row_n[5] 1.08fF
C14438 col_n[6] row_n[8] 0.37fF
C14439 col_n[12] row_n[11] 0.37fF
C14440 sample row_n[4] 0.92fF
C14441 col_n[4] row_n[7] 0.37fF
C14442 VDD rowon_n[3] 4.61fF
C14443 col_n[20] row_n[15] 0.37fF
C14444 col_n[2] row_n[6] 0.37fF
C14445 col_n[18] row_n[14] 0.37fF
C14446 col_n[16] row_n[13] 0.37fF
C14447 col_n[1] rowon_n[5] 0.17fF
C14448 col_n[0] rowon_n[4] 0.17fF
C14449 col_n[10] row_n[10] 0.37fF
C14450 col_n[19] rowon_n[14] 0.17fF
C14451 col_n[8] row_n[9] 0.37fF
C14452 col_n[17] rowon_n[13] 0.17fF
C14453 col_n[3] rowon_n[6] 0.17fF
C14454 col_n[21] rowon_n[15] 0.17fF
C14455 col_n[5] rowon_n[7] 0.17fF
C14456 col_n[13] rowon_n[11] 0.17fF
C14457 col_n[14] row_n[12] 0.37fF
C14458 col_n[7] rowon_n[8] 0.17fF
C14459 col_n[9] rowon_n[9] 0.17fF
C14460 col_n[11] rowon_n[10] 0.17fF
C14461 col_n[15] rowon_n[12] 0.17fF
C14462 a_2475_13198# col[11] 0.22fF
C14463 a_2161_10186# a_2275_10186# 0.17fF
C14464 a_2475_10186# a_2966_10162# 0.65fF
C14465 a_2475_2154# col[16] 0.22fF
C14466 col_n[23] rowoff_n[11] 0.17fF
C14467 a_2275_15206# a_24354_15222# 0.15fF
C14468 a_2475_15206# a_26970_15182# 0.41fF
C14469 m2_34864_13998# VDD 1.58fF
C14470 a_2475_8178# m2_34864_7974# 0.56fF
C14471 a_12914_18194# vcm 0.18fF
C14472 a_8990_8154# VDD 3.82fF
C14473 a_2275_8178# col_n[23] 0.17fF
C14474 a_16018_6146# col_n[13] 0.34fF
C14475 a_32082_8154# a_33086_8154# 0.86fF
C14476 a_30074_13174# rowon_n[11] 0.45fF
C14477 a_2275_12194# a_17934_12170# 0.17fF
C14478 a_15014_3134# vcm 0.89fF
C14479 a_21950_17190# a_22042_17190# 0.45fF
C14480 a_2275_16210# col[8] 0.17fF
C14481 a_2275_5166# col[13] 0.17fF
C14482 a_15014_11166# m2_15212_11414# 0.19fF
C14483 a_7986_13174# row_n[11] 0.43fF
C14484 a_24050_12170# VDD 2.27fF
C14485 m3_4876_18146# m3_5880_18146# 0.21fF
C14486 a_2475_9182# a_9994_9158# 0.68fF
C14487 a_23046_10162# a_23046_9158# 0.84fF
C14488 a_7894_17190# rowon_n[15] 0.14fF
C14489 col_n[7] rowoff_n[12] 0.29fF
C14490 a_2475_15206# col[28] 0.22fF
C14491 a_2275_14202# a_32994_14178# 0.17fF
C14492 a_18026_3134# row_n[1] 0.43fF
C14493 a_3970_3134# rowoff_n[1] 2.57fF
C14494 a_30074_7150# vcm 0.89fF
C14495 a_17934_7150# rowon_n[5] 0.14fF
C14496 a_24962_14178# rowoff_n[12] 0.49fF
C14497 a_34090_7150# m2_34288_7398# 0.19fF
C14498 a_4974_15182# VDD 4.23fF
C14499 a_2475_11190# a_25054_11166# 0.68fF
C14500 a_13006_11166# a_14010_11166# 0.86fF
C14501 a_4974_4138# col_n[2] 0.34fF
C14502 a_31382_5182# col_n[28] 0.11fF
C14503 a_20338_1166# vcm 0.24fF
C14504 a_15014_16186# col_n[12] 0.34fF
C14505 a_10998_10162# vcm 0.89fF
C14506 a_2275_7174# col[30] 0.17fF
C14507 a_31990_4138# a_32082_4138# 0.45fF
C14508 a_5978_9158# m2_6176_9406# 0.19fF
C14509 a_2275_8178# a_16018_8154# 0.71fF
C14510 a_3970_13174# a_3970_12170# 0.84fF
C14511 row_n[2] rowoff_n[2] 0.64fF
C14512 ctop rowoff_n[9] 0.28fF
C14513 a_2275_4162# vcm 7.71fF
C14514 a_25054_3134# col[22] 0.38fF
C14515 a_25054_5142# m2_25252_5390# 0.19fF
C14516 m2_1732_12994# rowon_n[11] 0.43fF
C14517 a_26058_14178# vcm 0.89fF
C14518 a_22954_4138# VDD 0.29fF
C14519 a_2475_5166# a_8898_5142# 0.41fF
C14520 a_2275_5166# a_6282_5182# 0.15fF
C14521 a_2966_8154# ctop 4.82fF
C14522 a_2275_18218# a_4882_18194# 0.17fF
C14523 a_2275_10186# a_31078_10162# 0.71fF
C14524 a_16018_10162# row_n[8] 0.43fF
C14525 a_5886_9158# rowoff_n[7] 0.70fF
C14526 a_15926_14178# rowon_n[12] 0.14fF
C14527 a_28066_15182# a_29070_15182# 0.86fF
C14528 a_20338_3174# col_n[17] 0.11fF
C14529 a_16322_8194# vcm 0.24fF
C14530 a_12914_15182# rowoff_n[13] 0.63fF
C14531 a_30378_15222# col_n[27] 0.11fF
C14532 a_3970_14178# col_n[1] 0.34fF
C14533 a_25966_4138# rowon_n[2] 0.14fF
C14534 a_2475_11190# col[5] 0.22fF
C14535 a_6982_17190# vcm 0.89fF
C14536 a_29070_3134# ctop 4.91fF
C14537 m2_11772_18014# m3_11904_18146# 4.41fF
C14538 a_14922_7150# rowoff_n[5] 0.60fF
C14539 a_2475_7174# a_23958_7150# 0.41fF
C14540 a_2275_7174# a_21342_7190# 0.15fF
C14541 a_12914_7150# a_13006_7150# 0.45fF
C14542 a_2275_17214# col_n[12] 0.17fF
C14543 a_9902_2130# vcm 0.18fF
C14544 a_19030_17190# a_19030_16186# 0.84fF
C14545 a_2275_6170# col_n[17] 0.17fF
C14546 a_16018_3134# m2_16216_3382# 0.19fF
C14547 a_31382_12210# vcm 0.24fF
C14548 a_23958_5142# rowoff_n[3] 0.50fF
C14549 a_2275_18218# VDD 31.58fF
C14550 a_2874_8154# rowon_n[6] 0.14fF
C14551 a_2275_4162# a_14922_4138# 0.17fF
C14552 a_9994_6146# ctop 4.91fF
C14553 a_24050_13174# col[21] 0.38fF
C14554 a_18938_11166# VDD 0.29fF
C14555 a_2966_9158# a_2966_8154# 0.84fF
C14556 a_2275_14202# col[2] 0.17fF
C14557 a_2275_3158# col[7] 0.17fF
C14558 a_32994_3134# rowoff_n[1] 0.40fF
C14559 a_24962_6146# vcm 0.18fF
C14560 col_n[16] rowon_n[7] 0.17fF
C14561 col_n[14] rowon_n[6] 0.17fF
C14562 a_9294_1166# col_n[6] 0.11fF
C14563 col_n[21] row_n[10] 0.37fF
C14564 col_n[30] rowon_n[14] 0.17fF
C14565 col_n[12] rowon_n[5] 0.17fF
C14566 col_n[19] row_n[9] 0.37fF
C14567 col_n[28] rowon_n[13] 0.17fF
C14568 col_n[10] rowon_n[4] 0.17fF
C14569 col_n[17] row_n[8] 0.37fF
C14570 col_n[1] row_n[0] 0.37fF
C14571 col_n[23] row_n[11] 0.37fF
C14572 col_n[8] rowon_n[3] 0.17fF
C14573 col_n[15] row_n[7] 0.37fF
C14574 col_n[6] rowon_n[2] 0.17fF
C14575 col_n[31] row_n[15] 0.37fF
C14576 col_n[13] row_n[6] 0.37fF
C14577 col_n[20] rowon_n[9] 0.17fF
C14578 VDD en_C0_n 0.37fF
C14579 col_n[18] rowon_n[8] 0.17fF
C14580 col_n[24] rowon_n[11] 0.17fF
C14581 col_n[25] row_n[12] 0.37fF
C14582 col_n[22] rowon_n[10] 0.17fF
C14583 col_n[3] row_n[1] 0.37fF
C14584 col_n[5] row_n[2] 0.37fF
C14585 vcm sw 0.10fF
C14586 col_n[26] rowon_n[12] 0.17fF
C14587 col_n[7] row_n[3] 0.37fF
C14588 col_n[9] row_n[4] 0.37fF
C14589 col_n[27] row_n[13] 0.37fF
C14590 col_n[2] rowon_n[0] 0.17fF
C14591 col_n[11] row_n[5] 0.37fF
C14592 col_n[29] row_n[14] 0.37fF
C14593 col_n[4] rowon_n[1] 0.17fF
C14594 a_12306_15222# vcm 0.24fF
C14595 a_2475_18218# a_17934_18194# 0.41fF
C14596 a_2475_13198# col[22] 0.22fF
C14597 a_19334_13214# col_n[16] 0.11fF
C14598 a_2275_6170# a_29982_6146# 0.17fF
C14599 a_25054_10162# ctop 4.91fF
C14600 a_14010_17190# row_n[15] 0.43fF
C14601 a_2475_2154# col[27] 0.22fF
C14602 a_33998_15182# VDD 0.29fF
C14603 a_27974_11166# a_28066_11166# 0.45fF
C14604 m2_31852_18014# vcm 0.71fF
C14605 a_24050_7150# row_n[5] 0.43fF
C14606 a_2275_15206# a_7986_15182# 0.71fF
C14607 a_23958_11166# rowon_n[9] 0.14fF
C14608 a_5886_9158# vcm 0.18fF
C14609 a_2475_3158# a_22042_3134# 0.68fF
C14610 a_29070_4138# a_29070_3134# 0.84fF
C14611 a_2475_1150# m2_24824_946# 0.62fF
C14612 m3_27968_1078# ctop 0.21fF
C14613 a_5978_13174# ctop 4.91fF
C14614 a_13006_11166# col[10] 0.38fF
C14615 a_14922_18194# VDD 0.50fF
C14616 a_2275_16210# col[19] 0.17fF
C14617 m2_34864_1950# m2_35292_2378# 0.19fF
C14618 a_2275_5166# col[24] 0.17fF
C14619 a_25054_11166# rowoff_n[9] 1.54fF
C14620 a_2275_17214# a_23046_17190# 0.71fF
C14621 m2_14784_18014# m2_15212_18442# 0.19fF
C14622 a_28066_7150# col_n[25] 0.34fF
C14623 a_20946_13174# vcm 0.18fF
C14624 a_17022_3134# VDD 2.99fF
C14625 col_n[18] rowoff_n[12] 0.21fF
C14626 a_19030_5142# a_20034_5142# 0.86fF
C14627 a_10998_5142# rowon_n[3] 0.45fF
C14628 a_2275_18218# a_33086_18194# 0.14fF
C14629 a_8290_11206# col_n[5] 0.11fF
C14630 a_21038_17190# ctop 4.93fF
C14631 a_34090_9158# rowoff_n[7] 1.10fF
C14632 a_2475_14202# a_15926_14178# 0.41fF
C14633 a_2275_14202# a_13310_14218# 0.15fF
C14634 a_8898_14178# a_8990_14178# 0.45fF
C14635 a_2275_2154# a_28066_2130# 0.71fF
C14636 a_34394_17230# vcm 0.24fF
C14637 a_32082_7150# VDD 1.44fF
C14638 a_9994_7150# a_9994_6146# 0.84fF
C14639 m2_33860_946# sw_n 0.69fF
C14640 a_2275_11190# a_6890_11166# 0.17fF
C14641 a_22042_14178# row_n[12] 0.43fF
C14642 a_3970_1126# vcm 0.89fF
C14643 a_2275_16210# a_28370_16226# 0.15fF
C14644 a_2475_16210# a_30986_16186# 0.41fF
C14645 a_32082_4138# row_n[2] 0.43fF
C14646 col_n[2] rowoff_n[13] 0.32fF
C14647 a_31990_8154# rowon_n[6] 0.14fF
C14648 a_17022_5142# col_n[14] 0.34fF
C14649 a_13006_10162# VDD 3.40fF
C14650 a_27062_17190# col_n[24] 0.34fF
C14651 col[5] rowoff_n[9] 0.31fF
C14652 col[0] rowoff_n[4] 0.34fF
C14653 col[1] rowoff_n[5] 0.34fF
C14654 col[2] rowoff_n[6] 0.33fF
C14655 col[3] rowoff_n[7] 0.33fF
C14656 col[4] rowoff_n[8] 0.32fF
C14657 a_2275_15206# col_n[6] 0.17fF
C14658 a_2275_4162# col_n[11] 0.17fF
C14659 a_2275_13198# a_21950_13174# 0.17fF
C14660 a_19030_5142# vcm 0.89fF
C14661 a_13006_12170# rowoff_n[10] 2.13fF
C14662 a_23958_18194# a_24050_18194# 0.11fF
C14663 a_2275_18218# m2_15788_18014# 0.51fF
C14664 a_18938_1126# a_19030_1126# 0.48fF
C14665 a_2275_1150# a_35398_1166# 0.15fF
C14666 a_8990_12170# rowon_n[10] 0.45fF
C14667 a_2275_1150# col[1] 0.17fF
C14668 m2_11772_18014# col[9] 0.37fF
C14669 a_28066_14178# VDD 1.85fF
C14670 a_25054_11166# a_25054_10162# 0.84fF
C14671 a_2475_10186# a_14010_10162# 0.68fF
C14672 a_4974_2130# rowoff_n[0] 2.52fF
C14673 a_19030_2130# rowon_n[0] 0.45fF
C14674 m2_34864_15002# vcm 0.72fF
C14675 a_2475_11190# col[16] 0.22fF
C14676 a_34090_9158# vcm 0.89fF
C14677 a_29070_16186# rowoff_n[14] 1.35fF
C14678 a_28978_1126# m2_28840_946# 0.31fF
C14679 a_2275_7174# a_4974_7150# 0.71fF
C14680 a_3878_7150# a_3970_7150# 0.45fF
C14681 a_5978_3134# col_n[3] 0.34fF
C14682 a_32386_4178# col_n[29] 0.11fF
C14683 a_8990_17190# VDD 3.82fF
C14684 a_2275_17214# col_n[23] 0.17fF
C14685 a_2475_12194# a_29070_12170# 0.68fF
C14686 a_15014_12170# a_16018_12170# 0.86fF
C14687 a_16018_15182# col_n[13] 0.34fF
C14688 a_2275_6170# col_n[28] 0.17fF
C14689 a_2275_18218# col_n[8] 0.17fF
C14690 a_24354_3174# vcm 0.24fF
C14691 a_30074_11166# row_n[9] 0.43fF
C14692 a_29982_15182# rowon_n[13] 0.14fF
C14693 a_2475_3158# m2_1732_2954# 0.16fF
C14694 a_15014_12170# vcm 0.89fF
C14695 a_11910_2130# VDD 0.29fF
C14696 a_33998_5142# a_34090_5142# 0.45fF
C14697 a_2275_14202# col[13] 0.17fF
C14698 a_2275_3158# col[18] 0.17fF
C14699 a_2275_9182# a_20034_9158# 0.71fF
C14700 a_5978_14178# a_5978_13174# 0.84fF
C14701 col_n[12] row_n[0] 0.37fF
C14702 col_n[31] rowon_n[9] 0.17fF
C14703 vcm col[3] 6.66fF
C14704 a_26058_2130# col[23] 0.38fF
C14705 col_n[29] rowon_n[8] 0.17fF
C14706 col_n[27] rowon_n[7] 0.17fF
C14707 col_n[25] rowon_n[6] 0.17fF
C14708 VDD col[6] 11.94fF
C14709 col_n[23] rowon_n[5] 0.17fF
C14710 col_n[30] row_n[9] 0.37fF
C14711 col_n[16] row_n[2] 0.37fF
C14712 col_n[14] row_n[1] 0.37fF
C14713 col_n[18] row_n[3] 0.37fF
C14714 col_n[20] row_n[4] 0.37fF
C14715 col_n[13] rowon_n[0] 0.17fF
C14716 col_n[22] row_n[5] 0.37fF
C14717 col_n[15] rowon_n[1] 0.17fF
C14718 col_n[24] row_n[6] 0.37fF
C14719 col_n[17] rowon_n[2] 0.17fF
C14720 col_n[26] row_n[7] 0.37fF
C14721 col_n[19] rowon_n[3] 0.17fF
C14722 col_n[28] row_n[8] 0.37fF
C14723 col_n[1] col[2] 6.24fF
C14724 col_n[21] rowon_n[4] 0.17fF
C14725 m2_27836_18014# col_n[25] 0.34fF
C14726 a_5278_6186# vcm 0.24fF
C14727 a_2874_18194# a_2966_18194# 0.11fF
C14728 a_30074_16186# vcm 0.89fF
C14729 a_18026_1126# ctop 1.30fF
C14730 a_26970_6146# VDD 0.29fF
C14731 a_2475_6170# a_12914_6146# 0.41fF
C14732 a_2275_6170# a_10298_6186# 0.15fF
C14733 a_30074_14178# m2_30272_14426# 0.19fF
C14734 a_17022_9158# rowon_n[7] 0.45fF
C14735 a_6890_8154# rowoff_n[6] 0.69fF
C14736 a_2275_11190# a_35094_11166# 0.14fF
C14737 a_21342_2170# col_n[18] 0.11fF
C14738 a_32994_1126# vcm 0.18fF
C14739 a_30074_16186# a_31078_16186# 0.86fF
C14740 a_31382_14218# col_n[28] 0.11fF
C14741 a_4974_13174# col_n[2] 0.34fF
C14742 m2_1732_5966# sample 0.31fF
C14743 a_20338_10202# vcm 0.24fF
C14744 a_17022_17190# rowoff_n[15] 1.94fF
C14745 m2_1732_17010# VDD 5.46fF
C14746 a_15926_6146# rowoff_n[4] 0.59fF
C14747 a_2874_3134# a_2966_3134# 0.45fF
C14748 a_33086_5142# ctop 4.91fF
C14749 a_7894_9158# VDD 0.29fF
C14750 m3_23952_18146# ctop 0.21fF
C14751 a_2275_16210# col[30] 0.17fF
C14752 a_2275_8178# a_25358_8194# 0.15fF
C14753 a_2475_8178# a_27974_8154# 0.41fF
C14754 a_1957_16210# m2_1732_16006# 0.33fF
C14755 a_14922_8154# a_15014_8154# 0.45fF
C14756 a_13918_4138# vcm 0.18fF
C14757 a_24962_4138# rowoff_n[2] 0.49fF
C14758 a_4882_3134# rowon_n[1] 0.14fF
C14759 a_2475_17214# a_5978_17190# 0.68fF
C14760 col_n[29] rowoff_n[12] 0.13fF
C14761 a_2275_13198# vcm 7.71fF
C14762 a_25054_12170# col[22] 0.38fF
C14763 a_2275_2154# col_n[5] 0.17fF
C14764 a_2275_5166# a_18938_5142# 0.17fF
C14765 a_21038_12170# m2_21236_12418# 0.19fF
C14766 a_14010_8154# ctop 4.91fF
C14767 a_22954_13174# VDD 0.29fF
C14768 a_2966_17190# ctop 4.83fF
C14769 a_33998_2130# rowoff_n[0] 0.39fF
C14770 a_28978_8154# vcm 0.18fF
C14771 a_20338_12210# col_n[17] 0.11fF
C14772 a_2475_2154# a_10998_2130# 0.68fF
C14773 a_5978_2130# a_6982_2130# 0.86fF
C14774 a_16322_17230# vcm 0.24fF
C14775 a_15014_16186# rowon_n[14] 0.45fF
C14776 a_2275_7174# a_33998_7150# 0.17fF
C14777 a_29070_12170# ctop 4.91fF
C14778 a_2475_9182# col[10] 0.22fF
C14779 a_29982_12170# a_30074_12170# 0.45fF
C14780 a_25054_6146# rowon_n[4] 0.45fF
C14781 col_n[13] rowoff_n[13] 0.24fF
C14782 a_2275_16210# a_12002_16186# 0.71fF
C14783 m2_1732_15002# m2_2160_15430# 0.19fF
C14784 a_9902_11166# vcm 0.18fF
C14785 a_5978_1126# VDD 0.15fF
C14786 col[7] rowoff_n[0] 0.30fF
C14787 col[8] rowoff_n[1] 0.29fF
C14788 col[9] rowoff_n[2] 0.29fF
C14789 col[10] rowoff_n[3] 0.28fF
C14790 col[11] rowoff_n[4] 0.27fF
C14791 col[12] rowoff_n[5] 0.27fF
C14792 col[13] rowoff_n[6] 0.26fF
C14793 col[14] rowoff_n[7] 0.25fF
C14794 col[15] rowoff_n[8] 0.25fF
C14795 col[16] rowoff_n[9] 0.24fF
C14796 a_2275_15206# col_n[17] 0.17fF
C14797 a_2475_4162# a_26058_4138# 0.68fF
C14798 a_31078_5142# a_31078_4138# 0.84fF
C14799 a_12002_10162# m2_12200_10410# 0.19fF
C14800 a_2275_4162# col_n[22] 0.17fF
C14801 m2_1732_1950# row_n[0] 0.44fF
C14802 a_14010_10162# col[11] 0.38fF
C14803 a_9994_15182# ctop 4.91fF
C14804 a_2475_13198# a_4882_13174# 0.41fF
C14805 a_2275_13198# a_3878_13174# 0.17fF
C14806 a_26058_10162# rowoff_n[8] 1.50fF
C14807 a_29070_6146# col_n[26] 0.34fF
C14808 a_2275_12194# col[7] 0.17fF
C14809 a_29982_13174# rowoff_n[11] 0.43fF
C14810 a_2275_1150# a_17022_1126# 0.14fF
C14811 a_31078_6146# m2_31276_6394# 0.19fF
C14812 a_2275_1150# col[12] 0.17fF
C14813 a_24962_15182# vcm 0.18fF
C14814 a_21038_5142# VDD 2.58fF
C14815 m2_22816_946# VDD 4.30fF
C14816 a_9294_10202# col_n[6] 0.11fF
C14817 a_21038_6146# a_22042_6146# 0.86fF
C14818 a_2475_11190# col[27] 0.22fF
C14819 VDD rowoff_n[14] 87.22fF
C14820 a_10906_15182# a_10998_15182# 0.45fF
C14821 a_2475_15206# a_19942_15182# 0.41fF
C14822 a_2275_15206# a_17326_15222# 0.15fF
C14823 col[0] rowoff_n[10] 0.34fF
C14824 a_2275_3158# a_32082_3134# 0.71fF
C14825 a_5886_18194# vcm 0.18fF
C14826 m2_14784_946# col[12] 0.51fF
C14827 a_2475_8178# VDD 41.96fF
C14828 a_12002_8154# a_12002_7150# 0.84fF
C14829 a_23046_13174# rowon_n[11] 0.45fF
C14830 a_2275_18218# col_n[19] 0.17fF
C14831 a_2275_12194# a_10906_12170# 0.17fF
C14832 a_7986_3134# vcm 0.89fF
C14833 m2_34864_4962# rowoff_n[3] 1.01fF
C14834 a_33086_3134# rowon_n[1] 0.45fF
C14835 a_2275_17214# a_32386_17230# 0.15fF
C14836 a_2475_17214# a_35002_17190# 0.41fF
C14837 a_2275_14202# col[24] 0.17fF
C14838 a_22042_4138# m2_22240_4386# 0.19fF
C14839 a_18026_4138# col_n[15] 0.34fF
C14840 a_2275_3158# col[29] 0.17fF
C14841 a_28066_16186# col_n[25] 0.34fF
C14842 a_17022_12170# VDD 2.99fF
C14843 a_1957_9182# a_2275_9182# 0.19fF
C14844 a_2475_9182# a_2874_9158# 0.41fF
C14845 col_n[31] row_n[4] 0.37fF
C14846 col_n[29] row_n[3] 0.37fF
C14847 col_n[27] row_n[2] 0.37fF
C14848 col_n[25] row_n[1] 0.37fF
C14849 col_n[23] row_n[0] 0.37fF
C14850 col_n[26] rowon_n[1] 0.17fF
C14851 VDD col[17] 9.20fF
C14852 col_n[24] rowon_n[0] 0.17fF
C14853 col_n[28] rowon_n[2] 0.17fF
C14854 col_n[7] col[7] 0.50fF
C14855 vcm col[14] 6.66fF
C14856 col_n[30] rowon_n[3] 0.17fF
C14857 a_2275_14202# a_25966_14178# 0.17fF
C14858 a_10998_3134# row_n[1] 0.43fF
C14859 a_23046_7150# vcm 0.89fF
C14860 a_10906_7150# rowon_n[5] 0.14fF
C14861 a_17934_14178# rowoff_n[12] 0.57fF
C14862 a_20946_2130# a_21038_2130# 0.45fF
C14863 a_32082_16186# VDD 1.44fF
C14864 a_27062_12170# a_27062_11166# 0.84fF
C14865 a_2475_11190# a_18026_11166# 0.68fF
C14866 a_13310_1166# vcm 0.25fF
C14867 a_3970_10162# vcm 0.89fF
C14868 a_2475_7174# col[4] 0.22fF
C14869 a_6982_2130# col_n[4] 0.34fF
C14870 a_33390_3174# col_n[30] 0.11fF
C14871 a_2275_8178# a_8990_8154# 0.71fF
C14872 a_17022_14178# col_n[14] 0.34fF
C14873 a_31078_10162# rowon_n[8] 0.45fF
C14874 a_17022_13174# a_18026_13174# 0.86fF
C14875 a_2475_13198# a_33086_13174# 0.68fF
C14876 a_2275_13198# col_n[11] 0.17fF
C14877 a_28370_5182# vcm 0.24fF
C14878 a_2275_2154# col_n[16] 0.17fF
C14879 a_19030_14178# vcm 0.89fF
C14880 a_15926_4138# VDD 0.29fF
C14881 a_2275_10186# a_24050_10162# 0.71fF
C14882 a_2275_10186# col[1] 0.17fF
C14883 a_8990_10162# row_n[8] 0.43fF
C14884 a_8898_14178# rowon_n[12] 0.14fF
C14885 a_7986_15182# a_7986_14178# 0.84fF
C14886 a_9294_8194# vcm 0.24fF
C14887 a_5886_15182# rowoff_n[13] 0.70fF
C14888 a_18938_4138# rowon_n[2] 0.14fF
C14889 a_22042_3134# ctop 4.91fF
C14890 a_34090_18194# vcm 0.15fF
C14891 a_2475_9182# col[21] 0.22fF
C14892 a_30986_8154# VDD 0.29fF
C14893 a_7894_7150# rowoff_n[5] 0.68fF
C14894 a_2275_7174# a_14314_7190# 0.15fF
C14895 a_2475_7174# a_16930_7150# 0.41fF
C14896 a_22346_1166# col_n[19] 0.11fF
C14897 col_n[24] rowoff_n[13] 0.16fF
C14898 a_32386_13214# col_n[29] 0.11fF
C14899 a_5978_12170# col_n[3] 0.34fF
C14900 a_32082_17190# a_33086_17190# 0.86fF
C14901 col[27] rowoff_n[9] 0.17fF
C14902 col[26] rowoff_n[8] 0.17fF
C14903 col[25] rowoff_n[7] 0.18fF
C14904 col[24] rowoff_n[6] 0.19fF
C14905 col[23] rowoff_n[5] 0.19fF
C14906 col[22] rowoff_n[4] 0.20fF
C14907 col[21] rowoff_n[3] 0.21fF
C14908 col[20] rowoff_n[2] 0.21fF
C14909 col[19] rowoff_n[1] 0.22fF
C14910 col[18] rowoff_n[0] 0.23fF
C14911 a_2275_15206# col_n[28] 0.17fF
C14912 a_2966_3134# m2_2736_1950# 0.84fF
C14913 a_24354_12210# vcm 0.24fF
C14914 a_16930_5142# rowoff_n[3] 0.58fF
C14915 a_2275_4162# a_7894_4138# 0.17fF
C14916 a_11910_11166# VDD 0.29fF
C14917 a_29070_17190# rowon_n[15] 0.45fF
C14918 a_2275_9182# a_29374_9198# 0.15fF
C14919 a_2475_9182# a_31990_9158# 0.41fF
C14920 a_16930_9158# a_17022_9158# 0.45fF
C14921 a_2275_12194# col[18] 0.17fF
C14922 a_25966_3134# rowoff_n[1] 0.48fF
C14923 a_2275_1150# col[23] 0.17fF
C14924 a_17934_6146# vcm 0.18fF
C14925 a_26058_11166# col[23] 0.38fF
C14926 a_18026_2130# a_18026_1126# 0.84fF
C14927 a_5278_15222# vcm 0.24fF
C14928 a_2475_18218# a_10906_18194# 0.41fF
C14929 a_2966_5142# VDD 4.45fF
C14930 a_2275_6170# a_22954_6146# 0.17fF
C14931 a_18026_10162# ctop 4.91fF
C14932 a_6982_17190# row_n[15] 0.43fF
C14933 col_n[8] rowoff_n[14] 0.28fF
C14934 a_26970_15182# VDD 0.29fF
C14935 col[11] rowoff_n[10] 0.27fF
C14936 m2_17796_18014# vcm 0.71fF
C14937 a_17022_7150# row_n[5] 0.43fF
C14938 a_16930_11166# rowon_n[9] 0.14fF
C14939 a_21342_11206# col_n[18] 0.11fF
C14940 a_32994_10162# vcm 0.18fF
C14941 a_2475_3158# a_15014_3134# 0.68fF
C14942 a_7986_3134# a_8990_3134# 0.86fF
C14943 a_2275_18218# col_n[30] 0.17fF
C14944 a_2275_1150# m2_7756_946# 0.51fF
C14945 m3_2868_2082# ctop 0.43fF
C14946 a_33086_14178# ctop 4.91fF
C14947 a_7894_18194# VDD 0.50fF
C14948 a_31990_13174# a_32082_13174# 0.45fF
C14949 a_18026_11166# rowoff_n[9] 1.89fF
C14950 a_2275_17214# a_16018_17190# 0.71fF
C14951 m2_7756_18014# m2_8184_18442# 0.19fF
C14952 a_13918_13174# vcm 0.18fF
C14953 a_9994_3134# VDD 3.71fF
C14954 rowon_n[7] row_n[7] 21.02fF
C14955 col_n[31] ctop 0.31fF
C14956 vcm col[25] 6.66fF
C14957 col_n[12] col[13] 6.22fF
C14958 a_15014_9158# col[12] 0.38fF
C14959 VDD col[28] 6.51fF
C14960 a_33086_6146# a_33086_5142# 0.84fF
C14961 a_2475_5166# a_30074_5142# 0.68fF
C14962 a_3970_5142# rowon_n[3] 0.45fF
C14963 a_2275_18218# a_26058_18194# 0.14fF
C14964 a_2275_11190# col_n[5] 0.17fF
C14965 m2_10768_946# m2_11772_946# 0.86fF
C14966 a_14010_17190# ctop 4.93fF
C14967 a_27062_9158# rowoff_n[7] 1.45fF
C14968 a_30074_5142# col_n[27] 0.34fF
C14969 a_2475_14202# a_8898_14178# 0.41fF
C14970 a_2275_14202# a_6282_14218# 0.15fF
C14971 a_34090_15182# rowoff_n[13] 1.10fF
C14972 a_2275_2154# a_21038_2130# 0.71fF
C14973 a_28978_17190# vcm 0.18fF
C14974 a_10298_9198# col_n[7] 0.11fF
C14975 a_25054_7150# VDD 2.16fF
C14976 a_23046_7150# a_24050_7150# 0.86fF
C14977 a_15014_14178# row_n[12] 0.43fF
C14978 a_31078_2130# vcm 0.89fF
C14979 a_2275_16210# a_21342_16226# 0.15fF
C14980 a_2475_16210# a_23958_16186# 0.41fF
C14981 a_12914_16186# a_13006_16186# 0.45fF
C14982 a_2475_7174# col[15] 0.22fF
C14983 a_25054_4138# row_n[2] 0.43fF
C14984 a_24962_8154# rowon_n[6] 0.14fF
C14985 a_5978_10162# VDD 4.13fF
C14986 a_14010_9158# a_14010_8154# 0.84fF
C14987 a_7986_17190# m2_8184_17438# 0.19fF
C14988 a_3970_7150# col[1] 0.38fF
C14989 a_2275_13198# col_n[22] 0.17fF
C14990 a_2275_2154# col_n[27] 0.17fF
C14991 a_2275_13198# a_14922_13174# 0.17fF
C14992 a_12002_5142# vcm 0.89fF
C14993 a_5978_12170# rowoff_n[10] 2.47fF
C14994 a_19030_3134# col_n[16] 0.34fF
C14995 a_2275_18218# m2_1732_18014# 0.27fF
C14996 a_2475_1150# a_28978_1126# 0.41fF
C14997 a_2275_1150# a_26362_1166# 0.15fF
C14998 a_29070_15182# col_n[26] 0.34fF
C14999 a_2475_12194# rowon_n[10] 0.40fF
C15000 a_2275_10186# col[12] 0.17fF
C15001 m3_18932_18146# VDD 0.10fF
C15002 a_27062_13174# m2_27260_13422# 0.19fF
C15003 a_21038_14178# VDD 2.58fF
C15004 a_2475_10186# a_6982_10162# 0.68fF
C15005 a_3970_10162# a_4974_10162# 0.86fF
C15006 a_12002_2130# rowon_n[0] 0.45fF
C15007 a_2275_15206# a_29982_15182# 0.17fF
C15008 a_27062_9158# vcm 0.89fF
C15009 a_22042_16186# rowoff_n[14] 1.69fF
C15010 a_22954_3134# a_23046_3134# 0.45fF
C15011 a_2475_17214# VDD 41.97fF
C15012 sample_n rowoff_n[3] 0.55fF
C15013 col[31] rowoff_n[2] 0.14fF
C15014 col[30] rowoff_n[1] 0.15fF
C15015 col[29] rowoff_n[0] 0.15fF
C15016 a_29070_13174# a_29070_12170# 0.84fF
C15017 a_2475_12194# a_22042_12170# 0.68fF
C15018 a_17326_3174# vcm 0.24fF
C15019 a_23046_11166# row_n[9] 0.43fF
C15020 a_22954_15182# rowon_n[13] 0.14fF
C15021 a_7986_12170# vcm 0.89fF
C15022 a_4882_2130# VDD 0.29fF
C15023 a_18026_11166# m2_18224_11414# 0.19fF
C15024 a_18026_13174# col_n[15] 0.34fF
C15025 a_32994_5142# rowon_n[3] 0.14fF
C15026 a_2275_12194# col[29] 0.17fF
C15027 a_2275_9182# a_13006_9158# 0.71fF
C15028 a_2475_18218# m2_27836_18014# 0.62fF
C15029 a_19030_14178# a_20034_14178# 0.86fF
C15030 a_32386_7190# vcm 0.24fF
C15031 a_2275_9182# col_n[0] 0.17fF
C15032 m2_24824_946# col[22] 0.51fF
C15033 col_n[19] rowoff_n[14] 0.20fF
C15034 a_23046_16186# vcm 0.89fF
C15035 a_19942_6146# VDD 0.29fF
C15036 a_2275_6170# a_3270_6186# 0.15fF
C15037 a_2475_6170# a_5886_6146# 0.41fF
C15038 a_9994_9158# rowon_n[7] 0.45fF
C15039 col[22] rowoff_n[10] 0.20fF
C15040 a_2275_11190# a_28066_11166# 0.71fF
C15041 a_25966_1126# vcm 0.18fF
C15042 a_9994_16186# a_9994_15182# 0.84fF
C15043 m2_1732_3958# rowon_n[2] 0.43fF
C15044 a_13310_10202# vcm 0.24fF
C15045 a_9994_17190# rowoff_n[15] 2.28fF
C15046 m2_21812_18014# VDD 3.33fF
C15047 a_8898_6146# rowoff_n[4] 0.67fF
C15048 a_8990_9158# m2_9188_9406# 0.19fF
C15049 a_26058_5142# ctop 4.91fF
C15050 a_35002_10162# VDD 0.36fF
C15051 a_2475_16210# col[4] 0.22fF
C15052 a_2275_8178# a_18330_8194# 0.15fF
C15053 a_2475_8178# a_20946_8154# 0.41fF
C15054 a_2475_5166# col[9] 0.22fF
C15055 a_33390_12210# col_n[30] 0.11fF
C15056 a_6982_11166# col_n[4] 0.34fF
C15057 m2_2736_1950# m2_3164_2378# 0.19fF
C15058 a_6890_4138# vcm 0.18fF
C15059 a_35002_12170# rowoff_n[10] 0.38fF
C15060 a_17934_4138# rowoff_n[2] 0.57fF
C15061 col_n[3] rowoff_n[15] 0.32fF
C15062 rowon_n[10] ctop 0.37fF
C15063 col_n[18] col[18] 0.50fF
C15064 a_28066_5142# m2_28264_5390# 0.19fF
C15065 a_31078_8154# row_n[6] 0.43fF
C15066 a_28370_14218# vcm 0.24fF
C15067 a_30986_12170# rowon_n[10] 0.14fF
C15068 a_2275_11190# col_n[16] 0.17fF
C15069 a_2275_5166# a_11910_5142# 0.17fF
C15070 a_6982_8154# ctop 4.91fF
C15071 col[6] rowoff_n[11] 0.31fF
C15072 a_15926_13174# VDD 0.29fF
C15073 a_18938_10162# a_19030_10162# 0.45fF
C15074 a_2275_10186# a_33390_10202# 0.15fF
C15075 a_26970_2130# rowoff_n[0] 0.47fF
C15076 a_27062_10162# col[24] 0.38fF
C15077 a_2275_8178# col[6] 0.17fF
C15078 a_21950_8154# vcm 0.18fF
C15079 a_2275_2154# a_2966_2130# 0.14fF
C15080 a_2475_2154# a_3970_2130# 0.68fF
C15081 a_20034_3134# a_20034_2130# 0.84fF
C15082 a_9294_17230# vcm 0.24fF
C15083 a_7986_16186# rowon_n[14] 0.45fF
C15084 m2_16792_18014# m3_16924_18146# 4.41fF
C15085 a_2275_7174# a_26970_7150# 0.17fF
C15086 a_22042_12170# ctop 4.91fF
C15087 a_30986_17190# VDD 0.29fF
C15088 a_2475_7174# col[26] 0.22fF
C15089 a_18026_6146# rowon_n[4] 0.45fF
C15090 a_22346_10202# col_n[19] 0.11fF
C15091 a_2275_16210# a_4974_16186# 0.71fF
C15092 a_3878_16186# a_3970_16186# 0.45fF
C15093 a_19030_3134# m2_19228_3382# 0.19fF
C15094 a_33086_2130# VDD 1.34fF
C15095 a_2475_4162# a_19030_4138# 0.68fF
C15096 a_9994_4138# a_10998_4138# 0.86fF
C15097 a_33998_14178# a_34090_14178# 0.45fF
C15098 a_19030_10162# rowoff_n[8] 1.84fF
C15099 m2_1732_4962# m2_1732_3958# 0.84fF
C15100 a_29070_15182# row_n[13] 0.43fF
C15101 a_22954_13174# rowoff_n[11] 0.51fF
C15102 a_2275_10186# col[23] 0.17fF
C15103 a_2275_1150# a_9994_1126# 0.14fF
C15104 a_16018_8154# col[13] 0.38fF
C15105 a_17934_15182# vcm 0.18fF
C15106 a_14010_5142# VDD 3.30fF
C15107 a_2475_6170# a_34090_6146# 0.68fF
C15108 a_28066_8154# rowoff_n[6] 1.40fF
C15109 a_2966_14178# VDD 4.45fF
C15110 a_31078_4138# col_n[28] 0.34fF
C15111 a_2275_15206# a_10298_15222# 0.15fF
C15112 a_2475_15206# a_12914_15182# 0.41fF
C15113 a_11302_8194# col_n[8] 0.11fF
C15114 a_2275_3158# a_25054_3134# 0.71fF
C15115 a_11910_1126# m2_11772_946# 0.31fF
C15116 a_2275_1150# m2_30848_946# 0.51fF
C15117 a_29070_9158# VDD 1.75fF
C15118 a_25054_8154# a_26058_8154# 0.86fF
C15119 a_16018_13174# rowon_n[11] 0.45fF
C15120 a_2874_12170# a_2966_12170# 0.45fF
C15121 a_35094_4138# vcm 0.15fF
C15122 a_26058_3134# rowon_n[1] 0.45fF
C15123 a_2275_17214# a_25358_17230# 0.15fF
C15124 a_2475_17214# a_27974_17190# 0.41fF
C15125 a_14922_17190# a_15014_17190# 0.45fF
C15126 m2_1732_18014# m2_1732_17010# 0.84fF
C15127 a_2475_3158# col[3] 0.22fF
C15128 a_4974_6146# col[2] 0.38fF
C15129 a_9994_12170# VDD 3.71fF
C15130 a_16018_10162# a_16018_9158# 0.84fF
C15131 a_2275_14202# a_18938_14178# 0.17fF
C15132 a_3970_3134# row_n[1] 0.43fF
C15133 a_2275_9182# col_n[10] 0.17fF
C15134 a_20034_2130# col_n[17] 0.33fF
C15135 col_n[30] rowoff_n[14] 0.12fF
C15136 a_16018_7150# vcm 0.89fF
C15137 a_10906_14178# rowoff_n[12] 0.65fF
C15138 a_30074_14178# col_n[27] 0.34fF
C15139 a_2275_2154# a_30378_2170# 0.15fF
C15140 a_2475_2154# a_32994_2130# 0.41fF
C15141 a_35398_7190# VDD 0.12fF
C15142 a_10298_18234# col_n[7] 0.11fF
C15143 a_25054_16186# VDD 2.16fF
C15144 a_2275_6170# col[0] 0.16fF
C15145 a_5978_11166# a_6982_11166# 0.86fF
C15146 a_2475_11190# a_10998_11166# 0.68fF
C15147 a_6282_1166# vcm 0.25fF
C15148 a_2275_16210# a_33998_16186# 0.17fF
C15149 a_31078_11166# vcm 0.89fF
C15150 a_2475_16210# col[15] 0.22fF
C15151 a_27974_1126# VDD 0.73fF
C15152 a_24962_4138# a_25054_4138# 0.45fF
C15153 a_2475_5166# col[20] 0.22fF
C15154 a_1957_8178# a_2161_8178# 0.11fF
C15155 a_2475_8178# a_2275_8178# 2.96fF
C15156 a_2475_13198# a_26058_13174# 0.68fF
C15157 a_31078_14178# a_31078_13174# 0.84fF
C15158 a_24050_10162# rowon_n[8] 0.45fF
C15159 a_3970_16186# col[1] 0.38fF
C15160 row_n[5] ctop 0.28fF
C15161 col_n[23] col[24] 6.22fF
C15162 col_n[14] rowoff_n[15] 0.24fF
C15163 a_21342_5182# vcm 0.24fF
C15164 a_2275_11190# col_n[27] 0.17fF
C15165 col[17] rowoff_n[11] 0.23fF
C15166 a_12002_14178# vcm 0.89fF
C15167 a_8898_4138# VDD 0.29fF
C15168 a_19030_12170# col_n[16] 0.34fF
C15169 a_2275_10186# a_17022_10162# 0.71fF
C15170 a_2475_10186# row_n[8] 0.48fF
C15171 a_2275_8178# col[17] 0.17fF
C15172 a_21038_15182# a_22042_15182# 0.86fF
C15173 a_3878_8154# vcm 0.18fF
C15174 a_11910_4138# rowon_n[2] 0.14fF
C15175 a_15014_3134# ctop 4.91fF
C15176 a_27062_18194# vcm 0.15fF
C15177 a_23958_8154# VDD 0.29fF
C15178 a_33390_1166# col_n[30] 0.11fF
C15179 a_2275_7174# a_7286_7190# 0.15fF
C15180 a_2475_7174# a_9902_7150# 0.41fF
C15181 a_5886_7150# a_5978_7150# 0.45fF
C15182 a_2275_12194# a_32082_12170# 0.71fF
C15183 a_29982_3134# vcm 0.18fF
C15184 a_12002_17190# a_12002_16186# 0.84fF
C15185 col[1] rowoff_n[12] 0.34fF
C15186 a_9902_5142# rowoff_n[3] 0.66fF
C15187 a_17326_12210# vcm 0.24fF
C15188 a_30074_7150# ctop 4.91fF
C15189 a_4882_11166# VDD 0.29fF
C15190 m3_33992_18146# m3_34996_18146# 0.21fF
C15191 m2_23820_946# m3_23952_1078# 4.41fF
C15192 a_7986_10162# col_n[5] 0.34fF
C15193 a_22042_17190# rowon_n[15] 0.45fF
C15194 a_2275_9182# a_22346_9198# 0.15fF
C15195 a_2475_9182# a_24962_9158# 0.41fF
C15196 a_18938_3134# rowoff_n[1] 0.56fF
C15197 a_10906_6146# vcm 0.18fF
C15198 a_32082_7150# rowon_n[5] 0.45fF
C15199 a_31078_2130# a_32082_2130# 0.86fF
C15200 a_32386_16226# vcm 0.24fF
C15201 a_2275_6170# a_15926_6146# 0.17fF
C15202 a_33086_14178# m2_33284_14426# 0.19fF
C15203 a_10998_10162# ctop 4.91fF
C15204 a_19942_15182# VDD 0.29fF
C15205 a_2275_7174# col_n[4] 0.17fF
C15206 a_20946_11166# a_21038_11166# 0.45fF
C15207 a_28066_9158# col[25] 0.38fF
C15208 m2_3740_18014# vcm 0.71fF
C15209 a_9994_7150# row_n[5] 0.43fF
C15210 a_9902_11166# rowon_n[9] 0.14fF
C15211 a_25966_10162# vcm 0.18fF
C15212 m2_5748_18014# col[3] 0.39fF
C15213 a_22042_4138# a_22042_3134# 0.84fF
C15214 a_2475_3158# a_7986_3134# 0.68fF
C15215 a_2275_4162# ctop 0.14fF
C15216 a_23046_2130# m2_22816_946# 0.84fF
C15217 m3_34996_16138# ctop 0.22fF
C15218 a_4974_16186# m2_5172_16434# 0.19fF
C15219 a_2275_8178# a_30986_8154# 0.17fF
C15220 a_26058_14178# ctop 4.91fF
C15221 a_23350_9198# col_n[20] 0.11fF
C15222 a_2475_14202# col[9] 0.22fF
C15223 a_10998_11166# rowoff_n[9] 2.23fF
C15224 a_2475_3158# col[14] 0.22fF
C15225 a_2275_17214# a_8990_17190# 0.71fF
C15226 a_6890_13174# vcm 0.18fF
C15227 a_2475_18218# col[0] 0.20fF
C15228 a_2874_3134# VDD 0.29fF
C15229 a_24050_12170# m2_24248_12418# 0.19fF
C15230 a_2475_5166# a_23046_5142# 0.68fF
C15231 a_12002_5142# a_13006_5142# 0.86fF
C15232 a_2275_18218# a_19030_18194# 0.14fF
C15233 a_2275_9182# col_n[21] 0.17fF
C15234 a_6982_17190# ctop 4.93fF
C15235 a_20034_9158# rowoff_n[7] 1.79fF
C15236 a_30074_14178# rowon_n[12] 0.45fF
C15237 a_27062_15182# rowoff_n[13] 1.45fF
C15238 a_17022_7150# col[14] 0.38fF
C15239 a_2475_7174# m2_34864_6970# 0.56fF
C15240 a_2275_2154# a_14010_2130# 0.71fF
C15241 a_2275_17214# col[6] 0.17fF
C15242 a_21950_17190# vcm 0.18fF
C15243 a_18026_7150# VDD 2.89fF
C15244 a_29070_7150# rowoff_n[5] 1.35fF
C15245 a_2275_6170# col[11] 0.17fF
C15246 a_32082_3134# col_n[29] 0.34fF
C15247 m2_21812_18014# col_n[19] 0.34fF
C15248 a_7986_14178# row_n[12] 0.43fF
C15249 a_24050_2130# vcm 0.89fF
C15250 a_2475_16210# col[26] 0.22fF
C15251 a_2475_16210# a_16930_16186# 0.41fF
C15252 a_2275_16210# a_14314_16226# 0.15fF
C15253 a_12306_7190# col_n[9] 0.11fF
C15254 a_2475_5166# col[31] 0.22fF
C15255 a_18026_4138# row_n[2] 0.43fF
C15256 a_17934_8154# rowon_n[6] 0.14fF
C15257 a_15014_10162# m2_15212_10410# 0.19fF
C15258 a_2275_4162# a_29070_4138# 0.71fF
C15259 a_33086_11166# VDD 1.34fF
C15260 m3_23952_1078# m3_24956_1078# 0.21fF
C15261 sw ctop 0.54fF
C15262 col_n[25] rowoff_n[15] 0.16fF
C15263 col_n[29] col[29] 0.55fF
C15264 a_27062_9158# a_28066_9158# 0.86fF
C15265 a_2275_17214# m2_1732_17010# 0.27fF
C15266 a_2275_13198# a_7894_13174# 0.17fF
C15267 col[28] rowoff_n[11] 0.16fF
C15268 a_4974_5142# vcm 0.89fF
C15269 a_16930_18194# a_17022_18194# 0.11fF
C15270 a_34090_6146# m2_34288_6394# 0.19fF
C15271 a_2475_1150# a_21950_1126# 0.41fF
C15272 a_2275_1150# a_19334_1166# 0.19fF
C15273 a_11910_1126# a_12002_1126# 0.11fF
C15274 a_5978_5142# col[3] 0.38fF
C15275 a_16018_17190# col[13] 0.38fF
C15276 a_2275_8178# col[28] 0.17fF
C15277 a_14010_14178# VDD 3.30fF
C15278 a_18026_11166# a_18026_10162# 0.84fF
C15279 a_4974_2130# rowon_n[0] 0.45fF
C15280 a_2275_15206# a_22954_15182# 0.17fF
C15281 a_31078_13174# col_n[28] 0.34fF
C15282 a_20034_9158# vcm 0.89fF
C15283 a_15014_16186# rowoff_n[14] 2.03fF
C15284 a_5978_8154# m2_6176_8402# 0.19fF
C15285 a_2275_3158# a_35398_3174# 0.15fF
C15286 a_19030_1126# m2_19228_1374# 0.19fF
C15287 a_11302_17230# col_n[8] 0.11fF
C15288 m2_1732_9982# rowoff_n[8] 2.46fF
C15289 col[12] rowoff_n[12] 0.27fF
C15290 a_7986_12170# a_8990_12170# 0.86fF
C15291 a_2475_12194# a_15014_12170# 0.68fF
C15292 a_10298_3174# vcm 0.24fF
C15293 a_16018_11166# row_n[9] 0.43fF
C15294 a_15926_15182# rowon_n[13] 0.14fF
C15295 a_25054_4138# m2_25252_4386# 0.19fF
C15296 a_35094_13174# vcm 0.15fF
C15297 a_31990_3134# VDD 0.29fF
C15298 a_26970_5142# a_27062_5142# 0.45fF
C15299 a_25966_5142# rowon_n[3] 0.14fF
C15300 a_2475_12194# col[3] 0.22fF
C15301 a_2275_9182# a_5978_9158# 0.71fF
C15302 a_5886_18194# m2_5748_18014# 0.34fF
C15303 a_2475_1150# col[8] 0.22fF
C15304 a_4974_15182# col[2] 0.38fF
C15305 a_2475_18218# m2_13780_18014# 0.62fF
C15306 a_2475_14202# a_30074_14178# 0.68fF
C15307 a_33086_15182# a_33086_14178# 0.84fF
C15308 a_25358_7190# vcm 0.24fF
C15309 a_20034_11166# col_n[17] 0.34fF
C15310 a_3970_1126# ctop 0.63fF
C15311 a_16018_16186# vcm 0.89fF
C15312 a_2275_7174# col_n[15] 0.17fF
C15313 a_12914_6146# VDD 0.29fF
C15314 a_2874_9158# rowon_n[7] 0.14fF
C15315 a_35398_16226# VDD 0.12fF
C15316 a_2275_11190# a_21038_11166# 0.71fF
C15317 a_18938_1126# vcm 0.19fF
C15318 a_2275_15206# col[0] 0.16fF
C15319 a_23046_16186# a_24050_16186# 0.86fF
C15320 a_2275_4162# col[5] 0.17fF
C15321 a_6282_10202# vcm 0.24fF
C15322 a_2874_17190# rowoff_n[15] 0.74fF
C15323 m2_7756_18014# VDD 4.79fF
C15324 a_19030_5142# ctop 4.91fF
C15325 a_27974_10162# VDD 0.29fF
C15326 a_7894_8154# a_7986_8154# 0.45fF
C15327 a_2275_8178# a_11302_8194# 0.15fF
C15328 a_2475_8178# a_13918_8154# 0.41fF
C15329 a_2475_14202# col[20] 0.22fF
C15330 a_2475_3158# col[25] 0.22fF
C15331 a_33998_5142# vcm 0.18fF
C15332 a_2475_18218# col[11] 0.22fF
C15333 a_27974_12170# rowoff_n[10] 0.46fF
C15334 a_10906_4138# rowoff_n[2] 0.65fF
C15335 m2_8760_946# col[6] 0.51fF
C15336 a_24050_8154# row_n[6] 0.43fF
C15337 a_21342_14218# vcm 0.24fF
C15338 a_23958_12170# rowon_n[10] 0.14fF
C15339 a_8990_9158# col_n[6] 0.34fF
C15340 a_2275_5166# a_4882_5142# 0.17fF
C15341 a_2966_5142# a_3970_5142# 0.86fF
C15342 a_34090_9158# ctop 4.80fF
C15343 a_8898_13174# VDD 0.29fF
C15344 a_2275_10186# a_26362_10202# 0.15fF
C15345 a_2475_10186# a_28978_10162# 0.41fF
C15346 a_33998_2130# rowon_n[0] 0.14fF
C15347 a_19942_2130# rowoff_n[0] 0.55fF
C15348 a_1957_9182# rowoff_n[7] 0.14fF
C15349 m2_34864_9982# m2_35292_10410# 0.19fF
C15350 a_2275_17214# col[17] 0.17fF
C15351 a_14922_8154# vcm 0.18fF
C15352 a_2275_6170# col[22] 0.17fF
C15353 a_33086_3134# a_34090_3134# 0.86fF
C15354 a_2275_18218# col[2] 0.17fF
C15355 a_3878_17190# vcm 0.18fF
C15356 a_2275_7174# a_19942_7150# 0.17fF
C15357 a_15014_12170# ctop 4.91fF
C15358 a_23958_17190# VDD 0.29fF
C15359 a_29070_8154# col[26] 0.38fF
C15360 a_22954_12170# a_23046_12170# 0.45fF
C15361 a_10998_6146# rowon_n[4] 0.45fF
C15362 a_29982_12170# vcm 0.18fF
C15363 a_26058_2130# VDD 2.06fF
C15364 row_n[13] sample_n 0.16fF
C15365 ctop col[3] 0.13fF
C15366 a_24050_5142# a_24050_4138# 0.84fF
C15367 a_2475_4162# a_12002_4138# 0.68fF
C15368 m3_34996_8106# m3_34996_7102# 0.20fF
C15369 a_2275_9182# a_35002_9158# 0.17fF
C15370 a_24962_18194# m2_24824_18014# 0.35fF
C15371 a_24354_8194# col_n[21] 0.11fF
C15372 a_30074_16186# ctop 4.91fF
C15373 a_12002_10162# rowoff_n[8] 2.18fF
C15374 a_22042_15182# row_n[13] 0.43fF
C15375 a_15926_13174# rowoff_n[11] 0.59fF
C15376 m2_2736_1950# VDD 4.43fF
C15377 a_2475_1150# a_3878_1126# 0.44fF
C15378 a_2275_1150# a_2874_1126# 0.17fF
C15379 a_10906_15182# vcm 0.18fF
C15380 a_6982_5142# VDD 4.02fF
C15381 a_32082_5142# row_n[3] 0.43fF
C15382 a_14010_6146# a_15014_6146# 0.86fF
C15383 a_2475_6170# a_27062_6146# 0.68fF
C15384 a_31990_9158# rowon_n[7] 0.14fF
C15385 a_21038_8154# rowoff_n[6] 1.74fF
C15386 a_2275_16210# col_n[4] 0.17fF
C15387 a_2475_15206# a_5886_15182# 0.41fF
C15388 a_2275_15206# a_3270_15222# 0.15fF
C15389 a_18026_6146# col[15] 0.38fF
C15390 a_2275_5166# col_n[9] 0.17fF
C15391 a_1957_9182# vcm 0.16fF
C15392 a_31990_17190# rowoff_n[15] 0.41fF
C15393 a_30074_6146# rowoff_n[4] 1.30fF
C15394 a_2275_3158# a_18026_3134# 0.71fF
C15395 a_2475_1150# m2_16792_946# 0.62fF
C15396 a_33086_2130# col_n[30] 0.34fF
C15397 a_22042_9158# VDD 2.47fF
C15398 m3_14916_1078# ctop 0.21fF
C15399 col[23] rowoff_n[12] 0.19fF
C15400 a_4974_8154# a_4974_7150# 0.84fF
C15401 a_8990_13174# rowon_n[11] 0.45fF
C15402 a_2275_13198# ctop 0.14fF
C15403 a_13310_6186# col_n[10] 0.11fF
C15404 a_28066_4138# vcm 0.89fF
C15405 a_19030_3134# rowon_n[1] 0.45fF
C15406 a_2475_17214# a_20946_17190# 0.41fF
C15407 a_2275_17214# a_18330_17230# 0.15fF
C15408 a_23350_18234# col_n[20] 0.11fF
C15409 a_2475_12194# col[14] 0.22fF
C15410 a_2275_5166# a_33086_5142# 0.71fF
C15411 a_2475_1150# col[19] 0.22fF
C15412 a_2874_12170# VDD 0.29fF
C15413 a_2275_18218# a_28370_18234# 0.15fF
C15414 m2_14784_946# m2_15212_1374# 0.19fF
C15415 a_29070_10162# a_30074_10162# 0.86fF
C15416 a_2275_14202# a_11910_14178# 0.17fF
C15417 a_2275_7174# col_n[26] 0.17fF
C15418 a_8990_7150# vcm 0.89fF
C15419 a_6982_4138# col[4] 0.38fF
C15420 a_30074_12170# row_n[10] 0.43fF
C15421 a_2275_2154# a_23350_2170# 0.15fF
C15422 a_2475_2154# a_25966_2130# 0.41fF
C15423 a_13918_2130# a_14010_2130# 0.45fF
C15424 col[7] rowoff_n[13] 0.30fF
C15425 a_17022_16186# col[14] 0.38fF
C15426 a_29982_16186# rowon_n[14] 0.14fF
C15427 a_18026_16186# VDD 2.89fF
C15428 a_2275_15206# col[11] 0.17fF
C15429 a_2275_11190# a_2966_11166# 0.67fF
C15430 a_2475_11190# a_3970_11166# 0.68fF
C15431 a_20034_12170# a_20034_11166# 0.84fF
C15432 a_2275_4162# col[16] 0.17fF
C15433 a_32082_12170# col_n[29] 0.34fF
C15434 a_33390_2170# vcm 0.24fF
C15435 a_2275_16210# a_26970_16186# 0.17fF
C15436 a_2475_2154# m2_1732_1950# 0.16fF
C15437 a_24050_11166# vcm 0.89fF
C15438 a_20946_1126# VDD 0.81fF
C15439 a_12306_16226# col_n[9] 0.11fF
C15440 a_2475_14202# col[31] 0.22fF
C15441 a_10998_17190# m2_11196_17438# 0.19fF
C15442 a_21038_17190# m2_20808_18014# 0.84fF
C15443 a_2475_18218# col[22] 0.22fF
C15444 a_17022_10162# rowon_n[8] 0.45fF
C15445 a_2475_13198# a_19030_13174# 0.68fF
C15446 a_9994_13174# a_10998_13174# 0.86fF
C15447 a_14314_5182# vcm 0.24fF
C15448 m2_10768_946# vcm 0.71fF
C15449 a_2275_1150# a_31990_1126# 0.17fF
C15450 a_4974_14178# vcm 0.89fF
C15451 a_28978_6146# a_29070_6146# 0.45fF
C15452 a_30074_13174# m2_30272_13422# 0.19fF
C15453 a_5978_14178# col[3] 0.38fF
C15454 a_2275_10186# a_9994_10162# 0.71fF
C15455 a_2275_17214# col[28] 0.17fF
C15456 a_2475_15206# a_34090_15182# 0.68fF
C15457 a_2275_18218# col[13] 0.17fF
C15458 a_21038_10162# col_n[18] 0.34fF
C15459 a_29374_9198# vcm 0.24fF
C15460 a_4882_4138# rowon_n[2] 0.14fF
C15461 a_7986_3134# ctop 4.91fF
C15462 a_20034_18194# vcm 0.15fF
C15463 a_16930_8154# VDD 0.29fF
C15464 a_1957_15206# m2_1732_15002# 0.33fF
C15465 a_2275_3158# col_n[3] 0.17fF
C15466 a_2275_12194# a_25054_12170# 0.71fF
C15467 a_22954_3134# vcm 0.18fF
C15468 a_25054_17190# a_26058_17190# 0.86fF
C15469 ctop col[14] 0.13fF
C15470 rowon_n[7] sample_n 0.15fF
C15471 a_2161_5166# rowoff_n[3] 0.14fF
C15472 a_10298_12210# vcm 0.24fF
C15473 a_21038_11166# m2_21236_11414# 0.19fF
C15474 a_23046_7150# ctop 4.91fF
C15475 a_31990_12170# VDD 0.29fF
C15476 m3_19936_18146# m3_20940_18146# 0.21fF
C15477 a_9902_9158# a_9994_9158# 0.45fF
C15478 a_15014_17190# rowon_n[15] 0.45fF
C15479 a_2275_9182# a_15318_9198# 0.15fF
C15480 a_2475_9182# a_17934_9158# 0.41fF
C15481 a_11910_3134# rowoff_n[1] 0.64fF
C15482 a_2475_10186# col[8] 0.22fF
C15483 a_25054_7150# rowon_n[5] 0.45fF
C15484 a_32082_14178# rowoff_n[12] 1.20fF
C15485 a_9994_8154# col_n[7] 0.34fF
C15486 a_25358_16226# vcm 0.24fF
C15487 a_2275_6170# a_8898_6146# 0.17fF
C15488 a_3970_10162# ctop 4.91fF
C15489 a_2275_16210# col_n[15] 0.17fF
C15490 a_2966_8154# rowoff_n[6] 2.62fF
C15491 a_12914_15182# VDD 0.29fF
C15492 a_2275_5166# col_n[20] 0.17fF
C15493 a_2475_11190# a_32994_11166# 0.41fF
C15494 a_2275_11190# a_30378_11206# 0.15fF
C15495 a_18938_10162# vcm 0.18fF
C15496 a_12002_9158# m2_12200_9406# 0.19fF
C15497 a_2275_13198# col[5] 0.17fF
C15498 m3_10900_18146# ctop 0.21fF
C15499 a_2275_2154# col[10] 0.17fF
C15500 a_34394_9198# col_n[31] 0.11fF
C15501 a_2275_8178# a_23958_8154# 0.17fF
C15502 a_30074_7150# col[27] 0.38fF
C15503 a_19030_14178# ctop 4.91fF
C15504 a_24962_13174# a_25054_13174# 0.45fF
C15505 a_2475_12194# col[25] 0.22fF
C15506 a_3970_11166# rowoff_n[9] 2.57fF
C15507 a_1957_17214# a_2161_17214# 0.11fF
C15508 a_2475_17214# a_2275_17214# 2.96fF
C15509 a_2475_1150# col[30] 0.22fF
C15510 a_31078_5142# m2_31276_5390# 0.19fF
C15511 a_33998_14178# vcm 0.18fF
C15512 a_30074_4138# VDD 1.65fF
C15513 a_26058_6146# a_26058_5142# 0.84fF
C15514 a_2475_5166# a_16018_5142# 0.68fF
C15515 a_25358_7190# col_n[22] 0.11fF
C15516 a_2275_18218# a_12002_18194# 0.14fF
C15517 a_13006_9158# rowoff_n[7] 2.13fF
C15518 a_23046_14178# rowon_n[12] 0.45fF
C15519 col[18] rowoff_n[13] 0.23fF
C15520 a_20034_15182# rowoff_n[13] 1.79fF
C15521 m2_34864_9982# VDD 1.58fF
C15522 a_33086_4138# rowon_n[2] 0.45fF
C15523 a_2275_2154# a_6982_2130# 0.71fF
C15524 a_14922_17190# vcm 0.18fF
C15525 col_n[1] rowoff_n[9] 0.33fF
C15526 sample rowoff_n[6] 0.22fF
C15527 m2_21812_18014# m3_21944_18146# 4.42fF
C15528 VDD rowoff_n[5] 87.22fF
C15529 vcm rowoff_n[8] 2.43fF
C15530 col_n[0] rowoff_n[7] 0.34fF
C15531 a_2275_15206# col[22] 0.17fF
C15532 a_10998_7150# VDD 3.61fF
C15533 a_22042_7150# rowoff_n[5] 1.69fF
C15534 a_16018_7150# a_17022_7150# 0.86fF
C15535 a_2475_7174# a_31078_7150# 0.68fF
C15536 a_2275_4162# col[27] 0.17fF
C15537 a_19030_5142# col[16] 0.38fF
C15538 a_17022_2130# vcm 0.89fF
C15539 a_2475_16210# a_9902_16186# 0.41fF
C15540 a_2275_16210# a_7286_16226# 0.15fF
C15541 a_5886_16186# a_5978_16186# 0.45fF
C15542 a_29070_17190# col[26] 0.38fF
C15543 a_22042_3134# m2_22240_3382# 0.19fF
C15544 a_31078_5142# rowoff_n[3] 1.25fF
C15545 a_10998_4138# row_n[2] 0.43fF
C15546 a_2275_1150# VDD 30.20fF
C15547 a_10906_8154# rowon_n[6] 0.14fF
C15548 a_2275_4162# a_22042_4138# 0.71fF
C15549 a_26058_11166# VDD 2.06fF
C15550 m3_9896_1078# m3_10900_1078# 0.21fF
C15551 a_6982_9158# a_6982_8154# 0.84fF
C15552 a_14314_5182# col_n[11] 0.11fF
C15553 a_24354_17230# col_n[21] 0.11fF
C15554 col[2] rowoff_n[14] 0.33fF
C15555 a_32082_6146# vcm 0.89fF
C15556 a_2475_1150# a_14922_1126# 0.41fF
C15557 a_2275_1150# a_12306_1166# 0.15fF
C15558 m2_14784_946# VDD 5.50fF
C15559 a_2475_8178# col[2] 0.22fF
C15560 a_6982_14178# VDD 4.02fF
C15561 a_31078_11166# a_32082_11166# 0.86fF
C15562 a_2275_18218# col[24] 0.17fF
C15563 a_2275_15206# a_15926_15182# 0.17fF
C15564 a_7986_3134# col[5] 0.38fF
C15565 a_31078_11166# rowon_n[9] 0.45fF
C15566 a_13006_9158# vcm 0.89fF
C15567 a_7986_16186# rowoff_n[14] 2.38fF
C15568 a_2275_14202# col_n[9] 0.17fF
C15569 a_18026_15182# col[15] 0.38fF
C15570 a_15926_3134# a_16018_3134# 0.45fF
C15571 a_2275_3158# a_27366_3174# 0.15fF
C15572 a_2475_3158# a_29982_3134# 0.41fF
C15573 a_2275_3158# col_n[14] 0.17fF
C15574 a_33086_11166# col_n[30] 0.34fF
C15575 col_n[0] vcm 3.22fF
C15576 VDD col_n[2] 15.94fF
C15577 row_n[2] sample_n 0.16fF
C15578 ctop col[25] 0.13fF
C15579 a_2475_12194# a_7986_12170# 0.68fF
C15580 a_22042_13174# a_22042_12170# 0.84fF
C15581 a_8990_11166# row_n[9] 0.43fF
C15582 a_3270_3174# vcm 0.24fF
C15583 a_32994_11166# rowoff_n[9] 0.40fF
C15584 a_2275_17214# a_30986_17190# 0.17fF
C15585 a_13310_15222# col_n[10] 0.11fF
C15586 a_8898_15182# rowon_n[13] 0.14fF
C15587 a_28066_13174# vcm 0.89fF
C15588 a_24962_3134# VDD 0.29fF
C15589 a_18938_5142# rowon_n[3] 0.14fF
C15590 m2_26832_946# m2_27836_946# 0.86fF
C15591 a_2475_10186# col[19] 0.22fF
C15592 a_2475_14202# a_23046_14178# 0.68fF
C15593 a_12002_14178# a_13006_14178# 0.86fF
C15594 a_18330_7190# vcm 0.24fF
C15595 a_2275_2154# a_34394_2170# 0.15fF
C15596 a_31078_2130# ctop 4.93fF
C15597 a_2275_16210# col_n[26] 0.17fF
C15598 a_8990_16186# vcm 0.89fF
C15599 a_5886_6146# VDD 0.29fF
C15600 a_6982_13174# col[4] 0.38fF
C15601 a_2275_5166# col_n[31] 0.17fF
C15602 a_30986_7150# a_31078_7150# 0.45fF
C15603 a_2275_11190# a_14010_11166# 0.71fF
C15604 a_22042_9158# col_n[19] 0.34fF
C15605 a_11910_1126# vcm 0.18fF
C15606 a_2275_13198# col[16] 0.17fF
C15607 a_33390_11206# vcm 0.24fF
C15608 a_2275_2154# col[21] 0.17fF
C15609 a_31478_1488# VDD 0.12fF
C15610 a_12002_5142# ctop 4.91fF
C15611 a_5978_2130# m2_5748_946# 0.84fF
C15612 a_20946_10162# VDD 0.29fF
C15613 a_2475_8178# a_6890_8154# 0.41fF
C15614 a_2275_8178# a_4274_8194# 0.15fF
C15615 a_2275_13198# a_29070_13174# 0.71fF
C15616 a_26970_5142# vcm 0.18fF
C15617 a_20946_12170# rowoff_n[10] 0.54fF
C15618 m2_1732_946# a_2275_1150# 0.27fF
C15619 m2_33860_946# vcm 0.42fF
C15620 a_2275_18218# m2_30848_18014# 0.51fF
C15621 a_17022_8154# row_n[6] 0.43fF
C15622 a_14314_14218# vcm 0.24fF
C15623 a_16930_12170# rowon_n[10] 0.14fF
C15624 a_27062_9158# ctop 4.91fF
C15625 a_2475_10186# a_21950_10162# 0.41fF
C15626 a_2275_10186# a_19334_10202# 0.15fF
C15627 a_11910_10162# a_12002_10162# 0.45fF
C15628 a_12914_2130# rowoff_n[0] 0.63fF
C15629 a_26970_2130# rowon_n[0] 0.14fF
C15630 col[29] rowoff_n[13] 0.15fF
C15631 m2_1732_16006# sample_n 0.12fF
C15632 col_n[5] rowoff_n[2] 0.30fF
C15633 col_n[8] rowoff_n[5] 0.28fF
C15634 col_n[11] rowoff_n[8] 0.26fF
C15635 col_n[4] rowoff_n[1] 0.31fF
C15636 col_n[12] rowoff_n[9] 0.25fF
C15637 col_n[9] rowoff_n[6] 0.27fF
C15638 col_n[6] rowoff_n[3] 0.29fF
C15639 a_7894_8154# vcm 0.18fF
C15640 col_n[3] rowoff_n[0] 0.32fF
C15641 col_n[10] rowoff_n[7] 0.27fF
C15642 col_n[7] rowoff_n[4] 0.29fF
C15643 a_1957_15206# rowoff_n[13] 0.14fF
C15644 a_10998_7150# col_n[8] 0.34fF
C15645 a_13006_3134# a_13006_2130# 0.84fF
C15646 a_29374_18234# vcm 0.25fF
C15647 a_2275_7174# a_12914_7150# 0.17fF
C15648 a_7986_12170# ctop 4.91fF
C15649 a_16930_17190# VDD 0.29fF
C15650 a_2275_12194# a_35398_12210# 0.15fF
C15651 a_3970_6146# rowon_n[4] 0.45fF
C15652 a_2275_12194# col_n[3] 0.17fF
C15653 a_2275_1150# col_n[8] 0.17fF
C15654 a_22954_12170# vcm 0.18fF
C15655 a_19030_2130# VDD 2.78fF
C15656 a_2475_4162# a_4974_4138# 0.68fF
C15657 a_31078_6146# col[28] 0.38fF
C15658 m3_34996_15134# m3_34996_14130# 0.20fF
C15659 m2_28840_946# m3_28972_1078# 4.41fF
C15660 a_2275_9182# a_27974_9158# 0.17fF
C15661 col[13] rowoff_n[14] 0.26fF
C15662 a_23046_16186# ctop 4.91fF
C15663 a_26970_14178# a_27062_14178# 0.45fF
C15664 a_4974_10162# rowoff_n[8] 2.52fF
C15665 a_15014_15182# row_n[13] 0.43fF
C15666 a_8898_13174# rowoff_n[11] 0.67fF
C15667 a_2475_8178# col[13] 0.22fF
C15668 a_34090_6146# VDD 1.23fF
C15669 a_26362_6186# col_n[23] 0.11fF
C15670 a_25054_5142# row_n[3] 0.43fF
C15671 a_2475_6170# a_20034_6146# 0.68fF
C15672 a_28066_7150# a_28066_6146# 0.84fF
C15673 a_9994_17190# col_n[7] 0.34fF
C15674 a_24962_9158# rowon_n[7] 0.14fF
C15675 a_14010_8154# rowoff_n[6] 2.08fF
C15676 a_2275_14202# col_n[20] 0.17fF
C15677 a_2275_3158# col_n[25] 0.17fF
C15678 a_24962_17190# rowoff_n[15] 0.49fF
C15679 a_2275_3158# a_10998_3134# 0.71fF
C15680 a_23046_6146# rowoff_n[4] 1.64fF
C15681 a_15014_9158# VDD 3.20fF
C15682 m3_1864_8106# ctop 0.22fF
C15683 VDD col_n[13] 13.21fF
C15684 vcm col_n[10] 3.22fF
C15685 analog_in col[31] 0.14fF
C15686 a_7986_16186# m2_8184_16434# 0.19fF
C15687 a_18026_8154# a_19030_8154# 0.86fF
C15688 a_2475_13198# rowon_n[11] 0.40fF
C15689 a_20034_4138# col[17] 0.38fF
C15690 a_2275_11190# col[10] 0.17fF
C15691 a_34394_18234# col_n[31] 0.11fF
C15692 a_30074_16186# col[27] 0.38fF
C15693 a_21038_4138# vcm 0.89fF
C15694 a_12002_3134# rowon_n[1] 0.45fF
C15695 a_32082_4138# rowoff_n[2] 1.20fF
C15696 a_7894_17190# a_7986_17190# 0.45fF
C15697 a_2475_17214# a_13918_17190# 0.41fF
C15698 a_2275_17214# a_11302_17230# 0.15fF
C15699 a_2475_10186# col[30] 0.22fF
C15700 a_27062_12170# m2_27260_12418# 0.19fF
C15701 a_2275_5166# a_26058_5142# 0.71fF
C15702 a_30074_13174# VDD 1.65fF
C15703 a_2275_18218# a_21342_18234# 0.15fF
C15704 m2_7756_946# m2_8184_1374# 0.19fF
C15705 a_15318_4178# col_n[12] 0.11fF
C15706 a_8990_10162# a_8990_9158# 0.84fF
C15707 a_25358_16226# col_n[22] 0.11fF
C15708 m2_34864_10986# vcm 0.72fF
C15709 a_2275_14202# a_4882_14178# 0.17fF
C15710 a_2966_14178# a_3970_14178# 0.86fF
C15711 a_2475_7174# vcm 1.32fF
C15712 a_23046_12170# row_n[10] 0.43fF
C15713 a_2275_2154# a_16322_2170# 0.15fF
C15714 a_2475_2154# a_18938_2130# 0.41fF
C15715 a_22954_16186# rowon_n[14] 0.14fF
C15716 a_10998_16186# VDD 3.61fF
C15717 a_33086_2130# row_n[0] 0.43fF
C15718 a_33086_12170# a_34090_12170# 0.86fF
C15719 a_32994_6146# rowon_n[4] 0.14fF
C15720 a_2275_13198# col[27] 0.17fF
C15721 a_8990_2130# col[6] 0.38fF
C15722 a_26362_2170# vcm 0.24fF
C15723 a_2275_16210# a_19942_16186# 0.17fF
C15724 a_19030_14178# col[16] 0.38fF
C15725 a_17022_11166# vcm 0.89fF
C15726 a_13918_1126# VDD 0.89fF
C15727 a_17934_4138# a_18026_4138# 0.45fF
C15728 a_18026_10162# m2_18224_10410# 0.19fF
C15729 a_2475_4162# a_33998_4138# 0.41fF
C15730 a_2275_4162# a_31382_4178# 0.15fF
C15731 a_2275_10186# VDD 3.18fF
C15732 a_34090_10162# col_n[31] 0.34fF
C15733 a_4274_2170# col_n[1] 0.11fF
C15734 a_24050_14178# a_24050_13174# 0.84fF
C15735 a_2475_13198# a_12002_13174# 0.68fF
C15736 a_9994_10162# rowon_n[8] 0.45fF
C15737 a_33998_10162# rowoff_n[8] 0.39fF
C15738 a_14314_14218# col_n[11] 0.11fF
C15739 a_7286_5182# vcm 0.24fF
C15740 a_2275_12194# rowoff_n[10] 0.81fF
C15741 a_2275_1150# a_24962_1126# 0.17fF
C15742 a_32082_15182# vcm 0.89fF
C15743 a_28978_5142# VDD 0.29fF
C15744 a_2475_10186# a_3878_10162# 0.41fF
C15745 a_2275_10186# a_2874_10162# 0.17fF
C15746 a_2475_17214# col[2] 0.22fF
C15747 col_n[17] rowoff_n[3] 0.21fF
C15748 col_n[20] rowoff_n[6] 0.19fF
C15749 col_n[23] rowoff_n[9] 0.17fF
C15750 col_n[16] rowoff_n[2] 0.22fF
C15751 col_n[19] rowoff_n[5] 0.20fF
C15752 col_n[14] rowoff_n[0] 0.24fF
C15753 col_n[21] rowoff_n[7] 0.19fF
C15754 col_n[18] rowoff_n[4] 0.21fF
C15755 col_n[15] rowoff_n[1] 0.23fF
C15756 col_n[22] rowoff_n[8] 0.18fF
C15757 a_2475_6170# col[7] 0.22fF
C15758 a_14010_15182# a_15014_15182# 0.86fF
C15759 a_2475_15206# a_27062_15182# 0.68fF
C15760 m2_1732_1950# sample 0.31fF
C15761 a_22346_9198# vcm 0.24fF
C15762 m2_1732_12994# VDD 5.46fF
C15763 a_7986_12170# col[5] 0.38fF
C15764 a_8990_8154# m2_9188_8402# 0.19fF
C15765 a_13006_18194# vcm 0.15fF
C15766 a_9902_8154# VDD 0.29fF
C15767 a_31078_9158# row_n[7] 0.43fF
C15768 a_32994_8154# a_33086_8154# 0.45fF
C15769 a_30986_13174# rowon_n[11] 0.14fF
C15770 a_2275_12194# col_n[14] 0.17fF
C15771 a_2275_1150# col_n[19] 0.17fF
C15772 a_23046_8154# col_n[20] 0.34fF
C15773 a_2275_12194# a_18026_12170# 0.71fF
C15774 a_15926_3134# vcm 0.18fF
C15775 a_4974_17190# a_4974_16186# 0.84fF
C15776 m2_32856_18014# m2_33860_18014# 0.86fF
C15777 a_28066_4138# m2_28264_4386# 0.19fF
C15778 a_3270_12210# vcm 0.24fF
C15779 a_35494_3496# VDD 0.13fF
C15780 a_2275_9182# col[4] 0.17fF
C15781 col[24] rowoff_n[14] 0.19fF
C15782 m2_15788_18014# col_n[13] 0.34fF
C15783 a_16018_7150# ctop 4.91fF
C15784 a_24962_12170# VDD 0.29fF
C15785 m3_5880_18146# m3_6884_18146# 0.21fF
C15786 a_7986_17190# rowon_n[15] 0.45fF
C15787 a_2475_9182# a_10906_9158# 0.41fF
C15788 a_2275_9182# a_8290_9198# 0.15fF
C15789 col_n[7] rowoff_n[10] 0.29fF
C15790 a_2275_14202# a_33086_14178# 0.71fF
C15791 a_4882_3134# rowoff_n[1] 0.72fF
C15792 a_2475_8178# col[24] 0.22fF
C15793 a_18026_7150# rowon_n[5] 0.45fF
C15794 a_30986_7150# vcm 0.18fF
C15795 a_25054_14178# rowoff_n[12] 1.54fF
C15796 a_24050_2130# a_25054_2130# 0.86fF
C15797 a_18330_16226# vcm 0.24fF
C15798 a_31078_11166# ctop 4.91fF
C15799 a_5886_15182# VDD 0.29fF
C15800 a_2275_14202# col_n[31] 0.17fF
C15801 a_2475_11190# a_25966_11166# 0.41fF
C15802 a_2275_11190# a_23350_11206# 0.15fF
C15803 a_13918_11166# a_14010_11166# 0.45fF
C15804 a_12002_6146# col_n[9] 0.34fF
C15805 m2_1732_12994# m2_2160_13422# 0.19fF
C15806 a_11910_10162# vcm 0.18fF
C15807 VDD col_n[24] 10.49fF
C15808 vcm col_n[21] 3.22fF
C15809 col[8] rowoff_n[15] 0.29fF
C15810 a_29070_16186# row_n[14] 0.43fF
C15811 a_15014_4138# a_15014_3134# 0.84fF
C15812 a_2275_11190# col[21] 0.17fF
C15813 a_2275_8178# a_16930_8154# 0.17fF
C15814 a_12002_14178# ctop 4.91fF
C15815 a_2966_4138# vcm 0.89fF
C15816 a_26970_14178# vcm 0.18fF
C15817 a_23046_4138# VDD 2.37fF
C15818 a_32082_5142# col[29] 0.38fF
C15819 a_4974_5142# a_5978_5142# 0.86fF
C15820 a_2475_5166# a_8990_5142# 0.68fF
C15821 a_2275_18218# a_4974_18194# 0.14fF
C15822 a_2275_10186# a_31990_10162# 0.17fF
C15823 a_5978_9158# rowoff_n[7] 2.47fF
C15824 a_16018_14178# rowon_n[12] 0.45fF
C15825 a_28978_15182# a_29070_15182# 0.45fF
C15826 a_13006_15182# rowoff_n[13] 2.13fF
C15827 a_27366_5182# col_n[24] 0.11fF
C15828 a_26058_4138# rowon_n[2] 0.45fF
C15829 a_7894_17190# vcm 0.18fF
C15830 a_10998_16186# col_n[8] 0.34fF
C15831 a_3970_7150# VDD 4.33fF
C15832 a_15014_7150# rowoff_n[5] 2.03fF
C15833 a_2475_7174# a_24050_7150# 0.68fF
C15834 a_30074_8154# a_30074_7150# 0.84fF
C15835 a_2475_4162# col[1] 0.22fF
C15836 a_9994_2130# vcm 0.89fF
C15837 m2_34864_17010# m2_34864_16006# 0.84fF
C15838 a_24050_5142# rowoff_n[3] 1.59fF
C15839 a_3970_4138# row_n[2] 0.43fF
C15840 a_2275_10186# col_n[8] 0.17fF
C15841 a_2275_4162# a_15014_4138# 0.71fF
C15842 a_19030_11166# VDD 2.78fF
C15843 a_21038_3134# col[18] 0.38fF
C15844 a_20034_9158# a_21038_9158# 0.86fF
C15845 a_31078_15182# col[28] 0.38fF
C15846 a_33086_3134# rowoff_n[1] 1.15fF
C15847 a_25054_6146# vcm 0.89fF
C15848 a_9902_18194# a_9994_18194# 0.11fF
C15849 a_4882_1126# a_4974_1126# 0.11fF
C15850 a_2275_1150# a_5278_1166# 0.15fF
C15851 a_2475_1150# a_7894_1126# 0.41fF
C15852 a_16322_3174# col_n[13] 0.11fF
C15853 a_2275_6170# a_30074_6146# 0.71fF
C15854 a_2475_17214# col[13] 0.22fF
C15855 col_n[25] rowoff_n[0] 0.16fF
C15856 col_n[28] rowoff_n[3] 0.14fF
C15857 col_n[31] rowoff_n[6] 0.11fF
C15858 col_n[26] rowoff_n[1] 0.15fF
C15859 col_n[29] rowoff_n[4] 0.13fF
C15860 col_n[30] rowoff_n[5] 0.12fF
C15861 col_n[27] rowoff_n[2] 0.14fF
C15862 a_34090_15182# VDD 1.23fF
C15863 a_26362_15222# col_n[23] 0.11fF
C15864 a_2475_6170# col[18] 0.22fF
C15865 a_10998_11166# a_10998_10162# 0.84fF
C15866 m2_32856_18014# vcm 0.71fF
C15867 a_2275_15206# a_8898_15182# 0.17fF
C15868 a_24050_11166# rowon_n[9] 0.45fF
C15869 a_5978_9158# vcm 0.89fF
C15870 a_2275_12194# col_n[25] 0.17fF
C15871 a_2475_3158# a_22954_3134# 0.41fF
C15872 a_2275_3158# a_20338_3174# 0.15fF
C15873 a_2475_1150# m2_25828_946# 0.62fF
C15874 m3_29976_1078# ctop 0.21fF
C15875 a_2275_1150# col_n[30] 0.18fF
C15876 a_20034_13174# col[17] 0.38fF
C15877 a_2475_11190# row_n[9] 0.48fF
C15878 a_30378_4178# vcm 0.24fF
C15879 a_25966_11166# rowoff_n[9] 0.48fF
C15880 a_2275_17214# a_23958_17190# 0.17fF
C15881 a_2275_9182# col[15] 0.17fF
C15882 a_21038_13174# vcm 0.89fF
C15883 a_17934_3134# VDD 0.29fF
C15884 col_n[18] rowoff_n[10] 0.21fF
C15885 a_19942_5142# a_20034_5142# 0.45fF
C15886 a_11910_5142# rowon_n[3] 0.14fF
C15887 a_2275_18218# a_33998_18194# 0.17fF
C15888 a_5278_1166# col_n[2] 0.11fF
C15889 a_35002_9158# rowoff_n[7] 0.38fF
C15890 a_15318_13214# col_n[12] 0.11fF
C15891 a_26058_15182# a_26058_14178# 0.84fF
C15892 a_2475_14202# a_16018_14178# 0.68fF
C15893 a_11302_7190# vcm 0.24fF
C15894 m2_34864_8978# row_n[7] 0.38fF
C15895 a_2275_2154# a_28978_2130# 0.17fF
C15896 a_2475_16210# vcm 1.32fF
C15897 a_24050_2130# ctop 4.93fF
C15898 a_32994_7150# VDD 0.29fF
C15899 a_2275_11190# a_6982_11166# 0.71fF
C15900 col_n[0] row_n[15] 0.37fF
C15901 vcm rowon_n[15] 0.91fF
C15902 sample rowon_n[14] 0.10fF
C15903 VDD row_n[14] 4.64fF
C15904 a_4882_1126# vcm 0.18fF
C15905 col[19] rowoff_n[15] 0.22fF
C15906 a_16018_16186# a_17022_16186# 0.86fF
C15907 a_2475_16210# a_31078_16186# 0.68fF
C15908 a_26362_11206# vcm 0.24fF
C15909 a_8990_11166# col[6] 0.38fF
C15910 a_24450_1488# VDD 0.14fF
C15911 col_n[2] rowoff_n[11] 0.32fF
C15912 a_32082_8154# rowon_n[6] 0.45fF
C15913 a_4974_5142# ctop 4.91fF
C15914 a_13918_10162# VDD 0.29fF
C15915 a_35002_9158# a_35094_9158# 0.11fF
C15916 a_14010_17190# m2_14208_17438# 0.19fF
C15917 a_24050_7150# col_n[21] 0.34fF
C15918 a_2275_13198# a_22042_13174# 0.71fF
C15919 a_2275_8178# col_n[2] 0.17fF
C15920 a_19942_5142# vcm 0.18fF
C15921 a_13918_12170# rowoff_n[10] 0.61fF
C15922 a_4274_11206# col_n[1] 0.11fF
C15923 a_2275_18218# m2_16792_18014# 0.51fF
C15924 a_1957_1150# sample 0.35fF
C15925 a_9994_8154# row_n[6] 0.43fF
C15926 a_7286_14218# vcm 0.24fF
C15927 a_9902_12170# rowon_n[10] 0.14fF
C15928 a_33086_13174# m2_33284_13422# 0.19fF
C15929 a_20034_9158# ctop 4.91fF
C15930 a_28978_14178# VDD 0.29fF
C15931 a_2475_10186# a_14922_10162# 0.41fF
C15932 a_2275_10186# a_12306_10202# 0.15fF
C15933 a_5886_2130# rowoff_n[0] 0.70fF
C15934 a_19942_2130# rowon_n[0] 0.14fF
C15935 m2_1732_13998# vcm 1.11fF
C15936 a_35002_9158# vcm 0.18fF
C15937 a_29982_16186# rowoff_n[14] 0.43fF
C15938 a_2475_15206# col[7] 0.22fF
C15939 a_2475_4162# col[12] 0.22fF
C15940 a_26058_3134# a_27062_3134# 0.86fF
C15941 a_22346_18234# vcm 0.25fF
C15942 a_4974_15182# m2_5172_15430# 0.19fF
C15943 a_2275_7174# a_5886_7150# 0.17fF
C15944 a_9902_17190# VDD 0.29fF
C15945 a_2275_12194# a_27366_12210# 0.15fF
C15946 a_2475_12194# a_29982_12170# 0.41fF
C15947 a_15926_12170# a_16018_12170# 0.45fF
C15948 a_13006_5142# col_n[10] 0.34fF
C15949 a_2275_10186# col_n[19] 0.17fF
C15950 a_23046_17190# col_n[20] 0.34fF
C15951 a_30074_15182# rowon_n[13] 0.45fF
C15952 a_15926_12170# vcm 0.18fF
C15953 a_12002_2130# VDD 3.51fF
C15954 a_24050_11166# m2_24248_11414# 0.19fF
C15955 a_17022_5142# a_17022_4138# 0.84fF
C15956 a_35494_12532# VDD 0.13fF
C15957 a_2275_9182# a_20946_9158# 0.17fF
C15958 a_16018_16186# ctop 4.91fF
C15959 a_2275_7174# col[9] 0.17fF
C15960 a_7986_15182# row_n[13] 0.43fF
C15961 a_33086_4138# col[30] 0.38fF
C15962 a_2475_17214# col[24] 0.22fF
C15963 a_2475_6170# m2_34864_5966# 0.56fF
C15964 row_n[9] rowoff_n[9] 0.64fF
C15965 a_30986_16186# vcm 0.18fF
C15966 m2_30848_18014# col[28] 0.39fF
C15967 a_2475_6170# col[29] 0.22fF
C15968 a_27062_6146# VDD 1.96fF
C15969 a_18026_5142# row_n[3] 0.43fF
C15970 a_2475_6170# a_13006_6146# 0.68fF
C15971 a_6982_6146# a_7986_6146# 0.86fF
C15972 a_17934_9158# rowon_n[7] 0.14fF
C15973 a_6982_8154# rowoff_n[6] 2.42fF
C15974 m2_34864_11990# rowoff_n[10] 1.02fF
C15975 a_2275_11190# a_34394_11206# 0.15fF
C15976 a_33086_1126# vcm 0.15fF
C15977 a_30986_16186# a_31078_16186# 0.45fF
C15978 a_28370_4178# col_n[25] 0.11fF
C15979 a_17934_17190# rowoff_n[15] 0.57fF
C15980 a_12002_15182# col_n[9] 0.34fF
C15981 a_16018_6146# rowoff_n[4] 1.98fF
C15982 a_15014_9158# m2_15212_9406# 0.19fF
C15983 a_2275_3158# a_3970_3134# 0.71fF
C15984 a_7986_9158# VDD 3.92fF
C15985 m3_25960_18146# ctop 0.21fF
C15986 a_2275_16210# m2_1732_16006# 0.27fF
C15987 a_2475_8178# a_28066_8154# 0.68fF
C15988 a_32082_9158# a_32082_8154# 0.84fF
C15989 a_2275_9182# col[26] 0.17fF
C15990 a_14010_4138# vcm 0.89fF
C15991 a_25054_4138# rowoff_n[2] 1.54fF
C15992 a_4974_3134# rowon_n[1] 0.45fF
C15993 a_2275_17214# a_4274_17230# 0.15fF
C15994 a_2475_17214# a_6890_17190# 0.41fF
C15995 col_n[29] rowoff_n[10] 0.13fF
C15996 a_34090_5142# m2_34288_5390# 0.19fF
C15997 a_2966_13174# vcm 0.89fF
C15998 a_22042_2130# col[19] 0.38fF
C15999 a_2275_5166# a_19030_5142# 0.71fF
C16000 a_23046_13174# VDD 2.37fF
C16001 a_32082_14178# col[29] 0.38fF
C16002 a_2275_18218# a_14314_18234# 0.15fF
C16003 a_22042_10162# a_23046_10162# 0.86fF
C16004 a_34090_2130# rowoff_n[0] 1.10fF
C16005 a_29070_8154# vcm 0.89fF
C16006 a_16018_12170# row_n[10] 0.43fF
C16007 a_6890_2130# a_6982_2130# 0.45fF
C16008 a_5978_7150# m2_6176_7398# 0.19fF
C16009 a_2475_2154# a_11910_2130# 0.41fF
C16010 a_2275_2154# a_9294_2170# 0.15fF
C16011 a_17326_2170# col_n[14] 0.11fF
C16012 m2_26832_18014# m3_26964_18146# 4.44fF
C16013 a_15926_16186# rowon_n[14] 0.14fF
C16014 a_27366_14218# col_n[24] 0.11fF
C16015 a_2275_7174# a_34090_7150# 0.71fF
C16016 col_n[10] row_n[15] 0.37fF
C16017 col_n[8] row_n[14] 0.37fF
C16018 col_n[6] row_n[13] 0.37fF
C16019 col_n[5] rowon_n[12] 0.17fF
C16020 col_n[7] rowon_n[13] 0.17fF
C16021 col_n[1] rowon_n[10] 0.17fF
C16022 col_n[0] rowon_n[9] 0.17fF
C16023 col_n[2] row_n[11] 0.37fF
C16024 col_n[9] rowon_n[14] 0.17fF
C16025 col_n[11] rowon_n[15] 0.17fF
C16026 VDD rowon_n[8] 4.61fF
C16027 col_n[3] rowon_n[11] 0.17fF
C16028 col_n[4] row_n[12] 0.37fF
C16029 sample row_n[9] 0.92fF
C16030 vcm row_n[10] 1.08fF
C16031 a_3970_16186# VDD 4.33fF
C16032 a_26058_2130# row_n[0] 0.43fF
C16033 col[30] rowoff_n[15] 0.15fF
C16034 m2_34864_17010# rowoff_n[15] 1.01fF
C16035 a_13006_12170# a_13006_11166# 0.84fF
C16036 a_25966_6146# rowon_n[4] 0.14fF
C16037 a_2475_13198# col[1] 0.22fF
C16038 a_19334_2170# vcm 0.24fF
C16039 a_2475_2154# col[6] 0.22fF
C16040 col_n[13] rowoff_n[11] 0.24fF
C16041 a_2275_16210# a_12914_16186# 0.17fF
C16042 a_25054_3134# m2_25252_3382# 0.19fF
C16043 a_9994_11166# vcm 0.89fF
C16044 a_6890_1126# VDD 0.97fF
C16045 a_2475_4162# a_26970_4138# 0.41fF
C16046 a_2275_4162# a_24354_4178# 0.15fF
C16047 m2_2736_1950# row_n[0] 0.39fF
C16048 a_2275_8178# col_n[13] 0.17fF
C16049 a_21038_12170# col[18] 0.38fF
C16050 a_2874_10162# rowon_n[8] 0.14fF
C16051 a_2475_13198# a_4974_13174# 0.68fF
C16052 a_26970_10162# rowoff_n[8] 0.47fF
C16053 a_35398_6186# vcm 0.24fF
C16054 a_30074_13174# rowoff_n[11] 1.30fF
C16055 a_3270_8194# col_n[0] 0.11fF
C16056 a_2275_1150# a_17934_1126# 0.17fF
C16057 a_25054_15182# vcm 0.89fF
C16058 a_21950_5142# VDD 0.29fF
C16059 a_2275_5166# col[3] 0.17fF
C16060 m2_23820_946# VDD 4.15fF
C16061 a_21950_6146# a_22042_6146# 0.45fF
C16062 a_16322_12210# col_n[13] 0.11fF
C16063 VDD rowoff_n[12] 87.22fF
C16064 a_2475_15206# col[18] 0.22fF
C16065 a_2475_15206# a_20034_15182# 0.68fF
C16066 a_28066_16186# a_28066_15182# 0.84fF
C16067 a_2475_4162# col[23] 0.22fF
C16068 a_15318_9198# vcm 0.24fF
C16069 a_2275_3158# a_32994_3134# 0.17fF
C16070 a_28066_4138# ctop 4.91fF
C16071 a_5978_18194# vcm 0.15fF
C16072 a_16930_1126# m2_16792_946# 0.31fF
C16073 a_2161_8178# VDD 0.23fF
C16074 a_24050_9158# row_n[7] 0.43fF
C16075 a_23958_13174# rowon_n[11] 0.14fF
C16076 a_2275_10186# col_n[30] 0.17fF
C16077 a_2275_12194# a_10998_12170# 0.71fF
C16078 a_8898_3134# vcm 0.18fF
C16079 a_9994_10162# col[7] 0.38fF
C16080 a_33998_3134# rowon_n[1] 0.14fF
C16081 a_18026_17190# a_19030_17190# 0.86fF
C16082 m2_25828_18014# m2_26832_18014# 0.86fF
C16083 a_30378_13214# vcm 0.24fF
C16084 a_2275_7174# col[20] 0.17fF
C16085 a_8990_7150# ctop 4.91fF
C16086 a_25054_6146# col_n[22] 0.34fF
C16087 a_17934_12170# VDD 0.29fF
C16088 m2_30848_946# m2_31276_1374# 0.19fF
C16089 a_2275_14202# a_26058_14178# 0.71fF
C16090 a_5278_10202# col_n[2] 0.11fF
C16091 rowon_n[5] rowoff_n[5] 20.66fF
C16092 a_23958_7150# vcm 0.18fF
C16093 a_10998_7150# rowon_n[5] 0.45fF
C16094 a_18026_14178# rowoff_n[12] 1.89fF
C16095 a_3970_2130# a_3970_1126# 0.84fF
C16096 a_11302_16226# vcm 0.24fF
C16097 a_24050_11166# ctop 4.91fF
C16098 a_32994_16186# VDD 0.29fF
C16099 m2_1732_12994# rowoff_n[11] 2.46fF
C16100 a_2275_11190# a_16322_11206# 0.15fF
C16101 a_2475_11190# a_18938_11166# 0.41fF
C16102 a_4882_10162# vcm 0.18fF
C16103 a_22042_16186# row_n[14] 0.43fF
C16104 m2_1046_19620# VDD 0.70fF
C16105 a_28066_4138# a_29070_4138# 0.86fF
C16106 a_2275_8178# a_9902_8154# 0.17fF
C16107 a_4974_14178# ctop 4.91fF
C16108 a_32082_6146# row_n[4] 0.43fF
C16109 a_14010_4138# col_n[11] 0.34fF
C16110 a_31990_10162# rowon_n[8] 0.14fF
C16111 a_2275_13198# a_31382_13214# 0.15fF
C16112 a_2475_13198# a_33998_13174# 0.41fF
C16113 a_17934_13174# a_18026_13174# 0.45fF
C16114 a_24050_16186# col_n[21] 0.34fF
C16115 m2_1732_2954# m2_1732_1950# 0.84fF
C16116 m2_28840_946# col_n[26] 0.49fF
C16117 a_2275_17214# col_n[2] 0.17fF
C16118 a_19942_14178# vcm 0.18fF
C16119 a_2275_6170# col_n[7] 0.17fF
C16120 a_16018_4138# VDD 3.09fF
C16121 a_1957_10186# sample 0.35fF
C16122 a_19030_6146# a_19030_5142# 0.84fF
C16123 a_2275_10186# a_24962_10162# 0.17fF
C16124 a_8990_14178# rowon_n[12] 0.45fF
C16125 a_34090_3134# col[31] 0.38fF
C16126 a_5978_15182# rowoff_n[13] 2.47fF
C16127 a_19030_4138# rowon_n[2] 0.45fF
C16128 a_35002_18194# vcm 0.18fF
C16129 col_n[20] rowon_n[14] 0.17fF
C16130 col_n[2] rowon_n[5] 0.17fF
C16131 col_n[9] row_n[9] 0.37fF
C16132 col_n[18] rowon_n[13] 0.17fF
C16133 col_n[7] row_n[8] 0.37fF
C16134 col_n[13] row_n[11] 0.37fF
C16135 col_n[5] row_n[7] 0.37fF
C16136 col_n[21] row_n[15] 0.37fF
C16137 col_n[3] row_n[6] 0.37fF
C16138 col_n[19] row_n[14] 0.37fF
C16139 col_n[17] row_n[13] 0.37fF
C16140 col_n[14] rowon_n[11] 0.17fF
C16141 vcm rowon_n[4] 0.91fF
C16142 col_n[6] rowon_n[7] 0.17fF
C16143 col_n[22] rowon_n[15] 0.17fF
C16144 sample rowon_n[3] 0.10fF
C16145 col_n[11] row_n[10] 0.37fF
C16146 col_n[4] rowon_n[6] 0.17fF
C16147 col_n[15] row_n[12] 0.37fF
C16148 col_n[8] rowon_n[8] 0.17fF
C16149 col_n[0] row_n[4] 0.37fF
C16150 col_n[1] row_n[5] 0.37fF
C16151 col_n[10] rowon_n[9] 0.17fF
C16152 col_n[12] rowon_n[10] 0.17fF
C16153 VDD row_n[3] 4.64fF
C16154 col_n[16] rowon_n[12] 0.17fF
C16155 a_31078_8154# VDD 1.54fF
C16156 a_7986_7150# rowoff_n[5] 2.38fF
C16157 a_2475_13198# col[12] 0.22fF
C16158 a_2475_7174# a_17022_7150# 0.68fF
C16159 a_8990_7150# a_9994_7150# 0.86fF
C16160 a_2475_2154# col[17] 0.22fF
C16161 col_n[24] rowoff_n[11] 0.16fF
C16162 a_2874_2130# vcm 0.18fF
C16163 a_29374_3174# col_n[26] 0.11fF
C16164 a_32994_17190# a_33086_17190# 0.45fF
C16165 a_13006_14178# col_n[10] 0.34fF
C16166 a_17022_5142# rowoff_n[3] 1.94fF
C16167 a_2275_8178# col_n[24] 0.17fF
C16168 a_2275_4162# a_7986_4138# 0.71fF
C16169 a_30074_13174# row_n[11] 0.43fF
C16170 a_12002_11166# VDD 3.51fF
C16171 m2_33860_946# m3_33992_1078# 1.28fF
C16172 a_29982_17190# rowon_n[15] 0.14fF
C16173 a_34090_10162# a_34090_9158# 0.84fF
C16174 a_2475_9182# a_32082_9158# 0.68fF
C16175 m2_34864_10986# rowon_n[9] 0.42fF
C16176 a_26058_3134# rowoff_n[1] 1.50fF
C16177 a_2275_16210# col[9] 0.17fF
C16178 a_18026_6146# vcm 0.89fF
C16179 a_2275_5166# col[14] 0.17fF
C16180 a_3878_5142# VDD 0.29fF
C16181 a_33086_13174# col[30] 0.38fF
C16182 a_2275_6170# a_23046_6146# 0.71fF
C16183 col_n[8] rowoff_n[12] 0.28fF
C16184 a_2475_15206# col[29] 0.22fF
C16185 a_27062_15182# VDD 1.96fF
C16186 a_24050_11166# a_25054_11166# 0.86fF
C16187 m2_18800_18014# vcm 0.71fF
C16188 a_17022_11166# rowon_n[9] 0.45fF
C16189 a_33086_10162# vcm 0.89fF
C16190 a_28370_13214# col_n[25] 0.11fF
C16191 a_2475_3158# a_15926_3134# 0.41fF
C16192 a_2275_3158# a_13310_3174# 0.15fF
C16193 a_8898_3134# a_8990_3134# 0.45fF
C16194 a_28066_2130# m2_27836_946# 0.84fF
C16195 a_2275_1150# m2_8760_946# 0.51fF
C16196 a_10998_16186# m2_11196_16434# 0.19fF
C16197 a_15014_13174# a_15014_12170# 0.84fF
C16198 a_23350_4178# vcm 0.24fF
C16199 a_18938_11166# rowoff_n[9] 0.56fF
C16200 a_2275_17214# a_16930_17190# 0.17fF
C16201 a_2275_7174# col[31] 0.17fF
C16202 a_14010_13174# vcm 0.89fF
C16203 a_10906_3134# VDD 0.29fF
C16204 a_2475_5166# a_30986_5142# 0.41fF
C16205 a_2275_5166# a_28370_5182# 0.15fF
C16206 a_30074_12170# m2_30272_12418# 0.19fF
C16207 a_4882_5142# rowon_n[3] 0.14fF
C16208 a_2275_18218# a_26970_18194# 0.17fF
C16209 a_22042_11166# col[19] 0.38fF
C16210 ctop rowoff_n[8] 0.28fF
C16211 a_27974_9158# rowoff_n[7] 0.46fF
C16212 a_2275_4162# col_n[1] 0.17fF
C16213 a_2475_14202# a_8990_14178# 0.68fF
C16214 a_4974_14178# a_5978_14178# 0.86fF
C16215 a_4274_7190# vcm 0.24fF
C16216 m2_1732_12994# row_n[11] 0.44fF
C16217 a_35002_15182# rowoff_n[13] 0.38fF
C16218 a_2275_2154# a_21950_2130# 0.17fF
C16219 a_17022_2130# ctop 4.93fF
C16220 a_29070_17190# vcm 0.89fF
C16221 a_25966_7150# VDD 0.29fF
C16222 a_1957_14202# m2_1732_13998# 0.33fF
C16223 a_23958_7150# a_24050_7150# 0.45fF
C16224 a_17326_11206# col_n[14] 0.11fF
C16225 a_31990_2130# vcm 0.18fF
C16226 a_2475_16210# a_24050_16186# 0.68fF
C16227 a_30074_17190# a_30074_16186# 0.84fF
C16228 a_19334_11206# vcm 0.24fF
C16229 a_2475_11190# col[6] 0.22fF
C16230 a_17422_1488# VDD 0.15fF
C16231 a_25054_8154# rowon_n[6] 0.45fF
C16232 a_21038_10162# m2_21236_10410# 0.19fF
C16233 a_32082_6146# ctop 4.91fF
C16234 a_6890_10162# VDD 0.29fF
C16235 a_2275_17214# col_n[13] 0.17fF
C16236 a_2275_13198# a_15014_13174# 0.71fF
C16237 a_10998_9158# col[8] 0.38fF
C16238 a_2275_6170# col_n[18] 0.17fF
C16239 a_12914_5142# vcm 0.18fF
C16240 a_6890_12170# rowoff_n[10] 0.69fF
C16241 a_2275_18218# m2_2736_18014# 0.48fF
C16242 a_35398_15222# vcm 0.24fF
C16243 a_26058_5142# col_n[23] 0.34fF
C16244 a_3270_17230# col_n[0] 0.11fF
C16245 a_13006_9158# ctop 4.91fF
C16246 a_2275_14202# col[3] 0.17fF
C16247 a_21950_14178# VDD 0.29fF
C16248 a_2275_10186# a_5278_10202# 0.15fF
C16249 a_2475_10186# a_7894_10162# 0.41fF
C16250 a_4882_10162# a_4974_10162# 0.45fF
C16251 a_2275_3158# col[8] 0.17fF
C16252 a_12914_2130# rowon_n[0] 0.14fF
C16253 a_6282_9198# col_n[3] 0.11fF
C16254 a_2275_15206# a_30074_15182# 0.71fF
C16255 col_n[19] rowon_n[8] 0.17fF
C16256 col_n[26] row_n[12] 0.37fF
C16257 col_n[25] rowon_n[11] 0.17fF
C16258 col_n[17] rowon_n[7] 0.17fF
C16259 col_n[15] rowon_n[6] 0.17fF
C16260 col_n[22] row_n[10] 0.37fF
C16261 a_27974_9158# vcm 0.18fF
C16262 col_n[31] rowon_n[14] 0.17fF
C16263 col_n[13] rowon_n[5] 0.17fF
C16264 col_n[20] row_n[9] 0.37fF
C16265 col_n[29] rowon_n[13] 0.17fF
C16266 col_n[11] rowon_n[4] 0.17fF
C16267 col_n[18] row_n[8] 0.37fF
C16268 col_n[24] row_n[11] 0.37fF
C16269 col_n[9] rowon_n[3] 0.17fF
C16270 col_n[4] row_n[1] 0.37fF
C16271 col_n[23] rowon_n[10] 0.17fF
C16272 col_n[2] row_n[0] 0.37fF
C16273 col_n[21] rowon_n[9] 0.17fF
C16274 col_n[6] row_n[2] 0.37fF
C16275 col_n[27] rowon_n[12] 0.17fF
C16276 col_n[8] row_n[3] 0.37fF
C16277 rowon_n[15] row_n[15] 21.02fF
C16278 col_n[10] row_n[4] 0.37fF
C16279 col_n[28] row_n[13] 0.37fF
C16280 col_n[3] rowon_n[0] 0.17fF
C16281 col_n[12] row_n[5] 0.37fF
C16282 col_n[30] row_n[14] 0.37fF
C16283 col_n[5] rowon_n[1] 0.17fF
C16284 VDD en_bit_n[1] 0.35fF
C16285 col_n[14] row_n[6] 0.37fF
C16286 col_n[7] rowon_n[2] 0.17fF
C16287 col_n[16] row_n[7] 0.37fF
C16288 a_22954_16186# rowoff_n[14] 0.51fF
C16289 a_2475_13198# col[23] 0.22fF
C16290 a_12002_8154# m2_12200_8402# 0.19fF
C16291 a_5978_3134# a_5978_2130# 0.84fF
C16292 a_15318_18234# vcm 0.25fF
C16293 a_2475_2154# col[28] 0.22fF
C16294 a_28066_13174# ctop 4.91fF
C16295 a_2161_17214# VDD 0.23fF
C16296 a_2275_12194# a_20338_12210# 0.15fF
C16297 a_2475_12194# a_22954_12170# 0.41fF
C16298 a_23046_15182# rowon_n[13] 0.45fF
C16299 a_31078_4138# m2_31276_4386# 0.19fF
C16300 a_8898_12170# vcm 0.18fF
C16301 a_4974_2130# VDD 4.23fF
C16302 a_30074_5142# a_31078_5142# 0.86fF
C16303 a_33086_5142# rowon_n[3] 0.45fF
C16304 a_15014_3134# col_n[12] 0.34fF
C16305 a_10906_18194# m2_10768_18014# 0.34fF
C16306 a_2275_9182# a_13918_9158# 0.17fF
C16307 a_2275_16210# col[20] 0.17fF
C16308 a_8990_16186# ctop 4.91fF
C16309 a_25054_15182# col_n[22] 0.34fF
C16310 a_2275_5166# col[25] 0.17fF
C16311 a_2475_18218# m2_28840_18014# 0.62fF
C16312 a_19942_14178# a_20034_14178# 0.45fF
C16313 a_2966_9158# col_n[0] 0.34fF
C16314 a_23958_16186# vcm 0.18fF
C16315 col_n[19] rowoff_n[12] 0.20fF
C16316 a_20034_6146# VDD 2.68fF
C16317 a_10998_5142# row_n[3] 0.43fF
C16318 a_2475_6170# a_5978_6146# 0.68fF
C16319 a_21038_7150# a_21038_6146# 0.84fF
C16320 a_10906_9158# rowon_n[7] 0.14fF
C16321 a_2275_11190# a_28978_11166# 0.17fF
C16322 a_26058_1126# vcm 0.15fF
C16323 a_10906_17190# rowoff_n[15] 0.65fF
C16324 m2_22816_18014# VDD 3.26fF
C16325 a_8990_6146# rowoff_n[4] 2.33fF
C16326 m2_33860_946# ctop 0.95fF
C16327 a_2475_8178# a_21038_8154# 0.68fF
C16328 a_10998_8154# a_12002_8154# 0.86fF
C16329 a_30378_2170# col_n[27] 0.11fF
C16330 a_3970_1126# col_n[1] 0.39fF
C16331 a_2475_9182# col[0] 0.20fF
C16332 a_14010_13174# col_n[11] 0.34fF
C16333 a_6982_4138# vcm 0.89fF
C16334 a_18026_4138# rowoff_n[2] 1.89fF
C16335 a_35002_18194# a_35094_18194# 0.11fF
C16336 col_n[3] rowoff_n[13] 0.32fF
C16337 a_29982_1126# a_30074_1126# 0.11fF
C16338 a_31078_12170# rowon_n[10] 0.45fF
C16339 a_2275_5166# a_12002_5142# 0.71fF
C16340 col[4] rowoff_n[7] 0.32fF
C16341 col[3] rowoff_n[6] 0.33fF
C16342 col[2] rowoff_n[5] 0.33fF
C16343 col[1] rowoff_n[4] 0.34fF
C16344 col[0] rowoff_n[3] 0.34fF
C16345 col[5] rowoff_n[8] 0.31fF
C16346 col[6] rowoff_n[9] 0.31fF
C16347 a_2275_15206# col_n[7] 0.17fF
C16348 a_16018_13174# VDD 3.09fF
C16349 a_2275_18218# a_7286_18234# 0.15fF
C16350 a_2275_4162# col_n[12] 0.17fF
C16351 a_27062_2130# rowoff_n[0] 1.45fF
C16352 a_22042_8154# vcm 0.89fF
C16353 m2_9764_18014# col_n[7] 0.34fF
C16354 a_8990_12170# row_n[10] 0.43fF
C16355 a_34090_12170# col[31] 0.38fF
C16356 a_2475_2154# a_4882_2130# 0.41fF
C16357 a_2275_2154# a_3878_2130# 0.17fF
C16358 a_2275_1150# col[2] 0.16fF
C16359 a_8898_16186# rowon_n[14] 0.14fF
C16360 a_2275_7174# a_27062_7150# 0.71fF
C16361 a_19030_2130# row_n[0] 0.43fF
C16362 a_31078_17190# VDD 1.54fF
C16363 a_26058_12170# a_27062_12170# 0.86fF
C16364 a_18938_6146# rowon_n[4] 0.14fF
C16365 a_2475_11190# col[17] 0.22fF
C16366 a_12306_2170# vcm 0.24fF
C16367 a_2275_16210# a_5886_16186# 0.17fF
C16368 a_2874_11166# vcm 0.18fF
C16369 a_29374_12210# col_n[26] 0.11fF
C16370 a_33998_2130# VDD 0.27fF
C16371 a_2475_4162# a_19942_4138# 0.41fF
C16372 a_2275_4162# a_17326_4178# 0.15fF
C16373 a_10906_4138# a_10998_4138# 0.45fF
C16374 a_2275_17214# col_n[24] 0.17fF
C16375 a_29982_18194# m2_29844_18014# 0.34fF
C16376 a_6982_17190# m2_6752_18014# 0.84fF
C16377 a_2275_6170# col_n[29] 0.17fF
C16378 a_2275_18218# col_n[9] 0.17fF
C16379 a_17022_14178# a_17022_13174# 0.84fF
C16380 a_19942_10162# rowoff_n[8] 0.55fF
C16381 a_27366_6186# vcm 0.24fF
C16382 a_23046_13174# rowoff_n[11] 1.64fF
C16383 a_2275_1150# a_10906_1126# 0.17fF
C16384 a_18026_15182# vcm 0.89fF
C16385 a_2275_14202# col[14] 0.17fF
C16386 a_14922_5142# VDD 0.29fF
C16387 a_1957_18218# vcm 0.16fF
C16388 a_2275_3158# col[19] 0.17fF
C16389 a_2275_6170# a_32386_6186# 0.15fF
C16390 a_2475_6170# a_35002_6146# 0.41fF
C16391 a_23046_10162# col[20] 0.38fF
C16392 a_28978_8154# rowoff_n[6] 0.44fF
C16393 a_3878_14178# VDD 0.29fF
C16394 col_n[17] row_n[2] 0.37fF
C16395 col_n[15] row_n[1] 0.37fF
C16396 col_n[2] col[2] 0.50fF
C16397 col_n[13] row_n[0] 0.37fF
C16398 col_n[30] rowon_n[8] 0.17fF
C16399 col_n[28] rowon_n[7] 0.17fF
C16400 col_n[14] rowon_n[0] 0.17fF
C16401 col_n[21] row_n[4] 0.37fF
C16402 col_n[19] row_n[3] 0.37fF
C16403 col_n[23] row_n[5] 0.37fF
C16404 col_n[16] rowon_n[1] 0.17fF
C16405 VDD col[7] 11.70fF
C16406 col_n[25] row_n[6] 0.37fF
C16407 col_n[18] rowon_n[2] 0.17fF
C16408 col_n[27] row_n[7] 0.37fF
C16409 col_n[20] rowon_n[3] 0.17fF
C16410 col_n[29] row_n[8] 0.37fF
C16411 col_n[22] rowon_n[4] 0.17fF
C16412 vcm col[4] 6.66fF
C16413 col_n[31] row_n[9] 0.37fF
C16414 col_n[24] rowon_n[5] 0.17fF
C16415 col_n[26] rowon_n[6] 0.17fF
C16416 a_6982_15182# a_7986_15182# 0.86fF
C16417 a_2475_15206# a_13006_15182# 0.68fF
C16418 a_8290_9198# vcm 0.24fF
C16419 a_2275_3158# a_25966_3134# 0.17fF
C16420 a_21038_4138# ctop 4.91fF
C16421 a_2275_1150# m2_31852_946# 0.51fF
C16422 a_18330_10202# col_n[15] 0.11fF
C16423 a_17022_9158# row_n[7] 0.43fF
C16424 a_29982_9158# VDD 0.29fF
C16425 a_25966_8154# a_26058_8154# 0.45fF
C16426 a_16930_13174# rowon_n[11] 0.14fF
C16427 a_2275_12194# a_3970_12170# 0.71fF
C16428 a_34394_4178# vcm 0.24fF
C16429 a_26970_3134# rowon_n[1] 0.14fF
C16430 a_2475_17214# a_28066_17190# 0.68fF
C16431 m2_1732_17010# sample 0.31fF
C16432 m2_18800_18014# m2_19804_18014# 0.86fF
C16433 a_23350_13214# vcm 0.24fF
C16434 a_2275_16210# col[31] 0.17fF
C16435 a_10906_12170# VDD 0.29fF
C16436 m2_23820_946# m2_24248_1374# 0.19fF
C16437 a_12002_8154# col[9] 0.38fF
C16438 a_2275_14202# a_19030_14178# 0.71fF
C16439 m2_34864_7974# m2_35292_8402# 0.19fF
C16440 col_n[30] rowoff_n[12] 0.12fF
C16441 a_16930_7150# vcm 0.18fF
C16442 a_3970_7150# rowon_n[5] 0.45fF
C16443 a_2275_13198# col_n[1] 0.17fF
C16444 a_10998_14178# rowoff_n[12] 2.23fF
C16445 a_27062_4138# col_n[24] 0.34fF
C16446 a_2475_2154# a_33086_2130# 0.68fF
C16447 a_17022_2130# a_18026_2130# 0.86fF
C16448 a_2275_2154# col_n[6] 0.17fF
C16449 a_4274_16226# vcm 0.24fF
C16450 a_1957_6170# VDD 0.28fF
C16451 a_17022_11166# ctop 4.91fF
C16452 a_25966_16186# VDD 0.29fF
C16453 a_7286_8194# col_n[4] 0.11fF
C16454 a_2275_11190# a_9294_11206# 0.15fF
C16455 a_2475_11190# a_11910_11166# 0.41fF
C16456 a_6890_11166# a_6982_11166# 0.45fF
C16457 a_2966_6146# col[0] 0.38fF
C16458 a_2275_16210# a_34090_16186# 0.71fF
C16459 a_31990_11166# vcm 0.18fF
C16460 a_15014_16186# row_n[14] 0.43fF
C16461 a_7986_4138# a_7986_3134# 0.84fF
C16462 a_2475_9182# col[11] 0.22fF
C16463 a_17022_17190# m2_17220_17438# 0.19fF
C16464 a_26058_17190# m2_25828_18014# 0.84fF
C16465 a_2161_8178# a_2275_8178# 0.17fF
C16466 a_2475_8178# a_2966_8154# 0.65fF
C16467 a_32082_15182# ctop 4.91fF
C16468 a_25054_6146# row_n[4] 0.43fF
C16469 a_24962_10162# rowon_n[8] 0.14fF
C16470 a_2475_13198# a_26970_13174# 0.41fF
C16471 a_2275_13198# a_24354_13214# 0.15fF
C16472 col_n[14] rowoff_n[13] 0.24fF
C16473 m2_34864_1950# a_34090_2130# 0.86fF
C16474 col[17] rowoff_n[9] 0.23fF
C16475 col[16] rowoff_n[8] 0.24fF
C16476 col[15] rowoff_n[7] 0.25fF
C16477 col[14] rowoff_n[6] 0.25fF
C16478 col[13] rowoff_n[5] 0.26fF
C16479 col[12] rowoff_n[4] 0.27fF
C16480 col[11] rowoff_n[3] 0.27fF
C16481 col[10] rowoff_n[2] 0.28fF
C16482 col[9] rowoff_n[1] 0.29fF
C16483 col[8] rowoff_n[0] 0.29fF
C16484 a_20034_1126# a_20338_1166# 0.10fF
C16485 a_2275_15206# col_n[18] 0.17fF
C16486 a_12914_14178# vcm 0.18fF
C16487 a_8990_4138# VDD 3.82fF
C16488 a_2275_4162# col_n[23] 0.17fF
C16489 a_32082_6146# a_33086_6146# 0.86fF
C16490 a_16018_2130# col_n[13] 0.34fF
C16491 a_26058_14178# col_n[23] 0.34fF
C16492 a_2275_10186# a_17934_10162# 0.17fF
C16493 a_2475_14202# rowon_n[12] 0.40fF
C16494 a_21950_15182# a_22042_15182# 0.45fF
C16495 a_2275_12194# col[8] 0.17fF
C16496 a_6282_18234# col_n[3] 0.11fF
C16497 a_2275_1150# col[13] 0.17fF
C16498 a_12002_4138# rowon_n[2] 0.45fF
C16499 a_27974_18194# vcm 0.18fF
C16500 a_24050_8154# VDD 2.27fF
C16501 a_7986_15182# m2_8184_15430# 0.19fF
C16502 a_23046_8154# a_23046_7150# 0.84fF
C16503 a_2475_7174# a_9994_7150# 0.68fF
C16504 a_2475_11190# col[28] 0.22fF
C16505 sample rowoff_n[14] 0.22fF
C16506 a_2275_12194# a_32994_12170# 0.17fF
C16507 m2_12776_946# col_n[10] 0.45fF
C16508 a_30074_3134# vcm 0.89fF
C16509 col[1] rowoff_n[10] 0.34fF
C16510 a_9994_5142# rowoff_n[3] 2.28fF
C16511 a_27062_11166# m2_27260_11414# 0.19fF
C16512 a_23046_13174# row_n[11] 0.43fF
C16513 a_2275_18218# col_n[20] 0.17fF
C16514 a_4974_11166# VDD 4.23fF
C16515 a_22954_17190# rowon_n[15] 0.14fF
C16516 a_2475_9182# a_25054_9158# 0.68fF
C16517 a_13006_9158# a_14010_9158# 0.86fF
C16518 a_31382_1166# col_n[28] 0.11fF
C16519 m2_1732_15002# rowon_n[13] 0.43fF
C16520 a_15014_12170# col_n[12] 0.34fF
C16521 a_19030_3134# rowoff_n[1] 1.84fF
C16522 a_33086_3134# row_n[1] 0.43fF
C16523 a_10998_6146# vcm 0.89fF
C16524 a_2275_14202# col[25] 0.17fF
C16525 a_32994_7150# rowon_n[5] 0.14fF
C16526 a_2275_3158# col[30] 0.17fF
C16527 a_31990_2130# a_32082_2130# 0.45fF
C16528 a_2275_6170# a_16018_6146# 0.71fF
C16529 col_n[27] rowon_n[1] 0.17fF
C16530 col_n[25] rowon_n[0] 0.17fF
C16531 col_n[30] row_n[3] 0.37fF
C16532 vcm col[15] 6.67fF
C16533 col_n[7] col[8] 6.22fF
C16534 col_n[28] row_n[2] 0.37fF
C16535 col_n[26] row_n[1] 0.37fF
C16536 col_n[24] row_n[0] 0.37fF
C16537 VDD col[18] 8.95fF
C16538 col_n[31] rowon_n[3] 0.17fF
C16539 col_n[29] rowon_n[2] 0.17fF
C16540 col_n[17] en_bit_n[0] 0.19fF
C16541 a_20034_15182# VDD 2.68fF
C16542 a_3970_11166# a_3970_10162# 0.84fF
C16543 m2_4744_18014# vcm 0.71fF
C16544 a_9994_11166# rowon_n[9] 0.45fF
C16545 a_26058_10162# vcm 0.89fF
C16546 a_18026_9158# m2_18224_9406# 0.19fF
C16547 a_2475_3158# a_8898_3134# 0.41fF
C16548 a_2275_3158# a_6282_3174# 0.15fF
C16549 a_2966_4138# ctop 4.82fF
C16550 m3_34996_15134# ctop 0.22fF
C16551 a_2275_8178# a_31078_8154# 0.71fF
C16552 a_28066_13174# a_29070_13174# 0.86fF
C16553 a_16322_4178# vcm 0.24fF
C16554 a_30378_11206# col_n[27] 0.11fF
C16555 a_3970_10162# col_n[1] 0.34fF
C16556 a_11910_11166# rowoff_n[9] 0.64fF
C16557 a_2275_17214# a_9902_17190# 0.17fF
C16558 a_2475_7174# col[5] 0.22fF
C16559 a_6982_13174# vcm 0.89fF
C16560 a_2275_5166# a_21342_5182# 0.15fF
C16561 a_2475_5166# a_23958_5142# 0.41fF
C16562 a_12914_5142# a_13006_5142# 0.45fF
C16563 a_2275_18218# a_19942_18194# 0.17fF
C16564 a_31078_10162# row_n[8] 0.43fF
C16565 a_20946_9158# rowoff_n[7] 0.54fF
C16566 a_2275_13198# col_n[12] 0.17fF
C16567 a_30986_14178# rowon_n[12] 0.14fF
C16568 a_19030_15182# a_19030_14178# 0.84fF
C16569 a_2275_2154# col_n[17] 0.17fF
C16570 a_31382_8194# vcm 0.24fF
C16571 a_27974_15182# rowoff_n[13] 0.46fF
C16572 m2_1732_6970# rowoff_n[5] 2.46fF
C16573 a_8990_7150# m2_9188_7398# 0.19fF
C16574 a_2275_2154# a_14922_2130# 0.17fF
C16575 a_9994_2130# ctop 4.93fF
C16576 a_22042_17190# vcm 0.89fF
C16577 m2_31852_18014# m3_31984_18146# 4.43fF
C16578 a_24050_9158# col[21] 0.38fF
C16579 a_18938_7150# VDD 0.29fF
C16580 a_29982_7150# rowoff_n[5] 0.43fF
C16581 a_2966_7150# a_2966_6146# 0.84fF
C16582 a_2275_10186# col[2] 0.17fF
C16583 a_24962_2130# vcm 0.18fF
C16584 a_2475_16210# a_17022_16186# 0.68fF
C16585 a_8990_16186# a_9994_16186# 0.86fF
C16586 m2_24824_18014# col[22] 0.37fF
C16587 a_28066_3134# m2_28264_3382# 0.19fF
C16588 a_12306_11206# vcm 0.24fF
C16589 a_2475_9182# col[22] 0.22fF
C16590 a_10394_1488# VDD 0.17fF
C16591 a_19334_9198# col_n[16] 0.11fF
C16592 a_18026_8154# rowon_n[6] 0.45fF
C16593 a_2275_4162# a_29982_4138# 0.17fF
C16594 a_25054_6146# ctop 4.91fF
C16595 a_33998_11166# VDD 0.29fF
C16596 m3_24956_1078# m3_25960_1078# 0.21fF
C16597 col_n[25] rowoff_n[13] 0.16fF
C16598 a_2966_17190# m2_1732_17010# 0.86fF
C16599 a_27974_9158# a_28066_9158# 0.45fF
C16600 a_2275_13198# a_7986_13174# 0.71fF
C16601 col[19] rowoff_n[0] 0.22fF
C16602 col[20] rowoff_n[1] 0.21fF
C16603 col[21] rowoff_n[2] 0.21fF
C16604 col[22] rowoff_n[3] 0.20fF
C16605 col[23] rowoff_n[4] 0.19fF
C16606 col[24] rowoff_n[5] 0.19fF
C16607 col[25] rowoff_n[6] 0.18fF
C16608 col[26] rowoff_n[7] 0.17fF
C16609 col[27] rowoff_n[8] 0.17fF
C16610 col[28] rowoff_n[9] 0.16fF
C16611 a_2275_15206# col_n[29] 0.17fF
C16612 a_5886_5142# vcm 0.18fF
C16613 m2_20232_2378# a_20034_2130# 0.19fF
C16614 a_27366_15222# vcm 0.24fF
C16615 a_2475_18218# a_32994_18194# 0.41fF
C16616 a_5978_9158# ctop 4.91fF
C16617 a_29070_17190# row_n[15] 0.43fF
C16618 a_13006_7150# col[10] 0.38fF
C16619 a_14922_14178# VDD 0.29fF
C16620 a_2275_12194# col[19] 0.17fF
C16621 a_5886_2130# rowon_n[0] 0.14fF
C16622 a_2275_1150# col[24] 0.17fF
C16623 a_2275_15206# a_23046_15182# 0.71fF
C16624 a_28066_3134# col_n[25] 0.34fF
C16625 a_20946_9158# vcm 0.18fF
C16626 a_15926_16186# rowoff_n[14] 0.59fF
C16627 a_19030_3134# a_20034_3134# 0.86fF
C16628 a_8290_18234# vcm 0.25fF
C16629 col_n[9] rowoff_n[14] 0.27fF
C16630 a_8290_7190# col_n[5] 0.11fF
C16631 a_21038_13174# ctop 4.91fF
C16632 a_29982_18194# VDD 0.50fF
C16633 col[12] rowoff_n[10] 0.27fF
C16634 a_8898_12170# a_8990_12170# 0.45fF
C16635 a_2275_12194# a_13310_12210# 0.15fF
C16636 a_2475_12194# a_15926_12170# 0.41fF
C16637 a_16018_15182# rowon_n[13] 0.45fF
C16638 m2_29844_18014# m2_30272_18442# 0.19fF
C16639 a_34394_13214# vcm 0.24fF
C16640 a_2275_18218# col_n[31] 0.17fF
C16641 a_32082_3134# VDD 1.44fF
C16642 a_9994_5142# a_9994_4138# 0.84fF
C16643 a_26058_5142# rowon_n[3] 0.45fF
C16644 a_2275_9182# a_6890_9158# 0.17fF
C16645 a_2475_18218# m2_14784_18014# 0.62fF
C16646 a_2275_14202# a_28370_14218# 0.15fF
C16647 a_2475_14202# a_30986_14178# 0.41fF
C16648 a_12002_17190# col[9] 0.38fF
C16649 m2_34864_5966# VDD 1.58fF
C16650 col_n[13] col[13] 0.50fF
C16651 VDD col[29] 6.26fF
C16652 vcm col[26] 6.66fF
C16653 rowon_n[15] ctop 0.37fF
C16654 a_16930_16186# vcm 0.18fF
C16655 a_13006_6146# VDD 3.40fF
C16656 a_3970_5142# row_n[3] 0.43fF
C16657 a_27062_13174# col_n[24] 0.34fF
C16658 a_2275_11190# col_n[6] 0.17fF
C16659 a_1957_15206# VDD 0.28fF
C16660 a_2275_11190# a_21950_11166# 0.17fF
C16661 a_7286_17230# col_n[4] 0.11fF
C16662 a_19030_1126# vcm 0.89fF
C16663 a_2966_15182# col[0] 0.38fF
C16664 a_23958_16186# a_24050_16186# 0.45fF
C16665 m2_8760_18014# VDD 4.61fF
C16666 a_2475_6170# rowoff_n[4] 4.75fF
C16667 a_10998_2130# m2_10768_946# 0.84fF
C16668 a_28066_10162# VDD 1.85fF
C16669 a_25054_9158# a_25054_8154# 0.84fF
C16670 a_2475_8178# a_14010_8154# 0.68fF
C16671 a_2475_7174# col[16] 0.22fF
C16672 a_34090_5142# vcm 0.89fF
C16673 a_28066_12170# rowoff_n[10] 1.40fF
C16674 a_10998_4138# rowoff_n[2] 2.23fF
C16675 a_24050_12170# rowon_n[10] 0.45fF
C16676 a_2275_5166# a_4974_5142# 0.71fF
C16677 a_3878_5142# a_3970_5142# 0.45fF
C16678 a_8990_13174# VDD 3.82fF
C16679 a_2275_13198# col_n[23] 0.17fF
C16680 a_16018_11166# col_n[13] 0.34fF
C16681 a_15014_10162# a_16018_10162# 0.86fF
C16682 a_2475_10186# a_29070_10162# 0.68fF
C16683 a_2275_2154# col_n[28] 0.17fF
C16684 a_34090_2130# rowon_n[0] 0.45fF
C16685 a_20034_2130# rowoff_n[0] 1.79fF
C16686 a_2275_9182# rowoff_n[7] 0.81fF
C16687 a_2475_18218# a_2874_18194# 0.41fF
C16688 a_15014_8154# vcm 0.89fF
C16689 a_2475_12194# row_n[10] 0.48fF
C16690 a_33998_3134# a_34090_3134# 0.45fF
C16691 a_2275_10186# col[13] 0.17fF
C16692 a_19030_1126# m3_18932_1078# 2.16fF
C16693 a_2275_7174# a_20034_7150# 0.71fF
C16694 a_12002_2130# row_n[0] 0.43fF
C16695 a_24050_17190# VDD 2.27fF
C16696 a_5978_12170# a_5978_11166# 0.84fF
C16697 a_11910_6146# rowon_n[4] 0.14fF
C16698 a_5278_2170# vcm 0.24fF
C16699 a_30074_12170# vcm 0.89fF
C16700 a_26970_2130# VDD 0.29fF
C16701 rowon_n[13] rowoff_n[13] 20.66fF
C16702 a_2275_4162# a_10298_4178# 0.15fF
C16703 a_2475_4162# a_12914_4138# 0.41fF
C16704 m3_1864_7102# m3_1864_6098# 0.20fF
C16705 a_2275_9182# a_35094_9158# 0.14fF
C16706 col[30] rowoff_n[0] 0.15fF
C16707 col[31] rowoff_n[1] 0.14fF
C16708 sample_n rowoff_n[2] 0.55fF
C16709 a_30074_14178# a_31078_14178# 0.86fF
C16710 a_12914_10162# rowoff_n[8] 0.63fF
C16711 a_31382_10202# col_n[28] 0.11fF
C16712 a_4974_9158# col_n[2] 0.34fF
C16713 a_20338_6186# vcm 0.24fF
C16714 a_16018_13174# rowoff_n[11] 1.98fF
C16715 a_2874_1126# a_2966_1126# 0.11fF
C16716 a_10998_15182# vcm 0.89fF
C16717 a_7894_5142# VDD 0.29fF
C16718 a_2275_12194# col[30] 0.17fF
C16719 a_2275_6170# a_25358_6186# 0.15fF
C16720 a_2475_6170# a_27974_6146# 0.41fF
C16721 a_14922_6146# a_15014_6146# 0.45fF
C16722 a_32082_9158# rowon_n[7] 0.45fF
C16723 a_21950_8154# rowoff_n[6] 0.52fF
C16724 m2_22816_946# col_n[20] 0.45fF
C16725 a_21038_16186# a_21038_15182# 0.84fF
C16726 a_2475_15206# a_5978_15182# 0.68fF
C16727 a_2275_9182# vcm 7.71fF
C16728 col_n[20] rowoff_n[14] 0.19fF
C16729 a_32082_17190# rowoff_n[15] 1.20fF
C16730 a_25054_8154# col[22] 0.38fF
C16731 a_2275_3158# a_18938_3134# 0.17fF
C16732 a_30986_6146# rowoff_n[4] 0.42fF
C16733 a_14010_4138# ctop 4.91fF
C16734 a_9994_9158# row_n[7] 0.43fF
C16735 m3_16924_1078# ctop 0.21fF
C16736 a_22954_9158# VDD 0.29fF
C16737 col[23] rowoff_n[10] 0.19fF
C16738 a_14010_16186# m2_14208_16434# 0.19fF
C16739 a_9902_13174# rowon_n[11] 0.14fF
C16740 a_2966_13174# ctop 4.82fF
C16741 a_28978_4138# vcm 0.18fF
C16742 m2_1732_3958# row_n[2] 0.44fF
C16743 a_19942_3134# rowon_n[1] 0.14fF
C16744 a_2475_17214# a_21038_17190# 0.68fF
C16745 a_10998_17190# a_12002_17190# 0.86fF
C16746 a_20338_8194# col_n[17] 0.11fF
C16747 m2_11772_18014# m2_12776_18014# 0.86fF
C16748 a_16322_13214# vcm 0.24fF
C16749 a_33086_12170# m2_33284_12418# 0.19fF
C16750 a_2275_5166# a_33998_5142# 0.17fF
C16751 a_2475_16210# col[5] 0.22fF
C16752 a_29070_8154# ctop 4.91fF
C16753 a_2475_5166# col[10] 0.22fF
C16754 a_29982_10162# a_30074_10162# 0.45fF
C16755 m2_1732_11990# sample_n 0.12fF
C16756 a_2275_14202# a_12002_14178# 0.71fF
C16757 col_n[18] col[19] 6.22fF
C16758 rowon_n[4] row_n[4] 21.02fF
C16759 row_n[10] ctop 0.28fF
C16760 col_n[4] rowoff_n[15] 0.31fF
C16761 a_9902_7150# vcm 0.18fF
C16762 a_3970_14178# rowoff_n[12] 2.57fF
C16763 a_2275_11190# col_n[17] 0.17fF
C16764 a_31078_3134# a_31078_2130# 0.84fF
C16765 a_2475_2154# a_26058_2130# 0.68fF
C16766 a_31382_17230# vcm 0.24fF
C16767 col[7] rowoff_n[11] 0.30fF
C16768 a_30074_16186# rowon_n[14] 0.45fF
C16769 a_14010_6146# col[11] 0.38fF
C16770 a_4974_14178# m2_5172_14426# 0.19fF
C16771 a_9994_11166# ctop 4.91fF
C16772 a_18938_16186# VDD 0.29fF
C16773 a_2275_11190# a_3878_11166# 0.17fF
C16774 a_2475_11190# a_4882_11166# 0.41fF
C16775 a_29070_2130# col_n[26] 0.34fF
C16776 a_2275_8178# col[7] 0.17fF
C16777 a_2275_16210# a_27062_16186# 0.71fF
C16778 a_2475_2154# m2_2736_1950# 0.59fF
C16779 a_24962_11166# vcm 0.18fF
C16780 a_21038_1126# VDD 0.11fF
C16781 a_7986_16186# row_n[14] 0.43fF
C16782 a_24050_10162# m2_24248_10410# 0.19fF
C16783 a_21038_4138# a_22042_4138# 0.86fF
C16784 a_9294_6186# col_n[6] 0.11fF
C16785 a_19334_18234# col_n[16] 0.11fF
C16786 a_2475_7174# col[27] 0.22fF
C16787 a_25054_15182# ctop 4.91fF
C16788 a_18026_6146# row_n[4] 0.43fF
C16789 a_2275_13198# a_17326_13214# 0.15fF
C16790 a_10906_13174# a_10998_13174# 0.45fF
C16791 a_2475_13198# a_19942_13174# 0.41fF
C16792 a_17934_10162# rowon_n[8] 0.14fF
C16793 m2_11772_946# vcm 0.71fF
C16794 a_2475_5166# m2_34864_4962# 0.56fF
C16795 a_2275_1150# a_32082_1126# 0.14fF
C16796 a_5886_14178# vcm 0.18fF
C16797 a_2475_4162# VDD 41.96fF
C16798 a_12002_6146# a_12002_5142# 0.84fF
C16799 a_2275_10186# a_10906_10162# 0.17fF
C16800 a_1957_2154# rowoff_n[0] 0.14fF
C16801 a_13006_16186# col[10] 0.38fF
C16802 a_2475_15206# a_35002_15182# 0.41fF
C16803 a_2275_15206# a_32386_15222# 0.15fF
C16804 a_2275_10186# col[24] 0.17fF
C16805 a_15014_8154# m2_15212_8402# 0.19fF
C16806 a_28066_12170# col_n[25] 0.34fF
C16807 a_4974_4138# rowon_n[2] 0.45fF
C16808 a_20946_18194# vcm 0.18fF
C16809 a_17022_8154# VDD 2.99fF
C16810 a_2475_7174# a_2874_7150# 0.41fF
C16811 a_1957_7174# a_2275_7174# 0.19fF
C16812 a_2275_15206# m2_1732_15002# 0.27fF
C16813 a_8290_16226# col_n[5] 0.11fF
C16814 a_2275_12194# a_25966_12170# 0.17fF
C16815 a_23046_3134# vcm 0.89fF
C16816 a_25966_17190# a_26058_17190# 0.45fF
C16817 a_34090_4138# m2_34288_4386# 0.19fF
C16818 a_2874_5142# rowoff_n[3] 0.74fF
C16819 a_16018_13174# row_n[11] 0.43fF
C16820 a_32082_12170# VDD 1.44fF
C16821 m3_20940_18146# m3_21944_18146# 0.21fF
C16822 a_15926_17190# rowon_n[15] 0.14fF
C16823 a_27062_10162# a_27062_9158# 0.84fF
C16824 a_2475_9182# a_18026_9158# 0.68fF
C16825 m2_34864_6970# vcm 0.72fF
C16826 a_12002_3134# rowoff_n[1] 2.18fF
C16827 a_26058_3134# row_n[1] 0.43fF
C16828 a_3970_6146# vcm 0.89fF
C16829 a_25966_7150# rowon_n[5] 0.14fF
C16830 a_32994_14178# rowoff_n[12] 0.40fF
C16831 a_2475_3158# col[4] 0.22fF
C16832 a_5978_6146# m2_6176_6394# 0.19fF
C16833 a_2275_6170# a_8990_6146# 0.71fF
C16834 a_17022_10162# col_n[14] 0.34fF
C16835 a_3878_8154# rowoff_n[6] 0.73fF
C16836 a_13006_15182# VDD 3.40fF
C16837 a_17022_11166# a_18026_11166# 0.86fF
C16838 a_2475_11190# a_33086_11166# 0.68fF
C16839 a_2275_9182# col_n[11] 0.17fF
C16840 col_n[31] rowoff_n[14] 0.11fF
C16841 a_28370_1166# vcm 0.25fF
C16842 a_2874_11166# rowon_n[9] 0.14fF
C16843 a_19030_10162# vcm 0.89fF
C16844 m3_12908_18146# ctop 0.21fF
C16845 a_2275_8178# a_24050_8154# 0.71fF
C16846 a_34090_17190# m2_34864_17010# 0.86fF
C16847 a_2275_6170# col[1] 0.17fF
C16848 a_7986_13174# a_7986_12170# 0.84fF
C16849 a_9294_4178# vcm 0.24fF
C16850 a_4882_11166# rowoff_n[9] 0.72fF
C16851 a_2161_17214# a_2275_17214# 0.17fF
C16852 a_2475_17214# a_2966_17190# 0.65fF
C16853 a_2475_16210# col[16] 0.22fF
C16854 a_34090_14178# vcm 0.89fF
C16855 a_2475_5166# col[21] 0.22fF
C16856 a_30986_4138# VDD 0.29fF
C16857 a_2275_5166# a_14314_5182# 0.15fF
C16858 a_2475_5166# a_16930_5142# 0.41fF
C16859 a_2275_18218# a_12914_18194# 0.17fF
C16860 a_24050_10162# row_n[8] 0.43fF
C16861 rowon_n[4] ctop 0.37fF
C16862 a_32386_9198# col_n[29] 0.11fF
C16863 col_n[24] col[24] 0.50fF
C16864 a_5978_8154# col_n[3] 0.34fF
C16865 col_n[15] rowoff_n[15] 0.23fF
C16866 a_13918_9158# rowoff_n[7] 0.61fF
C16867 a_23958_14178# rowon_n[12] 0.14fF
C16868 a_32082_15182# a_33086_15182# 0.86fF
C16869 a_2275_11190# col_n[28] 0.17fF
C16870 col[18] rowoff_n[11] 0.23fF
C16871 a_24354_8194# vcm 0.24fF
C16872 a_20946_15182# rowoff_n[13] 0.54fF
C16873 m2_1732_8978# VDD 5.46fF
C16874 a_33998_4138# rowon_n[2] 0.14fF
C16875 a_2275_2154# a_7894_2130# 0.17fF
C16876 a_15014_17190# vcm 0.89fF
C16877 a_11910_7150# VDD 0.29fF
C16878 a_22954_7150# rowoff_n[5] 0.51fF
C16879 a_16930_7150# a_17022_7150# 0.45fF
C16880 a_2275_7174# a_29374_7190# 0.15fF
C16881 a_2475_7174# a_31990_7150# 0.41fF
C16882 a_2275_8178# col[18] 0.17fF
C16883 a_17934_2130# vcm 0.18fF
C16884 a_23046_17190# a_23046_16186# 0.84fF
C16885 a_2475_16210# a_9994_16186# 0.68fF
C16886 a_26058_7150# col[23] 0.38fF
C16887 a_31990_5142# rowoff_n[3] 0.41fF
C16888 a_5278_11206# vcm 0.24fF
C16889 a_2966_1126# VDD 0.15fF
C16890 a_10998_8154# rowon_n[6] 0.45fF
C16891 a_2275_4162# a_22954_4138# 0.17fF
C16892 a_18026_6146# ctop 4.91fF
C16893 a_26970_11166# VDD 0.29fF
C16894 m3_10900_1078# m3_11904_1078# 0.21fF
C16895 col[2] rowoff_n[12] 0.33fF
C16896 a_21342_7190# col_n[18] 0.11fF
C16897 a_32994_6146# vcm 0.18fF
C16898 a_20338_15222# vcm 0.24fF
C16899 a_2475_18218# a_25966_18194# 0.41fF
C16900 m2_15788_946# VDD 5.35fF
C16901 a_33086_10162# ctop 4.91fF
C16902 a_22042_17190# row_n[15] 0.43fF
C16903 a_7894_14178# VDD 0.29fF
C16904 a_31990_11166# a_32082_11166# 0.45fF
C16905 a_32082_7150# row_n[5] 0.43fF
C16906 a_2275_15206# a_16018_15182# 0.71fF
C16907 m2_1732_10986# m2_2160_11414# 0.19fF
C16908 a_31990_11166# rowon_n[9] 0.14fF
C16909 a_13918_9158# vcm 0.18fF
C16910 a_8898_16186# rowoff_n[14] 0.67fF
C16911 a_15014_5142# col[12] 0.38fF
C16912 a_33086_4138# a_33086_3134# 0.84fF
C16913 a_2475_3158# a_30074_3134# 0.68fF
C16914 a_25054_17190# col[22] 0.38fF
C16915 a_2275_7174# col_n[5] 0.17fF
C16916 a_14010_13174# ctop 4.91fF
C16917 a_22954_18194# VDD 0.50fF
C16918 m2_3740_18014# col_n[1] 0.33fF
C16919 a_2475_12194# a_8898_12170# 0.41fF
C16920 a_2275_12194# a_6282_12210# 0.15fF
C16921 a_33086_11166# rowoff_n[9] 1.15fF
C16922 a_2275_17214# a_31078_17190# 0.71fF
C16923 a_8990_15182# rowon_n[13] 0.45fF
C16924 m2_22816_18014# m2_23244_18442# 0.19fF
C16925 a_10298_5182# col_n[7] 0.11fF
C16926 a_28978_13174# vcm 0.18fF
C16927 a_25054_3134# VDD 2.16fF
C16928 a_20338_17230# col_n[17] 0.11fF
C16929 a_23046_5142# a_24050_5142# 0.86fF
C16930 a_19030_5142# rowon_n[3] 0.45fF
C16931 a_29070_17190# ctop 4.93fF
C16932 a_2475_14202# col[10] 0.22fF
C16933 a_2475_14202# a_23958_14178# 0.41fF
C16934 a_2275_14202# a_21342_14218# 0.15fF
C16935 a_12914_14178# a_13006_14178# 0.45fF
C16936 a_2475_3158# col[15] 0.22fF
C16937 a_2475_18218# col[1] 0.22fF
C16938 a_9902_16186# vcm 0.18fF
C16939 a_5978_6146# VDD 4.13fF
C16940 a_14010_7150# a_14010_6146# 0.84fF
C16941 a_3970_3134# col[1] 0.38fF
C16942 a_2275_9182# col_n[22] 0.17fF
C16943 a_14010_15182# col[11] 0.38fF
C16944 a_30074_14178# row_n[12] 0.43fF
C16945 a_2275_11190# a_14922_11166# 0.17fF
C16946 a_12002_1126# vcm 0.15fF
C16947 a_2966_16186# a_2966_15182# 0.84fF
C16948 m2_34864_15002# m2_34864_13998# 0.84fF
C16949 a_29070_11166# col_n[26] 0.34fF
C16950 a_2275_17214# col[7] 0.17fF
C16951 a_2275_6170# col[12] 0.17fF
C16952 a_21038_10162# VDD 2.58fF
C16953 a_3970_8154# a_4974_8154# 0.86fF
C16954 a_2475_8178# a_6982_8154# 0.68fF
C16955 a_20034_17190# m2_20232_17438# 0.19fF
C16956 a_9294_15222# col_n[6] 0.11fF
C16957 a_2275_13198# a_29982_13174# 0.17fF
C16958 a_2475_16210# col[27] 0.22fF
C16959 a_27062_5142# vcm 0.89fF
C16960 a_21038_12170# rowoff_n[10] 1.74fF
C16961 a_3970_4138# rowoff_n[2] 2.57fF
C16962 a_27974_18194# a_28066_18194# 0.11fF
C16963 a_2275_18218# m2_31852_18014# 0.51fF
C16964 a_22954_1126# a_23046_1126# 0.11fF
C16965 a_17022_12170# rowon_n[10] 0.45fF
C16966 col_n[29] col[30] 6.16fF
C16967 sw_n ctop 0.60fF
C16968 col_n[26] rowoff_n[15] 0.15fF
C16969 a_2475_13198# VDD 41.96fF
C16970 a_2475_10186# a_22042_10162# 0.68fF
C16971 a_29070_11166# a_29070_10162# 0.84fF
C16972 a_27062_2130# rowon_n[0] 0.45fF
C16973 a_13006_2130# rowoff_n[0] 2.13fF
C16974 col[29] rowoff_n[11] 0.15fF
C16975 a_7986_8154# vcm 0.89fF
C16976 a_2275_15206# rowoff_n[13] 0.81fF
C16977 a_18026_9158# col_n[15] 0.34fF
C16978 a_2275_8178# col[29] 0.17fF
C16979 a_2275_7174# a_13006_7150# 0.71fF
C16980 a_10998_15182# m2_11196_15430# 0.19fF
C16981 m2_1732_5966# rowon_n[4] 0.43fF
C16982 a_17022_17190# VDD 2.99fF
C16983 a_4974_2130# row_n[0] 0.43fF
C16984 a_19030_12170# a_20034_12170# 0.86fF
C16985 a_4882_6146# rowon_n[4] 0.14fF
C16986 a_32386_3174# vcm 0.24fF
C16987 a_2275_5166# col_n[0] 0.17fF
C16988 a_23046_12170# vcm 0.89fF
C16989 a_19942_2130# VDD 0.29fF
C16990 a_2275_4162# a_3270_4178# 0.15fF
C16991 a_2475_4162# a_5886_4138# 0.41fF
C16992 a_30074_11166# m2_30272_11414# 0.19fF
C16993 m3_1864_14130# m3_1864_13126# 0.20fF
C16994 a_2275_9182# a_28066_9158# 0.71fF
C16995 col[13] rowoff_n[12] 0.26fF
C16996 a_9994_14178# a_9994_13174# 0.84fF
C16997 a_5886_10162# rowoff_n[8] 0.70fF
C16998 a_13310_6186# vcm 0.24fF
C16999 a_8990_13174# rowoff_n[11] 2.33fF
C17000 a_3970_15182# vcm 0.89fF
C17001 a_35002_6146# VDD 0.36fF
C17002 a_2475_12194# col[4] 0.22fF
C17003 a_1957_13198# m2_1732_12994# 0.33fF
C17004 a_2275_6170# a_18330_6186# 0.15fF
C17005 a_2475_6170# a_20946_6146# 0.41fF
C17006 a_2475_1150# col[9] 0.22fF
C17007 a_25054_9158# rowon_n[7] 0.45fF
C17008 a_33390_8194# col_n[30] 0.11fF
C17009 a_6982_7150# col_n[4] 0.34fF
C17010 a_14922_8154# rowoff_n[6] 0.60fF
C17011 a_28370_10202# vcm 0.24fF
C17012 a_25054_17190# rowoff_n[15] 1.54fF
C17013 a_3970_1126# en_C0_n 0.28fF
C17014 a_2275_7174# col_n[16] 0.17fF
C17015 a_2275_3158# a_11910_3134# 0.17fF
C17016 a_21038_9158# m2_21236_9406# 0.19fF
C17017 a_23958_6146# rowoff_n[4] 0.50fF
C17018 a_6982_4138# ctop 4.91fF
C17019 a_15926_9158# VDD 0.29fF
C17020 m3_1864_7102# ctop 0.22fF
C17021 a_18938_8154# a_19030_8154# 0.45fF
C17022 a_2275_8178# a_33390_8194# 0.15fF
C17023 a_2275_15206# col[1] 0.17fF
C17024 a_27062_6146# col[24] 0.38fF
C17025 a_2275_4162# col[6] 0.17fF
C17026 a_21950_4138# vcm 0.18fF
C17027 a_12914_3134# rowon_n[1] 0.14fF
C17028 a_32994_4138# rowoff_n[2] 0.40fF
C17029 a_2475_17214# a_14010_17190# 0.68fF
C17030 m2_4744_18014# m2_5748_18014# 0.86fF
C17031 a_9294_13214# vcm 0.24fF
C17032 a_2275_5166# a_26970_5142# 0.17fF
C17033 a_22042_8154# ctop 4.91fF
C17034 a_2475_14202# col[21] 0.22fF
C17035 a_30986_13174# VDD 0.29fF
C17036 m2_6752_946# col_n[4] 0.45fF
C17037 a_2475_3158# col[26] 0.22fF
C17038 a_22346_6186# col_n[19] 0.11fF
C17039 m2_1732_9982# vcm 1.11fF
C17040 a_2475_18218# col[12] 0.22fF
C17041 a_2275_14202# a_4974_14178# 0.71fF
C17042 a_3878_14178# a_3970_14178# 0.45fF
C17043 a_32386_18234# col_n[29] 0.11fF
C17044 a_5978_17190# col_n[3] 0.34fF
C17045 a_2475_2154# a_19030_2130# 0.68fF
C17046 a_12002_7150# m2_12200_7398# 0.19fF
C17047 a_9994_2130# a_10998_2130# 0.86fF
C17048 a_24354_17230# vcm 0.24fF
C17049 a_23046_16186# rowon_n[14] 0.45fF
C17050 a_11910_16186# VDD 0.29fF
C17051 a_33998_12170# a_34090_12170# 0.45fF
C17052 a_33086_6146# rowon_n[4] 0.45fF
C17053 a_2275_17214# col[18] 0.17fF
C17054 a_2275_16210# a_20034_16186# 0.71fF
C17055 a_2275_6170# col[23] 0.17fF
C17056 a_31078_3134# m2_31276_3382# 0.19fF
C17057 a_16018_4138# col[13] 0.38fF
C17058 a_17934_11166# vcm 0.18fF
C17059 a_2275_18218# col[3] 0.17fF
C17060 a_14010_1126# VDD 0.13fF
C17061 a_26058_16186# col[23] 0.38fF
C17062 a_2475_4162# a_34090_4138# 0.68fF
C17063 a_2966_10162# VDD 4.45fF
C17064 a_18026_15182# ctop 4.91fF
C17065 a_10998_6146# row_n[4] 0.43fF
C17066 a_10906_10162# rowon_n[8] 0.14fF
C17067 a_2275_13198# a_10298_13214# 0.15fF
C17068 a_2475_13198# a_12914_13174# 0.41fF
C17069 a_34090_10162# rowoff_n[8] 1.10fF
C17070 a_2966_12170# rowoff_n[10] 2.62fF
C17071 a_11302_4178# col_n[8] 0.11fF
C17072 m2_23244_2378# a_23046_2130# 0.19fF
C17073 ctop col[4] 0.13fF
C17074 rowon_n[12] sample_n 0.15fF
C17075 a_21342_16226# col_n[18] 0.11fF
C17076 a_2275_1150# a_25054_1126# 0.14fF
C17077 a_32994_15182# vcm 0.18fF
C17078 a_29070_5142# VDD 1.75fF
C17079 a_25054_6146# a_26058_6146# 0.86fF
C17080 a_2874_10162# a_2966_10162# 0.45fF
C17081 a_2475_15206# a_27974_15182# 0.41fF
C17082 a_2275_15206# a_25358_15222# 0.15fF
C17083 a_14922_15182# a_15014_15182# 0.45fF
C17084 a_13918_18194# vcm 0.18fF
C17085 a_4974_2130# col[2] 0.38fF
C17086 a_9994_8154# VDD 3.71fF
C17087 a_16018_8154# a_16018_7150# 0.84fF
C17088 a_15014_14178# col[12] 0.38fF
C17089 a_31078_13174# rowon_n[11] 0.45fF
C17090 a_2275_16210# col_n[5] 0.17fF
C17091 a_2275_12194# a_18938_12170# 0.17fF
C17092 a_2275_5166# col_n[10] 0.17fF
C17093 a_16018_3134# vcm 0.89fF
C17094 a_30074_10162# col_n[27] 0.34fF
C17095 a_35398_3174# VDD 0.12fF
C17096 col[24] rowoff_n[12] 0.19fF
C17097 a_10298_14218# col_n[7] 0.11fF
C17098 a_8990_13174# row_n[11] 0.43fF
C17099 a_25054_12170# VDD 2.16fF
C17100 m3_6884_18146# m3_7888_18146# 0.21fF
C17101 m2_4744_946# m3_4876_1078# 4.41fF
C17102 a_5978_9158# a_6982_9158# 0.86fF
C17103 a_2275_2154# col[0] 0.16fF
C17104 a_2475_9182# a_10998_9158# 0.68fF
C17105 a_8898_17190# rowon_n[15] 0.14fF
C17106 m2_18800_18014# col[16] 0.39fF
C17107 a_2275_14202# a_33998_14178# 0.17fF
C17108 a_19030_3134# row_n[1] 0.43fF
C17109 a_4974_3134# rowoff_n[1] 2.52fF
C17110 a_18938_7150# rowon_n[5] 0.14fF
C17111 a_31078_7150# vcm 0.89fF
C17112 a_25966_14178# rowoff_n[12] 0.48fF
C17113 a_2475_12194# col[15] 0.22fF
C17114 a_24962_2130# a_25054_2130# 0.45fF
C17115 a_2475_1150# col[20] 0.22fF
C17116 a_2475_6170# a_2275_6170# 2.96fF
C17117 a_1957_6170# a_2161_6170# 0.11fF
C17118 a_5978_15182# VDD 4.13fF
C17119 a_2475_11190# a_26058_11166# 0.68fF
C17120 a_31078_12170# a_31078_11166# 0.84fF
C17121 a_3970_12170# col[1] 0.38fF
C17122 a_21342_1166# vcm 0.25fF
C17123 a_2275_7174# col_n[27] 0.17fF
C17124 a_12002_10162# vcm 0.89fF
C17125 a_19030_8154# col_n[16] 0.34fF
C17126 col[8] rowoff_n[13] 0.29fF
C17127 a_2275_15206# col[12] 0.17fF
C17128 a_2275_8178# a_17022_8154# 0.71fF
C17129 a_2275_4162# col[17] 0.17fF
C17130 a_21038_13174# a_22042_13174# 0.86fF
C17131 a_3878_4138# vcm 0.18fF
C17132 a_27062_14178# vcm 0.89fF
C17133 a_23958_4138# VDD 0.29fF
C17134 a_5886_5142# a_5978_5142# 0.45fF
C17135 a_2275_5166# a_7286_5182# 0.15fF
C17136 a_2475_5166# a_9902_5142# 0.41fF
C17137 a_2275_18218# a_5886_18194# 0.17fF
C17138 a_2475_18218# col[23] 0.22fF
C17139 a_2275_10186# a_32082_10162# 0.71fF
C17140 a_17022_10162# row_n[8] 0.43fF
C17141 a_6890_9158# rowoff_n[7] 0.69fF
C17142 a_16930_14178# rowon_n[12] 0.14fF
C17143 a_12002_15182# a_12002_14178# 0.84fF
C17144 a_17326_8194# vcm 0.24fF
C17145 a_13918_15182# rowoff_n[13] 0.61fF
C17146 a_26970_4138# rowon_n[2] 0.14fF
C17147 a_7986_17190# vcm 0.89fF
C17148 a_30074_3134# ctop 4.91fF
C17149 a_4882_7150# VDD 0.29fF
C17150 a_15926_7150# rowoff_n[5] 0.59fF
C17151 a_7986_6146# col_n[5] 0.34fF
C17152 a_2475_7174# a_24962_7150# 0.41fF
C17153 a_2275_7174# a_22346_7190# 0.15fF
C17154 a_2275_17214# col[29] 0.17fF
C17155 a_2275_18218# col[14] 0.17fF
C17156 a_10906_2130# vcm 0.18fF
C17157 a_2475_16210# a_2874_16186# 0.41fF
C17158 a_1957_16210# a_2275_16210# 0.19fF
C17159 a_24962_5142# rowoff_n[3] 0.49fF
C17160 a_32386_12210# vcm 0.24fF
C17161 a_3970_8154# rowon_n[6] 0.45fF
C17162 a_2275_4162# a_15926_4138# 0.17fF
C17163 a_2275_14202# col_n[0] 0.17fF
C17164 a_10998_6146# ctop 4.91fF
C17165 a_2275_3158# col_n[4] 0.17fF
C17166 a_19942_11166# VDD 0.29fF
C17167 a_20946_9158# a_21038_9158# 0.45fF
C17168 a_28066_5142# col[25] 0.38fF
C17169 a_33998_3134# rowoff_n[1] 0.39fF
C17170 row_n[7] sample_n 0.16fF
C17171 ctop col[15] 0.13fF
C17172 a_25966_6146# vcm 0.18fF
C17173 a_13310_15222# vcm 0.24fF
C17174 a_2475_18218# a_18938_18194# 0.41fF
C17175 a_2275_6170# a_30986_6146# 0.17fF
C17176 a_15014_17190# row_n[15] 0.43fF
C17177 a_26058_10162# ctop 4.91fF
C17178 a_35002_15182# VDD 0.36fF
C17179 a_23350_5182# col_n[20] 0.11fF
C17180 a_2475_10186# col[9] 0.22fF
C17181 a_33390_17230# col_n[30] 0.11fF
C17182 a_6982_16186# col_n[4] 0.34fF
C17183 m2_33860_18014# vcm 0.71fF
C17184 a_25054_7150# row_n[5] 0.43fF
C17185 a_2275_15206# a_8990_15182# 0.71fF
C17186 a_24962_11166# rowon_n[9] 0.14fF
C17187 a_6890_9158# vcm 0.18fF
C17188 a_12002_3134# a_13006_3134# 0.86fF
C17189 a_2475_3158# a_23046_3134# 0.68fF
C17190 a_2475_1150# m2_26832_946# 0.62fF
C17191 a_33086_2130# m2_32856_946# 0.84fF
C17192 m3_31984_1078# ctop 0.21fF
C17193 a_2275_16210# col_n[16] 0.17fF
C17194 a_17022_16186# m2_17220_16434# 0.19fF
C17195 a_2275_5166# col_n[21] 0.17fF
C17196 a_6982_13174# ctop 4.91fF
C17197 a_15926_18194# VDD 0.50fF
C17198 m2_1732_946# m2_2160_1374# 0.19fF
C17199 a_26058_11166# rowoff_n[9] 1.50fF
C17200 a_17022_3134# col[14] 0.38fF
C17201 a_2275_17214# a_24050_17190# 0.71fF
C17202 a_2475_15206# rowon_n[13] 0.40fF
C17203 a_27062_15182# col[24] 0.38fF
C17204 m2_15788_18014# m2_16216_18442# 0.19fF
C17205 a_21950_13174# vcm 0.18fF
C17206 a_2275_13198# col[6] 0.17fF
C17207 a_18026_3134# VDD 2.89fF
C17208 a_2275_2154# col[11] 0.17fF
C17209 a_12002_5142# rowon_n[3] 0.45fF
C17210 a_2275_18218# a_34090_18194# 0.14fF
C17211 a_22042_17190# ctop 4.93fF
C17212 a_2475_12194# col[26] 0.22fF
C17213 a_2475_14202# a_16930_14178# 0.41fF
C17214 a_2275_14202# a_14314_14218# 0.15fF
C17215 a_12306_3174# col_n[9] 0.11fF
C17216 a_22346_15222# col_n[19] 0.11fF
C17217 a_2275_2154# a_29070_2130# 0.71fF
C17218 a_33086_7150# VDD 1.34fF
C17219 a_7986_14178# m2_8184_14426# 0.19fF
C17220 a_27062_7150# a_28066_7150# 0.86fF
C17221 a_23046_14178# row_n[12] 0.43fF
C17222 a_2275_11190# a_7894_11166# 0.17fF
C17223 a_4974_1126# vcm 0.15fF
C17224 col[19] rowoff_n[13] 0.22fF
C17225 a_16930_16186# a_17022_16186# 0.45fF
C17226 a_2475_16210# a_31990_16186# 0.41fF
C17227 a_2275_16210# a_29374_16226# 0.15fF
C17228 a_4974_2130# m2_5172_2378# 0.19fF
C17229 a_33086_4138# row_n[2] 0.43fF
C17230 col_n[0] rowoff_n[6] 0.34fF
C17231 vcm rowoff_n[7] 2.43fF
C17232 VDD rowoff_n[4] 87.22fF
C17233 sample rowoff_n[5] 0.22fF
C17234 col_n[2] rowoff_n[9] 0.32fF
C17235 col_n[1] rowoff_n[8] 0.33fF
C17236 a_32994_8154# rowon_n[6] 0.14fF
C17237 a_2275_15206# col[23] 0.17fF
C17238 a_27062_10162# m2_27260_10410# 0.19fF
C17239 a_16018_13174# col[13] 0.38fF
C17240 a_2275_4162# col[28] 0.17fF
C17241 a_14010_10162# VDD 3.30fF
C17242 a_18026_9158# a_18026_8154# 0.84fF
C17243 a_2275_13198# a_22954_13174# 0.17fF
C17244 a_31078_9158# col_n[28] 0.34fF
C17245 a_20034_5142# vcm 0.89fF
C17246 a_14010_12170# rowoff_n[10] 2.08fF
C17247 a_2275_18218# m2_17796_18014# 0.51fF
C17248 m2_20808_946# vcm 0.71fF
C17249 a_11302_13214# col_n[8] 0.11fF
C17250 a_9994_12170# rowon_n[10] 0.45fF
C17251 a_29070_14178# VDD 1.75fF
C17252 a_2475_10186# a_15014_10162# 0.68fF
C17253 a_7986_10162# a_8990_10162# 0.86fF
C17254 a_5978_2130# rowoff_n[0] 2.47fF
C17255 a_20034_2130# rowon_n[0] 0.45fF
C17256 col[3] rowoff_n[14] 0.33fF
C17257 a_35094_9158# vcm 0.15fF
C17258 a_30074_16186# rowoff_n[14] 1.30fF
C17259 a_26970_3134# a_27062_3134# 0.45fF
C17260 a_18026_8154# m2_18224_8402# 0.19fF
C17261 a_2475_8178# col[3] 0.22fF
C17262 a_2275_7174# a_5978_7150# 0.71fF
C17263 a_4974_11166# col[2] 0.38fF
C17264 a_2275_18218# col[25] 0.17fF
C17265 a_9994_17190# VDD 3.72fF
C17266 a_2475_12194# a_30074_12170# 0.68fF
C17267 a_33086_13174# a_33086_12170# 0.84fF
C17268 a_25358_3174# vcm 0.24fF
C17269 a_31078_11166# row_n[9] 0.43fF
C17270 a_30986_15182# rowon_n[13] 0.14fF
C17271 a_20034_7150# col_n[17] 0.34fF
C17272 a_2275_14202# col_n[10] 0.17fF
C17273 a_16018_12170# vcm 0.89fF
C17274 a_2275_3158# col_n[15] 0.17fF
C17275 a_12914_2130# VDD 0.29fF
C17276 a_35398_12210# VDD 0.12fF
C17277 VDD col_n[3] 15.69fF
C17278 a_15926_18194# m2_15788_18014# 0.34fF
C17279 a_2275_9182# a_21038_9158# 0.71fF
C17280 ctop col[26] 0.13fF
C17281 rowon_n[1] sample_n 0.15fF
C17282 a_2275_11190# col[0] 0.16fF
C17283 a_23046_14178# a_24050_14178# 0.86fF
C17284 a_6282_6186# vcm 0.24fF
C17285 a_2475_13198# rowoff_n[11] 4.75fF
C17286 a_8990_6146# m2_9188_6394# 0.19fF
C17287 a_19030_1126# ctop 2.45fF
C17288 a_31078_16186# vcm 0.89fF
C17289 a_27974_6146# VDD 0.29fF
C17290 a_7894_6146# a_7986_6146# 0.45fF
C17291 a_2475_6170# a_13918_6146# 0.41fF
C17292 a_2275_6170# a_11302_6186# 0.15fF
C17293 a_2475_10186# col[20] 0.22fF
C17294 a_18026_9158# rowon_n[7] 0.45fF
C17295 a_7894_8154# rowoff_n[6] 0.68fF
C17296 a_35002_1126# vcm 0.17fF
C17297 a_14010_16186# a_14010_15182# 0.84fF
C17298 a_21342_10202# vcm 0.24fF
C17299 a_18026_17190# rowoff_n[15] 1.89fF
C17300 a_2275_16210# col_n[27] 0.17fF
C17301 a_8990_5142# col_n[6] 0.34fF
C17302 a_2966_3134# a_3970_3134# 0.86fF
C17303 a_2275_3158# a_4882_3134# 0.17fF
C17304 a_16930_6146# rowoff_n[4] 0.58fF
C17305 a_34090_5142# ctop 4.80fF
C17306 a_8898_9158# VDD 0.29fF
C17307 m3_27968_18146# ctop 0.21fF
C17308 a_19030_17190# col_n[16] 0.34fF
C17309 a_2475_8178# a_28978_8154# 0.41fF
C17310 a_2275_8178# a_26362_8194# 0.15fF
C17311 a_2966_16186# m2_1732_16006# 0.86fF
C17312 a_2275_13198# col[17] 0.17fF
C17313 a_14922_4138# vcm 0.18fF
C17314 a_5886_3134# rowon_n[1] 0.14fF
C17315 a_25966_4138# rowoff_n[2] 0.48fF
C17316 a_3970_17190# a_4974_17190# 0.86fF
C17317 a_2475_17214# a_6982_17190# 0.68fF
C17318 a_2275_2154# col[22] 0.17fF
C17319 a_3878_13174# vcm 0.18fF
C17320 a_2275_5166# a_19942_5142# 0.17fF
C17321 a_15014_8154# ctop 4.91fF
C17322 a_23958_13174# VDD 0.29fF
C17323 a_29070_4138# col[26] 0.38fF
C17324 a_22954_10162# a_23046_10162# 0.45fF
C17325 a_35002_2130# rowoff_n[0] 0.38fF
C17326 a_29982_8154# vcm 0.18fF
C17327 a_24050_3134# a_24050_2130# 0.84fF
C17328 a_2475_2154# a_12002_2130# 0.68fF
C17329 a_17326_17230# vcm 0.24fF
C17330 a_16018_16186# rowon_n[14] 0.45fF
C17331 a_2275_7174# a_35002_7150# 0.17fF
C17332 a_24354_4178# col_n[21] 0.11fF
C17333 a_30074_12170# ctop 4.91fF
C17334 a_4882_16186# VDD 0.29fF
C17335 col[30] rowoff_n[13] 0.15fF
C17336 a_7986_15182# col_n[5] 0.34fF
C17337 a_26058_6146# rowon_n[4] 0.45fF
C17338 col_n[13] rowoff_n[9] 0.24fF
C17339 col_n[6] rowoff_n[2] 0.29fF
C17340 col_n[9] rowoff_n[5] 0.27fF
C17341 col_n[12] rowoff_n[8] 0.25fF
C17342 col_n[7] rowoff_n[3] 0.29fF
C17343 col_n[10] rowoff_n[6] 0.27fF
C17344 col_n[4] rowoff_n[0] 0.31fF
C17345 col_n[11] rowoff_n[7] 0.26fF
C17346 col_n[8] rowoff_n[4] 0.28fF
C17347 col_n[5] rowoff_n[1] 0.30fF
C17348 a_2275_16210# a_13006_16186# 0.71fF
C17349 a_10906_11166# vcm 0.18fF
C17350 a_6982_1126# VDD 0.14fF
C17351 a_14010_4138# a_15014_4138# 0.86fF
C17352 a_2475_4162# a_27062_4138# 0.68fF
C17353 a_35002_18194# m2_34864_18014# 0.33fF
C17354 a_12002_17190# m2_11772_18014# 0.84fF
C17355 a_10998_15182# ctop 4.91fF
C17356 a_3970_6146# row_n[4] 0.43fF
C17357 a_2275_12194# col_n[4] 0.17fF
C17358 a_2275_13198# a_3270_13214# 0.15fF
C17359 a_2475_13198# a_5886_13174# 0.41fF
C17360 a_18026_2130# col[15] 0.38fF
C17361 a_2275_1150# col_n[9] 0.17fF
C17362 a_27062_10162# rowoff_n[8] 1.45fF
C17363 a_1957_5166# vcm 0.16fF
C17364 a_28066_14178# col[25] 0.38fF
C17365 a_30986_13174# rowoff_n[11] 0.42fF
C17366 a_2275_1150# a_18026_1126# 0.79fF
C17367 a_25966_15182# vcm 0.18fF
C17368 a_22042_5142# VDD 2.47fF
C17369 m2_24824_946# VDD 4.00fF
C17370 a_4974_6146# a_4974_5142# 0.84fF
C17371 a_2275_9182# ctop 0.14fF
C17372 col[14] rowoff_n[14] 0.25fF
C17373 a_13310_2170# col_n[10] 0.11fF
C17374 VDD rowoff_n[10] 87.22fF
C17375 a_23350_14218# col_n[20] 0.11fF
C17376 a_2275_15206# a_18330_15222# 0.15fF
C17377 a_2475_15206# a_20946_15182# 0.41fF
C17378 a_2475_8178# col[14] 0.22fF
C17379 a_2275_3158# a_33086_3134# 0.71fF
C17380 a_6890_18194# vcm 0.18fF
C17381 a_2874_8154# VDD 0.29fF
C17382 a_29070_8154# a_30074_8154# 0.86fF
C17383 a_24050_13174# rowon_n[11] 0.45fF
C17384 a_2275_12194# a_11910_12170# 0.17fF
C17385 a_2275_14202# col_n[21] 0.17fF
C17386 a_8990_3134# vcm 0.89fF
C17387 a_2275_3158# col_n[26] 0.17fF
C17388 a_34090_3134# rowon_n[1] 0.45fF
C17389 a_18938_17190# a_19030_17190# 0.45fF
C17390 a_2275_17214# a_33390_17230# 0.15fF
C17391 m2_2736_1950# m3_2868_2082# 4.41fF
C17392 a_17022_12170# col[14] 0.38fF
C17393 VDD col_n[14] 12.96fF
C17394 vcm col_n[11] 3.22fF
C17395 a_2475_13198# row_n[11] 0.48fF
C17396 a_18026_12170# VDD 2.89fF
C17397 a_2275_11190# col[11] 0.17fF
C17398 a_3878_18194# m2_3740_18014# 0.34fF
C17399 a_2275_9182# a_2966_9158# 0.67fF
C17400 a_2475_9182# a_3970_9158# 0.68fF
C17401 a_20034_10162# a_20034_9158# 0.84fF
C17402 a_32082_8154# col_n[29] 0.34fF
C17403 a_2275_14202# a_26970_14178# 0.17fF
C17404 a_12002_3134# row_n[1] 0.43fF
C17405 a_11910_7150# rowon_n[5] 0.14fF
C17406 a_24050_7150# vcm 0.89fF
C17407 a_18938_14178# rowoff_n[12] 0.56fF
C17408 a_12306_12210# col_n[9] 0.11fF
C17409 a_2475_10186# col[31] 0.22fF
C17410 a_33086_16186# VDD 1.34fF
C17411 a_2475_11190# a_19030_11166# 0.68fF
C17412 a_9994_11166# a_10998_11166# 0.86fF
C17413 a_14314_1166# vcm 0.25fF
C17414 a_4974_10162# vcm 0.89fF
C17415 a_28978_4138# a_29070_4138# 0.45fF
C17416 a_5978_10162# col[3] 0.38fF
C17417 a_31078_17190# m2_30848_18014# 0.84fF
C17418 a_23046_17190# m2_23244_17438# 0.19fF
C17419 a_2275_8178# a_9994_8154# 0.71fF
C17420 a_2275_13198# col[28] 0.17fF
C17421 a_32082_10162# rowon_n[8] 0.45fF
C17422 a_2475_13198# a_34090_13174# 0.68fF
C17423 a_21038_6146# col_n[18] 0.34fF
C17424 a_29374_5182# vcm 0.24fF
C17425 a_20034_14178# vcm 0.89fF
C17426 a_16930_4138# VDD 0.29fF
C17427 m2_31852_946# col[29] 0.52fF
C17428 a_2275_10186# a_25054_10162# 0.71fF
C17429 a_9994_10162# row_n[8] 0.43fF
C17430 a_9902_14178# rowon_n[12] 0.14fF
C17431 a_25054_15182# a_26058_15182# 0.86fF
C17432 a_10298_8194# vcm 0.24fF
C17433 a_6890_15182# rowoff_n[13] 0.69fF
C17434 a_19942_4138# rowon_n[2] 0.14fF
C17435 a_23046_3134# ctop 4.91fF
C17436 a_35094_18194# vcm 0.15fF
C17437 m2_3740_18014# m3_3872_18146# 4.42fF
C17438 a_31990_8154# VDD 0.29fF
C17439 a_8898_7150# rowoff_n[5] 0.67fF
C17440 a_14010_15182# m2_14208_15430# 0.19fF
C17441 a_2475_7174# a_17934_7150# 0.41fF
C17442 a_2275_7174# a_15318_7190# 0.15fF
C17443 a_9902_7150# a_9994_7150# 0.45fF
C17444 a_2475_17214# col[3] 0.22fF
C17445 col_n[15] rowoff_n[0] 0.23fF
C17446 col_n[18] rowoff_n[3] 0.21fF
C17447 col_n[21] rowoff_n[6] 0.19fF
C17448 col_n[24] rowoff_n[9] 0.16fF
C17449 col_n[17] rowoff_n[2] 0.21fF
C17450 col_n[22] rowoff_n[7] 0.18fF
C17451 col_n[19] rowoff_n[4] 0.20fF
C17452 col_n[16] rowoff_n[1] 0.22fF
C17453 col_n[23] rowoff_n[8] 0.17fF
C17454 col_n[20] rowoff_n[5] 0.19fF
C17455 a_2475_6170# col[8] 0.22fF
C17456 a_16018_17190# a_16018_16186# 0.84fF
C17457 m2_1732_12994# sample 0.31fF
C17458 a_25358_12210# vcm 0.24fF
C17459 a_9994_4138# col_n[7] 0.34fF
C17460 a_17934_5142# rowoff_n[3] 0.57fF
C17461 a_20034_16186# col_n[17] 0.34fF
C17462 a_33086_11166# m2_33284_11414# 0.19fF
C17463 a_2275_4162# a_8898_4138# 0.17fF
C17464 a_3970_6146# ctop 4.91fF
C17465 a_2275_12194# col_n[15] 0.17fF
C17466 a_12914_11166# VDD 0.29fF
C17467 a_2275_1150# col_n[20] 0.17fF
C17468 a_2475_9182# a_32994_9158# 0.41fF
C17469 a_2275_9182# a_30378_9198# 0.15fF
C17470 a_30074_17190# rowon_n[15] 0.45fF
C17471 a_26970_3134# rowoff_n[1] 0.47fF
C17472 m2_34864_5966# m2_35292_6394# 0.19fF
C17473 a_18938_6146# vcm 0.18fF
C17474 a_2275_9182# col[5] 0.17fF
C17475 a_6282_15222# vcm 0.24fF
C17476 col[25] rowoff_n[14] 0.18fF
C17477 a_2475_18218# a_11910_18194# 0.41fF
C17478 a_34394_5182# col_n[31] 0.11fF
C17479 a_4974_13174# m2_5172_13422# 0.19fF
C17480 a_2275_6170# a_23958_6146# 0.17fF
C17481 a_30074_3134# col[27] 0.38fF
C17482 a_19030_10162# ctop 4.91fF
C17483 a_7986_17190# row_n[15] 0.43fF
C17484 col_n[8] rowoff_n[10] 0.28fF
C17485 a_27974_15182# VDD 0.29fF
C17486 a_24962_11166# a_25054_11166# 0.45fF
C17487 m2_19804_18014# vcm 0.71fF
C17488 a_2475_8178# col[25] 0.22fF
C17489 a_18026_7150# row_n[5] 0.43fF
C17490 a_2475_15206# a_2275_15206# 2.96fF
C17491 a_1957_15206# a_2161_15206# 0.11fF
C17492 a_17934_11166# rowon_n[9] 0.14fF
C17493 a_33998_10162# vcm 0.18fF
C17494 a_24050_9158# m2_24248_9406# 0.19fF
C17495 a_2475_3158# a_16018_3134# 0.68fF
C17496 a_26058_4138# a_26058_3134# 0.84fF
C17497 a_2275_1150# m2_9764_946# 0.51fF
C17498 a_25358_3174# col_n[22] 0.11fF
C17499 m3_3872_1078# ctop 0.33fF
C17500 a_8990_14178# col_n[6] 0.34fF
C17501 a_34090_14178# ctop 4.80fF
C17502 a_8898_18194# VDD 0.50fF
C17503 a_19030_11166# rowoff_n[9] 1.84fF
C17504 a_2275_17214# a_17022_17190# 0.71fF
C17505 VDD col_n[25] 10.24fF
C17506 vcm col_n[22] 3.22fF
C17507 col[9] rowoff_n[15] 0.29fF
C17508 m2_8760_18014# m2_9188_18442# 0.19fF
C17509 a_2475_4162# m2_34864_3958# 0.56fF
C17510 a_14922_13174# vcm 0.18fF
C17511 a_10998_3134# VDD 3.61fF
C17512 a_2275_11190# col[22] 0.17fF
C17513 a_2475_5166# a_31078_5142# 0.68fF
C17514 a_16018_5142# a_17022_5142# 0.86fF
C17515 a_4974_5142# rowon_n[3] 0.45fF
C17516 a_2275_18218# a_27062_18194# 0.14fF
C17517 m2_11772_946# m2_12776_946# 0.86fF
C17518 a_15014_17190# ctop 4.93fF
C17519 a_28066_9158# rowoff_n[7] 1.40fF
C17520 a_19030_1126# col[16] 0.53fF
C17521 a_29070_13174# col[26] 0.38fF
C17522 a_2475_14202# a_9902_14178# 0.41fF
C17523 a_2275_14202# a_7286_14218# 0.15fF
C17524 a_5886_14178# a_5978_14178# 0.45fF
C17525 a_15014_7150# m2_15212_7398# 0.19fF
C17526 a_2275_2154# a_22042_2130# 0.71fF
C17527 a_29982_17190# vcm 0.18fF
C17528 a_26058_7150# VDD 2.06fF
C17529 a_2275_14202# m2_1732_13998# 0.27fF
C17530 a_6982_7150# a_6982_6146# 0.84fF
C17531 a_14314_1166# col_n[11] 0.11fF
C17532 a_16018_14178# row_n[12] 0.43fF
C17533 a_24354_13214# col_n[21] 0.11fF
C17534 a_32082_2130# vcm 0.89fF
C17535 a_2475_16210# a_24962_16186# 0.41fF
C17536 a_2275_16210# a_22346_16226# 0.15fF
C17537 a_34090_3134# m2_34288_3382# 0.19fF
C17538 a_26058_4138# row_n[2] 0.43fF
C17539 a_25966_8154# rowon_n[6] 0.14fF
C17540 a_2475_4162# col[2] 0.22fF
C17541 a_6982_10162# VDD 4.02fF
C17542 a_31078_9158# a_32082_9158# 0.86fF
C17543 a_2275_13198# a_15926_13174# 0.17fF
C17544 a_13006_5142# vcm 0.89fF
C17545 a_6982_12170# rowoff_n[10] 2.42fF
C17546 m2_26256_2378# a_26058_2130# 0.19fF
C17547 a_20946_18194# a_21038_18194# 0.11fF
C17548 a_18026_11166# col[15] 0.38fF
C17549 a_2275_10186# col_n[9] 0.17fF
C17550 a_2275_18218# m2_3740_18014# 0.51fF
C17551 a_15926_1126# a_16018_1126# 0.11fF
C17552 a_2275_1150# a_27366_1166# 0.15fF
C17553 a_2475_1150# a_29982_1126# 0.41fF
C17554 a_5978_5142# m2_6176_5390# 0.19fF
C17555 a_1957_14202# vcm 0.16fF
C17556 a_2874_12170# rowon_n[10] 0.14fF
C17557 m3_22948_18146# VDD 0.11fF
C17558 a_33086_7150# col_n[30] 0.34fF
C17559 a_22042_14178# VDD 2.47fF
C17560 a_2475_10186# a_7986_10162# 0.68fF
C17561 a_22042_11166# a_22042_10162# 0.84fF
C17562 a_13006_2130# rowon_n[0] 0.45fF
C17563 a_2275_15206# a_30986_15182# 0.17fF
C17564 a_13310_11206# col_n[10] 0.11fF
C17565 a_28066_9158# vcm 0.89fF
C17566 a_23046_16186# rowoff_n[14] 1.64fF
C17567 a_24962_1126# m2_24824_946# 0.31fF
C17568 a_2475_17214# col[14] 0.22fF
C17569 col_n[30] rowoff_n[4] 0.12fF
C17570 col_n[26] rowoff_n[0] 0.15fF
C17571 col_n[29] rowoff_n[3] 0.13fF
C17572 col_n[27] rowoff_n[1] 0.14fF
C17573 col_n[31] rowoff_n[5] 0.11fF
C17574 col_n[28] rowoff_n[2] 0.14fF
C17575 a_2475_6170# col[19] 0.22fF
C17576 a_34090_16186# m2_34864_16006# 0.86fF
C17577 a_2874_17190# VDD 0.29fF
C17578 a_2475_12194# a_23046_12170# 0.68fF
C17579 a_12002_12170# a_13006_12170# 0.86fF
C17580 a_24050_11166# row_n[9] 0.43fF
C17581 a_18330_3174# vcm 0.24fF
C17582 a_23958_15182# rowon_n[13] 0.14fF
C17583 a_8990_12170# vcm 0.89fF
C17584 a_2275_12194# col_n[26] 0.17fF
C17585 a_5886_2130# VDD 0.29fF
C17586 a_2275_1150# col_n[31] 0.19fF
C17587 a_6982_9158# col[4] 0.38fF
C17588 a_30986_5142# a_31078_5142# 0.45fF
C17589 a_33998_5142# rowon_n[3] 0.14fF
C17590 m2_9764_946# m3_9896_1078# 4.41fF
C17591 a_2275_9182# a_14010_9158# 0.71fF
C17592 a_22042_5142# col_n[19] 0.34fF
C17593 a_2475_18218# m2_29844_18014# 0.62fF
C17594 a_2275_9182# col[16] 0.17fF
C17595 a_32082_17190# col_n[29] 0.34fF
C17596 a_33390_7190# vcm 0.24fF
C17597 col_n[19] rowoff_n[10] 0.20fF
C17598 a_24050_16186# vcm 0.89fF
C17599 a_20946_6146# VDD 0.29fF
C17600 a_2475_6170# a_6890_6146# 0.41fF
C17601 a_2275_6170# a_4274_6186# 0.15fF
C17602 a_10998_9158# rowon_n[7] 0.45fF
C17603 a_2275_11190# a_29070_11166# 0.71fF
C17604 a_26970_1126# vcm 0.18fF
C17605 a_27062_16186# a_28066_16186# 0.86fF
C17606 a_14314_10202# vcm 0.24fF
C17607 a_10998_17190# rowoff_n[15] 2.23fF
C17608 m2_23820_18014# VDD 3.15fF
C17609 a_9902_6146# rowoff_n[4] 0.66fF
C17610 a_27062_5142# ctop 4.91fF
C17611 a_16018_2130# m2_15788_946# 0.84fF
C17612 a_2475_8178# a_21950_8154# 0.41fF
C17613 a_2275_8178# a_19334_8194# 0.15fF
C17614 a_11910_8154# a_12002_8154# 0.45fF
C17615 col_n[1] rowon_n[15] 0.17fF
C17616 col_n[0] rowon_n[14] 0.17fF
C17617 VDD rowon_n[13] 4.61fF
C17618 sample row_n[14] 0.92fF
C17619 vcm row_n[15] 1.08fF
C17620 col[20] rowoff_n[15] 0.21fF
C17621 a_7894_4138# vcm 0.18fF
C17622 a_10998_3134# col_n[8] 0.34fF
C17623 a_18938_4138# rowoff_n[2] 0.56fF
C17624 col_n[3] rowoff_n[11] 0.32fF
C17625 a_21038_15182# col_n[18] 0.34fF
C17626 a_32082_8154# row_n[6] 0.43fF
C17627 a_29374_14218# vcm 0.24fF
C17628 a_31990_12170# rowon_n[10] 0.14fF
C17629 a_2275_5166# a_12914_5142# 0.17fF
C17630 a_7986_8154# ctop 4.91fF
C17631 a_16930_13174# VDD 0.29fF
C17632 a_2275_10186# a_35398_10202# 0.15fF
C17633 a_27974_2130# rowoff_n[0] 0.46fF
C17634 a_2275_8178# col_n[3] 0.17fF
C17635 a_22954_8154# vcm 0.18fF
C17636 a_2475_2154# a_4974_2130# 0.68fF
C17637 a_10298_17230# vcm 0.24fF
C17638 a_8990_16186# rowon_n[14] 0.45fF
C17639 a_31078_2130# col[28] 0.38fF
C17640 m2_12776_18014# col[10] 0.37fF
C17641 a_2275_7174# a_27974_7150# 0.17fF
C17642 a_23046_12170# ctop 4.91fF
C17643 a_31990_17190# VDD 0.29fF
C17644 a_26970_12170# a_27062_12170# 0.45fF
C17645 a_19030_6146# rowon_n[4] 0.45fF
C17646 a_2275_16210# a_5978_16186# 0.71fF
C17647 a_2475_15206# col[8] 0.22fF
C17648 a_2475_4162# col[13] 0.22fF
C17649 a_34090_2130# VDD 1.39fF
C17650 a_26362_2170# col_n[23] 0.11fF
C17651 a_2475_4162# a_20034_4138# 0.68fF
C17652 a_28066_5142# a_28066_4138# 0.84fF
C17653 a_9994_13174# col_n[7] 0.34fF
C17654 a_3970_15182# ctop 4.91fF
C17655 a_2275_10186# col_n[20] 0.17fF
C17656 a_20034_10162# rowoff_n[8] 1.79fF
C17657 a_30074_15182# row_n[13] 0.43fF
C17658 a_23958_13174# rowoff_n[11] 0.50fF
C17659 a_2275_1150# a_10998_1126# 0.14fF
C17660 a_18938_15182# vcm 0.18fF
C17661 a_15014_5142# VDD 3.20fF
C17662 a_18026_6146# a_19030_6146# 0.86fF
C17663 a_2275_7174# col[10] 0.17fF
C17664 a_29070_8154# rowoff_n[6] 1.35fF
C17665 a_34394_14218# col_n[31] 0.11fF
C17666 a_30074_12170# col[27] 0.38fF
C17667 m2_28840_18014# col_n[26] 0.33fF
C17668 a_7894_15182# a_7986_15182# 0.45fF
C17669 a_2475_15206# a_13918_15182# 0.41fF
C17670 a_2275_15206# a_11302_15222# 0.15fF
C17671 a_2475_17214# col[25] 0.22fF
C17672 a_2475_6170# col[30] 0.22fF
C17673 a_2275_3158# a_26058_3134# 0.71fF
C17674 a_2475_1150# m2_34864_946# 0.58fF
C17675 a_2275_1150# m2_32856_946# 0.52fF
C17676 a_30074_9158# VDD 1.65fF
C17677 a_20034_16186# m2_20232_16434# 0.19fF
C17678 a_8990_8154# a_8990_7150# 0.84fF
C17679 a_17022_13174# rowon_n[11] 0.45fF
C17680 a_25358_12210# col_n[22] 0.11fF
C17681 a_2275_12194# a_4882_12170# 0.17fF
C17682 a_2966_12170# a_3970_12170# 0.86fF
C17683 a_2475_3158# vcm 1.32fF
C17684 a_27062_3134# rowon_n[1] 0.45fF
C17685 a_2275_17214# a_26362_17230# 0.15fF
C17686 a_2475_17214# a_28978_17190# 0.41fF
C17687 a_10998_12170# VDD 3.61fF
C17688 a_33086_10162# a_34090_10162# 0.86fF
C17689 a_2275_9182# col[27] 0.17fF
C17690 a_2275_14202# a_19942_14178# 0.17fF
C17691 a_4974_3134# row_n[1] 0.43fF
C17692 a_19030_10162# col[16] 0.38fF
C17693 col_n[30] rowoff_n[10] 0.12fF
C17694 a_17022_7150# vcm 0.89fF
C17695 a_4882_7150# rowon_n[5] 0.14fF
C17696 a_11910_14178# rowoff_n[12] 0.64fF
C17697 a_2475_2154# a_33998_2130# 0.41fF
C17698 a_2275_2154# a_31382_2170# 0.15fF
C17699 a_17934_2130# a_18026_2130# 0.45fF
C17700 a_2275_6170# VDD 3.18fF
C17701 a_34090_6146# col_n[31] 0.34fF
C17702 a_10998_14178# m2_11196_14426# 0.19fF
C17703 a_26058_16186# VDD 2.06fF
C17704 a_24050_12170# a_24050_11166# 0.84fF
C17705 a_2475_11190# a_12002_11166# 0.68fF
C17706 a_14314_10202# col_n[11] 0.11fF
C17707 a_7286_1166# vcm 0.25fF
C17708 a_2275_16210# a_35002_16186# 0.17fF
C17709 a_7986_2130# m2_8184_2378# 0.19fF
C17710 a_32082_11166# vcm 0.89fF
C17711 a_28978_1126# VDD 0.72fF
C17712 a_30074_10162# m2_30272_10410# 0.19fF
C17713 col_n[3] row_n[11] 0.37fF
C17714 VDD row_n[8] 4.64fF
C17715 col_n[11] row_n[15] 0.37fF
C17716 col_n[9] row_n[14] 0.37fF
C17717 col_n[7] row_n[13] 0.37fF
C17718 col_n[1] row_n[10] 0.37fF
C17719 col_n[0] row_n[9] 0.37fF
C17720 vcm rowon_n[9] 0.91fF
C17721 col_n[6] rowon_n[12] 0.17fF
C17722 col_n[10] rowon_n[14] 0.17fF
C17723 col_n[8] rowon_n[13] 0.17fF
C17724 col_n[12] rowon_n[15] 0.17fF
C17725 col_n[4] rowon_n[11] 0.17fF
C17726 col_n[5] row_n[12] 0.37fF
C17727 col_n[2] rowon_n[10] 0.17fF
C17728 sample rowon_n[8] 0.10fF
C17729 col[31] rowoff_n[15] 0.14fF
C17730 a_2475_8178# a_3878_8154# 0.41fF
C17731 a_2275_8178# a_2874_8154# 0.17fF
C17732 a_2475_13198# col[2] 0.22fF
C17733 a_2475_2154# col[7] 0.22fF
C17734 a_25054_10162# rowon_n[8] 0.45fF
C17735 a_2475_13198# a_27062_13174# 0.68fF
C17736 a_14010_13174# a_15014_13174# 0.86fF
C17737 col_n[14] rowoff_n[11] 0.24fF
C17738 a_22346_5182# vcm 0.24fF
C17739 m2_34864_1950# a_35002_2130# 0.33fF
C17740 a_7986_8154# col[5] 0.38fF
C17741 a_13006_14178# vcm 0.89fF
C17742 a_9902_4138# VDD 0.29fF
C17743 a_1957_12194# m2_1732_11990# 0.33fF
C17744 a_32994_6146# a_33086_6146# 0.45fF
C17745 a_2275_8178# col_n[14] 0.17fF
C17746 a_2275_10186# a_18026_10162# 0.71fF
C17747 a_23046_4138# col_n[20] 0.34fF
C17748 a_33086_16186# col_n[30] 0.34fF
C17749 a_4974_15182# a_4974_14178# 0.84fF
C17750 a_3270_8194# vcm 0.24fF
C17751 a_2275_5166# col[4] 0.17fF
C17752 a_21038_8154# m2_21236_8402# 0.19fF
C17753 a_12914_4138# rowon_n[2] 0.14fF
C17754 a_16018_3134# ctop 4.91fF
C17755 a_28066_18194# vcm 0.15fF
C17756 a_24962_8154# VDD 0.29fF
C17757 a_2475_7174# a_10906_7150# 0.41fF
C17758 a_2275_7174# a_8290_7190# 0.15fF
C17759 sample rowoff_n[12] 0.22fF
C17760 a_2475_15206# col[19] 0.22fF
C17761 a_2275_12194# a_33086_12170# 0.71fF
C17762 a_2475_4162# col[24] 0.22fF
C17763 a_30986_3134# vcm 0.18fF
C17764 a_29070_17190# a_30074_17190# 0.86fF
C17765 a_18330_12210# vcm 0.24fF
C17766 a_10906_5142# rowoff_n[3] 0.65fF
C17767 m2_15788_946# col[13] 0.51fF
C17768 a_31078_7150# ctop 4.91fF
C17769 a_5886_11166# VDD 0.29fF
C17770 a_2275_10186# col_n[31] 0.17fF
C17771 a_23046_17190# rowon_n[15] 0.45fF
C17772 a_2275_9182# a_23350_9198# 0.15fF
C17773 a_2475_9182# a_25966_9158# 0.41fF
C17774 a_13918_9158# a_14010_9158# 0.45fF
C17775 m2_1732_7974# sample_n 0.12fF
C17776 m2_1732_3958# rowoff_n[2] 2.46fF
C17777 a_12002_2130# col_n[9] 0.34fF
C17778 a_19942_3134# rowoff_n[1] 0.55fF
C17779 a_1957_10186# rowoff_n[8] 0.14fF
C17780 a_11910_6146# vcm 0.18fF
C17781 a_33086_7150# rowon_n[5] 0.45fF
C17782 a_22042_14178# col_n[19] 0.34fF
C17783 a_12002_6146# m2_12200_6394# 0.19fF
C17784 a_33390_16226# vcm 0.24fF
C17785 a_2475_18218# a_4882_18194# 0.41fF
C17786 a_2275_7174# col[21] 0.17fF
C17787 a_2275_6170# a_16930_6146# 0.17fF
C17788 a_12002_10162# ctop 4.91fF
C17789 a_20946_15182# VDD 0.29fF
C17790 m2_5748_18014# vcm 0.71fF
C17791 row_n[5] rowoff_n[5] 0.64fF
C17792 a_10998_7150# row_n[5] 0.43fF
C17793 a_10906_11166# rowon_n[9] 0.14fF
C17794 a_26970_10162# vcm 0.18fF
C17795 a_2475_3158# a_8990_3134# 0.68fF
C17796 a_4974_3134# a_5978_3134# 0.86fF
C17797 m3_34996_14130# ctop 0.22fF
C17798 a_2275_8178# a_31990_8154# 0.17fF
C17799 a_27062_14178# ctop 4.91fF
C17800 a_28978_13174# a_29070_13174# 0.45fF
C17801 a_2475_18218# VDD 42.20fF
C17802 a_12002_11166# rowoff_n[9] 2.18fF
C17803 a_2275_17214# a_9994_17190# 0.71fF
C17804 a_27366_1166# col_n[24] 0.11fF
C17805 m2_1732_18014# m2_2160_18442# 0.19fF
C17806 a_7894_13174# vcm 0.18fF
C17807 a_10998_12170# col_n[8] 0.34fF
C17808 a_3970_3134# VDD 4.33fF
C17809 a_2475_5166# a_24050_5142# 0.68fF
C17810 a_30074_6146# a_30074_5142# 0.84fF
C17811 a_2275_18218# a_20034_18194# 0.14fF
C17812 m2_4744_946# m2_5748_946# 0.86fF
C17813 a_7986_17190# ctop 4.93fF
C17814 a_21038_9158# rowoff_n[7] 1.74fF
C17815 a_31078_14178# rowon_n[12] 0.45fF
C17816 a_2275_17214# col_n[3] 0.17fF
C17817 a_28066_15182# rowoff_n[13] 1.40fF
C17818 a_2275_6170# col_n[8] 0.17fF
C17819 m2_34864_1950# m3_34996_2082# 4.42fF
C17820 a_2275_2154# a_15014_2130# 0.71fF
C17821 a_22954_17190# vcm 0.18fF
C17822 a_19030_7150# VDD 2.78fF
C17823 a_30074_7150# rowoff_n[5] 1.30fF
C17824 a_20034_7150# a_21038_7150# 0.86fF
C17825 a_31078_11166# col[28] 0.38fF
C17826 a_8990_14178# row_n[12] 0.43fF
C17827 a_25054_2130# vcm 0.89fF
C17828 a_9902_16186# a_9994_16186# 0.45fF
C17829 a_2275_16210# a_15318_16226# 0.15fF
C17830 a_2475_16210# a_17934_16186# 0.41fF
C17831 a_19030_4138# row_n[2] 0.43fF
C17832 col_n[7] rowon_n[7] 0.17fF
C17833 col_n[23] rowon_n[15] 0.17fF
C17834 col_n[5] rowon_n[6] 0.17fF
C17835 col_n[12] row_n[10] 0.37fF
C17836 col_n[21] rowon_n[14] 0.17fF
C17837 col_n[3] rowon_n[5] 0.17fF
C17838 col_n[10] row_n[9] 0.37fF
C17839 col_n[19] rowon_n[13] 0.17fF
C17840 col_n[8] row_n[8] 0.37fF
C17841 col_n[14] row_n[11] 0.37fF
C17842 vcm row_n[4] 1.08fF
C17843 col_n[6] row_n[7] 0.37fF
C17844 col_n[22] row_n[15] 0.37fF
C17845 sample row_n[3] 0.92fF
C17846 col_n[4] row_n[6] 0.37fF
C17847 VDD rowon_n[2] 4.61fF
C17848 col_n[11] rowon_n[9] 0.17fF
C17849 col_n[9] rowon_n[8] 0.17fF
C17850 col_n[16] row_n[12] 0.37fF
C17851 col_n[15] rowon_n[11] 0.17fF
C17852 col_n[13] rowon_n[10] 0.17fF
C17853 col_n[0] rowon_n[3] 0.17fF
C17854 col_n[17] rowon_n[12] 0.17fF
C17855 col_n[1] rowon_n[4] 0.17fF
C17856 col_n[18] row_n[13] 0.37fF
C17857 col_n[2] row_n[5] 0.37fF
C17858 col_n[20] row_n[14] 0.37fF
C17859 a_18938_8154# rowon_n[6] 0.14fF
C17860 a_2275_4162# a_30074_4138# 0.71fF
C17861 a_2475_13198# col[13] 0.22fF
C17862 a_26362_11206# col_n[23] 0.11fF
C17863 a_34090_11166# VDD 1.23fF
C17864 m3_25960_1078# m3_26964_1078# 0.21fF
C17865 a_2475_2154# col[18] 0.22fF
C17866 a_2966_17190# m2_3164_17438# 0.19fF
C17867 a_10998_9158# a_10998_8154# 0.84fF
C17868 col_n[25] rowoff_n[11] 0.16fF
C17869 m2_34864_2954# vcm 0.72fF
C17870 a_2275_13198# a_8898_13174# 0.17fF
C17871 a_5978_5142# vcm 0.89fF
C17872 a_2475_1150# a_22954_1126# 0.41fF
C17873 a_2275_8178# col_n[25] 0.17fF
C17874 a_2275_1150# a_20338_1166# 0.19fF
C17875 a_15014_14178# VDD 3.20fF
C17876 m2_34864_10986# row_n[9] 0.38fF
C17877 a_5978_2130# rowon_n[0] 0.45fF
C17878 a_20034_9158# col[17] 0.38fF
C17879 a_2275_16210# col[10] 0.17fF
C17880 a_2275_15206# a_23958_15182# 0.17fF
C17881 a_2275_5166# col[15] 0.17fF
C17882 a_21038_9158# vcm 0.89fF
C17883 a_16018_16186# rowoff_n[14] 1.98fF
C17884 a_19942_3134# a_20034_3134# 0.45fF
C17885 col_n[9] rowoff_n[12] 0.27fF
C17886 a_2475_15206# col[30] 0.22fF
C17887 a_15318_9198# col_n[12] 0.11fF
C17888 a_26058_13174# a_26058_12170# 0.84fF
C17889 a_2475_12194# a_16018_12170# 0.68fF
C17890 a_11302_3174# vcm 0.24fF
C17891 a_17022_11166# row_n[9] 0.43fF
C17892 a_16930_15182# rowon_n[13] 0.14fF
C17893 a_2475_12194# vcm 1.32fF
C17894 a_32994_3134# VDD 0.29fF
C17895 a_26970_5142# rowon_n[3] 0.14fF
C17896 a_2275_9182# a_6982_9158# 0.71fF
C17897 a_2475_18218# m2_15788_18014# 0.62fF
C17898 a_16018_14178# a_17022_14178# 0.86fF
C17899 a_2475_14202# a_31078_14178# 0.68fF
C17900 a_26362_7190# vcm 0.24fF
C17901 a_8990_7150# col[6] 0.38fF
C17902 m2_1732_4962# VDD 5.46fF
C17903 a_17022_16186# vcm 0.89fF
C17904 a_13918_6146# VDD 0.29fF
C17905 a_35002_7150# a_35094_7150# 0.11fF
C17906 a_24050_3134# col_n[21] 0.34fF
C17907 a_3970_9158# rowon_n[7] 0.45fF
C17908 rowon_n[1] rowoff_n[1] 20.66fF
C17909 a_2275_15206# VDD 3.18fF
C17910 ctop rowoff_n[7] 0.28fF
C17911 a_34090_15182# col_n[31] 0.34fF
C17912 a_2275_11190# a_22042_11166# 0.71fF
C17913 a_2275_4162# col_n[2] 0.17fF
C17914 a_19942_1126# vcm 0.18fF
C17915 a_4274_7190# col_n[1] 0.11fF
C17916 a_6982_16186# a_6982_15182# 0.84fF
C17917 a_7286_10202# vcm 0.24fF
C17918 a_3970_17190# rowoff_n[15] 2.57fF
C17919 m2_9764_18014# VDD 4.55fF
C17920 a_2161_6170# rowoff_n[4] 0.14fF
C17921 a_20034_5142# ctop 4.91fF
C17922 a_28978_10162# VDD 0.29fF
C17923 a_26058_17190# m2_26256_17438# 0.19fF
C17924 a_2275_8178# a_12306_8194# 0.15fF
C17925 a_2475_8178# a_14922_8154# 0.41fF
C17926 a_35002_5142# vcm 0.18fF
C17927 a_2475_11190# col[7] 0.22fF
C17928 a_11910_4138# rowoff_n[2] 0.64fF
C17929 a_28978_12170# rowoff_n[10] 0.44fF
C17930 a_25054_8154# row_n[6] 0.43fF
C17931 a_22346_14218# vcm 0.24fF
C17932 a_24962_12170# rowon_n[10] 0.14fF
C17933 a_7986_17190# col[5] 0.38fF
C17934 a_2275_5166# a_5886_5142# 0.17fF
C17935 a_9902_13174# VDD 0.29fF
C17936 a_2275_10186# a_27366_10202# 0.15fF
C17937 a_2475_10186# a_29982_10162# 0.41fF
C17938 a_15926_10162# a_16018_10162# 0.45fF
C17939 a_2275_17214# col_n[14] 0.17fF
C17940 a_2966_9158# rowoff_n[7] 2.62fF
C17941 a_20946_2130# rowoff_n[0] 0.54fF
C17942 a_35002_2130# rowon_n[0] 0.14fF
C17943 a_2275_6170# col_n[19] 0.17fF
C17944 a_23046_13174# col_n[20] 0.34fF
C17945 a_2275_18218# col_n[0] 0.17fF
C17946 m2_1732_8978# m2_2160_9406# 0.19fF
C17947 a_15926_8154# vcm 0.18fF
C17948 a_17022_3134# a_17022_2130# 0.84fF
C17949 a_3270_17230# vcm 0.24fF
C17950 m2_8760_18014# m3_8892_18146# 4.41fF
C17951 a_2475_16210# rowon_n[14] 0.40fF
C17952 a_35494_8516# VDD 0.13fF
C17953 a_2275_14202# col[4] 0.17fF
C17954 a_17022_15182# m2_17220_15430# 0.19fF
C17955 a_2275_7174# a_20946_7150# 0.17fF
C17956 a_16018_12170# ctop 4.91fF
C17957 a_2275_3158# col[9] 0.17fF
C17958 a_24962_17190# VDD 0.29fF
C17959 a_12002_6146# rowon_n[4] 0.45fF
C17960 col_n[24] rowon_n[10] 0.17fF
C17961 col_n[3] row_n[0] 0.37fF
C17962 col_n[22] rowon_n[9] 0.17fF
C17963 col_n[20] rowon_n[8] 0.17fF
C17964 col_n[27] row_n[12] 0.37fF
C17965 col_n[26] rowon_n[11] 0.17fF
C17966 col_n[18] rowon_n[7] 0.17fF
C17967 col_n[16] rowon_n[6] 0.17fF
C17968 col_n[23] row_n[10] 0.37fF
C17969 col_n[14] rowon_n[5] 0.17fF
C17970 col_n[21] row_n[9] 0.37fF
C17971 col_n[28] rowon_n[12] 0.17fF
C17972 col_n[7] row_n[2] 0.37fF
C17973 col_n[5] row_n[1] 0.37fF
C17974 col_n[9] row_n[3] 0.37fF
C17975 col_n[11] row_n[4] 0.37fF
C17976 col_n[29] row_n[13] 0.37fF
C17977 col_n[4] rowon_n[0] 0.17fF
C17978 col_n[13] row_n[5] 0.37fF
C17979 col_n[31] row_n[14] 0.37fF
C17980 col_n[6] rowon_n[1] 0.17fF
C17981 VDD en_bit_n[2] 0.34fF
C17982 col_n[15] row_n[6] 0.37fF
C17983 col_n[8] rowon_n[2] 0.17fF
C17984 col_n[17] row_n[7] 0.37fF
C17985 col_n[10] rowon_n[3] 0.17fF
C17986 col_n[25] row_n[11] 0.37fF
C17987 vcm ctop 2.09fF
C17988 col_n[19] row_n[8] 0.37fF
C17989 col_n[12] rowon_n[4] 0.17fF
C17990 col_n[30] rowon_n[13] 0.17fF
C17991 a_2475_13198# col[24] 0.22fF
C17992 a_30986_12170# vcm 0.18fF
C17993 a_2475_2154# col[29] 0.22fF
C17994 a_27062_2130# VDD 1.96fF
C17995 a_2475_4162# a_13006_4138# 0.68fF
C17996 a_6982_4138# a_7986_4138# 0.86fF
C17997 m3_34996_7102# m3_34996_6098# 0.20fF
C17998 a_2275_9182# a_34394_9198# 0.15fF
C17999 a_31078_16186# ctop 4.91fF
C18000 a_30986_14178# a_31078_14178# 0.45fF
C18001 a_13006_10162# rowoff_n[8] 2.13fF
C18002 a_23046_15182# row_n[13] 0.43fF
C18003 a_16930_13174# rowoff_n[11] 0.58fF
C18004 a_12002_11166# col_n[9] 0.34fF
C18005 a_2275_1150# a_3970_1126# 0.79fF
C18006 a_11910_15182# vcm 0.18fF
C18007 a_7986_5142# VDD 3.92fF
C18008 a_33086_5142# row_n[3] 0.43fF
C18009 a_32082_7150# a_32082_6146# 0.84fF
C18010 a_2475_6170# a_28066_6146# 0.68fF
C18011 a_7986_13174# m2_8184_13422# 0.19fF
C18012 a_32994_9158# rowon_n[7] 0.14fF
C18013 a_2275_16210# col[21] 0.17fF
C18014 a_22042_8154# rowoff_n[6] 1.69fF
C18015 a_2275_5166# col[26] 0.17fF
C18016 a_2275_15206# a_4274_15222# 0.15fF
C18017 a_2475_15206# a_6890_15182# 0.41fF
C18018 m2_34864_12994# m2_34864_11990# 0.84fF
C18019 a_2966_9158# vcm 0.89fF
C18020 m2_25828_946# col[23] 0.51fF
C18021 col_n[20] rowoff_n[12] 0.19fF
C18022 a_32994_17190# rowoff_n[15] 0.40fF
C18023 a_31078_6146# rowoff_n[4] 1.25fF
C18024 a_27062_9158# m2_27260_9406# 0.19fF
C18025 a_2275_3158# a_19030_3134# 0.71fF
C18026 a_7894_1126# m2_7756_946# 0.31fF
C18027 m3_18932_1078# ctop 0.29fF
C18028 a_23046_9158# VDD 2.37fF
C18029 a_32082_10162# col[29] 0.38fF
C18030 a_22042_8154# a_23046_8154# 0.86fF
C18031 a_9994_13174# rowon_n[11] 0.45fF
C18032 a_29070_4138# vcm 0.89fF
C18033 a_20034_3134# rowon_n[1] 0.45fF
C18034 a_2275_17214# a_19334_17230# 0.15fF
C18035 a_2475_17214# a_21950_17190# 0.41fF
C18036 a_11910_17190# a_12002_17190# 0.45fF
C18037 a_27366_10202# col_n[24] 0.11fF
C18038 a_2275_5166# a_34090_5142# 0.71fF
C18039 a_2275_18218# a_29374_18234# 0.15fF
C18040 a_3970_12170# VDD 4.33fF
C18041 m2_15788_946# m2_16216_1374# 0.19fF
C18042 a_13006_10162# a_13006_9158# 0.84fF
C18043 a_2475_9182# col[1] 0.22fF
C18044 a_2275_14202# a_12914_14178# 0.17fF
C18045 col_n[4] rowoff_n[13] 0.31fF
C18046 a_9994_7150# vcm 0.89fF
C18047 a_4882_14178# rowoff_n[12] 0.72fF
C18048 a_31078_12170# row_n[10] 0.43fF
C18049 a_18026_7150# m2_18224_7398# 0.19fF
C18050 a_2475_2154# a_26970_2130# 0.41fF
C18051 a_2275_2154# a_24354_2170# 0.15fF
C18052 a_30986_16186# rowon_n[14] 0.14fF
C18053 col[7] rowoff_n[9] 0.30fF
C18054 col[6] rowoff_n[8] 0.31fF
C18055 col[5] rowoff_n[7] 0.31fF
C18056 col[0] rowoff_n[2] 0.34fF
C18057 col[1] rowoff_n[3] 0.34fF
C18058 col[2] rowoff_n[4] 0.33fF
C18059 col[3] rowoff_n[5] 0.33fF
C18060 col[4] rowoff_n[6] 0.32fF
C18061 a_2275_15206# col_n[8] 0.17fF
C18062 a_2275_4162# col_n[13] 0.17fF
C18063 a_19030_16186# VDD 2.78fF
C18064 a_21038_8154# col[18] 0.38fF
C18065 a_2475_11190# a_4974_11166# 0.68fF
C18066 a_35398_2170# vcm 0.24fF
C18067 a_2275_16210# a_27974_16186# 0.17fF
C18068 a_3270_4178# col_n[0] 0.11fF
C18069 a_25054_11166# vcm 0.89fF
C18070 a_2275_1150# col[3] 0.17fF
C18071 a_21950_1126# VDD 0.80fF
C18072 a_21950_4138# a_22042_4138# 0.45fF
C18073 a_16322_8194# col_n[13] 0.11fF
C18074 a_2475_11190# col[18] 0.22fF
C18075 a_18026_10162# rowon_n[8] 0.45fF
C18076 a_2475_13198# a_20034_13174# 0.68fF
C18077 a_28066_14178# a_28066_13174# 0.84fF
C18078 a_15318_5182# vcm 0.24fF
C18079 m2_29268_2378# a_29070_2130# 0.19fF
C18080 m2_12776_946# vcm 0.71fF
C18081 a_8990_5142# m2_9188_5390# 0.19fF
C18082 a_2275_1150# a_32994_1126# 0.17fF
C18083 a_5978_14178# vcm 0.89fF
C18084 a_2161_4162# VDD 0.23fF
C18085 a_2275_17214# col_n[25] 0.17fF
C18086 a_2275_6170# col_n[30] 0.17fF
C18087 a_2275_10186# a_10998_10162# 0.71fF
C18088 a_2275_18218# col_n[10] 0.17fF
C18089 a_2275_2154# rowoff_n[0] 0.81fF
C18090 a_9994_6146# col[7] 0.38fF
C18091 a_18026_15182# a_19030_15182# 0.86fF
C18092 a_30378_9198# vcm 0.24fF
C18093 a_2275_14202# col[15] 0.17fF
C18094 a_5886_4138# rowon_n[2] 0.14fF
C18095 a_8990_3134# ctop 4.91fF
C18096 a_2275_3158# col[20] 0.17fF
C18097 a_21038_18194# vcm 0.15fF
C18098 a_25054_2130# col_n[22] 0.34fF
C18099 a_17934_8154# VDD 0.29fF
C18100 a_2966_15182# m2_1732_15002# 0.86fF
C18101 col_n[20] row_n[3] 0.37fF
C18102 col_n[18] row_n[2] 0.37fF
C18103 VDD col[8] 11.45fF
C18104 col_n[16] row_n[1] 0.37fF
C18105 rowon_n[12] row_n[12] 21.02fF
C18106 col_n[14] row_n[0] 0.37fF
C18107 col_n[31] rowon_n[8] 0.17fF
C18108 col_n[17] rowon_n[1] 0.17fF
C18109 col_n[24] row_n[5] 0.37fF
C18110 col_n[22] row_n[4] 0.37fF
C18111 col_n[15] rowon_n[0] 0.17fF
C18112 vcm col[5] 6.66fF
C18113 col_n[26] row_n[6] 0.37fF
C18114 col_n[19] rowon_n[2] 0.17fF
C18115 col_n[28] row_n[7] 0.37fF
C18116 col_n[21] rowon_n[3] 0.17fF
C18117 col_n[30] row_n[8] 0.37fF
C18118 col_n[23] rowon_n[4] 0.17fF
C18119 col_n[25] rowon_n[5] 0.17fF
C18120 col_n[2] col[3] 6.22fF
C18121 col_n[27] rowon_n[6] 0.17fF
C18122 col_n[29] rowon_n[7] 0.17fF
C18123 a_2275_12194# a_26058_12170# 0.71fF
C18124 a_5278_6186# col_n[2] 0.11fF
C18125 a_23958_3134# vcm 0.18fF
C18126 a_15318_18234# col_n[12] 0.11fF
C18127 a_8990_17190# a_8990_16186# 0.84fF
C18128 a_18026_1126# en_bit_n[1] 0.28fF
C18129 a_11302_12210# vcm 0.24fF
C18130 a_24050_7150# ctop 4.91fF
C18131 a_32994_12170# VDD 0.29fF
C18132 m2_14784_946# m3_14916_1078# 4.41fF
C18133 m3_21944_18146# m3_22948_18146# 0.21fF
C18134 a_16018_17190# rowon_n[15] 0.45fF
C18135 a_2275_9182# a_16322_9198# 0.15fF
C18136 a_2475_9182# a_18938_9158# 0.41fF
C18137 m2_1732_5966# vcm 1.11fF
C18138 a_12914_3134# rowoff_n[1] 0.63fF
C18139 a_4882_6146# vcm 0.18fF
C18140 a_26058_7150# rowon_n[5] 0.45fF
C18141 a_33086_14178# rowoff_n[12] 1.15fF
C18142 a_28066_2130# a_29070_2130# 0.86fF
C18143 a_26362_16226# vcm 0.24fF
C18144 a_8990_16186# col[6] 0.38fF
C18145 a_2275_6170# a_9902_6146# 0.17fF
C18146 a_4974_10162# ctop 4.91fF
C18147 a_13918_15182# VDD 0.29fF
C18148 a_17934_11166# a_18026_11166# 0.45fF
C18149 a_2275_11190# a_31382_11206# 0.15fF
C18150 a_2475_11190# a_33998_11166# 0.41fF
C18151 a_24050_12170# col_n[21] 0.34fF
C18152 col_n[31] rowoff_n[12] 0.11fF
C18153 a_3970_7150# row_n[5] 0.43fF
C18154 a_2275_13198# col_n[2] 0.17fF
C18155 a_19942_10162# vcm 0.18fF
C18156 a_2275_2154# col_n[7] 0.17fF
C18157 a_4274_16226# col_n[1] 0.11fF
C18158 a_1957_6170# sample 0.35fF
C18159 a_19030_4138# a_19030_3134# 0.84fF
C18160 m3_14916_18146# ctop 0.21fF
C18161 a_2275_8178# a_24962_8154# 0.17fF
C18162 a_35002_17190# m2_34864_17010# 0.33fF
C18163 a_20034_14178# ctop 4.91fF
C18164 a_4974_11166# rowoff_n[9] 2.52fF
C18165 a_2475_17214# a_3878_17190# 0.41fF
C18166 a_2275_17214# a_2874_17190# 0.17fF
C18167 m2_34864_12994# rowon_n[11] 0.42fF
C18168 a_35002_14178# vcm 0.18fF
C18169 a_31078_4138# VDD 1.54fF
C18170 a_2475_9182# col[12] 0.22fF
C18171 a_2475_5166# a_17022_5142# 0.68fF
C18172 a_8990_5142# a_9994_5142# 0.86fF
C18173 a_2275_18218# a_13006_18194# 0.14fF
C18174 col_n[15] rowoff_n[13] 0.23fF
C18175 a_14010_9158# rowoff_n[7] 2.08fF
C18176 a_24050_14178# rowon_n[12] 0.45fF
C18177 a_32994_15182# a_33086_15182# 0.45fF
C18178 a_13006_10162# col_n[10] 0.34fF
C18179 a_2275_15206# col_n[19] 0.17fF
C18180 col[9] rowoff_n[0] 0.29fF
C18181 col[10] rowoff_n[1] 0.28fF
C18182 col[11] rowoff_n[2] 0.27fF
C18183 col[12] rowoff_n[3] 0.27fF
C18184 col[13] rowoff_n[4] 0.26fF
C18185 col[14] rowoff_n[5] 0.25fF
C18186 col[15] rowoff_n[6] 0.25fF
C18187 col[16] rowoff_n[7] 0.24fF
C18188 col[17] rowoff_n[8] 0.23fF
C18189 col[18] rowoff_n[9] 0.23fF
C18190 a_21038_15182# rowoff_n[13] 1.74fF
C18191 a_2275_4162# col_n[24] 0.17fF
C18192 a_34090_4138# rowon_n[2] 0.45fF
C18193 a_2275_2154# a_7986_2130# 0.71fF
C18194 a_15926_17190# vcm 0.18fF
C18195 a_12002_7150# VDD 3.51fF
C18196 a_23046_7150# rowoff_n[5] 1.64fF
C18197 a_34090_8154# a_34090_7150# 0.84fF
C18198 a_2475_7174# a_32082_7150# 0.68fF
C18199 a_35494_17552# VDD 0.13fF
C18200 a_2475_14202# row_n[12] 0.48fF
C18201 a_2275_12194# col[9] 0.17fF
C18202 a_18026_2130# vcm 0.89fF
C18203 a_2275_1150# col[14] 0.17fF
C18204 a_2275_16210# a_8290_16226# 0.15fF
C18205 a_2475_16210# a_10906_16186# 0.41fF
C18206 a_12002_4138# row_n[2] 0.43fF
C18207 a_32082_5142# rowoff_n[3] 1.20fF
C18208 a_3878_1126# VDD 0.90fF
C18209 a_33086_9158# col[30] 0.38fF
C18210 a_11910_8154# rowon_n[6] 0.14fF
C18211 a_2275_4162# a_23046_4138# 0.71fF
C18212 a_27062_11166# VDD 1.96fF
C18213 a_2475_11190# col[29] 0.22fF
C18214 m3_11904_1078# m3_12908_1078# 0.21fF
C18215 col_n[0] rowoff_n[14] 0.34fF
C18216 a_24050_9158# a_25054_9158# 0.86fF
C18217 col[2] rowoff_n[10] 0.33fF
C18218 a_33086_6146# vcm 0.89fF
C18219 a_13918_18194# a_14010_18194# 0.11fF
C18220 a_28370_9198# col_n[25] 0.11fF
C18221 a_8898_1126# a_8990_1126# 0.11fF
C18222 a_2475_1150# a_15926_1126# 0.41fF
C18223 a_2275_1150# a_13310_1166# 0.15fF
C18224 a_2275_18218# col_n[21] 0.17fF
C18225 m2_16792_946# VDD 5.20fF
C18226 m2_1732_15002# row_n[13] 0.44fF
C18227 a_7986_14178# VDD 3.92fF
C18228 a_15014_11166# a_15014_10162# 0.84fF
C18229 a_2275_14202# col[26] 0.17fF
C18230 a_2275_15206# a_16930_15182# 0.17fF
C18231 a_2275_3158# col[31] 0.17fF
C18232 a_32082_11166# rowon_n[9] 0.45fF
C18233 a_14010_9158# vcm 0.89fF
C18234 a_8990_16186# rowoff_n[14] 2.33fF
C18235 a_2275_3158# a_28370_3174# 0.15fF
C18236 a_2475_3158# a_30986_3134# 0.41fF
C18237 col_n[30] rowon_n[2] 0.17fF
C18238 col_n[28] rowon_n[1] 0.17fF
C18239 col_n[26] rowon_n[0] 0.17fF
C18240 col_n[31] row_n[3] 0.37fF
C18241 col_n[8] col[8] 0.50fF
C18242 col_n[29] row_n[2] 0.37fF
C18243 VDD col[19] 8.73fF
C18244 vcm col[16] 6.66fF
C18245 col_n[25] row_n[0] 0.37fF
C18246 col_n[27] row_n[1] 0.37fF
C18247 a_23046_16186# m2_23244_16434# 0.19fF
C18248 a_22042_7150# col[19] 0.38fF
C18249 a_4974_12170# a_5978_12170# 0.86fF
C18250 a_2475_12194# a_8990_12170# 0.68fF
C18251 a_4274_3174# vcm 0.24fF
C18252 a_9994_11166# row_n[9] 0.43fF
C18253 a_33998_11166# rowoff_n[9] 0.39fF
C18254 a_2275_17214# a_31990_17190# 0.17fF
C18255 m2_6752_18014# col[4] 0.39fF
C18256 a_9902_15182# rowon_n[13] 0.14fF
C18257 a_29070_13174# vcm 0.89fF
C18258 a_25966_3134# VDD 0.29fF
C18259 a_23958_5142# a_24050_5142# 0.45fF
C18260 a_17326_7190# col_n[14] 0.11fF
C18261 a_19942_5142# rowon_n[3] 0.14fF
C18262 m2_27836_946# m2_28840_946# 0.86fF
C18263 a_2475_18218# m2_1732_18014# 0.17fF
C18264 a_2475_14202# a_24050_14178# 0.68fF
C18265 a_30074_15182# a_30074_14178# 0.84fF
C18266 a_2475_7174# col[6] 0.22fF
C18267 a_19334_7190# vcm 0.24fF
C18268 a_32082_2130# ctop 4.93fF
C18269 a_9994_16186# vcm 0.89fF
C18270 m2_1732_15002# m3_1864_15134# 4.42fF
C18271 a_6890_6146# VDD 0.29fF
C18272 a_14010_14178# m2_14208_14426# 0.19fF
C18273 a_2275_11190# a_15014_11166# 0.71fF
C18274 a_2275_13198# col_n[13] 0.17fF
C18275 a_10998_5142# col[8] 0.38fF
C18276 a_2275_2154# col_n[18] 0.17fF
C18277 a_12914_1126# vcm 0.18fF
C18278 a_21038_17190# col[18] 0.38fF
C18279 a_20034_16186# a_21038_16186# 0.86fF
C18280 a_10998_2130# m2_11196_2378# 0.19fF
C18281 a_35398_11206# vcm 0.24fF
C18282 a_32482_1488# VDD 0.12fF
C18283 a_33086_10162# m2_33284_10410# 0.19fF
C18284 a_3270_13214# col_n[0] 0.11fF
C18285 a_13006_5142# ctop 4.91fF
C18286 a_2275_10186# col[3] 0.17fF
C18287 a_21950_10162# VDD 0.29fF
C18288 a_2275_8178# a_5278_8194# 0.15fF
C18289 a_2475_8178# a_7894_8154# 0.41fF
C18290 m2_22816_18014# col_n[20] 0.32fF
C18291 a_4882_8154# a_4974_8154# 0.45fF
C18292 a_6282_5182# col_n[3] 0.11fF
C18293 a_16322_17230# col_n[13] 0.11fF
C18294 a_2275_13198# a_30074_13174# 0.71fF
C18295 a_27974_5142# vcm 0.18fF
C18296 a_21950_12170# rowoff_n[10] 0.52fF
C18297 a_4882_4138# rowoff_n[2] 0.72fF
C18298 a_2275_18218# m2_32856_18014# 0.51fF
C18299 a_2475_9182# col[23] 0.22fF
C18300 a_18026_8154# row_n[6] 0.43fF
C18301 a_15318_14218# vcm 0.24fF
C18302 a_17934_12170# rowon_n[10] 0.14fF
C18303 a_4974_12170# m2_5172_12418# 0.19fF
C18304 a_28066_9158# ctop 4.91fF
C18305 col_n[26] rowoff_n[13] 0.15fF
C18306 a_2161_13198# VDD 0.23fF
C18307 a_2275_10186# a_20338_10202# 0.15fF
C18308 a_2475_10186# a_22954_10162# 0.41fF
C18309 a_27974_2130# rowon_n[0] 0.14fF
C18310 a_13918_2130# rowoff_n[0] 0.61fF
C18311 col[29] rowoff_n[9] 0.15fF
C18312 col[28] rowoff_n[8] 0.16fF
C18313 col[27] rowoff_n[7] 0.17fF
C18314 col[26] rowoff_n[6] 0.17fF
C18315 col[25] rowoff_n[5] 0.18fF
C18316 col[24] rowoff_n[4] 0.19fF
C18317 col[23] rowoff_n[3] 0.19fF
C18318 col[22] rowoff_n[2] 0.20fF
C18319 col[21] rowoff_n[1] 0.21fF
C18320 col[20] rowoff_n[0] 0.21fF
C18321 a_2275_15206# col_n[30] 0.17fF
C18322 a_8898_8154# vcm 0.18fF
C18323 a_9994_15182# col[7] 0.38fF
C18324 a_2966_15182# rowoff_n[13] 2.62fF
C18325 a_24050_8154# m2_24248_8402# 0.19fF
C18326 a_30074_3134# a_31078_3134# 0.86fF
C18327 a_30378_18234# vcm 0.25fF
C18328 a_2275_7174# a_13918_7150# 0.17fF
C18329 a_8990_12170# ctop 4.91fF
C18330 a_2275_12194# col[20] 0.17fF
C18331 a_25054_11166# col_n[22] 0.34fF
C18332 a_17934_17190# VDD 0.29fF
C18333 a_2275_1150# col[25] 0.17fF
C18334 a_19942_12170# a_20034_12170# 0.45fF
C18335 a_4974_6146# rowon_n[4] 0.45fF
C18336 a_5278_15222# col_n[2] 0.11fF
C18337 a_2475_3158# m2_34864_2954# 0.56fF
C18338 a_2966_5142# col_n[0] 0.34fF
C18339 a_23958_12170# vcm 0.18fF
C18340 a_20034_2130# VDD 2.68fF
C18341 col_n[10] rowoff_n[14] 0.27fF
C18342 a_21038_5142# a_21038_4138# 0.84fF
C18343 a_2475_4162# a_5978_4138# 0.68fF
C18344 m3_34996_14130# m3_34996_13126# 0.20fF
C18345 a_2275_9182# a_28978_9158# 0.17fF
C18346 a_20946_18194# m2_20808_18014# 0.34fF
C18347 col[13] rowoff_n[10] 0.26fF
C18348 a_24050_16186# ctop 4.91fF
C18349 a_5978_10162# rowoff_n[8] 2.47fF
C18350 a_16018_15182# row_n[13] 0.43fF
C18351 a_9902_13174# rowoff_n[11] 0.66fF
C18352 a_15014_6146# m2_15212_6394# 0.19fF
C18353 a_4882_15182# vcm 0.18fF
C18354 m2_1732_11990# m3_1864_12122# 4.42fF
C18355 a_26058_5142# row_n[3] 0.43fF
C18356 a_2475_6170# a_21038_6146# 0.68fF
C18357 a_2275_13198# m2_1732_12994# 0.27fF
C18358 a_10998_6146# a_12002_6146# 0.86fF
C18359 a_25966_9158# rowon_n[7] 0.14fF
C18360 a_15014_8154# rowoff_n[6] 2.03fF
C18361 a_2475_5166# col[0] 0.20fF
C18362 a_14010_9158# col_n[11] 0.34fF
C18363 a_35002_16186# a_35094_16186# 0.11fF
C18364 vcm col[27] 6.66fF
C18365 row_n[15] ctop 0.27fF
C18366 VDD col[30] 6.01fF
C18367 col_n[13] col[14] 6.22fF
C18368 a_25966_17190# rowoff_n[15] 0.48fF
C18369 m2_34864_17010# VDD 1.59fF
C18370 a_2275_3158# a_12002_3134# 0.71fF
C18371 a_24050_6146# rowoff_n[4] 1.59fF
C18372 a_2275_11190# col_n[7] 0.17fF
C18373 a_2475_1150# m2_4744_946# 0.62fF
C18374 m3_1864_6098# ctop 0.22fF
C18375 a_16018_9158# VDD 3.09fF
C18376 a_1957_15206# sample 0.35fF
C18377 a_2874_13174# rowon_n[11] 0.14fF
C18378 a_22042_4138# vcm 0.89fF
C18379 a_13006_3134# rowon_n[1] 0.45fF
C18380 a_33086_4138# rowoff_n[2] 1.15fF
C18381 a_2475_17214# a_14922_17190# 0.41fF
C18382 a_2275_17214# a_12306_17230# 0.15fF
C18383 a_5978_4138# m2_6176_4386# 0.19fF
C18384 a_34090_8154# col[31] 0.38fF
C18385 a_2275_5166# a_27062_5142# 0.71fF
C18386 a_31078_13174# VDD 1.54fF
C18387 a_2275_18218# a_22346_18234# 0.15fF
C18388 m2_8760_946# m2_9188_1374# 0.19fF
C18389 a_26058_10162# a_27062_10162# 0.86fF
C18390 a_2475_7174# col[17] 0.22fF
C18391 a_2275_14202# a_5886_14178# 0.17fF
C18392 m2_9764_946# col[7] 0.51fF
C18393 a_29374_8194# col_n[26] 0.11fF
C18394 a_2874_7150# vcm 0.18fF
C18395 a_24050_12170# row_n[10] 0.43fF
C18396 a_2275_2154# a_17326_2170# 0.15fF
C18397 a_2475_2154# a_19942_2130# 0.41fF
C18398 a_10906_2130# a_10998_2130# 0.45fF
C18399 a_23958_16186# rowon_n[14] 0.14fF
C18400 a_2275_13198# col_n[24] 0.17fF
C18401 a_34090_15182# m2_34864_15002# 0.86fF
C18402 a_2275_2154# col_n[29] 0.17fF
C18403 a_34090_2130# row_n[0] 0.43fF
C18404 a_12002_16186# VDD 3.51fF
C18405 a_17022_12170# a_17022_11166# 0.84fF
C18406 a_33998_6146# rowon_n[4] 0.14fF
C18407 a_27366_2170# vcm 0.24fF
C18408 a_2275_16210# a_20946_16186# 0.17fF
C18409 a_18026_11166# vcm 0.89fF
C18410 a_2275_10186# col[14] 0.17fF
C18411 a_14922_1126# VDD 0.88fF
C18412 a_2275_4162# a_32386_4178# 0.15fF
C18413 a_2475_4162# a_35002_4138# 0.41fF
C18414 a_23046_6146# col[20] 0.38fF
C18415 a_3878_10162# VDD 0.29fF
C18416 a_17022_17190# m2_16792_18014# 0.84fF
C18417 a_2475_13198# a_13006_13174# 0.68fF
C18418 a_6982_13174# a_7986_13174# 0.86fF
C18419 a_10998_10162# rowon_n[8] 0.45fF
C18420 a_35002_10162# rowoff_n[8] 0.38fF
C18421 a_8290_5182# vcm 0.24fF
C18422 a_3878_12170# rowoff_n[10] 0.73fF
C18423 a_2275_1150# a_25966_1126# 0.17fF
C18424 row_n[13] rowoff_n[13] 0.64fF
C18425 a_33086_15182# vcm 0.89fF
C18426 a_18330_6186# col_n[15] 0.11fF
C18427 m2_1732_8978# m3_1864_9110# 4.42fF
C18428 a_29982_5142# VDD 0.29fF
C18429 a_25966_6146# a_26058_6146# 0.45fF
C18430 a_28370_18234# col_n[25] 0.11fF
C18431 sample_n rowoff_n[1] 0.55fF
C18432 col[31] rowoff_n[0] 0.14fF
C18433 a_2275_10186# a_3970_10162# 0.71fF
C18434 a_32082_16186# a_32082_15182# 0.84fF
C18435 a_2475_15206# a_28066_15182# 0.68fF
C18436 a_23350_9198# vcm 0.24fF
C18437 a_2275_12194# col[31] 0.17fF
C18438 a_14010_18194# vcm 0.15fF
C18439 a_32082_9158# row_n[7] 0.43fF
C18440 a_10906_8154# VDD 0.29fF
C18441 a_31990_13174# rowon_n[11] 0.14fF
C18442 a_12002_4138# col[9] 0.38fF
C18443 a_22042_16186# col[19] 0.38fF
C18444 a_2275_12194# a_19030_12170# 0.71fF
C18445 a_16930_3134# vcm 0.18fF
C18446 a_2275_9182# col_n[1] 0.17fF
C18447 a_22042_17190# a_23046_17190# 0.86fF
C18448 col_n[21] rowoff_n[14] 0.19fF
C18449 m2_33860_18014# m2_34864_18014# 0.86fF
C18450 a_4274_12210# vcm 0.24fF
C18451 a_1957_2154# VDD 0.28fF
C18452 col[24] rowoff_n[10] 0.19fF
C18453 a_17022_7150# ctop 4.91fF
C18454 a_7286_4178# col_n[4] 0.11fF
C18455 a_25966_12170# VDD 0.29fF
C18456 m3_7888_18146# m3_8892_18146# 0.21fF
C18457 a_6890_9158# a_6982_9158# 0.45fF
C18458 a_8990_17190# rowon_n[15] 0.45fF
C18459 a_2275_9182# a_9294_9198# 0.15fF
C18460 a_2475_9182# a_11910_9158# 0.41fF
C18461 a_17326_16226# col_n[14] 0.11fF
C18462 a_2275_14202# a_34090_14178# 0.71fF
C18463 a_5886_3134# rowoff_n[1] 0.70fF
C18464 a_19030_7150# rowon_n[5] 0.45fF
C18465 a_31990_7150# vcm 0.18fF
C18466 a_26058_14178# rowoff_n[12] 1.50fF
C18467 a_2475_16210# col[6] 0.22fF
C18468 a_19334_16226# vcm 0.24fF
C18469 a_2475_5166# col[11] 0.22fF
C18470 a_2475_6170# a_2966_6146# 0.65fF
C18471 a_2161_6170# a_2275_6170# 0.17fF
C18472 a_32082_11166# ctop 4.91fF
C18473 a_6890_15182# VDD 0.29fF
C18474 a_2475_11190# a_26970_11166# 0.41fF
C18475 a_2275_11190# a_24354_11206# 0.15fF
C18476 col_n[19] col[19] 0.50fF
C18477 rowon_n[9] ctop 0.37fF
C18478 col_n[5] rowoff_n[15] 0.30fF
C18479 a_10998_14178# col[8] 0.38fF
C18480 a_2275_11190# col_n[18] 0.17fF
C18481 a_12914_10162# vcm 0.18fF
C18482 col[8] rowoff_n[11] 0.29fF
C18483 a_30074_16186# row_n[14] 0.43fF
C18484 a_32082_4138# a_33086_4138# 0.86fF
C18485 a_26058_10162# col_n[23] 0.34fF
C18486 a_2275_8178# a_17934_8154# 0.17fF
C18487 a_29070_17190# m2_29268_17438# 0.19fF
C18488 a_13006_14178# ctop 4.91fF
C18489 a_21950_13174# a_22042_13174# 0.45fF
C18490 a_2275_8178# col[8] 0.17fF
C18491 a_6282_14218# col_n[3] 0.11fF
C18492 m2_1732_17010# rowon_n[15] 0.43fF
C18493 a_27974_14178# vcm 0.18fF
C18494 m2_1732_5966# m3_1864_6098# 4.42fF
C18495 a_24050_4138# VDD 2.27fF
C18496 a_23046_6146# a_23046_5142# 0.84fF
C18497 a_2475_5166# a_9994_5142# 0.68fF
C18498 a_2475_7174# col[28] 0.22fF
C18499 a_2275_18218# a_5978_18194# 0.14fF
C18500 a_2275_10186# a_32994_10162# 0.17fF
C18501 a_6982_9158# rowoff_n[7] 2.42fF
C18502 a_17022_14178# rowon_n[12] 0.45fF
C18503 a_14010_15182# rowoff_n[13] 2.08fF
C18504 a_27062_4138# rowon_n[2] 0.45fF
C18505 a_8898_17190# vcm 0.18fF
C18506 m2_13780_18014# m3_13912_18146# 4.41fF
C18507 a_4974_7150# VDD 4.23fF
C18508 a_16018_7150# rowoff_n[5] 1.98fF
C18509 a_13006_7150# a_14010_7150# 0.86fF
C18510 a_2475_7174# a_25054_7150# 0.68fF
C18511 a_20034_15182# m2_20232_15430# 0.19fF
C18512 a_15014_8154# col_n[12] 0.34fF
C18513 a_10998_2130# vcm 0.89fF
C18514 a_2275_10186# col[25] 0.17fF
C18515 m2_1732_16006# m2_1732_15002# 0.84fF
C18516 a_4974_4138# row_n[2] 0.43fF
C18517 a_25054_5142# rowoff_n[3] 1.54fF
C18518 a_4882_8154# rowon_n[6] 0.14fF
C18519 a_2275_4162# a_16018_4138# 0.71fF
C18520 a_2966_14178# col_n[0] 0.34fF
C18521 a_20034_11166# VDD 2.68fF
C18522 a_3970_9158# a_3970_8154# 0.84fF
C18523 a_34090_3134# rowoff_n[1] 1.10fF
C18524 a_26058_6146# vcm 0.89fF
C18525 m2_34864_1950# a_2275_2154# 0.51fF
C18526 a_2475_1150# a_8898_1126# 0.41fF
C18527 a_2275_1150# a_6282_1166# 0.15fF
C18528 a_2275_6170# a_31078_6146# 0.71fF
C18529 a_10998_13174# m2_11196_13422# 0.19fF
C18530 a_28066_11166# a_29070_11166# 0.86fF
C18531 m2_34864_18014# vcm 0.73fF
C18532 a_3970_6146# col_n[1] 0.34fF
C18533 a_30378_7190# col_n[27] 0.11fF
C18534 a_2275_15206# a_9902_15182# 0.17fF
C18535 a_2475_14202# col[0] 0.20fF
C18536 a_2475_3158# col[5] 0.22fF
C18537 a_25054_11166# rowon_n[9] 0.45fF
C18538 a_6982_9158# vcm 0.89fF
C18539 a_2475_16210# rowoff_n[14] 4.75fF
C18540 a_2275_3158# a_21342_3174# 0.15fF
C18541 a_2475_3158# a_23958_3134# 0.41fF
C18542 a_30074_9158# m2_30272_9406# 0.19fF
C18543 a_12914_3134# a_13006_3134# 0.45fF
C18544 a_2475_1150# m2_27836_946# 0.62fF
C18545 m3_33992_1078# ctop 0.34fF
C18546 a_2275_9182# col_n[12] 0.17fF
C18547 a_19030_13174# a_19030_12170# 0.84fF
C18548 a_31382_4178# vcm 0.24fF
C18549 a_26970_11166# rowoff_n[9] 0.47fF
C18550 a_2275_17214# a_24962_17190# 0.17fF
C18551 a_22042_13174# vcm 0.89fF
C18552 a_24050_5142# col[21] 0.38fF
C18553 m2_1732_2954# m3_1864_3086# 4.42fF
C18554 a_18938_3134# VDD 0.29fF
C18555 a_34090_17190# col[31] 0.38fF
C18556 a_1957_11190# m2_1732_10986# 0.33fF
C18557 a_2966_5142# a_2966_4138# 0.84fF
C18558 a_2275_6170# col[2] 0.17fF
C18559 a_12914_5142# rowon_n[3] 0.14fF
C18560 a_2275_18218# a_35002_18194# 0.17fF
C18561 m2_20808_946# m2_21812_946# 0.86fF
C18562 a_2475_14202# a_17022_14178# 0.68fF
C18563 a_8990_14178# a_9994_14178# 0.86fF
C18564 a_2475_16210# col[17] 0.22fF
C18565 a_12306_7190# vcm 0.24fF
C18566 a_19334_5182# col_n[16] 0.11fF
C18567 a_2475_5166# col[22] 0.22fF
C18568 a_2275_2154# a_29982_2130# 0.17fF
C18569 a_21038_7150# m2_21236_7398# 0.19fF
C18570 a_29374_17230# col_n[26] 0.11fF
C18571 a_25054_2130# ctop 4.93fF
C18572 a_2874_16186# vcm 0.18fF
C18573 a_33998_7150# VDD 0.29fF
C18574 a_27974_7150# a_28066_7150# 0.45fF
C18575 col_n[24] col[25] 6.22fF
C18576 col_n[16] rowoff_n[15] 0.22fF
C18577 rowon_n[1] row_n[1] 21.02fF
C18578 row_n[4] ctop 0.28fF
C18579 a_2275_11190# a_7986_11166# 0.71fF
C18580 a_2275_11190# col_n[29] 0.17fF
C18581 a_5886_1126# vcm 0.18fF
C18582 col[19] rowoff_n[11] 0.22fF
C18583 a_34090_17190# a_34090_16186# 0.84fF
C18584 a_2475_16210# a_32082_16186# 0.68fF
C18585 m2_1732_8978# sample 0.31fF
C18586 a_27366_11206# vcm 0.24fF
C18587 a_25454_1488# VDD 0.13fF
C18588 a_33086_8154# rowon_n[6] 0.45fF
C18589 a_5978_5142# ctop 4.91fF
C18590 a_13006_3134# col[10] 0.38fF
C18591 a_14922_10162# VDD 0.29fF
C18592 a_2275_8178# col[19] 0.17fF
C18593 a_23046_15182# col[20] 0.38fF
C18594 a_2275_13198# a_23046_13174# 0.71fF
C18595 m2_34864_3958# m2_35292_4386# 0.19fF
C18596 a_20946_5142# vcm 0.18fF
C18597 a_14922_12170# rowoff_n[10] 0.60fF
C18598 m2_32280_2378# a_32082_2130# 0.19fF
C18599 m2_21812_946# vcm 0.71fF
C18600 a_2275_18218# m2_18800_18014# 0.51fF
C18601 a_10998_8154# row_n[6] 0.43fF
C18602 a_12002_5142# m2_12200_5390# 0.19fF
C18603 a_19030_1126# a_20034_1126# 0.86fF
C18604 a_8290_14218# vcm 0.24fF
C18605 a_10906_12170# rowon_n[10] 0.14fF
C18606 a_8290_3174# col_n[5] 0.11fF
C18607 a_21038_9158# ctop 4.91fF
C18608 a_18330_15222# col_n[15] 0.11fF
C18609 a_29982_14178# VDD 0.29fF
C18610 a_8898_10162# a_8990_10162# 0.45fF
C18611 a_2475_10186# a_15926_10162# 0.41fF
C18612 a_2275_10186# a_13310_10202# 0.15fF
C18613 a_20946_2130# rowon_n[0] 0.14fF
C18614 a_6890_2130# rowoff_n[0] 0.69fF
C18615 col[3] rowoff_n[12] 0.33fF
C18616 a_34394_9198# vcm 0.24fF
C18617 a_30986_16186# rowoff_n[14] 0.42fF
C18618 a_9994_3134# a_9994_2130# 0.84fF
C18619 a_23350_18234# vcm 0.25fF
C18620 a_29982_1126# m2_29844_946# 0.31fF
C18621 a_2275_7174# a_6890_7150# 0.17fF
C18622 a_10906_17190# VDD 0.29fF
C18623 a_2475_12194# a_30986_12170# 0.41fF
C18624 a_2275_12194# a_28370_12210# 0.15fF
C18625 a_12002_13174# col[9] 0.38fF
C18626 a_31078_15182# rowon_n[13] 0.45fF
C18627 a_16930_12170# vcm 0.18fF
C18628 a_13006_2130# VDD 3.40fF
C18629 a_27062_9158# col_n[24] 0.34fF
C18630 a_2275_7174# col_n[6] 0.17fF
C18631 a_1957_11190# VDD 0.28fF
C18632 m2_20808_946# m3_20940_1078# 4.41fF
C18633 a_2275_9182# a_21950_9158# 0.17fF
C18634 a_17022_16186# ctop 4.91fF
C18635 a_7286_13214# col_n[4] 0.11fF
C18636 a_23958_14178# a_24050_14178# 0.45fF
C18637 a_2966_11166# col[0] 0.38fF
C18638 a_8990_15182# row_n[13] 0.43fF
C18639 a_2161_13198# rowoff_n[11] 0.14fF
C18640 a_31990_16186# vcm 0.18fF
C18641 a_28066_6146# VDD 1.85fF
C18642 a_19030_5142# row_n[3] 0.43fF
C18643 a_25054_7150# a_25054_6146# 0.84fF
C18644 a_2475_6170# a_14010_6146# 0.68fF
C18645 a_18938_9158# rowon_n[7] 0.14fF
C18646 a_7986_8154# rowoff_n[6] 2.38fF
C18647 a_2475_14202# col[11] 0.22fF
C18648 a_2475_3158# col[16] 0.22fF
C18649 a_35094_1126# vcm 0.15fF
C18650 a_2475_18218# col[2] 0.22fF
C18651 m2_34864_3958# rowon_n[2] 0.42fF
C18652 a_18938_17190# rowoff_n[15] 0.56fF
C18653 a_2275_3158# a_4974_3134# 0.71fF
C18654 a_3878_3134# a_3970_3134# 0.45fF
C18655 a_17022_6146# rowoff_n[4] 1.94fF
C18656 a_2275_9182# col_n[23] 0.17fF
C18657 a_8990_9158# VDD 3.82fF
C18658 m3_29976_18146# ctop 0.21fF
C18659 a_16018_7150# col_n[13] 0.34fF
C18660 a_15014_8154# a_16018_8154# 0.86fF
C18661 a_2966_16186# m2_3164_16434# 0.19fF
C18662 a_2475_8178# a_29070_8154# 0.68fF
C18663 a_15014_4138# vcm 0.89fF
C18664 a_5978_3134# rowon_n[1] 0.45fF
C18665 a_26058_4138# rowoff_n[2] 1.50fF
C18666 a_2275_17214# a_5278_17230# 0.15fF
C18667 a_2475_17214# a_7894_17190# 0.41fF
C18668 a_4882_17190# a_4974_17190# 0.45fF
C18669 a_2275_17214# col[8] 0.17fF
C18670 a_35002_1126# a_35094_1126# 0.11fF
C18671 a_2275_6170# col[13] 0.17fF
C18672 a_2275_5166# a_20034_5142# 0.71fF
C18673 a_24050_13174# VDD 2.27fF
C18674 a_2275_18218# a_15318_18234# 0.15fF
C18675 a_5978_10162# a_5978_9158# 0.84fF
C18676 a_2475_16210# col[28] 0.22fF
C18677 a_30074_8154# vcm 0.89fF
C18678 a_17022_12170# row_n[10] 0.43fF
C18679 a_2275_2154# a_10298_2170# 0.15fF
C18680 a_2475_2154# a_12914_2130# 0.41fF
C18681 col_n[27] rowoff_n[15] 0.14fF
C18682 col_n[30] col[30] 0.63fF
C18683 a_16930_16186# rowon_n[14] 0.14fF
C18684 a_2275_7174# a_35094_7150# 0.14fF
C18685 a_27062_2130# row_n[0] 0.43fF
C18686 a_4974_16186# VDD 4.23fF
C18687 col[30] rowoff_n[11] 0.15fF
C18688 a_30074_12170# a_31078_12170# 0.86fF
C18689 a_26970_6146# rowon_n[4] 0.14fF
C18690 a_31382_6186# col_n[28] 0.11fF
C18691 a_4974_5142# col_n[2] 0.34fF
C18692 a_20338_2170# vcm 0.24fF
C18693 a_15014_17190# col_n[12] 0.34fF
C18694 a_2275_16210# a_13918_16186# 0.17fF
C18695 a_10998_11166# vcm 0.89fF
C18696 a_7894_1126# VDD 0.95fF
C18697 a_2275_8178# col[30] 0.17fF
C18698 a_14922_4138# a_15014_4138# 0.45fF
C18699 a_2275_4162# a_25358_4178# 0.15fF
C18700 a_2475_4162# a_27974_4138# 0.41fF
C18701 m2_1732_5966# row_n[4] 0.44fF
C18702 a_3970_10162# rowon_n[8] 0.45fF
C18703 a_2475_13198# a_5978_13174# 0.68fF
C18704 a_21038_14178# a_21038_13174# 0.84fF
.ends

