magic
tech sky130A
timestamp 1659692990
<< metal2 >>
rect 14 623 628 628
rect 14 595 19 623
rect 47 595 67 623
rect 95 595 115 623
rect 143 595 163 623
rect 191 595 211 623
rect 239 595 259 623
rect 287 595 307 623
rect 335 595 355 623
rect 383 595 403 623
rect 431 595 451 623
rect 479 595 499 623
rect 527 595 547 623
rect 575 595 595 623
rect 623 595 628 623
rect 14 575 628 595
rect 14 547 19 575
rect 47 547 163 575
rect 191 547 307 575
rect 335 547 451 575
rect 479 547 595 575
rect 623 547 628 575
rect 14 527 628 547
rect 14 499 19 527
rect 47 499 163 527
rect 191 499 307 527
rect 335 499 451 527
rect 479 499 595 527
rect 623 499 628 527
rect 14 479 628 499
rect 14 451 19 479
rect 47 451 67 479
rect 95 451 115 479
rect 143 451 163 479
rect 191 451 211 479
rect 239 451 259 479
rect 287 451 307 479
rect 335 451 355 479
rect 383 451 403 479
rect 431 451 451 479
rect 479 451 499 479
rect 527 451 547 479
rect 575 451 595 479
rect 623 451 628 479
rect 14 431 628 451
rect 14 403 19 431
rect 47 403 163 431
rect 191 403 307 431
rect 335 403 451 431
rect 479 403 595 431
rect 623 403 628 431
rect 14 383 628 403
rect 14 355 19 383
rect 47 355 163 383
rect 191 355 307 383
rect 335 355 451 383
rect 479 355 595 383
rect 623 355 628 383
rect 14 335 628 355
rect 14 307 19 335
rect 47 307 67 335
rect 95 307 115 335
rect 143 307 163 335
rect 191 307 211 335
rect 239 307 259 335
rect 287 307 307 335
rect 335 307 355 335
rect 383 307 403 335
rect 431 307 451 335
rect 479 307 499 335
rect 527 307 547 335
rect 575 307 595 335
rect 623 307 628 335
rect 14 287 628 307
rect 14 259 19 287
rect 47 259 163 287
rect 191 259 307 287
rect 335 259 451 287
rect 479 259 595 287
rect 623 259 628 287
rect 14 239 628 259
rect 14 211 19 239
rect 47 211 163 239
rect 191 211 307 239
rect 335 211 451 239
rect 479 211 595 239
rect 623 211 628 239
rect 14 191 628 211
rect 14 163 19 191
rect 47 163 67 191
rect 95 163 115 191
rect 143 163 163 191
rect 191 163 211 191
rect 239 163 259 191
rect 287 163 307 191
rect 335 163 355 191
rect 383 163 403 191
rect 431 163 451 191
rect 479 163 499 191
rect 527 163 547 191
rect 575 163 595 191
rect 623 163 628 191
rect 14 143 628 163
rect 14 115 19 143
rect 47 115 163 143
rect 191 115 307 143
rect 335 115 451 143
rect 479 115 595 143
rect 623 115 628 143
rect 14 95 628 115
rect 14 67 19 95
rect 47 67 163 95
rect 191 67 307 95
rect 335 67 451 95
rect 479 67 595 95
rect 623 67 628 95
rect 14 47 628 67
rect 14 19 19 47
rect 47 19 67 47
rect 95 19 115 47
rect 143 19 163 47
rect 191 19 211 47
rect 239 19 259 47
rect 287 19 307 47
rect 335 19 355 47
rect 383 19 403 47
rect 431 19 451 47
rect 479 19 499 47
rect 527 19 547 47
rect 575 19 595 47
rect 623 19 628 47
rect 14 14 628 19
<< via2 >>
rect 19 595 47 623
rect 67 595 95 623
rect 115 595 143 623
rect 163 595 191 623
rect 211 595 239 623
rect 259 595 287 623
rect 307 595 335 623
rect 355 595 383 623
rect 403 595 431 623
rect 451 595 479 623
rect 499 595 527 623
rect 547 595 575 623
rect 595 595 623 623
rect 19 547 47 575
rect 163 547 191 575
rect 307 547 335 575
rect 451 547 479 575
rect 595 547 623 575
rect 19 499 47 527
rect 163 499 191 527
rect 307 499 335 527
rect 451 499 479 527
rect 595 499 623 527
rect 19 451 47 479
rect 67 451 95 479
rect 115 451 143 479
rect 163 451 191 479
rect 211 451 239 479
rect 259 451 287 479
rect 307 451 335 479
rect 355 451 383 479
rect 403 451 431 479
rect 451 451 479 479
rect 499 451 527 479
rect 547 451 575 479
rect 595 451 623 479
rect 19 403 47 431
rect 163 403 191 431
rect 307 403 335 431
rect 451 403 479 431
rect 595 403 623 431
rect 19 355 47 383
rect 163 355 191 383
rect 307 355 335 383
rect 451 355 479 383
rect 595 355 623 383
rect 19 307 47 335
rect 67 307 95 335
rect 115 307 143 335
rect 163 307 191 335
rect 211 307 239 335
rect 259 307 287 335
rect 307 307 335 335
rect 355 307 383 335
rect 403 307 431 335
rect 451 307 479 335
rect 499 307 527 335
rect 547 307 575 335
rect 595 307 623 335
rect 19 259 47 287
rect 163 259 191 287
rect 307 259 335 287
rect 451 259 479 287
rect 595 259 623 287
rect 19 211 47 239
rect 163 211 191 239
rect 307 211 335 239
rect 451 211 479 239
rect 595 211 623 239
rect 19 163 47 191
rect 67 163 95 191
rect 115 163 143 191
rect 163 163 191 191
rect 211 163 239 191
rect 259 163 287 191
rect 307 163 335 191
rect 355 163 383 191
rect 403 163 431 191
rect 451 163 479 191
rect 499 163 527 191
rect 547 163 575 191
rect 595 163 623 191
rect 19 115 47 143
rect 163 115 191 143
rect 307 115 335 143
rect 451 115 479 143
rect 595 115 623 143
rect 19 67 47 95
rect 163 67 191 95
rect 307 67 335 95
rect 451 67 479 95
rect 595 67 623 95
rect 19 19 47 47
rect 67 19 95 47
rect 115 19 143 47
rect 163 19 191 47
rect 211 19 239 47
rect 259 19 287 47
rect 307 19 335 47
rect 355 19 383 47
rect 403 19 431 47
rect 451 19 479 47
rect 499 19 527 47
rect 547 19 575 47
rect 595 19 623 47
<< metal3 >>
rect 16 623 626 626
rect 16 595 19 623
rect 47 595 67 623
rect 95 595 115 623
rect 143 595 163 623
rect 191 595 211 623
rect 239 595 259 623
rect 287 595 307 623
rect 335 595 355 623
rect 383 595 403 623
rect 431 595 451 623
rect 479 595 499 623
rect 527 595 547 623
rect 575 595 595 623
rect 623 595 626 623
rect 16 592 626 595
rect 16 575 50 592
rect 16 547 19 575
rect 47 547 50 575
rect 160 575 194 592
rect 16 527 50 547
rect 16 499 19 527
rect 47 499 50 527
rect 80 554 130 562
rect 80 520 88 554
rect 122 520 130 554
rect 80 512 130 520
rect 160 547 163 575
rect 191 547 194 575
rect 304 575 338 592
rect 160 527 194 547
rect 16 482 50 499
rect 160 499 163 527
rect 191 499 194 527
rect 224 554 274 562
rect 224 520 232 554
rect 266 520 274 554
rect 224 512 274 520
rect 304 547 307 575
rect 335 547 338 575
rect 448 575 482 592
rect 304 527 338 547
rect 160 482 194 499
rect 304 499 307 527
rect 335 499 338 527
rect 368 554 418 562
rect 368 520 376 554
rect 410 520 418 554
rect 368 512 418 520
rect 448 547 451 575
rect 479 547 482 575
rect 592 575 626 592
rect 448 527 482 547
rect 304 482 338 499
rect 448 499 451 527
rect 479 499 482 527
rect 512 554 562 562
rect 512 520 520 554
rect 554 520 562 554
rect 512 512 562 520
rect 592 547 595 575
rect 623 547 626 575
rect 592 527 626 547
rect 448 482 482 499
rect 592 499 595 527
rect 623 499 626 527
rect 592 482 626 499
rect 16 479 626 482
rect 16 451 19 479
rect 47 451 67 479
rect 95 451 115 479
rect 143 451 163 479
rect 191 451 211 479
rect 239 451 259 479
rect 287 451 307 479
rect 335 451 355 479
rect 383 451 403 479
rect 431 451 451 479
rect 479 451 499 479
rect 527 451 547 479
rect 575 451 595 479
rect 623 451 626 479
rect 16 448 626 451
rect 16 431 50 448
rect 16 403 19 431
rect 47 403 50 431
rect 160 431 194 448
rect 16 383 50 403
rect 16 355 19 383
rect 47 355 50 383
rect 80 410 130 418
rect 80 376 88 410
rect 122 376 130 410
rect 80 368 130 376
rect 160 403 163 431
rect 191 403 194 431
rect 304 431 338 448
rect 160 383 194 403
rect 16 338 50 355
rect 160 355 163 383
rect 191 355 194 383
rect 224 410 274 418
rect 224 376 232 410
rect 266 376 274 410
rect 224 368 274 376
rect 304 403 307 431
rect 335 403 338 431
rect 448 431 482 448
rect 304 383 338 403
rect 160 338 194 355
rect 304 355 307 383
rect 335 355 338 383
rect 368 410 418 418
rect 368 376 376 410
rect 410 376 418 410
rect 368 368 418 376
rect 448 403 451 431
rect 479 403 482 431
rect 592 431 626 448
rect 448 383 482 403
rect 304 338 338 355
rect 448 355 451 383
rect 479 355 482 383
rect 512 410 562 418
rect 512 376 520 410
rect 554 376 562 410
rect 512 368 562 376
rect 592 403 595 431
rect 623 403 626 431
rect 592 383 626 403
rect 448 338 482 355
rect 592 355 595 383
rect 623 355 626 383
rect 592 338 626 355
rect 16 335 626 338
rect 16 307 19 335
rect 47 307 67 335
rect 95 307 115 335
rect 143 307 163 335
rect 191 307 211 335
rect 239 307 259 335
rect 287 307 307 335
rect 335 307 355 335
rect 383 307 403 335
rect 431 307 451 335
rect 479 307 499 335
rect 527 307 547 335
rect 575 307 595 335
rect 623 307 626 335
rect 16 304 626 307
rect 16 287 50 304
rect 16 259 19 287
rect 47 259 50 287
rect 160 287 194 304
rect 16 239 50 259
rect 16 211 19 239
rect 47 211 50 239
rect 80 266 130 274
rect 80 232 88 266
rect 122 232 130 266
rect 80 224 130 232
rect 160 259 163 287
rect 191 259 194 287
rect 304 287 338 304
rect 160 239 194 259
rect 16 194 50 211
rect 160 211 163 239
rect 191 211 194 239
rect 224 266 274 274
rect 224 232 232 266
rect 266 232 274 266
rect 224 224 274 232
rect 304 259 307 287
rect 335 259 338 287
rect 448 287 482 304
rect 304 239 338 259
rect 160 194 194 211
rect 304 211 307 239
rect 335 211 338 239
rect 368 266 418 274
rect 368 232 376 266
rect 410 232 418 266
rect 368 224 418 232
rect 448 259 451 287
rect 479 259 482 287
rect 592 287 626 304
rect 448 239 482 259
rect 304 194 338 211
rect 448 211 451 239
rect 479 211 482 239
rect 512 266 562 274
rect 512 232 520 266
rect 554 232 562 266
rect 512 224 562 232
rect 592 259 595 287
rect 623 259 626 287
rect 592 239 626 259
rect 448 194 482 211
rect 592 211 595 239
rect 623 211 626 239
rect 592 194 626 211
rect 16 191 626 194
rect 16 163 19 191
rect 47 163 67 191
rect 95 163 115 191
rect 143 163 163 191
rect 191 163 211 191
rect 239 163 259 191
rect 287 163 307 191
rect 335 163 355 191
rect 383 163 403 191
rect 431 163 451 191
rect 479 163 499 191
rect 527 163 547 191
rect 575 163 595 191
rect 623 163 626 191
rect 16 160 626 163
rect 16 143 50 160
rect 16 115 19 143
rect 47 115 50 143
rect 160 143 194 160
rect 16 95 50 115
rect 16 67 19 95
rect 47 67 50 95
rect 80 122 130 130
rect 80 88 88 122
rect 122 88 130 122
rect 80 80 130 88
rect 160 115 163 143
rect 191 115 194 143
rect 304 143 338 160
rect 160 95 194 115
rect 16 50 50 67
rect 160 67 163 95
rect 191 67 194 95
rect 224 122 274 130
rect 224 88 232 122
rect 266 88 274 122
rect 224 80 274 88
rect 304 115 307 143
rect 335 115 338 143
rect 448 143 482 160
rect 304 95 338 115
rect 160 50 194 67
rect 304 67 307 95
rect 335 67 338 95
rect 368 122 418 130
rect 368 88 376 122
rect 410 88 418 122
rect 368 80 418 88
rect 448 115 451 143
rect 479 115 482 143
rect 592 143 626 160
rect 448 95 482 115
rect 304 50 338 67
rect 448 67 451 95
rect 479 67 482 95
rect 512 122 562 130
rect 512 88 520 122
rect 554 88 562 122
rect 512 80 562 88
rect 592 115 595 143
rect 623 115 626 143
rect 592 95 626 115
rect 448 50 482 67
rect 592 67 595 95
rect 623 67 626 95
rect 592 50 626 67
rect 16 47 626 50
rect 16 19 19 47
rect 47 19 67 47
rect 95 19 115 47
rect 143 19 163 47
rect 191 19 211 47
rect 239 19 259 47
rect 287 19 307 47
rect 335 19 355 47
rect 383 19 403 47
rect 431 19 451 47
rect 479 19 499 47
rect 527 19 547 47
rect 575 19 595 47
rect 623 19 626 47
rect 16 16 626 19
<< via3 >>
rect 88 520 122 554
rect 232 520 266 554
rect 376 520 410 554
rect 520 520 554 554
rect 88 376 122 410
rect 232 376 266 410
rect 376 376 410 410
rect 520 376 554 410
rect 88 232 122 266
rect 232 232 266 266
rect 376 232 410 266
rect 520 232 554 266
rect 88 88 122 122
rect 232 88 266 122
rect 376 88 410 122
rect 520 88 554 122
<< metal4 >>
rect 90 562 120 609
rect 234 562 264 609
rect 378 562 408 609
rect 522 562 552 609
rect 80 554 130 562
rect 80 552 88 554
rect 33 522 88 552
rect 80 520 88 522
rect 122 552 130 554
rect 224 554 274 562
rect 224 552 232 554
rect 122 522 232 552
rect 122 520 130 522
rect 80 512 130 520
rect 224 520 232 522
rect 266 552 274 554
rect 368 554 418 562
rect 368 552 376 554
rect 266 522 376 552
rect 266 520 274 522
rect 224 512 274 520
rect 368 520 376 522
rect 410 552 418 554
rect 512 554 562 562
rect 512 552 520 554
rect 410 522 520 552
rect 410 520 418 522
rect 368 512 418 520
rect 512 520 520 522
rect 554 552 562 554
rect 554 522 609 552
rect 554 520 562 522
rect 512 512 562 520
rect 90 418 120 512
rect 234 418 264 512
rect 378 418 408 512
rect 522 418 552 512
rect 80 410 130 418
rect 80 408 88 410
rect 33 378 88 408
rect 80 376 88 378
rect 122 408 130 410
rect 224 410 274 418
rect 224 408 232 410
rect 122 378 232 408
rect 122 376 130 378
rect 80 368 130 376
rect 224 376 232 378
rect 266 408 274 410
rect 368 410 418 418
rect 368 408 376 410
rect 266 378 376 408
rect 266 376 274 378
rect 224 368 274 376
rect 368 376 376 378
rect 410 408 418 410
rect 512 410 562 418
rect 512 408 520 410
rect 410 378 520 408
rect 410 376 418 378
rect 368 368 418 376
rect 512 376 520 378
rect 554 408 562 410
rect 554 378 609 408
rect 554 376 562 378
rect 512 368 562 376
rect 90 274 120 368
rect 234 274 264 368
rect 378 274 408 368
rect 522 274 552 368
rect 80 266 130 274
rect 80 264 88 266
rect 33 234 88 264
rect 80 232 88 234
rect 122 264 130 266
rect 224 266 274 274
rect 224 264 232 266
rect 122 234 232 264
rect 122 232 130 234
rect 80 224 130 232
rect 224 232 232 234
rect 266 264 274 266
rect 368 266 418 274
rect 368 264 376 266
rect 266 234 376 264
rect 266 232 274 234
rect 224 224 274 232
rect 368 232 376 234
rect 410 264 418 266
rect 512 266 562 274
rect 512 264 520 266
rect 410 234 520 264
rect 410 232 418 234
rect 368 224 418 232
rect 512 232 520 234
rect 554 264 562 266
rect 554 234 609 264
rect 554 232 562 234
rect 512 224 562 232
rect 90 130 120 224
rect 234 130 264 224
rect 378 130 408 224
rect 522 130 552 224
rect 80 122 130 130
rect 80 120 88 122
rect 33 90 88 120
rect 80 88 88 90
rect 122 120 130 122
rect 224 122 274 130
rect 224 120 232 122
rect 122 90 232 120
rect 122 88 130 90
rect 80 80 130 88
rect 224 88 232 90
rect 266 120 274 122
rect 368 122 418 130
rect 368 120 376 122
rect 266 90 376 120
rect 266 88 274 90
rect 224 80 274 88
rect 368 88 376 90
rect 410 120 418 122
rect 512 122 562 130
rect 512 120 520 122
rect 410 90 520 120
rect 410 88 418 90
rect 368 80 418 88
rect 512 88 520 90
rect 554 120 562 122
rect 554 90 609 120
rect 554 88 562 90
rect 512 80 562 88
rect 90 33 120 80
rect 234 33 264 80
rect 378 33 408 80
rect 522 33 552 80
<< comment >>
rect 0 628 14 642
rect 628 628 642 642
rect 0 0 14 14
rect 628 0 642 14
<< end >>
