* SPICE3 file created from adc_array_wafflecap_16.ext - technology: sky130A

.subckt adc_array_wafflecap_16 ctop cbot
C0 ctop cbot 8.71fF
C1 cbot VSUBS 2.76fF
.ends
