magic
tech sky130A
timestamp 1658401033
<< metal2 >>
rect 7 669 675 674
rect 7 641 12 669
rect 40 641 64 669
rect 92 641 116 669
rect 144 641 168 669
rect 198 641 222 669
rect 250 641 274 669
rect 302 641 326 669
rect 356 641 380 669
rect 408 641 432 669
rect 460 641 484 669
rect 514 641 538 669
rect 566 641 590 669
rect 618 641 642 669
rect 672 641 675 669
rect 7 617 675 641
rect 7 589 12 617
rect 40 589 168 617
rect 198 589 326 617
rect 356 589 484 617
rect 514 589 642 617
rect 672 589 675 617
rect 7 565 675 589
rect 7 537 12 565
rect 40 537 168 565
rect 198 537 326 565
rect 356 537 484 565
rect 514 537 642 565
rect 672 537 675 565
rect 7 513 675 537
rect 7 483 12 513
rect 40 483 64 513
rect 92 483 116 513
rect 144 483 168 513
rect 198 483 222 513
rect 250 483 274 513
rect 302 483 326 513
rect 356 483 380 513
rect 408 483 432 513
rect 460 483 484 513
rect 514 483 538 513
rect 566 483 590 513
rect 618 483 642 513
rect 672 483 675 513
rect 7 459 675 483
rect 7 431 12 459
rect 40 431 168 459
rect 198 431 326 459
rect 356 431 484 459
rect 514 431 642 459
rect 672 431 675 459
rect 7 407 675 431
rect 7 379 12 407
rect 40 379 168 407
rect 198 379 326 407
rect 356 379 484 407
rect 514 379 642 407
rect 672 379 675 407
rect 7 355 675 379
rect 7 325 12 355
rect 40 325 64 355
rect 92 325 116 355
rect 144 325 168 355
rect 198 325 222 355
rect 250 325 274 355
rect 302 325 326 355
rect 356 325 380 355
rect 408 325 432 355
rect 460 325 484 355
rect 514 325 538 355
rect 566 325 590 355
rect 618 325 642 355
rect 672 325 675 355
rect 7 301 675 325
rect 7 273 12 301
rect 40 273 168 301
rect 198 273 326 301
rect 356 273 484 301
rect 514 273 642 301
rect 672 273 675 301
rect 7 249 675 273
rect 7 221 12 249
rect 40 221 168 249
rect 198 221 326 249
rect 356 221 484 249
rect 514 221 642 249
rect 672 221 675 249
rect 7 197 675 221
rect 7 167 12 197
rect 40 167 64 197
rect 92 167 116 197
rect 144 167 168 197
rect 198 167 222 197
rect 250 167 274 197
rect 302 167 326 197
rect 356 167 380 197
rect 408 167 432 197
rect 460 167 484 197
rect 514 167 538 197
rect 566 167 590 197
rect 618 167 642 197
rect 672 167 675 197
rect 7 143 675 167
rect 7 115 12 143
rect 40 115 168 143
rect 198 115 326 143
rect 356 115 484 143
rect 514 115 642 143
rect 672 115 675 143
rect 7 91 675 115
rect 7 63 12 91
rect 40 63 168 91
rect 198 63 326 91
rect 356 63 484 91
rect 514 63 642 91
rect 672 63 675 91
rect 7 39 675 63
rect 7 11 12 39
rect 40 11 64 39
rect 92 11 116 39
rect 144 11 168 39
rect 198 11 222 39
rect 250 11 274 39
rect 302 11 326 39
rect 356 11 380 39
rect 408 11 432 39
rect 460 11 484 39
rect 514 11 538 39
rect 566 11 590 39
rect 618 11 642 39
rect 672 11 675 39
rect 7 6 675 11
<< via2 >>
rect 12 641 40 669
rect 64 641 92 669
rect 116 641 144 669
rect 168 641 198 669
rect 222 641 250 669
rect 274 641 302 669
rect 326 641 356 669
rect 380 641 408 669
rect 432 641 460 669
rect 484 641 514 669
rect 538 641 566 669
rect 590 641 618 669
rect 642 641 672 669
rect 12 589 40 617
rect 168 589 198 617
rect 326 589 356 617
rect 484 589 514 617
rect 642 589 672 617
rect 12 537 40 565
rect 168 537 198 565
rect 326 537 356 565
rect 484 537 514 565
rect 642 537 672 565
rect 12 483 40 513
rect 64 483 92 513
rect 116 483 144 513
rect 168 483 198 513
rect 222 483 250 513
rect 274 483 302 513
rect 326 483 356 513
rect 380 483 408 513
rect 432 483 460 513
rect 484 483 514 513
rect 538 483 566 513
rect 590 483 618 513
rect 642 483 672 513
rect 12 431 40 459
rect 168 431 198 459
rect 326 431 356 459
rect 484 431 514 459
rect 642 431 672 459
rect 12 379 40 407
rect 168 379 198 407
rect 326 379 356 407
rect 484 379 514 407
rect 642 379 672 407
rect 12 325 40 355
rect 64 325 92 355
rect 116 325 144 355
rect 168 325 198 355
rect 222 325 250 355
rect 274 325 302 355
rect 326 325 356 355
rect 380 325 408 355
rect 432 325 460 355
rect 484 325 514 355
rect 538 325 566 355
rect 590 325 618 355
rect 642 325 672 355
rect 12 273 40 301
rect 168 273 198 301
rect 326 273 356 301
rect 484 273 514 301
rect 642 273 672 301
rect 12 221 40 249
rect 168 221 198 249
rect 326 221 356 249
rect 484 221 514 249
rect 642 221 672 249
rect 12 167 40 197
rect 64 167 92 197
rect 116 167 144 197
rect 168 167 198 197
rect 222 167 250 197
rect 274 167 302 197
rect 326 167 356 197
rect 380 167 408 197
rect 432 167 460 197
rect 484 167 514 197
rect 538 167 566 197
rect 590 167 618 197
rect 642 167 672 197
rect 12 115 40 143
rect 168 115 198 143
rect 326 115 356 143
rect 484 115 514 143
rect 642 115 672 143
rect 12 63 40 91
rect 168 63 198 91
rect 326 63 356 91
rect 484 63 514 91
rect 642 63 672 91
rect 12 11 40 39
rect 64 11 92 39
rect 116 11 144 39
rect 168 11 198 39
rect 222 11 250 39
rect 274 11 302 39
rect 326 11 356 39
rect 380 11 408 39
rect 432 11 460 39
rect 484 11 514 39
rect 538 11 566 39
rect 590 11 618 39
rect 642 11 672 39
<< metal3 >>
rect 7 669 675 674
rect 7 641 12 669
rect 40 641 64 669
rect 92 641 116 669
rect 144 641 168 669
rect 198 641 222 669
rect 250 641 274 669
rect 302 641 326 669
rect 356 641 380 669
rect 408 641 432 669
rect 460 641 484 669
rect 514 641 538 669
rect 566 641 590 669
rect 618 641 642 669
rect 672 641 675 669
rect 7 638 675 641
rect 7 617 43 638
rect 7 589 12 617
rect 40 589 43 617
rect 165 617 201 638
rect 7 565 43 589
rect 7 537 12 565
rect 40 537 43 565
rect 79 593 129 602
rect 79 561 88 593
rect 120 561 129 593
rect 79 552 129 561
rect 165 589 168 617
rect 198 589 201 617
rect 323 617 359 638
rect 165 565 201 589
rect 7 516 43 537
rect 165 537 168 565
rect 198 537 201 565
rect 237 593 287 602
rect 237 561 246 593
rect 278 561 287 593
rect 237 552 287 561
rect 323 589 326 617
rect 356 589 359 617
rect 481 617 517 638
rect 323 565 359 589
rect 165 516 201 537
rect 323 537 326 565
rect 356 537 359 565
rect 395 593 445 602
rect 395 561 404 593
rect 436 561 445 593
rect 395 552 445 561
rect 481 589 484 617
rect 514 589 517 617
rect 639 617 675 638
rect 481 565 517 589
rect 323 516 359 537
rect 481 537 484 565
rect 514 537 517 565
rect 553 593 603 602
rect 553 561 562 593
rect 594 561 603 593
rect 553 552 603 561
rect 639 589 642 617
rect 672 589 675 617
rect 639 565 675 589
rect 481 516 517 537
rect 639 537 642 565
rect 672 537 675 565
rect 639 516 675 537
rect 7 513 675 516
rect 7 483 12 513
rect 40 483 64 513
rect 92 483 116 513
rect 144 483 168 513
rect 198 483 222 513
rect 250 483 274 513
rect 302 483 326 513
rect 356 483 380 513
rect 408 483 432 513
rect 460 483 484 513
rect 514 483 538 513
rect 566 483 590 513
rect 618 483 642 513
rect 672 483 675 513
rect 7 480 675 483
rect 7 459 43 480
rect 7 431 12 459
rect 40 431 43 459
rect 165 459 201 480
rect 7 407 43 431
rect 7 379 12 407
rect 40 379 43 407
rect 79 435 129 444
rect 79 403 88 435
rect 120 403 129 435
rect 79 394 129 403
rect 165 431 168 459
rect 198 431 201 459
rect 323 459 359 480
rect 165 407 201 431
rect 7 358 43 379
rect 165 379 168 407
rect 198 379 201 407
rect 237 435 287 444
rect 237 403 246 435
rect 278 403 287 435
rect 237 394 287 403
rect 323 431 326 459
rect 356 431 359 459
rect 481 459 517 480
rect 323 407 359 431
rect 165 358 201 379
rect 323 379 326 407
rect 356 379 359 407
rect 395 435 445 444
rect 395 403 404 435
rect 436 403 445 435
rect 395 394 445 403
rect 481 431 484 459
rect 514 431 517 459
rect 639 459 675 480
rect 481 407 517 431
rect 323 358 359 379
rect 481 379 484 407
rect 514 379 517 407
rect 553 435 603 444
rect 553 403 562 435
rect 594 403 603 435
rect 553 394 603 403
rect 639 431 642 459
rect 672 431 675 459
rect 639 407 675 431
rect 481 358 517 379
rect 639 379 642 407
rect 672 379 675 407
rect 639 358 675 379
rect 7 355 675 358
rect 7 325 12 355
rect 40 325 64 355
rect 92 325 116 355
rect 144 325 168 355
rect 198 325 222 355
rect 250 325 274 355
rect 302 325 326 355
rect 356 325 380 355
rect 408 325 432 355
rect 460 325 484 355
rect 514 325 538 355
rect 566 325 590 355
rect 618 325 642 355
rect 672 325 675 355
rect 7 322 675 325
rect 7 301 43 322
rect 7 273 12 301
rect 40 273 43 301
rect 165 301 201 322
rect 7 249 43 273
rect 7 221 12 249
rect 40 221 43 249
rect 79 277 129 286
rect 79 245 88 277
rect 120 245 129 277
rect 79 236 129 245
rect 165 273 168 301
rect 198 273 201 301
rect 323 301 359 322
rect 165 249 201 273
rect 7 200 43 221
rect 165 221 168 249
rect 198 221 201 249
rect 237 277 287 286
rect 237 245 246 277
rect 278 245 287 277
rect 237 236 287 245
rect 323 273 326 301
rect 356 273 359 301
rect 481 301 517 322
rect 323 249 359 273
rect 165 200 201 221
rect 323 221 326 249
rect 356 221 359 249
rect 395 277 445 286
rect 395 245 404 277
rect 436 245 445 277
rect 395 236 445 245
rect 481 273 484 301
rect 514 273 517 301
rect 639 301 675 322
rect 481 249 517 273
rect 323 200 359 221
rect 481 221 484 249
rect 514 221 517 249
rect 553 277 603 286
rect 553 245 562 277
rect 594 245 603 277
rect 553 236 603 245
rect 639 273 642 301
rect 672 273 675 301
rect 639 249 675 273
rect 481 200 517 221
rect 639 221 642 249
rect 672 221 675 249
rect 639 200 675 221
rect 7 197 675 200
rect 7 167 12 197
rect 40 167 64 197
rect 92 167 116 197
rect 144 167 168 197
rect 198 167 222 197
rect 250 167 274 197
rect 302 167 326 197
rect 356 167 380 197
rect 408 167 432 197
rect 460 167 484 197
rect 514 167 538 197
rect 566 167 590 197
rect 618 167 642 197
rect 672 167 675 197
rect 7 164 675 167
rect 7 143 43 164
rect 7 115 12 143
rect 40 115 43 143
rect 165 143 201 164
rect 7 91 43 115
rect 7 63 12 91
rect 40 63 43 91
rect 79 119 129 128
rect 79 87 88 119
rect 120 87 129 119
rect 79 78 129 87
rect 165 115 168 143
rect 198 115 201 143
rect 323 143 359 164
rect 165 91 201 115
rect 7 42 43 63
rect 165 63 168 91
rect 198 63 201 91
rect 237 119 287 128
rect 237 87 246 119
rect 278 87 287 119
rect 237 78 287 87
rect 323 115 326 143
rect 356 115 359 143
rect 481 143 517 164
rect 323 91 359 115
rect 165 42 201 63
rect 323 63 326 91
rect 356 63 359 91
rect 395 119 445 128
rect 395 87 404 119
rect 436 87 445 119
rect 395 78 445 87
rect 481 115 484 143
rect 514 115 517 143
rect 639 143 675 164
rect 481 91 517 115
rect 323 42 359 63
rect 481 63 484 91
rect 514 63 517 91
rect 553 119 603 128
rect 553 87 562 119
rect 594 87 603 119
rect 553 78 603 87
rect 639 115 642 143
rect 672 115 675 143
rect 639 91 675 115
rect 481 42 517 63
rect 639 63 642 91
rect 672 63 675 91
rect 639 42 675 63
rect 7 39 675 42
rect 7 11 12 39
rect 40 11 64 39
rect 92 11 116 39
rect 144 11 168 39
rect 198 11 222 39
rect 250 11 274 39
rect 302 11 326 39
rect 356 11 380 39
rect 408 11 432 39
rect 460 11 484 39
rect 514 11 538 39
rect 566 11 590 39
rect 618 11 642 39
rect 672 11 675 39
rect 7 6 675 11
<< via3 >>
rect 88 561 120 593
rect 246 561 278 593
rect 404 561 436 593
rect 562 561 594 593
rect 88 403 120 435
rect 246 403 278 435
rect 404 403 436 435
rect 562 403 594 435
rect 88 245 120 277
rect 246 245 278 277
rect 404 245 436 277
rect 562 245 594 277
rect 88 87 120 119
rect 246 87 278 119
rect 404 87 436 119
rect 562 87 594 119
<< metal4 >>
rect 89 608 119 656
rect 247 608 277 656
rect 405 608 435 656
rect 563 608 593 656
rect 73 593 135 608
rect 73 592 88 593
rect 25 562 88 592
rect 73 561 88 562
rect 120 592 135 593
rect 231 593 293 608
rect 231 592 246 593
rect 120 562 246 592
rect 120 561 135 562
rect 73 546 135 561
rect 231 561 246 562
rect 278 592 293 593
rect 389 593 451 608
rect 389 592 404 593
rect 278 562 404 592
rect 278 561 293 562
rect 231 546 293 561
rect 389 561 404 562
rect 436 592 451 593
rect 547 593 609 608
rect 547 592 562 593
rect 436 562 562 592
rect 436 561 451 562
rect 389 546 451 561
rect 547 561 562 562
rect 594 592 609 593
rect 594 562 657 592
rect 594 561 609 562
rect 547 546 609 561
rect 89 450 119 546
rect 247 450 277 546
rect 405 450 435 546
rect 563 450 593 546
rect 73 435 135 450
rect 73 434 88 435
rect 25 404 88 434
rect 73 403 88 404
rect 120 434 135 435
rect 231 435 293 450
rect 231 434 246 435
rect 120 404 246 434
rect 120 403 135 404
rect 73 388 135 403
rect 231 403 246 404
rect 278 434 293 435
rect 389 435 451 450
rect 389 434 404 435
rect 278 404 404 434
rect 278 403 293 404
rect 231 388 293 403
rect 389 403 404 404
rect 436 434 451 435
rect 547 435 609 450
rect 547 434 562 435
rect 436 404 562 434
rect 436 403 451 404
rect 389 388 451 403
rect 547 403 562 404
rect 594 434 609 435
rect 594 404 657 434
rect 594 403 609 404
rect 547 388 609 403
rect 89 292 119 388
rect 247 292 277 388
rect 405 292 435 388
rect 563 292 593 388
rect 73 277 135 292
rect 73 276 88 277
rect 25 246 88 276
rect 73 245 88 246
rect 120 276 135 277
rect 231 277 293 292
rect 231 276 246 277
rect 120 246 246 276
rect 120 245 135 246
rect 73 230 135 245
rect 231 245 246 246
rect 278 276 293 277
rect 389 277 451 292
rect 389 276 404 277
rect 278 246 404 276
rect 278 245 293 246
rect 231 230 293 245
rect 389 245 404 246
rect 436 276 451 277
rect 547 277 609 292
rect 547 276 562 277
rect 436 246 562 276
rect 436 245 451 246
rect 389 230 451 245
rect 547 245 562 246
rect 594 276 609 277
rect 594 246 657 276
rect 594 245 609 246
rect 547 230 609 245
rect 89 134 119 230
rect 247 134 277 230
rect 405 134 435 230
rect 563 134 593 230
rect 73 119 135 134
rect 73 118 88 119
rect 24 88 88 118
rect 73 87 88 88
rect 120 118 135 119
rect 231 119 293 134
rect 231 118 246 119
rect 120 88 246 118
rect 120 87 135 88
rect 73 72 135 87
rect 231 87 246 88
rect 278 118 293 119
rect 389 119 451 134
rect 389 118 404 119
rect 278 88 404 118
rect 278 87 293 88
rect 231 72 293 87
rect 389 87 404 88
rect 436 118 451 119
rect 547 119 609 134
rect 547 118 562 119
rect 436 88 562 118
rect 436 87 451 88
rect 389 72 451 87
rect 547 87 562 88
rect 594 118 609 119
rect 594 88 657 118
rect 594 87 609 88
rect 547 72 609 87
rect 89 24 119 72
rect 247 24 277 72
rect 405 24 435 72
rect 563 24 593 72
use adc_array_circuit  adc_array_circuit_0
timestamp 1658400657
transform 1 0 1 0 1 0
box 0 0 680 680
<< labels >>
rlabel metal4 25 576 25 576 7 CTOP
port 1 w
<< end >>
