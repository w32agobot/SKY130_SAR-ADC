magic
tech sky130A
magscale 1 2
timestamp 1662367448
<< nwell >>
rect -10 48 408 452
<< nmos >>
rect 88 -216 118 -116
rect 184 -216 214 -116
rect 280 -216 310 -116
<< pmos >>
rect 88 110 118 310
rect 184 110 214 310
rect 280 110 310 310
<< ndiff >>
rect 26 -128 88 -116
rect 26 -204 38 -128
rect 72 -204 88 -128
rect 26 -216 88 -204
rect 118 -128 184 -116
rect 118 -204 134 -128
rect 168 -204 184 -128
rect 118 -216 184 -204
rect 214 -128 280 -116
rect 214 -204 230 -128
rect 264 -204 280 -128
rect 214 -216 280 -204
rect 310 -128 372 -116
rect 310 -204 326 -128
rect 360 -204 372 -128
rect 310 -216 372 -204
<< pdiff >>
rect 26 298 88 310
rect 26 122 38 298
rect 72 122 88 298
rect 26 110 88 122
rect 118 298 184 310
rect 118 122 134 298
rect 168 122 184 298
rect 118 110 184 122
rect 214 298 280 310
rect 214 122 230 298
rect 264 122 280 298
rect 214 110 280 122
rect 310 298 372 310
rect 310 122 326 298
rect 360 122 372 298
rect 310 110 372 122
<< ndiffc >>
rect 38 -204 72 -128
rect 134 -204 168 -128
rect 230 -204 264 -128
rect 326 -204 360 -128
<< pdiffc >>
rect 38 122 72 298
rect 134 122 168 298
rect 230 122 264 298
rect 326 122 360 298
<< psubdiff >>
rect 26 -304 52 -270
rect 86 -304 120 -270
rect 154 -304 188 -270
rect 222 -304 256 -270
rect 290 -304 324 -270
rect 358 -304 382 -270
rect 26 -322 382 -304
<< nsubdiff >>
rect 26 378 50 416
rect 88 378 126 416
rect 164 378 202 416
rect 240 378 278 416
rect 316 378 372 416
<< psubdiffcont >>
rect 52 -304 86 -270
rect 120 -304 154 -270
rect 188 -304 222 -270
rect 256 -304 290 -270
rect 324 -304 358 -270
<< nsubdiffcont >>
rect 50 378 88 416
rect 126 378 164 416
rect 202 378 240 416
rect 278 378 316 416
<< poly >>
rect 184 336 310 366
rect 88 310 118 336
rect 184 310 214 336
rect 280 310 310 336
rect 88 84 118 110
rect 76 60 118 84
rect -42 -30 22 -18
rect 76 -30 108 60
rect 184 28 214 110
rect 280 84 310 110
rect -42 -66 108 -30
rect 150 11 214 28
rect 150 -23 160 11
rect 194 -23 214 11
rect 150 -40 214 -23
rect -42 -74 22 -66
rect 76 -68 108 -66
rect 76 -92 118 -68
rect 88 -116 118 -92
rect 184 -70 214 -40
rect 184 -100 310 -70
rect 184 -116 214 -100
rect 280 -116 310 -100
rect 88 -242 118 -216
rect 184 -242 214 -216
rect 280 -242 310 -216
<< polycont >>
rect 160 -23 194 11
<< locali >>
rect -42 378 50 416
rect 88 378 126 416
rect 164 378 202 416
rect 240 378 278 416
rect 316 378 408 416
rect 38 298 72 314
rect 38 28 72 122
rect 134 298 168 378
rect 134 106 168 122
rect 230 298 264 314
rect 38 11 196 28
rect 38 -23 160 11
rect 194 -23 196 11
rect 38 -40 196 -23
rect 230 -8 264 122
rect 326 298 360 378
rect 326 106 360 122
rect 38 -128 72 -40
rect 230 -46 408 -8
rect 38 -220 72 -204
rect 134 -128 168 -112
rect 134 -270 168 -204
rect 230 -128 264 -46
rect 230 -220 264 -204
rect 326 -128 360 -112
rect 326 -270 360 -204
rect 26 -288 52 -270
rect -42 -304 52 -288
rect 86 -304 120 -270
rect 154 -304 188 -270
rect 222 -304 256 -270
rect 290 -304 324 -270
rect 358 -304 382 -270
rect -42 -326 382 -304
<< comment >>
rect 134 88 168 102
rect 326 90 360 104
rect 134 -108 168 -96
rect 326 -108 360 -96
<< labels >>
rlabel locali -42 -326 -42 -288 7 VSS
port 2 w
rlabel locali -42 378 -42 416 7 VDD
port 1 w
rlabel locali 408 -46 408 -8 3 out
port 4 e
rlabel poly -42 -74 -42 -18 7 in
port 5 w
<< end >>
