VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO delay_macrocell
  CLASS CORE ;
  FOREIGN delay_macrocell ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.660 BY 2.720 ;
  SITE unithd ;
  PIN in
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.880000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.990 0.500 1.320 ;
    END
  END in
  PIN out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.366000 ;
    ANTENNADIFFAREA 0.361800 ;
    PORT
      LAYER li1 ;
        RECT 6.550 1.460 6.720 2.300 ;
        RECT 6.960 1.010 7.130 1.340 ;
        RECT 8.855 0.980 9.085 1.290 ;
        RECT 6.660 0.380 6.830 0.890 ;
      LAYER mcon ;
        RECT 6.550 1.540 6.720 1.820 ;
        RECT 6.960 1.090 7.130 1.260 ;
        RECT 8.885 1.100 9.055 1.270 ;
        RECT 6.660 0.720 6.830 0.890 ;
      LAYER met1 ;
        RECT 6.520 1.240 6.750 1.970 ;
        RECT 6.930 1.240 7.160 1.320 ;
        RECT 8.825 1.240 9.115 1.300 ;
        RECT 6.520 1.100 9.115 1.240 ;
        RECT 6.630 1.030 7.160 1.100 ;
        RECT 8.825 1.070 9.115 1.100 ;
        RECT 6.630 0.660 6.860 1.030 ;
    END
  END out
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.635 9.660 2.805 ;
        RECT 0.750 1.395 0.920 2.235 ;
        RECT 5.590 1.460 5.760 2.635 ;
        RECT 7.300 1.290 7.470 2.635 ;
        RECT 7.300 1.120 7.850 1.290 ;
        RECT 7.680 0.380 7.850 1.120 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 0.750 1.475 0.920 2.155 ;
      LAYER met1 ;
        RECT 0.000 2.480 9.660 2.960 ;
        RECT 0.720 1.415 0.950 2.480 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 8.150 1.180 8.320 2.300 ;
        RECT 8.150 1.010 8.670 1.180 ;
        RECT 0.750 0.455 0.920 0.915 ;
        RECT 5.700 0.085 5.870 0.840 ;
        RECT 8.500 0.085 8.670 1.010 ;
        RECT 0.000 -0.085 9.660 0.085 ;
      LAYER mcon ;
        RECT 0.750 0.535 0.920 0.835 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
      LAYER met1 ;
        RECT 0.720 0.240 0.950 0.910 ;
        RECT 5.020 0.240 5.540 0.680 ;
        RECT 0.000 -0.240 9.660 0.240 ;
      LAYER via ;
        RECT 5.120 0.290 5.440 0.640 ;
      LAYER met2 ;
        RECT 5.020 0.240 5.540 0.680 ;
      LAYER via2 ;
        RECT 5.120 0.300 5.440 0.670 ;
      LAYER met3 ;
        RECT 1.210 0.700 4.890 2.480 ;
        RECT 6.090 0.700 8.360 2.480 ;
        RECT 1.210 0.270 8.360 0.700 ;
    END
  END VGND
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.235 9.850 2.910 ;
    END
  END VPB
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 -0.085 9.655 1.070 ;
    END
  END VNB
  OBS
      LAYER li1 ;
        RECT 5.040 1.180 5.210 2.235 ;
        RECT 6.070 1.460 6.240 2.300 ;
        RECT 7.640 1.460 7.840 2.300 ;
        RECT 8.630 1.460 8.830 2.300 ;
        RECT 5.630 1.180 5.990 1.290 ;
        RECT 5.040 1.010 5.990 1.180 ;
        RECT 5.040 0.365 5.210 1.010 ;
        RECT 6.180 0.380 6.350 0.840 ;
        RECT 7.200 0.380 7.370 0.840 ;
        RECT 8.160 0.380 8.330 0.840 ;
      LAYER mcon ;
        RECT 5.040 1.475 5.210 2.085 ;
        RECT 6.070 1.540 6.240 2.220 ;
        RECT 7.670 1.640 7.840 2.220 ;
        RECT 8.630 1.640 8.800 2.220 ;
        RECT 5.630 1.070 5.910 1.240 ;
        RECT 6.180 0.460 6.350 0.760 ;
        RECT 7.200 0.460 7.370 0.660 ;
        RECT 8.160 0.460 8.330 0.660 ;
      LAYER met1 ;
        RECT 5.010 1.290 5.240 2.195 ;
        RECT 6.040 2.110 8.830 2.280 ;
        RECT 6.040 1.480 6.270 2.110 ;
        RECT 7.640 1.580 7.870 2.110 ;
        RECT 8.600 1.580 8.830 2.110 ;
        RECT 5.010 1.010 5.990 1.290 ;
        RECT 6.150 0.520 6.380 0.820 ;
        RECT 7.170 0.520 7.400 0.720 ;
        RECT 8.130 0.520 8.360 0.720 ;
        RECT 6.150 0.380 8.360 0.520 ;
      LAYER via ;
        RECT 5.630 1.020 5.910 1.280 ;
      LAYER met2 ;
        RECT 5.260 0.840 5.990 1.430 ;
      LAYER met4 ;
        RECT 5.250 1.340 5.660 1.430 ;
        RECT 4.330 0.970 6.690 1.340 ;
        RECT 5.250 0.840 5.660 0.970 ;
  END
END delay_macrocell
END LIBRARY

