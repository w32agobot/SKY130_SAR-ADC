magic
tech sky130A
magscale 1 2
timestamp 1671366669
<< nwell >>
rect 0 506 1004 880
<< nmos >>
rect 232 252 262 336
rect 328 252 358 336
rect 616 254 646 338
rect 712 254 742 338
<< pmos >>
rect 232 542 262 702
rect 328 542 358 702
rect 616 544 646 704
rect 712 544 742 704
<< ndiff >>
rect 170 324 232 336
rect 170 264 182 324
rect 216 264 232 324
rect 170 252 232 264
rect 262 324 328 336
rect 262 264 278 324
rect 312 264 328 324
rect 262 252 328 264
rect 358 324 420 336
rect 358 264 374 324
rect 408 264 420 324
rect 358 252 420 264
rect 554 326 616 338
rect 554 266 566 326
rect 600 266 616 326
rect 554 254 616 266
rect 646 326 712 338
rect 646 266 662 326
rect 696 266 712 326
rect 646 254 712 266
rect 742 326 804 338
rect 742 266 758 326
rect 792 266 804 326
rect 742 254 804 266
<< pdiff >>
rect 170 690 232 702
rect 170 554 182 690
rect 216 554 232 690
rect 170 542 232 554
rect 262 690 328 702
rect 262 554 278 690
rect 312 554 328 690
rect 262 542 328 554
rect 358 690 420 702
rect 358 554 374 690
rect 408 554 420 690
rect 358 542 420 554
rect 554 692 616 704
rect 554 556 566 692
rect 600 556 616 692
rect 554 544 616 556
rect 646 692 712 704
rect 646 556 662 692
rect 696 556 712 692
rect 646 544 712 556
rect 742 692 804 704
rect 742 556 758 692
rect 792 556 804 692
rect 742 544 804 556
<< ndiffc >>
rect 182 264 216 324
rect 278 264 312 324
rect 374 264 408 324
rect 566 266 600 326
rect 662 266 696 326
rect 758 266 792 326
<< pdiffc >>
rect 182 554 216 690
rect 278 554 312 690
rect 374 554 408 690
rect 566 556 600 692
rect 662 556 696 692
rect 758 556 792 692
<< psubdiff >>
rect 182 148 230 182
rect 264 148 326 182
rect 360 148 430 182
rect 464 148 534 182
rect 568 148 628 182
rect 662 148 726 182
rect 760 148 792 182
<< nsubdiff >>
rect 302 838 806 844
rect 302 804 326 838
rect 360 804 430 838
rect 464 804 534 838
rect 568 804 630 838
rect 664 804 724 838
rect 758 804 806 838
rect 302 798 806 804
<< psubdiffcont >>
rect 230 148 264 182
rect 326 148 360 182
rect 430 148 464 182
rect 534 148 568 182
rect 628 148 662 182
rect 726 148 760 182
<< nsubdiffcont >>
rect 326 804 360 838
rect 430 804 464 838
rect 534 804 568 838
rect 630 804 664 838
rect 724 804 758 838
<< poly >>
rect 212 818 280 828
rect 212 782 228 818
rect 264 782 280 818
rect 212 748 280 782
rect 212 718 358 748
rect 232 702 262 718
rect 328 702 358 718
rect 616 704 646 730
rect 712 704 742 730
rect 232 336 262 542
rect 328 336 358 542
rect 616 430 646 544
rect 410 428 646 430
rect 712 428 742 544
rect 410 418 742 428
rect 410 384 426 418
rect 460 400 742 418
rect 460 384 498 400
rect 410 374 498 384
rect 616 374 742 400
rect 616 338 646 374
rect 712 338 742 374
rect 232 226 262 252
rect 328 226 358 252
rect 616 228 646 254
rect 712 228 742 254
<< polycont >>
rect 228 782 264 818
rect 426 384 460 418
<< locali >>
rect 34 922 148 1004
rect 34 888 48 922
rect 136 888 148 922
rect 34 102 148 888
rect 856 922 970 1004
rect 856 888 868 922
rect 954 888 970 922
rect 856 881 970 888
rect 302 838 806 844
rect 228 818 264 834
rect 302 804 326 838
rect 360 804 430 838
rect 464 804 534 838
rect 568 804 630 838
rect 664 804 724 838
rect 758 804 806 838
rect 302 798 806 804
rect 228 772 264 782
rect 228 738 230 772
rect 182 690 216 706
rect 182 538 216 554
rect 278 690 312 706
rect 182 324 216 340
rect 182 182 216 264
rect 278 334 312 554
rect 374 690 408 798
rect 374 538 408 554
rect 566 692 600 798
rect 566 540 600 556
rect 662 692 696 708
rect 356 418 476 420
rect 356 408 426 418
rect 394 384 426 408
rect 460 384 476 418
rect 394 374 476 384
rect 278 248 312 264
rect 374 324 408 340
rect 374 182 408 264
rect 566 326 600 342
rect 566 182 600 266
rect 662 326 696 556
rect 758 692 792 798
rect 758 540 792 556
rect 662 250 696 266
rect 758 326 792 342
rect 758 182 792 266
rect 182 148 230 182
rect 264 148 326 182
rect 360 148 430 182
rect 464 148 534 182
rect 568 148 628 182
rect 662 148 726 182
rect 760 148 792 182
rect 854 340 970 881
rect 854 292 868 340
rect 956 292 970 340
rect 854 108 970 292
rect 34 68 46 102
rect 136 68 148 102
rect 34 0 148 68
rect 856 102 970 108
rect 856 68 868 102
rect 956 68 970 102
rect 856 0 970 68
<< viali >>
rect 48 888 136 922
rect 868 888 954 922
rect 326 804 360 838
rect 430 804 464 838
rect 534 804 568 838
rect 630 804 664 838
rect 724 804 758 838
rect 230 738 264 772
rect 182 638 216 684
rect 374 638 408 684
rect 662 636 696 691
rect 356 374 394 408
rect 278 324 312 334
rect 278 298 312 324
rect 230 148 264 182
rect 326 148 360 182
rect 430 148 464 182
rect 534 148 568 182
rect 628 148 662 182
rect 726 148 760 182
rect 868 292 956 340
rect 46 68 136 102
rect 868 68 956 102
<< metal1 >>
rect 34 922 148 1004
rect 34 888 48 922
rect 136 888 148 922
rect 34 882 148 888
rect 856 922 970 1004
rect 856 888 868 922
rect 954 888 970 922
rect 856 882 970 888
rect 0 838 1004 854
rect 0 806 326 838
rect 0 798 196 806
rect 298 804 326 806
rect 360 804 430 838
rect 464 804 534 838
rect 568 804 630 838
rect 664 804 724 838
rect 758 804 1004 838
rect 298 798 1004 804
rect 218 772 276 778
rect 218 770 230 772
rect 0 740 230 770
rect 218 738 230 740
rect 264 738 276 772
rect 218 732 276 738
rect 654 740 1004 770
rect 654 691 702 740
rect 170 684 420 690
rect 170 638 182 684
rect 216 638 374 684
rect 408 638 420 684
rect 170 632 420 638
rect 654 636 662 691
rect 696 636 702 691
rect 654 624 702 636
rect 0 568 1004 596
rect 0 512 1004 540
rect 156 458 856 484
rect 0 456 1004 458
rect 0 430 194 456
rect 808 430 1004 456
rect 344 408 406 416
rect 344 402 356 408
rect 0 374 356 402
rect 394 374 406 408
rect 344 364 406 374
rect 488 374 1004 402
rect 270 334 318 346
rect 270 298 278 334
rect 312 322 318 334
rect 488 322 518 374
rect 312 298 518 322
rect 270 286 518 298
rect 854 340 970 346
rect 854 292 868 340
rect 956 292 970 340
rect 854 286 970 292
rect 0 220 1004 258
rect 0 182 1004 192
rect 0 148 230 182
rect 264 148 326 182
rect 360 148 430 182
rect 464 148 534 182
rect 568 148 628 182
rect 662 148 726 182
rect 760 148 1004 182
rect 0 136 1004 148
rect 34 102 148 108
rect 34 68 46 102
rect 136 68 148 102
rect 34 0 148 68
rect 856 102 970 108
rect 856 68 868 102
rect 956 68 970 102
rect 856 0 970 68
<< metal2 >>
rect 32 962 972 972
rect 32 906 42 962
rect 98 906 138 962
rect 194 906 234 962
rect 290 906 330 962
rect 386 906 426 962
rect 482 906 522 962
rect 578 906 618 962
rect 674 906 714 962
rect 770 906 810 962
rect 866 906 906 962
rect 962 906 972 962
rect 32 866 972 906
rect 32 810 42 866
rect 98 810 330 866
rect 386 810 618 866
rect 674 810 906 866
rect 962 810 972 866
rect 32 770 972 810
rect 32 714 42 770
rect 98 714 330 770
rect 386 714 618 770
rect 674 714 906 770
rect 962 714 972 770
rect 32 674 972 714
rect 32 618 42 674
rect 98 618 138 674
rect 194 618 234 674
rect 290 618 330 674
rect 386 618 426 674
rect 482 618 522 674
rect 578 618 618 674
rect 674 618 714 674
rect 770 618 810 674
rect 866 618 906 674
rect 962 618 972 674
rect 32 608 972 618
rect 32 578 396 608
rect 32 522 42 578
rect 98 522 330 578
rect 386 522 396 578
rect 608 578 972 608
rect 32 482 396 522
rect 32 426 42 482
rect 98 426 330 482
rect 386 426 396 482
rect 460 460 544 544
rect 608 522 618 578
rect 674 522 906 578
rect 962 522 972 578
rect 608 482 972 522
rect 32 396 396 426
rect 608 426 618 482
rect 674 426 906 482
rect 962 426 972 482
rect 608 396 972 426
rect 32 386 972 396
rect 32 330 42 386
rect 98 330 138 386
rect 194 330 234 386
rect 290 330 330 386
rect 386 330 426 386
rect 482 330 522 386
rect 578 330 618 386
rect 674 330 714 386
rect 770 330 810 386
rect 866 330 906 386
rect 962 330 972 386
rect 32 290 972 330
rect 32 234 42 290
rect 98 234 330 290
rect 386 234 618 290
rect 674 234 906 290
rect 962 234 972 290
rect 32 194 972 234
rect 32 138 42 194
rect 98 138 330 194
rect 386 138 618 194
rect 674 138 906 194
rect 962 138 972 194
rect 32 98 972 138
rect 32 42 42 98
rect 98 42 138 98
rect 194 42 234 98
rect 290 42 330 98
rect 386 42 426 98
rect 482 42 522 98
rect 578 42 618 98
rect 674 42 714 98
rect 770 42 810 98
rect 866 42 906 98
rect 962 42 972 98
rect 32 32 972 42
<< via2 >>
rect 42 906 98 962
rect 138 906 194 962
rect 234 906 290 962
rect 330 906 386 962
rect 426 906 482 962
rect 522 906 578 962
rect 618 906 674 962
rect 714 906 770 962
rect 810 906 866 962
rect 906 906 962 962
rect 42 810 98 866
rect 330 810 386 866
rect 618 810 674 866
rect 906 810 962 866
rect 42 714 98 770
rect 330 714 386 770
rect 618 714 674 770
rect 906 714 962 770
rect 42 618 98 674
rect 138 618 194 674
rect 234 618 290 674
rect 330 618 386 674
rect 426 618 482 674
rect 522 618 578 674
rect 618 618 674 674
rect 714 618 770 674
rect 810 618 866 674
rect 906 618 962 674
rect 42 522 98 578
rect 330 522 386 578
rect 42 426 98 482
rect 330 426 386 482
rect 618 522 674 578
rect 906 522 962 578
rect 618 426 674 482
rect 906 426 962 482
rect 42 330 98 386
rect 138 330 194 386
rect 234 330 290 386
rect 330 330 386 386
rect 426 330 482 386
rect 522 330 578 386
rect 618 330 674 386
rect 714 330 770 386
rect 810 330 866 386
rect 906 330 962 386
rect 42 234 98 290
rect 330 234 386 290
rect 618 234 674 290
rect 906 234 962 290
rect 42 138 98 194
rect 330 138 386 194
rect 618 138 674 194
rect 906 138 962 194
rect 42 42 98 98
rect 138 42 194 98
rect 234 42 290 98
rect 330 42 386 98
rect 426 42 482 98
rect 522 42 578 98
rect 618 42 674 98
rect 714 42 770 98
rect 810 42 866 98
rect 906 42 962 98
<< metal3 >>
rect 36 962 968 968
rect 36 906 42 962
rect 98 906 138 962
rect 194 906 234 962
rect 290 906 330 962
rect 386 906 426 962
rect 482 906 522 962
rect 578 906 618 962
rect 674 906 714 962
rect 770 906 810 962
rect 866 906 906 962
rect 962 906 968 962
rect 36 900 968 906
rect 36 866 104 900
rect 36 810 42 866
rect 98 810 104 866
rect 324 866 392 900
rect 36 770 104 810
rect 36 714 42 770
rect 98 714 104 770
rect 164 824 264 840
rect 164 756 180 824
rect 248 756 264 824
rect 164 740 264 756
rect 324 810 330 866
rect 386 810 392 866
rect 612 866 680 900
rect 324 770 392 810
rect 36 680 104 714
rect 324 714 330 770
rect 386 714 392 770
rect 452 824 552 840
rect 452 756 468 824
rect 536 756 552 824
rect 452 740 552 756
rect 612 810 618 866
rect 674 810 680 866
rect 900 866 968 900
rect 612 770 680 810
rect 324 680 392 714
rect 612 714 618 770
rect 674 714 680 770
rect 740 824 840 840
rect 740 756 756 824
rect 824 756 840 824
rect 740 740 840 756
rect 900 810 906 866
rect 962 810 968 866
rect 900 770 968 810
rect 612 680 680 714
rect 900 714 906 770
rect 962 714 968 770
rect 900 680 968 714
rect 36 674 968 680
rect 36 618 42 674
rect 98 618 138 674
rect 194 618 234 674
rect 290 618 330 674
rect 386 618 426 674
rect 482 618 522 674
rect 578 618 618 674
rect 674 618 714 674
rect 770 618 810 674
rect 866 618 906 674
rect 962 618 968 674
rect 36 612 968 618
rect 36 578 104 612
rect 36 522 42 578
rect 98 522 104 578
rect 324 578 392 612
rect 36 482 104 522
rect 36 426 42 482
rect 98 426 104 482
rect 164 536 264 552
rect 164 468 180 536
rect 248 468 264 536
rect 164 452 264 468
rect 324 522 330 578
rect 386 522 392 578
rect 324 482 392 522
rect 36 392 104 426
rect 324 426 330 482
rect 386 426 392 482
rect 324 392 392 426
rect 612 578 680 612
rect 612 522 618 578
rect 674 522 680 578
rect 900 578 968 612
rect 612 482 680 522
rect 612 426 618 482
rect 674 426 680 482
rect 740 536 840 552
rect 740 468 756 536
rect 824 468 840 536
rect 740 452 840 468
rect 900 522 906 578
rect 962 522 968 578
rect 900 482 968 522
rect 612 392 680 426
rect 900 426 906 482
rect 962 426 968 482
rect 900 392 968 426
rect 36 386 968 392
rect 36 330 42 386
rect 98 330 138 386
rect 194 330 234 386
rect 290 330 330 386
rect 386 330 426 386
rect 482 330 522 386
rect 578 330 618 386
rect 674 330 714 386
rect 770 330 810 386
rect 866 330 906 386
rect 962 330 968 386
rect 36 324 968 330
rect 36 290 104 324
rect 36 234 42 290
rect 98 234 104 290
rect 324 290 392 324
rect 36 194 104 234
rect 36 138 42 194
rect 98 138 104 194
rect 164 248 264 264
rect 164 180 180 248
rect 248 180 264 248
rect 164 164 264 180
rect 324 234 330 290
rect 386 234 392 290
rect 612 290 680 324
rect 324 194 392 234
rect 36 104 104 138
rect 324 138 330 194
rect 386 138 392 194
rect 452 248 552 264
rect 452 180 468 248
rect 536 180 552 248
rect 452 164 552 180
rect 612 234 618 290
rect 674 234 680 290
rect 900 290 968 324
rect 612 194 680 234
rect 324 104 392 138
rect 612 138 618 194
rect 674 138 680 194
rect 740 248 840 264
rect 740 180 756 248
rect 824 180 840 248
rect 740 164 840 180
rect 900 234 906 290
rect 962 234 968 290
rect 900 194 968 234
rect 612 104 680 138
rect 900 138 906 194
rect 962 138 968 194
rect 900 104 968 138
rect 36 98 968 104
rect 36 42 42 98
rect 98 42 138 98
rect 194 42 234 98
rect 290 42 330 98
rect 386 42 426 98
rect 482 42 522 98
rect 578 42 618 98
rect 674 42 714 98
rect 770 42 810 98
rect 866 42 906 98
rect 962 42 968 98
rect 36 36 968 42
<< via3 >>
rect 180 756 248 824
rect 468 756 536 824
rect 756 756 824 824
rect 180 468 248 536
rect 756 468 824 536
rect 180 180 248 248
rect 468 180 536 248
rect 756 180 824 248
<< metal4 >>
rect 184 840 244 934
rect 472 840 532 934
rect 760 840 820 934
rect 164 824 264 840
rect 164 820 180 824
rect 70 760 180 820
rect 164 756 180 760
rect 248 820 264 824
rect 452 824 552 840
rect 452 820 468 824
rect 248 760 468 820
rect 248 756 264 760
rect 164 740 264 756
rect 452 756 468 760
rect 536 820 552 824
rect 740 824 840 840
rect 740 820 756 824
rect 536 760 756 820
rect 536 756 552 760
rect 452 740 552 756
rect 740 756 756 760
rect 824 820 840 824
rect 824 760 934 820
rect 824 756 840 760
rect 740 740 840 756
rect 184 552 244 740
rect 472 646 532 740
rect 760 552 820 740
rect 164 536 264 552
rect 164 532 180 536
rect 70 472 180 532
rect 164 468 180 472
rect 248 532 264 536
rect 740 536 840 552
rect 740 532 756 536
rect 248 472 358 532
rect 646 472 756 532
rect 248 468 264 472
rect 164 452 264 468
rect 740 468 756 472
rect 824 532 840 536
rect 824 472 934 532
rect 824 468 840 472
rect 740 452 840 468
rect 184 264 244 452
rect 472 264 532 358
rect 760 264 820 452
rect 164 248 264 264
rect 164 244 180 248
rect 70 184 180 244
rect 164 180 180 184
rect 248 244 264 248
rect 452 248 552 264
rect 452 244 468 248
rect 248 184 468 244
rect 248 180 264 184
rect 164 164 264 180
rect 452 180 468 184
rect 536 244 552 248
rect 740 248 840 264
rect 740 244 756 248
rect 536 184 756 244
rect 536 180 552 184
rect 452 164 552 180
rect 740 180 756 184
rect 824 244 840 248
rect 824 184 934 244
rect 824 180 840 184
rect 740 164 840 180
rect 184 70 244 164
rect 472 70 532 164
rect 760 70 820 164
<< comment >>
rect 0 972 32 1004
rect 972 972 1004 1004
rect 138 750 308 798
rect 430 756 562 804
rect 138 260 194 750
rect 312 690 368 750
rect 358 428 406 688
rect 430 562 478 756
rect 564 716 606 762
rect 598 608 632 716
rect 576 604 632 608
rect 558 602 632 604
rect 558 576 608 602
rect 544 562 600 576
rect 430 558 600 562
rect 430 544 576 558
rect 430 514 558 544
rect 430 460 478 514
rect 560 478 602 522
rect 560 476 636 478
rect 428 428 478 460
rect 358 396 428 428
rect 300 260 356 318
rect 358 314 406 396
rect 138 258 356 260
rect 138 212 306 258
rect 430 206 478 428
rect 602 198 636 476
rect 670 198 716 802
rect 0 0 32 32
rect 972 0 1004 32
<< labels >>
flabel metal1 0 798 167 854 0 FreeSans 160 0 0 0 VDD
port 1 w power bidirectional
flabel metal1 837 798 1004 854 0 FreeSans 160 0 0 0 VDD
port 1 e power bidirectional
flabel metal1 0 136 1004 192 0 FreeSans 320 0 0 0 VSS
port 2 nsew ground bidirectional
flabel metal1 0 220 1004 258 0 FreeSans 320 0 0 0 vcom
port 3 nsew
flabel metal4 472 874 532 934 1 FreeSans 160 0 0 0 ctop
port 4 n
flabel metal1 34 0 148 108 5 FreeSans 320 0 0 0 col
port 5 s
flabel metal1 34 882 148 1004 1 FreeSans 320 0 0 0 col
port 5 n
flabel metal1 856 0 970 108 1 FreeSans 320 0 0 0 col_n
port 6 s
flabel metal1 856 882 970 1004 1 FreeSans 320 0 0 0 col_n
port 6 n
flabel metal1 0 430 158 458 0 FreeSans 160 0 0 0 row_n
port 7 w
flabel metal1 846 430 1004 458 0 FreeSans 160 0 0 0 row_n
port 7 e
flabel metal1 0 512 155 540 0 FreeSans 160 0 0 0 rowon_n
port 8 w
flabel metal1 849 512 1004 540 0 FreeSans 160 0 0 0 rowon_n
port 8 e
flabel metal1 0 374 158 402 0 FreeSans 160 0 0 0 sample_i
port 9 w
flabel metal1 846 374 1004 402 0 FreeSans 160 0 0 0 sample_o
port 10 e
flabel metal1 0 740 158 770 0 FreeSans 160 0 0 0 sample_n_i
port 11 nsew
flabel metal1 846 740 1004 770 0 FreeSans 160 0 0 0 sample_n_o
port 12 nsew
flabel metal1 0 568 156 596 7 FreeSans 160 0 0 0 off_n
port 13 w
flabel metal1 848 568 1004 596 3 FreeSans 160 0 0 0 off_n
port 13 e
rlabel metal2 500 972 500 972 1 cbot
<< end >>
