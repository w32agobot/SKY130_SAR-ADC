MACRO sky130_mm_sc_hd_dlyPoly5ns
  CLASS CORE ;
  FOREIGN sky130_mm_sc_hd_dlyPoly5ns ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.500 BY 2.720 ;
  SITE unithd ;
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.635 11.500 2.805 ;
        RECT 0.195 2.000 0.365 2.235 ;
        RECT 0.190 1.805 0.365 2.000 ;
        RECT 8.515 1.625 8.685 2.635 ;
        RECT 9.815 1.480 9.985 2.635 ;
        RECT 9.815 1.310 10.395 1.480 ;
        RECT 10.225 0.345 10.395 1.310 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 11.185 2.635 11.355 2.805 ;
        RECT 0.195 1.895 0.365 2.155 ;
      LAYER met1 ;
        RECT 0.000 2.480 11.500 2.960 ;
        RECT 0.165 1.810 0.395 2.480 ;
        RECT 0.190 1.805 0.365 1.810 ;
    END
  END VPWR
  PIN in
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.672600 ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.215 0.375 1.320 ;
        RECT 0.105 1.045 4.925 1.215 ;
        RECT 0.105 0.990 0.375 1.045 ;
    END
  END in
  PIN out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.366000 ;
    ANTENNADIFFAREA 0.361800 ;
    PORT
      LAYER li1 ;
        RECT 9.475 1.140 9.645 2.455 ;
        RECT 10.570 1.155 10.905 1.325 ;
        RECT 9.475 1.050 9.910 1.140 ;
        RECT 9.180 0.965 9.910 1.050 ;
        RECT 10.675 0.965 10.905 1.155 ;
        RECT 9.180 0.880 9.645 0.965 ;
        RECT 9.180 0.345 9.350 0.880 ;
    END
  END out
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 5.130 1.680 5.300 1.750 ;
        RECT 7.670 1.680 7.840 1.755 ;
        RECT 0.195 0.455 0.365 0.790 ;
        RECT 4.745 0.085 4.915 0.090 ;
        RECT 5.120 0.085 7.840 1.680 ;
        RECT 8.170 1.340 8.340 1.565 ;
        RECT 10.665 1.545 10.835 2.455 ;
        RECT 8.170 1.175 8.390 1.340 ;
        RECT 8.220 0.085 8.390 1.175 ;
        RECT 0.000 -0.085 11.500 0.085 ;
      LAYER mcon ;
        RECT 0.195 0.535 0.365 0.710 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.090 ;
        RECT 10.665 1.705 10.835 1.945 ;
        RECT 8.170 1.395 8.340 1.565 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
        RECT 11.185 -0.085 11.355 0.085 ;
      LAYER met1 ;
        RECT 8.110 1.570 8.370 1.600 ;
        RECT 10.635 1.570 10.865 2.010 ;
        RECT 8.110 1.375 10.865 1.570 ;
        RECT 8.110 1.365 8.370 1.375 ;
        RECT 0.165 0.240 0.395 0.775 ;
        RECT 0.000 -0.240 11.500 0.240 ;
    END
  END VGND
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 2.070 11.690 2.910 ;
        RECT -0.190 1.235 4.730 2.070 ;
        RECT 8.240 1.235 11.690 2.070 ;
    END
  END VPB
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 4.730 1.070 8.240 2.070 ;
        RECT 0.005 -0.085 11.495 1.070 ;
    END
  END VNB
  OBS
      LAYER li1 ;
        RECT 4.315 1.445 4.485 2.235 ;
        RECT 5.475 1.870 7.495 2.125 ;
        RECT 8.995 1.625 9.165 2.455 ;
        RECT 10.155 1.915 10.355 2.455 ;
        RECT 11.145 1.625 11.345 2.455 ;
        RECT 8.560 1.010 8.915 1.180 ;
        RECT 4.315 0.365 4.485 0.875 ;
        RECT 8.700 0.345 8.870 0.795 ;
        RECT 9.745 0.345 9.915 0.715 ;
        RECT 10.705 0.345 10.875 0.795 ;
      LAYER mcon ;
        RECT 4.315 1.525 4.485 2.085 ;
        RECT 6.140 1.920 6.320 2.090 ;
        RECT 6.630 1.920 6.810 2.090 ;
        RECT 8.995 1.770 9.165 2.225 ;
        RECT 10.185 2.060 10.355 2.255 ;
        RECT 11.145 1.805 11.315 2.215 ;
        RECT 8.615 1.010 8.835 1.180 ;
        RECT 4.315 0.535 4.485 0.715 ;
        RECT 8.700 0.525 8.870 0.715 ;
        RECT 9.745 0.495 9.915 0.665 ;
        RECT 10.705 0.525 10.875 0.695 ;
      LAYER met1 ;
        RECT 4.285 1.580 4.515 2.195 ;
        RECT 8.965 2.150 11.345 2.290 ;
        RECT 6.080 1.890 6.870 2.120 ;
        RECT 6.365 1.680 6.590 1.890 ;
        RECT 8.965 1.710 9.195 2.150 ;
        RECT 10.155 2.000 10.385 2.150 ;
        RECT 11.115 1.745 11.345 2.150 ;
        RECT 5.050 1.580 7.940 1.680 ;
        RECT 4.285 1.425 7.940 1.580 ;
        RECT 4.910 1.115 7.940 1.425 ;
        RECT 8.465 1.115 8.915 1.210 ;
        RECT 4.910 0.920 8.915 1.115 ;
        RECT 4.910 0.785 7.940 0.920 ;
        RECT 4.280 0.475 7.940 0.785 ;
        RECT 5.050 0.465 7.940 0.475 ;
        RECT 8.670 0.605 8.900 0.775 ;
        RECT 9.685 0.605 9.975 0.695 ;
        RECT 10.645 0.605 10.935 0.735 ;
        RECT 8.670 0.565 10.935 0.605 ;
        RECT 8.670 0.465 10.905 0.565 ;
  END
END sky130_mm_sc_hd_dlyPoly5ns
END LIBRARY

