* SPICE3 file created from adc_array_wafflecap_16(1)x300aF_28um2.ext - technology: sky130A

.subckt adc_array_wafflecap_16(1)x300aF_28um2 cbot ctop
C0 cbot ctop 0.30fF
C1 cfloating cbot 4.40fF
C2 cfloating ctop 0.60fF
C3 cbot VSUBS 2.17fF
C4 cfloating VSUBS 0.71fF
.ends
