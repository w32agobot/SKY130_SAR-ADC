VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO adc_comp_latch
  CLASS BLOCK ;
  FOREIGN adc_comp_latch ;
  ORIGIN 0.000 0.000 ;
  SIZE 42.000 BY 129.000 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 38.730 50.000 40.330 77.980 ;
    END
    PORT
      LAYER met4 ;
        RECT 8.240 50.000 9.840 77.980 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 36.780 50.000 38.380 77.980 ;
    END
    PORT
      LAYER met4 ;
        RECT 10.220 50.000 11.820 77.980 ;
    END
  END VSS
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 8.010 61.890 13.390 62.030 ;
    END
  END clk
  PIN inp
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 8.010 65.410 18.920 65.550 ;
    END
  END inp
  PIN inn
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 8.010 65.130 16.960 65.270 ;
    END
  END inn
  PIN comp_trig
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 34.520 62.590 40.330 62.730 ;
    END
  END comp_trig
  PIN latch_qn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 35.320 65.540 40.330 65.680 ;
    END
  END latch_qn
  PIN latch_q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 34.000 65.880 40.330 66.020 ;
    END
  END latch_q
  OBS
      LAYER li1 ;
        RECT 12.150 50.000 36.540 77.980 ;
      LAYER met1 ;
        RECT 8.010 66.300 40.330 76.890 ;
        RECT 8.010 65.830 33.720 66.300 ;
        RECT 19.200 65.600 33.720 65.830 ;
        RECT 19.200 65.260 35.040 65.600 ;
        RECT 19.200 65.130 40.330 65.260 ;
        RECT 17.240 64.850 40.330 65.130 ;
        RECT 8.010 63.010 40.330 64.850 ;
        RECT 8.010 62.310 34.240 63.010 ;
        RECT 13.670 61.610 40.330 62.310 ;
        RECT 8.010 51.040 40.330 61.610 ;
      LAYER met2 ;
        RECT 8.240 51.040 40.330 76.890 ;
      LAYER met3 ;
        RECT 8.240 51.040 40.330 76.890 ;
      LAYER met4 ;
        RECT 12.220 51.040 35.030 76.890 ;
  END
END adc_comp_latch
END LIBRARY

