magic
tech sky130A
magscale 1 2
timestamp 1663595907
<< nwell >>
rect 3118 6400 4700 6404
rect 760 5996 4700 6400
rect 760 5978 3052 5996
rect 1286 5976 1528 5978
rect 1894 5628 3052 5978
rect 3690 5948 4700 5996
rect 288 5210 730 5608
rect 3850 5256 4364 5308
rect 3154 4852 4364 5256
<< pwell >>
rect 906 7994 1386 8174
rect 3486 7994 3966 8174
rect 446 7914 1696 7994
rect 2346 7914 2526 7994
rect 3176 7914 4426 7994
rect 446 6854 4426 7914
rect 446 6774 1696 6854
rect 2346 6774 2526 6854
rect 3176 6774 4426 6854
rect 906 6594 1386 6774
rect 3486 6594 3966 6774
rect 906 4404 1386 4584
rect 3486 4404 3966 4584
rect 446 4324 1696 4404
rect 2346 4324 2526 4404
rect 3176 4324 4426 4404
rect 446 3264 4426 4324
rect 446 3184 1696 3264
rect 2346 3184 2526 3264
rect 3176 3184 4426 3264
rect 906 3004 1386 3184
rect 3486 3004 3966 3184
<< nmos >>
rect 596 6994 4276 7774
rect 3252 5732 3282 5832
rect 3348 5732 3378 5832
rect 3444 5732 3474 5832
rect 3788 5796 3818 5880
rect 3884 5796 3914 5880
rect 4284 5796 4314 5880
rect 4380 5796 4410 5880
rect 860 5264 890 5664
rect 956 5264 986 5664
rect 1052 5264 1082 5664
rect 1148 5264 1178 5664
rect 1244 5264 1274 5664
rect 1340 5264 1370 5664
rect 1436 5264 1466 5664
rect 1532 5264 1562 5664
rect 350 5054 434 5084
rect 584 5054 668 5084
rect 860 5004 890 5104
rect 956 5004 986 5104
rect 1052 5004 1082 5104
rect 1148 5004 1178 5104
rect 1244 5004 1274 5104
rect 1340 5004 1370 5104
rect 1436 5004 1466 5104
rect 1532 5004 1562 5104
rect 2314 4998 2344 5398
rect 2410 4998 2440 5398
rect 2506 4998 2536 5398
rect 2602 4998 2632 5398
rect 3252 5420 3282 5520
rect 3348 5420 3378 5520
rect 3444 5420 3474 5520
rect 3948 5376 3978 5460
rect 4044 5376 4074 5460
rect 596 3404 4276 4184
<< pmos >>
rect 860 6078 890 6178
rect 956 6078 986 6178
rect 1052 6078 1082 6178
rect 1148 6078 1178 6178
rect 1244 6078 1274 6178
rect 1340 6078 1370 6178
rect 1436 6078 1466 6178
rect 1532 6078 1562 6178
rect 1992 5728 2022 6128
rect 2088 5728 2118 6128
rect 2314 5728 2344 6128
rect 2410 5728 2440 6128
rect 2506 5728 2536 6128
rect 2602 5728 2632 6128
rect 2828 5728 2858 6128
rect 2924 5728 2954 6128
rect 3252 6058 3282 6258
rect 3348 6058 3378 6258
rect 3444 6058 3474 6258
rect 3788 6050 3818 6210
rect 3884 6050 3914 6210
rect 3980 6050 4010 6210
rect 4076 6050 4106 6210
rect 4284 6050 4314 6210
rect 4380 6050 4410 6210
rect 4476 6050 4506 6210
rect 4572 6050 4602 6210
rect 350 5396 438 5426
rect 584 5396 672 5426
rect 350 5304 438 5334
rect 584 5304 672 5334
rect 3252 4994 3282 5194
rect 3348 4994 3378 5194
rect 3444 4994 3474 5194
rect 3948 5046 3978 5206
rect 4044 5046 4074 5206
rect 4140 5046 4170 5206
rect 4236 5046 4266 5206
<< ndiff >>
rect 596 7894 4276 7914
rect 596 7794 606 7894
rect 726 7794 766 7894
rect 886 7794 926 7894
rect 1046 7794 1086 7894
rect 1206 7794 1246 7894
rect 1366 7794 1406 7894
rect 1526 7794 1566 7894
rect 1686 7794 3186 7894
rect 3306 7794 3346 7894
rect 3466 7794 3506 7894
rect 3626 7794 3666 7894
rect 3786 7794 3826 7894
rect 3946 7794 3986 7894
rect 4106 7794 4146 7894
rect 4266 7794 4276 7894
rect 596 7774 4276 7794
rect 596 6974 4276 6994
rect 596 6874 606 6974
rect 726 6874 766 6974
rect 886 6874 926 6974
rect 1046 6874 1086 6974
rect 1206 6874 1246 6974
rect 1366 6874 1406 6974
rect 1526 6874 1566 6974
rect 1686 6874 3186 6974
rect 3306 6874 3346 6974
rect 3466 6874 3506 6974
rect 3626 6874 3666 6974
rect 3786 6874 3826 6974
rect 3946 6874 3986 6974
rect 4106 6874 4146 6974
rect 4266 6874 4276 6974
rect 596 6854 4276 6874
rect 3190 5820 3252 5832
rect 3190 5744 3202 5820
rect 3236 5744 3252 5820
rect 3190 5732 3252 5744
rect 3282 5820 3348 5832
rect 3282 5744 3298 5820
rect 3332 5744 3348 5820
rect 3282 5732 3348 5744
rect 3378 5820 3444 5832
rect 3378 5744 3394 5820
rect 3428 5744 3444 5820
rect 3378 5732 3444 5744
rect 3474 5820 3536 5832
rect 3474 5744 3490 5820
rect 3524 5744 3536 5820
rect 3474 5732 3536 5744
rect 3726 5868 3788 5880
rect 3726 5808 3738 5868
rect 3772 5808 3788 5868
rect 3726 5796 3788 5808
rect 3818 5868 3884 5880
rect 3818 5808 3834 5868
rect 3868 5808 3884 5868
rect 3818 5796 3884 5808
rect 3914 5868 3976 5880
rect 3914 5808 3930 5868
rect 3964 5808 3976 5868
rect 3914 5796 3976 5808
rect 4222 5868 4284 5880
rect 4222 5808 4234 5868
rect 4268 5808 4284 5868
rect 4222 5796 4284 5808
rect 4314 5868 4380 5880
rect 4314 5808 4330 5868
rect 4364 5808 4380 5868
rect 4314 5796 4380 5808
rect 4410 5868 4472 5880
rect 4410 5808 4426 5868
rect 4460 5808 4472 5868
rect 4410 5796 4472 5808
rect 798 5652 860 5664
rect 798 5276 810 5652
rect 844 5276 860 5652
rect 798 5264 860 5276
rect 890 5652 956 5664
rect 890 5276 906 5652
rect 940 5276 956 5652
rect 890 5264 956 5276
rect 986 5652 1052 5664
rect 986 5276 1002 5652
rect 1036 5276 1052 5652
rect 986 5264 1052 5276
rect 1082 5652 1148 5664
rect 1082 5276 1098 5652
rect 1132 5276 1148 5652
rect 1082 5264 1148 5276
rect 1178 5652 1244 5664
rect 1178 5276 1194 5652
rect 1228 5276 1244 5652
rect 1178 5264 1244 5276
rect 1274 5652 1340 5664
rect 1274 5276 1290 5652
rect 1324 5276 1340 5652
rect 1274 5264 1340 5276
rect 1370 5652 1436 5664
rect 1370 5276 1386 5652
rect 1420 5276 1436 5652
rect 1370 5264 1436 5276
rect 1466 5652 1532 5664
rect 1466 5276 1482 5652
rect 1516 5276 1532 5652
rect 1466 5264 1532 5276
rect 1562 5652 1624 5664
rect 1562 5276 1578 5652
rect 1612 5276 1624 5652
rect 1562 5264 1624 5276
rect 2252 5386 2314 5398
rect 350 5130 434 5142
rect 350 5096 362 5130
rect 422 5096 434 5130
rect 350 5084 434 5096
rect 584 5130 668 5142
rect 584 5096 596 5130
rect 656 5096 668 5130
rect 584 5084 668 5096
rect 798 5092 860 5104
rect 350 5042 434 5054
rect 350 5008 362 5042
rect 422 5008 434 5042
rect 350 4996 434 5008
rect 584 5042 668 5054
rect 584 5008 596 5042
rect 656 5008 668 5042
rect 584 4996 668 5008
rect 798 5016 810 5092
rect 844 5016 860 5092
rect 798 5004 860 5016
rect 890 5092 956 5104
rect 890 5016 906 5092
rect 940 5016 956 5092
rect 890 5004 956 5016
rect 986 5092 1052 5104
rect 986 5016 1002 5092
rect 1036 5016 1052 5092
rect 986 5004 1052 5016
rect 1082 5092 1148 5104
rect 1082 5016 1098 5092
rect 1132 5016 1148 5092
rect 1082 5004 1148 5016
rect 1178 5092 1244 5104
rect 1178 5016 1194 5092
rect 1228 5016 1244 5092
rect 1178 5004 1244 5016
rect 1274 5092 1340 5104
rect 1274 5016 1290 5092
rect 1324 5016 1340 5092
rect 1274 5004 1340 5016
rect 1370 5092 1436 5104
rect 1370 5016 1386 5092
rect 1420 5016 1436 5092
rect 1370 5004 1436 5016
rect 1466 5092 1532 5104
rect 1466 5016 1482 5092
rect 1516 5016 1532 5092
rect 1466 5004 1532 5016
rect 1562 5092 1624 5104
rect 1562 5016 1578 5092
rect 1612 5016 1624 5092
rect 1562 5004 1624 5016
rect 2252 5010 2264 5386
rect 2298 5010 2314 5386
rect 2252 4998 2314 5010
rect 2344 5386 2410 5398
rect 2344 5010 2360 5386
rect 2394 5010 2410 5386
rect 2344 4998 2410 5010
rect 2440 5386 2506 5398
rect 2440 5010 2456 5386
rect 2490 5010 2506 5386
rect 2440 4998 2506 5010
rect 2536 5386 2602 5398
rect 2536 5010 2552 5386
rect 2586 5010 2602 5386
rect 2536 4998 2602 5010
rect 2632 5386 2694 5398
rect 2632 5010 2648 5386
rect 2682 5010 2694 5386
rect 3190 5508 3252 5520
rect 3190 5432 3202 5508
rect 3236 5432 3252 5508
rect 3190 5420 3252 5432
rect 3282 5508 3348 5520
rect 3282 5432 3298 5508
rect 3332 5432 3348 5508
rect 3282 5420 3348 5432
rect 3378 5508 3444 5520
rect 3378 5432 3394 5508
rect 3428 5432 3444 5508
rect 3378 5420 3444 5432
rect 3474 5508 3536 5520
rect 3474 5432 3490 5508
rect 3524 5432 3536 5508
rect 3474 5420 3536 5432
rect 3886 5448 3948 5460
rect 3886 5388 3898 5448
rect 3932 5388 3948 5448
rect 3886 5376 3948 5388
rect 3978 5448 4044 5460
rect 3978 5388 3994 5448
rect 4028 5388 4044 5448
rect 3978 5376 4044 5388
rect 4074 5448 4136 5460
rect 4074 5388 4090 5448
rect 4124 5388 4136 5448
rect 4074 5376 4136 5388
rect 2632 4998 2694 5010
rect 596 4304 4276 4324
rect 596 4204 606 4304
rect 726 4204 766 4304
rect 886 4204 926 4304
rect 1046 4204 1086 4304
rect 1206 4204 1246 4304
rect 1366 4204 1406 4304
rect 1526 4204 1566 4304
rect 1686 4204 3186 4304
rect 3306 4204 3346 4304
rect 3466 4204 3506 4304
rect 3626 4204 3666 4304
rect 3786 4204 3826 4304
rect 3946 4204 3986 4304
rect 4106 4204 4146 4304
rect 4266 4204 4276 4304
rect 596 4184 4276 4204
rect 596 3384 4276 3404
rect 596 3284 606 3384
rect 726 3284 766 3384
rect 886 3284 926 3384
rect 1046 3284 1086 3384
rect 1206 3284 1246 3384
rect 1366 3284 1406 3384
rect 1526 3284 1566 3384
rect 1686 3284 3186 3384
rect 3306 3284 3346 3384
rect 3466 3284 3506 3384
rect 3626 3284 3666 3384
rect 3786 3284 3826 3384
rect 3946 3284 3986 3384
rect 4106 3284 4146 3384
rect 4266 3284 4276 3384
rect 596 3264 4276 3284
<< pdiff >>
rect 3190 6246 3252 6258
rect 798 6166 860 6178
rect 798 6090 810 6166
rect 844 6090 860 6166
rect 798 6078 860 6090
rect 890 6166 956 6178
rect 890 6090 906 6166
rect 940 6090 956 6166
rect 890 6078 956 6090
rect 986 6166 1052 6178
rect 986 6090 1002 6166
rect 1036 6090 1052 6166
rect 986 6078 1052 6090
rect 1082 6166 1148 6178
rect 1082 6090 1098 6166
rect 1132 6090 1148 6166
rect 1082 6078 1148 6090
rect 1178 6166 1244 6178
rect 1178 6090 1194 6166
rect 1228 6090 1244 6166
rect 1178 6078 1244 6090
rect 1274 6166 1340 6178
rect 1274 6090 1290 6166
rect 1324 6090 1340 6166
rect 1274 6078 1340 6090
rect 1370 6166 1436 6178
rect 1370 6090 1386 6166
rect 1420 6090 1436 6166
rect 1370 6078 1436 6090
rect 1466 6166 1532 6178
rect 1466 6090 1482 6166
rect 1516 6090 1532 6166
rect 1466 6078 1532 6090
rect 1562 6166 1624 6178
rect 1562 6090 1578 6166
rect 1612 6090 1624 6166
rect 1562 6078 1624 6090
rect 1930 6116 1992 6128
rect 1930 5740 1942 6116
rect 1976 5740 1992 6116
rect 1930 5728 1992 5740
rect 2022 6116 2088 6128
rect 2022 5740 2038 6116
rect 2072 5740 2088 6116
rect 2022 5728 2088 5740
rect 2118 6116 2180 6128
rect 2118 5740 2134 6116
rect 2168 5740 2180 6116
rect 2118 5728 2180 5740
rect 2252 6116 2314 6128
rect 2252 5740 2264 6116
rect 2298 5740 2314 6116
rect 2252 5728 2314 5740
rect 2344 6116 2410 6128
rect 2344 5740 2360 6116
rect 2394 5740 2410 6116
rect 2344 5728 2410 5740
rect 2440 6116 2506 6128
rect 2440 5740 2456 6116
rect 2490 5740 2506 6116
rect 2440 5728 2506 5740
rect 2536 6116 2602 6128
rect 2536 5740 2552 6116
rect 2586 5740 2602 6116
rect 2536 5728 2602 5740
rect 2632 6116 2694 6128
rect 2632 5740 2648 6116
rect 2682 5740 2694 6116
rect 2632 5728 2694 5740
rect 2766 6116 2828 6128
rect 2766 5740 2778 6116
rect 2812 5740 2828 6116
rect 2766 5728 2828 5740
rect 2858 6116 2924 6128
rect 2858 5740 2874 6116
rect 2908 5740 2924 6116
rect 2858 5728 2924 5740
rect 2954 6116 3016 6128
rect 2954 5740 2970 6116
rect 3004 5740 3016 6116
rect 3190 6070 3202 6246
rect 3236 6070 3252 6246
rect 3190 6058 3252 6070
rect 3282 6246 3348 6258
rect 3282 6070 3298 6246
rect 3332 6070 3348 6246
rect 3282 6058 3348 6070
rect 3378 6246 3444 6258
rect 3378 6070 3394 6246
rect 3428 6070 3444 6246
rect 3378 6058 3444 6070
rect 3474 6246 3536 6258
rect 3474 6070 3490 6246
rect 3524 6070 3536 6246
rect 3474 6058 3536 6070
rect 3726 6198 3788 6210
rect 3726 6062 3738 6198
rect 3772 6062 3788 6198
rect 3726 6050 3788 6062
rect 3818 6198 3884 6210
rect 3818 6062 3834 6198
rect 3868 6062 3884 6198
rect 3818 6050 3884 6062
rect 3914 6198 3980 6210
rect 3914 6062 3930 6198
rect 3964 6062 3980 6198
rect 3914 6050 3980 6062
rect 4010 6198 4076 6210
rect 4010 6062 4026 6198
rect 4060 6062 4076 6198
rect 4010 6050 4076 6062
rect 4106 6198 4168 6210
rect 4106 6062 4122 6198
rect 4156 6062 4168 6198
rect 4106 6050 4168 6062
rect 4222 6198 4284 6210
rect 4222 6062 4234 6198
rect 4268 6062 4284 6198
rect 4222 6050 4284 6062
rect 4314 6198 4380 6210
rect 4314 6062 4330 6198
rect 4364 6062 4380 6198
rect 4314 6050 4380 6062
rect 4410 6198 4476 6210
rect 4410 6062 4426 6198
rect 4460 6062 4476 6198
rect 4410 6050 4476 6062
rect 4506 6198 4572 6210
rect 4506 6062 4522 6198
rect 4556 6062 4572 6198
rect 4506 6050 4572 6062
rect 4602 6198 4664 6210
rect 4602 6062 4618 6198
rect 4652 6062 4664 6198
rect 4602 6050 4664 6062
rect 2954 5728 3016 5740
rect 350 5474 438 5482
rect 350 5440 362 5474
rect 422 5440 438 5474
rect 350 5426 438 5440
rect 584 5474 672 5482
rect 584 5440 596 5474
rect 656 5440 672 5474
rect 584 5426 672 5440
rect 350 5382 438 5396
rect 350 5348 362 5382
rect 422 5348 438 5382
rect 350 5334 438 5348
rect 584 5382 672 5396
rect 584 5348 596 5382
rect 656 5348 672 5382
rect 584 5334 672 5348
rect 350 5292 438 5304
rect 350 5258 362 5292
rect 422 5258 438 5292
rect 350 5246 438 5258
rect 584 5292 672 5304
rect 584 5258 596 5292
rect 656 5258 672 5292
rect 584 5246 672 5258
rect 3886 5194 3948 5206
rect 3190 5182 3252 5194
rect 3190 5006 3202 5182
rect 3236 5006 3252 5182
rect 3190 4994 3252 5006
rect 3282 5182 3348 5194
rect 3282 5006 3298 5182
rect 3332 5006 3348 5182
rect 3282 4994 3348 5006
rect 3378 5182 3444 5194
rect 3378 5006 3394 5182
rect 3428 5006 3444 5182
rect 3378 4994 3444 5006
rect 3474 5182 3536 5194
rect 3474 5006 3490 5182
rect 3524 5006 3536 5182
rect 3886 5058 3898 5194
rect 3932 5058 3948 5194
rect 3886 5046 3948 5058
rect 3978 5194 4044 5206
rect 3978 5058 3994 5194
rect 4028 5058 4044 5194
rect 3978 5046 4044 5058
rect 4074 5194 4140 5206
rect 4074 5058 4090 5194
rect 4124 5058 4140 5194
rect 4074 5046 4140 5058
rect 4170 5194 4236 5206
rect 4170 5058 4186 5194
rect 4220 5058 4236 5194
rect 4170 5046 4236 5058
rect 4266 5194 4328 5206
rect 4266 5058 4282 5194
rect 4316 5058 4328 5194
rect 4266 5046 4328 5058
rect 3474 4994 3536 5006
<< ndiffc >>
rect 606 7794 726 7894
rect 766 7794 886 7894
rect 926 7794 1046 7894
rect 1086 7794 1206 7894
rect 1246 7794 1366 7894
rect 1406 7794 1526 7894
rect 1566 7794 1686 7894
rect 3186 7794 3306 7894
rect 3346 7794 3466 7894
rect 3506 7794 3626 7894
rect 3666 7794 3786 7894
rect 3826 7794 3946 7894
rect 3986 7794 4106 7894
rect 4146 7794 4266 7894
rect 606 6874 726 6974
rect 766 6874 886 6974
rect 926 6874 1046 6974
rect 1086 6874 1206 6974
rect 1246 6874 1366 6974
rect 1406 6874 1526 6974
rect 1566 6874 1686 6974
rect 3186 6874 3306 6974
rect 3346 6874 3466 6974
rect 3506 6874 3626 6974
rect 3666 6874 3786 6974
rect 3826 6874 3946 6974
rect 3986 6874 4106 6974
rect 4146 6874 4266 6974
rect 3202 5744 3236 5820
rect 3298 5744 3332 5820
rect 3394 5744 3428 5820
rect 3490 5744 3524 5820
rect 3738 5808 3772 5868
rect 3834 5808 3868 5868
rect 3930 5808 3964 5868
rect 4234 5808 4268 5868
rect 4330 5808 4364 5868
rect 4426 5808 4460 5868
rect 810 5276 844 5652
rect 906 5276 940 5652
rect 1002 5276 1036 5652
rect 1098 5276 1132 5652
rect 1194 5276 1228 5652
rect 1290 5276 1324 5652
rect 1386 5276 1420 5652
rect 1482 5276 1516 5652
rect 1578 5276 1612 5652
rect 362 5096 422 5130
rect 596 5096 656 5130
rect 362 5008 422 5042
rect 596 5008 656 5042
rect 810 5016 844 5092
rect 906 5016 940 5092
rect 1002 5016 1036 5092
rect 1098 5016 1132 5092
rect 1194 5016 1228 5092
rect 1290 5016 1324 5092
rect 1386 5016 1420 5092
rect 1482 5016 1516 5092
rect 1578 5016 1612 5092
rect 2264 5010 2298 5386
rect 2360 5010 2394 5386
rect 2456 5010 2490 5386
rect 2552 5010 2586 5386
rect 2648 5010 2682 5386
rect 3202 5432 3236 5508
rect 3298 5432 3332 5508
rect 3394 5432 3428 5508
rect 3490 5432 3524 5508
rect 3898 5388 3932 5448
rect 3994 5388 4028 5448
rect 4090 5388 4124 5448
rect 606 4204 726 4304
rect 766 4204 886 4304
rect 926 4204 1046 4304
rect 1086 4204 1206 4304
rect 1246 4204 1366 4304
rect 1406 4204 1526 4304
rect 1566 4204 1686 4304
rect 3186 4204 3306 4304
rect 3346 4204 3466 4304
rect 3506 4204 3626 4304
rect 3666 4204 3786 4304
rect 3826 4204 3946 4304
rect 3986 4204 4106 4304
rect 4146 4204 4266 4304
rect 606 3284 726 3384
rect 766 3284 886 3384
rect 926 3284 1046 3384
rect 1086 3284 1206 3384
rect 1246 3284 1366 3384
rect 1406 3284 1526 3384
rect 1566 3284 1686 3384
rect 3186 3284 3306 3384
rect 3346 3284 3466 3384
rect 3506 3284 3626 3384
rect 3666 3284 3786 3384
rect 3826 3284 3946 3384
rect 3986 3284 4106 3384
rect 4146 3284 4266 3384
<< pdiffc >>
rect 810 6090 844 6166
rect 906 6090 940 6166
rect 1002 6090 1036 6166
rect 1098 6090 1132 6166
rect 1194 6090 1228 6166
rect 1290 6090 1324 6166
rect 1386 6090 1420 6166
rect 1482 6090 1516 6166
rect 1578 6090 1612 6166
rect 1942 5740 1976 6116
rect 2038 5740 2072 6116
rect 2134 5740 2168 6116
rect 2264 5740 2298 6116
rect 2360 5740 2394 6116
rect 2456 5740 2490 6116
rect 2552 5740 2586 6116
rect 2648 5740 2682 6116
rect 2778 5740 2812 6116
rect 2874 5740 2908 6116
rect 2970 5740 3004 6116
rect 3202 6070 3236 6246
rect 3298 6070 3332 6246
rect 3394 6070 3428 6246
rect 3490 6070 3524 6246
rect 3738 6062 3772 6198
rect 3834 6062 3868 6198
rect 3930 6062 3964 6198
rect 4026 6062 4060 6198
rect 4122 6062 4156 6198
rect 4234 6062 4268 6198
rect 4330 6062 4364 6198
rect 4426 6062 4460 6198
rect 4522 6062 4556 6198
rect 4618 6062 4652 6198
rect 362 5440 422 5474
rect 596 5440 656 5474
rect 362 5348 422 5382
rect 596 5348 656 5382
rect 362 5258 422 5292
rect 596 5258 656 5292
rect 3202 5006 3236 5182
rect 3298 5006 3332 5182
rect 3394 5006 3428 5182
rect 3490 5006 3524 5182
rect 3898 5058 3932 5194
rect 3994 5058 4028 5194
rect 4090 5058 4124 5194
rect 4186 5058 4220 5194
rect 4282 5058 4316 5194
<< psubdiff >>
rect 430 8336 552 8362
rect 430 8262 454 8336
rect 528 8262 552 8336
rect 430 8238 552 8262
rect 978 8336 1100 8362
rect 978 8262 1002 8336
rect 1076 8262 1100 8336
rect 978 8238 1100 8262
rect 1526 8336 1648 8362
rect 1526 8262 1550 8336
rect 1624 8262 1648 8336
rect 1526 8238 1648 8262
rect 2074 8336 2196 8362
rect 2074 8262 2098 8336
rect 2172 8262 2196 8336
rect 2074 8238 2196 8262
rect 2622 8336 2744 8362
rect 2622 8262 2646 8336
rect 2720 8262 2744 8336
rect 2622 8238 2744 8262
rect 3152 8336 3274 8362
rect 3152 8262 3176 8336
rect 3250 8262 3274 8336
rect 3152 8238 3274 8262
rect 3700 8336 3822 8362
rect 3700 8262 3724 8336
rect 3798 8262 3822 8336
rect 3700 8238 3822 8262
rect 4250 8336 4372 8362
rect 4250 8262 4274 8336
rect 4348 8262 4372 8336
rect 4250 8238 4372 8262
rect 64 8194 186 8220
rect 64 8120 88 8194
rect 162 8120 186 8194
rect 64 8096 186 8120
rect 4746 8124 4868 8150
rect 916 8074 1376 8094
rect 916 8024 946 8074
rect 1346 8024 1376 8074
rect 916 8004 1376 8024
rect 3496 8074 3956 8094
rect 3496 8024 3526 8074
rect 3926 8024 3956 8074
rect 4746 8050 4770 8124
rect 4844 8050 4868 8124
rect 4746 8026 4868 8050
rect 3496 8004 3956 8024
rect 64 7720 186 7746
rect 64 7646 88 7720
rect 162 7646 186 7720
rect 64 7622 186 7646
rect 64 7246 186 7272
rect 64 7172 88 7246
rect 162 7172 186 7246
rect 64 7148 186 7172
rect 4746 7648 4868 7674
rect 4746 7574 4770 7648
rect 4844 7574 4868 7648
rect 4746 7550 4868 7574
rect 4746 7174 4868 7200
rect 4746 7100 4770 7174
rect 4844 7100 4868 7174
rect 4746 7076 4868 7100
rect 64 6772 186 6798
rect 64 6698 88 6772
rect 162 6698 186 6772
rect 64 6674 186 6698
rect 916 6744 1376 6764
rect 916 6694 946 6744
rect 1346 6694 1376 6744
rect 916 6674 1376 6694
rect 3496 6744 3956 6764
rect 3496 6694 3526 6744
rect 3926 6694 3956 6744
rect 3496 6674 3956 6694
rect 4744 6700 4866 6726
rect 4744 6626 4768 6700
rect 4842 6626 4866 6700
rect 4744 6608 4866 6626
rect 64 6086 186 6112
rect 64 6012 88 6086
rect 162 6012 186 6086
rect 64 5988 186 6012
rect 4744 6088 4866 6114
rect 4744 6014 4768 6088
rect 4842 6014 4866 6088
rect 4744 5990 4866 6014
rect 56 5560 178 5586
rect 56 5486 80 5560
rect 154 5486 178 5560
rect 56 5462 178 5486
rect 3810 5708 3834 5742
rect 3868 5708 3896 5742
rect 4306 5708 4330 5742
rect 4364 5708 4392 5742
rect 3190 5644 3216 5678
rect 3250 5644 3284 5678
rect 3318 5644 3352 5678
rect 3386 5644 3420 5678
rect 3454 5644 3488 5678
rect 3522 5644 3546 5678
rect 3190 5608 3546 5644
rect 3190 5574 3216 5608
rect 3250 5574 3284 5608
rect 3318 5574 3352 5608
rect 3386 5574 3420 5608
rect 3454 5574 3488 5608
rect 3522 5574 3546 5608
rect 4744 5614 4866 5640
rect 56 5086 178 5112
rect 56 5012 80 5086
rect 154 5012 178 5086
rect 56 4988 178 5012
rect 3970 5514 3994 5548
rect 4028 5514 4056 5548
rect 4744 5540 4768 5614
rect 4842 5540 4866 5614
rect 4744 5516 4866 5540
rect 350 4908 374 4942
rect 410 4908 434 4942
rect 350 4902 434 4908
rect 584 4908 608 4942
rect 644 4908 668 4942
rect 4744 5140 4866 5166
rect 4744 5066 4768 5140
rect 4842 5066 4866 5140
rect 4744 5042 4866 5066
rect 584 4902 668 4908
rect 2258 4850 2282 4886
rect 2318 4850 2374 4886
rect 2410 4850 2466 4886
rect 2502 4850 2558 4886
rect 2594 4850 2650 4886
rect 2686 4850 2710 4886
rect 2258 4848 2710 4850
rect 792 4842 1610 4844
rect 792 4806 816 4842
rect 852 4806 934 4842
rect 970 4806 1052 4842
rect 1088 4806 1170 4842
rect 1206 4806 1288 4842
rect 1324 4806 1406 4842
rect 1442 4806 1524 4842
rect 1560 4806 1610 4842
rect 792 4802 1610 4806
rect 916 4484 1376 4504
rect 70 4434 192 4460
rect 70 4360 94 4434
rect 168 4360 192 4434
rect 916 4434 946 4484
rect 1346 4434 1376 4484
rect 916 4414 1376 4434
rect 3496 4484 3956 4504
rect 3496 4434 3526 4484
rect 3926 4434 3956 4484
rect 3496 4414 3956 4434
rect 70 4336 192 4360
rect 4744 4404 4866 4430
rect 4744 4330 4768 4404
rect 4842 4330 4866 4404
rect 4744 4306 4866 4330
rect 70 3960 192 3986
rect 70 3886 94 3960
rect 168 3886 192 3960
rect 70 3862 192 3886
rect 70 3486 192 3512
rect 70 3412 94 3486
rect 168 3412 192 3486
rect 70 3388 192 3412
rect 4744 3930 4866 3956
rect 4744 3856 4768 3930
rect 4842 3856 4866 3930
rect 4744 3832 4866 3856
rect 4744 3456 4866 3482
rect 4744 3382 4768 3456
rect 4842 3382 4866 3456
rect 4744 3358 4866 3382
rect 916 3154 1376 3174
rect 916 3104 946 3154
rect 1346 3104 1376 3154
rect 916 3084 1376 3104
rect 3496 3154 3956 3174
rect 3496 3104 3526 3154
rect 3926 3104 3956 3154
rect 3496 3084 3956 3104
rect 600 2926 722 2952
rect 600 2852 624 2926
rect 698 2852 722 2926
rect 600 2828 722 2852
rect 1148 2926 1270 2952
rect 1148 2852 1172 2926
rect 1246 2852 1270 2926
rect 1148 2828 1270 2852
rect 1696 2926 1818 2952
rect 1696 2852 1720 2926
rect 1794 2852 1818 2926
rect 1696 2828 1818 2852
rect 2244 2926 2366 2952
rect 2244 2852 2268 2926
rect 2342 2852 2366 2926
rect 2244 2828 2366 2852
rect 2792 2926 2914 2952
rect 2792 2852 2816 2926
rect 2890 2852 2914 2926
rect 2792 2828 2914 2852
rect 3340 2926 3462 2952
rect 3340 2852 3364 2926
rect 3438 2852 3462 2926
rect 3340 2828 3462 2852
rect 3890 2926 4012 2952
rect 3890 2852 3914 2926
rect 3988 2852 4012 2926
rect 3890 2828 4012 2852
<< nsubdiff >>
rect 3190 6326 3214 6364
rect 3252 6326 3290 6364
rect 3328 6326 3366 6364
rect 3404 6326 3442 6364
rect 3480 6326 3536 6364
rect 3764 6334 3794 6368
rect 3828 6334 3862 6368
rect 3896 6334 3930 6368
rect 3964 6334 3998 6368
rect 4032 6334 4066 6368
rect 4100 6334 4142 6368
rect 4260 6334 4290 6368
rect 4324 6334 4358 6368
rect 4392 6334 4426 6368
rect 4460 6334 4494 6368
rect 4528 6334 4562 6368
rect 4596 6334 4638 6368
rect 2098 6284 2822 6292
rect 798 6274 1654 6282
rect 798 6240 828 6274
rect 862 6240 912 6274
rect 946 6240 996 6274
rect 1030 6240 1080 6274
rect 1114 6240 1164 6274
rect 1198 6240 1248 6274
rect 1282 6240 1332 6274
rect 1366 6240 1416 6274
rect 1450 6240 1500 6274
rect 1534 6240 1590 6274
rect 1624 6240 1654 6274
rect 2098 6250 2136 6284
rect 2170 6250 2220 6284
rect 2254 6250 2304 6284
rect 2338 6250 2388 6284
rect 2422 6250 2472 6284
rect 2506 6250 2556 6284
rect 2590 6250 2640 6284
rect 2674 6250 2724 6284
rect 2758 6250 2822 6284
rect 2098 6244 2822 6250
rect 798 6234 1654 6240
rect 350 5536 374 5572
rect 410 5536 434 5572
rect 584 5536 608 5572
rect 644 5536 668 5572
rect 3190 4888 3214 4926
rect 3252 4888 3290 4926
rect 3328 4888 3366 4926
rect 3404 4888 3442 4926
rect 3480 4888 3536 4926
rect 3924 4888 3954 4922
rect 3988 4888 4022 4922
rect 4056 4888 4090 4922
rect 4124 4888 4158 4922
rect 4192 4888 4226 4922
rect 4260 4888 4302 4922
<< psubdiffcont >>
rect 454 8262 528 8336
rect 1002 8262 1076 8336
rect 1550 8262 1624 8336
rect 2098 8262 2172 8336
rect 2646 8262 2720 8336
rect 3176 8262 3250 8336
rect 3724 8262 3798 8336
rect 4274 8262 4348 8336
rect 88 8120 162 8194
rect 946 8024 1346 8074
rect 3526 8024 3926 8074
rect 4770 8050 4844 8124
rect 88 7646 162 7720
rect 88 7172 162 7246
rect 4770 7574 4844 7648
rect 4770 7100 4844 7174
rect 88 6698 162 6772
rect 946 6694 1346 6744
rect 3526 6694 3926 6744
rect 4768 6626 4842 6700
rect 88 6012 162 6086
rect 4768 6014 4842 6088
rect 80 5486 154 5560
rect 3834 5708 3868 5742
rect 4330 5708 4364 5742
rect 3216 5644 3250 5678
rect 3284 5644 3318 5678
rect 3352 5644 3386 5678
rect 3420 5644 3454 5678
rect 3488 5644 3522 5678
rect 3216 5574 3250 5608
rect 3284 5574 3318 5608
rect 3352 5574 3386 5608
rect 3420 5574 3454 5608
rect 3488 5574 3522 5608
rect 80 5012 154 5086
rect 3994 5514 4028 5548
rect 4768 5540 4842 5614
rect 374 4908 410 4942
rect 608 4908 644 4942
rect 4768 5066 4842 5140
rect 2282 4850 2318 4886
rect 2374 4850 2410 4886
rect 2466 4850 2502 4886
rect 2558 4850 2594 4886
rect 2650 4850 2686 4886
rect 816 4806 852 4842
rect 934 4806 970 4842
rect 1052 4806 1088 4842
rect 1170 4806 1206 4842
rect 1288 4806 1324 4842
rect 1406 4806 1442 4842
rect 1524 4806 1560 4842
rect 94 4360 168 4434
rect 946 4434 1346 4484
rect 3526 4434 3926 4484
rect 4768 4330 4842 4404
rect 94 3886 168 3960
rect 94 3412 168 3486
rect 4768 3856 4842 3930
rect 4768 3382 4842 3456
rect 946 3104 1346 3154
rect 3526 3104 3926 3154
rect 624 2852 698 2926
rect 1172 2852 1246 2926
rect 1720 2852 1794 2926
rect 2268 2852 2342 2926
rect 2816 2852 2890 2926
rect 3364 2852 3438 2926
rect 3914 2852 3988 2926
<< nsubdiffcont >>
rect 3214 6326 3252 6364
rect 3290 6326 3328 6364
rect 3366 6326 3404 6364
rect 3442 6326 3480 6364
rect 3794 6334 3828 6368
rect 3862 6334 3896 6368
rect 3930 6334 3964 6368
rect 3998 6334 4032 6368
rect 4066 6334 4100 6368
rect 4290 6334 4324 6368
rect 4358 6334 4392 6368
rect 4426 6334 4460 6368
rect 4494 6334 4528 6368
rect 4562 6334 4596 6368
rect 828 6240 862 6274
rect 912 6240 946 6274
rect 996 6240 1030 6274
rect 1080 6240 1114 6274
rect 1164 6240 1198 6274
rect 1248 6240 1282 6274
rect 1332 6240 1366 6274
rect 1416 6240 1450 6274
rect 1500 6240 1534 6274
rect 1590 6240 1624 6274
rect 2136 6250 2170 6284
rect 2220 6250 2254 6284
rect 2304 6250 2338 6284
rect 2388 6250 2422 6284
rect 2472 6250 2506 6284
rect 2556 6250 2590 6284
rect 2640 6250 2674 6284
rect 2724 6250 2758 6284
rect 374 5536 410 5572
rect 608 5536 644 5572
rect 3214 4888 3252 4926
rect 3290 4888 3328 4926
rect 3366 4888 3404 4926
rect 3442 4888 3480 4926
rect 3954 4888 3988 4922
rect 4022 4888 4056 4922
rect 4090 4888 4124 4922
rect 4158 4888 4192 4922
rect 4226 4888 4260 4922
<< poly >>
rect 476 7644 596 7774
rect 476 7594 506 7644
rect 556 7594 596 7644
rect 476 7554 596 7594
rect 476 7504 506 7554
rect 556 7504 596 7554
rect 476 7464 596 7504
rect 476 7414 506 7464
rect 556 7414 596 7464
rect 476 7364 596 7414
rect 476 7314 506 7364
rect 556 7314 596 7364
rect 476 7274 596 7314
rect 476 7224 506 7274
rect 556 7224 596 7274
rect 476 7184 596 7224
rect 476 7134 506 7184
rect 556 7134 596 7184
rect 476 6994 596 7134
rect 4276 7634 4386 7774
rect 4276 7584 4316 7634
rect 4366 7584 4386 7634
rect 4276 7544 4386 7584
rect 4276 7494 4316 7544
rect 4366 7494 4386 7544
rect 4276 7454 4386 7494
rect 4276 7404 4316 7454
rect 4366 7424 4386 7454
rect 4366 7404 4396 7424
rect 4276 7354 4396 7404
rect 4276 7304 4316 7354
rect 4366 7344 4396 7354
rect 4366 7304 4386 7344
rect 4276 7264 4386 7304
rect 4276 7214 4316 7264
rect 4366 7214 4386 7264
rect 4276 7174 4386 7214
rect 4276 7124 4316 7174
rect 4366 7124 4386 7174
rect 4276 6994 4386 7124
rect 3348 6284 3474 6314
rect 3252 6258 3282 6284
rect 3348 6258 3378 6284
rect 3444 6258 3474 6284
rect 3744 6292 4010 6308
rect 3744 6258 3754 6292
rect 3788 6278 4010 6292
rect 3788 6258 3818 6278
rect 860 6178 890 6204
rect 956 6178 986 6204
rect 1052 6178 1082 6204
rect 1148 6178 1178 6204
rect 1244 6178 1274 6204
rect 1340 6178 1370 6204
rect 1436 6178 1466 6204
rect 1532 6178 1562 6204
rect 1992 6128 2022 6154
rect 2088 6128 2118 6154
rect 2314 6128 2344 6154
rect 2410 6128 2440 6154
rect 2506 6128 2536 6154
rect 2602 6128 2632 6154
rect 2828 6128 2858 6154
rect 2924 6128 2954 6154
rect 860 6052 890 6078
rect 956 6052 986 6078
rect 1052 6052 1082 6078
rect 1148 6052 1178 6078
rect 1244 6052 1274 6078
rect 1340 6052 1370 6078
rect 1436 6052 1466 6078
rect 1532 6052 1562 6078
rect 860 6020 1562 6052
rect 1182 5978 1240 6020
rect 702 5968 1240 5978
rect 702 5934 718 5968
rect 752 5942 1240 5968
rect 752 5934 768 5942
rect 702 5920 768 5934
rect 1368 5890 1440 5900
rect 1368 5850 1384 5890
rect 1424 5850 1440 5890
rect 976 5840 1048 5850
rect 1368 5840 1440 5850
rect 1816 5880 1884 5890
rect 1816 5844 1832 5880
rect 1868 5844 1884 5880
rect 976 5800 992 5840
rect 1032 5800 1048 5840
rect 976 5790 1048 5800
rect 1000 5720 1038 5790
rect 1384 5720 1422 5840
rect 1816 5806 1884 5844
rect 1816 5770 1832 5806
rect 1868 5770 1884 5806
rect 1816 5732 1884 5770
rect 860 5690 1178 5720
rect 860 5664 890 5690
rect 956 5664 986 5690
rect 1052 5664 1082 5690
rect 1148 5664 1178 5690
rect 1244 5690 1562 5720
rect 1244 5664 1274 5690
rect 1340 5664 1370 5690
rect 1436 5664 1466 5690
rect 1532 5664 1562 5690
rect 1816 5696 1832 5732
rect 1868 5712 1884 5732
rect 3744 6242 3818 6258
rect 3788 6210 3818 6242
rect 3884 6210 3914 6236
rect 3980 6210 4010 6278
rect 4240 6292 4506 6308
rect 4240 6258 4250 6292
rect 4284 6278 4506 6292
rect 4284 6258 4314 6278
rect 4240 6242 4314 6258
rect 4076 6210 4106 6236
rect 4284 6210 4314 6242
rect 4380 6210 4410 6236
rect 4476 6210 4506 6278
rect 4572 6210 4602 6236
rect 3252 6032 3282 6058
rect 3240 6008 3282 6032
rect 3112 5970 3186 5986
rect 3112 5936 3126 5970
rect 3162 5936 3186 5970
rect 3112 5918 3186 5936
rect 3240 5918 3272 6008
rect 3348 5976 3378 6058
rect 3444 6032 3474 6058
rect 3112 5898 3272 5918
rect 3314 5959 3378 5976
rect 3314 5925 3324 5959
rect 3358 5925 3378 5959
rect 3788 5936 3818 6050
rect 3884 6018 3914 6050
rect 3980 6024 4010 6050
rect 3860 6002 3914 6018
rect 3860 5968 3870 6002
rect 3904 5982 3914 6002
rect 4076 5982 4106 6050
rect 3904 5968 4106 5982
rect 3860 5952 4106 5968
rect 3314 5908 3378 5925
rect 3112 5864 3126 5898
rect 3162 5882 3272 5898
rect 3162 5864 3186 5882
rect 3112 5848 3186 5864
rect 3240 5880 3272 5882
rect 3240 5856 3282 5880
rect 3252 5832 3282 5856
rect 3348 5878 3378 5908
rect 3680 5904 3818 5936
rect 3348 5848 3474 5878
rect 3348 5832 3378 5848
rect 3444 5832 3474 5848
rect 3680 5744 3710 5904
rect 3788 5880 3818 5904
rect 3884 5880 3914 5952
rect 4284 5880 4314 6050
rect 4380 6018 4410 6050
rect 4476 6024 4506 6050
rect 4356 6002 4410 6018
rect 4356 5968 4366 6002
rect 4400 5982 4410 6002
rect 4572 5982 4602 6050
rect 4400 5968 4602 5982
rect 4356 5952 4602 5968
rect 4380 5880 4410 5952
rect 3788 5770 3818 5796
rect 3884 5770 3914 5796
rect 4284 5770 4314 5796
rect 4380 5770 4410 5796
rect 1992 5712 2022 5728
rect 2088 5712 2118 5728
rect 1868 5696 2118 5712
rect 1816 5682 2118 5696
rect 2314 5712 2344 5728
rect 2410 5712 2440 5728
rect 2314 5682 2440 5712
rect 304 5396 350 5426
rect 438 5396 464 5426
rect 538 5396 584 5426
rect 672 5396 698 5426
rect 304 5334 334 5396
rect 538 5334 568 5396
rect 304 5304 350 5334
rect 438 5304 464 5334
rect 538 5304 584 5334
rect 672 5304 698 5334
rect 304 5220 334 5304
rect 538 5220 568 5304
rect 2406 5616 2440 5682
rect 2374 5606 2440 5616
rect 2374 5572 2390 5606
rect 2424 5572 2440 5606
rect 2374 5562 2440 5572
rect 2314 5398 2344 5424
rect 2410 5398 2440 5562
rect 2506 5712 2536 5728
rect 2602 5712 2632 5728
rect 2506 5682 2632 5712
rect 2828 5712 2858 5728
rect 2924 5712 2954 5728
rect 2828 5682 2954 5712
rect 3252 5706 3282 5732
rect 3348 5706 3378 5732
rect 3444 5706 3474 5732
rect 3680 5726 3754 5744
rect 2506 5548 2540 5682
rect 2506 5538 2766 5548
rect 2506 5504 2524 5538
rect 2558 5504 2766 5538
rect 2920 5506 2954 5682
rect 3680 5692 3710 5726
rect 3744 5692 3754 5726
rect 3680 5676 3754 5692
rect 3252 5520 3282 5546
rect 3348 5520 3378 5546
rect 3444 5520 3474 5546
rect 2506 5494 2766 5504
rect 2506 5398 2536 5494
rect 2602 5398 2632 5424
rect 860 5236 890 5264
rect 956 5236 986 5264
rect 1052 5236 1082 5264
rect 1148 5236 1178 5264
rect 1244 5236 1274 5264
rect 1340 5236 1370 5264
rect 1436 5236 1466 5264
rect 1532 5236 1562 5264
rect 262 5204 334 5220
rect 262 5170 278 5204
rect 312 5170 334 5204
rect 262 5154 334 5170
rect 496 5204 568 5220
rect 496 5170 512 5204
rect 546 5170 568 5204
rect 496 5154 568 5170
rect 304 5084 334 5154
rect 538 5084 568 5154
rect 710 5170 776 5180
rect 710 5136 726 5170
rect 760 5160 776 5170
rect 760 5136 1562 5160
rect 710 5130 1562 5136
rect 710 5126 776 5130
rect 860 5104 890 5130
rect 956 5104 986 5130
rect 1052 5104 1082 5130
rect 1148 5104 1178 5130
rect 1244 5104 1274 5130
rect 1340 5104 1370 5130
rect 1436 5104 1466 5130
rect 1532 5104 1562 5130
rect 304 5054 350 5084
rect 434 5054 460 5084
rect 538 5054 584 5084
rect 668 5054 694 5084
rect 860 4978 890 5004
rect 956 4978 986 5004
rect 1052 4978 1082 5004
rect 1148 4978 1178 5004
rect 1244 4978 1274 5004
rect 1340 4978 1370 5004
rect 1436 4978 1466 5004
rect 1532 4978 1562 5004
rect 2710 5378 2766 5494
rect 2824 5490 2954 5506
rect 2824 5454 2834 5490
rect 2870 5454 2908 5490
rect 2944 5454 2954 5490
rect 2824 5438 2954 5454
rect 3948 5460 3978 5486
rect 4044 5460 4074 5486
rect 3252 5396 3282 5420
rect 2710 5370 3186 5378
rect 3240 5372 3282 5396
rect 3348 5404 3378 5420
rect 3444 5404 3474 5420
rect 3348 5374 3474 5404
rect 3240 5370 3272 5372
rect 2710 5334 3272 5370
rect 3348 5344 3378 5374
rect 2710 5322 3186 5334
rect 3240 5244 3272 5334
rect 3314 5327 3378 5344
rect 3314 5293 3324 5327
rect 3358 5293 3378 5327
rect 3314 5276 3378 5293
rect 3240 5220 3282 5244
rect 3252 5194 3282 5220
rect 3348 5194 3378 5276
rect 3444 5194 3474 5220
rect 3948 5206 3978 5376
rect 4044 5304 4074 5376
rect 4020 5288 4266 5304
rect 4020 5254 4030 5288
rect 4064 5274 4266 5288
rect 4064 5254 4074 5274
rect 4020 5238 4074 5254
rect 4044 5206 4074 5238
rect 4140 5206 4170 5232
rect 4236 5206 4266 5274
rect 2314 4930 2344 4998
rect 2410 4972 2440 4998
rect 2506 4972 2536 4998
rect 2602 4930 2632 4998
rect 3948 5014 3978 5046
rect 4044 5020 4074 5046
rect 3904 4998 3978 5014
rect 3252 4968 3282 4994
rect 3348 4968 3378 4994
rect 3444 4968 3474 4994
rect 3348 4938 3474 4968
rect 3904 4964 3914 4998
rect 3948 4978 3978 4998
rect 4140 4978 4170 5046
rect 4236 5020 4266 5046
rect 3948 4964 4170 4978
rect 3904 4948 4170 4964
rect 2078 4920 2632 4930
rect 2078 4886 2094 4920
rect 2128 4886 2172 4920
rect 2206 4900 2632 4920
rect 2206 4886 2222 4900
rect 2078 4876 2222 4886
rect 476 4054 596 4184
rect 476 4004 506 4054
rect 556 4004 596 4054
rect 476 3964 596 4004
rect 476 3914 506 3964
rect 556 3914 596 3964
rect 476 3874 596 3914
rect 476 3824 506 3874
rect 556 3824 596 3874
rect 476 3774 596 3824
rect 476 3724 506 3774
rect 556 3724 596 3774
rect 476 3684 596 3724
rect 476 3634 506 3684
rect 556 3634 596 3684
rect 476 3594 596 3634
rect 476 3544 506 3594
rect 556 3544 596 3594
rect 476 3404 596 3544
rect 4276 4044 4386 4184
rect 4276 3994 4316 4044
rect 4366 3994 4386 4044
rect 4276 3954 4386 3994
rect 4276 3904 4316 3954
rect 4366 3904 4386 3954
rect 4276 3864 4386 3904
rect 4276 3814 4316 3864
rect 4366 3834 4386 3864
rect 4366 3814 4396 3834
rect 4276 3764 4396 3814
rect 4276 3714 4316 3764
rect 4366 3754 4396 3764
rect 4366 3714 4386 3754
rect 4276 3674 4386 3714
rect 4276 3624 4316 3674
rect 4366 3624 4386 3674
rect 4276 3584 4386 3624
rect 4276 3534 4316 3584
rect 4366 3534 4386 3584
rect 4276 3404 4386 3534
<< polycont >>
rect 506 7594 556 7644
rect 506 7504 556 7554
rect 506 7414 556 7464
rect 506 7314 556 7364
rect 506 7224 556 7274
rect 506 7134 556 7184
rect 4316 7584 4366 7634
rect 4316 7494 4366 7544
rect 4316 7404 4366 7454
rect 4316 7304 4366 7354
rect 4316 7214 4366 7264
rect 4316 7124 4366 7174
rect 3754 6258 3788 6292
rect 718 5934 752 5968
rect 1384 5850 1424 5890
rect 1832 5844 1868 5880
rect 992 5800 1032 5840
rect 1832 5770 1868 5806
rect 1832 5696 1868 5732
rect 4250 6258 4284 6292
rect 3126 5936 3162 5970
rect 3324 5925 3358 5959
rect 3870 5968 3904 6002
rect 3126 5864 3162 5898
rect 4366 5968 4400 6002
rect 2390 5572 2424 5606
rect 2524 5504 2558 5538
rect 3710 5692 3744 5726
rect 278 5170 312 5204
rect 512 5170 546 5204
rect 726 5136 760 5170
rect 2834 5454 2870 5490
rect 2908 5454 2944 5490
rect 3324 5293 3358 5327
rect 4030 5254 4064 5288
rect 3914 4964 3948 4998
rect 2094 4886 2128 4920
rect 2172 4886 2206 4920
rect 506 4004 556 4054
rect 506 3914 556 3964
rect 506 3824 556 3874
rect 506 3724 556 3774
rect 506 3634 556 3684
rect 506 3544 556 3594
rect 4316 3994 4366 4044
rect 4316 3904 4366 3954
rect 4316 3814 4366 3864
rect 4316 3714 4366 3764
rect 4316 3624 4366 3674
rect 4316 3534 4366 3584
<< locali >>
rect 30 8336 4908 8392
rect 30 8262 454 8336
rect 528 8262 1002 8336
rect 1076 8262 1550 8336
rect 1624 8262 2098 8336
rect 2172 8262 2646 8336
rect 2720 8262 3176 8336
rect 3250 8262 3724 8336
rect 3798 8262 4274 8336
rect 4348 8262 4908 8336
rect 30 8194 4908 8262
rect 30 8144 88 8194
rect 162 8144 266 8194
rect 30 7744 66 8144
rect 196 7744 266 8144
rect 916 8094 1376 8194
rect 3496 8094 3956 8194
rect 4710 8124 4908 8194
rect 30 7720 266 7744
rect 30 7646 88 7720
rect 162 7704 266 7720
rect 346 8074 4526 8094
rect 346 8024 946 8074
rect 1346 8024 3526 8074
rect 3926 8024 4526 8074
rect 346 8014 4526 8024
rect 162 7646 228 7704
rect 30 7604 228 7646
rect 30 7164 50 7604
rect 186 7164 228 7604
rect 30 7044 228 7164
rect 30 6614 50 7044
rect 206 6614 228 7044
rect 346 6754 426 8014
rect 916 8004 1376 8014
rect 3496 8004 3956 8014
rect 586 7794 606 7894
rect 726 7794 766 7894
rect 886 7794 926 7894
rect 1046 7794 1086 7894
rect 1206 7794 1246 7894
rect 1366 7794 1406 7894
rect 1526 7794 1566 7894
rect 1686 7794 3186 7894
rect 3306 7794 3346 7894
rect 3466 7794 3506 7894
rect 3626 7794 3666 7894
rect 3786 7794 3826 7894
rect 3946 7794 3986 7894
rect 4106 7794 4146 7894
rect 4266 7794 4286 7894
rect 586 7774 4286 7794
rect 506 7694 1066 7734
rect 506 7644 616 7694
rect 1106 7654 1176 7774
rect 556 7594 616 7644
rect 656 7614 1176 7654
rect 506 7574 616 7594
rect 506 7554 1066 7574
rect 576 7534 1066 7554
rect 576 7504 616 7534
rect 506 7464 616 7504
rect 1106 7494 1176 7614
rect 576 7414 616 7464
rect 656 7454 1176 7494
rect 1216 7424 1256 7734
rect 1296 7474 1336 7774
rect 1376 7424 1416 7734
rect 1456 7474 1496 7774
rect 1536 7424 1576 7734
rect 1616 7474 1656 7774
rect 1696 7424 1736 7734
rect 1776 7474 1816 7774
rect 1856 7424 1896 7734
rect 1936 7474 1976 7774
rect 2016 7424 2056 7734
rect 2096 7474 2136 7774
rect 2176 7424 2216 7734
rect 2256 7474 2296 7774
rect 2336 7424 2376 7734
rect 2416 7474 2456 7774
rect 2496 7424 2536 7734
rect 2576 7474 2616 7774
rect 2656 7424 2696 7734
rect 2736 7474 2776 7774
rect 2816 7424 2856 7734
rect 2896 7474 2936 7774
rect 2976 7424 3016 7734
rect 3056 7474 3096 7774
rect 3136 7424 3176 7734
rect 3216 7474 3256 7774
rect 3296 7424 3336 7734
rect 3376 7474 3416 7774
rect 3456 7424 3496 7734
rect 3536 7474 3576 7774
rect 3616 7424 3656 7734
rect 3696 7654 3766 7774
rect 3806 7694 4366 7734
rect 3696 7614 4216 7654
rect 4256 7634 4366 7694
rect 3696 7494 3766 7614
rect 4256 7584 4316 7634
rect 4256 7574 4366 7584
rect 3806 7544 4366 7574
rect 3806 7534 4296 7544
rect 4256 7494 4296 7534
rect 3696 7454 4206 7494
rect 4256 7454 4366 7494
rect 1216 7414 3656 7424
rect 4256 7414 4296 7454
rect 506 7404 4296 7414
rect 506 7364 4366 7404
rect 576 7354 4366 7364
rect 576 7314 616 7354
rect 1216 7344 3656 7354
rect 506 7274 616 7314
rect 656 7274 1176 7314
rect 576 7234 616 7274
rect 576 7224 1066 7234
rect 506 7194 1066 7224
rect 506 7184 616 7194
rect 556 7134 616 7184
rect 1106 7154 1176 7274
rect 506 7074 616 7134
rect 656 7114 1176 7154
rect 506 7034 1066 7074
rect 1106 6994 1176 7114
rect 1216 7034 1256 7344
rect 1296 6994 1336 7294
rect 1376 7034 1416 7344
rect 1456 6994 1496 7294
rect 1536 7034 1576 7344
rect 1616 6994 1656 7294
rect 1696 7034 1736 7344
rect 1776 6994 1816 7294
rect 1856 7034 1896 7344
rect 1936 6994 1976 7294
rect 2016 7034 2056 7344
rect 2096 6994 2136 7294
rect 2176 7034 2216 7344
rect 2256 6994 2296 7294
rect 2336 7044 2376 7344
rect 2416 6994 2456 7294
rect 2496 7044 2536 7344
rect 2576 6994 2616 7294
rect 2656 7034 2696 7344
rect 2736 6994 2776 7294
rect 2816 7034 2856 7344
rect 2896 6994 2936 7294
rect 2976 7034 3016 7344
rect 3056 6994 3096 7294
rect 3136 7034 3176 7344
rect 3216 6994 3256 7294
rect 3296 7034 3336 7344
rect 3376 6994 3416 7294
rect 3456 7034 3496 7344
rect 3536 6994 3576 7294
rect 3616 7034 3656 7344
rect 3696 7274 4206 7314
rect 4256 7304 4296 7354
rect 3696 7154 3766 7274
rect 4256 7264 4366 7304
rect 4256 7234 4296 7264
rect 3806 7214 4296 7234
rect 3806 7194 4366 7214
rect 4256 7174 4366 7194
rect 3696 7114 4216 7154
rect 4256 7124 4316 7174
rect 3696 6994 3766 7114
rect 4256 7074 4366 7124
rect 3806 7034 4366 7074
rect 586 6974 4286 6994
rect 586 6874 606 6974
rect 726 6874 766 6974
rect 886 6874 926 6974
rect 1046 6874 1086 6974
rect 1206 6874 1246 6974
rect 1366 6874 1406 6974
rect 1526 6874 1566 6974
rect 1686 6874 3186 6974
rect 3306 6874 3346 6974
rect 3466 6874 3506 6974
rect 3626 6874 3666 6974
rect 3786 6874 3826 6974
rect 3946 6874 3986 6974
rect 4106 6874 4146 6974
rect 4266 6874 4286 6974
rect 916 6754 1376 6764
rect 3496 6754 3956 6764
rect 4446 6754 4526 8014
rect 346 6744 4526 6754
rect 346 6694 946 6744
rect 1346 6694 3526 6744
rect 3926 6694 4526 6744
rect 346 6674 4526 6694
rect 4710 8050 4770 8124
rect 4844 8050 4908 8124
rect 4710 7648 4908 8050
rect 4710 7574 4770 7648
rect 4844 7574 4908 7648
rect 4710 7174 4908 7574
rect 4710 7100 4770 7174
rect 4844 7100 4908 7174
rect 4710 6700 4908 7100
rect 30 6086 228 6614
rect 916 6594 1376 6674
rect 3496 6594 3956 6674
rect 4710 6626 4768 6700
rect 4842 6626 4908 6700
rect 3120 6404 3668 6424
rect 3120 6368 3214 6404
rect 3250 6368 3290 6404
rect 3326 6368 3366 6404
rect 3402 6368 3442 6404
rect 3478 6368 3518 6404
rect 3554 6368 3594 6404
rect 3630 6368 3668 6404
rect 3120 6364 3668 6368
rect 3120 6326 3214 6364
rect 3252 6326 3290 6364
rect 3328 6326 3366 6364
rect 3404 6326 3442 6364
rect 3480 6326 3668 6364
rect 3778 6334 3794 6368
rect 3828 6334 3862 6368
rect 3896 6334 3930 6368
rect 3964 6334 3998 6368
rect 4032 6334 4066 6368
rect 4100 6334 4290 6368
rect 4324 6334 4358 6368
rect 4392 6334 4426 6368
rect 4460 6334 4494 6368
rect 4528 6334 4562 6368
rect 4596 6334 4624 6368
rect 2098 6284 2822 6292
rect 30 6012 88 6086
rect 162 6012 228 6086
rect 30 5560 228 6012
rect 582 6276 1654 6282
rect 582 6240 594 6276
rect 628 6240 672 6276
rect 706 6240 744 6276
rect 778 6274 1654 6276
rect 778 6240 828 6274
rect 862 6240 912 6274
rect 946 6240 996 6274
rect 1030 6240 1080 6274
rect 1114 6240 1164 6274
rect 1198 6240 1248 6274
rect 1282 6240 1332 6274
rect 1366 6240 1416 6274
rect 1450 6240 1500 6274
rect 1534 6240 1590 6274
rect 1624 6240 1654 6274
rect 2098 6250 2136 6284
rect 2170 6250 2220 6284
rect 2254 6250 2304 6284
rect 2338 6250 2388 6284
rect 2422 6250 2472 6284
rect 2506 6250 2556 6284
rect 2590 6250 2640 6284
rect 2674 6250 2724 6284
rect 2758 6250 2822 6284
rect 2098 6244 2822 6250
rect 3202 6246 3236 6262
rect 582 6234 1654 6240
rect 582 5608 668 6234
rect 810 6216 1612 6234
rect 810 6166 844 6216
rect 810 6074 844 6090
rect 906 6166 940 6182
rect 906 6014 940 6090
rect 1002 6166 1036 6216
rect 1002 6074 1036 6090
rect 1098 6166 1132 6182
rect 1098 6014 1132 6090
rect 1194 6166 1228 6216
rect 1194 6074 1228 6090
rect 1290 6166 1324 6182
rect 906 5980 1132 6014
rect 1290 6014 1324 6090
rect 1386 6166 1420 6216
rect 1386 6074 1420 6090
rect 1482 6166 1516 6182
rect 1482 6014 1516 6090
rect 1578 6166 1612 6216
rect 1578 6074 1612 6090
rect 1706 6224 1896 6244
rect 1706 6074 1726 6224
rect 1876 6074 1896 6224
rect 2434 6210 2524 6244
rect 1706 6054 1896 6074
rect 1942 6166 2168 6200
rect 1942 6116 1976 6166
rect 1290 5980 1516 6014
rect 702 5968 768 5978
rect 702 5934 718 5968
rect 752 5934 768 5968
rect 702 5920 768 5934
rect 30 5486 80 5560
rect 154 5486 228 5560
rect 30 5086 228 5486
rect 262 5574 374 5608
rect 410 5574 608 5608
rect 644 5574 668 5608
rect 262 5572 668 5574
rect 262 5568 374 5572
rect 262 5384 298 5568
rect 350 5536 374 5568
rect 410 5568 608 5572
rect 410 5536 434 5568
rect 350 5476 438 5482
rect 346 5474 442 5476
rect 346 5440 362 5474
rect 422 5440 442 5474
rect 346 5438 442 5440
rect 488 5384 532 5568
rect 584 5536 608 5568
rect 644 5536 668 5572
rect 584 5476 672 5482
rect 580 5474 676 5476
rect 580 5440 596 5474
rect 656 5440 676 5474
rect 580 5438 676 5440
rect 262 5382 442 5384
rect 262 5348 362 5382
rect 422 5348 442 5382
rect 262 5346 442 5348
rect 488 5382 676 5384
rect 488 5348 596 5382
rect 656 5348 676 5382
rect 488 5346 676 5348
rect 346 5258 362 5292
rect 422 5258 442 5292
rect 580 5258 596 5292
rect 656 5258 676 5292
rect 350 5246 438 5258
rect 584 5246 672 5258
rect 262 5204 316 5220
rect 262 5170 278 5204
rect 312 5170 316 5204
rect 262 5154 316 5170
rect 350 5210 434 5246
rect 496 5210 550 5220
rect 350 5204 550 5210
rect 350 5170 512 5204
rect 546 5170 550 5204
rect 350 5164 550 5170
rect 350 5130 434 5164
rect 496 5154 550 5164
rect 584 5210 668 5246
rect 722 5210 768 5920
rect 906 5756 940 5980
rect 976 5840 1048 5850
rect 976 5800 992 5840
rect 1032 5800 1048 5840
rect 976 5790 1048 5800
rect 1084 5810 1132 5816
rect 1084 5774 1090 5810
rect 1126 5774 1132 5810
rect 1084 5756 1132 5774
rect 906 5722 1132 5756
rect 584 5180 768 5210
rect 810 5652 844 5668
rect 810 5226 844 5276
rect 906 5652 940 5722
rect 906 5260 940 5276
rect 1002 5652 1036 5668
rect 1002 5226 1036 5276
rect 1098 5652 1132 5722
rect 1290 5758 1324 5980
rect 1368 5890 1440 5900
rect 1368 5850 1384 5890
rect 1424 5850 1440 5890
rect 1368 5840 1440 5850
rect 1812 5880 1888 6054
rect 1812 5844 1832 5880
rect 1868 5844 1888 5880
rect 1812 5806 1888 5844
rect 1812 5770 1832 5806
rect 1868 5770 1888 5806
rect 1290 5724 1766 5758
rect 1098 5260 1132 5276
rect 1194 5652 1228 5668
rect 1194 5226 1228 5276
rect 1290 5652 1324 5724
rect 1290 5260 1324 5276
rect 1386 5652 1420 5668
rect 1386 5226 1420 5276
rect 1482 5652 1516 5724
rect 1482 5260 1516 5276
rect 1578 5652 1612 5668
rect 1690 5634 1766 5724
rect 1812 5732 1888 5770
rect 1812 5696 1832 5732
rect 1868 5696 1888 5732
rect 1812 5668 1888 5696
rect 1690 5622 1888 5634
rect 1690 5586 1832 5622
rect 1868 5586 1888 5622
rect 1942 5606 1976 5740
rect 2038 6116 2072 6132
rect 2038 5674 2072 5740
rect 2134 6116 2168 6166
rect 2134 5724 2168 5740
rect 2264 6176 2682 6210
rect 2264 6116 2298 6176
rect 2264 5724 2298 5740
rect 2360 6116 2394 6132
rect 2360 5674 2394 5740
rect 2456 6116 2490 6176
rect 2456 5724 2490 5740
rect 2552 6116 2586 6132
rect 2038 5640 2394 5674
rect 2552 5674 2586 5740
rect 2648 6116 2682 6176
rect 2648 5724 2682 5740
rect 2778 6166 3004 6200
rect 2778 6116 2812 6166
rect 2778 5724 2812 5740
rect 2874 6116 2908 6132
rect 2874 5674 2908 5740
rect 2552 5640 2908 5674
rect 2970 6116 3004 6166
rect 3004 5970 3168 5986
rect 3004 5936 3126 5970
rect 3162 5936 3168 5970
rect 3004 5898 3168 5936
rect 3004 5864 3126 5898
rect 3162 5864 3168 5898
rect 3004 5848 3168 5864
rect 3202 5976 3236 6070
rect 3298 6246 3332 6326
rect 3298 6054 3332 6070
rect 3394 6246 3428 6262
rect 3202 5959 3360 5976
rect 3202 5925 3324 5959
rect 3358 5925 3360 5959
rect 3202 5908 3360 5925
rect 3394 5940 3428 6070
rect 3490 6246 3524 6326
rect 3490 6054 3524 6070
rect 3502 5940 3562 5950
rect 3394 5938 3576 5940
rect 2970 5606 3004 5740
rect 3202 5820 3236 5908
rect 3394 5902 3508 5938
rect 3544 5902 3576 5938
rect 3202 5728 3236 5744
rect 3298 5820 3332 5836
rect 3298 5678 3332 5744
rect 3394 5820 3428 5902
rect 3502 5890 3562 5902
rect 3394 5728 3428 5744
rect 3490 5820 3524 5836
rect 3490 5678 3524 5744
rect 3190 5660 3216 5678
rect 3054 5644 3216 5660
rect 3250 5644 3284 5678
rect 3318 5644 3352 5678
rect 3386 5644 3420 5678
rect 3454 5644 3488 5678
rect 3522 5644 3546 5678
rect 3054 5608 3546 5644
rect 1690 5546 1888 5586
rect 1926 5572 2338 5606
rect 2374 5572 2390 5606
rect 2424 5572 3016 5606
rect 3054 5592 3216 5608
rect 1690 5510 1832 5546
rect 1868 5510 1888 5546
rect 1690 5472 1888 5510
rect 2304 5538 2338 5572
rect 2304 5504 2524 5538
rect 2558 5504 2574 5538
rect 1690 5436 1832 5472
rect 1868 5436 1888 5472
rect 1690 5422 1888 5436
rect 1578 5226 1612 5276
rect 810 5190 1612 5226
rect 584 5170 776 5180
rect 584 5164 726 5170
rect 584 5130 668 5164
rect 710 5136 726 5164
rect 760 5136 776 5170
rect 346 5096 362 5130
rect 422 5096 438 5130
rect 580 5096 596 5130
rect 656 5096 672 5130
rect 710 5126 776 5136
rect 350 5090 434 5096
rect 584 5090 668 5096
rect 810 5092 844 5190
rect 30 5012 80 5086
rect 154 5012 228 5086
rect 30 4952 228 5012
rect 346 5008 362 5042
rect 422 5008 438 5042
rect 580 5008 596 5042
rect 656 5008 672 5042
rect 30 4918 46 4952
rect 80 4918 118 4952
rect 152 4918 190 4952
rect 224 4918 228 4952
rect 30 4880 228 4918
rect 350 4942 434 5008
rect 350 4908 374 4942
rect 410 4908 434 4942
rect 350 4902 434 4908
rect 584 4942 668 5008
rect 810 5000 844 5016
rect 906 5092 940 5110
rect 584 4908 608 4942
rect 644 4908 668 4942
rect 584 4902 668 4908
rect 30 4846 46 4880
rect 80 4846 118 4880
rect 152 4846 190 4880
rect 224 4846 228 4880
rect 30 4808 228 4846
rect 906 4858 940 5016
rect 1002 5092 1036 5190
rect 1002 5000 1036 5016
rect 1098 5092 1132 5108
rect 1098 4858 1132 5016
rect 1194 5092 1228 5190
rect 1194 5000 1228 5016
rect 1290 5092 1324 5108
rect 1290 4858 1324 5016
rect 1386 5092 1420 5190
rect 1386 5000 1420 5016
rect 1482 5092 1516 5108
rect 1482 4858 1516 5016
rect 1578 5092 1612 5190
rect 1812 5164 1888 5422
rect 2264 5386 2298 5402
rect 1578 5000 1612 5016
rect 1806 5144 1996 5164
rect 1806 4994 1826 5144
rect 1976 4994 1996 5144
rect 1806 4974 1996 4994
rect 2078 4920 2222 4930
rect 2078 4886 2094 4920
rect 2128 4886 2172 4920
rect 2206 4886 2222 4920
rect 2264 4886 2298 5010
rect 2360 5386 2394 5504
rect 2618 5470 2652 5572
rect 2552 5436 2652 5470
rect 2828 5490 2950 5506
rect 2828 5454 2834 5490
rect 2870 5454 2908 5490
rect 2944 5454 2950 5490
rect 2828 5438 2950 5454
rect 2360 4994 2394 5010
rect 2456 5386 2490 5402
rect 2456 4886 2490 5010
rect 2552 5386 2586 5436
rect 2552 4994 2586 5010
rect 2648 5386 2682 5402
rect 3054 5266 3122 5592
rect 3190 5574 3216 5592
rect 3250 5574 3284 5608
rect 3318 5574 3352 5608
rect 3386 5574 3420 5608
rect 3454 5574 3488 5608
rect 3522 5574 3546 5608
rect 2648 4886 2682 5010
rect 2984 5198 3122 5266
rect 3202 5508 3236 5524
rect 3202 5344 3236 5432
rect 3298 5508 3332 5574
rect 3298 5416 3332 5432
rect 3394 5508 3428 5524
rect 3394 5350 3428 5432
rect 3490 5508 3524 5574
rect 3490 5416 3524 5432
rect 3506 5350 3566 5360
rect 3394 5348 3578 5350
rect 3202 5327 3360 5344
rect 3202 5293 3324 5327
rect 3358 5293 3360 5327
rect 3202 5276 3360 5293
rect 3394 5312 3512 5348
rect 3548 5312 3578 5348
rect 2078 4876 2222 4886
rect 906 4844 1516 4858
rect 2258 4850 2282 4886
rect 2318 4850 2374 4886
rect 2410 4850 2466 4886
rect 2502 4850 2558 4886
rect 2594 4850 2650 4886
rect 2686 4850 2710 4886
rect 2258 4848 2710 4850
rect 2984 4848 3064 5198
rect 3202 5182 3236 5276
rect 3202 4990 3236 5006
rect 3298 5182 3332 5198
rect 3298 4926 3332 5006
rect 3394 5182 3428 5312
rect 3506 5300 3566 5312
rect 3394 4990 3428 5006
rect 3490 5182 3524 5198
rect 3490 4926 3524 5006
rect 3612 4926 3668 6326
rect 3738 6292 3804 6300
rect 3738 6258 3754 6292
rect 3788 6258 3804 6292
rect 3738 6248 3804 6258
rect 3738 6198 3772 6214
rect 3738 5868 3772 6062
rect 3834 6198 3868 6214
rect 3834 6046 3868 6062
rect 3930 6198 3964 6334
rect 4234 6294 4300 6300
rect 4234 6258 4250 6294
rect 4284 6258 4300 6294
rect 4234 6248 4300 6258
rect 3930 6046 3964 6062
rect 4026 6198 4060 6214
rect 4026 6046 4060 6062
rect 4122 6198 4156 6214
rect 3854 6002 3920 6010
rect 3854 5968 3870 6002
rect 3904 5968 3920 6002
rect 3854 5958 3920 5968
rect 4122 5952 4156 6062
rect 4234 6198 4268 6214
rect 4122 5946 4170 5952
rect 4122 5942 4130 5946
rect 3950 5912 4130 5942
rect 4164 5912 4170 5946
rect 3950 5904 4170 5912
rect 3950 5884 3984 5904
rect 3738 5792 3772 5808
rect 3834 5868 3868 5884
rect 3834 5744 3868 5808
rect 3930 5868 3984 5884
rect 3964 5808 3984 5868
rect 3930 5792 3984 5808
rect 4234 5868 4268 6062
rect 4330 6198 4364 6214
rect 4330 6046 4364 6062
rect 4426 6198 4460 6334
rect 4426 6046 4460 6062
rect 4522 6198 4556 6214
rect 4522 6046 4556 6062
rect 4618 6198 4652 6214
rect 4350 6002 4416 6010
rect 4350 5968 4366 6002
rect 4400 5968 4416 6002
rect 4350 5958 4416 5968
rect 4618 5942 4652 6062
rect 4710 6088 4908 6626
rect 4710 6014 4768 6088
rect 4842 6014 4908 6088
rect 4446 5936 4676 5942
rect 4446 5904 4554 5936
rect 4446 5884 4480 5904
rect 4542 5900 4554 5904
rect 4590 5900 4628 5936
rect 4664 5900 4676 5936
rect 4542 5894 4676 5900
rect 4234 5792 4268 5808
rect 4330 5868 4364 5884
rect 4330 5744 4364 5808
rect 4426 5868 4480 5884
rect 4460 5808 4480 5868
rect 4426 5792 4480 5808
rect 4710 5744 4908 6014
rect 3808 5742 4908 5744
rect 3702 5726 3750 5742
rect 3702 5692 3710 5726
rect 3744 5692 3750 5726
rect 3808 5708 3834 5742
rect 3868 5708 4330 5742
rect 4364 5708 4908 5742
rect 3808 5692 4908 5708
rect 3702 5360 3750 5692
rect 3702 5324 3708 5360
rect 3744 5324 3750 5360
rect 3702 5008 3750 5324
rect 3784 5636 3832 5648
rect 3784 5600 3790 5636
rect 3826 5600 3832 5636
rect 3784 5300 3832 5600
rect 3970 5548 4056 5692
rect 3970 5514 3994 5548
rect 4028 5514 4056 5548
rect 4710 5614 4908 5692
rect 4710 5540 4768 5614
rect 4842 5540 4908 5614
rect 3784 5264 3790 5300
rect 3826 5264 3832 5300
rect 3784 5252 3832 5264
rect 3898 5448 3932 5464
rect 3898 5194 3932 5388
rect 3994 5448 4028 5514
rect 3994 5372 4028 5388
rect 4090 5448 4144 5464
rect 4124 5388 4144 5448
rect 4090 5372 4144 5388
rect 4110 5352 4144 5372
rect 4110 5346 4516 5352
rect 4110 5314 4392 5346
rect 4014 5288 4080 5298
rect 4014 5254 4030 5288
rect 4064 5254 4080 5288
rect 4014 5246 4080 5254
rect 3898 5042 3932 5058
rect 3994 5194 4028 5210
rect 3994 5042 4028 5058
rect 4090 5194 4124 5210
rect 3702 4998 3964 5008
rect 3702 4964 3914 4998
rect 3948 4964 3964 4998
rect 3702 4956 3964 4964
rect 3122 4888 3214 4926
rect 3252 4888 3290 4926
rect 3328 4888 3366 4926
rect 3404 4888 3442 4926
rect 3480 4922 3668 4926
rect 4090 4922 4124 5058
rect 4186 5194 4220 5210
rect 4186 5042 4220 5058
rect 4282 5194 4316 5314
rect 4380 5310 4392 5314
rect 4428 5310 4468 5346
rect 4504 5310 4516 5346
rect 4380 5304 4516 5310
rect 4282 5042 4316 5058
rect 4710 5140 4908 5540
rect 4710 5066 4768 5140
rect 4842 5066 4908 5140
rect 4710 4952 4908 5066
rect 3480 4888 3954 4922
rect 3988 4888 4022 4922
rect 4056 4888 4090 4922
rect 4124 4888 4158 4922
rect 4192 4888 4226 4922
rect 4260 4888 4288 4922
rect 4710 4918 4724 4952
rect 4758 4918 4796 4952
rect 4830 4918 4868 4952
rect 4902 4918 4908 4952
rect 4710 4880 4908 4918
rect 30 4774 46 4808
rect 80 4774 118 4808
rect 152 4774 190 4808
rect 224 4774 228 4808
rect 792 4842 1610 4844
rect 792 4806 816 4842
rect 852 4806 934 4842
rect 970 4806 1052 4842
rect 1088 4806 1170 4842
rect 1206 4806 1288 4842
rect 1324 4806 1406 4842
rect 1442 4806 1524 4842
rect 1560 4806 1610 4842
rect 792 4802 1610 4806
rect 2984 4830 3956 4848
rect 2984 4828 3066 4830
rect 30 4736 228 4774
rect 30 4702 46 4736
rect 80 4702 118 4736
rect 152 4702 190 4736
rect 224 4702 228 4736
rect 30 4664 228 4702
rect 30 4630 44 4664
rect 78 4630 116 4664
rect 150 4630 188 4664
rect 222 4630 228 4664
rect 30 4564 228 4630
rect 30 4134 48 4564
rect 206 4134 228 4564
rect 916 4504 1376 4802
rect 2984 4792 2992 4828
rect 3028 4794 3066 4828
rect 3102 4794 3146 4830
rect 3182 4794 3226 4830
rect 3262 4794 3306 4830
rect 3342 4794 3956 4830
rect 3028 4792 3956 4794
rect 2984 4778 3956 4792
rect 3496 4504 3956 4778
rect 4710 4846 4724 4880
rect 4758 4846 4796 4880
rect 4830 4846 4868 4880
rect 4902 4846 4908 4880
rect 4710 4808 4908 4846
rect 4710 4774 4724 4808
rect 4758 4774 4796 4808
rect 4830 4774 4868 4808
rect 4902 4774 4908 4808
rect 4710 4736 4908 4774
rect 4710 4702 4724 4736
rect 4758 4702 4796 4736
rect 4830 4702 4868 4736
rect 4902 4702 4908 4736
rect 4710 4664 4908 4702
rect 4710 4630 4724 4664
rect 4758 4630 4796 4664
rect 4830 4630 4868 4664
rect 4902 4630 4908 4664
rect 30 4014 228 4134
rect 30 3574 56 4014
rect 186 3574 228 4014
rect 30 3486 228 3574
rect 30 3444 94 3486
rect 168 3444 228 3486
rect 30 3034 56 3444
rect 216 3034 228 3444
rect 346 4484 4526 4504
rect 346 4434 946 4484
rect 1346 4434 3526 4484
rect 3926 4434 4526 4484
rect 346 4424 4526 4434
rect 346 3164 426 4424
rect 916 4414 1376 4424
rect 3496 4414 3956 4424
rect 586 4204 606 4304
rect 726 4204 766 4304
rect 886 4204 926 4304
rect 1046 4204 1086 4304
rect 1206 4204 1246 4304
rect 1366 4204 1406 4304
rect 1526 4204 1566 4304
rect 1686 4204 3186 4304
rect 3306 4204 3346 4304
rect 3466 4204 3506 4304
rect 3626 4204 3666 4304
rect 3786 4204 3826 4304
rect 3946 4204 3986 4304
rect 4106 4204 4146 4304
rect 4266 4204 4286 4304
rect 586 4184 4286 4204
rect 506 4104 1066 4144
rect 506 4054 616 4104
rect 1106 4064 1176 4184
rect 556 4004 616 4054
rect 656 4024 1176 4064
rect 506 3984 616 4004
rect 506 3964 1066 3984
rect 576 3944 1066 3964
rect 576 3914 616 3944
rect 506 3874 616 3914
rect 1106 3904 1176 4024
rect 576 3824 616 3874
rect 656 3864 1176 3904
rect 1216 3834 1256 4144
rect 1296 3884 1336 4184
rect 1376 3834 1416 4144
rect 1456 3884 1496 4184
rect 1536 3834 1576 4144
rect 1616 3884 1656 4184
rect 1696 3834 1736 4144
rect 1776 3884 1816 4184
rect 1856 3834 1896 4144
rect 1936 3884 1976 4184
rect 2016 3834 2056 4144
rect 2096 3884 2136 4184
rect 2176 3834 2216 4144
rect 2256 3884 2296 4184
rect 2336 3834 2376 4144
rect 2416 3884 2456 4184
rect 2496 3834 2536 4144
rect 2576 3884 2616 4184
rect 2656 3834 2696 4144
rect 2736 3884 2776 4184
rect 2816 3834 2856 4144
rect 2896 3884 2936 4184
rect 2976 3834 3016 4144
rect 3056 3884 3096 4184
rect 3136 3834 3176 4144
rect 3216 3884 3256 4184
rect 3296 3834 3336 4144
rect 3376 3884 3416 4184
rect 3456 3834 3496 4144
rect 3536 3884 3576 4184
rect 3616 3834 3656 4144
rect 3696 4064 3766 4184
rect 3806 4104 4366 4144
rect 3696 4024 4216 4064
rect 4256 4044 4366 4104
rect 3696 3904 3766 4024
rect 4256 3994 4316 4044
rect 4256 3984 4366 3994
rect 3806 3954 4366 3984
rect 3806 3944 4296 3954
rect 4256 3904 4296 3944
rect 3696 3864 4206 3904
rect 4256 3864 4366 3904
rect 1216 3824 3656 3834
rect 4256 3824 4296 3864
rect 506 3814 4296 3824
rect 506 3774 4366 3814
rect 576 3764 4366 3774
rect 576 3724 616 3764
rect 1216 3754 3656 3764
rect 506 3684 616 3724
rect 656 3684 1176 3724
rect 576 3644 616 3684
rect 576 3634 1066 3644
rect 506 3604 1066 3634
rect 506 3594 616 3604
rect 556 3544 616 3594
rect 1106 3564 1176 3684
rect 506 3484 616 3544
rect 656 3524 1176 3564
rect 506 3444 1066 3484
rect 1106 3404 1176 3524
rect 1216 3444 1256 3754
rect 1296 3404 1336 3704
rect 1376 3444 1416 3754
rect 1456 3404 1496 3704
rect 1536 3444 1576 3754
rect 1616 3404 1656 3704
rect 1696 3444 1736 3754
rect 1776 3404 1816 3704
rect 1856 3444 1896 3754
rect 1936 3404 1976 3704
rect 2016 3444 2056 3754
rect 2096 3404 2136 3704
rect 2176 3444 2216 3754
rect 2256 3404 2296 3704
rect 2336 3454 2376 3754
rect 2416 3404 2456 3704
rect 2496 3454 2536 3754
rect 2576 3404 2616 3704
rect 2656 3444 2696 3754
rect 2736 3404 2776 3704
rect 2816 3444 2856 3754
rect 2896 3404 2936 3704
rect 2976 3444 3016 3754
rect 3056 3404 3096 3704
rect 3136 3444 3176 3754
rect 3216 3404 3256 3704
rect 3296 3444 3336 3754
rect 3376 3404 3416 3704
rect 3456 3444 3496 3754
rect 3536 3404 3576 3704
rect 3616 3444 3656 3754
rect 3696 3684 4206 3724
rect 4256 3714 4296 3764
rect 3696 3564 3766 3684
rect 4256 3674 4366 3714
rect 4256 3644 4296 3674
rect 3806 3624 4296 3644
rect 3806 3604 4366 3624
rect 4256 3584 4366 3604
rect 3696 3524 4216 3564
rect 4256 3534 4316 3584
rect 3696 3404 3766 3524
rect 4256 3484 4366 3534
rect 3806 3444 4366 3484
rect 586 3384 4286 3404
rect 586 3284 606 3384
rect 726 3284 766 3384
rect 886 3284 926 3384
rect 1046 3284 1086 3384
rect 1206 3284 1246 3384
rect 1366 3284 1406 3384
rect 1526 3284 1566 3384
rect 1686 3284 3186 3384
rect 3306 3284 3346 3384
rect 3466 3284 3506 3384
rect 3626 3284 3666 3384
rect 3786 3284 3826 3384
rect 3946 3284 3986 3384
rect 4106 3284 4146 3384
rect 4266 3284 4286 3384
rect 916 3164 1376 3174
rect 3496 3164 3956 3174
rect 4446 3164 4526 4424
rect 346 3154 4526 3164
rect 346 3104 946 3154
rect 1346 3104 3526 3154
rect 3926 3104 4526 3154
rect 346 3084 4526 3104
rect 4710 4404 4908 4630
rect 4710 4330 4768 4404
rect 4842 4330 4908 4404
rect 4710 3930 4908 4330
rect 4710 3856 4768 3930
rect 4842 3856 4908 3930
rect 4710 3456 4908 3856
rect 4710 3382 4768 3456
rect 4842 3382 4908 3456
rect 30 2994 228 3034
rect 916 2994 1376 3084
rect 3496 2994 3956 3084
rect 4710 2994 4908 3382
rect 30 2926 4908 2994
rect 30 2852 624 2926
rect 698 2852 1172 2926
rect 1246 2852 1720 2926
rect 1794 2852 2268 2926
rect 2342 2852 2816 2926
rect 2890 2852 3364 2926
rect 3438 2852 3914 2926
rect 3988 2852 4908 2926
rect 30 2796 4908 2852
<< viali >>
rect 66 8120 88 8144
rect 88 8120 162 8144
rect 162 8120 196 8144
rect 66 7744 196 8120
rect 50 7246 186 7604
rect 50 7172 88 7246
rect 88 7172 162 7246
rect 162 7172 186 7246
rect 50 7164 186 7172
rect 50 6772 206 7044
rect 50 6698 88 6772
rect 88 6698 162 6772
rect 162 6698 206 6772
rect 50 6614 206 6698
rect 606 7794 726 7894
rect 766 7794 886 7894
rect 926 7794 1046 7894
rect 1086 7794 1206 7894
rect 3666 7794 3786 7894
rect 3826 7794 3946 7894
rect 3986 7794 4106 7894
rect 4146 7794 4266 7894
rect 526 7504 556 7554
rect 556 7504 576 7554
rect 526 7414 556 7464
rect 556 7414 576 7464
rect 4296 7494 4316 7544
rect 4316 7494 4346 7544
rect 4296 7404 4316 7454
rect 4316 7404 4346 7454
rect 526 7314 556 7364
rect 556 7314 576 7364
rect 526 7224 556 7274
rect 556 7224 576 7274
rect 4296 7304 4316 7354
rect 4316 7304 4346 7354
rect 4296 7214 4316 7264
rect 4316 7214 4346 7264
rect 606 6874 726 6974
rect 766 6874 886 6974
rect 926 6874 1046 6974
rect 1086 6874 1206 6974
rect 3666 6874 3786 6974
rect 3826 6874 3946 6974
rect 3986 6874 4106 6974
rect 4146 6874 4266 6974
rect 3214 6368 3250 6404
rect 3290 6368 3326 6404
rect 3366 6368 3402 6404
rect 3442 6368 3478 6404
rect 3518 6368 3554 6404
rect 3594 6368 3630 6404
rect 594 6240 628 6276
rect 672 6240 706 6276
rect 744 6240 778 6276
rect 828 6240 862 6274
rect 912 6240 946 6274
rect 996 6240 1030 6274
rect 1080 6240 1114 6274
rect 1164 6240 1198 6274
rect 1248 6240 1282 6274
rect 1332 6240 1366 6274
rect 1416 6240 1450 6274
rect 1500 6240 1534 6274
rect 1590 6240 1624 6274
rect 2136 6250 2170 6284
rect 2220 6250 2254 6284
rect 2304 6250 2338 6284
rect 2388 6250 2422 6284
rect 2472 6250 2506 6284
rect 2556 6250 2590 6284
rect 2640 6250 2674 6284
rect 2724 6250 2758 6284
rect 1726 6074 1876 6224
rect 374 5574 410 5608
rect 608 5574 644 5608
rect 362 5440 422 5474
rect 596 5440 656 5474
rect 362 5258 422 5292
rect 596 5258 656 5292
rect 278 5170 312 5204
rect 512 5170 546 5204
rect 992 5800 1032 5840
rect 1090 5774 1126 5810
rect 1384 5850 1424 5890
rect 1832 5844 1868 5880
rect 1832 5770 1868 5806
rect 1832 5696 1868 5732
rect 1832 5586 1868 5622
rect 3126 5936 3162 5970
rect 3126 5864 3162 5898
rect 3508 5902 3544 5938
rect 1832 5510 1868 5546
rect 1832 5436 1868 5472
rect 46 4918 80 4952
rect 118 4918 152 4952
rect 190 4918 224 4952
rect 374 4908 410 4942
rect 608 4908 644 4942
rect 46 4846 80 4880
rect 118 4846 152 4880
rect 190 4846 224 4880
rect 1826 4994 1976 5144
rect 2094 4886 2128 4920
rect 2172 4886 2206 4920
rect 2834 5454 2870 5490
rect 2908 5454 2944 5490
rect 3512 5312 3548 5348
rect 2282 4850 2318 4886
rect 2374 4850 2410 4886
rect 2466 4850 2502 4886
rect 2558 4850 2594 4886
rect 2650 4850 2686 4886
rect 4250 6292 4284 6294
rect 4250 6260 4284 6292
rect 3870 5968 3904 6002
rect 4130 5912 4164 5946
rect 3738 5808 3772 5868
rect 3930 5808 3964 5868
rect 4366 5968 4400 6002
rect 4554 5900 4590 5936
rect 4628 5900 4664 5936
rect 4234 5808 4268 5868
rect 4426 5808 4460 5868
rect 3708 5324 3744 5360
rect 3790 5600 3826 5636
rect 3790 5264 3826 5300
rect 3898 5388 3932 5448
rect 4090 5388 4124 5448
rect 4030 5254 4064 5288
rect 4392 5310 4428 5346
rect 4468 5310 4504 5346
rect 4724 4918 4758 4952
rect 4796 4918 4830 4952
rect 4868 4918 4902 4952
rect 46 4774 80 4808
rect 118 4774 152 4808
rect 190 4774 224 4808
rect 816 4806 852 4842
rect 934 4806 970 4842
rect 1052 4806 1088 4842
rect 1170 4806 1206 4842
rect 1288 4806 1324 4842
rect 1406 4806 1442 4842
rect 1524 4806 1560 4842
rect 46 4702 80 4736
rect 118 4702 152 4736
rect 190 4702 224 4736
rect 44 4630 78 4664
rect 116 4630 150 4664
rect 188 4630 222 4664
rect 48 4434 206 4564
rect 48 4360 94 4434
rect 94 4360 168 4434
rect 168 4360 206 4434
rect 48 4134 206 4360
rect 2992 4792 3028 4828
rect 3066 4794 3102 4830
rect 3146 4794 3182 4830
rect 3226 4794 3262 4830
rect 3306 4794 3342 4830
rect 4724 4846 4758 4880
rect 4796 4846 4830 4880
rect 4868 4846 4902 4880
rect 4724 4774 4758 4808
rect 4796 4774 4830 4808
rect 4868 4774 4902 4808
rect 4724 4702 4758 4736
rect 4796 4702 4830 4736
rect 4868 4702 4902 4736
rect 4724 4630 4758 4664
rect 4796 4630 4830 4664
rect 4868 4630 4902 4664
rect 56 3960 186 4014
rect 56 3886 94 3960
rect 94 3886 168 3960
rect 168 3886 186 3960
rect 56 3574 186 3886
rect 56 3412 94 3444
rect 94 3412 168 3444
rect 168 3412 216 3444
rect 56 3034 216 3412
rect 606 4204 726 4304
rect 766 4204 886 4304
rect 926 4204 1046 4304
rect 1086 4204 1206 4304
rect 3666 4204 3786 4304
rect 3826 4204 3946 4304
rect 3986 4204 4106 4304
rect 4146 4204 4266 4304
rect 526 3914 556 3964
rect 556 3914 576 3964
rect 526 3824 556 3874
rect 556 3824 576 3874
rect 4296 3904 4316 3954
rect 4316 3904 4346 3954
rect 4296 3814 4316 3864
rect 4316 3814 4346 3864
rect 526 3724 556 3774
rect 556 3724 576 3774
rect 526 3634 556 3684
rect 556 3634 576 3684
rect 4296 3714 4316 3764
rect 4316 3714 4346 3764
rect 4296 3624 4316 3674
rect 4316 3624 4346 3674
rect 606 3284 726 3384
rect 766 3284 886 3384
rect 926 3284 1046 3384
rect 1086 3284 1206 3384
rect 3666 3284 3786 3384
rect 3826 3284 3946 3384
rect 3986 3284 4106 3384
rect 4146 3284 4266 3384
<< metal1 >>
rect 30 8154 906 8174
rect 30 8144 286 8154
rect 30 7744 66 8144
rect 196 7954 286 8144
rect 486 7954 686 8154
rect 886 7954 906 8154
rect 196 7934 906 7954
rect 1386 8154 3486 8174
rect 1386 7954 1406 8154
rect 1606 7954 1626 8154
rect 1826 7954 2346 8154
rect 2526 7954 3046 8154
rect 3246 7954 3266 8154
rect 3466 7954 3486 8154
rect 1386 7934 3486 7954
rect 3966 8154 4606 8174
rect 3966 7954 3986 8154
rect 4186 7954 4386 8154
rect 4586 7954 4606 8154
rect 3966 7934 4606 7954
rect 196 7904 726 7934
rect 196 7894 2346 7904
rect 196 7834 606 7894
rect 196 7744 286 7834
rect 30 7704 286 7744
rect 266 7634 286 7704
rect 486 7794 606 7834
rect 726 7794 766 7894
rect 886 7794 926 7894
rect 1046 7794 1086 7894
rect 1206 7874 2346 7894
rect 1206 7794 1226 7874
rect 2376 7844 2496 7934
rect 4146 7904 4606 7934
rect 2526 7894 4606 7904
rect 2526 7874 3666 7894
rect 1256 7814 3616 7844
rect 486 7784 1226 7794
rect 486 7634 506 7784
rect 596 7774 2346 7784
rect 30 7604 206 7624
rect 266 7604 506 7634
rect 30 7164 50 7604
rect 186 7164 206 7604
rect 266 7554 596 7574
rect 266 7544 526 7554
rect 266 7434 286 7544
rect 486 7504 526 7544
rect 576 7504 596 7554
rect 626 7504 656 7774
rect 486 7464 596 7504
rect 486 7434 526 7464
rect 266 7414 526 7434
rect 576 7444 596 7464
rect 686 7444 716 7744
rect 746 7504 776 7774
rect 806 7444 836 7744
rect 866 7504 896 7774
rect 926 7444 956 7744
rect 986 7504 1016 7774
rect 1106 7754 2346 7774
rect 1046 7444 1076 7744
rect 1106 7664 1226 7754
rect 2376 7724 2496 7814
rect 3646 7794 3666 7874
rect 3786 7794 3826 7894
rect 3946 7794 3986 7894
rect 4106 7794 4146 7894
rect 4266 7834 4606 7894
rect 4266 7794 4386 7834
rect 3646 7784 4386 7794
rect 2526 7774 4276 7784
rect 2526 7754 3766 7774
rect 1256 7694 3616 7724
rect 1106 7634 2346 7664
rect 1106 7544 1226 7634
rect 2376 7604 2496 7694
rect 3646 7664 3766 7754
rect 2526 7634 3766 7664
rect 1256 7574 3616 7604
rect 1106 7514 2346 7544
rect 1106 7474 1226 7514
rect 2376 7484 2496 7574
rect 3646 7544 3766 7634
rect 2526 7514 3766 7544
rect 1256 7454 3616 7484
rect 3646 7474 3766 7514
rect 576 7424 1076 7444
rect 2376 7424 2496 7454
rect 3796 7444 3826 7744
rect 3856 7504 3886 7774
rect 3916 7444 3946 7744
rect 3976 7504 4006 7774
rect 4036 7444 4066 7744
rect 4096 7504 4126 7774
rect 4156 7444 4186 7744
rect 4216 7504 4246 7774
rect 4366 7634 4386 7784
rect 4586 7634 4606 7834
rect 4366 7604 4606 7634
rect 4276 7544 4606 7564
rect 4276 7494 4296 7544
rect 4346 7494 4386 7544
rect 4276 7454 4386 7494
rect 4276 7444 4296 7454
rect 3796 7424 4296 7444
rect 576 7414 4296 7424
rect 266 7404 4296 7414
rect 4346 7434 4386 7454
rect 4586 7434 4606 7544
rect 4346 7404 4606 7434
rect 266 7364 4606 7404
rect 266 7334 526 7364
rect 266 7224 286 7334
rect 486 7314 526 7334
rect 576 7354 4606 7364
rect 576 7314 4296 7354
rect 486 7304 4296 7314
rect 4346 7334 4606 7354
rect 4346 7304 4386 7334
rect 486 7284 4386 7304
rect 486 7274 596 7284
rect 486 7224 526 7274
rect 576 7224 596 7274
rect 266 7204 596 7224
rect 30 7144 206 7164
rect 266 7134 506 7164
rect 266 7064 286 7134
rect 30 7044 286 7064
rect 30 6614 50 7044
rect 206 6934 286 7044
rect 486 6984 506 7134
rect 626 6994 656 7254
rect 686 7024 716 7284
rect 746 6994 776 7254
rect 806 7024 836 7284
rect 866 6994 896 7254
rect 926 7024 956 7284
rect 986 6994 1016 7254
rect 1046 7024 1076 7284
rect 1106 7224 2346 7254
rect 1106 7134 1226 7224
rect 2376 7194 2496 7284
rect 2526 7224 3766 7254
rect 1256 7164 3616 7194
rect 1106 7104 2346 7134
rect 1106 7014 1226 7104
rect 2376 7074 2496 7164
rect 3646 7134 3766 7224
rect 2526 7104 3766 7134
rect 1256 7044 3616 7074
rect 1106 6994 2346 7014
rect 596 6984 2346 6994
rect 486 6974 1226 6984
rect 486 6934 606 6974
rect 206 6874 606 6934
rect 726 6874 766 6974
rect 886 6874 926 6974
rect 1046 6874 1086 6974
rect 1206 6894 1226 6974
rect 2376 6954 2496 7044
rect 3646 7014 3766 7104
rect 3796 7024 3826 7284
rect 2526 6994 3766 7014
rect 3856 6994 3886 7254
rect 3916 7024 3946 7284
rect 3976 6994 4006 7254
rect 4036 7024 4066 7284
rect 4096 6994 4126 7254
rect 4156 7024 4186 7284
rect 4276 7264 4386 7284
rect 4216 6994 4246 7254
rect 4276 7214 4296 7264
rect 4346 7224 4386 7264
rect 4586 7224 4606 7334
rect 4346 7214 4606 7224
rect 4276 7194 4606 7214
rect 4366 7134 4606 7164
rect 2526 6984 4276 6994
rect 4366 6984 4386 7134
rect 3646 6974 4386 6984
rect 1256 6924 3616 6954
rect 1206 6874 2346 6894
rect 206 6864 2346 6874
rect 206 6834 726 6864
rect 2376 6834 2496 6924
rect 3646 6894 3666 6974
rect 2526 6874 3666 6894
rect 3786 6874 3826 6974
rect 3946 6874 3986 6974
rect 4106 6874 4146 6974
rect 4266 6934 4386 6974
rect 4586 6934 4606 7134
rect 4266 6874 4606 6934
rect 2526 6864 4606 6874
rect 4146 6834 4606 6864
rect 206 6814 906 6834
rect 206 6614 286 6814
rect 486 6614 686 6814
rect 886 6614 906 6814
rect 30 6594 906 6614
rect 1386 6814 3486 6834
rect 1386 6614 1406 6814
rect 1606 6614 1626 6814
rect 1826 6614 2346 6814
rect 2526 6614 3046 6814
rect 3246 6614 3266 6814
rect 3466 6614 3486 6814
rect 1386 6594 3486 6614
rect 3966 6814 4606 6834
rect 3966 6614 3986 6814
rect 4186 6614 4386 6814
rect 4586 6614 4606 6814
rect 3966 6594 4606 6614
rect -558 6544 5426 6566
rect -558 6354 -494 6544
rect -334 6404 5246 6544
rect -334 6368 3214 6404
rect 3250 6368 3290 6404
rect 3326 6368 3366 6404
rect 3402 6368 3442 6404
rect 3478 6368 3518 6404
rect 3554 6368 3594 6404
rect 3630 6368 5246 6404
rect -334 6354 5246 6368
rect 5406 6354 5426 6544
rect -558 6336 5426 6354
rect 582 6276 1654 6336
rect 582 6240 594 6276
rect 628 6240 672 6276
rect 706 6240 744 6276
rect 778 6274 1654 6276
rect 778 6240 828 6274
rect 862 6240 912 6274
rect 946 6240 996 6274
rect 1030 6240 1080 6274
rect 1114 6240 1164 6274
rect 1198 6240 1248 6274
rect 1282 6240 1332 6274
rect 1366 6240 1416 6274
rect 1450 6240 1500 6274
rect 1534 6240 1590 6274
rect 1624 6240 1654 6274
rect 2098 6284 2822 6336
rect 2098 6250 2136 6284
rect 2170 6250 2220 6284
rect 2254 6250 2304 6284
rect 2338 6250 2388 6284
rect 2422 6250 2472 6284
rect 2506 6250 2556 6284
rect 2590 6250 2640 6284
rect 2674 6250 2724 6284
rect 2758 6250 2822 6284
rect 2098 6244 2822 6250
rect 3562 6300 3806 6306
rect 3562 6294 4296 6300
rect 3562 6272 4250 6294
rect 582 6234 1654 6240
rect 1706 6224 1896 6244
rect 1706 6074 1726 6224
rect 1876 6074 1896 6224
rect 1706 6054 1896 6074
rect 3112 5970 3168 5986
rect 3112 5936 3126 5970
rect 3162 5936 3168 5970
rect 3562 5950 3598 6272
rect 4234 6260 4250 6272
rect 4284 6260 4296 6294
rect 4234 6254 4296 6260
rect 3854 6006 3920 6010
rect 4350 6008 4416 6010
rect 4338 6006 4656 6008
rect 3722 6002 4080 6006
rect 3722 5970 3870 6002
rect 3854 5968 3870 5970
rect 3904 5970 4080 6002
rect 3904 5968 3920 5970
rect 3854 5958 3920 5968
rect -558 5890 1440 5906
rect 3112 5898 3168 5936
rect -558 5878 1384 5890
rect 1368 5850 1384 5878
rect 1424 5850 1440 5890
rect -558 5840 1048 5850
rect 1368 5840 1440 5850
rect 1820 5880 1880 5890
rect 1820 5844 1832 5880
rect 1868 5844 1880 5880
rect 3112 5864 3126 5898
rect 3162 5864 3168 5898
rect 3502 5938 3598 5950
rect 3502 5902 3508 5938
rect 3544 5902 3598 5938
rect 3502 5890 3598 5902
rect 3112 5846 3168 5864
rect -558 5822 992 5840
rect 976 5800 992 5822
rect 1032 5800 1048 5840
rect 976 5790 1048 5800
rect 1078 5812 1132 5816
rect 1820 5812 1880 5844
rect 1078 5810 1880 5812
rect 1078 5798 1090 5810
rect 1076 5774 1090 5798
rect 1126 5806 1880 5810
rect 1126 5774 1832 5806
rect 1076 5770 1832 5774
rect 1868 5770 1880 5806
rect 1076 5760 1880 5770
rect 1820 5732 1880 5760
rect 1820 5696 1832 5732
rect 1868 5696 1880 5732
rect 1820 5690 1880 5696
rect 3562 5648 3598 5890
rect 3732 5868 3778 5880
rect 3732 5808 3738 5868
rect 3772 5852 3778 5868
rect 3924 5868 3970 5880
rect 3924 5852 3930 5868
rect 3772 5824 3930 5852
rect 3772 5808 3778 5824
rect 3732 5796 3778 5808
rect 3924 5808 3930 5824
rect 3964 5808 3970 5868
rect 4044 5858 4080 5970
rect 4134 6002 4656 6006
rect 4134 5970 4366 6002
rect 4134 5958 4170 5970
rect 4350 5968 4366 5970
rect 4400 6000 4656 6002
rect 4400 5972 5452 6000
rect 4400 5968 4416 5972
rect 4350 5958 4416 5968
rect 4122 5946 4170 5958
rect 4122 5912 4130 5946
rect 4164 5912 4170 5946
rect 4122 5900 4170 5912
rect 4542 5936 4676 5942
rect 4542 5900 4554 5936
rect 4590 5900 4628 5936
rect 4664 5932 4676 5936
rect 4664 5904 5452 5932
rect 4664 5900 4676 5904
rect 4542 5894 4676 5900
rect 4228 5868 4274 5880
rect 4228 5858 4234 5868
rect 4044 5822 4234 5858
rect 3924 5796 3970 5808
rect 4228 5808 4234 5822
rect 4268 5852 4274 5868
rect 4420 5868 4466 5880
rect 4420 5852 4426 5868
rect 4268 5824 4426 5852
rect 4268 5808 4274 5824
rect 4228 5796 4274 5808
rect 4420 5808 4426 5824
rect 4460 5808 4466 5868
rect 4420 5796 4466 5808
rect 3562 5636 3832 5648
rect 1820 5622 1880 5628
rect 342 5608 440 5614
rect 342 5574 374 5608
rect 410 5574 440 5608
rect 342 5568 440 5574
rect 576 5608 674 5614
rect 576 5574 608 5608
rect 644 5574 674 5608
rect 576 5568 674 5574
rect 1820 5586 1832 5622
rect 1868 5586 1880 5622
rect 3562 5610 3790 5636
rect 3784 5600 3790 5610
rect 3826 5600 3832 5636
rect 3784 5588 3832 5600
rect 1820 5546 1880 5586
rect 1820 5510 1832 5546
rect 1868 5510 1880 5546
rect 354 5474 432 5488
rect 354 5440 362 5474
rect 422 5440 432 5474
rect 354 5292 432 5440
rect 354 5258 362 5292
rect 422 5258 432 5292
rect 354 5246 432 5258
rect 588 5474 666 5488
rect 588 5440 596 5474
rect 656 5440 666 5474
rect 588 5292 666 5440
rect 1820 5474 1880 5510
rect 2824 5490 2954 5506
rect 2824 5474 2834 5490
rect 1820 5472 2834 5474
rect 1820 5436 1832 5472
rect 1868 5454 2834 5472
rect 2870 5454 2908 5490
rect 2944 5454 2954 5490
rect 1868 5438 2954 5454
rect 3892 5448 3938 5460
rect 1868 5436 1880 5438
rect 1820 5430 1880 5436
rect 3892 5388 3898 5448
rect 3932 5432 3938 5448
rect 4084 5448 4130 5460
rect 4084 5432 4090 5448
rect 3932 5404 4090 5432
rect 3932 5388 3938 5404
rect 3892 5376 3938 5388
rect 4084 5388 4090 5404
rect 4124 5388 4130 5448
rect 4084 5376 4130 5388
rect 3702 5360 3750 5372
rect 3506 5350 3566 5360
rect 3702 5350 3708 5360
rect 3506 5348 3708 5350
rect 3506 5312 3512 5348
rect 3548 5324 3708 5348
rect 3744 5324 3750 5360
rect 3548 5312 3750 5324
rect 4380 5346 4516 5352
rect 3506 5300 3566 5312
rect 3784 5300 3832 5312
rect 4380 5310 4392 5346
rect 4428 5310 4468 5346
rect 4504 5342 4516 5346
rect 4504 5314 5452 5342
rect 4504 5310 4516 5314
rect 4380 5304 4516 5310
rect 588 5258 596 5292
rect 656 5258 666 5292
rect 588 5246 666 5258
rect 3784 5264 3790 5300
rect 3826 5286 3832 5300
rect 4014 5288 4080 5298
rect 4014 5286 4030 5288
rect 3826 5264 4030 5286
rect 3784 5254 4030 5264
rect 4064 5254 4080 5288
rect 3784 5250 4080 5254
rect 3784 5248 3882 5250
rect 4014 5246 4080 5250
rect 256 5204 318 5220
rect 256 5202 278 5204
rect -558 5174 278 5202
rect 256 5170 278 5174
rect 312 5170 318 5204
rect 256 5154 318 5170
rect 496 5204 552 5220
rect 496 5170 512 5204
rect 546 5186 552 5204
rect 546 5170 756 5186
rect 496 5154 756 5170
rect 30 4952 230 4972
rect 30 4918 46 4952
rect 80 4918 118 4952
rect 152 4918 190 4952
rect 224 4942 684 4952
rect 224 4918 374 4942
rect 30 4908 374 4918
rect 410 4908 608 4942
rect 644 4908 684 4942
rect 30 4880 684 4908
rect 30 4848 46 4880
rect -558 4846 46 4848
rect 80 4846 118 4880
rect 152 4846 190 4880
rect 224 4848 684 4880
rect 714 4930 756 5154
rect 1806 5144 1996 5164
rect 1806 4994 1826 5144
rect 1976 4994 1996 5144
rect 1806 4974 1996 4994
rect 4710 4952 4908 4972
rect 714 4920 2222 4930
rect 714 4886 2094 4920
rect 2128 4886 2172 4920
rect 2206 4886 2222 4920
rect 4710 4918 4724 4952
rect 4758 4918 4796 4952
rect 4830 4918 4868 4952
rect 4902 4918 4908 4952
rect 714 4876 2222 4886
rect 2258 4886 2710 4892
rect 2258 4850 2282 4886
rect 2318 4850 2374 4886
rect 2410 4850 2466 4886
rect 2502 4850 2558 4886
rect 2594 4850 2650 4886
rect 2686 4850 2710 4886
rect 2258 4848 2710 4850
rect 4710 4880 4908 4918
rect 4710 4848 4724 4880
rect 224 4846 4724 4848
rect 4758 4846 4796 4880
rect 4830 4846 4868 4880
rect 4902 4848 4908 4880
rect 4902 4846 5156 4848
rect -558 4842 5156 4846
rect -558 4824 816 4842
rect -558 4634 -214 4824
rect -54 4820 816 4824
rect -54 4808 286 4820
rect -54 4774 46 4808
rect 80 4774 118 4808
rect 152 4774 190 4808
rect 224 4774 286 4808
rect 852 4806 934 4842
rect 970 4806 1052 4842
rect 1088 4806 1170 4842
rect 1206 4806 1288 4842
rect 1324 4806 1406 4842
rect 1442 4806 1524 4842
rect 1560 4830 5156 4842
rect 1560 4828 3066 4830
rect 1560 4806 2992 4828
rect -54 4736 286 4774
rect -54 4702 46 4736
rect 80 4702 118 4736
rect 152 4702 190 4736
rect 224 4702 286 4736
rect -54 4664 286 4702
rect -54 4634 44 4664
rect -558 4630 44 4634
rect 78 4630 116 4664
rect 150 4630 188 4664
rect 222 4654 286 4664
rect 842 4792 2992 4806
rect 3028 4794 3066 4828
rect 3102 4794 3146 4830
rect 3182 4794 3226 4830
rect 3262 4794 3306 4830
rect 3342 4824 5156 4830
rect 3342 4808 4976 4824
rect 3342 4794 4724 4808
rect 3028 4792 4724 4794
rect 842 4774 4724 4792
rect 4758 4774 4796 4808
rect 4830 4774 4868 4808
rect 4902 4774 4976 4808
rect 842 4736 4976 4774
rect 842 4702 4724 4736
rect 4758 4702 4796 4736
rect 4830 4702 4868 4736
rect 4902 4702 4976 4736
rect 842 4664 4976 4702
rect 842 4654 4724 4664
rect 222 4630 4724 4654
rect 4758 4630 4796 4664
rect 4830 4630 4868 4664
rect 4902 4634 4976 4664
rect 5136 4634 5156 4824
rect 4902 4630 5156 4634
rect -558 4616 5156 4630
rect 28 4564 906 4584
rect 28 4134 48 4564
rect 206 4364 286 4564
rect 486 4364 686 4564
rect 886 4364 906 4564
rect 206 4344 906 4364
rect 1386 4564 3486 4584
rect 1386 4364 1406 4564
rect 1606 4364 1626 4564
rect 1826 4364 2346 4564
rect 2526 4364 3046 4564
rect 3246 4364 3266 4564
rect 3466 4364 3486 4564
rect 1386 4344 3486 4364
rect 3966 4564 4606 4584
rect 3966 4364 3986 4564
rect 4186 4364 4386 4564
rect 4586 4364 4606 4564
rect 3966 4344 4606 4364
rect 206 4314 726 4344
rect 206 4304 2346 4314
rect 206 4244 606 4304
rect 206 4134 286 4244
rect 28 4114 286 4134
rect 266 4044 286 4114
rect 486 4204 606 4244
rect 726 4204 766 4304
rect 886 4204 926 4304
rect 1046 4204 1086 4304
rect 1206 4284 2346 4304
rect 1206 4204 1226 4284
rect 2376 4254 2496 4344
rect 4146 4314 4606 4344
rect 2526 4304 4606 4314
rect 2526 4284 3666 4304
rect 1256 4224 3616 4254
rect 486 4194 1226 4204
rect 486 4044 506 4194
rect 596 4184 2346 4194
rect 30 4014 206 4034
rect 266 4014 506 4044
rect 30 3574 56 4014
rect 186 3574 206 4014
rect 266 3964 596 3984
rect 266 3954 526 3964
rect 266 3844 286 3954
rect 486 3914 526 3954
rect 576 3914 596 3964
rect 626 3914 656 4184
rect 486 3874 596 3914
rect 486 3844 526 3874
rect 266 3824 526 3844
rect 576 3854 596 3874
rect 686 3854 716 4154
rect 746 3914 776 4184
rect 806 3854 836 4154
rect 866 3914 896 4184
rect 926 3854 956 4154
rect 986 3914 1016 4184
rect 1106 4164 2346 4184
rect 1046 3854 1076 4154
rect 1106 4074 1226 4164
rect 2376 4134 2496 4224
rect 3646 4204 3666 4284
rect 3786 4204 3826 4304
rect 3946 4204 3986 4304
rect 4106 4204 4146 4304
rect 4266 4244 4606 4304
rect 4266 4204 4386 4244
rect 3646 4194 4386 4204
rect 2526 4184 4276 4194
rect 2526 4164 3766 4184
rect 1256 4104 3616 4134
rect 1106 4044 2346 4074
rect 1106 3954 1226 4044
rect 2376 4014 2496 4104
rect 3646 4074 3766 4164
rect 2526 4044 3766 4074
rect 1256 3984 3616 4014
rect 1106 3924 2346 3954
rect 1106 3884 1226 3924
rect 2376 3894 2496 3984
rect 3646 3954 3766 4044
rect 2526 3924 3766 3954
rect 1256 3864 3616 3894
rect 3646 3884 3766 3924
rect 576 3834 1076 3854
rect 2376 3834 2496 3864
rect 3796 3854 3826 4154
rect 3856 3914 3886 4184
rect 3916 3854 3946 4154
rect 3976 3914 4006 4184
rect 4036 3854 4066 4154
rect 4096 3914 4126 4184
rect 4156 3854 4186 4154
rect 4216 3914 4246 4184
rect 4366 4044 4386 4194
rect 4586 4044 4606 4244
rect 4366 4014 4606 4044
rect 4276 3954 4606 3974
rect 4276 3904 4296 3954
rect 4346 3904 4386 3954
rect 4276 3864 4386 3904
rect 4276 3854 4296 3864
rect 3796 3834 4296 3854
rect 576 3824 4296 3834
rect 266 3814 4296 3824
rect 4346 3844 4386 3864
rect 4586 3844 4606 3954
rect 4346 3814 4606 3844
rect 266 3774 4606 3814
rect 266 3744 526 3774
rect 266 3634 286 3744
rect 486 3724 526 3744
rect 576 3764 4606 3774
rect 576 3724 4296 3764
rect 486 3714 4296 3724
rect 4346 3744 4606 3764
rect 4346 3714 4386 3744
rect 486 3694 4386 3714
rect 486 3684 596 3694
rect 486 3634 526 3684
rect 576 3634 596 3684
rect 266 3614 596 3634
rect 30 3554 206 3574
rect 266 3544 506 3574
rect 266 3474 286 3544
rect 30 3444 286 3474
rect 30 3034 56 3444
rect 216 3344 286 3444
rect 486 3394 506 3544
rect 626 3404 656 3664
rect 686 3434 716 3694
rect 746 3404 776 3664
rect 806 3434 836 3694
rect 866 3404 896 3664
rect 926 3434 956 3694
rect 986 3404 1016 3664
rect 1046 3434 1076 3694
rect 1106 3634 2346 3664
rect 1106 3544 1226 3634
rect 2376 3604 2496 3694
rect 2526 3634 3766 3664
rect 1256 3574 3616 3604
rect 1106 3514 2346 3544
rect 1106 3424 1226 3514
rect 2376 3484 2496 3574
rect 3646 3544 3766 3634
rect 2526 3514 3766 3544
rect 1256 3454 3616 3484
rect 1106 3404 2346 3424
rect 596 3394 2346 3404
rect 486 3384 1226 3394
rect 486 3344 606 3384
rect 216 3284 606 3344
rect 726 3284 766 3384
rect 886 3284 926 3384
rect 1046 3284 1086 3384
rect 1206 3304 1226 3384
rect 2376 3364 2496 3454
rect 3646 3424 3766 3514
rect 3796 3434 3826 3694
rect 2526 3404 3766 3424
rect 3856 3404 3886 3664
rect 3916 3434 3946 3694
rect 3976 3404 4006 3664
rect 4036 3434 4066 3694
rect 4096 3404 4126 3664
rect 4156 3434 4186 3694
rect 4276 3674 4386 3694
rect 4216 3404 4246 3664
rect 4276 3624 4296 3674
rect 4346 3634 4386 3674
rect 4586 3634 4606 3744
rect 4346 3624 4606 3634
rect 4276 3604 4606 3624
rect 4366 3544 4606 3574
rect 2526 3394 4276 3404
rect 4366 3394 4386 3544
rect 3646 3384 4386 3394
rect 1256 3334 3616 3364
rect 1206 3284 2346 3304
rect 216 3274 2346 3284
rect 216 3244 726 3274
rect 2376 3244 2496 3334
rect 3646 3304 3666 3384
rect 2526 3284 3666 3304
rect 3786 3284 3826 3384
rect 3946 3284 3986 3384
rect 4106 3284 4146 3384
rect 4266 3344 4386 3384
rect 4586 3344 4606 3544
rect 4266 3284 4606 3344
rect 2526 3274 4606 3284
rect 4146 3244 4606 3274
rect 216 3224 906 3244
rect 216 3034 286 3224
rect 30 3024 286 3034
rect 486 3024 686 3224
rect 886 3024 906 3224
rect 30 3004 906 3024
rect 1386 3224 3486 3244
rect 1386 3024 1406 3224
rect 1606 3024 1626 3224
rect 1826 3024 2346 3224
rect 2526 3024 3046 3224
rect 3246 3024 3266 3224
rect 3466 3024 3486 3224
rect 1386 3004 3486 3024
rect 3966 3224 4606 3244
rect 3966 3024 3986 3224
rect 4186 3024 4386 3224
rect 4586 3024 4606 3224
rect 3966 3004 4606 3024
<< via1 >>
rect 66 7744 196 8144
rect 286 7954 486 8154
rect 686 7954 886 8154
rect 1406 7954 1606 8154
rect 1626 7954 1826 8154
rect 2346 7954 2526 8154
rect 3046 7954 3246 8154
rect 3266 7954 3466 8154
rect 3986 7954 4186 8154
rect 4386 7954 4586 8154
rect 286 7634 486 7834
rect 50 7164 186 7604
rect 286 7434 486 7544
rect 4386 7634 4586 7834
rect 4386 7434 4586 7544
rect 286 7224 486 7334
rect 286 6934 486 7134
rect 4386 7224 4586 7334
rect 4386 6934 4586 7134
rect 286 6614 486 6814
rect 686 6614 886 6814
rect 1406 6614 1606 6814
rect 1626 6614 1826 6814
rect 2346 6614 2526 6814
rect 3046 6614 3246 6814
rect 3266 6614 3466 6814
rect 3986 6614 4186 6814
rect 4386 6614 4586 6814
rect -494 6354 -334 6544
rect 5246 6354 5406 6544
rect 1726 6074 1876 6224
rect 1826 4994 1976 5144
rect -214 4634 -54 4824
rect 286 4806 816 4820
rect 816 4806 842 4820
rect 286 4654 842 4806
rect 4976 4634 5136 4824
rect 286 4364 486 4564
rect 686 4364 886 4564
rect 1406 4364 1606 4564
rect 1626 4364 1826 4564
rect 2346 4364 2526 4564
rect 3046 4364 3246 4564
rect 3266 4364 3466 4564
rect 3986 4364 4186 4564
rect 4386 4364 4586 4564
rect 286 4044 486 4244
rect 56 3574 186 4014
rect 286 3844 486 3954
rect 4386 4044 4586 4244
rect 4386 3844 4586 3954
rect 286 3634 486 3744
rect 56 3034 216 3444
rect 286 3344 486 3544
rect 4386 3634 4586 3744
rect 4386 3344 4586 3544
rect 286 3024 486 3224
rect 686 3024 886 3224
rect 1406 3024 1606 3224
rect 1626 3024 1826 3224
rect 2346 3024 2526 3224
rect 3046 3024 3246 3224
rect 3266 3024 3466 3224
rect 3986 3024 4186 3224
rect 4386 3024 4586 3224
<< metal2 >>
rect 30 8154 906 8174
rect 30 8144 286 8154
rect 30 7744 66 8144
rect 196 7954 286 8144
rect 486 7954 686 8154
rect 886 7954 906 8154
rect 196 7934 906 7954
rect 1386 8154 3486 8174
rect 1386 7954 1406 8154
rect 1606 7954 1626 8154
rect 1826 7954 2346 8154
rect 2526 7954 3046 8154
rect 3246 7954 3266 8154
rect 3466 7954 3486 8154
rect 196 7834 656 7934
rect 1386 7894 3486 7954
rect 3966 8154 4606 8174
rect 3966 7954 3986 8154
rect 4186 7954 4386 8154
rect 4586 7954 4606 8154
rect 3966 7934 4606 7954
rect 196 7744 286 7834
rect 30 7704 286 7744
rect 266 7634 286 7704
rect 486 7744 656 7834
rect 686 7774 4186 7894
rect 4216 7834 4606 7934
rect 486 7714 1056 7744
rect 486 7634 656 7714
rect 1086 7684 1146 7774
rect 686 7654 1146 7684
rect 266 7624 656 7634
rect 30 7604 206 7624
rect 266 7604 1056 7624
rect 30 7164 50 7604
rect 186 7164 206 7604
rect 546 7594 1056 7604
rect 266 7544 506 7564
rect 266 7434 286 7544
rect 486 7434 506 7544
rect 266 7334 506 7434
rect 266 7224 286 7334
rect 486 7224 506 7334
rect 266 7204 506 7224
rect 546 7474 656 7594
rect 1086 7564 1146 7654
rect 686 7534 1146 7564
rect 546 7414 1056 7474
rect 1086 7444 1146 7534
rect 1176 7414 1206 7744
rect 1236 7444 1266 7774
rect 1296 7414 1326 7744
rect 1356 7444 1386 7774
rect 1416 7414 1446 7744
rect 1476 7444 1506 7774
rect 1536 7414 1566 7744
rect 1596 7444 1626 7774
rect 1656 7414 1686 7744
rect 1716 7444 1746 7774
rect 1776 7414 1806 7744
rect 1836 7444 1866 7774
rect 1896 7414 1926 7744
rect 1956 7444 1986 7774
rect 2016 7414 2046 7744
rect 2076 7444 2106 7774
rect 2136 7414 2166 7744
rect 2196 7444 2226 7774
rect 2256 7414 2286 7744
rect 2316 7444 2346 7774
rect 2376 7414 2496 7744
rect 2526 7444 2556 7774
rect 2586 7414 2616 7744
rect 2646 7444 2676 7774
rect 2706 7414 2736 7744
rect 2766 7444 2796 7774
rect 2826 7414 2856 7744
rect 2886 7444 2916 7774
rect 2946 7414 2976 7744
rect 3006 7444 3036 7774
rect 3066 7414 3096 7744
rect 3126 7444 3156 7774
rect 3186 7414 3216 7744
rect 3246 7444 3276 7774
rect 3306 7414 3336 7744
rect 3366 7444 3396 7774
rect 3426 7414 3456 7744
rect 3486 7444 3516 7774
rect 3546 7414 3576 7744
rect 3606 7444 3636 7774
rect 3666 7414 3696 7744
rect 3726 7684 3786 7774
rect 4216 7744 4386 7834
rect 3816 7714 4386 7744
rect 3726 7654 4186 7684
rect 3726 7564 3786 7654
rect 4216 7634 4386 7714
rect 4586 7634 4606 7834
rect 4216 7624 4606 7634
rect 3816 7604 4606 7624
rect 3816 7594 4326 7604
rect 3726 7534 4186 7564
rect 3726 7444 3786 7534
rect 4216 7474 4326 7594
rect 3816 7414 4326 7474
rect 546 7354 4326 7414
rect 546 7264 1056 7354
rect 546 7174 656 7264
rect 1086 7234 1146 7324
rect 686 7204 1146 7234
rect 546 7164 1056 7174
rect 30 7144 206 7164
rect 266 7144 1056 7164
rect 266 7134 656 7144
rect 266 6934 286 7134
rect 486 7054 656 7134
rect 1086 7114 1146 7204
rect 686 7084 1146 7114
rect 486 7024 1056 7054
rect 486 6934 656 7024
rect 1086 6994 1146 7084
rect 1176 7024 1206 7354
rect 1236 6994 1266 7324
rect 1296 7024 1326 7354
rect 1356 6994 1386 7324
rect 1416 7024 1446 7354
rect 1476 6994 1506 7324
rect 1536 7024 1566 7354
rect 1596 6994 1626 7324
rect 1656 7024 1686 7354
rect 1716 6994 1746 7324
rect 1776 7024 1806 7354
rect 1836 6994 1866 7324
rect 1896 7024 1926 7354
rect 1956 6994 1986 7324
rect 2016 7024 2046 7354
rect 2076 6994 2106 7324
rect 2136 7024 2166 7354
rect 2196 6994 2226 7324
rect 2256 7024 2286 7354
rect 2316 6994 2346 7324
rect 2376 7024 2496 7354
rect 2526 6994 2556 7324
rect 2586 7024 2616 7354
rect 2646 6994 2676 7324
rect 2706 7024 2736 7354
rect 2766 6994 2796 7324
rect 2826 7024 2856 7354
rect 2886 6994 2916 7324
rect 2946 7024 2976 7354
rect 3006 6994 3036 7324
rect 3066 7024 3096 7354
rect 3126 6994 3156 7324
rect 3186 7024 3216 7354
rect 3246 6994 3276 7324
rect 3306 7024 3336 7354
rect 3366 6994 3396 7324
rect 3426 7024 3456 7354
rect 3486 6994 3516 7324
rect 3546 7024 3576 7354
rect 3606 6994 3636 7324
rect 3666 7024 3696 7354
rect 3726 7234 3786 7324
rect 3816 7264 4326 7354
rect 3726 7204 4186 7234
rect 3726 7114 3786 7204
rect 4216 7174 4326 7264
rect 4366 7544 4606 7564
rect 4366 7434 4386 7544
rect 4586 7434 4606 7544
rect 4366 7334 4606 7434
rect 4366 7224 4386 7334
rect 4586 7224 4606 7334
rect 4366 7204 4606 7224
rect 3816 7164 4326 7174
rect 3816 7144 4606 7164
rect 4216 7134 4606 7144
rect 3726 7084 4186 7114
rect 3726 6994 3786 7084
rect 4216 7054 4386 7134
rect 3816 7024 4386 7054
rect 266 6834 656 6934
rect 686 6874 4186 6994
rect 4216 6934 4386 7024
rect 4586 6934 4606 7134
rect 266 6814 906 6834
rect 266 6614 286 6814
rect 486 6614 686 6814
rect 886 6614 906 6814
rect 266 6594 906 6614
rect 1386 6814 3486 6874
rect 4216 6834 4606 6934
rect 1386 6614 1406 6814
rect 1606 6614 1626 6814
rect 1826 6614 2346 6814
rect 2526 6614 3046 6814
rect 3246 6614 3266 6814
rect 3466 6614 3486 6814
rect 1386 6594 3486 6614
rect 3966 6814 4606 6834
rect 3966 6614 3986 6814
rect 4186 6614 4386 6814
rect 4586 6614 4606 6814
rect 3966 6594 4606 6614
rect -512 6544 -312 6566
rect -512 6354 -494 6544
rect -334 6354 -312 6544
rect -512 6336 -312 6354
rect 1706 6224 1896 6594
rect 5226 6544 5426 6566
rect 5226 6354 5246 6544
rect 5406 6354 5426 6544
rect 5226 6336 5426 6354
rect 1706 6074 1726 6224
rect 1876 6074 1896 6224
rect 1706 6054 1896 6074
rect 1806 5144 1996 5164
rect 1806 4994 1826 5144
rect 1976 4994 1996 5144
rect -236 4824 -36 4848
rect -236 4634 -214 4824
rect -54 4634 -36 4824
rect 258 4820 888 4848
rect 258 4654 286 4820
rect 842 4654 888 4820
rect 258 4648 888 4654
rect -236 4616 -36 4634
rect 266 4584 896 4648
rect 1806 4584 1996 4994
rect 4956 4824 5156 4848
rect 4956 4634 4976 4824
rect 5136 4634 5156 4824
rect 4956 4616 5156 4634
rect 266 4564 906 4584
rect 266 4364 286 4564
rect 486 4364 686 4564
rect 886 4364 906 4564
rect 266 4344 906 4364
rect 1386 4564 3486 4584
rect 1386 4364 1406 4564
rect 1606 4364 1626 4564
rect 1826 4364 2346 4564
rect 2526 4364 3046 4564
rect 3246 4364 3266 4564
rect 3466 4364 3486 4564
rect 266 4244 656 4344
rect 1386 4304 3486 4364
rect 3966 4564 4606 4584
rect 3966 4364 3986 4564
rect 4186 4364 4386 4564
rect 4586 4364 4606 4564
rect 3966 4344 4606 4364
rect 266 4044 286 4244
rect 486 4154 656 4244
rect 686 4184 4186 4304
rect 4216 4244 4606 4344
rect 486 4124 1056 4154
rect 486 4044 656 4124
rect 1086 4094 1146 4184
rect 686 4064 1146 4094
rect 266 4034 656 4044
rect 30 4014 206 4034
rect 266 4014 1056 4034
rect 30 3574 56 4014
rect 186 3574 206 4014
rect 546 4004 1056 4014
rect 266 3954 506 3974
rect 266 3844 286 3954
rect 486 3844 506 3954
rect 266 3744 506 3844
rect 266 3634 286 3744
rect 486 3634 506 3744
rect 266 3614 506 3634
rect 546 3884 656 4004
rect 1086 3974 1146 4064
rect 686 3944 1146 3974
rect 546 3824 1056 3884
rect 1086 3854 1146 3944
rect 1176 3824 1206 4154
rect 1236 3854 1266 4184
rect 1296 3824 1326 4154
rect 1356 3854 1386 4184
rect 1416 3824 1446 4154
rect 1476 3854 1506 4184
rect 1536 3824 1566 4154
rect 1596 3854 1626 4184
rect 1656 3824 1686 4154
rect 1716 3854 1746 4184
rect 1776 3824 1806 4154
rect 1836 3854 1866 4184
rect 1896 3824 1926 4154
rect 1956 3854 1986 4184
rect 2016 3824 2046 4154
rect 2076 3854 2106 4184
rect 2136 3824 2166 4154
rect 2196 3854 2226 4184
rect 2256 3824 2286 4154
rect 2316 3854 2346 4184
rect 2376 3824 2496 4154
rect 2526 3854 2556 4184
rect 2586 3824 2616 4154
rect 2646 3854 2676 4184
rect 2706 3824 2736 4154
rect 2766 3854 2796 4184
rect 2826 3824 2856 4154
rect 2886 3854 2916 4184
rect 2946 3824 2976 4154
rect 3006 3854 3036 4184
rect 3066 3824 3096 4154
rect 3126 3854 3156 4184
rect 3186 3824 3216 4154
rect 3246 3854 3276 4184
rect 3306 3824 3336 4154
rect 3366 3854 3396 4184
rect 3426 3824 3456 4154
rect 3486 3854 3516 4184
rect 3546 3824 3576 4154
rect 3606 3854 3636 4184
rect 3666 3824 3696 4154
rect 3726 4094 3786 4184
rect 4216 4154 4386 4244
rect 3816 4124 4386 4154
rect 3726 4064 4186 4094
rect 3726 3974 3786 4064
rect 4216 4044 4386 4124
rect 4586 4044 4606 4244
rect 4216 4034 4606 4044
rect 3816 4014 4606 4034
rect 3816 4004 4326 4014
rect 3726 3944 4186 3974
rect 3726 3854 3786 3944
rect 4216 3884 4326 4004
rect 3816 3824 4326 3884
rect 546 3764 4326 3824
rect 546 3674 1056 3764
rect 546 3584 656 3674
rect 1086 3644 1146 3734
rect 686 3614 1146 3644
rect 546 3574 1056 3584
rect 30 3554 206 3574
rect 266 3554 1056 3574
rect 266 3544 656 3554
rect 266 3474 286 3544
rect 30 3444 286 3474
rect 30 3034 56 3444
rect 216 3344 286 3444
rect 486 3464 656 3544
rect 1086 3524 1146 3614
rect 686 3494 1146 3524
rect 486 3434 1056 3464
rect 486 3344 656 3434
rect 1086 3404 1146 3494
rect 1176 3434 1206 3764
rect 1236 3404 1266 3734
rect 1296 3434 1326 3764
rect 1356 3404 1386 3734
rect 1416 3434 1446 3764
rect 1476 3404 1506 3734
rect 1536 3434 1566 3764
rect 1596 3404 1626 3734
rect 1656 3434 1686 3764
rect 1716 3404 1746 3734
rect 1776 3434 1806 3764
rect 1836 3404 1866 3734
rect 1896 3434 1926 3764
rect 1956 3404 1986 3734
rect 2016 3434 2046 3764
rect 2076 3404 2106 3734
rect 2136 3434 2166 3764
rect 2196 3404 2226 3734
rect 2256 3434 2286 3764
rect 2316 3404 2346 3734
rect 2376 3434 2496 3764
rect 2526 3404 2556 3734
rect 2586 3434 2616 3764
rect 2646 3404 2676 3734
rect 2706 3434 2736 3764
rect 2766 3404 2796 3734
rect 2826 3434 2856 3764
rect 2886 3404 2916 3734
rect 2946 3434 2976 3764
rect 3006 3404 3036 3734
rect 3066 3434 3096 3764
rect 3126 3404 3156 3734
rect 3186 3434 3216 3764
rect 3246 3404 3276 3734
rect 3306 3434 3336 3764
rect 3366 3404 3396 3734
rect 3426 3434 3456 3764
rect 3486 3404 3516 3734
rect 3546 3434 3576 3764
rect 3606 3404 3636 3734
rect 3666 3434 3696 3764
rect 3726 3644 3786 3734
rect 3816 3674 4326 3764
rect 3726 3614 4186 3644
rect 3726 3524 3786 3614
rect 4216 3584 4326 3674
rect 4366 3954 4606 3974
rect 4366 3844 4386 3954
rect 4586 3844 4606 3954
rect 4366 3744 4606 3844
rect 4366 3634 4386 3744
rect 4586 3634 4606 3744
rect 4366 3614 4606 3634
rect 3816 3574 4326 3584
rect 3816 3554 4606 3574
rect 4216 3544 4606 3554
rect 3726 3494 4186 3524
rect 3726 3404 3786 3494
rect 4216 3464 4386 3544
rect 3816 3434 4386 3464
rect 216 3244 656 3344
rect 686 3284 4186 3404
rect 4216 3344 4386 3434
rect 4586 3344 4606 3544
rect 216 3224 906 3244
rect 216 3034 286 3224
rect 30 3024 286 3034
rect 486 3024 686 3224
rect 886 3024 906 3224
rect 30 3004 906 3024
rect 1386 3224 3486 3284
rect 4216 3244 4606 3344
rect 1386 3024 1406 3224
rect 1606 3024 1626 3224
rect 1826 3024 2346 3224
rect 2526 3024 3046 3224
rect 3246 3024 3266 3224
rect 3466 3024 3486 3224
rect 1386 3004 3486 3024
rect 3966 3224 4606 3244
rect 3966 3024 3986 3224
rect 4186 3024 4386 3224
rect 4586 3024 4606 3224
rect 3966 3004 4606 3024
<< via2 >>
rect 66 7744 196 8144
rect 50 7164 186 7604
rect -494 6354 -334 6544
rect 5246 6354 5406 6544
rect -214 4634 -54 4824
rect 286 4654 842 4820
rect 4976 4634 5136 4824
rect 56 3574 186 4014
rect 56 3034 216 3444
<< metal3 >>
rect 30 8154 906 8174
rect 30 8144 286 8154
rect 30 7744 66 8144
rect 196 7984 286 8144
rect 456 7984 706 8154
rect 876 7984 906 8154
rect 1386 8154 3486 8174
rect 1386 8024 1406 8154
rect 1536 8024 1566 8154
rect 1696 8024 3176 8154
rect 3306 8024 3336 8154
rect 3466 8024 3486 8154
rect 1386 8004 3486 8024
rect 3966 8154 4606 8174
rect 196 7924 906 7984
rect 3966 7984 3996 8154
rect 4166 7984 4416 8154
rect 4586 7984 4606 8154
rect 3966 7924 4606 7984
rect 196 7894 4606 7924
rect 196 7744 286 7894
rect 30 7724 286 7744
rect 456 7724 4416 7894
rect 4586 7724 4606 7894
rect 30 7704 4606 7724
rect 266 7694 4606 7704
rect 30 7604 206 7624
rect 30 7164 50 7604
rect 186 7164 206 7604
rect 30 7144 206 7164
rect 266 7604 436 7624
rect 266 7404 286 7604
rect 416 7404 436 7604
rect 266 7364 436 7404
rect 266 7164 286 7364
rect 416 7164 436 7364
rect 266 7144 436 7164
rect 516 7074 4356 7694
rect 4436 7604 4606 7624
rect 4436 7404 4456 7604
rect 4586 7404 4606 7604
rect 4436 7364 4606 7404
rect 4436 7164 4456 7364
rect 4586 7164 4606 7364
rect 4436 7144 4606 7164
rect 266 7044 4606 7074
rect 266 6874 286 7044
rect 456 6874 4416 7044
rect 4586 6874 4606 7044
rect 266 6844 4606 6874
rect 266 6784 906 6844
rect 266 6614 286 6784
rect 456 6614 706 6784
rect 876 6614 906 6784
rect 3966 6784 4606 6844
rect 266 6594 906 6614
rect 1386 6744 3486 6764
rect 1386 6614 1406 6744
rect 1536 6614 1566 6744
rect 1696 6614 3176 6744
rect 3306 6614 3336 6744
rect 3466 6614 3486 6744
rect 1386 6594 3486 6614
rect 3966 6614 3996 6784
rect 4166 6614 4416 6784
rect 4586 6614 4606 6784
rect 3966 6594 4606 6614
rect -512 6544 -312 6566
rect -512 6354 -494 6544
rect -334 6354 -312 6544
rect -512 6336 -312 6354
rect 5226 6544 5426 6566
rect 5226 6354 5246 6544
rect 5406 6354 5426 6544
rect 5226 6336 5426 6354
rect -236 4824 -36 4848
rect -236 4634 -214 4824
rect -54 4634 -36 4824
rect 258 4820 888 4848
rect 258 4654 286 4820
rect 842 4654 888 4820
rect 258 4648 888 4654
rect 4956 4824 5156 4848
rect -236 4616 -36 4634
rect 4956 4634 4976 4824
rect 5136 4634 5156 4824
rect 4956 4616 5156 4634
rect 266 4564 906 4584
rect 266 4394 286 4564
rect 456 4394 706 4564
rect 876 4394 906 4564
rect 1386 4564 3486 4584
rect 1386 4434 1406 4564
rect 1536 4434 1566 4564
rect 1696 4434 3176 4564
rect 3306 4434 3336 4564
rect 3466 4434 3486 4564
rect 1386 4414 3486 4434
rect 3966 4564 4606 4584
rect 266 4334 906 4394
rect 3966 4394 3996 4564
rect 4166 4394 4416 4564
rect 4586 4394 4606 4564
rect 3966 4334 4606 4394
rect 266 4304 4606 4334
rect 266 4134 286 4304
rect 456 4134 4416 4304
rect 4586 4134 4606 4304
rect 266 4104 4606 4134
rect 30 4014 206 4034
rect 30 3574 56 4014
rect 186 3574 206 4014
rect 30 3554 206 3574
rect 266 4014 436 4034
rect 266 3814 286 4014
rect 416 3814 436 4014
rect 266 3774 436 3814
rect 266 3574 286 3774
rect 416 3574 436 3774
rect 266 3554 436 3574
rect 516 3484 4356 4104
rect 4436 4014 4606 4034
rect 4436 3814 4456 4014
rect 4586 3814 4606 4014
rect 4436 3774 4606 3814
rect 4436 3574 4456 3774
rect 4586 3574 4606 3774
rect 4436 3554 4606 3574
rect 266 3474 4606 3484
rect 30 3454 4606 3474
rect 30 3444 286 3454
rect 30 3034 56 3444
rect 216 3284 286 3444
rect 456 3284 4416 3454
rect 4586 3284 4606 3454
rect 216 3254 4606 3284
rect 216 3194 906 3254
rect 216 3034 286 3194
rect 30 3024 286 3034
rect 456 3024 706 3194
rect 876 3024 906 3194
rect 3966 3194 4606 3254
rect 30 3004 906 3024
rect 1386 3154 3486 3174
rect 1386 3024 1406 3154
rect 1536 3024 1566 3154
rect 1696 3024 3176 3154
rect 3306 3024 3336 3154
rect 3466 3024 3486 3154
rect 1386 3004 3486 3024
rect 3966 3024 3996 3194
rect 4166 3024 4416 3194
rect 4586 3024 4606 3194
rect 3966 3004 4606 3024
<< via3 >>
rect 66 7744 196 8144
rect 286 7984 456 8154
rect 706 7984 876 8154
rect 1406 8024 1536 8154
rect 1566 8024 1696 8154
rect 3176 8024 3306 8154
rect 3336 8024 3466 8154
rect 3996 7984 4166 8154
rect 4416 7984 4586 8154
rect 286 7724 456 7894
rect 4416 7724 4586 7894
rect 50 7164 186 7604
rect 286 7404 416 7604
rect 286 7164 416 7364
rect 4456 7404 4586 7604
rect 4456 7164 4586 7364
rect 286 6874 456 7044
rect 4416 6874 4586 7044
rect 286 6614 456 6784
rect 706 6614 876 6784
rect 1406 6614 1536 6744
rect 1566 6614 1696 6744
rect 3176 6614 3306 6744
rect 3336 6614 3466 6744
rect 3996 6614 4166 6784
rect 4416 6614 4586 6784
rect -494 6354 -334 6544
rect 5246 6354 5406 6544
rect -214 4634 -54 4824
rect 4976 4634 5136 4824
rect 286 4394 456 4564
rect 706 4394 876 4564
rect 1406 4434 1536 4564
rect 1566 4434 1696 4564
rect 3176 4434 3306 4564
rect 3336 4434 3466 4564
rect 3996 4394 4166 4564
rect 4416 4394 4586 4564
rect 286 4134 456 4304
rect 4416 4134 4586 4304
rect 56 3574 186 4014
rect 286 3814 416 4014
rect 286 3574 416 3774
rect 4456 3814 4586 4014
rect 4456 3574 4586 3774
rect 56 3034 216 3444
rect 286 3284 456 3454
rect 4416 3284 4586 3454
rect 286 3024 456 3194
rect 706 3024 876 3194
rect 1406 3024 1536 3154
rect 1566 3024 1696 3154
rect 3176 3024 3306 3154
rect 3336 3024 3466 3154
rect 3996 3024 4166 3194
rect 4416 3024 4586 3194
<< mimcap >>
rect 546 7864 4326 7894
rect 546 6904 576 7864
rect 4296 6904 4326 7864
rect 546 6874 4326 6904
rect 546 4274 4326 4304
rect 546 3314 576 4274
rect 4296 3314 4326 4274
rect 546 3284 4326 3314
<< mimcapcontact >>
rect 576 6904 4296 7864
rect 576 3314 4296 4274
<< metal4 >>
rect -512 6544 -312 8392
rect -512 6354 -494 6544
rect -334 6354 -312 6544
rect -512 2796 -312 6354
rect -236 4824 -36 8392
rect 30 8154 896 8174
rect 30 8144 286 8154
rect 30 7744 66 8144
rect 196 7984 286 8144
rect 456 7984 706 8154
rect 876 7984 896 8154
rect 196 7964 896 7984
rect 1386 8154 3486 8174
rect 1386 8024 1406 8154
rect 1536 8024 1566 8154
rect 1696 8024 3176 8154
rect 3306 8024 3336 8154
rect 3466 8024 3486 8154
rect 196 7894 476 7964
rect 196 7744 286 7894
rect 30 7724 286 7744
rect 456 7724 476 7894
rect 1386 7884 3486 8024
rect 3976 8154 4606 8174
rect 3976 7984 3996 8154
rect 4166 7984 4416 8154
rect 4586 7984 4606 8154
rect 3976 7964 4606 7984
rect 4396 7894 4606 7964
rect 30 7704 476 7724
rect 556 7864 4316 7884
rect 556 7624 576 7864
rect 30 7604 576 7624
rect 30 7164 50 7604
rect 186 7404 286 7604
rect 416 7404 576 7604
rect 186 7364 576 7404
rect 186 7164 286 7364
rect 416 7164 576 7364
rect 30 7144 576 7164
rect 266 7044 476 7064
rect 266 6874 286 7044
rect 456 6874 476 7044
rect 556 6904 576 7144
rect 4296 7624 4316 7864
rect 4396 7724 4416 7894
rect 4586 7724 4606 7894
rect 4396 7704 4606 7724
rect 4296 7604 4606 7624
rect 4296 7404 4456 7604
rect 4586 7404 4606 7604
rect 4296 7364 4606 7404
rect 4296 7164 4456 7364
rect 4586 7164 4606 7364
rect 4296 7144 4606 7164
rect 4296 6904 4316 7144
rect 556 6884 4316 6904
rect 4396 7044 4606 7064
rect 266 6804 476 6874
rect 266 6784 896 6804
rect 266 6614 286 6784
rect 456 6614 706 6784
rect 876 6614 896 6784
rect 266 6594 896 6614
rect 1386 6744 3486 6884
rect 4396 6874 4416 7044
rect 4586 6874 4606 7044
rect 4396 6804 4606 6874
rect 1386 6614 1406 6744
rect 1536 6614 1566 6744
rect 1696 6614 3176 6744
rect 3306 6614 3336 6744
rect 3466 6614 3486 6744
rect 1386 6594 3486 6614
rect 3976 6784 4606 6804
rect 3976 6614 3996 6784
rect 4166 6614 4416 6784
rect 4586 6614 4606 6784
rect 3976 6594 4606 6614
rect -236 4634 -214 4824
rect -54 4634 -36 4824
rect -236 2796 -36 4634
rect 4956 4824 5156 8392
rect 4956 4634 4976 4824
rect 5136 4634 5156 4824
rect 266 4564 896 4584
rect 266 4394 286 4564
rect 456 4394 706 4564
rect 876 4394 896 4564
rect 266 4374 896 4394
rect 1386 4564 3486 4584
rect 1386 4434 1406 4564
rect 1536 4434 1566 4564
rect 1696 4434 3176 4564
rect 3306 4434 3336 4564
rect 3466 4434 3486 4564
rect 266 4304 476 4374
rect 266 4134 286 4304
rect 456 4134 476 4304
rect 1386 4294 3486 4434
rect 3976 4564 4606 4584
rect 3976 4394 3996 4564
rect 4166 4394 4416 4564
rect 4586 4394 4606 4564
rect 3976 4374 4606 4394
rect 4396 4304 4606 4374
rect 266 4114 476 4134
rect 556 4274 4316 4294
rect 556 4034 576 4274
rect 30 4014 576 4034
rect 30 3574 56 4014
rect 186 3814 286 4014
rect 416 3814 576 4014
rect 186 3774 576 3814
rect 186 3574 286 3774
rect 416 3574 576 3774
rect 30 3554 576 3574
rect 30 3454 476 3474
rect 30 3444 286 3454
rect 30 3034 56 3444
rect 216 3284 286 3444
rect 456 3284 476 3454
rect 556 3314 576 3554
rect 4296 4034 4316 4274
rect 4396 4134 4416 4304
rect 4586 4134 4606 4304
rect 4396 4114 4606 4134
rect 4296 4014 4606 4034
rect 4296 3814 4456 4014
rect 4586 3814 4606 4014
rect 4296 3774 4606 3814
rect 4296 3574 4456 3774
rect 4586 3574 4606 3774
rect 4296 3554 4606 3574
rect 4296 3314 4316 3554
rect 556 3294 4316 3314
rect 4396 3454 4606 3474
rect 216 3214 476 3284
rect 216 3194 896 3214
rect 216 3034 286 3194
rect 30 3024 286 3034
rect 456 3024 706 3194
rect 876 3024 896 3194
rect 30 3004 896 3024
rect 1386 3154 3486 3294
rect 4396 3284 4416 3454
rect 4586 3284 4606 3454
rect 4396 3214 4606 3284
rect 1386 3024 1406 3154
rect 1536 3024 1566 3154
rect 1696 3024 3176 3154
rect 3306 3024 3336 3154
rect 3466 3024 3486 3154
rect 1386 3004 3486 3024
rect 3976 3194 4606 3214
rect 3976 3024 3996 3194
rect 4166 3024 4416 3194
rect 4586 3024 4606 3194
rect 3976 3004 4606 3024
rect 4956 2796 5156 4634
rect 5226 6544 5426 8392
rect 5226 6354 5246 6544
rect 5406 6354 5426 6544
rect 5226 2796 5426 6354
<< comment >>
rect 810 6116 842 6158
rect 1006 6112 1038 6154
rect 1196 6110 1228 6152
rect 1388 6110 1420 6152
rect 1580 6112 1612 6154
rect 2048 5824 2066 6028
rect 2270 5836 2290 6056
rect 2464 5808 2484 6028
rect 2658 5866 2678 6086
rect 3820 6060 3840 6208
rect 3928 6060 3966 6196
rect 4054 6054 4074 6202
rect 4316 6060 4336 6208
rect 4424 6060 4462 6196
rect 4550 6054 4570 6202
rect 3298 6036 3332 6050
rect 3490 6038 3524 6052
rect 2884 5824 2902 6028
rect 3298 5840 3332 5852
rect 3490 5840 3524 5852
rect 3836 5814 3864 5862
rect 4332 5814 4360 5862
rect 816 5422 848 5464
rect 1004 5436 1036 5478
rect 1192 5438 1224 5480
rect 1396 5442 1428 5484
rect 1584 5450 1616 5492
rect 3298 5400 3332 5412
rect 3490 5400 3524 5412
rect 3996 5394 4024 5442
rect 2264 5118 2292 5286
rect 2458 5116 2486 5284
rect 2650 5102 2678 5270
rect 3298 5202 3332 5216
rect 3490 5200 3524 5214
rect 908 5034 940 5076
rect 1106 5032 1138 5074
rect 1294 5034 1326 5076
rect 1482 5034 1514 5076
rect 3980 5048 4000 5196
rect 4088 5060 4126 5196
rect 4214 5054 4234 5202
<< labels >>
flabel metal1 s -558 5174 -544 5202 7 FreeSans 160 0 0 0 clk
port 32 w
flabel metal1 s -558 5822 -544 5850 7 FreeSans 160 0 0 0 inn
port 30 w
flabel metal1 s -558 5878 -544 5906 7 FreeSans 160 0 0 0 inp
port 31 w
flabel metal1 s -558 6336 -530 6566 7 FreeSans 160 0 0 0 VDD
port 27 w
flabel metal1 s -558 4616 -536 4848 7 FreeSans 160 0 0 0 VSS
port 26 w
flabel metal1 s 5290 5972 5452 6000 3 FreeSans 160 0 0 0 latch_q
port 21 e
flabel metal1 s 5290 5904 5452 5932 3 FreeSans 160 0 0 0 latch_qn
port 22 e
flabel metal1 s 5290 5314 5452 5342 3 FreeSans 160 0 0 0 comp_trig
port 23 e
rlabel locali 496 5164 496 5210 7 inverter_1/in
rlabel locali 730 5164 730 5210 3 inverter_1/out
rlabel metal1 578 4902 578 4948 7 inverter_1/VSS
rlabel metal1 576 5568 576 5614 7 inverter_1/VDD
rlabel locali 262 5164 262 5210 7 inverter_0/in
rlabel locali 496 5164 496 5210 3 inverter_0/out
rlabel metal1 344 4902 344 4948 7 inverter_0/VSS
rlabel metal1 342 5568 342 5614 7 inverter_0/VDD
rlabel locali 1926 5572 1926 5606 7 adc_comp_circuit_0/bn
rlabel locali 3016 5572 3016 5606 3 adc_comp_circuit_0/bp
rlabel locali 3578 5312 3578 5350 3 adc_comp_circuit_0/outn
rlabel locali 3576 5902 3576 5940 3 adc_comp_circuit_0/outp
rlabel locali 1290 5724 1290 5756 7 adc_comp_circuit_0/on
rlabel locali 906 5724 906 5756 7 adc_comp_circuit_0/op
rlabel locali 2156 4876 2156 4930 7 adc_comp_circuit_0/nclk
rlabel locali 710 5130 710 5160 7 adc_comp_circuit_0/clk
flabel metal4 4956 2796 5156 8392 0 FreeSans 800 90 0 0 adc_comp_circuit_0/VSS
flabel metal4 5226 2796 5426 8392 0 FreeSans 800 90 0 0 adc_comp_circuit_0/VDD
flabel metal4 -236 2796 -36 8392 0 FreeSans 800 90 0 0 adc_comp_circuit_0/VSS
flabel metal4 -512 2796 -312 8392 0 FreeSans 800 90 0 0 adc_comp_circuit_0/VDD
rlabel metal1 -558 5878 -558 5906 7 adc_comp_circuit_0/inp
rlabel metal1 -558 5822 -558 5850 7 adc_comp_circuit_0/inn
rlabel metal1 -558 4690 -558 4848 7 adc_comp_circuit_0/VSS
rlabel metal1 -558 6336 -558 6474 7 adc_comp_circuit_0/VDD
flabel metal1 266 6594 906 6834 5 FreeSans 320 0 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_1/nmoscap_bot
flabel metal1 266 7934 906 8174 1 FreeSans 320 0 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_1/nmoscap_bot
flabel metal1 3966 6594 4606 6834 5 FreeSans 320 0 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_1/nmoscap_bot
flabel metal1 3966 7934 4606 8174 1 FreeSans 320 0 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_1/nmoscap_bot
flabel metal1 266 7604 506 8174 7 FreeSans 160 90 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_1/nmoscap_bot
flabel metal1 266 6594 506 7164 7 FreeSans 160 90 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_1/nmoscap_bot
flabel metal1 4366 6594 4606 7164 3 FreeSans 160 90 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_1/nmoscap_bot
flabel metal1 4366 7604 4606 8174 3 FreeSans 160 90 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_1/nmoscap_bot
flabel metal1 1386 6594 3486 6834 5 FreeSans 320 0 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_1/nmoscap_top
flabel metal1 1386 7934 3486 8174 1 FreeSans 320 0 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_1/nmoscap_top
flabel metal1 266 7204 506 7574 7 FreeSans 320 90 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_1/nmoscap_top
flabel metal1 4366 7194 4606 7564 3 FreeSans 320 90 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_1/nmoscap_top
flabel locali 916 6594 1376 6674 5 FreeSans 320 0 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_1/pwell
flabel locali 3496 6594 3956 6674 5 FreeSans 320 0 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_1/pwell
flabel locali 916 8094 1376 8174 1 FreeSans 320 0 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_1/pwell
flabel locali 3496 8094 3956 8174 1 FreeSans 320 0 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_1/pwell
flabel metal3 266 6594 906 6834 5 FreeSans 320 0 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_1/mimcap_bot
flabel metal3 3966 6594 4606 6834 5 FreeSans 320 0 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_1/mimcap_bot
flabel metal3 266 7934 906 8174 1 FreeSans 320 0 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_1/mimcap_bot
flabel metal3 3966 7934 4606 8174 1 FreeSans 320 0 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_1/mimcap_bot
flabel metal3 266 7694 516 8174 7 FreeSans 320 90 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_1/mimcap_bot
flabel metal3 266 6594 516 7074 7 FreeSans 320 90 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_1/mimcap_bot
flabel metal3 4356 6594 4606 7074 3 FreeSans 320 90 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_1/mimcap_bot
flabel metal3 4356 7694 4606 8174 3 FreeSans 320 90 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_1/mimcap_bot
flabel metal3 1386 6594 3486 6764 5 FreeSans 320 0 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_1/mimcap_top
flabel metal3 1386 8004 3486 8174 1 FreeSans 320 0 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_1/mimcap_top
flabel metal3 4436 7144 4606 7624 3 FreeSans 320 90 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_1/mimcap_top
flabel metal3 266 7144 436 7624 7 FreeSans 320 90 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_1/mimcap_top
flabel metal1 266 3004 906 3244 5 FreeSans 320 0 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_0/nmoscap_bot
flabel metal1 266 4344 906 4584 1 FreeSans 320 0 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_0/nmoscap_bot
flabel metal1 3966 3004 4606 3244 5 FreeSans 320 0 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_0/nmoscap_bot
flabel metal1 3966 4344 4606 4584 1 FreeSans 320 0 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_0/nmoscap_bot
flabel metal1 266 4014 506 4584 7 FreeSans 160 90 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_0/nmoscap_bot
flabel metal1 266 3004 506 3574 7 FreeSans 160 90 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_0/nmoscap_bot
flabel metal1 4366 3004 4606 3574 3 FreeSans 160 90 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_0/nmoscap_bot
flabel metal1 4366 4014 4606 4584 3 FreeSans 160 90 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_0/nmoscap_bot
flabel metal1 1386 3004 3486 3244 5 FreeSans 320 0 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_0/nmoscap_top
flabel metal1 1386 4344 3486 4584 1 FreeSans 320 0 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_0/nmoscap_top
flabel metal1 266 3614 506 3984 7 FreeSans 320 90 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_0/nmoscap_top
flabel metal1 4366 3604 4606 3974 3 FreeSans 320 90 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_0/nmoscap_top
flabel locali 916 3004 1376 3084 5 FreeSans 320 0 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_0/pwell
flabel locali 3496 3004 3956 3084 5 FreeSans 320 0 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_0/pwell
flabel locali 916 4504 1376 4584 1 FreeSans 320 0 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_0/pwell
flabel locali 3496 4504 3956 4584 1 FreeSans 320 0 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_0/pwell
flabel metal3 266 3004 906 3244 5 FreeSans 320 0 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_0/mimcap_bot
flabel metal3 3966 3004 4606 3244 5 FreeSans 320 0 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_0/mimcap_bot
flabel metal3 266 4344 906 4584 1 FreeSans 320 0 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_0/mimcap_bot
flabel metal3 3966 4344 4606 4584 1 FreeSans 320 0 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_0/mimcap_bot
flabel metal3 266 4104 516 4584 7 FreeSans 320 90 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_0/mimcap_bot
flabel metal3 266 3004 516 3484 7 FreeSans 320 90 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_0/mimcap_bot
flabel metal3 4356 3004 4606 3484 3 FreeSans 320 90 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_0/mimcap_bot
flabel metal3 4356 4104 4606 4584 3 FreeSans 320 90 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_0/mimcap_bot
flabel metal3 1386 3004 3486 3174 5 FreeSans 320 0 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_0/mimcap_top
flabel metal3 1386 4414 3486 4584 1 FreeSans 320 0 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_0/mimcap_top
flabel metal3 4436 3554 4606 4034 3 FreeSans 320 90 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_0/mimcap_top
flabel metal3 266 3554 436 4034 7 FreeSans 320 90 0 0 adc_comp_circuit_0/adc_noise_decoup_cell2_0/mimcap_top
rlabel locali 3122 5592 3122 5630 7 adc_comp_circuit_0/adc_comp_buffer_1/VSS
rlabel locali 3122 4888 3122 4926 7 adc_comp_circuit_0/adc_comp_buffer_1/VDD
rlabel locali 3572 5312 3572 5350 3 adc_comp_circuit_0/adc_comp_buffer_1/out
rlabel poly 3122 5322 3122 5378 7 adc_comp_circuit_0/adc_comp_buffer_1/in
rlabel locali 3122 5622 3122 5660 7 adc_comp_circuit_0/adc_comp_buffer_0/VSS
rlabel locali 3122 6326 3122 6364 7 adc_comp_circuit_0/adc_comp_buffer_0/VDD
rlabel locali 3572 5902 3572 5940 3 adc_comp_circuit_0/adc_comp_buffer_0/out
rlabel poly 3122 5874 3122 5930 7 adc_comp_circuit_0/adc_comp_buffer_0/in
rlabel locali 3938 4888 3938 4922 7 NOR_0/VDD
rlabel locali 4316 5314 4316 5352 3 NOR_0/Q
rlabel metal1 3882 5250 3882 5286 7 NOR_0/B
rlabel locali 3898 4956 3898 5008 7 NOR_0/A
rlabel locali 3970 5514 3970 5548 7 NOR_0/VSS
rlabel poly 3690 5904 3690 5936 7 NOR-Latch_0/R
rlabel metal1 3684 6274 3684 6306 7 NOR-Latch_0/S
rlabel locali 3778 6334 3778 6368 7 NOR-Latch_0/VDD
rlabel locali 4652 5904 4652 5944 3 NOR-Latch_0/QN
rlabel metal1 4656 5972 4656 6008 3 NOR-Latch_0/Q
rlabel locali 3808 5708 3808 5742 7 NOR-Latch_0/VSS
rlabel locali 4274 6334 4274 6368 7 NOR-Latch_0/NOR_1/VDD
rlabel locali 4652 5904 4652 5942 3 NOR-Latch_0/NOR_1/Q
rlabel metal1 4218 5970 4218 6006 7 NOR-Latch_0/NOR_1/B
rlabel locali 4234 6248 4234 6300 7 NOR-Latch_0/NOR_1/A
rlabel locali 4306 5708 4306 5742 7 NOR-Latch_0/NOR_1/VSS
rlabel locali 3778 6334 3778 6368 7 NOR-Latch_0/NOR_0/VDD
rlabel locali 4156 5904 4156 5942 3 NOR-Latch_0/NOR_0/Q
rlabel metal1 3722 5970 3722 6006 7 NOR-Latch_0/NOR_0/B
rlabel locali 3738 6248 3738 6300 7 NOR-Latch_0/NOR_0/A
rlabel locali 3810 5708 3810 5742 7 NOR-Latch_0/NOR_0/VSS
<< end >>
