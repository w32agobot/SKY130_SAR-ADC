* NGSPICE file created from adc_array_cap_16.ext - technology: sky130A

.subckt adc_array_circuit ROW_N COL_N COLON_N SAMPLE SAMPLE_N CBOT VCOM VDD VSS
X0 VINT2 COLON_N VDRV VSS sky130_fd_pr__nfet_01v8 ad=2.478e+11p pd=2.86e+06u as=2.52e+11p ps=2.88e+06u w=420000u l=180000u
X1 VINT2 ROW_N VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.26e+11p ps=1.44e+06u w=420000u l=180000u
X2 VSS COL_N VINT2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=180000u
X3 CBOT SAMPLE_N VCOM VDD sky130_fd_pr__pfet_01v8 ad=4.5e+11p pd=2.8e+06u as=4.5e+11p ps=2.8e+06u w=900000u l=180000u
X4 VDRV SAMPLE CBOT VDD sky130_fd_pr__pfet_01v8 ad=1.305e+12p pd=8.3e+06u as=0p ps=0u w=900000u l=180000u
X5 VINT COL_N VDRV VDD sky130_fd_pr__pfet_01v8 ad=4.5e+11p pd=2.8e+06u as=0p ps=0u w=900000u l=180000u
X6 CBOT SAMPLE_N VDRV VSS sky130_fd_pr__nfet_01v8 ad=1.26e+11p pd=1.44e+06u as=0p ps=0u w=420000u l=180000u
X7 VCOM SAMPLE CBOT VSS sky130_fd_pr__nfet_01v8 ad=1.26e+11p pd=1.44e+06u as=0p ps=0u w=420000u l=180000u
X8 VDD ROW_N VINT VDD sky130_fd_pr__pfet_01v8 ad=4.5e+11p pd=2.8e+06u as=0p ps=0u w=900000u l=180000u
X9 VDRV COLON_N VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=900000u l=180000u
.ends

.subckt adc_array_wafflecap_16x544aF_46um2 COL_N COLON_N CTOP ROW_N SAMPLE SAMPLE_N VCOM VDD CBOT VSS
Xadc_array_circuit_0 ROW_N COL_N COLON_N SAMPLE SAMPLE_N CBOT VCOM VDD VSS adc_array_circuit
.ends

