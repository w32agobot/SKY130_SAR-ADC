VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO delay_macrocell
  CLASS BLOCK ;
  FOREIGN delay_macrocell ;
  ORIGIN 0.190 0.240 ;
  SIZE 8.640 BY 3.210 ;
  PIN VPWR
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 8.260 2.810 ;
        RECT 0.050 1.500 0.220 2.380 ;
        RECT 4.890 1.520 5.060 2.630 ;
        RECT 6.600 1.350 6.770 2.630 ;
        RECT 6.600 1.180 7.150 1.350 ;
        RECT 6.980 0.380 7.150 1.180 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 0.050 1.580 0.220 2.300 ;
      LAYER met1 ;
        RECT 0.000 2.480 8.260 2.970 ;
        RECT 0.020 1.520 0.250 2.480 ;
    END
  END VPWR
  PIN in
    ANTENNAGATEAREA 5.040000 ;
    PORT
      LAYER li1 ;
        RECT -0.160 1.030 0.240 1.300 ;
    END
  END in
  PIN out
    ANTENNAGATEAREA 0.366000 ;
    ANTENNADIFFAREA 0.361800 ;
    PORT
      LAYER li1 ;
        RECT 5.850 1.520 6.020 2.360 ;
        RECT 6.260 1.010 6.430 1.340 ;
        RECT 5.960 0.380 6.130 0.890 ;
      LAYER mcon ;
        RECT 5.850 1.600 6.020 1.880 ;
        RECT 6.260 1.090 6.430 1.260 ;
        RECT 5.960 0.720 6.130 0.890 ;
      LAYER met1 ;
        RECT 5.820 1.240 6.050 2.030 ;
        RECT 6.230 1.240 6.460 1.320 ;
        RECT 5.820 1.100 8.260 1.240 ;
        RECT 5.930 1.030 6.460 1.100 ;
        RECT 5.930 0.660 6.160 1.030 ;
    END
  END out
  PIN VPB
    PORT
      LAYER nwell ;
        RECT -0.190 1.220 8.450 2.910 ;
    END
  END VPB
  PIN VGND
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 7.450 1.180 7.620 2.360 ;
        RECT 7.450 1.010 7.970 1.180 ;
        RECT 0.050 0.380 0.220 0.840 ;
        RECT 5.000 0.090 5.170 0.840 ;
        RECT 7.800 0.090 7.970 1.010 ;
        RECT 0.000 -0.090 8.260 0.090 ;
      LAYER mcon ;
        RECT 0.050 0.460 0.220 0.760 ;
        RECT 0.140 -0.090 0.320 0.090 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 6.825 -0.085 6.995 0.085 ;
        RECT 7.285 -0.085 7.455 0.085 ;
        RECT 7.745 -0.085 7.915 0.085 ;
      LAYER met1 ;
        RECT 0.020 0.240 0.250 0.820 ;
        RECT 4.320 0.240 4.840 0.590 ;
        RECT 0.000 -0.240 8.260 0.240 ;
      LAYER via ;
        RECT 4.420 0.290 4.740 0.550 ;
      LAYER met2 ;
        RECT 4.320 0.240 4.840 0.590 ;
      LAYER via2 ;
        RECT 4.420 0.300 4.740 0.580 ;
      LAYER met3 ;
        RECT 0.270 0.610 4.250 2.480 ;
        RECT 5.230 0.610 8.260 2.480 ;
        RECT 0.270 0.270 8.260 0.610 ;
    END
  END VGND
  PIN VNB
    ANTENNADIFFAREA 1.650000 ;
    PORT
      LAYER pwell ;
        RECT -0.190 -0.090 8.450 1.220 ;
    END
  END VNB
  OBS
      LAYER li1 ;
        RECT 4.340 1.290 4.510 2.380 ;
        RECT 5.370 1.520 5.540 2.360 ;
        RECT 6.940 1.520 7.140 2.360 ;
        RECT 7.930 1.520 8.130 2.360 ;
        RECT 4.340 1.010 4.930 1.290 ;
        RECT 4.340 0.380 4.510 1.010 ;
        RECT 5.480 0.380 5.650 0.840 ;
        RECT 6.500 0.380 6.670 0.840 ;
        RECT 7.460 0.380 7.630 0.840 ;
      LAYER mcon ;
        RECT 4.340 1.580 4.510 2.230 ;
        RECT 5.370 1.600 5.540 2.280 ;
        RECT 6.970 1.700 7.140 2.280 ;
        RECT 7.930 1.700 8.100 2.280 ;
        RECT 4.570 1.060 4.850 1.230 ;
        RECT 5.480 0.460 5.650 0.760 ;
        RECT 6.500 0.460 6.670 0.660 ;
        RECT 7.460 0.460 7.630 0.660 ;
      LAYER met1 ;
        RECT 4.310 1.290 4.540 2.340 ;
        RECT 5.340 2.170 8.130 2.340 ;
        RECT 5.340 1.540 5.570 2.170 ;
        RECT 6.940 1.640 7.170 2.170 ;
        RECT 7.900 1.640 8.130 2.170 ;
        RECT 4.310 1.010 4.930 1.290 ;
        RECT 5.450 0.520 5.680 0.820 ;
        RECT 6.470 0.520 6.700 0.720 ;
        RECT 7.430 0.520 7.660 0.720 ;
        RECT 5.450 0.380 7.660 0.520 ;
      LAYER via ;
        RECT 4.570 1.020 4.850 1.280 ;
      LAYER met2 ;
        RECT 4.550 1.290 4.920 1.450 ;
        RECT 4.490 1.010 4.920 1.290 ;
        RECT 4.550 0.840 4.920 1.010 ;
      LAYER via2 ;
        RECT 4.600 1.010 4.880 1.300 ;
      LAYER met3 ;
        RECT 4.550 0.910 4.930 1.590 ;
      LAYER via3 ;
        RECT 4.580 1.000 4.900 1.320 ;
      LAYER met4 ;
        RECT 4.550 1.340 4.960 1.450 ;
        RECT 3.660 0.970 5.990 1.340 ;
        RECT 4.550 0.840 4.960 0.970 ;
  END
END delay_macrocell
END LIBRARY

