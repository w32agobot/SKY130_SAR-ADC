VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO adc_clkgen_with_edgedetect
  CLASS BLOCK ;
  FOREIGN adc_clkgen_with_edgedetect ;
  ORIGIN 0.000 0.000 ;
  SIZE 171.000 BY 60.000 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 26.720 2.480 28.320 57.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 70.720 2.480 72.320 57.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 114.720 2.480 116.320 57.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 158.720 2.480 160.320 57.360 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 48.720 2.480 50.320 57.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 92.720 2.480 94.320 57.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 136.720 2.480 138.320 57.360 ;
    END
  END VSS
  PIN clk_comp_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 167.000 14.320 171.000 14.920 ;
    END
  END clk_comp_out
  PIN clk_dig_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.880 4.000 9.480 ;
    END
  END clk_dig_out
  PIN dlycontrol1_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.960 4.000 13.560 ;
    END
  END dlycontrol1_in[0]
  PIN dlycontrol1_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.000 4.000 15.600 ;
    END
  END dlycontrol1_in[1]
  PIN dlycontrol1_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END dlycontrol1_in[2]
  PIN dlycontrol1_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.080 4.000 19.680 ;
    END
  END dlycontrol1_in[3]
  PIN dlycontrol1_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.120 4.000 21.720 ;
    END
  END dlycontrol1_in[4]
  PIN dlycontrol2_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.160 4.000 23.760 ;
    END
  END dlycontrol2_in[0]
  PIN dlycontrol2_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.200 4.000 25.800 ;
    END
  END dlycontrol2_in[1]
  PIN dlycontrol2_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END dlycontrol2_in[2]
  PIN dlycontrol2_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.280 4.000 29.880 ;
    END
  END dlycontrol2_in[3]
  PIN dlycontrol2_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 31.320 4.000 31.920 ;
    END
  END dlycontrol2_in[4]
  PIN dlycontrol3_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 33.360 4.000 33.960 ;
    END
  END dlycontrol3_in[0]
  PIN dlycontrol3_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.400 4.000 36.000 ;
    END
  END dlycontrol3_in[1]
  PIN dlycontrol3_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END dlycontrol3_in[2]
  PIN dlycontrol3_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 39.480 4.000 40.080 ;
    END
  END dlycontrol3_in[3]
  PIN dlycontrol3_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 41.520 4.000 42.120 ;
    END
  END dlycontrol3_in[4]
  PIN dlycontrol4_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.560 4.000 44.160 ;
    END
  END dlycontrol4_in[0]
  PIN dlycontrol4_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 45.600 4.000 46.200 ;
    END
  END dlycontrol4_in[1]
  PIN dlycontrol4_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END dlycontrol4_in[2]
  PIN dlycontrol4_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.680 4.000 50.280 ;
    END
  END dlycontrol4_in[3]
  PIN dlycontrol4_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.720 4.000 52.320 ;
    END
  END dlycontrol4_in[4]
  PIN dlycontrol4_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.760 4.000 54.360 ;
    END
  END dlycontrol4_in[5]
  PIN ena_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.800 4.000 5.400 ;
    END
  END ena_in
  PIN enable_dlycontrol_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.920 4.000 11.520 ;
    END
  END enable_dlycontrol_in
  PIN ndecision_finish_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 167.000 44.240 171.000 44.840 ;
    END
  END ndecision_finish_in
  PIN nsample_n_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.810 0.000 107.090 4.000 ;
    END
  END nsample_n_in
  PIN nsample_n_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.590 0.000 149.870 4.000 ;
    END
  END nsample_n_out
  PIN nsample_p_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.810 56.000 107.090 60.000 ;
    END
  END nsample_p_in
  PIN nsample_p_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.590 56.000 149.870 60.000 ;
    END
  END nsample_p_out
  PIN sample_n_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.250 0.000 21.530 4.000 ;
    END
  END sample_n_in
  PIN sample_n_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.030 0.000 64.310 4.000 ;
    END
  END sample_n_out
  PIN sample_p_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.250 56.000 21.530 60.000 ;
    END
  END sample_p_in
  PIN sample_p_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.030 56.000 64.310 60.000 ;
    END
  END sample_p_out
  PIN start_conv_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END start_conv_in
  OBS
      LAYER li1 ;
        RECT 5.520 2.635 165.140 57.205 ;
      LAYER met1 ;
        RECT 5.520 0.040 165.140 59.800 ;
      LAYER met2 ;
        RECT 7.920 55.720 20.970 59.830 ;
        RECT 21.810 55.720 63.750 59.830 ;
        RECT 64.590 55.720 106.530 59.830 ;
        RECT 107.370 55.720 149.310 59.830 ;
        RECT 150.150 55.720 162.280 59.830 ;
        RECT 7.920 4.280 162.280 55.720 ;
        RECT 7.920 0.010 20.970 4.280 ;
        RECT 21.810 0.010 63.750 4.280 ;
        RECT 64.590 0.010 106.530 4.280 ;
        RECT 107.370 0.010 149.310 4.280 ;
        RECT 150.150 0.010 162.280 4.280 ;
      LAYER met3 ;
        RECT 4.000 54.760 167.000 59.665 ;
        RECT 4.400 53.360 167.000 54.760 ;
        RECT 4.000 52.720 167.000 53.360 ;
        RECT 4.400 51.320 167.000 52.720 ;
        RECT 4.000 50.680 167.000 51.320 ;
        RECT 4.400 49.280 167.000 50.680 ;
        RECT 4.000 48.640 167.000 49.280 ;
        RECT 4.400 47.240 167.000 48.640 ;
        RECT 4.000 46.600 167.000 47.240 ;
        RECT 4.400 45.240 167.000 46.600 ;
        RECT 4.400 45.200 166.600 45.240 ;
        RECT 4.000 44.560 166.600 45.200 ;
        RECT 4.400 43.840 166.600 44.560 ;
        RECT 4.400 43.160 167.000 43.840 ;
        RECT 4.000 42.520 167.000 43.160 ;
        RECT 4.400 41.120 167.000 42.520 ;
        RECT 4.000 40.480 167.000 41.120 ;
        RECT 4.400 39.080 167.000 40.480 ;
        RECT 4.000 38.440 167.000 39.080 ;
        RECT 4.400 37.040 167.000 38.440 ;
        RECT 4.000 36.400 167.000 37.040 ;
        RECT 4.400 35.000 167.000 36.400 ;
        RECT 4.000 34.360 167.000 35.000 ;
        RECT 4.400 32.960 167.000 34.360 ;
        RECT 4.000 32.320 167.000 32.960 ;
        RECT 4.400 30.920 167.000 32.320 ;
        RECT 4.000 30.280 167.000 30.920 ;
        RECT 4.400 28.880 167.000 30.280 ;
        RECT 4.000 28.240 167.000 28.880 ;
        RECT 4.400 26.840 167.000 28.240 ;
        RECT 4.000 26.200 167.000 26.840 ;
        RECT 4.400 24.800 167.000 26.200 ;
        RECT 4.000 24.160 167.000 24.800 ;
        RECT 4.400 22.760 167.000 24.160 ;
        RECT 4.000 22.120 167.000 22.760 ;
        RECT 4.400 20.720 167.000 22.120 ;
        RECT 4.000 20.080 167.000 20.720 ;
        RECT 4.400 18.680 167.000 20.080 ;
        RECT 4.000 18.040 167.000 18.680 ;
        RECT 4.400 16.640 167.000 18.040 ;
        RECT 4.000 16.000 167.000 16.640 ;
        RECT 4.400 15.320 167.000 16.000 ;
        RECT 4.400 14.600 166.600 15.320 ;
        RECT 4.000 13.960 166.600 14.600 ;
        RECT 4.400 13.920 166.600 13.960 ;
        RECT 4.400 12.560 167.000 13.920 ;
        RECT 4.000 11.920 167.000 12.560 ;
        RECT 4.400 10.520 167.000 11.920 ;
        RECT 4.000 9.880 167.000 10.520 ;
        RECT 4.400 8.480 167.000 9.880 ;
        RECT 4.000 7.840 167.000 8.480 ;
        RECT 4.400 6.440 167.000 7.840 ;
        RECT 4.000 5.800 167.000 6.440 ;
        RECT 4.400 4.400 167.000 5.800 ;
        RECT 4.000 0.175 167.000 4.400 ;
      LAYER met4 ;
        RECT 17.775 12.415 26.320 53.545 ;
        RECT 28.720 12.415 48.320 53.545 ;
        RECT 50.720 12.415 63.185 53.545 ;
  END
END adc_clkgen_with_edgedetect
END LIBRARY

