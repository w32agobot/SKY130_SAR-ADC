magic
tech sky130A
timestamp 1662366209
<< nwell >>
rect 0 89 104 288
<< nmos >>
rect 31 11 73 26
<< pmos >>
rect 31 182 75 197
rect 31 136 75 151
<< ndiff >>
rect 31 49 73 55
rect 31 32 37 49
rect 67 32 73 49
rect 31 26 73 32
rect 31 5 73 11
rect 31 -12 37 5
rect 67 -12 73 5
rect 31 -18 73 -12
<< pdiff >>
rect 31 221 75 225
rect 31 204 37 221
rect 67 204 75 221
rect 31 197 75 204
rect 31 175 75 182
rect 31 158 37 175
rect 67 158 75 175
rect 31 151 75 158
rect 31 130 75 136
rect 31 113 37 130
rect 67 113 75 130
rect 31 107 75 113
<< ndiffc >>
rect 37 32 67 49
rect 37 -12 67 5
<< pdiffc >>
rect 37 204 67 221
rect 37 158 67 175
rect 37 113 67 130
<< psubdiff >>
rect 31 -62 43 -45
rect 61 -62 73 -45
rect 31 -65 73 -62
<< nsubdiff >>
rect 31 252 43 270
rect 61 252 73 270
<< psubdiffcont >>
rect 43 -62 61 -45
<< nsubdiffcont >>
rect 43 252 61 270
<< poly >>
rect 8 182 31 197
rect 75 182 88 197
rect 8 151 23 182
rect 8 136 31 151
rect 75 136 88 151
rect 8 94 23 136
rect -13 86 23 94
rect -13 69 -5 86
rect 12 69 23 86
rect -13 61 23 69
rect 8 26 23 61
rect 8 11 31 26
rect 73 11 86 26
<< polycont >>
rect -5 69 12 86
<< locali >>
rect -13 271 43 288
rect 61 271 73 288
rect -13 270 73 271
rect -13 268 43 270
rect -13 176 5 268
rect 31 252 43 268
rect 61 252 73 270
rect 31 222 75 225
rect 29 221 77 222
rect 29 204 37 221
rect 67 204 77 221
rect 29 203 77 204
rect -13 175 77 176
rect -13 158 37 175
rect 67 158 77 175
rect -13 157 77 158
rect 29 113 37 130
rect 67 113 77 130
rect 31 107 75 113
rect -13 86 14 94
rect -13 69 -5 86
rect 12 69 14 86
rect -13 61 14 69
rect 31 89 73 107
rect 31 66 104 89
rect 31 49 73 66
rect 29 32 37 49
rect 67 32 75 49
rect 31 29 73 32
rect 29 -12 37 5
rect 67 -12 75 5
rect 31 -45 73 -12
rect 31 -62 43 -45
rect 61 -62 73 -45
rect 31 -65 73 -62
<< viali >>
rect 43 271 61 288
rect 37 204 67 221
rect 37 113 67 130
rect 43 -62 61 -45
<< metal1 >>
rect 27 288 76 291
rect 27 271 43 288
rect 61 271 76 288
rect 27 268 76 271
rect 33 221 72 228
rect 33 204 37 221
rect 67 204 72 221
rect 33 130 72 204
rect 33 113 37 130
rect 67 113 72 130
rect 33 107 72 113
rect 28 -45 76 -42
rect 28 -62 43 -45
rect 61 -62 76 -45
rect 28 -65 76 -62
<< labels >>
rlabel locali -13 66 -13 89 7 in
rlabel locali 104 66 104 89 3 out
rlabel metal1 28 -65 28 -42 7 VSS
port 2 w
rlabel metal1 27 268 27 291 7 VDD
port 1 w
<< end >>
