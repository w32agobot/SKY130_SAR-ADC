magic
tech sky130A
timestamp 1664529495
<< nwell >>
rect 0 253 502 440
<< nmos >>
rect 116 126 131 168
rect 164 126 179 168
rect 268 126 283 168
rect 316 126 331 168
rect 364 126 379 168
<< pmos >>
rect 116 271 131 351
rect 164 271 179 351
rect 268 287 283 367
rect 316 287 331 367
rect 364 287 379 367
<< ndiff >>
rect 85 162 116 168
rect 85 132 91 162
rect 108 132 116 162
rect 85 126 116 132
rect 131 162 164 168
rect 131 132 139 162
rect 156 132 164 162
rect 131 126 164 132
rect 179 162 210 168
rect 179 132 187 162
rect 204 132 210 162
rect 179 126 210 132
rect 237 162 268 168
rect 237 132 243 162
rect 260 132 268 162
rect 237 126 268 132
rect 283 162 316 168
rect 283 132 291 162
rect 308 132 316 162
rect 283 126 316 132
rect 331 162 364 168
rect 331 132 339 162
rect 356 132 364 162
rect 331 126 364 132
rect 379 162 410 168
rect 379 132 387 162
rect 404 132 410 162
rect 379 126 410 132
<< pdiff >>
rect 237 361 268 367
rect 85 345 116 351
rect 85 277 91 345
rect 108 277 116 345
rect 85 271 116 277
rect 131 345 164 351
rect 131 277 139 345
rect 156 277 164 345
rect 131 271 164 277
rect 179 345 210 351
rect 179 277 187 345
rect 204 277 210 345
rect 237 293 243 361
rect 260 293 268 361
rect 237 287 268 293
rect 283 361 316 367
rect 283 293 291 361
rect 308 293 316 361
rect 283 287 316 293
rect 331 361 364 367
rect 331 293 339 361
rect 356 293 364 361
rect 331 287 364 293
rect 379 361 410 367
rect 379 293 387 361
rect 404 293 410 361
rect 379 287 410 293
rect 179 271 210 277
<< ndiffc >>
rect 91 132 108 162
rect 139 132 156 162
rect 187 132 204 162
rect 243 132 260 162
rect 291 132 308 162
rect 339 132 356 162
rect 387 132 404 162
<< pdiffc >>
rect 91 277 108 345
rect 139 277 156 345
rect 187 277 204 345
rect 243 293 260 361
rect 291 293 308 361
rect 339 293 356 361
rect 387 293 404 361
<< psubdiff >>
rect 91 74 115 91
rect 132 74 163 91
rect 180 74 192 91
rect 339 74 363 91
rect 380 74 396 91
<< nsubdiff >>
rect 151 419 403 422
rect 151 402 163 419
rect 180 402 215 419
rect 232 402 267 419
rect 284 402 315 419
rect 332 402 362 419
rect 379 402 403 419
rect 151 399 403 402
<< psubdiffcont >>
rect 115 74 132 91
rect 163 74 180 91
rect 363 74 380 91
<< nsubdiffcont >>
rect 163 402 180 419
rect 215 402 232 419
rect 267 402 284 419
rect 315 402 332 419
rect 362 402 379 419
<< poly >>
rect 106 409 140 414
rect 106 391 114 409
rect 132 391 140 409
rect 106 359 140 391
rect 268 367 283 380
rect 316 367 331 380
rect 364 367 379 380
rect 116 351 131 359
rect 164 351 179 364
rect 116 168 131 271
rect 164 254 179 271
rect 268 268 283 287
rect 316 274 331 287
rect 364 279 379 287
rect 364 274 417 279
rect 164 244 198 254
rect 164 225 173 244
rect 190 225 198 244
rect 164 176 198 225
rect 247 199 283 268
rect 304 258 417 274
rect 304 240 338 258
rect 312 215 330 240
rect 383 238 417 258
rect 312 213 338 215
rect 268 196 283 199
rect 304 196 338 213
rect 268 181 379 196
rect 164 168 179 176
rect 268 168 283 181
rect 316 168 331 181
rect 364 168 379 181
rect 116 113 131 126
rect 164 113 179 126
rect 268 113 283 126
rect 316 113 331 126
rect 364 113 379 126
rect 268 103 331 113
rect 255 98 331 103
rect 253 81 261 98
rect 278 81 295 98
rect 312 81 320 98
rect 253 75 320 81
<< polycont >>
rect 114 391 132 409
rect 173 225 190 244
rect 261 81 278 98
rect 295 81 312 98
<< locali >>
rect 17 353 74 502
rect 427 460 485 502
rect 151 419 403 422
rect 114 409 132 417
rect 151 402 163 419
rect 180 402 215 419
rect 232 402 267 419
rect 284 402 315 419
rect 332 402 362 419
rect 379 402 403 419
rect 151 399 403 402
rect 114 386 132 391
rect 114 369 115 386
rect 187 361 260 369
rect 17 345 108 353
rect 17 277 91 345
rect 17 187 108 277
rect 139 345 156 353
rect 17 133 74 187
rect 17 116 57 133
rect 91 168 114 170
rect 91 162 97 168
rect 108 146 114 151
rect 139 162 156 277
rect 187 350 243 361
rect 187 345 216 350
rect 204 332 216 345
rect 233 332 243 350
rect 204 311 243 332
rect 204 293 216 311
rect 233 293 243 311
rect 204 285 260 293
rect 291 361 308 399
rect 291 285 308 293
rect 339 361 356 381
rect 204 277 238 285
rect 339 280 356 293
rect 387 361 404 369
rect 387 285 404 293
rect 187 269 238 277
rect 173 244 190 252
rect 173 207 190 225
rect 173 187 190 190
rect 207 187 238 269
rect 221 170 238 187
rect 91 124 108 132
rect 139 124 156 132
rect 187 162 204 170
rect 221 168 260 170
rect 221 151 229 168
rect 246 162 260 168
rect 221 150 243 151
rect 187 130 204 132
rect 17 0 74 116
rect 243 124 260 132
rect 291 162 308 170
rect 291 124 308 132
rect 339 162 356 170
rect 187 110 204 113
rect 261 98 278 103
rect 295 98 312 103
rect 91 74 115 91
rect 132 74 163 91
rect 180 74 192 91
rect 253 81 261 98
rect 278 81 295 98
rect 312 81 320 98
rect 339 91 356 132
rect 387 162 404 170
rect 387 124 404 132
rect 261 0 278 81
rect 295 75 312 81
rect 339 74 363 91
rect 380 74 396 91
rect 422 28 485 460
rect 427 0 485 28
<< viali >>
rect 163 402 180 419
rect 215 402 232 419
rect 267 402 284 419
rect 315 402 332 419
rect 362 402 379 419
rect 115 369 132 386
rect 139 326 156 344
rect 139 287 156 305
rect 57 116 74 133
rect 97 162 114 168
rect 97 151 108 162
rect 108 151 114 162
rect 216 332 233 350
rect 216 293 233 311
rect 387 332 404 350
rect 387 293 404 311
rect 173 190 190 207
rect 229 162 246 168
rect 229 151 243 162
rect 243 151 246 162
rect 187 113 204 130
rect 291 145 308 162
rect 115 74 132 91
rect 163 74 180 91
rect 387 145 404 162
rect 363 74 380 91
<< metal1 >>
rect 0 419 502 427
rect 0 403 163 419
rect 0 399 98 403
rect 149 402 163 403
rect 180 402 215 419
rect 232 402 267 419
rect 284 402 315 419
rect 332 402 362 419
rect 379 402 502 419
rect 149 399 502 402
rect 109 386 138 389
rect 109 385 115 386
rect 0 370 115 385
rect 109 369 115 370
rect 132 385 138 386
rect 132 370 502 385
rect 132 369 138 370
rect 109 366 138 369
rect 133 349 162 351
rect 213 350 236 356
rect 132 323 135 349
rect 161 323 164 349
rect 132 310 164 323
rect 132 284 135 310
rect 161 284 164 310
rect 213 332 216 350
rect 233 333 236 350
rect 384 350 407 356
rect 384 333 387 350
rect 233 332 387 333
rect 404 332 407 350
rect 213 319 407 332
rect 213 311 236 319
rect 213 293 216 311
rect 233 293 236 311
rect 213 287 236 293
rect 384 311 407 319
rect 384 293 387 311
rect 404 293 407 311
rect 384 287 407 293
rect 387 284 404 287
rect 0 256 502 270
rect 248 243 277 256
rect 83 229 225 239
rect 297 229 328 232
rect 385 229 415 242
rect 0 224 502 229
rect 0 215 97 224
rect 211 215 502 224
rect 167 207 196 210
rect 297 209 328 215
rect 167 201 173 207
rect 0 190 173 201
rect 190 201 196 207
rect 190 195 283 201
rect 368 195 502 201
rect 190 190 502 195
rect 0 187 502 190
rect 167 184 196 187
rect 265 181 408 187
rect 91 168 120 173
rect 91 151 97 168
rect 114 164 120 168
rect 223 168 252 173
rect 223 164 229 168
rect 114 151 229 164
rect 246 151 252 168
rect 91 150 252 151
rect 91 146 120 150
rect 223 146 252 150
rect 285 162 410 166
rect 285 145 291 162
rect 308 145 387 162
rect 404 145 410 162
rect 285 142 410 145
rect 54 133 77 139
rect 54 124 57 133
rect 0 116 57 124
rect 74 124 77 133
rect 184 130 208 136
rect 184 124 187 130
rect 74 116 187 124
rect 0 113 187 116
rect 204 124 208 130
rect 204 113 502 124
rect 0 110 502 113
rect 0 91 502 96
rect 0 74 115 91
rect 132 74 163 91
rect 180 74 363 91
rect 380 74 502 91
rect 0 68 502 74
<< via1 >>
rect 135 344 161 349
rect 135 326 139 344
rect 139 326 156 344
rect 156 326 161 344
rect 135 323 161 326
rect 135 305 161 310
rect 135 287 139 305
rect 139 287 156 305
rect 156 287 161 305
rect 135 284 161 287
<< metal2 >>
rect 16 481 486 486
rect 16 453 21 481
rect 49 453 69 481
rect 97 453 117 481
rect 145 453 165 481
rect 193 453 213 481
rect 241 453 261 481
rect 289 453 309 481
rect 337 453 357 481
rect 385 453 405 481
rect 433 453 453 481
rect 481 453 486 481
rect 16 433 486 453
rect 16 405 21 433
rect 49 405 165 433
rect 193 405 309 433
rect 337 405 453 433
rect 481 405 486 433
rect 16 385 486 405
rect 16 357 21 385
rect 49 357 165 385
rect 193 357 309 385
rect 337 357 453 385
rect 481 357 486 385
rect 16 349 486 357
rect 16 337 135 349
rect 161 337 486 349
rect 16 309 21 337
rect 49 309 69 337
rect 97 309 117 337
rect 161 323 165 337
rect 145 310 165 323
rect 161 309 165 310
rect 193 309 213 337
rect 241 309 261 337
rect 289 309 309 337
rect 337 309 357 337
rect 385 309 405 337
rect 433 309 453 337
rect 481 309 486 337
rect 16 289 135 309
rect 16 261 21 289
rect 49 284 135 289
rect 161 304 486 309
rect 161 289 198 304
rect 161 284 165 289
rect 49 261 165 284
rect 193 261 198 289
rect 304 289 486 304
rect 16 241 198 261
rect 16 213 21 241
rect 49 213 165 241
rect 193 213 198 241
rect 230 230 272 272
rect 304 261 309 289
rect 337 261 453 289
rect 481 261 486 289
rect 304 241 486 261
rect 16 198 198 213
rect 304 213 309 241
rect 337 213 453 241
rect 481 213 486 241
rect 304 198 486 213
rect 16 193 486 198
rect 16 165 21 193
rect 49 165 69 193
rect 97 165 117 193
rect 145 165 165 193
rect 193 165 213 193
rect 241 165 261 193
rect 289 165 309 193
rect 337 165 357 193
rect 385 165 405 193
rect 433 165 453 193
rect 481 165 486 193
rect 16 145 486 165
rect 16 117 21 145
rect 49 117 165 145
rect 193 117 309 145
rect 337 117 453 145
rect 481 117 486 145
rect 16 97 486 117
rect 16 69 21 97
rect 49 69 165 97
rect 193 69 309 97
rect 337 69 453 97
rect 481 69 486 97
rect 16 49 486 69
rect 16 21 21 49
rect 49 21 69 49
rect 97 21 117 49
rect 145 21 165 49
rect 193 21 213 49
rect 241 21 261 49
rect 289 21 309 49
rect 337 21 357 49
rect 385 21 405 49
rect 433 21 453 49
rect 481 21 486 49
rect 16 16 486 21
<< via2 >>
rect 21 453 49 481
rect 69 453 97 481
rect 117 453 145 481
rect 165 453 193 481
rect 213 453 241 481
rect 261 453 289 481
rect 309 453 337 481
rect 357 453 385 481
rect 405 453 433 481
rect 453 453 481 481
rect 21 405 49 433
rect 165 405 193 433
rect 309 405 337 433
rect 453 405 481 433
rect 21 357 49 385
rect 165 357 193 385
rect 309 357 337 385
rect 453 357 481 385
rect 21 309 49 337
rect 69 309 97 337
rect 117 323 135 337
rect 135 323 145 337
rect 117 310 145 323
rect 117 309 135 310
rect 135 309 145 310
rect 165 309 193 337
rect 213 309 241 337
rect 261 309 289 337
rect 309 309 337 337
rect 357 309 385 337
rect 405 309 433 337
rect 453 309 481 337
rect 21 261 49 289
rect 165 261 193 289
rect 21 213 49 241
rect 165 213 193 241
rect 309 261 337 289
rect 453 261 481 289
rect 309 213 337 241
rect 453 213 481 241
rect 21 165 49 193
rect 69 165 97 193
rect 117 165 145 193
rect 165 165 193 193
rect 213 165 241 193
rect 261 165 289 193
rect 309 165 337 193
rect 357 165 385 193
rect 405 165 433 193
rect 453 165 481 193
rect 21 117 49 145
rect 165 117 193 145
rect 309 117 337 145
rect 453 117 481 145
rect 21 69 49 97
rect 165 69 193 97
rect 309 69 337 97
rect 453 69 481 97
rect 21 21 49 49
rect 69 21 97 49
rect 117 21 145 49
rect 165 21 193 49
rect 213 21 241 49
rect 261 21 289 49
rect 309 21 337 49
rect 357 21 385 49
rect 405 21 433 49
rect 453 21 481 49
<< metal3 >>
rect 18 481 484 484
rect 18 453 21 481
rect 49 453 69 481
rect 97 453 117 481
rect 145 453 165 481
rect 193 453 213 481
rect 241 453 261 481
rect 289 453 309 481
rect 337 453 357 481
rect 385 453 405 481
rect 433 453 453 481
rect 481 453 484 481
rect 18 450 484 453
rect 18 433 52 450
rect 18 405 21 433
rect 49 405 52 433
rect 162 433 196 450
rect 18 385 52 405
rect 18 357 21 385
rect 49 357 52 385
rect 82 412 132 420
rect 82 378 90 412
rect 124 378 132 412
rect 82 370 132 378
rect 162 405 165 433
rect 193 405 196 433
rect 306 433 340 450
rect 162 385 196 405
rect 18 340 52 357
rect 162 357 165 385
rect 193 357 196 385
rect 226 412 276 420
rect 226 378 234 412
rect 268 378 276 412
rect 226 370 276 378
rect 306 405 309 433
rect 337 405 340 433
rect 450 433 484 450
rect 306 385 340 405
rect 162 340 196 357
rect 306 357 309 385
rect 337 357 340 385
rect 370 412 420 420
rect 370 378 378 412
rect 412 378 420 412
rect 370 370 420 378
rect 450 405 453 433
rect 481 405 484 433
rect 450 385 484 405
rect 306 340 340 357
rect 450 357 453 385
rect 481 357 484 385
rect 450 340 484 357
rect 18 337 484 340
rect 18 309 21 337
rect 49 309 69 337
rect 97 309 117 337
rect 145 309 165 337
rect 193 309 213 337
rect 241 309 261 337
rect 289 309 309 337
rect 337 309 357 337
rect 385 309 405 337
rect 433 309 453 337
rect 481 309 484 337
rect 18 306 484 309
rect 18 289 52 306
rect 18 261 21 289
rect 49 261 52 289
rect 162 289 196 306
rect 18 241 52 261
rect 18 213 21 241
rect 49 213 52 241
rect 82 268 132 276
rect 82 234 90 268
rect 124 234 132 268
rect 82 226 132 234
rect 162 261 165 289
rect 193 261 196 289
rect 162 241 196 261
rect 18 196 52 213
rect 162 213 165 241
rect 193 213 196 241
rect 162 196 196 213
rect 306 289 340 306
rect 306 261 309 289
rect 337 261 340 289
rect 450 289 484 306
rect 306 241 340 261
rect 306 213 309 241
rect 337 213 340 241
rect 370 268 420 276
rect 370 234 378 268
rect 412 234 420 268
rect 370 226 420 234
rect 450 261 453 289
rect 481 261 484 289
rect 450 241 484 261
rect 306 196 340 213
rect 450 213 453 241
rect 481 213 484 241
rect 450 196 484 213
rect 18 193 484 196
rect 18 165 21 193
rect 49 165 69 193
rect 97 165 117 193
rect 145 165 165 193
rect 193 165 213 193
rect 241 165 261 193
rect 289 165 309 193
rect 337 165 357 193
rect 385 165 405 193
rect 433 165 453 193
rect 481 165 484 193
rect 18 162 484 165
rect 18 145 52 162
rect 18 117 21 145
rect 49 117 52 145
rect 162 145 196 162
rect 18 97 52 117
rect 18 69 21 97
rect 49 69 52 97
rect 82 124 132 132
rect 82 90 90 124
rect 124 90 132 124
rect 82 82 132 90
rect 162 117 165 145
rect 193 117 196 145
rect 306 145 340 162
rect 162 97 196 117
rect 18 52 52 69
rect 162 69 165 97
rect 193 69 196 97
rect 226 124 276 132
rect 226 90 234 124
rect 268 90 276 124
rect 226 82 276 90
rect 306 117 309 145
rect 337 117 340 145
rect 450 145 484 162
rect 306 97 340 117
rect 162 52 196 69
rect 306 69 309 97
rect 337 69 340 97
rect 370 124 420 132
rect 370 90 378 124
rect 412 90 420 124
rect 370 82 420 90
rect 450 117 453 145
rect 481 117 484 145
rect 450 97 484 117
rect 306 52 340 69
rect 450 69 453 97
rect 481 69 484 97
rect 450 52 484 69
rect 18 49 484 52
rect 18 21 21 49
rect 49 21 69 49
rect 97 21 117 49
rect 145 21 165 49
rect 193 21 213 49
rect 241 21 261 49
rect 289 21 309 49
rect 337 21 357 49
rect 385 21 405 49
rect 433 21 453 49
rect 481 21 484 49
rect 18 18 484 21
<< via3 >>
rect 90 378 124 412
rect 234 378 268 412
rect 378 378 412 412
rect 90 234 124 268
rect 378 234 412 268
rect 90 90 124 124
rect 234 90 268 124
rect 378 90 412 124
<< metal4 >>
rect 92 420 122 467
rect 236 420 266 467
rect 380 420 410 467
rect 82 412 132 420
rect 82 410 90 412
rect 35 380 90 410
rect 82 378 90 380
rect 124 410 132 412
rect 226 412 276 420
rect 226 410 234 412
rect 124 380 234 410
rect 124 378 132 380
rect 82 370 132 378
rect 226 378 234 380
rect 268 410 276 412
rect 370 412 420 420
rect 268 380 323 410
rect 268 378 276 380
rect 226 370 276 378
rect 370 378 378 412
rect 412 410 420 412
rect 412 380 467 410
rect 412 378 420 380
rect 370 370 420 378
rect 92 323 122 370
rect 236 323 266 370
rect 380 276 410 370
rect 82 268 132 276
rect 82 266 90 268
rect 35 236 90 266
rect 82 234 90 236
rect 124 266 132 268
rect 370 268 420 276
rect 370 266 378 268
rect 124 236 179 266
rect 323 236 378 266
rect 124 234 132 236
rect 82 226 132 234
rect 370 234 378 236
rect 412 266 420 268
rect 412 236 467 266
rect 412 234 420 236
rect 370 226 420 234
rect 92 132 122 226
rect 236 132 266 179
rect 380 132 410 226
rect 82 124 132 132
rect 82 122 90 124
rect 35 92 90 122
rect 82 90 90 92
rect 124 122 132 124
rect 226 124 276 132
rect 226 122 234 124
rect 124 92 234 122
rect 124 90 132 92
rect 82 82 132 90
rect 226 90 234 92
rect 268 122 276 124
rect 370 124 420 132
rect 370 122 378 124
rect 268 92 378 122
rect 268 90 276 92
rect 226 82 276 90
rect 370 90 378 92
rect 412 122 420 124
rect 412 92 467 122
rect 412 90 420 92
rect 370 82 420 90
rect 92 35 122 82
rect 236 35 266 82
rect 380 35 410 82
<< comment >>
rect 0 486 16 502
rect 486 486 502 502
rect 288 288 304 304
rect 272 272 288 288
rect 214 214 230 230
rect 198 198 214 214
rect 0 0 16 16
rect 486 0 502 16
<< labels >>
rlabel metal1 0 399 0 427 7 VDD
port 1 w
rlabel metal1 0 370 0 385 7 sample_n
port 2 w
rlabel metal1 0 256 0 270 7 colon_n
port 3 w
rlabel metal1 0 215 0 229 7 col_n
port 4 w
rlabel metal1 0 187 0 201 7 sample
port 5 w
rlabel metal1 0 110 0 124 7 vcom
port 6 w
rlabel metal1 0 68 0 96 7 VSS
port 7 w
rlabel locali 427 0 485 0 5 row_n
port 8 s
rlabel locali 261 0 278 0 5 en_n
port 9 s
rlabel metal4 92 467 122 467 1 ctop
port 10 n
<< end >>
