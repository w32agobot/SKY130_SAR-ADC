magic
tech sky130A
magscale 1 2
timestamp 1658837386
<< nwell >>
rect -209 -116 209 116
<< pmos >>
rect -111 -80 -81 80
rect -15 -80 15 80
rect 81 -80 111 80
<< pdiff >>
rect -173 68 -111 80
rect -173 -68 -161 68
rect -127 -68 -111 68
rect -173 -80 -111 -68
rect -81 68 -15 80
rect -81 -68 -65 68
rect -31 -68 -15 68
rect -81 -80 -15 -68
rect 15 68 81 80
rect 15 -68 31 68
rect 65 -68 81 68
rect 15 -80 81 -68
rect 111 68 173 80
rect 111 -68 127 68
rect 161 -68 173 68
rect 111 -80 173 -68
<< pdiffc >>
rect -161 -68 -127 68
rect -65 -68 -31 68
rect 31 -68 65 68
rect 127 -68 161 68
<< poly >>
rect -111 80 -81 106
rect -15 80 15 106
rect 81 80 111 106
rect -111 -106 -81 -80
rect -15 -106 15 -80
rect 81 -106 111 -80
<< locali >>
rect -161 68 -127 84
rect -161 -84 -127 -68
rect -65 68 -31 84
rect -65 -84 -31 -68
rect 31 68 65 84
rect 31 -84 65 -68
rect 127 68 161 84
rect 127 -84 161 -68
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.8 l 0.15 m 1 nf 3 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
