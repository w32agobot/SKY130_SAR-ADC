magic
tech sky130A
magscale 1 2
timestamp 1673912611
<< error_s >>
rect 2997 276 3984 345
rect 185 -470 261 -461
rect 620 -468 695 -459
rect 185 -526 190 -470
rect 620 -524 634 -468
rect 185 -533 261 -526
rect 620 -531 695 -524
rect 3447 -970 3481 -936
rect 3519 -970 3553 -936
rect 3591 -970 3625 -936
rect 3663 -970 3697 -936
rect 3735 -970 3769 -936
rect 2926 -1202 3145 -984
rect 3180 -1202 3830 -1108
rect 2926 -1238 3866 -1202
rect 3145 -1312 3866 -1238
<< nwell >>
rect 878 186 3984 276
rect 878 177 3024 186
rect 3068 177 3984 186
rect 878 -73 2727 177
rect 3145 -65 3165 177
rect -676 -144 2727 -73
rect -676 -413 2656 -144
rect -676 -480 -190 -413
rect -674 -482 -190 -480
rect -674 -566 -218 -482
rect 2787 -1276 2825 -1238
rect 2863 -1276 2901 -1238
rect 2939 -1276 2977 -1238
rect 3015 -1276 3053 -1238
rect 3180 -1276 3830 -1238
<< nmos >>
rect 30 -1170 60 -1070
rect 118 -1170 148 -1070
rect 206 -1170 236 -1070
rect 294 -1170 324 -1070
rect 382 -1170 412 -1070
rect 470 -1170 500 -1070
rect 558 -1170 588 -1070
rect 646 -1170 676 -1070
rect 734 -1170 764 -1070
rect 822 -1170 852 -1070
rect 1525 -1188 1555 -788
rect 1617 -1188 1647 -788
rect 1713 -1188 1743 -788
rect 1809 -1188 1839 -788
rect 1905 -1188 1935 -788
rect 1997 -1188 2027 -788
<< pmos >>
rect 12 -343 42 -243
rect 104 -343 134 -243
rect 196 -343 226 -243
rect 288 -343 318 -243
rect 380 -343 410 -243
rect 472 -343 502 -243
rect 564 -343 594 -243
rect 656 -343 686 -243
rect 748 -343 778 -243
rect 840 -343 870 -243
rect 1148 -348 1178 52
rect 1236 -348 1266 52
rect 1324 -348 1354 52
rect 1412 -348 1442 52
rect 1500 -348 1530 52
rect 1588 -348 1618 52
rect 1935 -348 1965 52
rect 2023 -348 2053 52
rect 2111 -348 2141 52
rect 2199 -348 2229 52
rect 2287 -348 2317 52
rect 2375 -348 2405 52
<< nmoslvt >>
rect 30 -973 60 -573
rect 118 -973 148 -573
rect 206 -973 236 -573
rect 294 -973 324 -573
rect 382 -973 412 -573
rect 470 -973 500 -573
rect 558 -973 588 -573
rect 646 -973 676 -573
rect 734 -973 764 -573
rect 822 -973 852 -573
<< ndiff >>
rect -28 -585 30 -573
rect -28 -961 -16 -585
rect 18 -961 30 -585
rect -28 -973 30 -961
rect 60 -585 118 -573
rect 60 -961 72 -585
rect 106 -961 118 -585
rect 60 -973 118 -961
rect 148 -585 206 -573
rect 148 -961 160 -585
rect 194 -961 206 -585
rect 148 -973 206 -961
rect 236 -585 294 -573
rect 236 -961 248 -585
rect 282 -961 294 -585
rect 236 -973 294 -961
rect 324 -585 382 -573
rect 324 -961 336 -585
rect 370 -961 382 -585
rect 324 -973 382 -961
rect 412 -585 470 -573
rect 412 -961 424 -585
rect 458 -961 470 -585
rect 412 -973 470 -961
rect 500 -585 558 -573
rect 500 -961 512 -585
rect 546 -961 558 -585
rect 500 -973 558 -961
rect 588 -585 646 -573
rect 588 -961 600 -585
rect 634 -961 646 -585
rect 588 -973 646 -961
rect 676 -585 734 -573
rect 676 -961 688 -585
rect 722 -961 734 -585
rect 676 -973 734 -961
rect 764 -585 822 -573
rect 764 -961 776 -585
rect 810 -961 822 -585
rect 764 -973 822 -961
rect 852 -585 910 -573
rect 852 -961 864 -585
rect 898 -961 910 -585
rect 852 -973 910 -961
rect 1463 -800 1525 -788
rect -28 -1082 30 -1070
rect -28 -1158 -16 -1082
rect 18 -1158 30 -1082
rect -28 -1170 30 -1158
rect 60 -1082 118 -1070
rect 60 -1158 72 -1082
rect 106 -1158 118 -1082
rect 60 -1170 118 -1158
rect 148 -1082 206 -1070
rect 148 -1158 160 -1082
rect 194 -1158 206 -1082
rect 148 -1170 206 -1158
rect 236 -1082 294 -1070
rect 236 -1158 248 -1082
rect 282 -1158 294 -1082
rect 236 -1170 294 -1158
rect 324 -1082 382 -1070
rect 324 -1158 336 -1082
rect 370 -1158 382 -1082
rect 324 -1170 382 -1158
rect 412 -1082 470 -1070
rect 412 -1158 424 -1082
rect 458 -1158 470 -1082
rect 412 -1170 470 -1158
rect 500 -1082 558 -1070
rect 500 -1158 512 -1082
rect 546 -1158 558 -1082
rect 500 -1170 558 -1158
rect 588 -1082 646 -1070
rect 588 -1158 600 -1082
rect 634 -1158 646 -1082
rect 588 -1170 646 -1158
rect 676 -1082 734 -1070
rect 676 -1158 688 -1082
rect 722 -1158 734 -1082
rect 676 -1170 734 -1158
rect 764 -1082 822 -1070
rect 764 -1158 776 -1082
rect 810 -1158 822 -1082
rect 764 -1170 822 -1158
rect 852 -1082 910 -1070
rect 852 -1158 864 -1082
rect 898 -1158 910 -1082
rect 852 -1170 910 -1158
rect 1463 -1176 1475 -800
rect 1509 -1176 1525 -800
rect 1463 -1188 1525 -1176
rect 1555 -800 1617 -788
rect 1555 -1176 1567 -800
rect 1601 -1176 1617 -800
rect 1555 -1188 1617 -1176
rect 1647 -800 1713 -788
rect 1647 -1176 1663 -800
rect 1697 -1176 1713 -800
rect 1647 -1188 1713 -1176
rect 1743 -800 1809 -788
rect 1743 -1176 1759 -800
rect 1793 -1176 1809 -800
rect 1743 -1188 1809 -1176
rect 1839 -800 1905 -788
rect 1839 -1176 1855 -800
rect 1889 -1176 1905 -800
rect 1839 -1188 1905 -1176
rect 1935 -800 1997 -788
rect 1935 -1176 1951 -800
rect 1985 -1176 1997 -800
rect 1935 -1188 1997 -1176
rect 2027 -800 2089 -788
rect 2027 -1176 2043 -800
rect 2077 -1176 2089 -800
rect 2027 -1188 2089 -1176
<< pdiff >>
rect 1090 40 1148 52
rect -50 -255 12 -243
rect -50 -331 -38 -255
rect -4 -331 12 -255
rect -50 -343 12 -331
rect 42 -255 104 -243
rect 42 -331 54 -255
rect 88 -331 104 -255
rect 42 -343 104 -331
rect 134 -255 196 -243
rect 134 -331 148 -255
rect 182 -331 196 -255
rect 134 -343 196 -331
rect 226 -255 288 -243
rect 226 -331 240 -255
rect 274 -331 288 -255
rect 226 -343 288 -331
rect 318 -255 380 -243
rect 318 -331 332 -255
rect 366 -331 380 -255
rect 318 -343 380 -331
rect 410 -255 472 -243
rect 410 -331 424 -255
rect 458 -331 472 -255
rect 410 -343 472 -331
rect 502 -255 564 -243
rect 502 -331 516 -255
rect 550 -331 564 -255
rect 502 -343 564 -331
rect 594 -255 656 -243
rect 594 -331 608 -255
rect 642 -331 656 -255
rect 594 -343 656 -331
rect 686 -255 748 -243
rect 686 -331 700 -255
rect 734 -331 748 -255
rect 686 -343 748 -331
rect 778 -255 840 -243
rect 778 -331 794 -255
rect 828 -331 840 -255
rect 778 -343 840 -331
rect 870 -255 932 -243
rect 870 -331 886 -255
rect 920 -331 932 -255
rect 870 -343 932 -331
rect 1090 -336 1102 40
rect 1136 -336 1148 40
rect 1090 -348 1148 -336
rect 1178 40 1236 52
rect 1178 -336 1190 40
rect 1224 -336 1236 40
rect 1178 -348 1236 -336
rect 1266 40 1324 52
rect 1266 -336 1278 40
rect 1312 -336 1324 40
rect 1266 -348 1324 -336
rect 1354 40 1412 52
rect 1354 -336 1366 40
rect 1400 -336 1412 40
rect 1354 -348 1412 -336
rect 1442 40 1500 52
rect 1442 -336 1454 40
rect 1488 -336 1500 40
rect 1442 -348 1500 -336
rect 1530 40 1588 52
rect 1530 -336 1542 40
rect 1576 -336 1588 40
rect 1530 -348 1588 -336
rect 1618 40 1676 52
rect 1618 -336 1630 40
rect 1664 -336 1676 40
rect 1618 -348 1676 -336
rect 1877 40 1935 52
rect 1877 -336 1889 40
rect 1923 -336 1935 40
rect 1877 -348 1935 -336
rect 1965 40 2023 52
rect 1965 -336 1977 40
rect 2011 -336 2023 40
rect 1965 -348 2023 -336
rect 2053 40 2111 52
rect 2053 -336 2065 40
rect 2099 -336 2111 40
rect 2053 -348 2111 -336
rect 2141 40 2199 52
rect 2141 -336 2153 40
rect 2187 -336 2199 40
rect 2141 -348 2199 -336
rect 2229 40 2287 52
rect 2229 -336 2241 40
rect 2275 -336 2287 40
rect 2229 -348 2287 -336
rect 2317 40 2375 52
rect 2317 -336 2329 40
rect 2363 -336 2375 40
rect 2317 -348 2375 -336
rect 2405 40 2463 52
rect 2405 -336 2417 40
rect 2451 -336 2463 40
rect 2405 -348 2463 -336
<< ndiffc >>
rect -16 -961 18 -585
rect 72 -961 106 -585
rect 160 -961 194 -585
rect 248 -961 282 -585
rect 336 -961 370 -585
rect 424 -961 458 -585
rect 512 -961 546 -585
rect 600 -961 634 -585
rect 688 -961 722 -585
rect 776 -961 810 -585
rect 864 -961 898 -585
rect -16 -1158 18 -1082
rect 72 -1158 106 -1082
rect 160 -1158 194 -1082
rect 248 -1158 282 -1082
rect 336 -1158 370 -1082
rect 424 -1158 458 -1082
rect 512 -1158 546 -1082
rect 600 -1158 634 -1082
rect 688 -1158 722 -1082
rect 776 -1158 810 -1082
rect 864 -1158 898 -1082
rect 1475 -1176 1509 -800
rect 1567 -1176 1601 -800
rect 1663 -1176 1697 -800
rect 1759 -1176 1793 -800
rect 1855 -1176 1889 -800
rect 1951 -1176 1985 -800
rect 2043 -1176 2077 -800
<< pdiffc >>
rect -38 -331 -4 -255
rect 54 -331 88 -255
rect 148 -331 182 -255
rect 240 -331 274 -255
rect 332 -331 366 -255
rect 424 -331 458 -255
rect 516 -331 550 -255
rect 608 -331 642 -255
rect 700 -331 734 -255
rect 794 -331 828 -255
rect 886 -331 920 -255
rect 1102 -336 1136 40
rect 1190 -336 1224 40
rect 1278 -336 1312 40
rect 1366 -336 1400 40
rect 1454 -336 1488 40
rect 1542 -336 1576 40
rect 1630 -336 1664 40
rect 1889 -336 1923 40
rect 1977 -336 2011 40
rect 2065 -336 2099 40
rect 2153 -336 2187 40
rect 2241 -336 2275 40
rect 2329 -336 2363 40
rect 2417 -336 2451 40
<< psubdiff >>
rect -286 2162 -164 2188
rect -286 2088 -262 2162
rect -188 2088 -164 2162
rect -286 2064 -164 2088
rect 262 2162 384 2188
rect 262 2088 286 2162
rect 360 2088 384 2162
rect 262 2064 384 2088
rect 810 2162 932 2188
rect 810 2088 834 2162
rect 908 2088 932 2162
rect 810 2064 932 2088
rect 1358 2162 1480 2188
rect 1358 2088 1382 2162
rect 1456 2088 1480 2162
rect 1358 2064 1480 2088
rect 1906 2162 2028 2188
rect 1906 2088 1930 2162
rect 2004 2088 2028 2162
rect 1906 2064 2028 2088
rect 2436 2162 2558 2188
rect 2436 2088 2460 2162
rect 2534 2088 2558 2162
rect 2436 2064 2558 2088
rect 2984 2162 3106 2188
rect 2984 2088 3008 2162
rect 3082 2088 3106 2162
rect 2984 2064 3106 2088
rect 3534 2162 3656 2188
rect 3534 2088 3558 2162
rect 3632 2088 3656 2162
rect 3534 2064 3656 2088
rect -652 2020 -530 2046
rect -652 1946 -628 2020
rect -554 1946 -530 2020
rect -652 1922 -530 1946
rect 4353 1950 4475 1976
rect 4353 1876 4377 1950
rect 4451 1876 4475 1950
rect 4353 1852 4475 1876
rect -652 1546 -530 1572
rect -652 1472 -628 1546
rect -554 1472 -530 1546
rect -652 1448 -530 1472
rect 4353 1474 4475 1500
rect 4353 1400 4377 1474
rect 4451 1400 4475 1474
rect 4353 1376 4475 1400
rect -652 1072 -530 1098
rect -652 998 -628 1072
rect -554 998 -530 1072
rect -652 974 -530 998
rect 4353 1000 4475 1026
rect 4353 926 4377 1000
rect 4451 926 4475 1000
rect 4353 902 4475 926
rect -652 598 -530 624
rect -652 524 -628 598
rect -554 524 -530 598
rect -652 500 -530 524
rect 4351 526 4473 552
rect 4351 452 4375 526
rect 4449 452 4473 526
rect 4351 434 4473 452
rect -116 -642 -82 -569
rect 4351 -560 4473 -534
rect -116 -711 -82 -677
rect -116 -780 -82 -746
rect -116 -849 -82 -815
rect -116 -918 -82 -884
rect -116 -987 -82 -953
rect 964 -632 998 -569
rect 964 -701 998 -667
rect 964 -770 998 -736
rect 4351 -634 4375 -560
rect 4449 -634 4473 -560
rect 4351 -658 4473 -634
rect 964 -839 998 -805
rect 964 -908 998 -874
rect 964 -977 998 -943
rect -116 -1056 -82 -1022
rect 964 -1046 998 -1012
rect -116 -1125 -82 -1091
rect -116 -1194 -82 -1160
rect 964 -1115 998 -1081
rect -116 -1263 -82 -1229
rect 964 -1184 998 -1150
rect 964 -1253 998 -1219
rect -116 -1326 -82 -1298
rect 964 -1326 998 -1288
rect 1375 -843 1409 -809
rect 1375 -912 1409 -878
rect 1375 -981 1409 -947
rect 1375 -1050 1409 -1016
rect 1375 -1119 1409 -1085
rect 1375 -1188 1409 -1154
rect 2143 -843 2177 -809
rect 2143 -912 2177 -878
rect 2143 -981 2177 -947
rect 2143 -1050 2177 -1016
rect 2143 -1119 2177 -1085
rect 4351 -1034 4473 -1008
rect 4351 -1108 4375 -1034
rect 4449 -1108 4473 -1034
rect 4351 -1132 4473 -1108
rect 2143 -1188 2177 -1154
rect 1375 -1257 1409 -1223
rect 2143 -1257 2177 -1223
rect 1375 -1326 1409 -1292
rect 2143 -1326 2177 -1292
rect -116 -1332 1121 -1326
rect -116 -1368 100 -1332
rect 136 -1368 218 -1332
rect 254 -1368 336 -1332
rect 372 -1368 454 -1332
rect 490 -1368 572 -1332
rect 608 -1368 690 -1332
rect 726 -1368 808 -1332
rect 844 -1362 1121 -1332
rect 1157 -1362 1213 -1326
rect 1249 -1362 1305 -1326
rect 1341 -1362 1397 -1326
rect 1433 -1362 1489 -1326
rect 1525 -1362 1581 -1326
rect 1617 -1362 1673 -1326
rect 1709 -1362 1769 -1326
rect 1805 -1362 1857 -1326
rect 1893 -1362 1949 -1326
rect 1985 -1362 2041 -1326
rect 2077 -1362 2133 -1326
rect 2169 -1362 2193 -1326
rect 844 -1368 2193 -1362
rect -116 -1372 2193 -1368
rect -646 -1740 -524 -1714
rect -646 -1814 -622 -1740
rect -548 -1814 -524 -1740
rect -646 -1838 -524 -1814
rect 4351 -1770 4473 -1744
rect 4351 -1844 4375 -1770
rect 4449 -1844 4473 -1770
rect 4351 -1868 4473 -1844
rect -646 -2214 -524 -2188
rect -646 -2288 -622 -2214
rect -548 -2288 -524 -2214
rect -646 -2312 -524 -2288
rect 4351 -2244 4473 -2218
rect 4351 -2318 4375 -2244
rect 4449 -2318 4473 -2244
rect 4351 -2342 4473 -2318
rect -646 -2688 -524 -2662
rect -646 -2762 -622 -2688
rect -548 -2762 -524 -2688
rect -646 -2786 -524 -2762
rect 4351 -2718 4473 -2692
rect 4351 -2792 4375 -2718
rect 4449 -2792 4473 -2718
rect 4351 -2816 4473 -2792
rect -116 -3248 6 -3222
rect -116 -3322 -92 -3248
rect -18 -3322 6 -3248
rect -116 -3346 6 -3322
rect 432 -3248 554 -3222
rect 432 -3322 456 -3248
rect 530 -3322 554 -3248
rect 432 -3346 554 -3322
rect 980 -3248 1102 -3222
rect 980 -3322 1004 -3248
rect 1078 -3322 1102 -3248
rect 980 -3346 1102 -3322
rect 1528 -3248 1650 -3222
rect 1528 -3322 1552 -3248
rect 1626 -3322 1650 -3248
rect 1528 -3346 1650 -3322
rect 2076 -3248 2198 -3222
rect 2076 -3322 2100 -3248
rect 2174 -3322 2198 -3248
rect 2076 -3346 2198 -3322
rect 2624 -3248 2746 -3222
rect 2624 -3322 2648 -3248
rect 2722 -3322 2746 -3248
rect 2624 -3346 2746 -3322
rect 3174 -3248 3296 -3222
rect 3174 -3322 3198 -3248
rect 3272 -3322 3296 -3248
rect 3174 -3346 3296 -3322
<< nsubdiff >>
rect 935 226 3068 234
rect 935 210 1084 226
rect 935 176 939 210
rect 974 192 1084 210
rect 1118 192 1168 226
rect 1202 192 1252 226
rect 1286 192 1336 226
rect 1370 192 1420 226
rect 1454 192 1504 226
rect 1538 192 1588 226
rect 1622 192 1672 226
rect 1706 192 1840 226
rect 1874 192 1924 226
rect 1958 192 2008 226
rect 2042 192 2080 226
rect 2114 192 2164 226
rect 2198 192 2248 226
rect 2282 192 2320 226
rect 2354 192 2404 226
rect 2438 192 2476 226
rect 2510 192 2632 226
rect 2666 192 3068 226
rect 974 186 3068 192
rect 974 176 980 186
rect 935 127 980 176
rect 935 93 939 127
rect 974 93 980 127
rect 935 44 980 93
rect 1753 127 1799 186
rect 1753 93 1759 127
rect 1793 93 1799 127
rect 935 10 939 44
rect 974 10 980 44
rect 935 -39 980 10
rect 935 -73 939 -39
rect 974 -73 980 -39
rect 935 -122 980 -73
rect -640 -130 980 -122
rect -640 -164 -600 -130
rect -566 -164 -444 -130
rect -410 -164 -290 -130
rect -256 -164 -146 -130
rect -112 -164 -32 -130
rect 2 -164 82 -130
rect 116 -164 166 -130
rect 200 -164 250 -130
rect 284 -164 334 -130
rect 368 -164 418 -130
rect 452 -164 502 -130
rect 536 -164 586 -130
rect 620 -164 670 -130
rect 704 -164 754 -130
rect 788 -164 838 -130
rect 872 -164 922 -130
rect 956 -164 980 -130
rect -640 -177 980 -164
rect 1753 44 1799 93
rect 2573 127 2619 186
rect 2573 93 2579 127
rect 2613 93 2619 127
rect 1753 10 1759 44
rect 1793 10 1799 44
rect 1753 -39 1799 10
rect 1753 -73 1759 -39
rect 1793 -73 1799 -39
rect 1753 -127 1799 -73
rect 1753 -161 1759 -127
rect 1793 -161 1799 -127
rect 1753 -210 1799 -161
rect 1753 -244 1759 -210
rect 1793 -244 1799 -210
rect 1753 -293 1799 -244
rect 1753 -327 1759 -293
rect 1793 -327 1799 -293
rect 1753 -370 1799 -327
rect 2573 44 2619 93
rect 2573 10 2579 44
rect 2613 10 2619 44
rect 2573 -39 2619 10
rect 2573 -73 2579 -39
rect 2613 -73 2619 -39
rect 2573 -122 2619 -73
rect 2573 -156 2579 -122
rect 2613 -156 2619 -122
rect 2573 -191 2619 -156
rect 3180 -1276 3204 -1238
rect 3242 -1276 3280 -1238
rect 3318 -1276 3356 -1238
rect 3394 -1276 3432 -1238
rect 3470 -1276 3508 -1238
rect 3546 -1276 3584 -1238
rect 3622 -1276 3660 -1238
rect 3698 -1276 3736 -1238
rect 3774 -1276 3830 -1238
<< psubdiffcont >>
rect -262 2088 -188 2162
rect 286 2088 360 2162
rect 834 2088 908 2162
rect 1382 2088 1456 2162
rect 1930 2088 2004 2162
rect 2460 2088 2534 2162
rect 3008 2088 3082 2162
rect 3558 2088 3632 2162
rect -628 1946 -554 2020
rect 4377 1876 4451 1950
rect -628 1472 -554 1546
rect 4377 1400 4451 1474
rect -628 998 -554 1072
rect 4377 926 4451 1000
rect -628 524 -554 598
rect 4375 452 4449 526
rect -116 -677 -82 -642
rect -116 -746 -82 -711
rect -116 -815 -82 -780
rect -116 -884 -82 -849
rect -116 -953 -82 -918
rect 964 -667 998 -632
rect 964 -736 998 -701
rect 964 -805 998 -770
rect 4375 -634 4449 -560
rect 964 -874 998 -839
rect 964 -943 998 -908
rect -116 -1022 -82 -987
rect 964 -1012 998 -977
rect -116 -1091 -82 -1056
rect -116 -1160 -82 -1125
rect 964 -1081 998 -1046
rect 964 -1150 998 -1115
rect -116 -1229 -82 -1194
rect -116 -1298 -82 -1263
rect 964 -1219 998 -1184
rect 964 -1288 998 -1253
rect 1375 -878 1409 -843
rect 1375 -947 1409 -912
rect 1375 -1016 1409 -981
rect 1375 -1085 1409 -1050
rect 1375 -1154 1409 -1119
rect 2143 -878 2177 -843
rect 2143 -947 2177 -912
rect 2143 -1016 2177 -981
rect 2143 -1085 2177 -1050
rect 2143 -1154 2177 -1119
rect 4375 -1108 4449 -1034
rect 1375 -1223 1409 -1188
rect 2143 -1223 2177 -1188
rect 1375 -1292 1409 -1257
rect 2143 -1292 2177 -1257
rect 100 -1368 136 -1332
rect 218 -1368 254 -1332
rect 336 -1368 372 -1332
rect 454 -1368 490 -1332
rect 572 -1368 608 -1332
rect 690 -1368 726 -1332
rect 808 -1368 844 -1332
rect 1121 -1362 1157 -1326
rect 1213 -1362 1249 -1326
rect 1305 -1362 1341 -1326
rect 1397 -1362 1433 -1326
rect 1489 -1362 1525 -1326
rect 1581 -1362 1617 -1326
rect 1673 -1362 1709 -1326
rect 1769 -1362 1805 -1326
rect 1857 -1362 1893 -1326
rect 1949 -1362 1985 -1326
rect 2041 -1362 2077 -1326
rect 2133 -1362 2169 -1326
rect -622 -1814 -548 -1740
rect 4375 -1844 4449 -1770
rect -622 -2288 -548 -2214
rect 4375 -2318 4449 -2244
rect -622 -2762 -548 -2688
rect 4375 -2792 4449 -2718
rect -92 -3322 -18 -3248
rect 456 -3322 530 -3248
rect 1004 -3322 1078 -3248
rect 1552 -3322 1626 -3248
rect 2100 -3322 2174 -3248
rect 2648 -3322 2722 -3248
rect 3198 -3322 3272 -3248
<< nsubdiffcont >>
rect 939 176 974 210
rect 1084 192 1118 226
rect 1168 192 1202 226
rect 1252 192 1286 226
rect 1336 192 1370 226
rect 1420 192 1454 226
rect 1504 192 1538 226
rect 1588 192 1622 226
rect 1672 192 1706 226
rect 1840 192 1874 226
rect 1924 192 1958 226
rect 2008 192 2042 226
rect 2080 192 2114 226
rect 2164 192 2198 226
rect 2248 192 2282 226
rect 2320 192 2354 226
rect 2404 192 2438 226
rect 2476 192 2510 226
rect 2632 192 2666 226
rect 939 93 974 127
rect 1759 93 1793 127
rect 939 10 974 44
rect 939 -73 974 -39
rect -600 -164 -566 -130
rect -444 -164 -410 -130
rect -290 -164 -256 -130
rect -146 -164 -112 -130
rect -32 -164 2 -130
rect 82 -164 116 -130
rect 166 -164 200 -130
rect 250 -164 284 -130
rect 334 -164 368 -130
rect 418 -164 452 -130
rect 502 -164 536 -130
rect 586 -164 620 -130
rect 670 -164 704 -130
rect 754 -164 788 -130
rect 838 -164 872 -130
rect 922 -164 956 -130
rect 2579 93 2613 127
rect 1759 10 1793 44
rect 1759 -73 1793 -39
rect 1759 -161 1793 -127
rect 1759 -244 1793 -210
rect 1759 -327 1793 -293
rect 2579 10 2613 44
rect 2579 -73 2613 -39
rect 2579 -156 2613 -122
rect 2787 -1276 2825 -1238
rect 2863 -1276 2901 -1238
rect 2939 -1276 2977 -1238
rect 3015 -1276 3053 -1238
rect 3204 -1276 3242 -1238
rect 3280 -1276 3318 -1238
rect 3356 -1276 3394 -1238
rect 3432 -1276 3470 -1238
rect 3508 -1276 3546 -1238
rect 3584 -1276 3622 -1238
rect 3660 -1276 3698 -1238
rect 3736 -1276 3774 -1238
<< poly >>
rect 1148 52 1178 78
rect 1236 52 1266 78
rect 1324 52 1354 78
rect 1412 52 1442 78
rect 1500 52 1530 78
rect 1588 52 1618 78
rect 12 -243 42 -217
rect 104 -243 134 -217
rect 196 -243 226 -217
rect 288 -243 318 -217
rect 380 -243 410 -217
rect 472 -243 502 -217
rect 564 -243 594 -217
rect 656 -243 686 -217
rect 748 -243 778 -217
rect 840 -243 870 -217
rect 12 -369 42 -343
rect 104 -369 134 -343
rect 196 -369 226 -343
rect 288 -369 318 -343
rect 380 -369 410 -343
rect 12 -390 410 -369
rect 12 -430 22 -390
rect 69 -399 410 -390
rect 472 -369 502 -343
rect 564 -369 594 -343
rect 656 -369 686 -343
rect 748 -369 778 -343
rect 840 -369 870 -343
rect 1935 52 1965 78
rect 2023 52 2053 78
rect 2111 52 2141 78
rect 2199 52 2229 78
rect 2287 52 2317 78
rect 2375 52 2405 78
rect 472 -390 870 -369
rect 472 -399 807 -390
rect 69 -430 80 -399
rect 12 -446 80 -430
rect 797 -430 807 -399
rect 854 -399 870 -390
rect 1148 -374 1178 -348
rect 1236 -374 1266 -348
rect 1324 -374 1354 -348
rect 854 -430 865 -399
rect 1148 -402 1354 -374
rect 1148 -404 1190 -402
rect 797 -446 865 -430
rect 1174 -436 1190 -404
rect 1226 -404 1354 -402
rect 1412 -374 1442 -348
rect 1500 -374 1530 -348
rect 1588 -374 1618 -348
rect 1412 -404 1618 -374
rect 1226 -436 1244 -404
rect 1174 -446 1244 -436
rect 1530 -413 1618 -404
rect 1530 -447 1544 -413
rect 1606 -447 1618 -413
rect 1530 -463 1618 -447
rect 1935 -374 1965 -348
rect 2023 -374 2053 -348
rect 2111 -374 2141 -348
rect 1935 -404 2141 -374
rect 2199 -374 2229 -348
rect 2287 -370 2317 -348
rect 2375 -370 2405 -348
rect 2287 -374 2405 -370
rect 2199 -402 2405 -374
rect 2199 -404 2329 -402
rect 1935 -413 2023 -404
rect 1935 -447 1949 -413
rect 2011 -447 2023 -413
rect 2313 -436 2329 -404
rect 2363 -404 2405 -402
rect 2363 -436 2379 -404
rect 2313 -446 2379 -436
rect 1935 -463 2023 -447
rect 180 -492 260 -482
rect 180 -516 196 -492
rect 30 -526 196 -516
rect 244 -516 260 -492
rect 622 -490 702 -480
rect 622 -514 638 -490
rect 244 -526 412 -516
rect 30 -547 412 -526
rect 30 -573 60 -547
rect 118 -573 148 -547
rect 206 -573 236 -547
rect 294 -573 324 -547
rect 382 -573 412 -547
rect 470 -524 638 -514
rect 686 -514 702 -490
rect 686 -524 852 -514
rect 470 -545 852 -524
rect 470 -573 500 -545
rect 558 -573 588 -545
rect 646 -573 676 -545
rect 734 -573 764 -545
rect 822 -573 852 -545
rect 1649 -652 1743 -624
rect 1649 -705 1670 -652
rect 1718 -705 1743 -652
rect 1649 -719 1743 -705
rect 1525 -788 1555 -762
rect 1617 -788 1647 -762
rect 1713 -788 1743 -719
rect 1809 -652 1903 -624
rect 1809 -706 1836 -652
rect 1884 -706 1903 -652
rect 1809 -719 1903 -706
rect 1809 -788 1839 -719
rect 1905 -788 1935 -762
rect 1997 -788 2027 -762
rect 30 -1001 60 -973
rect 118 -1001 148 -973
rect 206 -1001 236 -973
rect 294 -1001 324 -973
rect 382 -1001 412 -973
rect 470 -1001 500 -973
rect 558 -1001 588 -973
rect 646 -1001 676 -973
rect 734 -1001 764 -973
rect 822 -1001 852 -973
rect 30 -1070 60 -1044
rect 118 -1070 148 -1044
rect 206 -1070 236 -1044
rect 294 -1070 324 -1044
rect 382 -1070 412 -1044
rect 470 -1070 500 -1044
rect 558 -1070 588 -1044
rect 646 -1070 676 -1044
rect 734 -1070 764 -1044
rect 822 -1070 852 -1044
rect 30 -1196 60 -1170
rect 118 -1196 148 -1170
rect 30 -1238 148 -1196
rect 30 -1272 68 -1238
rect 110 -1272 148 -1238
rect 30 -1298 148 -1272
rect 206 -1196 236 -1170
rect 294 -1196 324 -1170
rect 206 -1238 324 -1196
rect 206 -1272 244 -1238
rect 286 -1272 324 -1238
rect 206 -1298 324 -1272
rect 382 -1196 412 -1170
rect 470 -1196 500 -1170
rect 382 -1238 500 -1196
rect 382 -1272 420 -1238
rect 462 -1272 500 -1238
rect 382 -1298 500 -1272
rect 558 -1196 588 -1170
rect 646 -1196 676 -1170
rect 558 -1238 676 -1196
rect 558 -1272 596 -1238
rect 638 -1272 676 -1238
rect 558 -1298 676 -1272
rect 734 -1196 764 -1170
rect 822 -1196 852 -1170
rect 734 -1238 852 -1196
rect 734 -1272 772 -1238
rect 814 -1272 852 -1238
rect 734 -1298 852 -1272
rect 1525 -1227 1555 -1188
rect 1617 -1226 1647 -1188
rect 1713 -1214 1743 -1188
rect 1809 -1214 1839 -1188
rect 1905 -1226 1935 -1188
rect 1997 -1226 2027 -1188
rect 1462 -1237 1555 -1227
rect 1462 -1279 1478 -1237
rect 1539 -1279 1555 -1237
rect 1462 -1290 1555 -1279
rect 1611 -1242 1671 -1226
rect 1611 -1276 1621 -1242
rect 1655 -1276 1671 -1242
rect 1611 -1292 1671 -1276
rect 1883 -1242 1943 -1226
rect 1883 -1276 1893 -1242
rect 1927 -1276 1943 -1242
rect 1883 -1292 1943 -1276
rect 1997 -1236 2090 -1226
rect 1997 -1278 2013 -1236
rect 2074 -1278 2090 -1236
rect 1997 -1289 2090 -1278
<< polycont >>
rect 22 -430 69 -390
rect 807 -430 854 -390
rect 1190 -436 1226 -402
rect 1544 -447 1606 -413
rect 1949 -447 2011 -413
rect 2329 -436 2363 -402
rect 196 -526 244 -492
rect 638 -524 686 -490
rect 1670 -705 1718 -652
rect 1836 -706 1884 -652
rect 68 -1272 110 -1238
rect 244 -1272 286 -1238
rect 420 -1272 462 -1238
rect 596 -1272 638 -1238
rect 772 -1272 814 -1238
rect 1478 -1279 1539 -1237
rect 1621 -1276 1655 -1242
rect 1893 -1276 1927 -1242
rect 2013 -1278 2074 -1236
<< locali >>
rect -686 2162 4515 2218
rect -686 2088 -262 2162
rect -188 2088 286 2162
rect 360 2088 834 2162
rect 908 2088 1382 2162
rect 1456 2088 1930 2162
rect 2004 2088 2460 2162
rect 2534 2088 3008 2162
rect 3082 2088 3558 2162
rect 3632 2088 4515 2162
rect -686 2020 4515 2088
rect -686 1970 -628 2020
rect -554 1970 -450 2020
rect 200 2000 660 2020
rect 2780 2000 3240 2020
rect -686 1570 -650 1970
rect -520 1570 -450 1970
rect -686 1546 -450 1570
rect -686 1472 -628 1546
rect -554 1530 -450 1546
rect 4317 1950 4515 2020
rect 4317 1876 4377 1950
rect 4451 1876 4515 1950
rect -554 1472 -488 1530
rect -686 1430 -488 1472
rect -686 990 -666 1430
rect -530 990 -488 1430
rect 4317 1474 4515 1876
rect 4317 1400 4377 1474
rect 4451 1400 4515 1474
rect -686 870 -488 990
rect -686 440 -666 870
rect -510 440 -488 870
rect -686 420 -488 440
rect 4317 1000 4515 1400
rect 4317 926 4377 1000
rect 4451 926 4515 1000
rect 4317 526 4515 926
rect 4317 452 4375 526
rect 4449 452 4515 526
rect 935 227 4179 234
rect 935 226 3299 227
rect 935 210 1084 226
rect 935 176 939 210
rect 974 192 1084 210
rect 1118 192 1168 226
rect 1202 192 1252 226
rect 1286 192 1336 226
rect 1370 192 1420 226
rect 1454 192 1504 226
rect 1538 192 1588 226
rect 1622 192 1672 226
rect 1706 192 1840 226
rect 1874 192 1924 226
rect 1958 192 2008 226
rect 2042 192 2080 226
rect 2114 192 2164 226
rect 2198 192 2248 226
rect 2282 192 2320 226
rect 2354 192 2404 226
rect 2438 192 2476 226
rect 2510 192 2632 226
rect 2666 192 2716 226
rect 2750 192 2788 226
rect 2822 192 2917 226
rect 2951 192 2989 226
rect 3023 193 3299 226
rect 3333 193 3371 227
rect 3405 193 3443 227
rect 3477 193 3515 227
rect 3549 193 3587 227
rect 3621 193 3659 227
rect 3693 193 3732 227
rect 3766 193 3804 227
rect 3838 193 3876 227
rect 3910 193 3948 227
rect 3982 193 4020 227
rect 4054 193 4092 227
rect 4126 193 4179 227
rect 3023 192 4179 193
rect 974 186 4179 192
rect 974 176 980 186
rect 935 127 980 176
rect 935 93 939 127
rect 974 93 980 127
rect 935 44 980 93
rect 1753 127 1799 186
rect 1753 93 1759 127
rect 1793 93 1799 127
rect 935 10 939 44
rect 974 10 980 44
rect 935 -39 980 10
rect 935 -73 939 -39
rect 974 -73 980 -39
rect 935 -122 980 -73
rect -640 -130 980 -122
rect -640 -164 -600 -130
rect -566 -164 -444 -130
rect -410 -164 -290 -130
rect -256 -164 -146 -130
rect -112 -164 -32 -130
rect 2 -164 82 -130
rect 116 -164 166 -130
rect 200 -164 250 -130
rect 284 -164 334 -130
rect 368 -164 418 -130
rect 452 -164 502 -130
rect 536 -164 586 -130
rect 620 -164 670 -130
rect 704 -164 754 -130
rect 788 -164 838 -130
rect 872 -164 922 -130
rect 956 -164 980 -130
rect -640 -177 980 -164
rect 1102 40 1136 56
rect -38 -255 -4 -239
rect -38 -347 -4 -331
rect 54 -255 88 -239
rect 54 -347 88 -331
rect 148 -255 182 -239
rect 148 -347 182 -331
rect 240 -255 274 -239
rect 240 -347 274 -331
rect 332 -255 366 -239
rect 332 -347 366 -331
rect 424 -255 458 -239
rect 424 -347 458 -331
rect 516 -255 550 -239
rect 516 -347 550 -331
rect 608 -255 642 -239
rect 608 -347 642 -331
rect 700 -255 734 -239
rect 700 -347 734 -331
rect 794 -255 828 -239
rect 794 -347 828 -331
rect 886 -255 920 -239
rect 886 -347 920 -331
rect 1102 -352 1136 -336
rect 1190 40 1224 56
rect 1190 -352 1224 -336
rect 1278 40 1312 56
rect 1278 -352 1312 -336
rect 1366 40 1400 56
rect 1366 -352 1400 -336
rect 1454 40 1488 56
rect 1454 -352 1488 -336
rect 1542 40 1576 56
rect 1542 -352 1576 -336
rect 1630 40 1664 56
rect 1630 -352 1664 -336
rect 1753 44 1799 93
rect 2573 127 2619 186
rect 2573 93 2579 127
rect 2613 93 2619 127
rect 1753 10 1759 44
rect 1793 10 1799 44
rect 1753 -39 1799 10
rect 1753 -73 1759 -39
rect 1793 -73 1799 -39
rect 1753 -127 1799 -73
rect 1753 -161 1759 -127
rect 1793 -161 1799 -127
rect 1753 -210 1799 -161
rect 1753 -244 1759 -210
rect 1793 -244 1799 -210
rect 1753 -293 1799 -244
rect 1753 -327 1759 -293
rect 1793 -327 1799 -293
rect 6 -390 85 -389
rect 6 -430 22 -390
rect 69 -430 85 -390
rect 791 -430 807 -390
rect 854 -430 870 -390
rect 1174 -402 1244 -386
rect 6 -431 85 -430
rect 1174 -436 1190 -402
rect 1226 -436 1244 -402
rect 1174 -446 1244 -436
rect 1530 -413 1618 -397
rect 1753 -413 1799 -327
rect 1889 40 1923 56
rect 1889 -352 1923 -336
rect 1977 40 2011 56
rect 1977 -352 2011 -336
rect 2065 40 2099 56
rect 2065 -352 2099 -336
rect 2153 40 2187 56
rect 2153 -352 2187 -336
rect 2241 40 2275 56
rect 2241 -352 2275 -336
rect 2329 40 2363 56
rect 2329 -352 2363 -336
rect 2417 40 2451 56
rect 2573 44 2619 93
rect 2573 10 2579 44
rect 2613 10 2619 44
rect 2573 -39 2619 10
rect 2573 -73 2579 -39
rect 2613 -73 2619 -39
rect 2573 -122 2619 -73
rect 2573 -156 2579 -122
rect 2613 -156 2619 -122
rect 2573 -191 2619 -156
rect 2417 -352 2451 -336
rect 3429 -349 3803 -314
rect 3429 -350 3633 -349
rect 1935 -413 2023 -397
rect 1182 -448 1226 -446
rect 1530 -447 1544 -413
rect 1606 -447 1618 -413
rect 1530 -463 1618 -447
rect 1935 -447 1949 -413
rect 2011 -447 2023 -413
rect 2313 -402 2379 -386
rect 2313 -436 2329 -402
rect 2363 -436 2379 -402
rect 3429 -401 3463 -350
rect 3497 -401 3549 -350
rect 3583 -400 3633 -350
rect 3667 -350 3803 -349
rect 3667 -400 3717 -350
rect 3583 -401 3717 -400
rect 3751 -401 3803 -350
rect 3429 -436 3803 -401
rect 2313 -446 2379 -436
rect 1935 -463 2023 -447
rect 2325 -448 2367 -446
rect 180 -492 260 -482
rect 180 -526 196 -492
rect 244 -526 260 -492
rect 180 -533 260 -526
rect 622 -490 702 -480
rect 622 -524 638 -490
rect 686 -524 702 -490
rect 622 -531 702 -524
rect 2695 -500 3119 -462
rect 2695 -501 2806 -500
rect 2695 -552 2721 -501
rect 2755 -551 2806 -501
rect 2840 -501 2978 -500
rect 2840 -551 2890 -501
rect 2755 -552 2890 -551
rect 2924 -551 2978 -501
rect 3012 -551 3061 -500
rect 3095 -551 3119 -500
rect 2924 -552 3119 -551
rect -116 -642 -74 -569
rect -82 -677 -74 -642
rect -116 -711 -74 -677
rect -82 -746 -74 -711
rect -116 -780 -74 -746
rect -82 -815 -74 -780
rect -116 -849 -74 -815
rect -82 -884 -74 -849
rect -116 -918 -74 -884
rect -82 -953 -74 -918
rect -116 -987 -74 -953
rect -16 -585 18 -569
rect -16 -977 18 -961
rect 72 -585 106 -569
rect 72 -977 106 -961
rect 160 -585 194 -568
rect 160 -977 194 -961
rect 248 -585 282 -569
rect 248 -977 282 -961
rect 336 -585 370 -568
rect 424 -585 458 -569
rect 512 -585 546 -568
rect 336 -977 370 -961
rect 424 -977 458 -961
rect 512 -977 546 -961
rect 600 -585 634 -569
rect 600 -977 634 -961
rect 688 -585 722 -568
rect 688 -977 722 -961
rect 776 -585 810 -569
rect 776 -977 810 -961
rect 864 -585 898 -569
rect 864 -977 898 -961
rect 956 -632 998 -569
rect 2695 -590 3119 -552
rect 4317 -560 4515 452
rect 956 -667 964 -632
rect 4317 -634 4375 -560
rect 4449 -634 4515 -560
rect 956 -701 998 -667
rect 956 -736 964 -701
rect 1654 -707 1670 -652
rect 1718 -707 1734 -652
rect 1820 -707 1836 -652
rect 1884 -707 1900 -652
rect 956 -770 998 -736
rect 956 -805 964 -770
rect 956 -839 998 -805
rect 1475 -800 1509 -784
rect 956 -874 964 -839
rect 956 -908 998 -874
rect 956 -943 964 -908
rect 956 -977 998 -943
rect -82 -1022 -74 -987
rect -116 -1056 -74 -1022
rect -82 -1091 -74 -1056
rect 956 -1012 964 -977
rect 956 -1046 998 -1012
rect -116 -1125 -74 -1091
rect -82 -1160 -74 -1125
rect -116 -1194 -74 -1160
rect -16 -1082 18 -1064
rect -16 -1174 18 -1158
rect 72 -1082 106 -1064
rect 72 -1174 106 -1158
rect 160 -1082 194 -1064
rect -82 -1229 -74 -1194
rect -116 -1263 -74 -1229
rect -82 -1298 -74 -1263
rect 52 -1237 126 -1226
rect 52 -1272 68 -1237
rect 110 -1272 126 -1237
rect 52 -1282 126 -1272
rect -116 -1316 -74 -1298
rect 160 -1316 194 -1158
rect 248 -1082 282 -1064
rect 248 -1174 282 -1158
rect 336 -1082 370 -1064
rect 228 -1237 302 -1226
rect 228 -1272 244 -1237
rect 286 -1272 302 -1237
rect 228 -1282 302 -1272
rect 336 -1316 370 -1158
rect 424 -1082 458 -1064
rect 424 -1174 458 -1158
rect 512 -1082 546 -1064
rect 404 -1237 478 -1226
rect 404 -1272 420 -1237
rect 462 -1272 478 -1237
rect 404 -1282 478 -1272
rect 512 -1316 546 -1158
rect 600 -1082 634 -1064
rect 600 -1174 634 -1158
rect 688 -1082 722 -1064
rect 580 -1237 654 -1226
rect 580 -1272 596 -1237
rect 638 -1272 654 -1237
rect 580 -1282 654 -1272
rect 688 -1316 722 -1158
rect 776 -1082 810 -1064
rect 776 -1174 810 -1158
rect 864 -1082 898 -1064
rect 864 -1174 898 -1158
rect 956 -1081 964 -1046
rect 956 -1115 998 -1081
rect 956 -1150 964 -1115
rect 956 -1184 998 -1150
rect 956 -1219 964 -1184
rect 756 -1237 830 -1226
rect 756 -1272 772 -1237
rect 814 -1272 830 -1237
rect 756 -1282 830 -1272
rect 956 -1253 998 -1219
rect 956 -1288 964 -1253
rect 956 -1316 998 -1288
rect 1375 -843 1417 -809
rect 1409 -878 1417 -843
rect 1375 -912 1417 -878
rect 1409 -947 1417 -912
rect 1375 -981 1417 -947
rect 1409 -1016 1417 -981
rect 1375 -1050 1417 -1016
rect 1409 -1085 1417 -1050
rect 1375 -1119 1417 -1085
rect 1409 -1154 1417 -1119
rect 1375 -1188 1417 -1154
rect 1409 -1223 1417 -1188
rect 1475 -1192 1509 -1176
rect 1567 -800 1601 -784
rect 1567 -1192 1601 -1176
rect 1663 -800 1697 -784
rect 1663 -1192 1697 -1176
rect 1759 -800 1793 -784
rect 1759 -1192 1793 -1176
rect 1855 -800 1889 -784
rect 1855 -1192 1889 -1176
rect 1951 -800 1985 -784
rect 1951 -1192 1985 -1176
rect 2043 -800 2077 -784
rect 2043 -1192 2077 -1176
rect 2135 -843 2177 -809
rect 2135 -878 2143 -843
rect 2135 -912 2177 -878
rect 2135 -947 2143 -912
rect 2135 -981 2177 -947
rect 2135 -1016 2143 -981
rect 2135 -1050 2177 -1016
rect 2135 -1085 2143 -1050
rect 2135 -1119 2177 -1085
rect 2135 -1154 2143 -1119
rect 2135 -1188 2177 -1154
rect 1375 -1257 1417 -1223
rect 2135 -1223 2143 -1188
rect 1409 -1292 1417 -1257
rect 1375 -1316 1417 -1292
rect -116 -1326 1417 -1316
rect 1462 -1237 1555 -1227
rect 1462 -1279 1478 -1237
rect 1539 -1279 1555 -1237
rect 1462 -1326 1555 -1279
rect 1611 -1232 1697 -1226
rect 1611 -1242 1649 -1232
rect 1611 -1276 1621 -1242
rect 1611 -1278 1649 -1276
rect 1683 -1278 1697 -1232
rect 1611 -1292 1697 -1278
rect 1857 -1232 1943 -1226
rect 1857 -1278 1871 -1232
rect 1905 -1242 1943 -1232
rect 1927 -1276 1943 -1242
rect 1905 -1278 1943 -1276
rect 1857 -1292 1943 -1278
rect 1997 -1236 2090 -1226
rect 1997 -1278 2013 -1236
rect 2074 -1278 2090 -1236
rect 1997 -1326 2090 -1278
rect 2135 -1257 2177 -1223
rect 4317 -1034 4515 -634
rect 4317 -1108 4375 -1034
rect 4449 -1108 4515 -1034
rect 4317 -1222 4515 -1108
rect 2135 -1292 2143 -1257
rect 3104 -1276 3204 -1238
rect 3242 -1276 3280 -1238
rect 3318 -1276 3356 -1238
rect 3394 -1276 3432 -1238
rect 3470 -1276 3508 -1238
rect 3546 -1276 3584 -1238
rect 3622 -1276 3660 -1238
rect 3698 -1276 3736 -1238
rect 3774 -1276 3830 -1238
rect 4317 -1256 4331 -1222
rect 4365 -1256 4403 -1222
rect 4437 -1256 4475 -1222
rect 4509 -1256 4515 -1222
rect 2135 -1311 2177 -1292
rect 4317 -1294 4515 -1256
rect 2135 -1326 3240 -1311
rect -686 -1366 -488 -1326
rect -686 -1400 -670 -1366
rect -636 -1400 -598 -1366
rect -564 -1400 -526 -1366
rect -492 -1400 -488 -1366
rect -116 -1332 1121 -1326
rect -116 -1368 100 -1332
rect 136 -1368 218 -1332
rect 254 -1368 336 -1332
rect 372 -1368 454 -1332
rect 490 -1368 572 -1332
rect 608 -1368 690 -1332
rect 726 -1368 808 -1332
rect 844 -1368 1121 -1332
rect -116 -1376 1121 -1368
rect 1157 -1376 1213 -1326
rect 1249 -1376 1305 -1326
rect 1341 -1376 1397 -1326
rect 1433 -1376 1489 -1326
rect 1525 -1376 1581 -1326
rect 1617 -1376 1673 -1326
rect 1709 -1376 1769 -1326
rect 1805 -1376 1857 -1326
rect 1893 -1376 1949 -1326
rect 1985 -1376 2041 -1326
rect 2077 -1376 2133 -1326
rect 2169 -1344 3240 -1326
rect 2169 -1376 2286 -1344
rect -116 -1380 2286 -1376
rect 2322 -1380 2360 -1344
rect 2396 -1380 2440 -1344
rect 2476 -1380 2520 -1344
rect 2556 -1380 2595 -1344
rect 2631 -1380 2669 -1344
rect 2705 -1380 2749 -1344
rect 2785 -1380 2829 -1344
rect 2865 -1380 2903 -1344
rect 2939 -1380 2983 -1344
rect 3019 -1380 3063 -1344
rect 3099 -1380 3143 -1344
rect 3179 -1380 3240 -1344
rect -116 -1395 3240 -1380
rect -686 -1438 -488 -1400
rect -686 -1472 -670 -1438
rect -636 -1472 -598 -1438
rect -564 -1472 -526 -1438
rect -492 -1472 -488 -1438
rect -686 -1510 -488 -1472
rect -686 -1544 -672 -1510
rect -638 -1544 -600 -1510
rect -566 -1544 -528 -1510
rect -494 -1544 -488 -1510
rect -686 -1610 -488 -1544
rect 200 -1590 660 -1395
rect 2278 -1396 3240 -1395
rect 2780 -1590 3240 -1396
rect 4317 -1328 4331 -1294
rect 4365 -1328 4403 -1294
rect 4437 -1328 4475 -1294
rect 4509 -1328 4515 -1294
rect 4317 -1366 4515 -1328
rect 4317 -1400 4331 -1366
rect 4365 -1400 4403 -1366
rect 4437 -1400 4475 -1366
rect 4509 -1400 4515 -1366
rect 4317 -1438 4515 -1400
rect 4317 -1472 4331 -1438
rect 4365 -1472 4403 -1438
rect 4437 -1472 4475 -1438
rect 4509 -1472 4515 -1438
rect 4317 -1510 4515 -1472
rect 4317 -1544 4331 -1510
rect 4365 -1544 4403 -1510
rect 4437 -1544 4475 -1510
rect 4509 -1544 4515 -1510
rect -686 -2040 -668 -1610
rect -510 -2040 -488 -1610
rect -686 -2160 -488 -2040
rect -686 -2600 -660 -2160
rect -530 -2600 -488 -2160
rect 4317 -1770 4515 -1544
rect 4317 -1844 4375 -1770
rect 4449 -1844 4515 -1770
rect 4317 -2244 4515 -1844
rect 4317 -2318 4375 -2244
rect 4449 -2318 4515 -2244
rect -686 -2688 -488 -2600
rect -686 -2730 -622 -2688
rect -548 -2730 -488 -2688
rect -686 -3140 -660 -2730
rect -500 -3140 -488 -2730
rect -686 -3180 -488 -3140
rect 4317 -2718 4515 -2318
rect 4317 -2792 4375 -2718
rect 4449 -2792 4515 -2718
rect 200 -3180 660 -3170
rect 2780 -3180 3240 -3170
rect 4317 -3180 4515 -2792
rect -686 -3248 4515 -3180
rect -686 -3322 -92 -3248
rect -18 -3322 456 -3248
rect 530 -3322 1004 -3248
rect 1078 -3322 1552 -3248
rect 1626 -3322 2100 -3248
rect 2174 -3322 2648 -3248
rect 2722 -3322 3198 -3248
rect 3272 -3322 4515 -3248
rect -686 -3378 4515 -3322
<< viali >>
rect -650 1946 -628 1970
rect -628 1946 -554 1970
rect -554 1946 -520 1970
rect -650 1570 -520 1946
rect -666 1072 -530 1430
rect -666 998 -628 1072
rect -628 998 -554 1072
rect -554 998 -530 1072
rect -666 990 -530 998
rect 4048 1156 4147 1260
rect -666 598 -510 870
rect -666 524 -628 598
rect -628 524 -554 598
rect -554 524 -510 598
rect -666 440 -510 524
rect 939 176 974 210
rect 1084 192 1118 226
rect 1168 192 1202 226
rect 1252 192 1286 226
rect 1336 192 1370 226
rect 1420 192 1454 226
rect 1504 192 1538 226
rect 1588 192 1622 226
rect 1672 192 1706 226
rect 1840 192 1874 226
rect 1924 192 1958 226
rect 2008 192 2042 226
rect 2080 192 2114 226
rect 2164 192 2198 226
rect 2248 192 2282 226
rect 2320 192 2354 226
rect 2404 192 2438 226
rect 2476 192 2510 226
rect 2632 192 2666 226
rect 2716 192 2750 226
rect 2788 192 2822 226
rect 2917 192 2951 226
rect 2989 192 3023 226
rect 3299 193 3333 227
rect 3371 193 3405 227
rect 3443 193 3477 227
rect 3515 193 3549 227
rect 3587 193 3621 227
rect 3659 193 3693 227
rect 3732 193 3766 227
rect 3804 193 3838 227
rect 3876 193 3910 227
rect 3948 193 3982 227
rect 4020 193 4054 227
rect 4092 193 4126 227
rect 939 93 974 127
rect 939 10 974 44
rect 939 -73 974 -39
rect -600 -164 -566 -130
rect -444 -164 -410 -130
rect -290 -164 -256 -130
rect -146 -164 -112 -130
rect -32 -164 2 -130
rect 82 -164 116 -130
rect 166 -164 200 -130
rect 250 -164 284 -130
rect 334 -164 368 -130
rect 418 -164 452 -130
rect 502 -164 536 -130
rect 586 -164 620 -130
rect 670 -164 704 -130
rect 754 -164 788 -130
rect 838 -164 872 -130
rect 922 -164 956 -130
rect 1102 -78 1136 -28
rect -38 -331 -4 -255
rect 54 -331 88 -255
rect 148 -331 182 -289
rect 240 -331 274 -255
rect 332 -331 366 -289
rect 424 -331 458 -255
rect 516 -331 550 -289
rect 608 -331 642 -255
rect 700 -331 734 -289
rect 794 -331 828 -255
rect 886 -331 920 -255
rect 1190 -78 1224 -28
rect 1278 -310 1312 -260
rect 1366 -78 1400 -28
rect 1454 3 1488 37
rect 1542 -78 1576 -28
rect 1630 -78 1664 -28
rect 2579 93 2613 127
rect 22 -430 69 -390
rect 807 -430 854 -390
rect 1190 -436 1226 -402
rect 1889 -78 1923 -28
rect 1977 -78 2011 -28
rect 2065 0 2099 34
rect 2153 -78 2187 -28
rect 2241 -310 2275 -260
rect 2329 -78 2363 -28
rect 2417 -78 2451 -28
rect 2579 10 2613 44
rect 2579 -73 2613 -39
rect 2579 -156 2613 -122
rect 1544 -447 1606 -413
rect 1949 -447 2011 -413
rect 2329 -436 2363 -402
rect 3463 -401 3497 -350
rect 3549 -401 3583 -350
rect 3633 -400 3667 -349
rect 3717 -401 3751 -350
rect 196 -526 244 -492
rect 638 -524 686 -490
rect 2721 -552 2755 -501
rect 2806 -551 2840 -500
rect 2890 -552 2924 -501
rect 2978 -551 3012 -500
rect 3061 -551 3095 -500
rect -16 -961 18 -900
rect 72 -961 106 -900
rect 160 -620 194 -585
rect 248 -961 282 -900
rect 342 -620 370 -585
rect 370 -620 376 -585
rect 506 -620 512 -585
rect 512 -620 540 -585
rect 424 -961 458 -900
rect 600 -961 634 -900
rect 688 -620 722 -585
rect 776 -961 810 -900
rect 864 -961 898 -900
rect 1670 -705 1718 -652
rect 1670 -707 1718 -705
rect 1836 -706 1884 -652
rect 1836 -707 1884 -706
rect -16 -1158 18 -1082
rect 72 -1158 106 -1082
rect 160 -1158 194 -1082
rect 68 -1238 110 -1237
rect 68 -1272 110 -1238
rect 248 -1158 282 -1082
rect 336 -1158 370 -1082
rect 244 -1238 286 -1237
rect 244 -1272 286 -1238
rect 424 -1158 458 -1082
rect 512 -1158 546 -1082
rect 420 -1238 462 -1237
rect 420 -1272 462 -1238
rect 600 -1158 634 -1082
rect 688 -1158 722 -1082
rect 596 -1238 638 -1237
rect 596 -1272 638 -1238
rect 776 -1158 810 -1082
rect 864 -1158 898 -1082
rect 772 -1238 814 -1237
rect 772 -1272 814 -1238
rect 1475 -1176 1509 -1132
rect 1567 -1176 1601 -1132
rect 1663 -1057 1697 -1012
rect 1759 -1176 1793 -1132
rect 1855 -972 1889 -927
rect 1951 -1176 1985 -1132
rect 2043 -1176 2077 -1132
rect 3447 -970 3481 -936
rect 3519 -970 3553 -936
rect 3591 -970 3625 -936
rect 3663 -970 3697 -936
rect 3735 -970 3769 -936
rect 1649 -1242 1683 -1232
rect 1649 -1276 1655 -1242
rect 1655 -1276 1683 -1242
rect 1649 -1278 1683 -1276
rect 1871 -1242 1905 -1232
rect 1871 -1276 1893 -1242
rect 1893 -1276 1905 -1242
rect 1871 -1278 1905 -1276
rect 2789 -1274 2823 -1240
rect 2865 -1274 2899 -1240
rect 2941 -1274 2975 -1240
rect 3017 -1274 3051 -1240
rect 3206 -1274 3240 -1240
rect 3282 -1274 3316 -1240
rect 3358 -1274 3392 -1240
rect 3434 -1274 3468 -1240
rect 3510 -1274 3544 -1240
rect 3586 -1274 3620 -1240
rect 3662 -1274 3696 -1240
rect 3738 -1274 3772 -1240
rect 4331 -1256 4365 -1222
rect 4403 -1256 4437 -1222
rect 4475 -1256 4509 -1222
rect -670 -1400 -636 -1366
rect -598 -1400 -564 -1366
rect -526 -1400 -492 -1366
rect 100 -1368 136 -1332
rect 218 -1368 254 -1332
rect 336 -1368 372 -1332
rect 454 -1368 490 -1332
rect 572 -1368 608 -1332
rect 690 -1368 726 -1332
rect 808 -1368 844 -1332
rect 1121 -1362 1157 -1340
rect 1121 -1376 1157 -1362
rect 1213 -1362 1249 -1340
rect 1213 -1376 1249 -1362
rect 1305 -1362 1341 -1340
rect 1305 -1376 1341 -1362
rect 1397 -1362 1433 -1340
rect 1397 -1376 1433 -1362
rect 1489 -1362 1525 -1340
rect 1489 -1376 1525 -1362
rect 1581 -1362 1617 -1340
rect 1581 -1376 1617 -1362
rect 1673 -1362 1709 -1340
rect 1673 -1376 1709 -1362
rect 1769 -1362 1805 -1340
rect 1769 -1376 1805 -1362
rect 1857 -1362 1893 -1340
rect 1857 -1376 1893 -1362
rect 1949 -1362 1985 -1340
rect 1949 -1376 1985 -1362
rect 2041 -1362 2077 -1340
rect 2041 -1376 2077 -1362
rect 2133 -1362 2169 -1340
rect 2133 -1376 2169 -1362
rect 2286 -1380 2322 -1344
rect 2360 -1380 2396 -1344
rect 2440 -1380 2476 -1344
rect 2520 -1380 2556 -1344
rect 2595 -1380 2631 -1344
rect 2669 -1380 2705 -1344
rect 2749 -1380 2785 -1344
rect 2829 -1380 2865 -1344
rect 2903 -1380 2939 -1344
rect 2983 -1380 3019 -1344
rect 3063 -1380 3099 -1344
rect 3143 -1380 3179 -1344
rect -670 -1472 -636 -1438
rect -598 -1472 -564 -1438
rect -526 -1472 -492 -1438
rect -672 -1544 -638 -1510
rect -600 -1544 -566 -1510
rect -528 -1544 -494 -1510
rect 4331 -1328 4365 -1294
rect 4403 -1328 4437 -1294
rect 4475 -1328 4509 -1294
rect 4331 -1400 4365 -1366
rect 4403 -1400 4437 -1366
rect 4475 -1400 4509 -1366
rect 4331 -1472 4365 -1438
rect 4403 -1472 4437 -1438
rect 4475 -1472 4509 -1438
rect 4331 -1544 4365 -1510
rect 4403 -1544 4437 -1510
rect 4475 -1544 4509 -1510
rect -668 -1740 -510 -1610
rect -668 -1814 -622 -1740
rect -622 -1814 -548 -1740
rect -548 -1814 -510 -1740
rect -668 -2040 -510 -1814
rect -660 -2214 -530 -2160
rect -660 -2288 -622 -2214
rect -622 -2288 -548 -2214
rect -548 -2288 -530 -2214
rect -660 -2600 -530 -2288
rect 4048 -2434 4147 -2330
rect -660 -2762 -622 -2730
rect -622 -2762 -548 -2730
rect -548 -2762 -500 -2730
rect -660 -3140 -500 -2762
<< metal1 >>
rect -686 1970 -450 2000
rect -686 1570 -650 1970
rect -520 1570 -450 1970
rect -686 1530 -450 1570
rect 3890 1520 4154 1651
rect -686 1430 -510 1450
rect -686 990 -666 1430
rect -530 990 -510 1430
rect -686 970 -510 990
rect 4042 1260 4154 1520
rect 4042 1156 4048 1260
rect 4147 1156 4154 1260
rect 4042 900 4154 1156
rect -686 870 -450 890
rect -686 440 -666 870
rect -510 440 -450 870
rect 3890 769 4154 900
rect -686 420 -450 440
rect 809 370 4978 392
rect 809 227 4678 370
rect 809 226 3299 227
rect 809 210 1084 226
rect 809 176 939 210
rect 974 192 1084 210
rect 1118 192 1168 226
rect 1202 192 1252 226
rect 1286 192 1336 226
rect 1370 192 1420 226
rect 1454 192 1504 226
rect 1538 192 1588 226
rect 1622 192 1672 226
rect 1706 192 1840 226
rect 1874 192 1924 226
rect 1958 192 2008 226
rect 2042 192 2080 226
rect 2114 192 2164 226
rect 2198 192 2248 226
rect 2282 192 2320 226
rect 2354 192 2404 226
rect 2438 192 2476 226
rect 2510 192 2632 226
rect 2666 192 2716 226
rect 2750 192 2788 226
rect 2822 192 2917 226
rect 2951 192 2989 226
rect 3023 193 3299 226
rect 3333 193 3371 227
rect 3405 193 3443 227
rect 3477 193 3515 227
rect 3549 193 3587 227
rect 3621 193 3659 227
rect 3693 193 3732 227
rect 3766 193 3804 227
rect 3838 193 3876 227
rect 3910 193 3948 227
rect 3982 193 4020 227
rect 4054 193 4092 227
rect 4126 193 4678 227
rect 3023 192 4678 193
rect 974 186 4678 192
rect 4958 186 4978 370
rect 974 176 980 186
rect 809 127 980 176
rect 809 93 939 127
rect 974 93 980 127
rect 809 44 980 93
rect 809 10 939 44
rect 974 10 980 44
rect 809 -39 980 10
rect 1448 37 1494 186
rect 1448 3 1454 37
rect 1488 3 1494 37
rect 1448 -9 1494 3
rect 2059 34 2105 186
rect 2059 0 2065 34
rect 2099 0 2105 34
rect 2059 -12 2105 0
rect 2573 127 2619 186
rect 2573 93 2579 127
rect 2613 93 2619 127
rect 2573 44 2619 93
rect 2573 10 2579 44
rect 2613 10 2619 44
rect 809 -73 939 -39
rect 974 -73 980 -39
rect -641 -122 80 -101
rect 809 -122 980 -73
rect 1096 -28 1142 -16
rect 1096 -78 1102 -28
rect 1136 -41 1142 -28
rect 1184 -28 1230 -16
rect 1184 -41 1190 -28
rect 1136 -69 1190 -41
rect 1136 -78 1142 -69
rect 1096 -90 1142 -78
rect 1184 -78 1190 -69
rect 1224 -41 1230 -28
rect 1360 -28 1406 -16
rect 1360 -41 1366 -28
rect 1224 -69 1366 -41
rect 1224 -78 1230 -69
rect 1184 -90 1230 -78
rect 1360 -78 1366 -69
rect 1400 -41 1406 -28
rect 1536 -28 1582 -16
rect 1536 -41 1542 -28
rect 1400 -69 1542 -41
rect 1400 -78 1406 -69
rect 1360 -90 1406 -78
rect 1536 -78 1542 -69
rect 1576 -41 1582 -28
rect 1624 -28 1670 -16
rect 1624 -41 1630 -28
rect 1576 -69 1630 -41
rect 1576 -78 1582 -69
rect 1536 -90 1582 -78
rect 1624 -78 1630 -69
rect 1664 -78 1670 -28
rect 1624 -90 1670 -78
rect 1883 -28 1929 -16
rect 1883 -78 1889 -28
rect 1923 -41 1929 -28
rect 1971 -28 2017 -16
rect 1971 -41 1977 -28
rect 1923 -69 1977 -41
rect 1923 -78 1929 -69
rect 1883 -90 1929 -78
rect 1971 -78 1977 -69
rect 2011 -41 2017 -28
rect 2147 -28 2193 -16
rect 2147 -41 2153 -28
rect 2011 -69 2153 -41
rect 2011 -78 2017 -69
rect 1971 -90 2017 -78
rect 2147 -78 2153 -69
rect 2187 -41 2193 -28
rect 2323 -28 2369 -16
rect 2323 -41 2329 -28
rect 2187 -69 2329 -41
rect 2187 -78 2193 -69
rect 2147 -90 2193 -78
rect 2323 -78 2329 -69
rect 2363 -41 2369 -28
rect 2411 -28 2457 -16
rect 2411 -41 2417 -28
rect 2363 -69 2417 -41
rect 2363 -78 2369 -69
rect 2323 -90 2369 -78
rect 2411 -78 2417 -69
rect 2451 -78 2457 -28
rect 2411 -90 2457 -78
rect 2573 -39 2619 10
rect 2573 -73 2579 -39
rect 2613 -73 2619 -39
rect -641 -130 980 -122
rect -641 -164 -600 -130
rect -566 -164 -444 -130
rect -410 -164 -290 -130
rect -256 -164 -146 -130
rect -112 -164 -32 -130
rect 2 -164 82 -130
rect 116 -164 166 -130
rect 200 -164 250 -130
rect 284 -164 334 -130
rect 368 -164 418 -130
rect 452 -164 502 -130
rect 536 -164 586 -130
rect 620 -164 670 -130
rect 704 -164 754 -130
rect 788 -164 838 -130
rect 872 -164 922 -130
rect 956 -164 980 -130
rect -641 -177 980 -164
rect 2573 -122 2619 -73
rect 2573 -156 2579 -122
rect 2613 -156 2619 -122
rect 48 -239 94 -177
rect -44 -255 94 -239
rect 233 -253 280 -177
rect -44 -331 -38 -255
rect -4 -331 54 -255
rect 88 -331 94 -255
rect 234 -255 280 -253
rect -44 -347 94 -331
rect 142 -289 188 -277
rect 142 -331 148 -289
rect 182 -331 188 -289
rect 142 -375 188 -331
rect 234 -331 240 -255
rect 274 -331 280 -255
rect 418 -255 464 -177
rect 234 -347 280 -331
rect 326 -289 372 -277
rect 326 -331 332 -289
rect 366 -331 372 -289
rect 326 -375 372 -331
rect 418 -331 424 -255
rect 458 -331 464 -255
rect 602 -255 648 -177
rect 418 -347 464 -331
rect 510 -289 556 -277
rect 510 -331 516 -289
rect 550 -331 556 -289
rect -99 -437 -93 -383
rect -23 -390 81 -383
rect -23 -430 22 -390
rect 69 -430 81 -390
rect 142 -407 372 -375
rect -23 -437 81 -430
rect 327 -450 372 -407
rect 510 -379 556 -331
rect 602 -331 608 -255
rect 642 -331 648 -255
rect 788 -239 834 -177
rect 2573 -191 2619 -156
rect 2651 -212 2721 -184
rect 788 -255 926 -239
rect 602 -347 648 -331
rect 694 -289 740 -277
rect 694 -331 700 -289
rect 734 -331 740 -289
rect 694 -379 740 -331
rect 788 -331 794 -255
rect 828 -331 886 -255
rect 920 -331 926 -255
rect 1269 -260 1321 -240
rect 1269 -310 1278 -260
rect 1312 -310 1321 -260
rect 1269 -316 1321 -310
rect 2232 -260 2284 -241
rect 2232 -310 2241 -260
rect 2275 -310 2284 -260
rect 2232 -316 2284 -310
rect 788 -347 926 -331
rect 510 -407 740 -379
rect 795 -390 908 -383
rect 510 -450 555 -407
rect 795 -430 807 -390
rect 854 -430 908 -390
rect 795 -437 908 -430
rect 978 -437 984 -383
rect 1174 -396 1244 -386
rect 327 -456 383 -450
rect 180 -526 192 -474
rect 246 -526 260 -474
rect 180 -533 260 -526
rect 379 -508 383 -456
rect 154 -585 206 -568
rect 154 -620 160 -585
rect 194 -604 206 -585
rect 327 -585 383 -508
rect 327 -604 342 -585
rect 194 -620 342 -604
rect 376 -620 383 -585
rect 154 -632 383 -620
rect 499 -456 555 -450
rect 1174 -448 1180 -396
rect 1234 -448 1244 -396
rect 1174 -453 1244 -448
rect 499 -508 503 -456
rect 499 -585 555 -508
rect 622 -524 635 -472
rect 689 -524 702 -472
rect 622 -531 702 -524
rect 1272 -548 1318 -316
rect 1530 -413 1618 -397
rect 1530 -447 1544 -413
rect 1606 -430 1618 -413
rect 1935 -413 2023 -397
rect 1935 -430 1949 -413
rect 1606 -447 1684 -430
rect 1530 -463 1684 -447
rect 1678 -482 1684 -463
rect 1736 -482 1742 -430
rect 1811 -482 1817 -430
rect 1869 -447 1949 -430
rect 2011 -447 2023 -413
rect 1869 -463 2023 -447
rect 1869 -482 1875 -463
rect 1811 -548 1839 -482
rect 2235 -548 2281 -316
rect 2313 -396 2379 -386
rect 2651 -396 2679 -212
rect 2313 -448 2321 -396
rect 2373 -448 2379 -396
rect 2313 -454 2379 -448
rect 2637 -428 2679 -396
rect 3307 -349 4157 -314
rect 3307 -350 3633 -349
rect 3307 -401 3463 -350
rect 3497 -401 3549 -350
rect 3583 -400 3633 -350
rect 3667 -350 4157 -349
rect 3667 -400 3717 -350
rect 3583 -401 3717 -400
rect 3751 -361 4157 -350
rect 3751 -401 3981 -361
rect 3307 -413 3981 -401
rect 4033 -413 4060 -361
rect 4112 -413 4157 -361
rect 499 -620 506 -585
rect 540 -603 555 -585
rect 676 -585 728 -567
rect 1272 -576 1624 -548
rect 676 -603 688 -585
rect 540 -620 688 -603
rect 722 -620 728 -585
rect 1618 -600 1624 -576
rect 1676 -576 1839 -548
rect 1676 -600 1682 -576
rect 1867 -600 1873 -548
rect 1925 -576 2281 -548
rect 1925 -600 1931 -576
rect 499 -632 728 -620
rect 1654 -652 1734 -646
rect 1654 -707 1670 -652
rect 1718 -707 1734 -652
rect 1654 -708 1734 -707
rect 1654 -760 1670 -708
rect 1722 -760 1734 -708
rect 1654 -766 1734 -760
rect 1820 -652 1900 -646
rect 1820 -707 1836 -652
rect 1884 -707 1900 -652
rect 1820 -708 1900 -707
rect 1820 -760 1833 -708
rect 1885 -760 1900 -708
rect 1820 -766 1900 -760
rect -22 -900 24 -867
rect -486 -962 -398 -953
rect -486 -1018 -480 -962
rect -404 -1018 -398 -962
rect -486 -1027 -398 -1018
rect -22 -961 -16 -900
rect 18 -961 24 -900
rect -22 -1004 24 -961
rect 66 -900 112 -867
rect 66 -961 72 -900
rect 106 -961 112 -900
rect 66 -1004 112 -961
rect 242 -900 288 -867
rect 242 -961 248 -900
rect 282 -961 288 -900
rect 242 -1004 288 -961
rect 418 -900 464 -867
rect 418 -961 424 -900
rect 458 -961 464 -900
rect 418 -1004 464 -961
rect 594 -900 640 -867
rect 594 -961 600 -900
rect 634 -961 640 -900
rect 594 -1004 640 -961
rect 770 -900 816 -867
rect 770 -961 776 -900
rect 810 -961 816 -900
rect 770 -1004 816 -961
rect 858 -900 904 -867
rect 858 -961 864 -900
rect 898 -961 904 -900
rect 1648 -923 1712 -921
rect 1648 -950 1654 -923
rect 858 -1004 904 -961
rect 1353 -975 1654 -950
rect 1706 -950 1712 -923
rect 1839 -927 1903 -921
rect 1839 -950 1855 -927
rect 1706 -972 1855 -950
rect 1889 -950 1903 -927
rect 2637 -950 2665 -428
rect 3307 -436 4157 -413
rect 3307 -462 3367 -436
rect 2695 -500 3367 -462
rect 2695 -501 2806 -500
rect 2695 -552 2721 -501
rect 2755 -551 2806 -501
rect 2840 -501 2978 -500
rect 2840 -551 2890 -501
rect 2755 -552 2890 -551
rect 2924 -551 2978 -501
rect 3012 -551 3061 -500
rect 3095 -525 3367 -500
rect 3095 -551 3119 -525
rect 2924 -552 3119 -551
rect 2695 -590 3119 -552
rect 1889 -972 2665 -950
rect 1706 -975 2665 -972
rect 1353 -978 2665 -975
rect -22 -1036 904 -1004
rect 2693 -1006 2721 -840
rect 3407 -936 3825 -928
rect 3407 -970 3447 -936
rect 3481 -970 3519 -936
rect 3553 -970 3591 -936
rect 3625 -970 3663 -936
rect 3697 -970 3735 -936
rect 3769 -970 3825 -936
rect 3407 -978 3825 -970
rect 1353 -1008 2721 -1006
rect 1353 -1012 1845 -1008
rect 1353 -1034 1663 -1012
rect -22 -1082 24 -1036
rect -22 -1158 -16 -1082
rect 18 -1158 24 -1082
rect -22 -1174 24 -1158
rect 66 -1082 112 -1036
rect 66 -1158 72 -1082
rect 106 -1158 112 -1082
rect 66 -1174 112 -1158
rect 154 -1082 200 -1064
rect 154 -1158 160 -1082
rect 194 -1158 200 -1082
rect 154 -1174 200 -1158
rect 242 -1082 288 -1036
rect 242 -1158 248 -1082
rect 282 -1158 288 -1082
rect 242 -1174 288 -1158
rect 330 -1082 376 -1064
rect 330 -1158 336 -1082
rect 370 -1158 376 -1082
rect 330 -1174 376 -1158
rect 418 -1082 464 -1036
rect 418 -1158 424 -1082
rect 458 -1158 464 -1082
rect 418 -1174 464 -1158
rect 506 -1082 552 -1064
rect 506 -1158 512 -1082
rect 546 -1158 552 -1082
rect 506 -1174 552 -1158
rect 594 -1082 640 -1036
rect 594 -1158 600 -1082
rect 634 -1158 640 -1082
rect 594 -1174 640 -1158
rect 682 -1082 728 -1064
rect 682 -1158 688 -1082
rect 722 -1158 728 -1082
rect 682 -1174 728 -1158
rect 770 -1082 816 -1036
rect 770 -1158 776 -1082
rect 810 -1158 816 -1082
rect 770 -1174 816 -1158
rect 858 -1082 904 -1036
rect 1648 -1057 1663 -1034
rect 1697 -1034 1845 -1012
rect 1697 -1057 1712 -1034
rect 1648 -1063 1712 -1057
rect 1839 -1060 1845 -1034
rect 1897 -1034 2721 -1008
rect 3697 -979 3825 -978
rect 3697 -1032 3703 -979
rect 3755 -1032 3767 -979
rect 3819 -1032 3825 -979
rect 1897 -1060 1903 -1034
rect 1839 -1063 1903 -1060
rect 858 -1158 864 -1082
rect 898 -1158 904 -1082
rect 858 -1174 904 -1158
rect 1463 -1132 1607 -1118
rect 1463 -1176 1475 -1132
rect 1509 -1176 1567 -1132
rect 1601 -1176 1607 -1132
rect 1463 -1182 1607 -1176
rect 30 -1237 852 -1226
rect 30 -1244 68 -1237
rect -99 -1296 -92 -1244
rect -38 -1272 68 -1244
rect 110 -1272 244 -1237
rect 286 -1272 420 -1237
rect 462 -1272 596 -1237
rect 638 -1272 772 -1237
rect 814 -1244 852 -1237
rect 814 -1272 924 -1244
rect -38 -1296 924 -1272
rect 978 -1296 984 -1244
rect -99 -1298 984 -1296
rect 1561 -1326 1607 -1182
rect 1753 -1132 1799 -1118
rect 1753 -1176 1759 -1132
rect 1793 -1176 1799 -1132
rect 1635 -1226 1705 -1218
rect 1635 -1278 1643 -1226
rect 1697 -1278 1705 -1226
rect 1635 -1284 1705 -1278
rect 1753 -1326 1799 -1176
rect 1945 -1132 2089 -1118
rect 1945 -1176 1951 -1132
rect 1985 -1176 2043 -1132
rect 2077 -1176 2089 -1132
rect 1945 -1182 2089 -1176
rect 3681 -1168 3830 -1156
rect 1847 -1226 1917 -1218
rect 1847 -1278 1854 -1226
rect 1908 -1278 1917 -1226
rect 1847 -1284 1917 -1278
rect 1945 -1326 1991 -1182
rect 3681 -1234 3699 -1168
rect 2762 -1240 3699 -1234
rect 2762 -1274 2789 -1240
rect 2823 -1274 2865 -1240
rect 2899 -1274 2941 -1240
rect 2975 -1274 3017 -1240
rect 3051 -1274 3206 -1240
rect 3240 -1274 3282 -1240
rect 3316 -1274 3358 -1240
rect 3392 -1274 3434 -1240
rect 3468 -1274 3510 -1240
rect 3544 -1274 3586 -1240
rect 3620 -1274 3662 -1240
rect 3696 -1268 3699 -1240
rect 3814 -1268 3830 -1168
rect 3696 -1274 3738 -1268
rect 3772 -1274 3830 -1268
rect 2762 -1280 3830 -1274
rect 4317 -1222 4515 -1202
rect 4317 -1256 4331 -1222
rect 4365 -1256 4403 -1222
rect 4437 -1256 4475 -1222
rect 4509 -1256 4515 -1222
rect 4317 -1294 4515 -1256
rect 4317 -1326 4331 -1294
rect -686 -1328 4331 -1326
rect 4365 -1328 4403 -1294
rect 4437 -1328 4475 -1294
rect 4509 -1326 4515 -1294
rect 4509 -1328 4588 -1326
rect -686 -1332 4588 -1328
rect -686 -1354 100 -1332
rect -686 -1366 -422 -1354
rect -686 -1400 -670 -1366
rect -636 -1400 -598 -1366
rect -564 -1400 -526 -1366
rect -492 -1400 -422 -1366
rect 136 -1368 218 -1332
rect 254 -1368 336 -1332
rect 372 -1368 454 -1332
rect 490 -1368 572 -1332
rect 608 -1368 690 -1332
rect 726 -1368 808 -1332
rect 844 -1340 4588 -1332
rect 844 -1368 1121 -1340
rect -686 -1438 -422 -1400
rect -686 -1472 -670 -1438
rect -636 -1472 -598 -1438
rect -564 -1472 -526 -1438
rect -492 -1472 -422 -1438
rect -686 -1510 -422 -1472
rect -686 -1544 -672 -1510
rect -638 -1544 -600 -1510
rect -566 -1544 -528 -1510
rect -494 -1520 -422 -1510
rect 126 -1376 1121 -1368
rect 1157 -1376 1213 -1340
rect 1249 -1376 1305 -1340
rect 1341 -1376 1397 -1340
rect 1433 -1376 1489 -1340
rect 1525 -1376 1581 -1340
rect 1617 -1376 1673 -1340
rect 1709 -1376 1750 -1340
rect 1805 -1376 1857 -1340
rect 1893 -1376 1949 -1340
rect 1985 -1376 2041 -1340
rect 2077 -1376 2133 -1340
rect 2169 -1344 4588 -1340
rect 2169 -1376 2286 -1344
rect 126 -1392 1750 -1376
rect 1802 -1380 2286 -1376
rect 2322 -1380 2360 -1344
rect 2396 -1380 2440 -1344
rect 2476 -1380 2520 -1344
rect 2556 -1380 2595 -1344
rect 2631 -1380 2669 -1344
rect 2705 -1380 2749 -1344
rect 2785 -1380 2829 -1344
rect 2865 -1380 2903 -1344
rect 2939 -1380 2983 -1344
rect 3019 -1380 3063 -1344
rect 3099 -1380 3143 -1344
rect 3179 -1350 4588 -1344
rect 3179 -1366 4526 -1350
rect 3179 -1380 4331 -1366
rect 1802 -1392 4331 -1380
rect 126 -1400 4331 -1392
rect 4365 -1400 4403 -1366
rect 4437 -1400 4475 -1366
rect 4509 -1400 4526 -1366
rect 126 -1438 4526 -1400
rect 126 -1472 4331 -1438
rect 4365 -1472 4403 -1438
rect 4437 -1472 4475 -1438
rect 4509 -1472 4526 -1438
rect 126 -1510 4526 -1472
rect 126 -1520 4331 -1510
rect -494 -1544 4331 -1520
rect 4365 -1544 4403 -1510
rect 4437 -1544 4475 -1510
rect 4509 -1540 4526 -1510
rect 4578 -1540 4588 -1350
rect 4509 -1544 4588 -1540
rect -686 -1558 4588 -1544
rect -686 -1610 -450 -1590
rect -686 -2040 -668 -1610
rect -510 -2040 -450 -1610
rect -686 -2060 -450 -2040
rect 3890 -2070 4154 -1939
rect -686 -2160 -510 -2140
rect -686 -2600 -660 -2160
rect -530 -2600 -510 -2160
rect -686 -2620 -510 -2600
rect 4042 -2330 4154 -2070
rect 4042 -2434 4048 -2330
rect 4147 -2434 4154 -2330
rect 4042 -2690 4154 -2434
rect -686 -2730 -450 -2700
rect -686 -3140 -660 -2730
rect -500 -3140 -450 -2730
rect 3890 -2821 4154 -2690
rect -686 -3170 -450 -3140
<< via1 >>
rect -650 1570 -520 1970
rect -666 990 -530 1430
rect 4048 1156 4147 1260
rect 4678 186 4958 370
rect -93 -437 -23 -383
rect 908 -437 978 -383
rect 192 -492 246 -474
rect 192 -526 196 -492
rect 196 -526 244 -492
rect 244 -526 246 -492
rect 327 -508 379 -456
rect 1180 -402 1234 -396
rect 1180 -436 1190 -402
rect 1190 -436 1226 -402
rect 1226 -436 1234 -402
rect 1180 -448 1234 -436
rect 503 -508 555 -456
rect 635 -490 689 -472
rect 635 -524 638 -490
rect 638 -524 686 -490
rect 686 -524 689 -490
rect 1684 -482 1736 -430
rect 1817 -482 1869 -430
rect 2321 -402 2373 -396
rect 2321 -436 2329 -402
rect 2329 -436 2363 -402
rect 2363 -436 2373 -402
rect 2321 -448 2373 -436
rect 3981 -413 4033 -361
rect 4060 -413 4112 -361
rect 1624 -600 1676 -548
rect 1873 -600 1925 -548
rect 1670 -760 1722 -708
rect 1833 -760 1885 -708
rect -480 -1018 -404 -962
rect 1654 -975 1706 -923
rect 1845 -1060 1897 -1008
rect 3703 -1032 3755 -979
rect 3767 -1032 3819 -979
rect -92 -1296 -38 -1244
rect 924 -1296 978 -1244
rect 1643 -1232 1697 -1226
rect 1643 -1278 1649 -1232
rect 1649 -1278 1683 -1232
rect 1683 -1278 1697 -1232
rect 1854 -1232 1908 -1226
rect 1854 -1278 1871 -1232
rect 1871 -1278 1905 -1232
rect 1905 -1278 1908 -1232
rect 3699 -1240 3814 -1168
rect 3699 -1268 3738 -1240
rect 3738 -1268 3772 -1240
rect 3772 -1268 3814 -1240
rect -422 -1368 100 -1354
rect 100 -1368 126 -1354
rect -422 -1520 126 -1368
rect 1750 -1376 1769 -1340
rect 1769 -1376 1802 -1340
rect 1750 -1392 1802 -1376
rect 4526 -1540 4578 -1350
rect -660 -2600 -530 -2160
rect 4048 -2434 4147 -2330
rect -660 -3140 -528 -2730
<< metal2 >>
rect -686 1970 -450 2000
rect -686 1570 -650 1970
rect -520 1570 -450 1970
rect -686 1530 -450 1570
rect -686 1430 -510 1450
rect -686 990 -666 1430
rect -530 990 -510 1430
rect 4042 1260 4154 1265
rect 4042 1156 4048 1260
rect 4147 1156 4154 1260
rect 4042 1149 4154 1156
rect -686 970 -510 990
rect 1744 339 1808 420
rect 1744 266 1808 275
rect 4658 370 4978 392
rect 4658 180 4678 370
rect 4958 180 4978 370
rect 4658 162 4978 180
rect -99 -437 -93 -383
rect -23 -437 -17 -383
rect 902 -437 908 -383
rect 978 -437 984 -383
rect -486 -962 -398 -953
rect -486 -1018 -480 -962
rect -404 -1018 -398 -962
rect -486 -1027 -398 -1018
rect -99 -1244 -71 -437
rect 327 -456 383 -450
rect 179 -470 261 -460
rect 179 -526 190 -470
rect 246 -526 261 -470
rect 179 -533 261 -526
rect 379 -477 383 -456
rect 327 -542 383 -533
rect 499 -456 555 -450
rect 499 -477 503 -456
rect 620 -468 702 -458
rect 620 -524 634 -468
rect 690 -524 702 -468
rect 620 -531 702 -524
rect 499 -542 555 -533
rect 956 -1244 984 -437
rect 1174 -396 1244 -386
rect 1174 -448 1180 -396
rect 1234 -413 1244 -396
rect 2313 -396 2379 -386
rect 2313 -413 2321 -396
rect 1234 -422 1354 -413
rect 1234 -448 1298 -422
rect 1174 -453 1298 -448
rect 2198 -422 2321 -413
rect 1678 -454 1684 -430
rect 1298 -487 1354 -478
rect 1561 -482 1684 -454
rect 1736 -482 1742 -430
rect 1561 -708 1589 -482
rect 1710 -548 1742 -482
rect 1811 -482 1817 -430
rect 1869 -454 1875 -430
rect 1869 -482 1988 -454
rect 1811 -519 1839 -482
rect 1618 -600 1624 -548
rect 1676 -600 1682 -548
rect 1710 -576 1873 -548
rect 1867 -600 1873 -576
rect 1925 -600 1931 -548
rect 1960 -708 1988 -482
rect 2254 -448 2321 -422
rect 2373 -448 2379 -396
rect 3967 -419 3976 -361
rect 4033 -419 4060 -361
rect 4117 -419 4126 -361
rect 2254 -454 2379 -448
rect 2198 -487 2254 -478
rect 1561 -736 1670 -708
rect 1664 -760 1670 -736
rect 1722 -760 1728 -708
rect 1827 -760 1833 -708
rect 1885 -736 1988 -708
rect 1885 -760 1891 -736
rect 1678 -897 1706 -760
rect 1654 -923 1706 -897
rect 1654 -1066 1706 -975
rect 1845 -897 1873 -760
rect 1845 -1008 1897 -897
rect 1845 -1066 1897 -1060
rect 3681 -979 3830 -978
rect 3681 -1032 3703 -979
rect 3755 -1032 3767 -979
rect 3819 -1032 3830 -979
rect 1746 -1079 1806 -1070
rect 1746 -1135 1748 -1079
rect 1804 -1135 1806 -1079
rect -99 -1296 -92 -1244
rect -38 -1296 -31 -1244
rect -99 -1298 -31 -1296
rect 916 -1296 924 -1244
rect 978 -1296 984 -1244
rect 1633 -1222 1707 -1218
rect 1633 -1278 1642 -1222
rect 1698 -1278 1707 -1222
rect 1633 -1284 1707 -1278
rect 916 -1298 984 -1296
rect -450 -1354 190 -1326
rect -450 -1520 -422 -1354
rect 126 -1520 190 -1354
rect 1746 -1340 1806 -1135
rect 3681 -1105 3830 -1032
rect 3681 -1165 3698 -1105
rect 3813 -1165 3830 -1105
rect 3681 -1168 3830 -1165
rect 1844 -1222 1918 -1215
rect 1844 -1278 1853 -1222
rect 1909 -1278 1918 -1222
rect 1844 -1287 1918 -1278
rect 3681 -1268 3699 -1168
rect 3814 -1268 3830 -1168
rect 3681 -1280 3830 -1268
rect 1746 -1392 1750 -1340
rect 1802 -1392 1806 -1340
rect 1746 -1400 1806 -1392
rect 4268 -1350 4588 -1326
rect -450 -1590 190 -1520
rect 1744 -1443 1808 -1434
rect 1744 -1590 1808 -1507
rect 4268 -1540 4288 -1350
rect 4578 -1540 4588 -1350
rect 4268 -1558 4588 -1540
rect -686 -2160 -510 -2140
rect -686 -2600 -660 -2160
rect -530 -2600 -510 -2160
rect 4042 -2330 4154 -2325
rect 4042 -2434 4048 -2330
rect 4147 -2434 4154 -2330
rect 4042 -2441 4154 -2434
rect -686 -2620 -510 -2600
rect -686 -2730 -450 -2700
rect -686 -3140 -660 -2730
rect -528 -3140 -450 -2730
rect -686 -3170 -450 -3140
<< via2 >>
rect -650 1570 -520 1970
rect -666 990 -530 1430
rect 1744 275 1808 339
rect 4678 186 4958 370
rect 4678 180 4958 186
rect -480 -1018 -404 -962
rect 190 -474 246 -470
rect 190 -526 192 -474
rect 192 -526 246 -474
rect 327 -508 379 -477
rect 379 -508 383 -477
rect 327 -533 383 -508
rect 499 -508 503 -477
rect 503 -508 555 -477
rect 499 -533 555 -508
rect 634 -472 690 -468
rect 634 -524 635 -472
rect 635 -524 689 -472
rect 689 -524 690 -472
rect 1298 -478 1354 -422
rect 2198 -478 2254 -422
rect 3976 -413 3981 -361
rect 3981 -413 4033 -361
rect 3976 -419 4033 -413
rect 4060 -413 4112 -361
rect 4112 -413 4117 -361
rect 4060 -419 4117 -413
rect 1748 -1135 1804 -1079
rect 1642 -1226 1698 -1222
rect 1642 -1278 1643 -1226
rect 1643 -1278 1697 -1226
rect 1697 -1278 1698 -1226
rect -422 -1520 126 -1354
rect 3698 -1165 3813 -1105
rect 1853 -1226 1909 -1222
rect 1853 -1278 1854 -1226
rect 1854 -1278 1908 -1226
rect 1908 -1278 1909 -1226
rect 3699 -1268 3814 -1208
rect 1744 -1507 1808 -1443
rect 4288 -1540 4526 -1350
rect 4526 -1540 4578 -1350
rect -660 -2600 -530 -2160
rect -660 -3140 -528 -2730
<< metal3 >>
rect -686 1970 -512 2000
rect -686 1570 -650 1970
rect -520 1570 -512 1970
rect -686 1530 -512 1570
rect -686 1430 -510 1450
rect -686 990 -666 1430
rect -530 990 -510 1430
rect 3890 1258 4588 1265
rect 3890 1159 4291 1258
rect 4576 1159 4588 1258
rect 3890 1149 4588 1159
rect -686 970 -510 990
rect 4658 370 4978 392
rect 1724 339 1824 357
rect 1724 275 1744 339
rect 1808 275 1824 339
rect 1724 261 1824 275
rect 1291 -422 1361 -415
rect 185 -470 261 -461
rect 185 -526 190 -470
rect 246 -526 261 -470
rect 185 -533 261 -526
rect 322 -477 390 -459
rect 322 -533 327 -477
rect 383 -533 390 -477
rect 322 -560 390 -533
rect 320 -855 390 -560
rect 384 -919 390 -855
rect 320 -925 390 -919
rect 492 -477 560 -459
rect 492 -533 499 -477
rect 555 -533 560 -477
rect 620 -468 695 -459
rect 620 -524 634 -468
rect 690 -524 695 -468
rect 620 -531 695 -524
rect 1043 -483 1107 -470
rect 492 -560 560 -533
rect 492 -729 562 -560
rect 492 -793 498 -729
rect 492 -925 562 -793
rect 1043 -729 1107 -547
rect 1043 -925 1107 -793
rect 1167 -609 1231 -473
rect 1167 -855 1231 -673
rect 1291 -478 1298 -422
rect 1354 -478 1361 -422
rect 1746 -423 1806 201
rect 4658 180 4678 370
rect 4958 180 4978 370
rect 4658 162 4978 180
rect 3963 -358 4130 -356
rect 2191 -422 2261 -415
rect 1291 -483 1361 -478
rect 1291 -547 1294 -483
rect 1358 -547 1361 -483
rect 1291 -679 1361 -547
rect 1556 -733 1996 -423
rect 2191 -478 2198 -422
rect 2254 -478 2261 -422
rect 3963 -422 3969 -358
rect 4033 -422 4060 -358
rect 4124 -422 4130 -358
rect 3963 -424 4130 -422
rect 2191 -609 2261 -478
rect 2191 -673 2194 -609
rect 2258 -673 2261 -609
rect 2191 -679 2261 -673
rect 2322 -483 2386 -470
rect 2322 -729 2386 -547
rect 1167 -925 1231 -919
rect -486 -960 -398 -953
rect -486 -962 -165 -960
rect -486 -1018 -480 -962
rect -404 -1018 -165 -962
rect -486 -1020 -165 -1018
rect -486 -1027 -398 -1020
rect -230 -1204 -165 -1020
rect 1743 -1079 1809 -733
rect 2322 -925 2386 -793
rect 2448 -609 2512 -473
rect 2448 -855 2512 -673
rect 2448 -925 2512 -919
rect 1743 -1135 1748 -1079
rect 1804 -1135 1809 -1079
rect 4658 -1032 4978 -1022
rect 4658 -1087 4675 -1032
rect 1743 -1144 1809 -1135
rect 3681 -1105 4675 -1087
rect 3681 -1165 3698 -1105
rect 3813 -1145 4675 -1105
rect 4967 -1145 4978 -1032
rect 3813 -1156 4978 -1145
rect 3813 -1165 3830 -1156
rect -230 -1222 1918 -1204
rect -230 -1264 1642 -1222
rect 1630 -1278 1642 -1264
rect 1698 -1278 1853 -1222
rect 1909 -1278 1918 -1222
rect 1630 -1288 1918 -1278
rect 3681 -1208 3830 -1165
rect 3681 -1268 3699 -1208
rect 3814 -1268 3830 -1208
rect 3681 -1280 3830 -1268
rect -450 -1354 180 -1326
rect -450 -1520 -422 -1354
rect 126 -1520 180 -1354
rect 4268 -1350 4588 -1326
rect -450 -1526 180 -1520
rect 1724 -1443 1825 -1432
rect 1724 -1507 1744 -1443
rect 1808 -1507 1825 -1443
rect 1724 -1528 1825 -1507
rect 4268 -1540 4288 -1350
rect 4578 -1540 4588 -1350
rect 4268 -1558 4588 -1540
rect -686 -2160 -510 -2140
rect -686 -2600 -660 -2160
rect -530 -2600 -510 -2160
rect 3889 -2335 4588 -2325
rect 3889 -2434 4299 -2335
rect 4567 -2434 4588 -2335
rect 3889 -2442 4588 -2434
rect -686 -2620 -510 -2600
rect -686 -2730 -514 -2700
rect -686 -3140 -660 -2730
rect -528 -3140 -514 -2730
rect -686 -3170 -514 -3140
<< via3 >>
rect -650 1570 -520 1970
rect -666 990 -530 1430
rect 4291 1159 4576 1258
rect 1744 275 1808 339
rect 320 -919 384 -855
rect 1043 -547 1107 -483
rect 498 -793 562 -729
rect 1043 -793 1107 -729
rect 1167 -673 1231 -609
rect 4678 180 4958 370
rect 1294 -547 1358 -483
rect 3969 -361 4033 -358
rect 3969 -419 3976 -361
rect 3976 -419 4033 -361
rect 3969 -422 4033 -419
rect 4060 -361 4124 -358
rect 4060 -419 4117 -361
rect 4117 -419 4124 -361
rect 4060 -422 4124 -419
rect 2194 -673 2258 -609
rect 2322 -547 2386 -483
rect 1167 -919 1231 -855
rect 2322 -793 2386 -729
rect 2448 -673 2512 -609
rect 2448 -919 2512 -855
rect 4675 -1145 4967 -1032
rect 1744 -1507 1808 -1443
rect 4288 -1540 4578 -1350
rect -660 -2600 -530 -2160
rect 4299 -2434 4567 -2335
rect -660 -3140 -528 -2730
<< metal4 >>
rect -686 1970 -450 2000
rect -686 1570 -650 1970
rect -520 1570 -450 1970
rect 4268 1651 4588 2218
rect -686 1530 -450 1570
rect 3890 1530 4588 1651
rect -686 1430 -450 1450
rect -686 990 -666 1430
rect -530 990 -450 1430
rect -686 970 -450 990
rect 4268 1258 4588 1530
rect 4268 1159 4291 1258
rect 4576 1159 4588 1258
rect 4268 890 4588 1159
rect 3890 769 4588 890
rect 1743 339 1809 340
rect 1743 275 1744 339
rect 1808 275 1809 339
rect 1743 274 1809 275
rect 1042 -483 1108 -482
rect 1042 -547 1043 -483
rect 1107 -488 1108 -483
rect 1293 -483 1359 -482
rect 1293 -488 1294 -483
rect 1107 -547 1294 -488
rect 1358 -488 1359 -483
rect 1746 -488 1806 274
rect 4268 -356 4588 769
rect 3963 -358 4588 -356
rect 3963 -422 3969 -358
rect 4033 -422 4060 -358
rect 4124 -422 4588 -358
rect 3963 -424 4588 -422
rect 2195 -488 2261 -482
rect 2321 -483 2387 -482
rect 2321 -488 2322 -483
rect 1358 -547 2322 -488
rect 2386 -488 2387 -483
rect 2386 -547 2513 -488
rect 1042 -548 2513 -547
rect 1042 -609 2513 -608
rect 1042 -668 1167 -609
rect 1166 -673 1167 -668
rect 1231 -668 2194 -609
rect 1231 -673 1232 -668
rect 1166 -674 1232 -673
rect 319 -729 563 -728
rect 319 -734 498 -729
rect -156 -793 498 -734
rect 562 -734 563 -729
rect 1042 -729 1108 -728
rect 1042 -734 1043 -729
rect 562 -793 1043 -734
rect 1107 -734 1108 -729
rect 1107 -793 1232 -734
rect -156 -794 1232 -793
rect -156 -855 1232 -854
rect -156 -914 320 -855
rect 319 -919 320 -914
rect 384 -914 1167 -855
rect 384 -919 563 -914
rect 319 -920 563 -919
rect 1166 -919 1167 -914
rect 1231 -919 1232 -855
rect 1166 -920 1232 -919
rect 1746 -1437 1806 -668
rect 2193 -673 2194 -668
rect 2258 -668 2448 -609
rect 2258 -673 2259 -668
rect 2193 -674 2259 -673
rect 2447 -673 2448 -668
rect 2512 -673 2513 -609
rect 2447 -674 2513 -673
rect 2321 -729 2387 -728
rect 2321 -793 2322 -729
rect 2386 -734 2387 -729
rect 2386 -793 2513 -734
rect 2321 -794 2513 -793
rect 2321 -855 2513 -854
rect 2321 -914 2448 -855
rect 2447 -919 2448 -914
rect 2512 -919 2513 -855
rect 2447 -920 2513 -919
rect 4268 -1350 4588 -424
rect 1743 -1443 1809 -1437
rect 1743 -1507 1744 -1443
rect 1808 -1507 1809 -1443
rect 1743 -1509 1809 -1507
rect 4268 -1540 4288 -1350
rect 4578 -1540 4588 -1350
rect 4268 -1939 4588 -1540
rect 3890 -2060 4588 -1939
rect -686 -2160 -450 -2140
rect -686 -2600 -660 -2160
rect -530 -2600 -450 -2160
rect -686 -2620 -450 -2600
rect 4268 -2335 4588 -2060
rect 4268 -2434 4299 -2335
rect 4567 -2434 4588 -2335
rect 4268 -2700 4588 -2434
rect -686 -2730 -450 -2700
rect -686 -3140 -660 -2730
rect -528 -3140 -450 -2730
rect 3890 -2821 4588 -2700
rect -686 -3170 -450 -3140
rect 4268 -3378 4588 -2821
rect 4658 370 4978 2218
rect 4658 180 4678 370
rect 4958 180 4978 370
rect 4658 -1032 4978 180
rect 4658 -1145 4675 -1032
rect 4967 -1145 4978 -1032
rect 4658 -3378 4978 -1145
<< comment >>
rect 439 -972 443 -585
use adc_comp_buffer  adc_comp_buffer_0
timestamp 1673705348
transform 1 0 2737 0 1 -192
box -42 -306 408 452
use adc_comp_buffer  adc_comp_buffer_1
timestamp 1673705348
transform 1 0 2737 0 -1 -860
box -42 -306 408 452
use adc_noise_decoup_cell2  adc_noise_decoup_cell2_0
timestamp 1663247402
transform 1 0 -450 0 1 -3170
box 0 0 4340 1580
use adc_noise_decoup_cell2  adc_noise_decoup_cell2_1
timestamp 1663247402
transform 1 0 -450 0 1 420
box 0 0 4340 1580
<< labels >>
flabel metal4 s 4658 -3378 4978 2218 0 FreeSans 800 90 0 0 VPWR
port 1 nsew
flabel metal4 s 4268 -3378 4588 2218 0 FreeSans 800 90 0 0 VGND
port 2 nsew
flabel metal1 1272 -469 1318 -427 0 FreeSans 160 180 0 0 bp
flabel metal1 2235 -477 2281 -435 0 FreeSans 160 180 0 0 bn
flabel metal4 1427 -548 1487 -488 0 FreeSans 160 0 0 0 on
flabel metal4 1425 -668 1485 -608 0 FreeSans 160 0 0 0 op
<< end >>
