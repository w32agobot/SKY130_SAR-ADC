* NGSPICE file created from delay_macrocell.ext - technology: sky130A

.subckt delay_macrocell VPWR in out VGND VNB VPB
X0 cap_top VGND sky130_fd_pr__cap_mim_m3_1 l=1.93e+06u w=3.68e+06u
X1 VGND out a_1058_308# VPB sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=7.6e+11p ps=6.7e+06u w=800000u l=150000u
X2 a_1058_308# out VGND VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3 cap_top in VGND VNB sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=2.478e+11p ps=2.86e+06u w=420000u l=4e+06u
X4 cap_top in VPWR VPB sky130_fd_pr__pfet_01v8_lvt ad=2.436e+11p pd=2.26e+06u as=4.836e+11p ps=4.46e+06u w=840000u l=4e+06u
X5 a_1080_80# cap_top VGND VNB sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X6 out cap_top a_1058_308# VPB sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X7 a_1058_308# cap_top VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8 VPWR out a_1080_80# VNB sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X9 cap_top VGND sky130_fd_pr__cap_mim_m3_1 l=1.93e+06u w=2.63e+06u
X10 out cap_top a_1080_80# VNB sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X11 a_1080_80# out VPWR VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

