* NGSPICE file created from adc_clkgen_with_edgedetect.ext - technology: sky130A

.subckt sky130_fd_sc_hd__decap_4 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=4.524e+11p pd=4.52e+06u as=0p ps=0u w=870000u l=1.05e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=2.86e+11p pd=3.24e+06u as=0p ps=0u w=550000u l=1.05e+06u
.ends

.subckt sky130_fd_sc_hd__inv_2 A Y VPWR VGND VNB VPB
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=5.2e+11p ps=5.04e+06u w=1e+06u l=150000u
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=3.38e+11p pd=3.64e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__mux2_1 VGND VPWR S A1 A0 X VNB VPB
X0 VPWR a_505_21# a_535_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=4.553e+11p pd=4.29e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X1 a_505_21# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X2 a_218_374# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X3 VGND a_505_21# a_439_47# VNB sky130_fd_pr__nfet_01v8 ad=5.155e+11p pd=4.31e+06u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4 a_76_199# A0 a_218_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X5 a_505_21# S VGND VNB sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X6 a_439_47# A0 a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X7 a_535_374# A1 a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_76_199# A1 a_218_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X9 a_218_47# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VPWR VPB VNB
D0 VNB DIODE sky130_fd_pr__diode_pw2nd_05v5 pj=2.64e+06u area=4.347e+11p
.ends

.subckt sky130_fd_sc_hd__or2_1 A X B VGND VPWR VNB VPB
X0 VGND A a_68_297# VNB sky130_fd_pr__nfet_01v8 ad=3.097e+11p pd=3.33e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X1 a_68_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 X a_68_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X3 VPWR A a_150_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=2.915e+11p pd=2.67e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X4 X a_68_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=3.4e+11p pd=2.68e+06u as=0p ps=0u w=1e+06u l=150000u
X5 a_150_297# B a_68_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
.ends

.subckt sky130_mm_sc_hd_dlyPoly5ns VPWR in out VGND VNB VPB
X0 a_851_95# in VGND VNB sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=1.0453e+12p ps=9.52e+06u w=420000u l=3.83e+06u
X1 a_1724_71# a_851_95# VGND VNB sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=0p ps=0u w=420000u l=150000u
X2 VPWR out a_1724_71# VNB sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3 VGND out a_1783_329# VPB sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u
X4 a_1783_329# out VGND VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5 a_1724_71# out VPWR VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VGND a_851_95# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.375e+06u l=2.25e+06u
X7 a_1783_329# a_851_95# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.72e+11p ps=4.38e+06u w=800000u l=150000u
X8 out a_851_95# a_1783_329# VPB sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X9 a_851_95# in VPWR VPB sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.83e+06u
X10 out a_851_95# a_1724_71# VNB sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__decap_3 VPWR VGND VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=4.524e+11p pd=4.52e+06u as=0p ps=0u w=870000u l=590000u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=2.86e+11p pd=3.24e+06u as=0p ps=0u w=550000u l=590000u
.ends

.subckt sky130_fd_sc_hd__and2_1 VPWR VGND X B A VNB VPB
X0 VPWR B a_59_75# VPB sky130_fd_pr__pfet_01v8_hvt ad=4.507e+11p pd=4.18e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X1 X a_59_75# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=4.75e+11p pd=2.95e+06u as=0p ps=0u w=1e+06u l=150000u
X2 VGND B a_145_75# VNB sky130_fd_pr__nfet_01v8 ad=2.236e+11p pd=2.08e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X3 a_59_75# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 X a_59_75# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X5 a_145_75# A a_59_75# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__decap_6 VPWR VGND VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=4.524e+11p pd=4.52e+06u as=0p ps=0u w=870000u l=1.97e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=2.86e+11p pd=3.24e+06u as=0p ps=0u w=550000u l=1.97e+06u
.ends

.subckt sky130_fd_sc_hd__nor2b_1 B_N Y A VGND VPWR VNB VPB
X0 Y a_74_47# a_265_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X1 VPWR B_N a_74_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=3.146e+11p pd=2.78e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X2 a_265_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=3.695e+11p ps=3.79e+06u w=650000u l=150000u
X4 VGND B_N a_74_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X5 VGND a_74_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__decap_8 VPWR VGND VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=4.524e+11p pd=4.52e+06u as=0p ps=0u w=870000u l=2.89e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=2.86e+11p pd=3.24e+06u as=0p ps=0u w=550000u l=2.89e+06u
.ends

.subckt sky130_fd_sc_hd__and2b_1 X A_N B VGND VPWR VNB VPB
X0 VPWR B a_207_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=5.986e+11p pd=5e+06u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X1 X a_207_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X2 a_297_47# a_27_413# a_207_413# VNB sky130_fd_pr__nfet_01v8 ad=1.008e+11p pd=1.32e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X3 X a_207_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=3.118e+11p ps=3.34e+06u w=650000u l=150000u
X4 a_207_413# a_27_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VPWR A_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X6 VGND B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_27_413# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__buf_1 VGND VPWR X A VNB VPB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=2.291e+11p pd=2.16e+06u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X1 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=1.508e+11p ps=1.62e+06u w=520000u l=150000u
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X3 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
.ends

.subckt sky130_fd_sc_hd__dlymetal6s6s_1 VPWR VGND A X VNB VPB
X0 X a_629_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=5.82e+11p ps=5.85e+06u w=650000u l=150000u
X1 a_523_47# a_346_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X2 VGND a_240_47# a_346_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X3 a_240_47# a_63_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X4 VPWR a_240_47# a_346_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=8.445e+11p pd=7.95e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X5 VGND A a_63_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X6 VPWR A a_63_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X7 VPWR a_523_47# a_629_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X8 VGND a_523_47# a_629_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X9 a_523_47# a_346_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X10 a_240_47# a_63_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X11 X a_629_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__buf_4 VPWR VGND X A VNB VPB
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=8e+11p pd=7.6e+06u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=5.2e+11p ps=5.5e+06u w=650000u l=150000u
X5 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X9 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
.ends

.subckt adc_clkgen_with_edgedetect VGND VPWR clk_comp_out clk_dig_out dlycontrol1_in[0]
+ dlycontrol1_in[1] dlycontrol1_in[2] dlycontrol1_in[3] dlycontrol1_in[4] dlycontrol2_in[0]
+ dlycontrol2_in[1] dlycontrol2_in[2] dlycontrol2_in[3] dlycontrol2_in[4] dlycontrol3_in[0]
+ dlycontrol3_in[1] dlycontrol3_in[2] dlycontrol3_in[3] dlycontrol3_in[4] dlycontrol4_in[0]
+ dlycontrol4_in[1] dlycontrol4_in[2] dlycontrol4_in[3] dlycontrol4_in[4] dlycontrol4_in[5]
+ ena_in enable_dlycontrol_in ndecision_finish_in nsample_n_in nsample_n_out nsample_p_in
+ nsample_p_out sample_n_in sample_n_out sample_p_in sample_p_out start_conv_in
XFILLER_7_7 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_2.genblk1\[0\].control_invert dlycontrol2_in[0] clkgen.delay_155ns_2.genblk1\[0\].bypass_enable/B
+ VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_12_32 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_302 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_2.genblk1\[0\].dly_binary.out_mux VGND VPWR clkgen.delay_155ns_2.genblk1\[0\].bypass_enable/X
+ outbuf_1/A clkgen.delay_155ns_2.genblk1\[0\].dly_binary.out_mux/A0 clkgen.delay_155ns_2.genblk1\[0\].dly_binary.out_mux/X
+ VGND VPWR sky130_fd_sc_hd__mux2_1
Xclkgen.delay_155ns_2.genblk1\[2\].dly_binary.out_mux VGND VPWR clkgen.delay_155ns_2.genblk1\[2\].bypass_enable/X
+ clkgen.delay_155ns_2.genblk1\[1\].dly_binary.out_mux/X clkgen.delay_155ns_2.genblk1\[2\].dly_binary.out_mux/A0
+ clkgen.delay_155ns_2.genblk1\[2\].dly_binary.out_mux/X VGND VPWR sky130_fd_sc_hd__mux2_1
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.out_mux VGND VPWR clkgen.delay_155ns_2.genblk1\[4\].bypass_enable/X
+ clkgen.delay_155ns_2.genblk1\[3\].dly_binary.out_mux/X clkgen.delay_155ns_2.genblk1\[4\].dly_binary.out_mux/A0
+ clkgen.nor1/A VGND VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_clkgen.delay_155ns_1.genblk1\[2\].control_invert_A dlycontrol1_in[2] VGND
+ VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_20_275 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xedgedetect.or1 edgedetect.or1/A clkgen.nor1/B_N inbuf_1/X VGND VPWR VGND VPWR sky130_fd_sc_hd__or2_1
Xclkgen.delay_155ns_3.genblk1\[0\].dly_binary.genblk1\[0\].delay_unit VPWR clkgen.delay_155ns_3.genblk1\[0\].dly_binary.and_bypass_switch/X
+ clkgen.delay_155ns_3.genblk1\[0\].dly_binary.out_mux/A0 VGND VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_19_183 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xedgedetect.dly_315ns_1.genblk1\[1\].bypass_enable VPWR VGND edgedetect.dly_315ns_1.genblk1\[1\].bypass_enable/X
+ edgedetect.dly_315ns_1.genblk1\[1\].bypass_enable/B edgedetect.dly_315ns_1.enablebuffer/X
+ VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_3_282 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_315 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_164 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_230 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.delay_155ns_2.genblk1\[1\].control_invert_A dlycontrol2_in[1] VGND
+ VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit VPWR clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit/in
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_10_307 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.delay_155ns_2.genblk1\[1\].dly_binary.and_bypass_switch_A_N clkgen.delay_155ns_2.genblk1\[1\].bypass_enable/X
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_1.genblk1\[2\].bypass_enable VPWR VGND clkgen.delay_155ns_1.genblk1\[2\].bypass_enable/X
+ clkgen.delay_155ns_1.genblk1\[2\].bypass_enable/B clkgen.delay_155ns_1.enablebuffer/X
+ VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_2_314 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xclkgen.delay_155ns_2.genblk1\[3\].bypass_enable VPWR VGND clkgen.delay_155ns_2.genblk1\[3\].bypass_enable/X
+ clkgen.delay_155ns_2.genblk1\[3\].bypass_enable/B clkgen.delay_155ns_2.enablebuffer/X
+ VGND VPWR sky130_fd_sc_hd__and2_1
Xclkgen.delay_155ns_3.genblk1\[4\].bypass_enable VPWR VGND clkgen.delay_155ns_3.genblk1\[4\].bypass_enable/X
+ clkgen.delay_155ns_3.genblk1\[4\].bypass_enable/B clkgen.delay_155ns_3.enablebuffer/X
+ VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_15_229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.delay_155ns_3.genblk1\[0\].control_invert_A dlycontrol3_in[0] VGND
+ VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[3\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[3\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[4\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_sampledly04_A nsample_n_in VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_18_32 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_276 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_214 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit VPWR clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit/in
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[2\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[1\].control_invert dlycontrol4_in[1] edgedetect.dly_315ns_1.genblk1\[1\].bypass_enable/B
+ VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_3_294 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_275 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[8\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[8\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[9\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_9_106 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA_clkgen.delay_155ns_1.genblk1\[4\].dly_binary.and_bypass_switch_A_N clkgen.delay_155ns_1.genblk1\[4\].bypass_enable/X
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit VPWR clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit/in
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit VPWR clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit/in
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_5_120 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_175 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_274 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xedgedetect.nor1 inbuf_2/X edgedetect.or1/A edgedetect.nor1/A VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__nor2b_1
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[0\].delay_unit VPWR clkgen.delay_155ns_2.genblk1\[4\].dly_binary.and_bypass_switch/X
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_19_174 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[1\].control_invert dlycontrol3_in[1] clkgen.delay_155ns_3.genblk1\[1\].bypass_enable/B
+ VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_13_125 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_90 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit VPWR clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit/in
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_18_206 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit VPWR clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit/in
+ clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_5_110 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_143 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_187 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_124 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[10\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[9\].delay_unit/out
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[11\].delay_unit/in VGND
+ VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_11_234 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[10\].delay_unit VPWR clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit/out
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_edgedetect.dly_315ns_1.genblk1\[5\].bypass_enable_A edgedetect.dly_315ns_1.enablebuffer/X
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit/in VGND
+ VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit VPWR clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit/in
+ clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_0_244 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_211 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_288 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit VPWR clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit/in
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.and_bypass_switch_A_N edgedetect.dly_315ns_1.genblk1\[3\].bypass_enable/X
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[0\].delay_unit VPWR clkgen.delay_155ns_2.genblk1\[3\].dly_binary.and_bypass_switch/X
+ clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit VPWR clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit/in
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.out_mux/A0 VGND VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[15\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[15\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[16\].delay_unit/in VGND
+ VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_5_133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.nor1 clkgen.nor1/B_N clkgen.nor1/Y clkgen.nor1/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2b_1
XANTENNA_sampledly02_A sample_n_in VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit VPWR clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit/in
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit/out VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_1_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit VPWR clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit/in
+ clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_6_16 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_187 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_7 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_231 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[2\].dly_binary.genblk1\[1\].delay_unit VPWR clkgen.delay_155ns_3.genblk1\[2\].dly_binary.genblk1\[1\].delay_unit/in
+ clkgen.delay_155ns_3.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_1.genblk1\[2\].control_invert dlycontrol1_in[2] clkgen.delay_155ns_1.genblk1\[2\].bypass_enable/B
+ VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[22\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[22\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[23\].delay_unit/in VGND
+ VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_5_315 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_164 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA_edgedetect.dly_315ns_1.enablebuffer_A enable_dlycontrol_in VGND VPWR VPWR
+ VGND sky130_fd_sc_hd__diode_2
XFILLER_20_214 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_192 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[27\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[27\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[28\].delay_unit/in VGND
+ VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_clkgen.delay_155ns_1.genblk1\[1\].control_invert_A dlycontrol1_in[1] VGND
+ VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit VPWR clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit/in
+ clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_1_3 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkgen.delay_155ns_2.enablebuffer_A enable_dlycontrol_in VGND VPWR VPWR VGND
+ sky130_fd_sc_hd__diode_2
XANTENNA_inbuf_3_A ndecision_finish_in VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_20_59 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_317 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xclkgen.delay_155ns_2.genblk1\[2\].dly_binary.genblk1\[0\].delay_unit VPWR clkgen.delay_155ns_2.genblk1\[2\].dly_binary.and_bypass_switch/X
+ clkgen.delay_155ns_2.genblk1\[2\].dly_binary.genblk1\[1\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_19_144 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.clkdig_inverter clkgen.clkdig_inverter/A outbuf_1/A VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_3_243 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_276 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_191 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_0 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkgen.delay_155ns_2.genblk1\[0\].control_invert_A dlycontrol2_in[0] VGND
+ VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_2_308 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.out_mux/A0 VGND VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_4_94 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit VPWR clkgen.delay_155ns_3.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit/in
+ clkgen.delay_155ns_3.genblk1\[1\].dly_binary.out_mux/A0 VGND VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_18_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_315 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_307 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_288 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.delay_155ns_1.genblk1\[4\].dly_binary.out_mux_S clkgen.delay_155ns_1.genblk1\[4\].bypass_enable/X
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_16_148 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xedgedetect.dly_315ns_1.genblk1\[0\].dly_binary.out_mux VGND VPWR edgedetect.dly_315ns_1.genblk1\[0\].bypass_enable/X
+ inbuf_2/X edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.out_mux/A0 edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.out_mux/X
+ VGND VPWR sky130_fd_sc_hd__mux2_1
XPHY_1 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA_edgedetect.dly_315ns_1.genblk1\[0\].bypass_enable_A edgedetect.dly_315ns_1.enablebuffer/X
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xedgedetect.dly_315ns_1.genblk1\[2\].dly_binary.out_mux VGND VPWR edgedetect.dly_315ns_1.genblk1\[2\].bypass_enable/X
+ edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.out_mux/X edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.out_mux/A0
+ edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.out_mux/X VGND VPWR sky130_fd_sc_hd__mux2_1
Xedgedetect.dly_315ns_1.genblk1\[0\].dly_binary.and_bypass_switch edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.and_bypass_switch/X
+ edgedetect.dly_315ns_1.genblk1\[0\].bypass_enable/X inbuf_2/X VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__and2b_1
XFILLER_5_306 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xinbuf_1 VGND VPWR inbuf_1/X ena_in VGND VPWR sky130_fd_sc_hd__buf_1
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.out_mux VGND VPWR edgedetect.dly_315ns_1.genblk1\[4\].bypass_enable/X
+ edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.out_mux/X edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.out_mux/A0
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.out_mux/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_17_276 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_243 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xsampledly31 VPWR VGND sampledly31/A outbuf_3/A VGND VPWR sky130_fd_sc_hd__dlymetal6s6s_1
Xclkgen.delay_155ns_2.genblk1\[1\].dly_binary.genblk1\[0\].delay_unit VPWR clkgen.delay_155ns_2.genblk1\[1\].dly_binary.and_bypass_switch/X
+ clkgen.delay_155ns_2.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_4_62 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_183 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_227 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[2\].bypass_enable VPWR VGND edgedetect.dly_315ns_1.genblk1\[2\].bypass_enable/X
+ edgedetect.dly_315ns_1.genblk1\[2\].bypass_enable/B edgedetect.dly_315ns_1.enablebuffer/X
+ VGND VPWR sky130_fd_sc_hd__and2_1
Xclkgen.delay_155ns_2.genblk1\[3\].control_invert dlycontrol2_in[3] clkgen.delay_155ns_2.genblk1\[3\].bypass_enable/B
+ VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_6_275 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_63 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[10\].delay_unit VPWR clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit/out
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_10_94 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_212 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_116 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_2 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xclkgen.delay_155ns_1.genblk1\[3\].bypass_enable VPWR VGND clkgen.delay_155ns_1.genblk1\[3\].bypass_enable/X
+ clkgen.delay_155ns_1.genblk1\[3\].bypass_enable/B clkgen.delay_155ns_1.enablebuffer/X
+ VGND VPWR sky130_fd_sc_hd__and2_1
Xclkgen.delay_155ns_2.genblk1\[4\].bypass_enable VPWR VGND clkgen.delay_155ns_2.genblk1\[4\].bypass_enable/X
+ clkgen.delay_155ns_2.genblk1\[4\].bypass_enable/B clkgen.delay_155ns_2.enablebuffer/X
+ VGND VPWR sky130_fd_sc_hd__and2_1
Xinbuf_2 VGND VPWR inbuf_2/X start_conv_in VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_12_174 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit VPWR clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit/in
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.out_mux/A0 VGND VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
Xsampledly21 VPWR VGND sampledly21/A sampledly31/A VGND VPWR sky130_fd_sc_hd__dlymetal6s6s_1
Xsampledly32 VPWR VGND sampledly32/A outbuf_4/A VGND VPWR sky130_fd_sc_hd__dlymetal6s6s_1
Xclkgen.delay_155ns_1.genblk1\[0\].dly_binary.out_mux VGND VPWR clkgen.delay_155ns_1.genblk1\[0\].bypass_enable/X
+ inbuf_3/X clkgen.delay_155ns_1.genblk1\[0\].dly_binary.out_mux/A0 clkgen.delay_155ns_1.genblk1\[0\].dly_binary.out_mux/X
+ VGND VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_outbuf_2_A outbuf_2/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_1.genblk1\[2\].dly_binary.out_mux VGND VPWR clkgen.delay_155ns_1.genblk1\[2\].bypass_enable/X
+ clkgen.delay_155ns_1.genblk1\[1\].dly_binary.out_mux/X clkgen.delay_155ns_1.genblk1\[2\].dly_binary.out_mux/A0
+ clkgen.delay_155ns_1.genblk1\[2\].dly_binary.out_mux/X VGND VPWR sky130_fd_sc_hd__mux2_1
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.out_mux VGND VPWR clkgen.delay_155ns_1.genblk1\[4\].bypass_enable/X
+ clkgen.delay_155ns_1.genblk1\[3\].dly_binary.out_mux/X clkgen.delay_155ns_1.genblk1\[4\].dly_binary.out_mux/A0
+ clkgen.clkdig_inverter/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_1_31 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[1\].dly_binary.and_bypass_switch edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.and_bypass_switch/X
+ edgedetect.dly_315ns_1.genblk1\[1\].bypass_enable/X edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.out_mux/X
+ VGND VPWR VGND VPWR sky130_fd_sc_hd__and2b_1
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[4\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[4\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[5\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_inbuf_1_A ena_in VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_19_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_290 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_106 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[2\].delay_unit VPWR clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[2\].delay_unit/in
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_2.genblk1\[0\].dly_binary.genblk1\[0\].delay_unit VPWR clkgen.delay_155ns_2.genblk1\[0\].dly_binary.and_bypass_switch/X
+ clkgen.delay_155ns_2.genblk1\[0\].dly_binary.out_mux/A0 VGND VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_15_183 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_3 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xinbuf_3 VGND VPWR inbuf_3/X ndecision_finish_in VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_12_19 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_124 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_edgedetect.dly_315ns_1.genblk1\[5\].control_invert_A dlycontrol4_in[5] VGND
+ VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xsampledly33 VPWR VGND sampledly33/A outbuf_5/A VGND VPWR sky130_fd_sc_hd__dlymetal6s6s_1
Xsampledly11 VPWR VGND sampledly11/A sampledly21/A VGND VPWR sky130_fd_sc_hd__dlymetal6s6s_1
Xedgedetect.dly_315ns_1.genblk1\[4\].control_invert dlycontrol4_in[4] edgedetect.dly_315ns_1.genblk1\[4\].bypass_enable/B
+ VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
Xsampledly22 VPWR VGND sampledly22/A sampledly32/A VGND VPWR sky130_fd_sc_hd__dlymetal6s6s_1
XANTENNA_clkgen.delay_155ns_1.genblk1\[0\].dly_binary.out_mux_S clkgen.delay_155ns_1.genblk1\[0\].bypass_enable/X
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_1_311 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[9\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[9\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[9\].delay_unit/out VGND
+ VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_14_204 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.delay_155ns_2.genblk1\[0\].dly_binary.and_bypass_switch_B outbuf_1/A
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_20_218 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_218 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit VPWR clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit/in
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit VPWR clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit/in
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_19_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit VPWR clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit/in
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[2\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_3_203 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[0\].bypass_enable VPWR VGND clkgen.delay_155ns_3.genblk1\[0\].bypass_enable/X
+ clkgen.delay_155ns_3.genblk1\[0\].bypass_enable/B clkgen.delay_155ns_3.enablebuffer/X
+ VGND VPWR sky130_fd_sc_hd__and2_1
Xclkgen.delay_155ns_3.genblk1\[1\].dly_binary.out_mux VGND VPWR clkgen.delay_155ns_3.genblk1\[1\].bypass_enable/X
+ clkgen.delay_155ns_3.genblk1\[0\].dly_binary.out_mux/X clkgen.delay_155ns_3.genblk1\[1\].dly_binary.out_mux/A0
+ clkgen.delay_155ns_3.genblk1\[1\].dly_binary.out_mux/X VGND VPWR sky130_fd_sc_hd__mux2_1
XPHY_4 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_20 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[3\].dly_binary.out_mux VGND VPWR clkgen.delay_155ns_3.genblk1\[3\].bypass_enable/X
+ clkgen.delay_155ns_3.genblk1\[2\].dly_binary.out_mux/X clkgen.delay_155ns_3.genblk1\[3\].dly_binary.out_mux/A0
+ clkgen.delay_155ns_3.genblk1\[3\].dly_binary.out_mux/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_1_301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xsampledly23 VPWR VGND sampledly23/A sampledly33/A VGND VPWR sky130_fd_sc_hd__dlymetal6s6s_1
Xsampledly01 VPWR VGND sample_p_in sampledly11/A VGND VPWR sky130_fd_sc_hd__dlymetal6s6s_1
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_3.genblk1\[4\].control_invert dlycontrol3_in[4] clkgen.delay_155ns_3.genblk1\[4\].bypass_enable/B
+ VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
Xsampledly34 VPWR VGND sampledly34/A outbuf_6/A VGND VPWR sky130_fd_sc_hd__dlymetal6s6s_1
XFILLER_4_32 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xsampledly12 VPWR VGND sampledly12/A sampledly22/A VGND VPWR sky130_fd_sc_hd__dlymetal6s6s_1
XFILLER_13_63 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit VPWR clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit/in
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[2\].dly_binary.and_bypass_switch edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.and_bypass_switch/X
+ edgedetect.dly_315ns_1.genblk1\[2\].bypass_enable/X edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.out_mux/X
+ VGND VPWR VGND VPWR sky130_fd_sc_hd__and2b_1
Xclkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit VPWR clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit/in
+ clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_10_274 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[0\].delay_unit VPWR clkgen.delay_155ns_1.genblk1\[4\].dly_binary.and_bypass_switch/X
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_clkgen.delay_155ns_1.genblk1\[0\].control_invert_A dlycontrol1_in[0] VGND
+ VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_3_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_3 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_270 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[11\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[11\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[12\].delay_unit/in VGND
+ VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit VPWR clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit/in
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit/out VGND
+ VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
XPHY_5 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xclkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit VPWR clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit/in
+ clkgen.delay_155ns_3.genblk1\[3\].dly_binary.out_mux/A0 VGND VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit/in VGND
+ VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_17_214 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit VPWR clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit/in
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
Xsampledly13 VPWR VGND sampledly13/A sampledly23/A VGND VPWR sky130_fd_sc_hd__dlymetal6s6s_1
Xsampledly24 VPWR VGND sampledly24/A sampledly34/A VGND VPWR sky130_fd_sc_hd__dlymetal6s6s_1
Xsampledly02 VPWR VGND sample_n_in sampledly12/A VGND VPWR sky130_fd_sc_hd__dlymetal6s6s_1
Xclkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit VPWR clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit/in
+ clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_9_276 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_176 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[16\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[16\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[17\].delay_unit/in VGND
+ VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.and_bypass_switch_A_N edgedetect.dly_315ns_1.genblk1\[1\].bypass_enable/X
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_19_63 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_87 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_43 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.delay_155ns_2.genblk1\[2\].dly_binary.out_mux_S clkgen.delay_155ns_2.genblk1\[2\].bypass_enable/X
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_1.genblk1\[0\].control_invert dlycontrol1_in[0] clkgen.delay_155ns_1.genblk1\[0\].bypass_enable/B
+ VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
Xedgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XPHY_6 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xclkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit VPWR clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit/in
+ clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_12_167 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit VPWR clkgen.delay_155ns_3.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit/in
+ clkgen.delay_155ns_3.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[23\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[23\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[24\].delay_unit/in VGND
+ VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[3\].dly_binary.and_bypass_switch edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.and_bypass_switch/X
+ edgedetect.dly_315ns_1.genblk1\[3\].bypass_enable/X edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.out_mux/X
+ VGND VPWR VGND VPWR sky130_fd_sc_hd__and2b_1
XANTENNA_edgedetect.dly_315ns_1.genblk1\[3\].bypass_enable_A edgedetect.dly_315ns_1.enablebuffer/X
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xsampledly03 VPWR VGND nsample_p_in sampledly13/A VGND VPWR sky130_fd_sc_hd__dlymetal6s6s_1
Xsampledly14 VPWR VGND sampledly14/A sampledly24/A VGND VPWR sky130_fd_sc_hd__dlymetal6s6s_1
Xclkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[0\].delay_unit VPWR clkgen.delay_155ns_1.genblk1\[3\].dly_binary.and_bypass_switch/X
+ clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_4_152 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_174 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_76 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_3 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_199 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_166 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.out_mux_S edgedetect.dly_315ns_1.genblk1\[4\].bypass_enable/X
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_19_31 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[28\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[28\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[29\].delay_unit/in VGND
+ VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit VPWR clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit/in
+ clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_15_154 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[30\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[30\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[31\].delay_unit/in VGND
+ VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
XPHY_7 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xclkgen.delay_155ns_2.genblk1\[2\].dly_binary.genblk1\[1\].delay_unit VPWR clkgen.delay_155ns_2.genblk1\[2\].dly_binary.genblk1\[1\].delay_unit/in
+ clkgen.delay_155ns_2.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_12_124 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_183 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xsampledly04 VPWR VGND nsample_n_in sampledly14/A VGND VPWR sky130_fd_sc_hd__dlymetal6s6s_1
XFILLER_4_142 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_164 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_200 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_56 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_240 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_284 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.enablebuffer VPWR VGND edgedetect.dly_315ns_1.enablebuffer/X
+ enable_dlycontrol_in VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_12_317 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA_edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.out_mux_S edgedetect.dly_315ns_1.genblk1\[2\].bypass_enable/X
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_1.genblk1\[2\].dly_binary.genblk1\[0\].delay_unit VPWR clkgen.delay_155ns_1.genblk1\[2\].dly_binary.and_bypass_switch/X
+ clkgen.delay_155ns_1.genblk1\[2\].dly_binary.genblk1\[1\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.and_bypass_switch edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.and_bypass_switch/X
+ edgedetect.dly_315ns_1.genblk1\[4\].bypass_enable/X edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.out_mux/X
+ VGND VPWR VGND VPWR sky130_fd_sc_hd__and2b_1
XFILLER_16_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_8 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA_edgedetect.dly_315ns_1.genblk1\[4\].control_invert_A dlycontrol4_in[4] VGND
+ VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_1.enablebuffer VPWR VGND clkgen.delay_155ns_1.enablebuffer/X enable_dlycontrol_in
+ VGND VPWR sky130_fd_sc_hd__buf_4
Xedgedetect.dly_315ns_1.genblk1\[3\].bypass_enable VPWR VGND edgedetect.dly_315ns_1.genblk1\[3\].bypass_enable/X
+ edgedetect.dly_315ns_1.genblk1\[3\].bypass_enable/B edgedetect.dly_315ns_1.enablebuffer/X
+ VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_10_245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_2.genblk1\[1\].control_invert dlycontrol2_in[1] clkgen.delay_155ns_2.genblk1\[1\].bypass_enable/B
+ VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
Xclkgen.delay_155ns_2.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit VPWR clkgen.delay_155ns_2.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit/in
+ clkgen.delay_155ns_2.genblk1\[1\].dly_binary.out_mux/A0 VGND VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_15_315 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_219 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_164 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_252 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_296 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[4\].bypass_enable VPWR VGND clkgen.delay_155ns_1.genblk1\[4\].bypass_enable/X
+ clkgen.delay_155ns_1.genblk1\[4\].bypass_enable/B clkgen.delay_155ns_1.enablebuffer/X
+ VGND VPWR sky130_fd_sc_hd__and2_1
Xclkgen.delay_155ns_3.genblk1\[0\].dly_binary.and_bypass_switch clkgen.delay_155ns_3.genblk1\[0\].dly_binary.and_bypass_switch/X
+ clkgen.delay_155ns_3.genblk1\[0\].bypass_enable/X clkgen.nor1/Y VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__and2b_1
XPHY_9 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit VPWR clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit/in
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_clkgen.delay_155ns_1.enablebuffer_A enable_dlycontrol_in VGND VPWR VPWR VGND
+ sky130_fd_sc_hd__diode_2
XANTENNA_edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.out_mux_S edgedetect.dly_315ns_1.genblk1\[0\].bypass_enable/X
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_clkgen.delay_155ns_1.genblk1\[4\].dly_binary.out_mux_A0 clkgen.delay_155ns_1.genblk1\[4\].dly_binary.out_mux/A0
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_4_314 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA_clkgen.delay_155ns_2.genblk1\[2\].dly_binary.and_bypass_switch_A_N clkgen.delay_155ns_2.genblk1\[2\].bypass_enable/X
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[0\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.and_bypass_switch/X
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[1\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_13_276 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xclkgen.delay_155ns_1.genblk1\[1\].dly_binary.genblk1\[0\].delay_unit VPWR clkgen.delay_155ns_1.genblk1\[1\].dly_binary.and_bypass_switch/X
+ clkgen.delay_155ns_1.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_6_3 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.and_bypass_switch edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.and_bypass_switch/X
+ edgedetect.dly_315ns_1.genblk1\[5\].bypass_enable/X edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.out_mux/X
+ VGND VPWR VGND VPWR sky130_fd_sc_hd__and2b_1
XFILLER_2_264 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[5\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[5\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[6\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_7_120 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[2\].control_invert dlycontrol4_in[2] edgedetect.dly_315ns_1.genblk1\[2\].bypass_enable/B
+ VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit VPWR clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit/in
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_1_307 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_274 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_16 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_36 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_192 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_2.genblk1\[0\].bypass_enable VPWR VGND clkgen.delay_155ns_2.genblk1\[0\].bypass_enable/X
+ clkgen.delay_155ns_2.genblk1\[0\].bypass_enable/B clkgen.delay_155ns_2.enablebuffer/X
+ VGND VPWR sky130_fd_sc_hd__and2_1
Xclkgen.delay_155ns_3.genblk1\[1\].bypass_enable VPWR VGND clkgen.delay_155ns_3.genblk1\[1\].bypass_enable/X
+ clkgen.delay_155ns_3.genblk1\[1\].bypass_enable/B clkgen.delay_155ns_3.enablebuffer/X
+ VGND VPWR sky130_fd_sc_hd__and2_1
Xclkgen.delay_155ns_3.genblk1\[1\].dly_binary.and_bypass_switch clkgen.delay_155ns_3.genblk1\[1\].dly_binary.and_bypass_switch/X
+ clkgen.delay_155ns_3.genblk1\[1\].bypass_enable/X clkgen.delay_155ns_3.genblk1\[0\].dly_binary.out_mux/X
+ VGND VPWR VGND VPWR sky130_fd_sc_hd__and2b_1
XFILLER_2_276 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkgen.delay_155ns_3.genblk1\[4\].control_invert_A dlycontrol3_in[4] VGND
+ VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit VPWR clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit/in
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_15_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit VPWR clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit/in
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_2.genblk1\[0\].dly_binary.and_bypass_switch clkgen.delay_155ns_2.genblk1\[0\].dly_binary.and_bypass_switch/X
+ clkgen.delay_155ns_2.genblk1\[0\].bypass_enable/X outbuf_1/A VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__and2b_1
XFILLER_7_49 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[0\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.and_bypass_switch/X
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[2\].delay_unit VPWR clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[2\].delay_unit/in
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_14_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_154 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[0\].dly_binary.genblk1\[0\].delay_unit VPWR clkgen.delay_155ns_1.genblk1\[0\].dly_binary.and_bypass_switch/X
+ clkgen.delay_155ns_1.genblk1\[0\].dly_binary.out_mux/A0 VGND VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_clkgen.delay_155ns_1.genblk1\[0\].dly_binary.and_bypass_switch_A_N clkgen.delay_155ns_1.genblk1\[0\].bypass_enable/X
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_4_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[2\].control_invert dlycontrol3_in[2] clkgen.delay_155ns_3.genblk1\[2\].bypass_enable/B
+ VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_13_59 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_216 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_271 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_182 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_10_16 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit VPWR clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit/in
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_2_200 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_222 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit VPWR clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit/in
+ clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_2_94 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit VPWR clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit/in
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[2\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_16_59 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[12\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[12\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[13\].delay_unit/in VGND
+ VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_2.genblk1\[1\].dly_binary.out_mux VGND VPWR clkgen.delay_155ns_2.genblk1\[1\].bypass_enable/X
+ clkgen.delay_155ns_2.genblk1\[0\].dly_binary.out_mux/X clkgen.delay_155ns_2.genblk1\[1\].dly_binary.out_mux/A0
+ clkgen.delay_155ns_2.genblk1\[1\].dly_binary.out_mux/X VGND VPWR sky130_fd_sc_hd__mux2_1
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit VPWR clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit/in
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_2.genblk1\[3\].dly_binary.out_mux VGND VPWR clkgen.delay_155ns_2.genblk1\[3\].bypass_enable/X
+ clkgen.delay_155ns_2.genblk1\[2\].dly_binary.out_mux/X clkgen.delay_155ns_2.genblk1\[3\].dly_binary.out_mux/A0
+ clkgen.delay_155ns_2.genblk1\[3\].dly_binary.out_mux/X VGND VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.and_bypass_switch_A_N edgedetect.dly_315ns_1.genblk1\[4\].bypass_enable/X
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_13_49 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[2\].dly_binary.and_bypass_switch clkgen.delay_155ns_3.genblk1\[2\].dly_binary.and_bypass_switch/X
+ clkgen.delay_155ns_3.genblk1\[2\].bypass_enable/X clkgen.delay_155ns_3.genblk1\[1\].dly_binary.out_mux/X
+ VGND VPWR VGND VPWR sky130_fd_sc_hd__and2b_1
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit/in VGND
+ VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_18_316 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[0\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.and_bypass_switch/X
+ edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_2.genblk1\[1\].dly_binary.and_bypass_switch clkgen.delay_155ns_2.genblk1\[1\].dly_binary.and_bypass_switch/X
+ clkgen.delay_155ns_2.genblk1\[1\].bypass_enable/X clkgen.delay_155ns_2.genblk1\[0\].dly_binary.out_mux/X
+ VGND VPWR VGND VPWR sky130_fd_sc_hd__and2b_1
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit VPWR clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit/in
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit VPWR clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit/in
+ clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_2_234 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_124 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[17\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[17\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[18\].delay_unit/in VGND
+ VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_1.genblk1\[0\].dly_binary.and_bypass_switch clkgen.delay_155ns_1.genblk1\[0\].dly_binary.and_bypass_switch/X
+ clkgen.delay_155ns_1.genblk1\[0\].bypass_enable/X inbuf_3/X VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__and2b_1
XFILLER_11_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_315 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_16 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_152 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_94 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit VPWR clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit/in
+ clkgen.delay_155ns_2.genblk1\[3\].dly_binary.out_mux/A0 VGND VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_1.genblk1\[3\].control_invert dlycontrol1_in[3] clkgen.delay_155ns_1.genblk1\[3\].bypass_enable/B
+ VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XANTENNA_edgedetect.dly_315ns_1.genblk1\[3\].control_invert_A dlycontrol4_in[3] VGND
+ VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_13_214 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xclkgen.delay_155ns_3.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit VPWR clkgen.delay_155ns_3.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit/in
+ clkgen.delay_155ns_3.genblk1\[2\].dly_binary.out_mux/A0 VGND VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_0_173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[24\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[24\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[25\].delay_unit/in VGND
+ VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_8_284 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
Xclkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit VPWR clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit/in
+ clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_5_276 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_246 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[29\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[29\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[30\].delay_unit/in VGND
+ VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[2\].dly_binary.genblk1\[0\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.and_bypass_switch/X
+ edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.genblk1\[1\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_3.genblk1\[3\].dly_binary.and_bypass_switch clkgen.delay_155ns_3.genblk1\[3\].dly_binary.and_bypass_switch/X
+ clkgen.delay_155ns_3.genblk1\[3\].bypass_enable/X clkgen.delay_155ns_3.genblk1\[2\].dly_binary.out_mux/X
+ VGND VPWR VGND VPWR sky130_fd_sc_hd__and2b_1
Xclkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit VPWR clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit/in
+ clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_17_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_212 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[31\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[31\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.out_mux/A0 VGND VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_2.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit VPWR clkgen.delay_155ns_2.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit/in
+ clkgen.delay_155ns_2.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_0_300 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_3 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xclkgen.delay_155ns_2.genblk1\[2\].dly_binary.and_bypass_switch clkgen.delay_155ns_2.genblk1\[2\].dly_binary.and_bypass_switch/X
+ clkgen.delay_155ns_2.genblk1\[2\].bypass_enable/X clkgen.delay_155ns_2.genblk1\[1\].dly_binary.out_mux/X
+ VGND VPWR VGND VPWR sky130_fd_sc_hd__and2b_1
XFILLER_0_152 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_252 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_63 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[1\].dly_binary.and_bypass_switch clkgen.delay_155ns_1.genblk1\[1\].dly_binary.and_bypass_switch/X
+ clkgen.delay_155ns_1.genblk1\[1\].bypass_enable/X clkgen.delay_155ns_1.genblk1\[0\].dly_binary.out_mux/X
+ VGND VPWR VGND VPWR sky130_fd_sc_hd__and2b_1
XFILLER_14_94 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_244 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_edgedetect.dly_315ns_1.genblk1\[1\].bypass_enable_A edgedetect.dly_315ns_1.enablebuffer/X
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_2_214 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_258 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_84 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_195 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sampledly03_A nsample_p_in VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_20_121 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_276 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_187 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[2\].dly_binary.genblk1\[1\].delay_unit VPWR clkgen.delay_155ns_1.genblk1\[2\].dly_binary.genblk1\[1\].delay_unit/in
+ clkgen.delay_155ns_1.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[4\].bypass_enable VPWR VGND edgedetect.dly_315ns_1.genblk1\[4\].bypass_enable/X
+ edgedetect.dly_315ns_1.genblk1\[4\].bypass_enable/B edgedetect.dly_315ns_1.enablebuffer/X
+ VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_3_150 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_194 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_164 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_31 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.delay_155ns_2.genblk1\[4\].control_invert_A dlycontrol2_in[4] VGND
+ VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_14_62 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_2.enablebuffer VPWR VGND clkgen.delay_155ns_2.enablebuffer/X enable_dlycontrol_in
+ VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_17_182 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[1\].dly_binary.genblk1\[0\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.and_bypass_switch/X
+ edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_11_30 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.and_bypass_switch clkgen.delay_155ns_3.genblk1\[4\].dly_binary.and_bypass_switch/X
+ clkgen.delay_155ns_3.genblk1\[4\].bypass_enable/X clkgen.delay_155ns_3.genblk1\[3\].dly_binary.out_mux/X
+ VGND VPWR VGND VPWR sky130_fd_sc_hd__and2b_1
XFILLER_11_74 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.delay_155ns_3.genblk1\[3\].control_invert_A dlycontrol3_in[3] VGND
+ VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_2_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.out_mux_A0 edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.out_mux/A0
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_2.genblk1\[4\].control_invert dlycontrol2_in[4] clkgen.delay_155ns_2.genblk1\[4\].bypass_enable/B
+ VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
Xclkgen.delay_155ns_2.genblk1\[3\].dly_binary.and_bypass_switch clkgen.delay_155ns_2.genblk1\[3\].dly_binary.and_bypass_switch/X
+ clkgen.delay_155ns_2.genblk1\[3\].bypass_enable/X clkgen.delay_155ns_2.genblk1\[2\].dly_binary.out_mux/X
+ VGND VPWR VGND VPWR sky130_fd_sc_hd__and2b_1
XFILLER_16_203 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[2\].dly_binary.and_bypass_switch clkgen.delay_155ns_1.genblk1\[2\].dly_binary.and_bypass_switch/X
+ clkgen.delay_155ns_1.genblk1\[2\].bypass_enable/X clkgen.delay_155ns_1.genblk1\[1\].dly_binary.out_mux/X
+ VGND VPWR VGND VPWR sky130_fd_sc_hd__and2b_1
XFILLER_4_107 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit VPWR clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit/in
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_8_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_121 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[1\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[1\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[2\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XPHY_40 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_271 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit VPWR clkgen.delay_155ns_1.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit/in
+ clkgen.delay_155ns_1.genblk1\[1\].dly_binary.out_mux/A0 VGND VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_20_315 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_315 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_164 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_156 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_300 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[0\].control_invert dlycontrol4_in[0] edgedetect.dly_315ns_1.genblk1\[0\].bypass_enable/B
+ VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_17_63 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[6\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[6\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[7\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_1.genblk1\[0\].bypass_enable VPWR VGND clkgen.delay_155ns_1.genblk1\[0\].bypass_enable/X
+ clkgen.delay_155ns_1.genblk1\[0\].bypass_enable/B clkgen.delay_155ns_1.enablebuffer/X
+ VGND VPWR sky130_fd_sc_hd__and2_1
Xedgedetect.dly_315ns_1.genblk1\[0\].dly_binary.genblk1\[0\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.and_bypass_switch/X
+ edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.out_mux/A0 VGND VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_0_199 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_2.genblk1\[1\].bypass_enable VPWR VGND clkgen.delay_155ns_2.genblk1\[1\].bypass_enable/X
+ clkgen.delay_155ns_2.genblk1\[1\].bypass_enable/B clkgen.delay_155ns_2.enablebuffer/X
+ VGND VPWR sky130_fd_sc_hd__and2_1
Xclkgen.delay_155ns_3.genblk1\[2\].bypass_enable VPWR VGND clkgen.delay_155ns_3.genblk1\[2\].bypass_enable/X
+ clkgen.delay_155ns_3.genblk1\[2\].bypass_enable/B clkgen.delay_155ns_3.enablebuffer/X
+ VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_12_284 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_3 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit VPWR clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit/in
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_5_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[10\].delay_unit VPWR clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit/out
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[5\].control_invert dlycontrol4_in[5] edgedetect.dly_315ns_1.genblk1\[5\].bypass_enable/B
+ VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_2_228 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_41 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_30 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_313 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_283 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.and_bypass_switch clkgen.delay_155ns_2.genblk1\[4\].dly_binary.and_bypass_switch/X
+ clkgen.delay_155ns_2.genblk1\[4\].bypass_enable/X clkgen.delay_155ns_2.genblk1\[3\].dly_binary.out_mux/X
+ VGND VPWR VGND VPWR sky130_fd_sc_hd__and2b_1
XANTENNA_clkgen.delay_155ns_1.genblk1\[3\].dly_binary.and_bypass_switch_A_N clkgen.delay_155ns_1.genblk1\[3\].bypass_enable/X
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_1.genblk1\[3\].dly_binary.and_bypass_switch clkgen.delay_155ns_1.genblk1\[3\].dly_binary.and_bypass_switch/X
+ clkgen.delay_155ns_1.genblk1\[3\].bypass_enable/X clkgen.delay_155ns_1.genblk1\[2\].dly_binary.out_mux/X
+ VGND VPWR VGND VPWR sky130_fd_sc_hd__and2b_1
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit VPWR clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit/in
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit/out VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_6_183 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sampledly01_A sample_p_in VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit VPWR clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit/in
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.out_mux/A0 VGND VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_0_315 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[2\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_17_31 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[0\].control_invert dlycontrol3_in[0] clkgen.delay_155ns_3.genblk1\[0\].bypass_enable/B
+ VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit VPWR clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit/in
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_12_252 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_edgedetect.dly_315ns_1.genblk1\[2\].control_invert_A dlycontrol4_in[2] VGND
+ VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_8_223 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_32 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_215 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_207 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_31 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_20 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_306 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_295 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[1\].dly_binary.out_mux VGND VPWR edgedetect.dly_315ns_1.genblk1\[1\].bypass_enable/X
+ edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.out_mux/X edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.out_mux/A0
+ edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.out_mux/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_14_122 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit VPWR clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit/in
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_20_125 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xedgedetect.dly_315ns_1.genblk1\[3\].dly_binary.out_mux VGND VPWR edgedetect.dly_315ns_1.genblk1\[3\].bypass_enable/X
+ edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.out_mux/X edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.out_mux/A0
+ edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.out_mux/X VGND VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_inbuf_2_A start_conv_in VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.out_mux VGND VPWR edgedetect.dly_315ns_1.genblk1\[5\].bypass_enable/X
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.out_mux/X edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.out_mux/A0
+ edgedetect.nor1/A VGND VPWR sky130_fd_sc_hd__mux2_1
Xclkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit VPWR clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit/in
+ clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_0_3 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_280 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[2\].delay_unit VPWR clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[2\].delay_unit/in
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_3_143 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkgen.delay_155ns_1.genblk1\[3\].dly_binary.out_mux_S clkgen.delay_155ns_1.genblk1\[3\].bypass_enable/X
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[13\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[13\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[14\].delay_unit/in VGND
+ VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit VPWR clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit/in
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XPHY_32 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.and_bypass_switch clkgen.delay_155ns_1.genblk1\[4\].dly_binary.and_bypass_switch/X
+ clkgen.delay_155ns_1.genblk1\[4\].bypass_enable/X clkgen.delay_155ns_1.genblk1\[3\].dly_binary.out_mux/X
+ VGND VPWR VGND VPWR sky130_fd_sc_hd__and2b_1
XPHY_10 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit/in VGND
+ VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_17_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.and_bypass_switch_A_N edgedetect.dly_315ns_1.genblk1\[2\].bypass_enable/X
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_1_230 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
Xoutbuf_1 VPWR VGND clk_dig_out outbuf_1/A VGND VPWR sky130_fd_sc_hd__buf_4
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit VPWR clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit/in
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_edgedetect.dly_315ns_1.genblk1\[4\].bypass_enable_A edgedetect.dly_315ns_1.enablebuffer/X
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit VPWR clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit/in
+ clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[18\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[18\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[19\].delay_unit/in VGND
+ VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_clkgen.delay_155ns_1.genblk1\[4\].control_invert_A dlycontrol1_in[4] VGND
+ VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[20\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[20\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[21\].delay_unit/in VGND
+ VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_0_306 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_9 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[1\].control_invert dlycontrol1_in[1] clkgen.delay_155ns_1.genblk1\[1\].bypass_enable/B
+ VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_3_133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[1\].dly_binary.out_mux VGND VPWR clkgen.delay_155ns_1.genblk1\[1\].bypass_enable/X
+ clkgen.delay_155ns_1.genblk1\[0\].dly_binary.out_mux/X clkgen.delay_155ns_1.genblk1\[1\].dly_binary.out_mux/A0
+ clkgen.delay_155ns_1.genblk1\[1\].dly_binary.out_mux/X VGND VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_edgedetect.nor1_B_N inbuf_2/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xedgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_1.genblk1\[3\].dly_binary.out_mux VGND VPWR clkgen.delay_155ns_1.genblk1\[3\].bypass_enable/X
+ clkgen.delay_155ns_1.genblk1\[2\].dly_binary.out_mux/X clkgen.delay_155ns_1.genblk1\[3\].dly_binary.out_mux/A0
+ clkgen.delay_155ns_1.genblk1\[3\].dly_binary.out_mux/X VGND VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_clkgen.delay_155ns_2.genblk1\[3\].control_invert_A dlycontrol2_in[3] VGND
+ VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XPHY_33 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_90 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_242 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_59 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[25\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[25\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[26\].delay_unit/in VGND
+ VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit VPWR clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit/in
+ clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
Xoutbuf_2 VPWR VGND clk_comp_out outbuf_2/A VGND VPWR sky130_fd_sc_hd__buf_4
XANTENNA_clkgen.delay_155ns_3.genblk1\[2\].control_invert_A dlycontrol3_in[2] VGND
+ VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_3_315 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_3 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_171 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_266 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_259 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[2\].dly_binary.genblk1\[1\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.genblk1\[1\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit VPWR clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit/in
+ clkgen.delay_155ns_1.genblk1\[3\].dly_binary.out_mux/A0 VGND VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_2.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit VPWR clkgen.delay_155ns_2.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit/in
+ clkgen.delay_155ns_2.genblk1\[2\].dly_binary.out_mux/A0 VGND VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_4_284 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_12 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_16 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xoutbuf_3 VPWR VGND sample_p_out outbuf_3/A VGND VPWR sky130_fd_sc_hd__buf_4
Xclkgen.delay_155ns_3.genblk1\[0\].dly_binary.out_mux VGND VPWR clkgen.delay_155ns_3.genblk1\[0\].bypass_enable/X
+ clkgen.nor1/Y clkgen.delay_155ns_3.genblk1\[0\].dly_binary.out_mux/A0 clkgen.delay_155ns_3.genblk1\[0\].dly_binary.out_mux/X
+ VGND VPWR sky130_fd_sc_hd__mux2_1
Xclkgen.delay_155ns_3.genblk1\[2\].dly_binary.out_mux VGND VPWR clkgen.delay_155ns_3.genblk1\[2\].bypass_enable/X
+ clkgen.delay_155ns_3.genblk1\[1\].dly_binary.out_mux/X clkgen.delay_155ns_3.genblk1\[2\].dly_binary.out_mux/A0
+ clkgen.delay_155ns_3.genblk1\[2\].dly_binary.out_mux/X VGND VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_outbuf_1_A outbuf_1/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_19_217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].bypass_enable VPWR VGND edgedetect.dly_315ns_1.genblk1\[5\].bypass_enable/X
+ edgedetect.dly_315ns_1.genblk1\[5\].bypass_enable/B edgedetect.dly_315ns_1.enablebuffer/X
+ VGND VPWR sky130_fd_sc_hd__and2_1
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.out_mux VGND VPWR clkgen.delay_155ns_3.genblk1\[4\].bypass_enable/X
+ clkgen.delay_155ns_3.genblk1\[3\].dly_binary.out_mux/X clkgen.delay_155ns_3.genblk1\[4\].dly_binary.out_mux/A0
+ outbuf_2/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_8_59 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_220 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_179 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_212 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit VPWR clkgen.delay_155ns_1.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit/in
+ clkgen.delay_155ns_1.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_20_90 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_315 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_274 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_35 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_307 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_24 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_3 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_13 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xoutbuf_4 VPWR VGND sample_n_out outbuf_4/A VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_13_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.enablebuffer VPWR VGND clkgen.delay_155ns_3.enablebuffer/X enable_dlycontrol_in
+ VGND VPWR sky130_fd_sc_hd__buf_4
Xclkgen.delay_155ns_2.genblk1\[2\].control_invert dlycontrol2_in[2] clkgen.delay_155ns_2.genblk1\[2\].bypass_enable/B
+ VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_3_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.out_mux/A0 VGND VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_8_16 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_306 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.delay_155ns_2.genblk1\[4\].dly_binary.out_mux_A0 clkgen.delay_155ns_2.genblk1\[4\].dly_binary.out_mux/A0
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_15_276 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_191 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_206 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_edgedetect.dly_315ns_1.genblk1\[1\].control_invert_A dlycontrol4_in[1] VGND
+ VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit VPWR clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[13\].delay_unit/in
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_17_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_36 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_212 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_14 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xedgedetect.dly_315ns_1.genblk1\[0\].bypass_enable VPWR VGND edgedetect.dly_315ns_1.genblk1\[0\].bypass_enable/X
+ edgedetect.dly_315ns_1.genblk1\[0\].bypass_enable/B edgedetect.dly_315ns_1.enablebuffer/X
+ VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_1_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xoutbuf_5 VPWR VGND nsample_p_out outbuf_5/A VGND VPWR sky130_fd_sc_hd__buf_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[2\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[2\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[3\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.out_mux_S edgedetect.dly_315ns_1.genblk1\[5\].bypass_enable/X
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.and_bypass_switch_B inbuf_2/X
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_18_274 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[0\].delay_unit VPWR clkgen.delay_155ns_3.genblk1\[4\].dly_binary.and_bypass_switch/X
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[1\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_1.genblk1\[1\].bypass_enable VPWR VGND clkgen.delay_155ns_1.genblk1\[1\].bypass_enable/X
+ clkgen.delay_155ns_1.genblk1\[1\].bypass_enable/B clkgen.delay_155ns_1.enablebuffer/X
+ VGND VPWR sky130_fd_sc_hd__and2_1
Xclkgen.delay_155ns_2.genblk1\[2\].bypass_enable VPWR VGND clkgen.delay_155ns_2.genblk1\[2\].bypass_enable/X
+ clkgen.delay_155ns_2.genblk1\[2\].bypass_enable/B clkgen.delay_155ns_2.enablebuffer/X
+ VGND VPWR sky130_fd_sc_hd__and2_1
XANTENNA_clkgen.delay_155ns_2.genblk1\[1\].dly_binary.out_mux_S clkgen.delay_155ns_2.genblk1\[1\].bypass_enable/X
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_17_3 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xclkgen.delay_155ns_3.genblk1\[3\].bypass_enable VPWR VGND clkgen.delay_155ns_3.genblk1\[3\].bypass_enable/X
+ clkgen.delay_155ns_3.genblk1\[3\].bypass_enable/B clkgen.delay_155ns_3.enablebuffer/X
+ VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_12_203 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[7\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[7\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[8\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_14_16 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[3\].control_invert dlycontrol4_in[3] edgedetect.dly_315ns_1.genblk1\[3\].bypass_enable/B
+ VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XPHY_37 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_94 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_61 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_125 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit VPWR clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit/in
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[6\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_1_224 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit VPWR clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit/in
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[12\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
Xoutbuf_6 VPWR VGND nsample_n_out outbuf_6/A VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_13_172 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_187 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_164 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_124 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.out_mux_S edgedetect.dly_315ns_1.genblk1\[3\].bypass_enable/X
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_15_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkgen.delay_155ns_1.genblk1\[3\].control_invert_A dlycontrol1_in[3] VGND
+ VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_20_292 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_259 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.delay_155ns_2.genblk1\[0\].dly_binary.out_mux_A1 outbuf_1/A VGND VPWR
+ VPWR VGND sky130_fd_sc_hd__diode_2
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[2\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[2\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XPHY_38 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit VPWR clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit/in
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[5\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XPHY_16 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkgen.delay_155ns_2.genblk1\[2\].control_invert_A dlycontrol2_in[2] VGND
+ VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_15_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[0\].delay_unit VPWR clkgen.delay_155ns_3.genblk1\[3\].dly_binary.and_bypass_switch/X
+ clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[1\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_3.genblk1\[3\].control_invert dlycontrol3_in[3] clkgen.delay_155ns_3.genblk1\[3\].bypass_enable/B
+ VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_1_236 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_313 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_317 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkgen.delay_155ns_3.enablebuffer_A enable_dlycontrol_in VGND VPWR VPWR VGND
+ sky130_fd_sc_hd__diode_2
XFILLER_9_155 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_30 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_63 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkgen.delay_155ns_3.genblk1\[1\].control_invert_A dlycontrol3_in[1] VGND
+ VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_12_94 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[7\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit VPWR clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit/in
+ clkgen.delay_155ns_2.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit/out VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_2_161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit VPWR clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit/in
+ clkgen.delay_155ns_3.genblk1\[3\].dly_binary.genblk1\[6\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_edgedetect.dly_315ns_1.genblk1\[1\].dly_binary.out_mux_S edgedetect.dly_315ns_1.genblk1\[1\].bypass_enable/X
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[10\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit/out
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[11\].delay_unit/in VGND
+ VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
XANTENNA_edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.and_bypass_switch_A_N edgedetect.dly_315ns_1.genblk1\[5\].bypass_enable/X
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit VPWR clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[3\].delay_unit/in
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[4\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_4_212 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_28 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_17 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_259 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[14\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[14\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[15\].delay_unit/in VGND
+ VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_9_315 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit VPWR clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[14\].delay_unit/in
+ clkgen.delay_155ns_3.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_6_307 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xedgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.genblk1\[15\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[4\].dly_binary.out_mux/A0 VGND VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_12_62 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[2\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit VPWR clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[8\].delay_unit/in
+ clkgen.delay_155ns_1.genblk1\[4\].dly_binary.genblk1\[9\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit VPWR clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit/in
+ clkgen.delay_155ns_2.genblk1\[3\].dly_binary.genblk1\[5\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_0_32 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA_edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.and_bypass_switch_A_N edgedetect.dly_315ns_1.genblk1\[0\].bypass_enable/X
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xclkgen.delay_155ns_3.genblk1\[2\].dly_binary.genblk1\[0\].delay_unit VPWR clkgen.delay_155ns_3.genblk1\[2\].dly_binary.and_bypass_switch/X
+ clkgen.delay_155ns_3.genblk1\[2\].dly_binary.genblk1\[1\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_9_74 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_94 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[19\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[19\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[20\].delay_unit/in VGND
+ VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_7_243 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[21\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[21\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[22\].delay_unit/in VGND
+ VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_15_3 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_276 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_edgedetect.dly_315ns_1.genblk1\[0\].dly_binary.out_mux_A1 inbuf_2/X VGND
+ VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XPHY_29 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_18 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xedgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.genblk1\[7\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[3\].dly_binary.out_mux/A0 VGND VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_9_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[4\].control_invert dlycontrol1_in[4] clkgen.delay_155ns_1.genblk1\[4\].bypass_enable/B
+ VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_16_194 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[26\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[26\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[5\].dly_binary.genblk1\[27\].delay_unit/in VGND
+ VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
Xclkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit VPWR clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[3\].delay_unit/in
+ clkgen.delay_155ns_1.genblk1\[3\].dly_binary.genblk1\[4\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_9_31 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_62 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_edgedetect.dly_315ns_1.genblk1\[2\].bypass_enable_A edgedetect.dly_315ns_1.enablebuffer/X
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_4_203 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_edgedetect.dly_315ns_1.genblk1\[0\].control_invert_A dlycontrol4_in[0] VGND
+ VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_6_32 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_19 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_206 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xedgedetect.dly_315ns_1.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit VPWR edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.genblk1\[2\].delay_unit/in
+ edgedetect.dly_315ns_1.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_15_63 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_294 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_110 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xclkgen.delay_155ns_3.genblk1\[1\].dly_binary.genblk1\[0\].delay_unit VPWR clkgen.delay_155ns_3.genblk1\[1\].dly_binary.and_bypass_switch/X
+ clkgen.delay_155ns_3.genblk1\[1\].dly_binary.genblk1\[1\].delay_unit/in VGND VGND
+ VPWR sky130_mm_sc_hd_dlyPoly5ns
XFILLER_9_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_124 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_3 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_238 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_241 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_3 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_31 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_218 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkgen.delay_155ns_1.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit VPWR clkgen.delay_155ns_1.genblk1\[2\].dly_binary.genblk1\[3\].delay_unit/in
+ clkgen.delay_155ns_1.genblk1\[2\].dly_binary.out_mux/A0 VGND VGND VPWR sky130_mm_sc_hd_dlyPoly5ns
.ends

