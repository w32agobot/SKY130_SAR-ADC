magic
tech sky130A
timestamp 1661503936
<< nwell >>
rect 0 89 104 243
<< nmos >>
rect 31 11 73 26
<< pmos >>
rect 31 136 73 151
<< ndiff >>
rect 31 49 73 55
rect 31 32 37 49
rect 67 32 73 49
rect 31 26 73 32
rect 31 5 73 11
rect 31 -12 37 5
rect 67 -12 73 5
rect 31 -18 73 -12
<< pdiff >>
rect 31 174 73 180
rect 31 157 37 174
rect 67 157 73 174
rect 31 151 73 157
rect 31 130 73 136
rect 31 113 37 130
rect 67 113 73 130
rect 31 107 73 113
<< ndiffc >>
rect 37 32 67 49
rect 37 -12 67 5
<< pdiffc >>
rect 37 157 67 174
rect 37 113 67 130
<< psubdiff >>
rect 31 -62 43 -45
rect 61 -62 73 -45
rect 31 -65 73 -62
<< nsubdiff >>
rect 31 207 43 225
rect 61 207 73 225
<< psubdiffcont >>
rect 43 -62 61 -45
<< nsubdiffcont >>
rect 43 207 61 225
<< poly >>
rect 8 136 31 151
rect 73 136 86 151
rect 8 94 23 136
rect -13 86 23 94
rect -13 69 -5 86
rect 12 69 23 86
rect -13 61 23 69
rect 8 26 23 61
rect 8 11 31 26
rect 73 11 86 26
<< polycont >>
rect -5 69 12 86
<< locali >>
rect 31 226 43 243
rect 61 226 73 243
rect 31 225 73 226
rect 31 207 43 225
rect 61 207 73 225
rect 31 174 73 207
rect 29 157 37 174
rect 67 157 75 174
rect 29 113 37 130
rect 67 113 75 130
rect -13 86 14 94
rect -13 69 -5 86
rect 12 69 14 86
rect -13 61 14 69
rect 31 89 73 113
rect 31 66 104 89
rect 31 49 73 66
rect 29 32 37 49
rect 67 32 75 49
rect 31 29 73 32
rect 29 -12 37 5
rect 67 -12 75 5
rect 31 -45 73 -12
rect 31 -62 43 -45
rect 61 -62 73 -45
rect 31 -65 73 -62
<< viali >>
rect 43 226 61 243
rect 43 -62 61 -45
<< metal1 >>
rect 27 243 76 246
rect 27 226 43 243
rect 61 226 76 243
rect 27 223 76 226
rect 28 -45 76 -42
rect 28 -62 43 -45
rect 61 -62 76 -45
rect 28 -65 76 -62
<< labels >>
rlabel locali -13 66 -13 89 7 in
rlabel locali 104 66 104 89 3 out
rlabel metal1 27 223 27 246 7 VDD
port 1 w
rlabel metal1 28 -65 28 -42 7 VSS
port 2 w
<< end >>
