magic
tech sky130A
timestamp 1660641620
<< metal2 >>
rect 14 1430 628 1490
rect 14 1402 19 1430
rect 47 1402 83 1430
rect 111 1402 147 1430
rect 175 1402 211 1430
rect 239 1402 275 1430
rect 303 1402 339 1430
rect 367 1402 403 1430
rect 431 1402 467 1430
rect 495 1402 531 1430
rect 559 1402 595 1430
rect 623 1402 628 1430
rect 14 1344 628 1402
rect 14 1316 19 1344
rect 47 1316 83 1344
rect 111 1316 147 1344
rect 175 1316 211 1344
rect 239 1316 275 1344
rect 303 1316 339 1344
rect 367 1316 403 1344
rect 431 1316 467 1344
rect 495 1316 531 1344
rect 559 1316 595 1344
rect 623 1334 628 1344
rect 656 1430 1270 1490
rect 656 1402 661 1430
rect 689 1402 725 1430
rect 753 1402 789 1430
rect 817 1402 853 1430
rect 881 1402 917 1430
rect 945 1402 981 1430
rect 1009 1402 1045 1430
rect 1073 1402 1109 1430
rect 1137 1402 1173 1430
rect 1201 1402 1237 1430
rect 1265 1402 1270 1430
rect 656 1344 1270 1402
rect 656 1334 661 1344
rect 623 1317 661 1334
rect 623 1316 628 1317
rect 14 1258 628 1316
rect 14 1230 19 1258
rect 47 1230 83 1258
rect 111 1230 147 1258
rect 175 1230 211 1258
rect 239 1230 275 1258
rect 303 1230 339 1258
rect 367 1230 403 1258
rect 431 1230 467 1258
rect 495 1230 531 1258
rect 559 1230 595 1258
rect 623 1230 628 1258
rect 14 1170 628 1230
rect 656 1316 661 1317
rect 689 1316 725 1344
rect 753 1316 789 1344
rect 817 1316 853 1344
rect 881 1316 917 1344
rect 945 1316 981 1344
rect 1009 1316 1045 1344
rect 1073 1316 1109 1344
rect 1137 1316 1173 1344
rect 1201 1316 1237 1344
rect 1265 1334 1270 1344
rect 1298 1430 1912 1490
rect 1298 1402 1303 1430
rect 1331 1402 1367 1430
rect 1395 1402 1431 1430
rect 1459 1402 1495 1430
rect 1523 1402 1559 1430
rect 1587 1402 1623 1430
rect 1651 1402 1687 1430
rect 1715 1402 1751 1430
rect 1779 1402 1815 1430
rect 1843 1402 1879 1430
rect 1907 1402 1912 1430
rect 1298 1344 1912 1402
rect 1298 1334 1303 1344
rect 1265 1317 1303 1334
rect 1265 1316 1270 1317
rect 656 1258 1270 1316
rect 656 1230 661 1258
rect 689 1230 725 1258
rect 753 1230 789 1258
rect 817 1230 853 1258
rect 881 1230 917 1258
rect 945 1230 981 1258
rect 1009 1230 1045 1258
rect 1073 1230 1109 1258
rect 1137 1230 1173 1258
rect 1201 1230 1237 1258
rect 1265 1230 1270 1258
rect 656 1170 1270 1230
rect 1298 1316 1303 1317
rect 1331 1316 1367 1344
rect 1395 1316 1431 1344
rect 1459 1316 1495 1344
rect 1523 1316 1559 1344
rect 1587 1316 1623 1344
rect 1651 1316 1687 1344
rect 1715 1316 1751 1344
rect 1779 1316 1815 1344
rect 1843 1316 1879 1344
rect 1907 1334 1912 1344
rect 1940 1430 2554 1490
rect 1940 1402 1945 1430
rect 1973 1402 2009 1430
rect 2037 1402 2073 1430
rect 2101 1402 2137 1430
rect 2165 1402 2201 1430
rect 2229 1402 2265 1430
rect 2293 1402 2329 1430
rect 2357 1402 2393 1430
rect 2421 1402 2457 1430
rect 2485 1402 2521 1430
rect 2549 1402 2554 1430
rect 1940 1344 2554 1402
rect 1940 1334 1945 1344
rect 1907 1317 1945 1334
rect 1907 1316 1912 1317
rect 1298 1258 1912 1316
rect 1298 1230 1303 1258
rect 1331 1230 1367 1258
rect 1395 1230 1431 1258
rect 1459 1230 1495 1258
rect 1523 1230 1559 1258
rect 1587 1230 1623 1258
rect 1651 1230 1687 1258
rect 1715 1230 1751 1258
rect 1779 1230 1815 1258
rect 1843 1230 1879 1258
rect 1907 1230 1912 1258
rect 1298 1170 1912 1230
rect 1940 1316 1945 1317
rect 1973 1316 2009 1344
rect 2037 1316 2073 1344
rect 2101 1316 2137 1344
rect 2165 1316 2201 1344
rect 2229 1316 2265 1344
rect 2293 1316 2329 1344
rect 2357 1316 2393 1344
rect 2421 1316 2457 1344
rect 2485 1316 2521 1344
rect 2549 1334 2554 1344
rect 2582 1430 3196 1490
rect 2582 1402 2587 1430
rect 2615 1402 2651 1430
rect 2679 1402 2715 1430
rect 2743 1402 2779 1430
rect 2807 1402 2843 1430
rect 2871 1402 2907 1430
rect 2935 1402 2971 1430
rect 2999 1402 3035 1430
rect 3063 1402 3099 1430
rect 3127 1402 3163 1430
rect 3191 1402 3196 1430
rect 2582 1344 3196 1402
rect 2582 1334 2587 1344
rect 2549 1317 2587 1334
rect 2549 1316 2554 1317
rect 1940 1258 2554 1316
rect 1940 1230 1945 1258
rect 1973 1230 2009 1258
rect 2037 1230 2073 1258
rect 2101 1230 2137 1258
rect 2165 1230 2201 1258
rect 2229 1230 2265 1258
rect 2293 1230 2329 1258
rect 2357 1230 2393 1258
rect 2421 1230 2457 1258
rect 2485 1230 2521 1258
rect 2549 1230 2554 1258
rect 1940 1170 2554 1230
rect 2582 1316 2587 1317
rect 2615 1316 2651 1344
rect 2679 1316 2715 1344
rect 2743 1316 2779 1344
rect 2807 1316 2843 1344
rect 2871 1316 2907 1344
rect 2935 1316 2971 1344
rect 2999 1316 3035 1344
rect 3063 1316 3099 1344
rect 3127 1316 3163 1344
rect 3191 1334 3196 1344
rect 3224 1430 3838 1490
rect 3224 1402 3229 1430
rect 3257 1402 3293 1430
rect 3321 1402 3357 1430
rect 3385 1402 3421 1430
rect 3449 1402 3485 1430
rect 3513 1402 3549 1430
rect 3577 1402 3613 1430
rect 3641 1402 3677 1430
rect 3705 1402 3741 1430
rect 3769 1402 3805 1430
rect 3833 1402 3838 1430
rect 3224 1344 3838 1402
rect 3224 1334 3229 1344
rect 3191 1317 3229 1334
rect 3191 1316 3196 1317
rect 2582 1258 3196 1316
rect 2582 1230 2587 1258
rect 2615 1230 2651 1258
rect 2679 1230 2715 1258
rect 2743 1230 2779 1258
rect 2807 1230 2843 1258
rect 2871 1230 2907 1258
rect 2935 1230 2971 1258
rect 2999 1230 3035 1258
rect 3063 1230 3099 1258
rect 3127 1230 3163 1258
rect 3191 1230 3196 1258
rect 2582 1170 3196 1230
rect 3224 1316 3229 1317
rect 3257 1316 3293 1344
rect 3321 1316 3357 1344
rect 3385 1316 3421 1344
rect 3449 1316 3485 1344
rect 3513 1316 3549 1344
rect 3577 1316 3613 1344
rect 3641 1316 3677 1344
rect 3705 1316 3741 1344
rect 3769 1316 3805 1344
rect 3833 1334 3838 1344
rect 3866 1430 4480 1490
rect 3866 1402 3871 1430
rect 3899 1402 3935 1430
rect 3963 1402 3999 1430
rect 4027 1402 4063 1430
rect 4091 1402 4127 1430
rect 4155 1402 4191 1430
rect 4219 1402 4255 1430
rect 4283 1402 4319 1430
rect 4347 1402 4383 1430
rect 4411 1402 4447 1430
rect 4475 1402 4480 1430
rect 3866 1344 4480 1402
rect 3866 1334 3871 1344
rect 3833 1317 3871 1334
rect 3833 1316 3838 1317
rect 3224 1258 3838 1316
rect 3224 1230 3229 1258
rect 3257 1230 3293 1258
rect 3321 1230 3357 1258
rect 3385 1230 3421 1258
rect 3449 1230 3485 1258
rect 3513 1230 3549 1258
rect 3577 1230 3613 1258
rect 3641 1230 3677 1258
rect 3705 1230 3741 1258
rect 3769 1230 3805 1258
rect 3833 1230 3838 1258
rect 3224 1170 3838 1230
rect 3866 1316 3871 1317
rect 3899 1316 3935 1344
rect 3963 1316 3999 1344
rect 4027 1316 4063 1344
rect 4091 1316 4127 1344
rect 4155 1316 4191 1344
rect 4219 1316 4255 1344
rect 4283 1316 4319 1344
rect 4347 1316 4383 1344
rect 4411 1316 4447 1344
rect 4475 1334 4480 1344
rect 4508 1430 5122 1490
rect 4508 1402 4513 1430
rect 4541 1402 4577 1430
rect 4605 1402 4641 1430
rect 4669 1402 4705 1430
rect 4733 1402 4769 1430
rect 4797 1402 4833 1430
rect 4861 1402 4897 1430
rect 4925 1402 4961 1430
rect 4989 1402 5025 1430
rect 5053 1402 5089 1430
rect 5117 1402 5122 1430
rect 4508 1344 5122 1402
rect 4508 1334 4513 1344
rect 4475 1317 4513 1334
rect 4475 1316 4480 1317
rect 3866 1258 4480 1316
rect 3866 1230 3871 1258
rect 3899 1230 3935 1258
rect 3963 1230 3999 1258
rect 4027 1230 4063 1258
rect 4091 1230 4127 1258
rect 4155 1230 4191 1258
rect 4219 1230 4255 1258
rect 4283 1230 4319 1258
rect 4347 1230 4383 1258
rect 4411 1230 4447 1258
rect 4475 1230 4480 1258
rect 3866 1170 4480 1230
rect 4508 1316 4513 1317
rect 4541 1316 4577 1344
rect 4605 1316 4641 1344
rect 4669 1316 4705 1344
rect 4733 1316 4769 1344
rect 4797 1316 4833 1344
rect 4861 1316 4897 1344
rect 4925 1316 4961 1344
rect 4989 1316 5025 1344
rect 5053 1316 5089 1344
rect 5117 1334 5122 1344
rect 5150 1430 5764 1490
rect 5150 1402 5155 1430
rect 5183 1402 5219 1430
rect 5247 1402 5283 1430
rect 5311 1402 5347 1430
rect 5375 1402 5411 1430
rect 5439 1402 5475 1430
rect 5503 1402 5539 1430
rect 5567 1402 5603 1430
rect 5631 1402 5667 1430
rect 5695 1402 5731 1430
rect 5759 1402 5764 1430
rect 5150 1344 5764 1402
rect 5150 1334 5155 1344
rect 5117 1317 5155 1334
rect 5117 1316 5122 1317
rect 4508 1258 5122 1316
rect 4508 1230 4513 1258
rect 4541 1230 4577 1258
rect 4605 1230 4641 1258
rect 4669 1230 4705 1258
rect 4733 1230 4769 1258
rect 4797 1230 4833 1258
rect 4861 1230 4897 1258
rect 4925 1230 4961 1258
rect 4989 1230 5025 1258
rect 5053 1230 5089 1258
rect 5117 1230 5122 1258
rect 4508 1170 5122 1230
rect 5150 1316 5155 1317
rect 5183 1316 5219 1344
rect 5247 1316 5283 1344
rect 5311 1316 5347 1344
rect 5375 1316 5411 1344
rect 5439 1316 5475 1344
rect 5503 1316 5539 1344
rect 5567 1316 5603 1344
rect 5631 1316 5667 1344
rect 5695 1316 5731 1344
rect 5759 1334 5764 1344
rect 5792 1430 6406 1490
rect 5792 1402 5797 1430
rect 5825 1402 5861 1430
rect 5889 1402 5925 1430
rect 5953 1402 5989 1430
rect 6017 1402 6053 1430
rect 6081 1402 6117 1430
rect 6145 1402 6181 1430
rect 6209 1402 6245 1430
rect 6273 1402 6309 1430
rect 6337 1402 6373 1430
rect 6401 1402 6406 1430
rect 5792 1344 6406 1402
rect 5792 1334 5797 1344
rect 5759 1317 5797 1334
rect 5759 1316 5764 1317
rect 5150 1258 5764 1316
rect 5150 1230 5155 1258
rect 5183 1230 5219 1258
rect 5247 1230 5283 1258
rect 5311 1230 5347 1258
rect 5375 1230 5411 1258
rect 5439 1230 5475 1258
rect 5503 1230 5539 1258
rect 5567 1230 5603 1258
rect 5631 1230 5667 1258
rect 5695 1230 5731 1258
rect 5759 1230 5764 1258
rect 5150 1170 5764 1230
rect 5792 1316 5797 1317
rect 5825 1316 5861 1344
rect 5889 1316 5925 1344
rect 5953 1316 5989 1344
rect 6017 1316 6053 1344
rect 6081 1316 6117 1344
rect 6145 1316 6181 1344
rect 6209 1316 6245 1344
rect 6273 1316 6309 1344
rect 6337 1316 6373 1344
rect 6401 1334 6406 1344
rect 6434 1430 7048 1490
rect 6434 1402 6439 1430
rect 6467 1402 6503 1430
rect 6531 1402 6567 1430
rect 6595 1402 6631 1430
rect 6659 1402 6695 1430
rect 6723 1402 6759 1430
rect 6787 1402 6823 1430
rect 6851 1402 6887 1430
rect 6915 1402 6951 1430
rect 6979 1402 7015 1430
rect 7043 1402 7048 1430
rect 6434 1344 7048 1402
rect 6434 1334 6439 1344
rect 6401 1317 6439 1334
rect 6401 1316 6406 1317
rect 5792 1258 6406 1316
rect 5792 1230 5797 1258
rect 5825 1230 5861 1258
rect 5889 1230 5925 1258
rect 5953 1230 5989 1258
rect 6017 1230 6053 1258
rect 6081 1230 6117 1258
rect 6145 1230 6181 1258
rect 6209 1230 6245 1258
rect 6273 1230 6309 1258
rect 6337 1230 6373 1258
rect 6401 1230 6406 1258
rect 5792 1170 6406 1230
rect 6434 1316 6439 1317
rect 6467 1316 6503 1344
rect 6531 1316 6567 1344
rect 6595 1316 6631 1344
rect 6659 1316 6695 1344
rect 6723 1316 6759 1344
rect 6787 1316 6823 1344
rect 6851 1316 6887 1344
rect 6915 1316 6951 1344
rect 6979 1316 7015 1344
rect 7043 1334 7048 1344
rect 7076 1430 7690 1490
rect 7076 1402 7081 1430
rect 7109 1402 7145 1430
rect 7173 1402 7209 1430
rect 7237 1402 7273 1430
rect 7301 1402 7337 1430
rect 7365 1402 7401 1430
rect 7429 1402 7465 1430
rect 7493 1402 7529 1430
rect 7557 1402 7593 1430
rect 7621 1402 7657 1430
rect 7685 1402 7690 1430
rect 7076 1344 7690 1402
rect 7076 1334 7081 1344
rect 7043 1317 7081 1334
rect 7043 1316 7048 1317
rect 6434 1258 7048 1316
rect 6434 1230 6439 1258
rect 6467 1230 6503 1258
rect 6531 1230 6567 1258
rect 6595 1230 6631 1258
rect 6659 1230 6695 1258
rect 6723 1230 6759 1258
rect 6787 1230 6823 1258
rect 6851 1230 6887 1258
rect 6915 1230 6951 1258
rect 6979 1230 7015 1258
rect 7043 1230 7048 1258
rect 6434 1170 7048 1230
rect 7076 1316 7081 1317
rect 7109 1316 7145 1344
rect 7173 1316 7209 1344
rect 7237 1316 7273 1344
rect 7301 1316 7337 1344
rect 7365 1316 7401 1344
rect 7429 1316 7465 1344
rect 7493 1316 7529 1344
rect 7557 1316 7593 1344
rect 7621 1316 7657 1344
rect 7685 1334 7690 1344
rect 7718 1430 8332 1490
rect 7718 1402 7723 1430
rect 7751 1402 7787 1430
rect 7815 1402 7851 1430
rect 7879 1402 7915 1430
rect 7943 1402 7979 1430
rect 8007 1402 8043 1430
rect 8071 1402 8107 1430
rect 8135 1402 8171 1430
rect 8199 1402 8235 1430
rect 8263 1402 8299 1430
rect 8327 1402 8332 1430
rect 7718 1344 8332 1402
rect 7718 1334 7723 1344
rect 7685 1317 7723 1334
rect 7685 1316 7690 1317
rect 7076 1258 7690 1316
rect 7076 1230 7081 1258
rect 7109 1230 7145 1258
rect 7173 1230 7209 1258
rect 7237 1230 7273 1258
rect 7301 1230 7337 1258
rect 7365 1230 7401 1258
rect 7429 1230 7465 1258
rect 7493 1230 7529 1258
rect 7557 1230 7593 1258
rect 7621 1230 7657 1258
rect 7685 1230 7690 1258
rect 7076 1170 7690 1230
rect 7718 1316 7723 1317
rect 7751 1316 7787 1344
rect 7815 1316 7851 1344
rect 7879 1316 7915 1344
rect 7943 1316 7979 1344
rect 8007 1316 8043 1344
rect 8071 1316 8107 1344
rect 8135 1316 8171 1344
rect 8199 1316 8235 1344
rect 8263 1316 8299 1344
rect 8327 1334 8332 1344
rect 8360 1430 8974 1490
rect 8360 1402 8365 1430
rect 8393 1402 8429 1430
rect 8457 1402 8493 1430
rect 8521 1402 8557 1430
rect 8585 1402 8621 1430
rect 8649 1402 8685 1430
rect 8713 1402 8749 1430
rect 8777 1402 8813 1430
rect 8841 1402 8877 1430
rect 8905 1402 8941 1430
rect 8969 1402 8974 1430
rect 8360 1344 8974 1402
rect 8360 1334 8365 1344
rect 8327 1317 8365 1334
rect 8327 1316 8332 1317
rect 7718 1258 8332 1316
rect 7718 1230 7723 1258
rect 7751 1230 7787 1258
rect 7815 1230 7851 1258
rect 7879 1230 7915 1258
rect 7943 1230 7979 1258
rect 8007 1230 8043 1258
rect 8071 1230 8107 1258
rect 8135 1230 8171 1258
rect 8199 1230 8235 1258
rect 8263 1230 8299 1258
rect 8327 1230 8332 1258
rect 7718 1170 8332 1230
rect 8360 1316 8365 1317
rect 8393 1316 8429 1344
rect 8457 1316 8493 1344
rect 8521 1316 8557 1344
rect 8585 1316 8621 1344
rect 8649 1316 8685 1344
rect 8713 1316 8749 1344
rect 8777 1316 8813 1344
rect 8841 1316 8877 1344
rect 8905 1316 8941 1344
rect 8969 1334 8974 1344
rect 9002 1430 9616 1490
rect 9002 1402 9007 1430
rect 9035 1402 9071 1430
rect 9099 1402 9135 1430
rect 9163 1402 9199 1430
rect 9227 1402 9263 1430
rect 9291 1402 9327 1430
rect 9355 1402 9391 1430
rect 9419 1402 9455 1430
rect 9483 1402 9519 1430
rect 9547 1402 9583 1430
rect 9611 1402 9616 1430
rect 9002 1344 9616 1402
rect 9002 1334 9007 1344
rect 8969 1317 9007 1334
rect 8969 1316 8974 1317
rect 8360 1258 8974 1316
rect 8360 1230 8365 1258
rect 8393 1230 8429 1258
rect 8457 1230 8493 1258
rect 8521 1230 8557 1258
rect 8585 1230 8621 1258
rect 8649 1230 8685 1258
rect 8713 1230 8749 1258
rect 8777 1230 8813 1258
rect 8841 1230 8877 1258
rect 8905 1230 8941 1258
rect 8969 1230 8974 1258
rect 8360 1170 8974 1230
rect 9002 1316 9007 1317
rect 9035 1316 9071 1344
rect 9099 1316 9135 1344
rect 9163 1316 9199 1344
rect 9227 1316 9263 1344
rect 9291 1316 9327 1344
rect 9355 1316 9391 1344
rect 9419 1316 9455 1344
rect 9483 1316 9519 1344
rect 9547 1316 9583 1344
rect 9611 1334 9616 1344
rect 9644 1430 10258 1490
rect 9644 1402 9649 1430
rect 9677 1402 9713 1430
rect 9741 1402 9777 1430
rect 9805 1402 9841 1430
rect 9869 1402 9905 1430
rect 9933 1402 9969 1430
rect 9997 1402 10033 1430
rect 10061 1402 10097 1430
rect 10125 1402 10161 1430
rect 10189 1402 10225 1430
rect 10253 1402 10258 1430
rect 9644 1344 10258 1402
rect 9644 1334 9649 1344
rect 9611 1317 9649 1334
rect 9611 1316 9616 1317
rect 9002 1258 9616 1316
rect 9002 1230 9007 1258
rect 9035 1230 9071 1258
rect 9099 1230 9135 1258
rect 9163 1230 9199 1258
rect 9227 1230 9263 1258
rect 9291 1230 9327 1258
rect 9355 1230 9391 1258
rect 9419 1230 9455 1258
rect 9483 1230 9519 1258
rect 9547 1230 9583 1258
rect 9611 1230 9616 1258
rect 9002 1170 9616 1230
rect 9644 1316 9649 1317
rect 9677 1316 9713 1344
rect 9741 1316 9777 1344
rect 9805 1316 9841 1344
rect 9869 1316 9905 1344
rect 9933 1316 9969 1344
rect 9997 1316 10033 1344
rect 10061 1316 10097 1344
rect 10125 1316 10161 1344
rect 10189 1316 10225 1344
rect 10253 1334 10258 1344
rect 10286 1430 10900 1490
rect 10286 1402 10291 1430
rect 10319 1402 10355 1430
rect 10383 1402 10419 1430
rect 10447 1402 10483 1430
rect 10511 1402 10547 1430
rect 10575 1402 10611 1430
rect 10639 1402 10675 1430
rect 10703 1402 10739 1430
rect 10767 1402 10803 1430
rect 10831 1402 10867 1430
rect 10895 1402 10900 1430
rect 10286 1344 10900 1402
rect 10286 1334 10291 1344
rect 10253 1317 10291 1334
rect 10253 1316 10258 1317
rect 9644 1258 10258 1316
rect 9644 1230 9649 1258
rect 9677 1230 9713 1258
rect 9741 1230 9777 1258
rect 9805 1230 9841 1258
rect 9869 1230 9905 1258
rect 9933 1230 9969 1258
rect 9997 1230 10033 1258
rect 10061 1230 10097 1258
rect 10125 1230 10161 1258
rect 10189 1230 10225 1258
rect 10253 1230 10258 1258
rect 9644 1170 10258 1230
rect 10286 1316 10291 1317
rect 10319 1316 10355 1344
rect 10383 1316 10419 1344
rect 10447 1316 10483 1344
rect 10511 1316 10547 1344
rect 10575 1316 10611 1344
rect 10639 1316 10675 1344
rect 10703 1316 10739 1344
rect 10767 1316 10803 1344
rect 10831 1316 10867 1344
rect 10895 1334 10900 1344
rect 10928 1430 11542 1490
rect 10928 1402 10933 1430
rect 10961 1402 10997 1430
rect 11025 1402 11061 1430
rect 11089 1402 11125 1430
rect 11153 1402 11189 1430
rect 11217 1402 11253 1430
rect 11281 1402 11317 1430
rect 11345 1402 11381 1430
rect 11409 1402 11445 1430
rect 11473 1402 11509 1430
rect 11537 1402 11542 1430
rect 10928 1344 11542 1402
rect 10928 1334 10933 1344
rect 10895 1317 10933 1334
rect 10895 1316 10900 1317
rect 10286 1258 10900 1316
rect 10286 1230 10291 1258
rect 10319 1230 10355 1258
rect 10383 1230 10419 1258
rect 10447 1230 10483 1258
rect 10511 1230 10547 1258
rect 10575 1230 10611 1258
rect 10639 1230 10675 1258
rect 10703 1230 10739 1258
rect 10767 1230 10803 1258
rect 10831 1230 10867 1258
rect 10895 1230 10900 1258
rect 10286 1170 10900 1230
rect 10928 1316 10933 1317
rect 10961 1316 10997 1344
rect 11025 1316 11061 1344
rect 11089 1316 11125 1344
rect 11153 1316 11189 1344
rect 11217 1316 11253 1344
rect 11281 1316 11317 1344
rect 11345 1316 11381 1344
rect 11409 1316 11445 1344
rect 11473 1316 11509 1344
rect 11537 1334 11542 1344
rect 11570 1430 12184 1490
rect 11570 1402 11575 1430
rect 11603 1402 11639 1430
rect 11667 1402 11703 1430
rect 11731 1402 11767 1430
rect 11795 1402 11831 1430
rect 11859 1402 11895 1430
rect 11923 1402 11959 1430
rect 11987 1402 12023 1430
rect 12051 1402 12087 1430
rect 12115 1402 12151 1430
rect 12179 1402 12184 1430
rect 11570 1344 12184 1402
rect 11570 1334 11575 1344
rect 11537 1317 11575 1334
rect 11537 1316 11542 1317
rect 10928 1258 11542 1316
rect 10928 1230 10933 1258
rect 10961 1230 10997 1258
rect 11025 1230 11061 1258
rect 11089 1230 11125 1258
rect 11153 1230 11189 1258
rect 11217 1230 11253 1258
rect 11281 1230 11317 1258
rect 11345 1230 11381 1258
rect 11409 1230 11445 1258
rect 11473 1230 11509 1258
rect 11537 1230 11542 1258
rect 10928 1170 11542 1230
rect 11570 1316 11575 1317
rect 11603 1316 11639 1344
rect 11667 1316 11703 1344
rect 11731 1316 11767 1344
rect 11795 1316 11831 1344
rect 11859 1316 11895 1344
rect 11923 1316 11959 1344
rect 11987 1316 12023 1344
rect 12051 1316 12087 1344
rect 12115 1316 12151 1344
rect 12179 1334 12184 1344
rect 12212 1430 12826 1490
rect 12212 1402 12217 1430
rect 12245 1402 12281 1430
rect 12309 1402 12345 1430
rect 12373 1402 12409 1430
rect 12437 1402 12473 1430
rect 12501 1402 12537 1430
rect 12565 1402 12601 1430
rect 12629 1402 12665 1430
rect 12693 1402 12729 1430
rect 12757 1402 12793 1430
rect 12821 1402 12826 1430
rect 12212 1344 12826 1402
rect 12212 1334 12217 1344
rect 12179 1317 12217 1334
rect 12179 1316 12184 1317
rect 11570 1258 12184 1316
rect 11570 1230 11575 1258
rect 11603 1230 11639 1258
rect 11667 1230 11703 1258
rect 11731 1230 11767 1258
rect 11795 1230 11831 1258
rect 11859 1230 11895 1258
rect 11923 1230 11959 1258
rect 11987 1230 12023 1258
rect 12051 1230 12087 1258
rect 12115 1230 12151 1258
rect 12179 1230 12184 1258
rect 11570 1170 12184 1230
rect 12212 1316 12217 1317
rect 12245 1316 12281 1344
rect 12309 1316 12345 1344
rect 12373 1316 12409 1344
rect 12437 1316 12473 1344
rect 12501 1316 12537 1344
rect 12565 1316 12601 1344
rect 12629 1316 12665 1344
rect 12693 1316 12729 1344
rect 12757 1316 12793 1344
rect 12821 1316 12826 1344
rect 12212 1258 12826 1316
rect 12212 1230 12217 1258
rect 12245 1230 12281 1258
rect 12309 1230 12345 1258
rect 12373 1230 12409 1258
rect 12437 1230 12473 1258
rect 12501 1230 12537 1258
rect 12565 1230 12601 1258
rect 12629 1230 12665 1258
rect 12693 1230 12729 1258
rect 12757 1230 12793 1258
rect 12821 1230 12826 1258
rect 12212 1170 12826 1230
rect 315 1110 329 1170
rect 2877 1110 2891 1170
rect 3521 1110 3535 1170
rect 6089 1110 6103 1170
rect 6668 1110 6682 1170
rect 9299 1110 9313 1170
rect 9941 1110 9955 1170
rect 12507 1110 12521 1170
rect 14 1050 628 1110
rect 14 1022 19 1050
rect 47 1022 83 1050
rect 111 1022 147 1050
rect 175 1022 211 1050
rect 239 1022 275 1050
rect 303 1022 339 1050
rect 367 1022 403 1050
rect 431 1022 467 1050
rect 495 1022 531 1050
rect 559 1022 595 1050
rect 623 1022 628 1050
rect 14 964 628 1022
rect 14 936 19 964
rect 47 936 83 964
rect 111 936 147 964
rect 175 936 211 964
rect 239 936 275 964
rect 303 936 339 964
rect 367 936 403 964
rect 431 936 467 964
rect 495 936 531 964
rect 559 936 595 964
rect 623 936 628 964
rect 14 878 628 936
rect 14 850 19 878
rect 47 850 83 878
rect 111 850 147 878
rect 175 850 211 878
rect 239 850 275 878
rect 303 850 339 878
rect 367 850 403 878
rect 431 850 467 878
rect 495 850 531 878
rect 559 850 595 878
rect 623 850 628 878
rect 14 790 628 850
rect 656 1050 1270 1110
rect 656 1022 661 1050
rect 689 1022 725 1050
rect 753 1022 789 1050
rect 817 1022 853 1050
rect 881 1022 917 1050
rect 945 1022 981 1050
rect 1009 1022 1045 1050
rect 1073 1022 1109 1050
rect 1137 1022 1173 1050
rect 1201 1022 1237 1050
rect 1265 1022 1270 1050
rect 656 964 1270 1022
rect 656 936 661 964
rect 689 936 725 964
rect 753 936 789 964
rect 817 936 853 964
rect 881 936 917 964
rect 945 936 981 964
rect 1009 936 1045 964
rect 1073 936 1109 964
rect 1137 936 1173 964
rect 1201 936 1237 964
rect 1265 936 1270 964
rect 656 878 1270 936
rect 656 850 661 878
rect 689 850 725 878
rect 753 850 789 878
rect 817 850 853 878
rect 881 850 917 878
rect 945 850 981 878
rect 1009 850 1045 878
rect 1073 850 1109 878
rect 1137 850 1173 878
rect 1201 850 1237 878
rect 1265 850 1270 878
rect 656 804 1270 850
rect 1298 1050 1912 1110
rect 1298 1022 1303 1050
rect 1331 1022 1367 1050
rect 1395 1022 1431 1050
rect 1459 1022 1495 1050
rect 1523 1022 1559 1050
rect 1587 1022 1623 1050
rect 1651 1022 1687 1050
rect 1715 1022 1751 1050
rect 1779 1022 1815 1050
rect 1843 1022 1879 1050
rect 1907 1022 1912 1050
rect 1298 964 1912 1022
rect 1298 936 1303 964
rect 1331 936 1367 964
rect 1395 936 1431 964
rect 1459 936 1495 964
rect 1523 936 1559 964
rect 1587 936 1623 964
rect 1651 936 1687 964
rect 1715 936 1751 964
rect 1779 936 1815 964
rect 1843 936 1879 964
rect 1907 936 1912 964
rect 1298 878 1912 936
rect 1298 850 1303 878
rect 1331 850 1367 878
rect 1395 850 1431 878
rect 1459 850 1495 878
rect 1523 850 1559 878
rect 1587 850 1623 878
rect 1651 850 1687 878
rect 1715 850 1751 878
rect 1779 850 1815 878
rect 1843 850 1879 878
rect 1907 850 1912 878
rect 1298 806 1912 850
rect 1940 1050 2554 1110
rect 1940 1022 1945 1050
rect 1973 1022 2009 1050
rect 2037 1022 2073 1050
rect 2101 1022 2137 1050
rect 2165 1022 2201 1050
rect 2229 1022 2265 1050
rect 2293 1022 2329 1050
rect 2357 1022 2393 1050
rect 2421 1022 2457 1050
rect 2485 1022 2521 1050
rect 2549 1022 2554 1050
rect 1940 964 2554 1022
rect 1940 936 1945 964
rect 1973 936 2009 964
rect 2037 936 2073 964
rect 2101 936 2137 964
rect 2165 936 2201 964
rect 2229 936 2265 964
rect 2293 936 2329 964
rect 2357 936 2393 964
rect 2421 936 2457 964
rect 2485 936 2521 964
rect 2549 936 2554 964
rect 1940 878 2554 936
rect 1940 850 1945 878
rect 1973 850 2009 878
rect 2037 850 2073 878
rect 2101 850 2137 878
rect 2165 850 2201 878
rect 2229 850 2265 878
rect 2293 850 2329 878
rect 2357 850 2393 878
rect 2421 850 2457 878
rect 2485 850 2521 878
rect 2549 850 2554 878
rect 1940 806 2554 850
rect 1298 804 2554 806
rect 656 791 2554 804
rect 656 790 1912 791
rect 1940 790 2554 791
rect 2582 1050 3196 1110
rect 2582 1022 2587 1050
rect 2615 1022 2651 1050
rect 2679 1022 2715 1050
rect 2743 1022 2779 1050
rect 2807 1022 2843 1050
rect 2871 1022 2907 1050
rect 2935 1022 2971 1050
rect 2999 1022 3035 1050
rect 3063 1022 3099 1050
rect 3127 1022 3163 1050
rect 3191 1022 3196 1050
rect 2582 964 3196 1022
rect 2582 936 2587 964
rect 2615 936 2651 964
rect 2679 936 2715 964
rect 2743 936 2779 964
rect 2807 936 2843 964
rect 2871 936 2907 964
rect 2935 936 2971 964
rect 2999 936 3035 964
rect 3063 936 3099 964
rect 3127 936 3163 964
rect 3191 936 3196 964
rect 2582 878 3196 936
rect 2582 850 2587 878
rect 2615 850 2651 878
rect 2679 850 2715 878
rect 2743 850 2779 878
rect 2807 850 2843 878
rect 2871 850 2907 878
rect 2935 850 2971 878
rect 2999 850 3035 878
rect 3063 850 3099 878
rect 3127 850 3163 878
rect 3191 850 3196 878
rect 2582 790 3196 850
rect 3224 1050 3838 1110
rect 3224 1022 3229 1050
rect 3257 1022 3293 1050
rect 3321 1022 3357 1050
rect 3385 1022 3421 1050
rect 3449 1022 3485 1050
rect 3513 1022 3549 1050
rect 3577 1022 3613 1050
rect 3641 1022 3677 1050
rect 3705 1022 3741 1050
rect 3769 1022 3805 1050
rect 3833 1022 3838 1050
rect 3224 964 3838 1022
rect 3224 936 3229 964
rect 3257 936 3293 964
rect 3321 936 3357 964
rect 3385 936 3421 964
rect 3449 936 3485 964
rect 3513 936 3549 964
rect 3577 936 3613 964
rect 3641 936 3677 964
rect 3705 936 3741 964
rect 3769 936 3805 964
rect 3833 936 3838 964
rect 3224 878 3838 936
rect 3224 850 3229 878
rect 3257 850 3293 878
rect 3321 850 3357 878
rect 3385 850 3421 878
rect 3449 850 3485 878
rect 3513 850 3549 878
rect 3577 850 3613 878
rect 3641 850 3677 878
rect 3705 850 3741 878
rect 3769 850 3805 878
rect 3833 850 3838 878
rect 3224 790 3838 850
rect 3866 1050 4480 1110
rect 3866 1022 3871 1050
rect 3899 1022 3935 1050
rect 3963 1022 3999 1050
rect 4027 1022 4063 1050
rect 4091 1022 4127 1050
rect 4155 1022 4191 1050
rect 4219 1022 4255 1050
rect 4283 1022 4319 1050
rect 4347 1022 4383 1050
rect 4411 1022 4447 1050
rect 4475 1022 4480 1050
rect 3866 964 4480 1022
rect 3866 936 3871 964
rect 3899 936 3935 964
rect 3963 936 3999 964
rect 4027 936 4063 964
rect 4091 936 4127 964
rect 4155 936 4191 964
rect 4219 936 4255 964
rect 4283 936 4319 964
rect 4347 936 4383 964
rect 4411 936 4447 964
rect 4475 936 4480 964
rect 3866 878 4480 936
rect 3866 850 3871 878
rect 3899 850 3935 878
rect 3963 850 3999 878
rect 4027 850 4063 878
rect 4091 850 4127 878
rect 4155 850 4191 878
rect 4219 850 4255 878
rect 4283 850 4319 878
rect 4347 850 4383 878
rect 4411 850 4447 878
rect 4475 850 4480 878
rect 3866 807 4480 850
rect 4508 1050 5122 1110
rect 4508 1022 4513 1050
rect 4541 1022 4577 1050
rect 4605 1022 4641 1050
rect 4669 1022 4705 1050
rect 4733 1022 4769 1050
rect 4797 1022 4833 1050
rect 4861 1022 4897 1050
rect 4925 1022 4961 1050
rect 4989 1022 5025 1050
rect 5053 1022 5089 1050
rect 5117 1022 5122 1050
rect 4508 964 5122 1022
rect 4508 936 4513 964
rect 4541 936 4577 964
rect 4605 936 4641 964
rect 4669 936 4705 964
rect 4733 936 4769 964
rect 4797 936 4833 964
rect 4861 936 4897 964
rect 4925 936 4961 964
rect 4989 936 5025 964
rect 5053 936 5089 964
rect 5117 936 5122 964
rect 4508 878 5122 936
rect 4508 850 4513 878
rect 4541 850 4577 878
rect 4605 850 4641 878
rect 4669 850 4705 878
rect 4733 850 4769 878
rect 4797 850 4833 878
rect 4861 850 4897 878
rect 4925 850 4961 878
rect 4989 850 5025 878
rect 5053 850 5089 878
rect 5117 850 5122 878
rect 4508 807 5122 850
rect 3866 804 5122 807
rect 5150 1050 5764 1110
rect 5150 1022 5155 1050
rect 5183 1022 5219 1050
rect 5247 1022 5283 1050
rect 5311 1022 5347 1050
rect 5375 1022 5411 1050
rect 5439 1022 5475 1050
rect 5503 1022 5539 1050
rect 5567 1022 5603 1050
rect 5631 1022 5667 1050
rect 5695 1022 5731 1050
rect 5759 1022 5764 1050
rect 5150 964 5764 1022
rect 5150 936 5155 964
rect 5183 936 5219 964
rect 5247 936 5283 964
rect 5311 936 5347 964
rect 5375 936 5411 964
rect 5439 936 5475 964
rect 5503 936 5539 964
rect 5567 936 5603 964
rect 5631 936 5667 964
rect 5695 936 5731 964
rect 5759 936 5764 964
rect 5150 878 5764 936
rect 5150 850 5155 878
rect 5183 850 5219 878
rect 5247 850 5283 878
rect 5311 850 5347 878
rect 5375 850 5411 878
rect 5439 850 5475 878
rect 5503 850 5539 878
rect 5567 850 5603 878
rect 5631 850 5667 878
rect 5695 850 5731 878
rect 5759 850 5764 878
rect 5150 804 5764 850
rect 3866 792 5764 804
rect 3866 790 4480 792
rect 4508 790 5764 792
rect 5792 1050 6406 1110
rect 5792 1022 5797 1050
rect 5825 1022 5861 1050
rect 5889 1022 5925 1050
rect 5953 1022 5989 1050
rect 6017 1022 6053 1050
rect 6081 1022 6117 1050
rect 6145 1022 6181 1050
rect 6209 1022 6245 1050
rect 6273 1022 6309 1050
rect 6337 1022 6373 1050
rect 6401 1022 6406 1050
rect 5792 964 6406 1022
rect 5792 936 5797 964
rect 5825 936 5861 964
rect 5889 936 5925 964
rect 5953 936 5989 964
rect 6017 936 6053 964
rect 6081 936 6117 964
rect 6145 936 6181 964
rect 6209 936 6245 964
rect 6273 936 6309 964
rect 6337 936 6373 964
rect 6401 936 6406 964
rect 5792 878 6406 936
rect 5792 850 5797 878
rect 5825 850 5861 878
rect 5889 850 5925 878
rect 5953 850 5989 878
rect 6017 850 6053 878
rect 6081 850 6117 878
rect 6145 850 6181 878
rect 6209 850 6245 878
rect 6273 850 6309 878
rect 6337 850 6373 878
rect 6401 850 6406 878
rect 5792 790 6406 850
rect 6434 1050 7048 1110
rect 6434 1022 6439 1050
rect 6467 1022 6503 1050
rect 6531 1022 6567 1050
rect 6595 1022 6631 1050
rect 6659 1022 6695 1050
rect 6723 1022 6759 1050
rect 6787 1022 6823 1050
rect 6851 1022 6887 1050
rect 6915 1022 6951 1050
rect 6979 1022 7015 1050
rect 7043 1022 7048 1050
rect 6434 964 7048 1022
rect 6434 936 6439 964
rect 6467 936 6503 964
rect 6531 936 6567 964
rect 6595 936 6631 964
rect 6659 936 6695 964
rect 6723 936 6759 964
rect 6787 936 6823 964
rect 6851 936 6887 964
rect 6915 936 6951 964
rect 6979 936 7015 964
rect 7043 936 7048 964
rect 6434 878 7048 936
rect 6434 850 6439 878
rect 6467 850 6503 878
rect 6531 850 6567 878
rect 6595 850 6631 878
rect 6659 850 6695 878
rect 6723 850 6759 878
rect 6787 850 6823 878
rect 6851 850 6887 878
rect 6915 850 6951 878
rect 6979 850 7015 878
rect 7043 850 7048 878
rect 6434 790 7048 850
rect 7076 1050 7690 1110
rect 7076 1022 7081 1050
rect 7109 1022 7145 1050
rect 7173 1022 7209 1050
rect 7237 1022 7273 1050
rect 7301 1022 7337 1050
rect 7365 1022 7401 1050
rect 7429 1022 7465 1050
rect 7493 1022 7529 1050
rect 7557 1022 7593 1050
rect 7621 1022 7657 1050
rect 7685 1022 7690 1050
rect 7076 964 7690 1022
rect 7076 936 7081 964
rect 7109 936 7145 964
rect 7173 936 7209 964
rect 7237 936 7273 964
rect 7301 936 7337 964
rect 7365 936 7401 964
rect 7429 936 7465 964
rect 7493 936 7529 964
rect 7557 936 7593 964
rect 7621 936 7657 964
rect 7685 936 7690 964
rect 7076 878 7690 936
rect 7076 850 7081 878
rect 7109 850 7145 878
rect 7173 850 7209 878
rect 7237 850 7273 878
rect 7301 850 7337 878
rect 7365 850 7401 878
rect 7429 850 7465 878
rect 7493 850 7529 878
rect 7557 850 7593 878
rect 7621 850 7657 878
rect 7685 850 7690 878
rect 7076 805 7690 850
rect 7718 1050 8332 1110
rect 7718 1022 7723 1050
rect 7751 1022 7787 1050
rect 7815 1022 7851 1050
rect 7879 1022 7915 1050
rect 7943 1022 7979 1050
rect 8007 1022 8043 1050
rect 8071 1022 8107 1050
rect 8135 1022 8171 1050
rect 8199 1022 8235 1050
rect 8263 1022 8299 1050
rect 8327 1022 8332 1050
rect 7718 964 8332 1022
rect 7718 936 7723 964
rect 7751 936 7787 964
rect 7815 936 7851 964
rect 7879 936 7915 964
rect 7943 936 7979 964
rect 8007 936 8043 964
rect 8071 936 8107 964
rect 8135 936 8171 964
rect 8199 936 8235 964
rect 8263 936 8299 964
rect 8327 936 8332 964
rect 7718 878 8332 936
rect 7718 850 7723 878
rect 7751 850 7787 878
rect 7815 850 7851 878
rect 7879 850 7915 878
rect 7943 850 7979 878
rect 8007 850 8043 878
rect 8071 850 8107 878
rect 8135 850 8171 878
rect 8199 850 8235 878
rect 8263 850 8299 878
rect 8327 850 8332 878
rect 7718 805 8332 850
rect 7076 804 8332 805
rect 8360 1050 8974 1110
rect 8360 1022 8365 1050
rect 8393 1022 8429 1050
rect 8457 1022 8493 1050
rect 8521 1022 8557 1050
rect 8585 1022 8621 1050
rect 8649 1022 8685 1050
rect 8713 1022 8749 1050
rect 8777 1022 8813 1050
rect 8841 1022 8877 1050
rect 8905 1022 8941 1050
rect 8969 1022 8974 1050
rect 8360 964 8974 1022
rect 8360 936 8365 964
rect 8393 936 8429 964
rect 8457 936 8493 964
rect 8521 936 8557 964
rect 8585 936 8621 964
rect 8649 936 8685 964
rect 8713 936 8749 964
rect 8777 936 8813 964
rect 8841 936 8877 964
rect 8905 936 8941 964
rect 8969 936 8974 964
rect 8360 878 8974 936
rect 8360 850 8365 878
rect 8393 850 8429 878
rect 8457 850 8493 878
rect 8521 850 8557 878
rect 8585 850 8621 878
rect 8649 850 8685 878
rect 8713 850 8749 878
rect 8777 850 8813 878
rect 8841 850 8877 878
rect 8905 850 8941 878
rect 8969 850 8974 878
rect 8360 804 8974 850
rect 7076 790 8974 804
rect 9002 1050 9616 1110
rect 9002 1022 9007 1050
rect 9035 1022 9071 1050
rect 9099 1022 9135 1050
rect 9163 1022 9199 1050
rect 9227 1022 9263 1050
rect 9291 1022 9327 1050
rect 9355 1022 9391 1050
rect 9419 1022 9455 1050
rect 9483 1022 9519 1050
rect 9547 1022 9583 1050
rect 9611 1022 9616 1050
rect 9002 964 9616 1022
rect 9002 936 9007 964
rect 9035 936 9071 964
rect 9099 936 9135 964
rect 9163 936 9199 964
rect 9227 936 9263 964
rect 9291 936 9327 964
rect 9355 936 9391 964
rect 9419 936 9455 964
rect 9483 936 9519 964
rect 9547 936 9583 964
rect 9611 936 9616 964
rect 9002 878 9616 936
rect 9002 850 9007 878
rect 9035 850 9071 878
rect 9099 850 9135 878
rect 9163 850 9199 878
rect 9227 850 9263 878
rect 9291 850 9327 878
rect 9355 850 9391 878
rect 9419 850 9455 878
rect 9483 850 9519 878
rect 9547 850 9583 878
rect 9611 850 9616 878
rect 9002 790 9616 850
rect 9644 1050 10258 1110
rect 9644 1022 9649 1050
rect 9677 1022 9713 1050
rect 9741 1022 9777 1050
rect 9805 1022 9841 1050
rect 9869 1022 9905 1050
rect 9933 1022 9969 1050
rect 9997 1022 10033 1050
rect 10061 1022 10097 1050
rect 10125 1022 10161 1050
rect 10189 1022 10225 1050
rect 10253 1022 10258 1050
rect 9644 964 10258 1022
rect 9644 936 9649 964
rect 9677 936 9713 964
rect 9741 936 9777 964
rect 9805 936 9841 964
rect 9869 936 9905 964
rect 9933 936 9969 964
rect 9997 936 10033 964
rect 10061 936 10097 964
rect 10125 936 10161 964
rect 10189 936 10225 964
rect 10253 936 10258 964
rect 9644 878 10258 936
rect 9644 850 9649 878
rect 9677 850 9713 878
rect 9741 850 9777 878
rect 9805 850 9841 878
rect 9869 850 9905 878
rect 9933 850 9969 878
rect 9997 850 10033 878
rect 10061 850 10097 878
rect 10125 850 10161 878
rect 10189 850 10225 878
rect 10253 850 10258 878
rect 9644 790 10258 850
rect 10286 1050 10900 1110
rect 10286 1022 10291 1050
rect 10319 1022 10355 1050
rect 10383 1022 10419 1050
rect 10447 1022 10483 1050
rect 10511 1022 10547 1050
rect 10575 1022 10611 1050
rect 10639 1022 10675 1050
rect 10703 1022 10739 1050
rect 10767 1022 10803 1050
rect 10831 1022 10867 1050
rect 10895 1022 10900 1050
rect 10286 964 10900 1022
rect 10286 936 10291 964
rect 10319 936 10355 964
rect 10383 936 10419 964
rect 10447 936 10483 964
rect 10511 936 10547 964
rect 10575 936 10611 964
rect 10639 936 10675 964
rect 10703 936 10739 964
rect 10767 936 10803 964
rect 10831 936 10867 964
rect 10895 936 10900 964
rect 10286 878 10900 936
rect 10286 850 10291 878
rect 10319 850 10355 878
rect 10383 850 10419 878
rect 10447 850 10483 878
rect 10511 850 10547 878
rect 10575 850 10611 878
rect 10639 850 10675 878
rect 10703 850 10739 878
rect 10767 850 10803 878
rect 10831 850 10867 878
rect 10895 850 10900 878
rect 10286 806 10900 850
rect 10928 1050 11542 1110
rect 10928 1022 10933 1050
rect 10961 1022 10997 1050
rect 11025 1022 11061 1050
rect 11089 1022 11125 1050
rect 11153 1022 11189 1050
rect 11217 1022 11253 1050
rect 11281 1022 11317 1050
rect 11345 1022 11381 1050
rect 11409 1022 11445 1050
rect 11473 1022 11509 1050
rect 11537 1022 11542 1050
rect 10928 964 11542 1022
rect 10928 936 10933 964
rect 10961 936 10997 964
rect 11025 936 11061 964
rect 11089 936 11125 964
rect 11153 936 11189 964
rect 11217 936 11253 964
rect 11281 936 11317 964
rect 11345 936 11381 964
rect 11409 936 11445 964
rect 11473 936 11509 964
rect 11537 936 11542 964
rect 10928 878 11542 936
rect 10928 850 10933 878
rect 10961 850 10997 878
rect 11025 850 11061 878
rect 11089 850 11125 878
rect 11153 850 11189 878
rect 11217 850 11253 878
rect 11281 850 11317 878
rect 11345 850 11381 878
rect 11409 850 11445 878
rect 11473 850 11509 878
rect 11537 850 11542 878
rect 10928 806 11542 850
rect 10286 804 11542 806
rect 11570 1050 12184 1110
rect 11570 1022 11575 1050
rect 11603 1022 11639 1050
rect 11667 1022 11703 1050
rect 11731 1022 11767 1050
rect 11795 1022 11831 1050
rect 11859 1022 11895 1050
rect 11923 1022 11959 1050
rect 11987 1022 12023 1050
rect 12051 1022 12087 1050
rect 12115 1022 12151 1050
rect 12179 1022 12184 1050
rect 11570 964 12184 1022
rect 11570 936 11575 964
rect 11603 936 11639 964
rect 11667 936 11703 964
rect 11731 936 11767 964
rect 11795 936 11831 964
rect 11859 936 11895 964
rect 11923 936 11959 964
rect 11987 936 12023 964
rect 12051 936 12087 964
rect 12115 936 12151 964
rect 12179 936 12184 964
rect 11570 878 12184 936
rect 11570 850 11575 878
rect 11603 850 11639 878
rect 11667 850 11703 878
rect 11731 850 11767 878
rect 11795 850 11831 878
rect 11859 850 11895 878
rect 11923 850 11959 878
rect 11987 850 12023 878
rect 12051 850 12087 878
rect 12115 850 12151 878
rect 12179 850 12184 878
rect 11570 804 12184 850
rect 10286 791 12184 804
rect 10286 790 10900 791
rect 10928 790 12184 791
rect 12212 1050 12826 1110
rect 12212 1022 12217 1050
rect 12245 1022 12281 1050
rect 12309 1022 12345 1050
rect 12373 1022 12409 1050
rect 12437 1022 12473 1050
rect 12501 1022 12537 1050
rect 12565 1022 12601 1050
rect 12629 1022 12665 1050
rect 12693 1022 12729 1050
rect 12757 1022 12793 1050
rect 12821 1022 12826 1050
rect 12212 964 12826 1022
rect 12212 936 12217 964
rect 12245 936 12281 964
rect 12309 936 12345 964
rect 12373 936 12409 964
rect 12437 936 12473 964
rect 12501 936 12537 964
rect 12565 936 12601 964
rect 12629 936 12665 964
rect 12693 936 12729 964
rect 12757 936 12793 964
rect 12821 936 12826 964
rect 12212 878 12826 936
rect 12212 850 12217 878
rect 12245 850 12281 878
rect 12309 850 12345 878
rect 12373 850 12409 878
rect 12437 850 12473 878
rect 12501 850 12537 878
rect 12565 850 12601 878
rect 12629 850 12665 878
rect 12693 850 12729 878
rect 12757 850 12793 878
rect 12821 850 12826 878
rect 12212 790 12826 850
rect 315 730 329 790
rect 1260 789 1306 790
rect 1597 730 1612 790
rect 2877 730 2891 790
rect 3521 730 3535 790
rect 4867 730 4882 790
rect 6089 730 6103 790
rect 6668 730 6682 790
rect 8079 730 8094 790
rect 8323 789 8368 790
rect 9299 730 9313 790
rect 9941 730 9955 790
rect 11225 730 11240 790
rect 11536 789 11581 790
rect 12507 730 12521 790
rect 14 670 628 730
rect 14 642 19 670
rect 47 642 83 670
rect 111 642 147 670
rect 175 642 211 670
rect 239 642 275 670
rect 303 642 339 670
rect 367 642 403 670
rect 431 642 467 670
rect 495 642 531 670
rect 559 642 595 670
rect 623 642 628 670
rect 14 584 628 642
rect 14 556 19 584
rect 47 556 83 584
rect 111 556 147 584
rect 175 556 211 584
rect 239 556 275 584
rect 303 556 339 584
rect 367 556 403 584
rect 431 556 467 584
rect 495 556 531 584
rect 559 556 595 584
rect 623 556 628 584
rect 14 498 628 556
rect 14 470 19 498
rect 47 470 83 498
rect 111 470 147 498
rect 175 470 211 498
rect 239 470 275 498
rect 303 470 339 498
rect 367 470 403 498
rect 431 470 467 498
rect 495 470 531 498
rect 559 470 595 498
rect 623 470 628 498
rect 14 410 628 470
rect 656 670 1270 730
rect 656 642 661 670
rect 689 642 725 670
rect 753 642 789 670
rect 817 642 853 670
rect 881 642 917 670
rect 945 642 981 670
rect 1009 642 1045 670
rect 1073 642 1109 670
rect 1137 642 1173 670
rect 1201 642 1237 670
rect 1265 642 1270 670
rect 656 584 1270 642
rect 656 556 661 584
rect 689 556 725 584
rect 753 556 789 584
rect 817 556 853 584
rect 881 556 917 584
rect 945 556 981 584
rect 1009 556 1045 584
rect 1073 556 1109 584
rect 1137 556 1173 584
rect 1201 556 1237 584
rect 1265 556 1270 584
rect 656 498 1270 556
rect 656 470 661 498
rect 689 470 725 498
rect 753 470 789 498
rect 817 470 853 498
rect 881 470 917 498
rect 945 470 981 498
rect 1009 470 1045 498
rect 1073 470 1109 498
rect 1137 470 1173 498
rect 1201 470 1237 498
rect 1265 470 1270 498
rect 656 425 1270 470
rect 1298 670 1912 730
rect 1298 642 1303 670
rect 1331 642 1367 670
rect 1395 642 1431 670
rect 1459 642 1495 670
rect 1523 642 1559 670
rect 1587 642 1623 670
rect 1651 642 1687 670
rect 1715 642 1751 670
rect 1779 642 1815 670
rect 1843 642 1879 670
rect 1907 642 1912 670
rect 1298 584 1912 642
rect 1298 556 1303 584
rect 1331 556 1367 584
rect 1395 556 1431 584
rect 1459 556 1495 584
rect 1523 556 1559 584
rect 1587 556 1623 584
rect 1651 556 1687 584
rect 1715 556 1751 584
rect 1779 556 1815 584
rect 1843 556 1879 584
rect 1907 556 1912 584
rect 1298 498 1912 556
rect 1298 470 1303 498
rect 1331 470 1367 498
rect 1395 470 1431 498
rect 1459 470 1495 498
rect 1523 470 1559 498
rect 1587 470 1623 498
rect 1651 470 1687 498
rect 1715 470 1751 498
rect 1779 470 1815 498
rect 1843 470 1879 498
rect 1907 470 1912 498
rect 1298 425 1912 470
rect 1940 670 2554 730
rect 1940 642 1945 670
rect 1973 642 2009 670
rect 2037 642 2073 670
rect 2101 642 2137 670
rect 2165 642 2201 670
rect 2229 642 2265 670
rect 2293 642 2329 670
rect 2357 642 2393 670
rect 2421 642 2457 670
rect 2485 642 2521 670
rect 2549 642 2554 670
rect 1940 584 2554 642
rect 1940 556 1945 584
rect 1973 556 2009 584
rect 2037 556 2073 584
rect 2101 556 2137 584
rect 2165 556 2201 584
rect 2229 556 2265 584
rect 2293 556 2329 584
rect 2357 556 2393 584
rect 2421 556 2457 584
rect 2485 556 2521 584
rect 2549 556 2554 584
rect 1940 498 2554 556
rect 1940 470 1945 498
rect 1973 470 2009 498
rect 2037 470 2073 498
rect 2101 470 2137 498
rect 2165 470 2201 498
rect 2229 470 2265 498
rect 2293 470 2329 498
rect 2357 470 2393 498
rect 2421 470 2457 498
rect 2485 470 2521 498
rect 2549 470 2554 498
rect 1940 425 2554 470
rect 656 410 2554 425
rect 2582 670 3196 730
rect 2582 642 2587 670
rect 2615 642 2651 670
rect 2679 642 2715 670
rect 2743 642 2779 670
rect 2807 642 2843 670
rect 2871 642 2907 670
rect 2935 642 2971 670
rect 2999 642 3035 670
rect 3063 642 3099 670
rect 3127 642 3163 670
rect 3191 642 3196 670
rect 2582 584 3196 642
rect 2582 556 2587 584
rect 2615 556 2651 584
rect 2679 556 2715 584
rect 2743 556 2779 584
rect 2807 556 2843 584
rect 2871 556 2907 584
rect 2935 556 2971 584
rect 2999 556 3035 584
rect 3063 556 3099 584
rect 3127 556 3163 584
rect 3191 556 3196 584
rect 2582 498 3196 556
rect 2582 470 2587 498
rect 2615 470 2651 498
rect 2679 470 2715 498
rect 2743 470 2779 498
rect 2807 470 2843 498
rect 2871 470 2907 498
rect 2935 470 2971 498
rect 2999 470 3035 498
rect 3063 470 3099 498
rect 3127 470 3163 498
rect 3191 470 3196 498
rect 2582 410 3196 470
rect 3224 670 3838 730
rect 3224 642 3229 670
rect 3257 642 3293 670
rect 3321 642 3357 670
rect 3385 642 3421 670
rect 3449 642 3485 670
rect 3513 642 3549 670
rect 3577 642 3613 670
rect 3641 642 3677 670
rect 3705 642 3741 670
rect 3769 642 3805 670
rect 3833 642 3838 670
rect 3224 584 3838 642
rect 3224 556 3229 584
rect 3257 556 3293 584
rect 3321 556 3357 584
rect 3385 556 3421 584
rect 3449 556 3485 584
rect 3513 556 3549 584
rect 3577 556 3613 584
rect 3641 556 3677 584
rect 3705 556 3741 584
rect 3769 556 3805 584
rect 3833 556 3838 584
rect 3224 498 3838 556
rect 3224 470 3229 498
rect 3257 470 3293 498
rect 3321 470 3357 498
rect 3385 470 3421 498
rect 3449 470 3485 498
rect 3513 470 3549 498
rect 3577 470 3613 498
rect 3641 470 3677 498
rect 3705 470 3741 498
rect 3769 470 3805 498
rect 3833 470 3838 498
rect 3224 410 3838 470
rect 3866 670 4480 730
rect 3866 642 3871 670
rect 3899 642 3935 670
rect 3963 642 3999 670
rect 4027 642 4063 670
rect 4091 642 4127 670
rect 4155 642 4191 670
rect 4219 642 4255 670
rect 4283 642 4319 670
rect 4347 642 4383 670
rect 4411 642 4447 670
rect 4475 642 4480 670
rect 3866 584 4480 642
rect 3866 556 3871 584
rect 3899 556 3935 584
rect 3963 556 3999 584
rect 4027 556 4063 584
rect 4091 556 4127 584
rect 4155 556 4191 584
rect 4219 556 4255 584
rect 4283 556 4319 584
rect 4347 556 4383 584
rect 4411 556 4447 584
rect 4475 556 4480 584
rect 3866 498 4480 556
rect 3866 470 3871 498
rect 3899 470 3935 498
rect 3963 470 3999 498
rect 4027 470 4063 498
rect 4091 470 4127 498
rect 4155 470 4191 498
rect 4219 470 4255 498
rect 4283 470 4319 498
rect 4347 470 4383 498
rect 4411 470 4447 498
rect 4475 470 4480 498
rect 3866 423 4480 470
rect 4508 670 5122 730
rect 4508 642 4513 670
rect 4541 642 4577 670
rect 4605 642 4641 670
rect 4669 642 4705 670
rect 4733 642 4769 670
rect 4797 642 4833 670
rect 4861 642 4897 670
rect 4925 642 4961 670
rect 4989 642 5025 670
rect 5053 642 5089 670
rect 5117 642 5122 670
rect 4508 584 5122 642
rect 4508 556 4513 584
rect 4541 556 4577 584
rect 4605 556 4641 584
rect 4669 556 4705 584
rect 4733 556 4769 584
rect 4797 556 4833 584
rect 4861 556 4897 584
rect 4925 556 4961 584
rect 4989 556 5025 584
rect 5053 556 5089 584
rect 5117 556 5122 584
rect 4508 498 5122 556
rect 4508 470 4513 498
rect 4541 470 4577 498
rect 4605 470 4641 498
rect 4669 470 4705 498
rect 4733 470 4769 498
rect 4797 470 4833 498
rect 4861 470 4897 498
rect 4925 470 4961 498
rect 4989 470 5025 498
rect 5053 470 5089 498
rect 5117 470 5122 498
rect 4508 426 5122 470
rect 5150 670 5764 730
rect 5150 642 5155 670
rect 5183 642 5219 670
rect 5247 642 5283 670
rect 5311 642 5347 670
rect 5375 642 5411 670
rect 5439 642 5475 670
rect 5503 642 5539 670
rect 5567 642 5603 670
rect 5631 642 5667 670
rect 5695 642 5731 670
rect 5759 642 5764 670
rect 5150 584 5764 642
rect 5150 556 5155 584
rect 5183 556 5219 584
rect 5247 556 5283 584
rect 5311 556 5347 584
rect 5375 556 5411 584
rect 5439 556 5475 584
rect 5503 556 5539 584
rect 5567 556 5603 584
rect 5631 556 5667 584
rect 5695 556 5731 584
rect 5759 556 5764 584
rect 5150 498 5764 556
rect 5150 470 5155 498
rect 5183 470 5219 498
rect 5247 470 5283 498
rect 5311 470 5347 498
rect 5375 470 5411 498
rect 5439 470 5475 498
rect 5503 470 5539 498
rect 5567 470 5603 498
rect 5631 470 5667 498
rect 5695 470 5731 498
rect 5759 470 5764 498
rect 5150 426 5764 470
rect 4508 423 5764 426
rect 3866 411 5764 423
rect 3866 410 5122 411
rect 5150 410 5764 411
rect 5792 670 6406 730
rect 5792 642 5797 670
rect 5825 642 5861 670
rect 5889 642 5925 670
rect 5953 642 5989 670
rect 6017 642 6053 670
rect 6081 642 6117 670
rect 6145 642 6181 670
rect 6209 642 6245 670
rect 6273 642 6309 670
rect 6337 642 6373 670
rect 6401 642 6406 670
rect 5792 584 6406 642
rect 5792 556 5797 584
rect 5825 556 5861 584
rect 5889 556 5925 584
rect 5953 556 5989 584
rect 6017 556 6053 584
rect 6081 556 6117 584
rect 6145 556 6181 584
rect 6209 556 6245 584
rect 6273 556 6309 584
rect 6337 556 6373 584
rect 6401 556 6406 584
rect 5792 498 6406 556
rect 5792 470 5797 498
rect 5825 470 5861 498
rect 5889 470 5925 498
rect 5953 470 5989 498
rect 6017 470 6053 498
rect 6081 470 6117 498
rect 6145 470 6181 498
rect 6209 470 6245 498
rect 6273 470 6309 498
rect 6337 470 6373 498
rect 6401 470 6406 498
rect 5792 410 6406 470
rect 6434 670 7048 730
rect 6434 642 6439 670
rect 6467 642 6503 670
rect 6531 642 6567 670
rect 6595 642 6631 670
rect 6659 642 6695 670
rect 6723 642 6759 670
rect 6787 642 6823 670
rect 6851 642 6887 670
rect 6915 642 6951 670
rect 6979 642 7015 670
rect 7043 642 7048 670
rect 6434 584 7048 642
rect 6434 556 6439 584
rect 6467 556 6503 584
rect 6531 556 6567 584
rect 6595 556 6631 584
rect 6659 556 6695 584
rect 6723 556 6759 584
rect 6787 556 6823 584
rect 6851 556 6887 584
rect 6915 556 6951 584
rect 6979 556 7015 584
rect 7043 556 7048 584
rect 6434 498 7048 556
rect 6434 470 6439 498
rect 6467 470 6503 498
rect 6531 470 6567 498
rect 6595 470 6631 498
rect 6659 470 6695 498
rect 6723 470 6759 498
rect 6787 470 6823 498
rect 6851 470 6887 498
rect 6915 470 6951 498
rect 6979 470 7015 498
rect 7043 470 7048 498
rect 6434 410 7048 470
rect 7076 670 7690 730
rect 7076 642 7081 670
rect 7109 642 7145 670
rect 7173 642 7209 670
rect 7237 642 7273 670
rect 7301 642 7337 670
rect 7365 642 7401 670
rect 7429 642 7465 670
rect 7493 642 7529 670
rect 7557 642 7593 670
rect 7621 642 7657 670
rect 7685 642 7690 670
rect 7076 584 7690 642
rect 7076 556 7081 584
rect 7109 556 7145 584
rect 7173 556 7209 584
rect 7237 556 7273 584
rect 7301 556 7337 584
rect 7365 556 7401 584
rect 7429 556 7465 584
rect 7493 556 7529 584
rect 7557 556 7593 584
rect 7621 556 7657 584
rect 7685 556 7690 584
rect 7076 498 7690 556
rect 7076 470 7081 498
rect 7109 470 7145 498
rect 7173 470 7209 498
rect 7237 470 7273 498
rect 7301 470 7337 498
rect 7365 470 7401 498
rect 7429 470 7465 498
rect 7493 470 7529 498
rect 7557 470 7593 498
rect 7621 470 7657 498
rect 7685 470 7690 498
rect 7076 426 7690 470
rect 7718 670 8332 730
rect 7718 642 7723 670
rect 7751 642 7787 670
rect 7815 642 7851 670
rect 7879 642 7915 670
rect 7943 642 7979 670
rect 8007 642 8043 670
rect 8071 642 8107 670
rect 8135 642 8171 670
rect 8199 642 8235 670
rect 8263 642 8299 670
rect 8327 642 8332 670
rect 7718 584 8332 642
rect 7718 556 7723 584
rect 7751 556 7787 584
rect 7815 556 7851 584
rect 7879 556 7915 584
rect 7943 556 7979 584
rect 8007 556 8043 584
rect 8071 556 8107 584
rect 8135 556 8171 584
rect 8199 556 8235 584
rect 8263 556 8299 584
rect 8327 556 8332 584
rect 7718 498 8332 556
rect 7718 470 7723 498
rect 7751 470 7787 498
rect 7815 470 7851 498
rect 7879 470 7915 498
rect 7943 470 7979 498
rect 8007 470 8043 498
rect 8071 470 8107 498
rect 8135 470 8171 498
rect 8199 470 8235 498
rect 8263 470 8299 498
rect 8327 470 8332 498
rect 7718 426 8332 470
rect 8360 670 8974 730
rect 8360 642 8365 670
rect 8393 642 8429 670
rect 8457 642 8493 670
rect 8521 642 8557 670
rect 8585 642 8621 670
rect 8649 642 8685 670
rect 8713 642 8749 670
rect 8777 642 8813 670
rect 8841 642 8877 670
rect 8905 642 8941 670
rect 8969 642 8974 670
rect 8360 584 8974 642
rect 8360 556 8365 584
rect 8393 556 8429 584
rect 8457 556 8493 584
rect 8521 556 8557 584
rect 8585 556 8621 584
rect 8649 556 8685 584
rect 8713 556 8749 584
rect 8777 556 8813 584
rect 8841 556 8877 584
rect 8905 556 8941 584
rect 8969 556 8974 584
rect 8360 498 8974 556
rect 8360 470 8365 498
rect 8393 470 8429 498
rect 8457 470 8493 498
rect 8521 470 8557 498
rect 8585 470 8621 498
rect 8649 470 8685 498
rect 8713 470 8749 498
rect 8777 470 8813 498
rect 8841 470 8877 498
rect 8905 470 8941 498
rect 8969 470 8974 498
rect 8360 426 8974 470
rect 7076 411 8974 426
rect 7076 410 7690 411
rect 7718 410 8332 411
rect 8360 410 8974 411
rect 9002 670 9616 730
rect 9002 642 9007 670
rect 9035 642 9071 670
rect 9099 642 9135 670
rect 9163 642 9199 670
rect 9227 642 9263 670
rect 9291 642 9327 670
rect 9355 642 9391 670
rect 9419 642 9455 670
rect 9483 642 9519 670
rect 9547 642 9583 670
rect 9611 642 9616 670
rect 9002 584 9616 642
rect 9002 556 9007 584
rect 9035 556 9071 584
rect 9099 556 9135 584
rect 9163 556 9199 584
rect 9227 556 9263 584
rect 9291 556 9327 584
rect 9355 556 9391 584
rect 9419 556 9455 584
rect 9483 556 9519 584
rect 9547 556 9583 584
rect 9611 556 9616 584
rect 9002 498 9616 556
rect 9002 470 9007 498
rect 9035 470 9071 498
rect 9099 470 9135 498
rect 9163 470 9199 498
rect 9227 470 9263 498
rect 9291 470 9327 498
rect 9355 470 9391 498
rect 9419 470 9455 498
rect 9483 470 9519 498
rect 9547 470 9583 498
rect 9611 470 9616 498
rect 9002 410 9616 470
rect 9644 670 10258 730
rect 9644 642 9649 670
rect 9677 642 9713 670
rect 9741 642 9777 670
rect 9805 642 9841 670
rect 9869 642 9905 670
rect 9933 642 9969 670
rect 9997 642 10033 670
rect 10061 642 10097 670
rect 10125 642 10161 670
rect 10189 642 10225 670
rect 10253 642 10258 670
rect 9644 584 10258 642
rect 9644 556 9649 584
rect 9677 556 9713 584
rect 9741 556 9777 584
rect 9805 556 9841 584
rect 9869 556 9905 584
rect 9933 556 9969 584
rect 9997 556 10033 584
rect 10061 556 10097 584
rect 10125 556 10161 584
rect 10189 556 10225 584
rect 10253 556 10258 584
rect 9644 498 10258 556
rect 9644 470 9649 498
rect 9677 470 9713 498
rect 9741 470 9777 498
rect 9805 470 9841 498
rect 9869 470 9905 498
rect 9933 470 9969 498
rect 9997 470 10033 498
rect 10061 470 10097 498
rect 10125 470 10161 498
rect 10189 470 10225 498
rect 10253 470 10258 498
rect 9644 410 10258 470
rect 10286 670 10900 730
rect 10286 642 10291 670
rect 10319 642 10355 670
rect 10383 642 10419 670
rect 10447 642 10483 670
rect 10511 642 10547 670
rect 10575 642 10611 670
rect 10639 642 10675 670
rect 10703 642 10739 670
rect 10767 642 10803 670
rect 10831 642 10867 670
rect 10895 642 10900 670
rect 10286 584 10900 642
rect 10286 556 10291 584
rect 10319 556 10355 584
rect 10383 556 10419 584
rect 10447 556 10483 584
rect 10511 556 10547 584
rect 10575 556 10611 584
rect 10639 556 10675 584
rect 10703 556 10739 584
rect 10767 556 10803 584
rect 10831 556 10867 584
rect 10895 556 10900 584
rect 10286 498 10900 556
rect 10286 470 10291 498
rect 10319 470 10355 498
rect 10383 470 10419 498
rect 10447 470 10483 498
rect 10511 470 10547 498
rect 10575 470 10611 498
rect 10639 470 10675 498
rect 10703 470 10739 498
rect 10767 470 10803 498
rect 10831 470 10867 498
rect 10895 470 10900 498
rect 10286 425 10900 470
rect 10928 670 11542 730
rect 10928 642 10933 670
rect 10961 642 10997 670
rect 11025 642 11061 670
rect 11089 642 11125 670
rect 11153 642 11189 670
rect 11217 642 11253 670
rect 11281 642 11317 670
rect 11345 642 11381 670
rect 11409 642 11445 670
rect 11473 642 11509 670
rect 11537 642 11542 670
rect 10928 584 11542 642
rect 10928 556 10933 584
rect 10961 556 10997 584
rect 11025 556 11061 584
rect 11089 556 11125 584
rect 11153 556 11189 584
rect 11217 556 11253 584
rect 11281 556 11317 584
rect 11345 556 11381 584
rect 11409 556 11445 584
rect 11473 556 11509 584
rect 11537 556 11542 584
rect 10928 498 11542 556
rect 10928 470 10933 498
rect 10961 470 10997 498
rect 11025 470 11061 498
rect 11089 470 11125 498
rect 11153 470 11189 498
rect 11217 470 11253 498
rect 11281 470 11317 498
rect 11345 470 11381 498
rect 11409 470 11445 498
rect 11473 470 11509 498
rect 11537 470 11542 498
rect 10928 425 11542 470
rect 11570 670 12184 730
rect 11570 642 11575 670
rect 11603 642 11639 670
rect 11667 642 11703 670
rect 11731 642 11767 670
rect 11795 642 11831 670
rect 11859 642 11895 670
rect 11923 642 11959 670
rect 11987 642 12023 670
rect 12051 642 12087 670
rect 12115 642 12151 670
rect 12179 642 12184 670
rect 11570 584 12184 642
rect 11570 556 11575 584
rect 11603 556 11639 584
rect 11667 556 11703 584
rect 11731 556 11767 584
rect 11795 556 11831 584
rect 11859 556 11895 584
rect 11923 556 11959 584
rect 11987 556 12023 584
rect 12051 556 12087 584
rect 12115 556 12151 584
rect 12179 556 12184 584
rect 11570 498 12184 556
rect 11570 470 11575 498
rect 11603 470 11639 498
rect 11667 470 11703 498
rect 11731 470 11767 498
rect 11795 470 11831 498
rect 11859 470 11895 498
rect 11923 470 11959 498
rect 11987 470 12023 498
rect 12051 470 12087 498
rect 12115 470 12151 498
rect 12179 470 12184 498
rect 11570 425 12184 470
rect 10286 410 12184 425
rect 12212 670 12826 730
rect 12212 642 12217 670
rect 12245 642 12281 670
rect 12309 642 12345 670
rect 12373 642 12409 670
rect 12437 642 12473 670
rect 12501 642 12537 670
rect 12565 642 12601 670
rect 12629 642 12665 670
rect 12693 642 12729 670
rect 12757 642 12793 670
rect 12821 642 12826 670
rect 12212 584 12826 642
rect 12212 556 12217 584
rect 12245 556 12281 584
rect 12309 556 12345 584
rect 12373 556 12409 584
rect 12437 556 12473 584
rect 12501 556 12537 584
rect 12565 556 12601 584
rect 12629 556 12665 584
rect 12693 556 12729 584
rect 12757 556 12793 584
rect 12821 556 12826 584
rect 12212 498 12826 556
rect 12212 470 12217 498
rect 12245 470 12281 498
rect 12309 470 12345 498
rect 12373 470 12409 498
rect 12437 470 12473 498
rect 12501 470 12537 498
rect 12565 470 12601 498
rect 12629 470 12665 498
rect 12693 470 12729 498
rect 12757 470 12793 498
rect 12821 470 12826 498
rect 12212 410 12826 470
rect 315 350 329 410
rect 2877 350 2891 410
rect 3521 350 3535 410
rect 4469 408 4514 410
rect 5080 350 5095 410
rect 6089 350 6103 410
rect 6668 350 6682 410
rect 8296 350 8311 410
rect 9299 350 9313 410
rect 9941 350 9955 410
rect 11507 350 11522 410
rect 12507 350 12521 410
rect 14 290 628 350
rect 14 262 19 290
rect 47 262 83 290
rect 111 262 147 290
rect 175 262 211 290
rect 239 262 275 290
rect 303 262 339 290
rect 367 262 403 290
rect 431 262 467 290
rect 495 262 531 290
rect 559 262 595 290
rect 623 262 628 290
rect 14 204 628 262
rect 14 176 19 204
rect 47 176 83 204
rect 111 176 147 204
rect 175 176 211 204
rect 239 176 275 204
rect 303 176 339 204
rect 367 176 403 204
rect 431 176 467 204
rect 495 176 531 204
rect 559 176 595 204
rect 623 176 628 204
rect 14 173 628 176
rect 656 290 1270 350
rect 656 262 661 290
rect 689 262 725 290
rect 753 262 789 290
rect 817 262 853 290
rect 881 262 917 290
rect 945 262 981 290
rect 1009 262 1045 290
rect 1073 262 1109 290
rect 1137 262 1173 290
rect 1201 262 1237 290
rect 1265 262 1270 290
rect 656 204 1270 262
rect 656 176 661 204
rect 689 176 725 204
rect 753 176 789 204
rect 817 176 853 204
rect 881 176 917 204
rect 945 176 981 204
rect 1009 176 1045 204
rect 1073 176 1109 204
rect 1137 176 1173 204
rect 1201 176 1237 204
rect 1265 176 1270 204
rect 656 173 1270 176
rect 1298 290 1912 350
rect 1298 262 1303 290
rect 1331 262 1367 290
rect 1395 262 1431 290
rect 1459 262 1495 290
rect 1523 262 1559 290
rect 1587 262 1623 290
rect 1651 262 1687 290
rect 1715 262 1751 290
rect 1779 262 1815 290
rect 1843 262 1879 290
rect 1907 262 1912 290
rect 1298 204 1912 262
rect 1298 176 1303 204
rect 1331 176 1367 204
rect 1395 176 1431 204
rect 1459 176 1495 204
rect 1523 176 1559 204
rect 1587 176 1623 204
rect 1651 176 1687 204
rect 1715 176 1751 204
rect 1779 176 1815 204
rect 1843 176 1879 204
rect 1907 176 1912 204
rect 1298 173 1912 176
rect 1940 290 2554 350
rect 1940 262 1945 290
rect 1973 262 2009 290
rect 2037 262 2073 290
rect 2101 262 2137 290
rect 2165 262 2201 290
rect 2229 262 2265 290
rect 2293 262 2329 290
rect 2357 262 2393 290
rect 2421 262 2457 290
rect 2485 262 2521 290
rect 2549 262 2554 290
rect 1940 204 2554 262
rect 1940 176 1945 204
rect 1973 176 2009 204
rect 2037 176 2073 204
rect 2101 176 2137 204
rect 2165 176 2201 204
rect 2229 176 2265 204
rect 2293 176 2329 204
rect 2357 176 2393 204
rect 2421 176 2457 204
rect 2485 176 2521 204
rect 2549 176 2554 204
rect 1940 173 2554 176
rect 2582 290 3196 350
rect 2582 262 2587 290
rect 2615 262 2651 290
rect 2679 262 2715 290
rect 2743 262 2779 290
rect 2807 262 2843 290
rect 2871 262 2907 290
rect 2935 262 2971 290
rect 2999 262 3035 290
rect 3063 262 3099 290
rect 3127 262 3163 290
rect 3191 262 3196 290
rect 2582 204 3196 262
rect 2582 176 2587 204
rect 2615 176 2651 204
rect 2679 176 2715 204
rect 2743 176 2779 204
rect 2807 176 2843 204
rect 2871 176 2907 204
rect 2935 176 2971 204
rect 2999 176 3035 204
rect 3063 176 3099 204
rect 3127 176 3163 204
rect 3191 176 3196 204
rect 2582 173 3196 176
rect 3224 290 3838 350
rect 3224 262 3229 290
rect 3257 262 3293 290
rect 3321 262 3357 290
rect 3385 262 3421 290
rect 3449 262 3485 290
rect 3513 262 3549 290
rect 3577 262 3613 290
rect 3641 262 3677 290
rect 3705 262 3741 290
rect 3769 262 3805 290
rect 3833 262 3838 290
rect 3224 204 3838 262
rect 3224 176 3229 204
rect 3257 176 3293 204
rect 3321 176 3357 204
rect 3385 176 3421 204
rect 3449 176 3485 204
rect 3513 176 3549 204
rect 3577 176 3613 204
rect 3641 176 3677 204
rect 3705 176 3741 204
rect 3769 176 3805 204
rect 3833 176 3838 204
rect 3224 173 3838 176
rect 3866 290 4480 350
rect 3866 262 3871 290
rect 3899 262 3935 290
rect 3963 262 3999 290
rect 4027 262 4063 290
rect 4091 262 4127 290
rect 4155 262 4191 290
rect 4219 262 4255 290
rect 4283 262 4319 290
rect 4347 262 4383 290
rect 4411 262 4447 290
rect 4475 262 4480 290
rect 3866 204 4480 262
rect 3866 176 3871 204
rect 3899 176 3935 204
rect 3963 176 3999 204
rect 4027 176 4063 204
rect 4091 176 4127 204
rect 4155 176 4191 204
rect 4219 176 4255 204
rect 4283 176 4319 204
rect 4347 176 4383 204
rect 4411 176 4447 204
rect 4475 176 4480 204
rect 3866 173 4480 176
rect 14 156 4480 173
rect 14 118 628 156
rect 14 90 19 118
rect 47 90 83 118
rect 111 90 147 118
rect 175 90 211 118
rect 239 90 275 118
rect 303 90 339 118
rect 367 90 403 118
rect 431 90 467 118
rect 495 90 531 118
rect 559 90 595 118
rect 623 90 628 118
rect 14 30 628 90
rect 656 118 1270 156
rect 656 90 661 118
rect 689 90 725 118
rect 753 90 789 118
rect 817 90 853 118
rect 881 90 917 118
rect 945 90 981 118
rect 1009 90 1045 118
rect 1073 90 1109 118
rect 1137 90 1173 118
rect 1201 90 1237 118
rect 1265 90 1270 118
rect 656 30 1270 90
rect 1298 118 1912 156
rect 1298 90 1303 118
rect 1331 90 1367 118
rect 1395 90 1431 118
rect 1459 90 1495 118
rect 1523 90 1559 118
rect 1587 90 1623 118
rect 1651 90 1687 118
rect 1715 90 1751 118
rect 1779 90 1815 118
rect 1843 90 1879 118
rect 1907 90 1912 118
rect 1298 30 1912 90
rect 1940 118 2554 156
rect 1940 90 1945 118
rect 1973 90 2009 118
rect 2037 90 2073 118
rect 2101 90 2137 118
rect 2165 90 2201 118
rect 2229 90 2265 118
rect 2293 90 2329 118
rect 2357 90 2393 118
rect 2421 90 2457 118
rect 2485 90 2521 118
rect 2549 90 2554 118
rect 1940 30 2554 90
rect 2582 118 3196 156
rect 2582 90 2587 118
rect 2615 90 2651 118
rect 2679 90 2715 118
rect 2743 90 2779 118
rect 2807 90 2843 118
rect 2871 90 2907 118
rect 2935 90 2971 118
rect 2999 90 3035 118
rect 3063 90 3099 118
rect 3127 90 3163 118
rect 3191 90 3196 118
rect 2582 30 3196 90
rect 3224 118 3838 156
rect 3224 90 3229 118
rect 3257 90 3293 118
rect 3321 90 3357 118
rect 3385 90 3421 118
rect 3449 90 3485 118
rect 3513 90 3549 118
rect 3577 90 3613 118
rect 3641 90 3677 118
rect 3705 90 3741 118
rect 3769 90 3805 118
rect 3833 90 3838 118
rect 3224 30 3838 90
rect 3866 118 4480 156
rect 3866 90 3871 118
rect 3899 90 3935 118
rect 3963 90 3999 118
rect 4027 90 4063 118
rect 4091 90 4127 118
rect 4155 90 4191 118
rect 4219 90 4255 118
rect 4283 90 4319 118
rect 4347 90 4383 118
rect 4411 90 4447 118
rect 4475 90 4480 118
rect 3866 30 4480 90
rect 4508 290 5122 350
rect 4508 262 4513 290
rect 4541 262 4577 290
rect 4605 262 4641 290
rect 4669 262 4705 290
rect 4733 262 4769 290
rect 4797 262 4833 290
rect 4861 262 4897 290
rect 4925 262 4961 290
rect 4989 262 5025 290
rect 5053 262 5089 290
rect 5117 262 5122 290
rect 4508 204 5122 262
rect 4508 176 4513 204
rect 4541 176 4577 204
rect 4605 176 4641 204
rect 4669 176 4705 204
rect 4733 176 4769 204
rect 4797 176 4833 204
rect 4861 176 4897 204
rect 4925 176 4961 204
rect 4989 176 5025 204
rect 5053 176 5089 204
rect 5117 176 5122 204
rect 4508 118 5122 176
rect 4508 90 4513 118
rect 4541 90 4577 118
rect 4605 90 4641 118
rect 4669 90 4705 118
rect 4733 90 4769 118
rect 4797 90 4833 118
rect 4861 90 4897 118
rect 4925 90 4961 118
rect 4989 90 5025 118
rect 5053 90 5089 118
rect 5117 90 5122 118
rect 4508 30 5122 90
rect 5150 290 5764 350
rect 5150 262 5155 290
rect 5183 262 5219 290
rect 5247 262 5283 290
rect 5311 262 5347 290
rect 5375 262 5411 290
rect 5439 262 5475 290
rect 5503 262 5539 290
rect 5567 262 5603 290
rect 5631 262 5667 290
rect 5695 262 5731 290
rect 5759 262 5764 290
rect 5150 204 5764 262
rect 5150 176 5155 204
rect 5183 176 5219 204
rect 5247 176 5283 204
rect 5311 176 5347 204
rect 5375 176 5411 204
rect 5439 176 5475 204
rect 5503 176 5539 204
rect 5567 176 5603 204
rect 5631 176 5667 204
rect 5695 176 5731 204
rect 5759 180 5764 204
rect 5792 290 6406 350
rect 5792 262 5797 290
rect 5825 262 5861 290
rect 5889 262 5925 290
rect 5953 262 5989 290
rect 6017 262 6053 290
rect 6081 262 6117 290
rect 6145 262 6181 290
rect 6209 262 6245 290
rect 6273 262 6309 290
rect 6337 262 6373 290
rect 6401 262 6406 290
rect 5792 204 6406 262
rect 5792 180 5797 204
rect 5759 176 5797 180
rect 5825 176 5861 204
rect 5889 176 5925 204
rect 5953 176 5989 204
rect 6017 176 6053 204
rect 6081 176 6117 204
rect 6145 176 6181 204
rect 6209 176 6245 204
rect 6273 176 6309 204
rect 6337 176 6373 204
rect 6401 180 6406 204
rect 6434 290 7048 350
rect 6434 262 6439 290
rect 6467 262 6503 290
rect 6531 262 6567 290
rect 6595 262 6631 290
rect 6659 262 6695 290
rect 6723 262 6759 290
rect 6787 262 6823 290
rect 6851 262 6887 290
rect 6915 262 6951 290
rect 6979 262 7015 290
rect 7043 262 7048 290
rect 6434 204 7048 262
rect 6434 180 6439 204
rect 6401 176 6439 180
rect 6467 176 6503 204
rect 6531 176 6567 204
rect 6595 176 6631 204
rect 6659 176 6695 204
rect 6723 176 6759 204
rect 6787 176 6823 204
rect 6851 176 6887 204
rect 6915 176 6951 204
rect 6979 176 7015 204
rect 7043 180 7048 204
rect 7076 290 7690 350
rect 7076 262 7081 290
rect 7109 262 7145 290
rect 7173 262 7209 290
rect 7237 262 7273 290
rect 7301 262 7337 290
rect 7365 262 7401 290
rect 7429 262 7465 290
rect 7493 262 7529 290
rect 7557 262 7593 290
rect 7621 262 7657 290
rect 7685 262 7690 290
rect 7076 204 7690 262
rect 7076 180 7081 204
rect 7043 176 7081 180
rect 7109 176 7145 204
rect 7173 176 7209 204
rect 7237 176 7273 204
rect 7301 176 7337 204
rect 7365 176 7401 204
rect 7429 176 7465 204
rect 7493 176 7529 204
rect 7557 176 7593 204
rect 7621 176 7657 204
rect 7685 176 7690 204
rect 5150 163 7690 176
rect 5150 118 5764 163
rect 5150 90 5155 118
rect 5183 90 5219 118
rect 5247 90 5283 118
rect 5311 90 5347 118
rect 5375 90 5411 118
rect 5439 90 5475 118
rect 5503 90 5539 118
rect 5567 90 5603 118
rect 5631 90 5667 118
rect 5695 90 5731 118
rect 5759 90 5764 118
rect 5150 30 5764 90
rect 5792 118 6406 163
rect 5792 90 5797 118
rect 5825 90 5861 118
rect 5889 90 5925 118
rect 5953 90 5989 118
rect 6017 90 6053 118
rect 6081 90 6117 118
rect 6145 90 6181 118
rect 6209 90 6245 118
rect 6273 90 6309 118
rect 6337 90 6373 118
rect 6401 90 6406 118
rect 5792 30 6406 90
rect 6434 118 7048 163
rect 6434 90 6439 118
rect 6467 90 6503 118
rect 6531 90 6567 118
rect 6595 90 6631 118
rect 6659 90 6695 118
rect 6723 90 6759 118
rect 6787 90 6823 118
rect 6851 90 6887 118
rect 6915 90 6951 118
rect 6979 90 7015 118
rect 7043 90 7048 118
rect 6434 30 7048 90
rect 7076 118 7690 163
rect 7076 90 7081 118
rect 7109 90 7145 118
rect 7173 90 7209 118
rect 7237 90 7273 118
rect 7301 90 7337 118
rect 7365 90 7401 118
rect 7429 90 7465 118
rect 7493 90 7529 118
rect 7557 90 7593 118
rect 7621 90 7657 118
rect 7685 90 7690 118
rect 7076 30 7690 90
rect 7718 290 8332 350
rect 7718 262 7723 290
rect 7751 262 7787 290
rect 7815 262 7851 290
rect 7879 262 7915 290
rect 7943 262 7979 290
rect 8007 262 8043 290
rect 8071 262 8107 290
rect 8135 262 8171 290
rect 8199 262 8235 290
rect 8263 262 8299 290
rect 8327 262 8332 290
rect 7718 204 8332 262
rect 7718 176 7723 204
rect 7751 176 7787 204
rect 7815 176 7851 204
rect 7879 176 7915 204
rect 7943 176 7979 204
rect 8007 176 8043 204
rect 8071 176 8107 204
rect 8135 176 8171 204
rect 8199 176 8235 204
rect 8263 176 8299 204
rect 8327 176 8332 204
rect 7718 118 8332 176
rect 7718 90 7723 118
rect 7751 90 7787 118
rect 7815 90 7851 118
rect 7879 90 7915 118
rect 7943 90 7979 118
rect 8007 90 8043 118
rect 8071 90 8107 118
rect 8135 90 8171 118
rect 8199 90 8235 118
rect 8263 90 8299 118
rect 8327 90 8332 118
rect 7718 30 8332 90
rect 8360 290 8974 350
rect 8360 262 8365 290
rect 8393 262 8429 290
rect 8457 262 8493 290
rect 8521 262 8557 290
rect 8585 262 8621 290
rect 8649 262 8685 290
rect 8713 262 8749 290
rect 8777 262 8813 290
rect 8841 262 8877 290
rect 8905 262 8941 290
rect 8969 262 8974 290
rect 8360 204 8974 262
rect 8360 176 8365 204
rect 8393 176 8429 204
rect 8457 176 8493 204
rect 8521 176 8557 204
rect 8585 176 8621 204
rect 8649 176 8685 204
rect 8713 176 8749 204
rect 8777 176 8813 204
rect 8841 176 8877 204
rect 8905 176 8941 204
rect 8969 198 8974 204
rect 9002 290 9616 350
rect 9002 262 9007 290
rect 9035 262 9071 290
rect 9099 262 9135 290
rect 9163 262 9199 290
rect 9227 262 9263 290
rect 9291 262 9327 290
rect 9355 262 9391 290
rect 9419 262 9455 290
rect 9483 262 9519 290
rect 9547 262 9583 290
rect 9611 262 9616 290
rect 9002 204 9616 262
rect 9002 198 9007 204
rect 8969 181 9007 198
rect 8969 176 8974 181
rect 8360 118 8974 176
rect 8360 90 8365 118
rect 8393 90 8429 118
rect 8457 90 8493 118
rect 8521 90 8557 118
rect 8585 90 8621 118
rect 8649 90 8685 118
rect 8713 90 8749 118
rect 8777 90 8813 118
rect 8841 90 8877 118
rect 8905 90 8941 118
rect 8969 90 8974 118
rect 8360 30 8974 90
rect 9002 176 9007 181
rect 9035 176 9071 204
rect 9099 176 9135 204
rect 9163 176 9199 204
rect 9227 176 9263 204
rect 9291 176 9327 204
rect 9355 176 9391 204
rect 9419 176 9455 204
rect 9483 176 9519 204
rect 9547 176 9583 204
rect 9611 198 9616 204
rect 9644 290 10258 350
rect 9644 262 9649 290
rect 9677 262 9713 290
rect 9741 262 9777 290
rect 9805 262 9841 290
rect 9869 262 9905 290
rect 9933 262 9969 290
rect 9997 262 10033 290
rect 10061 262 10097 290
rect 10125 262 10161 290
rect 10189 262 10225 290
rect 10253 262 10258 290
rect 9644 204 10258 262
rect 9644 198 9649 204
rect 9611 181 9649 198
rect 9611 176 9616 181
rect 9002 118 9616 176
rect 9002 90 9007 118
rect 9035 90 9071 118
rect 9099 90 9135 118
rect 9163 90 9199 118
rect 9227 90 9263 118
rect 9291 90 9327 118
rect 9355 90 9391 118
rect 9419 90 9455 118
rect 9483 90 9519 118
rect 9547 90 9583 118
rect 9611 90 9616 118
rect 9002 30 9616 90
rect 9644 176 9649 181
rect 9677 176 9713 204
rect 9741 176 9777 204
rect 9805 176 9841 204
rect 9869 176 9905 204
rect 9933 176 9969 204
rect 9997 176 10033 204
rect 10061 176 10097 204
rect 10125 176 10161 204
rect 10189 176 10225 204
rect 10253 198 10258 204
rect 10286 290 10900 350
rect 10286 262 10291 290
rect 10319 262 10355 290
rect 10383 262 10419 290
rect 10447 262 10483 290
rect 10511 262 10547 290
rect 10575 262 10611 290
rect 10639 262 10675 290
rect 10703 262 10739 290
rect 10767 262 10803 290
rect 10831 262 10867 290
rect 10895 262 10900 290
rect 10286 204 10900 262
rect 10286 198 10291 204
rect 10253 181 10291 198
rect 10253 176 10258 181
rect 9644 118 10258 176
rect 9644 90 9649 118
rect 9677 90 9713 118
rect 9741 90 9777 118
rect 9805 90 9841 118
rect 9869 90 9905 118
rect 9933 90 9969 118
rect 9997 90 10033 118
rect 10061 90 10097 118
rect 10125 90 10161 118
rect 10189 90 10225 118
rect 10253 90 10258 118
rect 9644 30 10258 90
rect 10286 176 10291 181
rect 10319 176 10355 204
rect 10383 176 10419 204
rect 10447 176 10483 204
rect 10511 176 10547 204
rect 10575 176 10611 204
rect 10639 176 10675 204
rect 10703 176 10739 204
rect 10767 176 10803 204
rect 10831 176 10867 204
rect 10895 176 10900 204
rect 10286 118 10900 176
rect 10286 90 10291 118
rect 10319 90 10355 118
rect 10383 90 10419 118
rect 10447 90 10483 118
rect 10511 90 10547 118
rect 10575 90 10611 118
rect 10639 90 10675 118
rect 10703 90 10739 118
rect 10767 90 10803 118
rect 10831 90 10867 118
rect 10895 90 10900 118
rect 10286 30 10900 90
rect 10928 290 11542 350
rect 10928 262 10933 290
rect 10961 262 10997 290
rect 11025 262 11061 290
rect 11089 262 11125 290
rect 11153 262 11189 290
rect 11217 262 11253 290
rect 11281 262 11317 290
rect 11345 262 11381 290
rect 11409 262 11445 290
rect 11473 262 11509 290
rect 11537 262 11542 290
rect 10928 204 11542 262
rect 10928 176 10933 204
rect 10961 176 10997 204
rect 11025 176 11061 204
rect 11089 176 11125 204
rect 11153 176 11189 204
rect 11217 176 11253 204
rect 11281 176 11317 204
rect 11345 176 11381 204
rect 11409 176 11445 204
rect 11473 176 11509 204
rect 11537 176 11542 204
rect 10928 118 11542 176
rect 10928 90 10933 118
rect 10961 90 10997 118
rect 11025 90 11061 118
rect 11089 90 11125 118
rect 11153 90 11189 118
rect 11217 90 11253 118
rect 11281 90 11317 118
rect 11345 90 11381 118
rect 11409 90 11445 118
rect 11473 90 11509 118
rect 11537 90 11542 118
rect 10928 30 11542 90
rect 11570 290 12184 350
rect 11570 262 11575 290
rect 11603 262 11639 290
rect 11667 262 11703 290
rect 11731 262 11767 290
rect 11795 262 11831 290
rect 11859 262 11895 290
rect 11923 262 11959 290
rect 11987 262 12023 290
rect 12051 262 12087 290
rect 12115 262 12151 290
rect 12179 262 12184 290
rect 11570 204 12184 262
rect 11570 176 11575 204
rect 11603 176 11639 204
rect 11667 176 11703 204
rect 11731 176 11767 204
rect 11795 176 11831 204
rect 11859 176 11895 204
rect 11923 176 11959 204
rect 11987 176 12023 204
rect 12051 176 12087 204
rect 12115 176 12151 204
rect 12179 191 12184 204
rect 12212 290 12826 350
rect 12212 262 12217 290
rect 12245 262 12281 290
rect 12309 262 12345 290
rect 12373 262 12409 290
rect 12437 262 12473 290
rect 12501 262 12537 290
rect 12565 262 12601 290
rect 12629 262 12665 290
rect 12693 262 12729 290
rect 12757 262 12793 290
rect 12821 262 12826 290
rect 12212 204 12826 262
rect 12212 191 12217 204
rect 12179 176 12217 191
rect 12245 176 12281 204
rect 12309 176 12345 204
rect 12373 176 12409 204
rect 12437 176 12473 204
rect 12501 176 12537 204
rect 12565 176 12601 204
rect 12629 176 12665 204
rect 12693 176 12729 204
rect 12757 176 12793 204
rect 12821 176 12826 204
rect 11570 174 12826 176
rect 11570 118 12184 174
rect 11570 90 11575 118
rect 11603 90 11639 118
rect 11667 90 11703 118
rect 11731 90 11767 118
rect 11795 90 11831 118
rect 11859 90 11895 118
rect 11923 90 11959 118
rect 11987 90 12023 118
rect 12051 90 12087 118
rect 12115 90 12151 118
rect 12179 90 12184 118
rect 11570 30 12184 90
rect 12212 118 12826 174
rect 12212 90 12217 118
rect 12245 90 12281 118
rect 12309 90 12345 118
rect 12373 90 12409 118
rect 12437 90 12473 118
rect 12501 90 12537 118
rect 12565 90 12601 118
rect 12629 90 12665 118
rect 12693 90 12729 118
rect 12757 90 12793 118
rect 12821 90 12826 118
rect 12212 30 12826 90
<< via2 >>
rect 19 1402 47 1430
rect 83 1402 111 1430
rect 147 1402 175 1430
rect 211 1402 239 1430
rect 275 1402 303 1430
rect 339 1402 367 1430
rect 403 1402 431 1430
rect 467 1402 495 1430
rect 531 1402 559 1430
rect 595 1402 623 1430
rect 19 1316 47 1344
rect 83 1316 111 1344
rect 147 1316 175 1344
rect 211 1316 239 1344
rect 275 1316 303 1344
rect 339 1316 367 1344
rect 403 1316 431 1344
rect 467 1316 495 1344
rect 531 1316 559 1344
rect 595 1316 623 1344
rect 661 1402 689 1430
rect 725 1402 753 1430
rect 789 1402 817 1430
rect 853 1402 881 1430
rect 917 1402 945 1430
rect 981 1402 1009 1430
rect 1045 1402 1073 1430
rect 1109 1402 1137 1430
rect 1173 1402 1201 1430
rect 1237 1402 1265 1430
rect 19 1230 47 1258
rect 83 1230 111 1258
rect 147 1230 175 1258
rect 211 1230 239 1258
rect 275 1230 303 1258
rect 339 1230 367 1258
rect 403 1230 431 1258
rect 467 1230 495 1258
rect 531 1230 559 1258
rect 595 1230 623 1258
rect 661 1316 689 1344
rect 725 1316 753 1344
rect 789 1316 817 1344
rect 853 1316 881 1344
rect 917 1316 945 1344
rect 981 1316 1009 1344
rect 1045 1316 1073 1344
rect 1109 1316 1137 1344
rect 1173 1316 1201 1344
rect 1237 1316 1265 1344
rect 1303 1402 1331 1430
rect 1367 1402 1395 1430
rect 1431 1402 1459 1430
rect 1495 1402 1523 1430
rect 1559 1402 1587 1430
rect 1623 1402 1651 1430
rect 1687 1402 1715 1430
rect 1751 1402 1779 1430
rect 1815 1402 1843 1430
rect 1879 1402 1907 1430
rect 661 1230 689 1258
rect 725 1230 753 1258
rect 789 1230 817 1258
rect 853 1230 881 1258
rect 917 1230 945 1258
rect 981 1230 1009 1258
rect 1045 1230 1073 1258
rect 1109 1230 1137 1258
rect 1173 1230 1201 1258
rect 1237 1230 1265 1258
rect 1303 1316 1331 1344
rect 1367 1316 1395 1344
rect 1431 1316 1459 1344
rect 1495 1316 1523 1344
rect 1559 1316 1587 1344
rect 1623 1316 1651 1344
rect 1687 1316 1715 1344
rect 1751 1316 1779 1344
rect 1815 1316 1843 1344
rect 1879 1316 1907 1344
rect 1945 1402 1973 1430
rect 2009 1402 2037 1430
rect 2073 1402 2101 1430
rect 2137 1402 2165 1430
rect 2201 1402 2229 1430
rect 2265 1402 2293 1430
rect 2329 1402 2357 1430
rect 2393 1402 2421 1430
rect 2457 1402 2485 1430
rect 2521 1402 2549 1430
rect 1303 1230 1331 1258
rect 1367 1230 1395 1258
rect 1431 1230 1459 1258
rect 1495 1230 1523 1258
rect 1559 1230 1587 1258
rect 1623 1230 1651 1258
rect 1687 1230 1715 1258
rect 1751 1230 1779 1258
rect 1815 1230 1843 1258
rect 1879 1230 1907 1258
rect 1945 1316 1973 1344
rect 2009 1316 2037 1344
rect 2073 1316 2101 1344
rect 2137 1316 2165 1344
rect 2201 1316 2229 1344
rect 2265 1316 2293 1344
rect 2329 1316 2357 1344
rect 2393 1316 2421 1344
rect 2457 1316 2485 1344
rect 2521 1316 2549 1344
rect 2587 1402 2615 1430
rect 2651 1402 2679 1430
rect 2715 1402 2743 1430
rect 2779 1402 2807 1430
rect 2843 1402 2871 1430
rect 2907 1402 2935 1430
rect 2971 1402 2999 1430
rect 3035 1402 3063 1430
rect 3099 1402 3127 1430
rect 3163 1402 3191 1430
rect 1945 1230 1973 1258
rect 2009 1230 2037 1258
rect 2073 1230 2101 1258
rect 2137 1230 2165 1258
rect 2201 1230 2229 1258
rect 2265 1230 2293 1258
rect 2329 1230 2357 1258
rect 2393 1230 2421 1258
rect 2457 1230 2485 1258
rect 2521 1230 2549 1258
rect 2587 1316 2615 1344
rect 2651 1316 2679 1344
rect 2715 1316 2743 1344
rect 2779 1316 2807 1344
rect 2843 1316 2871 1344
rect 2907 1316 2935 1344
rect 2971 1316 2999 1344
rect 3035 1316 3063 1344
rect 3099 1316 3127 1344
rect 3163 1316 3191 1344
rect 3229 1402 3257 1430
rect 3293 1402 3321 1430
rect 3357 1402 3385 1430
rect 3421 1402 3449 1430
rect 3485 1402 3513 1430
rect 3549 1402 3577 1430
rect 3613 1402 3641 1430
rect 3677 1402 3705 1430
rect 3741 1402 3769 1430
rect 3805 1402 3833 1430
rect 2587 1230 2615 1258
rect 2651 1230 2679 1258
rect 2715 1230 2743 1258
rect 2779 1230 2807 1258
rect 2843 1230 2871 1258
rect 2907 1230 2935 1258
rect 2971 1230 2999 1258
rect 3035 1230 3063 1258
rect 3099 1230 3127 1258
rect 3163 1230 3191 1258
rect 3229 1316 3257 1344
rect 3293 1316 3321 1344
rect 3357 1316 3385 1344
rect 3421 1316 3449 1344
rect 3485 1316 3513 1344
rect 3549 1316 3577 1344
rect 3613 1316 3641 1344
rect 3677 1316 3705 1344
rect 3741 1316 3769 1344
rect 3805 1316 3833 1344
rect 3871 1402 3899 1430
rect 3935 1402 3963 1430
rect 3999 1402 4027 1430
rect 4063 1402 4091 1430
rect 4127 1402 4155 1430
rect 4191 1402 4219 1430
rect 4255 1402 4283 1430
rect 4319 1402 4347 1430
rect 4383 1402 4411 1430
rect 4447 1402 4475 1430
rect 3229 1230 3257 1258
rect 3293 1230 3321 1258
rect 3357 1230 3385 1258
rect 3421 1230 3449 1258
rect 3485 1230 3513 1258
rect 3549 1230 3577 1258
rect 3613 1230 3641 1258
rect 3677 1230 3705 1258
rect 3741 1230 3769 1258
rect 3805 1230 3833 1258
rect 3871 1316 3899 1344
rect 3935 1316 3963 1344
rect 3999 1316 4027 1344
rect 4063 1316 4091 1344
rect 4127 1316 4155 1344
rect 4191 1316 4219 1344
rect 4255 1316 4283 1344
rect 4319 1316 4347 1344
rect 4383 1316 4411 1344
rect 4447 1316 4475 1344
rect 4513 1402 4541 1430
rect 4577 1402 4605 1430
rect 4641 1402 4669 1430
rect 4705 1402 4733 1430
rect 4769 1402 4797 1430
rect 4833 1402 4861 1430
rect 4897 1402 4925 1430
rect 4961 1402 4989 1430
rect 5025 1402 5053 1430
rect 5089 1402 5117 1430
rect 3871 1230 3899 1258
rect 3935 1230 3963 1258
rect 3999 1230 4027 1258
rect 4063 1230 4091 1258
rect 4127 1230 4155 1258
rect 4191 1230 4219 1258
rect 4255 1230 4283 1258
rect 4319 1230 4347 1258
rect 4383 1230 4411 1258
rect 4447 1230 4475 1258
rect 4513 1316 4541 1344
rect 4577 1316 4605 1344
rect 4641 1316 4669 1344
rect 4705 1316 4733 1344
rect 4769 1316 4797 1344
rect 4833 1316 4861 1344
rect 4897 1316 4925 1344
rect 4961 1316 4989 1344
rect 5025 1316 5053 1344
rect 5089 1316 5117 1344
rect 5155 1402 5183 1430
rect 5219 1402 5247 1430
rect 5283 1402 5311 1430
rect 5347 1402 5375 1430
rect 5411 1402 5439 1430
rect 5475 1402 5503 1430
rect 5539 1402 5567 1430
rect 5603 1402 5631 1430
rect 5667 1402 5695 1430
rect 5731 1402 5759 1430
rect 4513 1230 4541 1258
rect 4577 1230 4605 1258
rect 4641 1230 4669 1258
rect 4705 1230 4733 1258
rect 4769 1230 4797 1258
rect 4833 1230 4861 1258
rect 4897 1230 4925 1258
rect 4961 1230 4989 1258
rect 5025 1230 5053 1258
rect 5089 1230 5117 1258
rect 5155 1316 5183 1344
rect 5219 1316 5247 1344
rect 5283 1316 5311 1344
rect 5347 1316 5375 1344
rect 5411 1316 5439 1344
rect 5475 1316 5503 1344
rect 5539 1316 5567 1344
rect 5603 1316 5631 1344
rect 5667 1316 5695 1344
rect 5731 1316 5759 1344
rect 5797 1402 5825 1430
rect 5861 1402 5889 1430
rect 5925 1402 5953 1430
rect 5989 1402 6017 1430
rect 6053 1402 6081 1430
rect 6117 1402 6145 1430
rect 6181 1402 6209 1430
rect 6245 1402 6273 1430
rect 6309 1402 6337 1430
rect 6373 1402 6401 1430
rect 5155 1230 5183 1258
rect 5219 1230 5247 1258
rect 5283 1230 5311 1258
rect 5347 1230 5375 1258
rect 5411 1230 5439 1258
rect 5475 1230 5503 1258
rect 5539 1230 5567 1258
rect 5603 1230 5631 1258
rect 5667 1230 5695 1258
rect 5731 1230 5759 1258
rect 5797 1316 5825 1344
rect 5861 1316 5889 1344
rect 5925 1316 5953 1344
rect 5989 1316 6017 1344
rect 6053 1316 6081 1344
rect 6117 1316 6145 1344
rect 6181 1316 6209 1344
rect 6245 1316 6273 1344
rect 6309 1316 6337 1344
rect 6373 1316 6401 1344
rect 6439 1402 6467 1430
rect 6503 1402 6531 1430
rect 6567 1402 6595 1430
rect 6631 1402 6659 1430
rect 6695 1402 6723 1430
rect 6759 1402 6787 1430
rect 6823 1402 6851 1430
rect 6887 1402 6915 1430
rect 6951 1402 6979 1430
rect 7015 1402 7043 1430
rect 5797 1230 5825 1258
rect 5861 1230 5889 1258
rect 5925 1230 5953 1258
rect 5989 1230 6017 1258
rect 6053 1230 6081 1258
rect 6117 1230 6145 1258
rect 6181 1230 6209 1258
rect 6245 1230 6273 1258
rect 6309 1230 6337 1258
rect 6373 1230 6401 1258
rect 6439 1316 6467 1344
rect 6503 1316 6531 1344
rect 6567 1316 6595 1344
rect 6631 1316 6659 1344
rect 6695 1316 6723 1344
rect 6759 1316 6787 1344
rect 6823 1316 6851 1344
rect 6887 1316 6915 1344
rect 6951 1316 6979 1344
rect 7015 1316 7043 1344
rect 7081 1402 7109 1430
rect 7145 1402 7173 1430
rect 7209 1402 7237 1430
rect 7273 1402 7301 1430
rect 7337 1402 7365 1430
rect 7401 1402 7429 1430
rect 7465 1402 7493 1430
rect 7529 1402 7557 1430
rect 7593 1402 7621 1430
rect 7657 1402 7685 1430
rect 6439 1230 6467 1258
rect 6503 1230 6531 1258
rect 6567 1230 6595 1258
rect 6631 1230 6659 1258
rect 6695 1230 6723 1258
rect 6759 1230 6787 1258
rect 6823 1230 6851 1258
rect 6887 1230 6915 1258
rect 6951 1230 6979 1258
rect 7015 1230 7043 1258
rect 7081 1316 7109 1344
rect 7145 1316 7173 1344
rect 7209 1316 7237 1344
rect 7273 1316 7301 1344
rect 7337 1316 7365 1344
rect 7401 1316 7429 1344
rect 7465 1316 7493 1344
rect 7529 1316 7557 1344
rect 7593 1316 7621 1344
rect 7657 1316 7685 1344
rect 7723 1402 7751 1430
rect 7787 1402 7815 1430
rect 7851 1402 7879 1430
rect 7915 1402 7943 1430
rect 7979 1402 8007 1430
rect 8043 1402 8071 1430
rect 8107 1402 8135 1430
rect 8171 1402 8199 1430
rect 8235 1402 8263 1430
rect 8299 1402 8327 1430
rect 7081 1230 7109 1258
rect 7145 1230 7173 1258
rect 7209 1230 7237 1258
rect 7273 1230 7301 1258
rect 7337 1230 7365 1258
rect 7401 1230 7429 1258
rect 7465 1230 7493 1258
rect 7529 1230 7557 1258
rect 7593 1230 7621 1258
rect 7657 1230 7685 1258
rect 7723 1316 7751 1344
rect 7787 1316 7815 1344
rect 7851 1316 7879 1344
rect 7915 1316 7943 1344
rect 7979 1316 8007 1344
rect 8043 1316 8071 1344
rect 8107 1316 8135 1344
rect 8171 1316 8199 1344
rect 8235 1316 8263 1344
rect 8299 1316 8327 1344
rect 8365 1402 8393 1430
rect 8429 1402 8457 1430
rect 8493 1402 8521 1430
rect 8557 1402 8585 1430
rect 8621 1402 8649 1430
rect 8685 1402 8713 1430
rect 8749 1402 8777 1430
rect 8813 1402 8841 1430
rect 8877 1402 8905 1430
rect 8941 1402 8969 1430
rect 7723 1230 7751 1258
rect 7787 1230 7815 1258
rect 7851 1230 7879 1258
rect 7915 1230 7943 1258
rect 7979 1230 8007 1258
rect 8043 1230 8071 1258
rect 8107 1230 8135 1258
rect 8171 1230 8199 1258
rect 8235 1230 8263 1258
rect 8299 1230 8327 1258
rect 8365 1316 8393 1344
rect 8429 1316 8457 1344
rect 8493 1316 8521 1344
rect 8557 1316 8585 1344
rect 8621 1316 8649 1344
rect 8685 1316 8713 1344
rect 8749 1316 8777 1344
rect 8813 1316 8841 1344
rect 8877 1316 8905 1344
rect 8941 1316 8969 1344
rect 9007 1402 9035 1430
rect 9071 1402 9099 1430
rect 9135 1402 9163 1430
rect 9199 1402 9227 1430
rect 9263 1402 9291 1430
rect 9327 1402 9355 1430
rect 9391 1402 9419 1430
rect 9455 1402 9483 1430
rect 9519 1402 9547 1430
rect 9583 1402 9611 1430
rect 8365 1230 8393 1258
rect 8429 1230 8457 1258
rect 8493 1230 8521 1258
rect 8557 1230 8585 1258
rect 8621 1230 8649 1258
rect 8685 1230 8713 1258
rect 8749 1230 8777 1258
rect 8813 1230 8841 1258
rect 8877 1230 8905 1258
rect 8941 1230 8969 1258
rect 9007 1316 9035 1344
rect 9071 1316 9099 1344
rect 9135 1316 9163 1344
rect 9199 1316 9227 1344
rect 9263 1316 9291 1344
rect 9327 1316 9355 1344
rect 9391 1316 9419 1344
rect 9455 1316 9483 1344
rect 9519 1316 9547 1344
rect 9583 1316 9611 1344
rect 9649 1402 9677 1430
rect 9713 1402 9741 1430
rect 9777 1402 9805 1430
rect 9841 1402 9869 1430
rect 9905 1402 9933 1430
rect 9969 1402 9997 1430
rect 10033 1402 10061 1430
rect 10097 1402 10125 1430
rect 10161 1402 10189 1430
rect 10225 1402 10253 1430
rect 9007 1230 9035 1258
rect 9071 1230 9099 1258
rect 9135 1230 9163 1258
rect 9199 1230 9227 1258
rect 9263 1230 9291 1258
rect 9327 1230 9355 1258
rect 9391 1230 9419 1258
rect 9455 1230 9483 1258
rect 9519 1230 9547 1258
rect 9583 1230 9611 1258
rect 9649 1316 9677 1344
rect 9713 1316 9741 1344
rect 9777 1316 9805 1344
rect 9841 1316 9869 1344
rect 9905 1316 9933 1344
rect 9969 1316 9997 1344
rect 10033 1316 10061 1344
rect 10097 1316 10125 1344
rect 10161 1316 10189 1344
rect 10225 1316 10253 1344
rect 10291 1402 10319 1430
rect 10355 1402 10383 1430
rect 10419 1402 10447 1430
rect 10483 1402 10511 1430
rect 10547 1402 10575 1430
rect 10611 1402 10639 1430
rect 10675 1402 10703 1430
rect 10739 1402 10767 1430
rect 10803 1402 10831 1430
rect 10867 1402 10895 1430
rect 9649 1230 9677 1258
rect 9713 1230 9741 1258
rect 9777 1230 9805 1258
rect 9841 1230 9869 1258
rect 9905 1230 9933 1258
rect 9969 1230 9997 1258
rect 10033 1230 10061 1258
rect 10097 1230 10125 1258
rect 10161 1230 10189 1258
rect 10225 1230 10253 1258
rect 10291 1316 10319 1344
rect 10355 1316 10383 1344
rect 10419 1316 10447 1344
rect 10483 1316 10511 1344
rect 10547 1316 10575 1344
rect 10611 1316 10639 1344
rect 10675 1316 10703 1344
rect 10739 1316 10767 1344
rect 10803 1316 10831 1344
rect 10867 1316 10895 1344
rect 10933 1402 10961 1430
rect 10997 1402 11025 1430
rect 11061 1402 11089 1430
rect 11125 1402 11153 1430
rect 11189 1402 11217 1430
rect 11253 1402 11281 1430
rect 11317 1402 11345 1430
rect 11381 1402 11409 1430
rect 11445 1402 11473 1430
rect 11509 1402 11537 1430
rect 10291 1230 10319 1258
rect 10355 1230 10383 1258
rect 10419 1230 10447 1258
rect 10483 1230 10511 1258
rect 10547 1230 10575 1258
rect 10611 1230 10639 1258
rect 10675 1230 10703 1258
rect 10739 1230 10767 1258
rect 10803 1230 10831 1258
rect 10867 1230 10895 1258
rect 10933 1316 10961 1344
rect 10997 1316 11025 1344
rect 11061 1316 11089 1344
rect 11125 1316 11153 1344
rect 11189 1316 11217 1344
rect 11253 1316 11281 1344
rect 11317 1316 11345 1344
rect 11381 1316 11409 1344
rect 11445 1316 11473 1344
rect 11509 1316 11537 1344
rect 11575 1402 11603 1430
rect 11639 1402 11667 1430
rect 11703 1402 11731 1430
rect 11767 1402 11795 1430
rect 11831 1402 11859 1430
rect 11895 1402 11923 1430
rect 11959 1402 11987 1430
rect 12023 1402 12051 1430
rect 12087 1402 12115 1430
rect 12151 1402 12179 1430
rect 10933 1230 10961 1258
rect 10997 1230 11025 1258
rect 11061 1230 11089 1258
rect 11125 1230 11153 1258
rect 11189 1230 11217 1258
rect 11253 1230 11281 1258
rect 11317 1230 11345 1258
rect 11381 1230 11409 1258
rect 11445 1230 11473 1258
rect 11509 1230 11537 1258
rect 11575 1316 11603 1344
rect 11639 1316 11667 1344
rect 11703 1316 11731 1344
rect 11767 1316 11795 1344
rect 11831 1316 11859 1344
rect 11895 1316 11923 1344
rect 11959 1316 11987 1344
rect 12023 1316 12051 1344
rect 12087 1316 12115 1344
rect 12151 1316 12179 1344
rect 12217 1402 12245 1430
rect 12281 1402 12309 1430
rect 12345 1402 12373 1430
rect 12409 1402 12437 1430
rect 12473 1402 12501 1430
rect 12537 1402 12565 1430
rect 12601 1402 12629 1430
rect 12665 1402 12693 1430
rect 12729 1402 12757 1430
rect 12793 1402 12821 1430
rect 11575 1230 11603 1258
rect 11639 1230 11667 1258
rect 11703 1230 11731 1258
rect 11767 1230 11795 1258
rect 11831 1230 11859 1258
rect 11895 1230 11923 1258
rect 11959 1230 11987 1258
rect 12023 1230 12051 1258
rect 12087 1230 12115 1258
rect 12151 1230 12179 1258
rect 12217 1316 12245 1344
rect 12281 1316 12309 1344
rect 12345 1316 12373 1344
rect 12409 1316 12437 1344
rect 12473 1316 12501 1344
rect 12537 1316 12565 1344
rect 12601 1316 12629 1344
rect 12665 1316 12693 1344
rect 12729 1316 12757 1344
rect 12793 1316 12821 1344
rect 12217 1230 12245 1258
rect 12281 1230 12309 1258
rect 12345 1230 12373 1258
rect 12409 1230 12437 1258
rect 12473 1230 12501 1258
rect 12537 1230 12565 1258
rect 12601 1230 12629 1258
rect 12665 1230 12693 1258
rect 12729 1230 12757 1258
rect 12793 1230 12821 1258
rect 19 1022 47 1050
rect 83 1022 111 1050
rect 147 1022 175 1050
rect 211 1022 239 1050
rect 275 1022 303 1050
rect 339 1022 367 1050
rect 403 1022 431 1050
rect 467 1022 495 1050
rect 531 1022 559 1050
rect 595 1022 623 1050
rect 19 936 47 964
rect 83 936 111 964
rect 147 936 175 964
rect 211 936 239 964
rect 275 936 303 964
rect 339 936 367 964
rect 403 936 431 964
rect 467 936 495 964
rect 531 936 559 964
rect 595 936 623 964
rect 19 850 47 878
rect 83 850 111 878
rect 147 850 175 878
rect 211 850 239 878
rect 275 850 303 878
rect 339 850 367 878
rect 403 850 431 878
rect 467 850 495 878
rect 531 850 559 878
rect 595 850 623 878
rect 661 1022 689 1050
rect 725 1022 753 1050
rect 789 1022 817 1050
rect 853 1022 881 1050
rect 917 1022 945 1050
rect 981 1022 1009 1050
rect 1045 1022 1073 1050
rect 1109 1022 1137 1050
rect 1173 1022 1201 1050
rect 1237 1022 1265 1050
rect 661 936 689 964
rect 725 936 753 964
rect 789 936 817 964
rect 853 936 881 964
rect 917 936 945 964
rect 981 936 1009 964
rect 1045 936 1073 964
rect 1109 936 1137 964
rect 1173 936 1201 964
rect 1237 936 1265 964
rect 661 850 689 878
rect 725 850 753 878
rect 789 850 817 878
rect 853 850 881 878
rect 917 850 945 878
rect 981 850 1009 878
rect 1045 850 1073 878
rect 1109 850 1137 878
rect 1173 850 1201 878
rect 1237 850 1265 878
rect 1303 1022 1331 1050
rect 1367 1022 1395 1050
rect 1431 1022 1459 1050
rect 1495 1022 1523 1050
rect 1559 1022 1587 1050
rect 1623 1022 1651 1050
rect 1687 1022 1715 1050
rect 1751 1022 1779 1050
rect 1815 1022 1843 1050
rect 1879 1022 1907 1050
rect 1303 936 1331 964
rect 1367 936 1395 964
rect 1431 936 1459 964
rect 1495 936 1523 964
rect 1559 936 1587 964
rect 1623 936 1651 964
rect 1687 936 1715 964
rect 1751 936 1779 964
rect 1815 936 1843 964
rect 1879 936 1907 964
rect 1303 850 1331 878
rect 1367 850 1395 878
rect 1431 850 1459 878
rect 1495 850 1523 878
rect 1559 850 1587 878
rect 1623 850 1651 878
rect 1687 850 1715 878
rect 1751 850 1779 878
rect 1815 850 1843 878
rect 1879 850 1907 878
rect 1945 1022 1973 1050
rect 2009 1022 2037 1050
rect 2073 1022 2101 1050
rect 2137 1022 2165 1050
rect 2201 1022 2229 1050
rect 2265 1022 2293 1050
rect 2329 1022 2357 1050
rect 2393 1022 2421 1050
rect 2457 1022 2485 1050
rect 2521 1022 2549 1050
rect 1945 936 1973 964
rect 2009 936 2037 964
rect 2073 936 2101 964
rect 2137 936 2165 964
rect 2201 936 2229 964
rect 2265 936 2293 964
rect 2329 936 2357 964
rect 2393 936 2421 964
rect 2457 936 2485 964
rect 2521 936 2549 964
rect 1945 850 1973 878
rect 2009 850 2037 878
rect 2073 850 2101 878
rect 2137 850 2165 878
rect 2201 850 2229 878
rect 2265 850 2293 878
rect 2329 850 2357 878
rect 2393 850 2421 878
rect 2457 850 2485 878
rect 2521 850 2549 878
rect 2587 1022 2615 1050
rect 2651 1022 2679 1050
rect 2715 1022 2743 1050
rect 2779 1022 2807 1050
rect 2843 1022 2871 1050
rect 2907 1022 2935 1050
rect 2971 1022 2999 1050
rect 3035 1022 3063 1050
rect 3099 1022 3127 1050
rect 3163 1022 3191 1050
rect 2587 936 2615 964
rect 2651 936 2679 964
rect 2715 936 2743 964
rect 2779 936 2807 964
rect 2843 936 2871 964
rect 2907 936 2935 964
rect 2971 936 2999 964
rect 3035 936 3063 964
rect 3099 936 3127 964
rect 3163 936 3191 964
rect 2587 850 2615 878
rect 2651 850 2679 878
rect 2715 850 2743 878
rect 2779 850 2807 878
rect 2843 850 2871 878
rect 2907 850 2935 878
rect 2971 850 2999 878
rect 3035 850 3063 878
rect 3099 850 3127 878
rect 3163 850 3191 878
rect 3229 1022 3257 1050
rect 3293 1022 3321 1050
rect 3357 1022 3385 1050
rect 3421 1022 3449 1050
rect 3485 1022 3513 1050
rect 3549 1022 3577 1050
rect 3613 1022 3641 1050
rect 3677 1022 3705 1050
rect 3741 1022 3769 1050
rect 3805 1022 3833 1050
rect 3229 936 3257 964
rect 3293 936 3321 964
rect 3357 936 3385 964
rect 3421 936 3449 964
rect 3485 936 3513 964
rect 3549 936 3577 964
rect 3613 936 3641 964
rect 3677 936 3705 964
rect 3741 936 3769 964
rect 3805 936 3833 964
rect 3229 850 3257 878
rect 3293 850 3321 878
rect 3357 850 3385 878
rect 3421 850 3449 878
rect 3485 850 3513 878
rect 3549 850 3577 878
rect 3613 850 3641 878
rect 3677 850 3705 878
rect 3741 850 3769 878
rect 3805 850 3833 878
rect 3871 1022 3899 1050
rect 3935 1022 3963 1050
rect 3999 1022 4027 1050
rect 4063 1022 4091 1050
rect 4127 1022 4155 1050
rect 4191 1022 4219 1050
rect 4255 1022 4283 1050
rect 4319 1022 4347 1050
rect 4383 1022 4411 1050
rect 4447 1022 4475 1050
rect 3871 936 3899 964
rect 3935 936 3963 964
rect 3999 936 4027 964
rect 4063 936 4091 964
rect 4127 936 4155 964
rect 4191 936 4219 964
rect 4255 936 4283 964
rect 4319 936 4347 964
rect 4383 936 4411 964
rect 4447 936 4475 964
rect 3871 850 3899 878
rect 3935 850 3963 878
rect 3999 850 4027 878
rect 4063 850 4091 878
rect 4127 850 4155 878
rect 4191 850 4219 878
rect 4255 850 4283 878
rect 4319 850 4347 878
rect 4383 850 4411 878
rect 4447 850 4475 878
rect 4513 1022 4541 1050
rect 4577 1022 4605 1050
rect 4641 1022 4669 1050
rect 4705 1022 4733 1050
rect 4769 1022 4797 1050
rect 4833 1022 4861 1050
rect 4897 1022 4925 1050
rect 4961 1022 4989 1050
rect 5025 1022 5053 1050
rect 5089 1022 5117 1050
rect 4513 936 4541 964
rect 4577 936 4605 964
rect 4641 936 4669 964
rect 4705 936 4733 964
rect 4769 936 4797 964
rect 4833 936 4861 964
rect 4897 936 4925 964
rect 4961 936 4989 964
rect 5025 936 5053 964
rect 5089 936 5117 964
rect 4513 850 4541 878
rect 4577 850 4605 878
rect 4641 850 4669 878
rect 4705 850 4733 878
rect 4769 850 4797 878
rect 4833 850 4861 878
rect 4897 850 4925 878
rect 4961 850 4989 878
rect 5025 850 5053 878
rect 5089 850 5117 878
rect 5155 1022 5183 1050
rect 5219 1022 5247 1050
rect 5283 1022 5311 1050
rect 5347 1022 5375 1050
rect 5411 1022 5439 1050
rect 5475 1022 5503 1050
rect 5539 1022 5567 1050
rect 5603 1022 5631 1050
rect 5667 1022 5695 1050
rect 5731 1022 5759 1050
rect 5155 936 5183 964
rect 5219 936 5247 964
rect 5283 936 5311 964
rect 5347 936 5375 964
rect 5411 936 5439 964
rect 5475 936 5503 964
rect 5539 936 5567 964
rect 5603 936 5631 964
rect 5667 936 5695 964
rect 5731 936 5759 964
rect 5155 850 5183 878
rect 5219 850 5247 878
rect 5283 850 5311 878
rect 5347 850 5375 878
rect 5411 850 5439 878
rect 5475 850 5503 878
rect 5539 850 5567 878
rect 5603 850 5631 878
rect 5667 850 5695 878
rect 5731 850 5759 878
rect 5797 1022 5825 1050
rect 5861 1022 5889 1050
rect 5925 1022 5953 1050
rect 5989 1022 6017 1050
rect 6053 1022 6081 1050
rect 6117 1022 6145 1050
rect 6181 1022 6209 1050
rect 6245 1022 6273 1050
rect 6309 1022 6337 1050
rect 6373 1022 6401 1050
rect 5797 936 5825 964
rect 5861 936 5889 964
rect 5925 936 5953 964
rect 5989 936 6017 964
rect 6053 936 6081 964
rect 6117 936 6145 964
rect 6181 936 6209 964
rect 6245 936 6273 964
rect 6309 936 6337 964
rect 6373 936 6401 964
rect 5797 850 5825 878
rect 5861 850 5889 878
rect 5925 850 5953 878
rect 5989 850 6017 878
rect 6053 850 6081 878
rect 6117 850 6145 878
rect 6181 850 6209 878
rect 6245 850 6273 878
rect 6309 850 6337 878
rect 6373 850 6401 878
rect 6439 1022 6467 1050
rect 6503 1022 6531 1050
rect 6567 1022 6595 1050
rect 6631 1022 6659 1050
rect 6695 1022 6723 1050
rect 6759 1022 6787 1050
rect 6823 1022 6851 1050
rect 6887 1022 6915 1050
rect 6951 1022 6979 1050
rect 7015 1022 7043 1050
rect 6439 936 6467 964
rect 6503 936 6531 964
rect 6567 936 6595 964
rect 6631 936 6659 964
rect 6695 936 6723 964
rect 6759 936 6787 964
rect 6823 936 6851 964
rect 6887 936 6915 964
rect 6951 936 6979 964
rect 7015 936 7043 964
rect 6439 850 6467 878
rect 6503 850 6531 878
rect 6567 850 6595 878
rect 6631 850 6659 878
rect 6695 850 6723 878
rect 6759 850 6787 878
rect 6823 850 6851 878
rect 6887 850 6915 878
rect 6951 850 6979 878
rect 7015 850 7043 878
rect 7081 1022 7109 1050
rect 7145 1022 7173 1050
rect 7209 1022 7237 1050
rect 7273 1022 7301 1050
rect 7337 1022 7365 1050
rect 7401 1022 7429 1050
rect 7465 1022 7493 1050
rect 7529 1022 7557 1050
rect 7593 1022 7621 1050
rect 7657 1022 7685 1050
rect 7081 936 7109 964
rect 7145 936 7173 964
rect 7209 936 7237 964
rect 7273 936 7301 964
rect 7337 936 7365 964
rect 7401 936 7429 964
rect 7465 936 7493 964
rect 7529 936 7557 964
rect 7593 936 7621 964
rect 7657 936 7685 964
rect 7081 850 7109 878
rect 7145 850 7173 878
rect 7209 850 7237 878
rect 7273 850 7301 878
rect 7337 850 7365 878
rect 7401 850 7429 878
rect 7465 850 7493 878
rect 7529 850 7557 878
rect 7593 850 7621 878
rect 7657 850 7685 878
rect 7723 1022 7751 1050
rect 7787 1022 7815 1050
rect 7851 1022 7879 1050
rect 7915 1022 7943 1050
rect 7979 1022 8007 1050
rect 8043 1022 8071 1050
rect 8107 1022 8135 1050
rect 8171 1022 8199 1050
rect 8235 1022 8263 1050
rect 8299 1022 8327 1050
rect 7723 936 7751 964
rect 7787 936 7815 964
rect 7851 936 7879 964
rect 7915 936 7943 964
rect 7979 936 8007 964
rect 8043 936 8071 964
rect 8107 936 8135 964
rect 8171 936 8199 964
rect 8235 936 8263 964
rect 8299 936 8327 964
rect 7723 850 7751 878
rect 7787 850 7815 878
rect 7851 850 7879 878
rect 7915 850 7943 878
rect 7979 850 8007 878
rect 8043 850 8071 878
rect 8107 850 8135 878
rect 8171 850 8199 878
rect 8235 850 8263 878
rect 8299 850 8327 878
rect 8365 1022 8393 1050
rect 8429 1022 8457 1050
rect 8493 1022 8521 1050
rect 8557 1022 8585 1050
rect 8621 1022 8649 1050
rect 8685 1022 8713 1050
rect 8749 1022 8777 1050
rect 8813 1022 8841 1050
rect 8877 1022 8905 1050
rect 8941 1022 8969 1050
rect 8365 936 8393 964
rect 8429 936 8457 964
rect 8493 936 8521 964
rect 8557 936 8585 964
rect 8621 936 8649 964
rect 8685 936 8713 964
rect 8749 936 8777 964
rect 8813 936 8841 964
rect 8877 936 8905 964
rect 8941 936 8969 964
rect 8365 850 8393 878
rect 8429 850 8457 878
rect 8493 850 8521 878
rect 8557 850 8585 878
rect 8621 850 8649 878
rect 8685 850 8713 878
rect 8749 850 8777 878
rect 8813 850 8841 878
rect 8877 850 8905 878
rect 8941 850 8969 878
rect 9007 1022 9035 1050
rect 9071 1022 9099 1050
rect 9135 1022 9163 1050
rect 9199 1022 9227 1050
rect 9263 1022 9291 1050
rect 9327 1022 9355 1050
rect 9391 1022 9419 1050
rect 9455 1022 9483 1050
rect 9519 1022 9547 1050
rect 9583 1022 9611 1050
rect 9007 936 9035 964
rect 9071 936 9099 964
rect 9135 936 9163 964
rect 9199 936 9227 964
rect 9263 936 9291 964
rect 9327 936 9355 964
rect 9391 936 9419 964
rect 9455 936 9483 964
rect 9519 936 9547 964
rect 9583 936 9611 964
rect 9007 850 9035 878
rect 9071 850 9099 878
rect 9135 850 9163 878
rect 9199 850 9227 878
rect 9263 850 9291 878
rect 9327 850 9355 878
rect 9391 850 9419 878
rect 9455 850 9483 878
rect 9519 850 9547 878
rect 9583 850 9611 878
rect 9649 1022 9677 1050
rect 9713 1022 9741 1050
rect 9777 1022 9805 1050
rect 9841 1022 9869 1050
rect 9905 1022 9933 1050
rect 9969 1022 9997 1050
rect 10033 1022 10061 1050
rect 10097 1022 10125 1050
rect 10161 1022 10189 1050
rect 10225 1022 10253 1050
rect 9649 936 9677 964
rect 9713 936 9741 964
rect 9777 936 9805 964
rect 9841 936 9869 964
rect 9905 936 9933 964
rect 9969 936 9997 964
rect 10033 936 10061 964
rect 10097 936 10125 964
rect 10161 936 10189 964
rect 10225 936 10253 964
rect 9649 850 9677 878
rect 9713 850 9741 878
rect 9777 850 9805 878
rect 9841 850 9869 878
rect 9905 850 9933 878
rect 9969 850 9997 878
rect 10033 850 10061 878
rect 10097 850 10125 878
rect 10161 850 10189 878
rect 10225 850 10253 878
rect 10291 1022 10319 1050
rect 10355 1022 10383 1050
rect 10419 1022 10447 1050
rect 10483 1022 10511 1050
rect 10547 1022 10575 1050
rect 10611 1022 10639 1050
rect 10675 1022 10703 1050
rect 10739 1022 10767 1050
rect 10803 1022 10831 1050
rect 10867 1022 10895 1050
rect 10291 936 10319 964
rect 10355 936 10383 964
rect 10419 936 10447 964
rect 10483 936 10511 964
rect 10547 936 10575 964
rect 10611 936 10639 964
rect 10675 936 10703 964
rect 10739 936 10767 964
rect 10803 936 10831 964
rect 10867 936 10895 964
rect 10291 850 10319 878
rect 10355 850 10383 878
rect 10419 850 10447 878
rect 10483 850 10511 878
rect 10547 850 10575 878
rect 10611 850 10639 878
rect 10675 850 10703 878
rect 10739 850 10767 878
rect 10803 850 10831 878
rect 10867 850 10895 878
rect 10933 1022 10961 1050
rect 10997 1022 11025 1050
rect 11061 1022 11089 1050
rect 11125 1022 11153 1050
rect 11189 1022 11217 1050
rect 11253 1022 11281 1050
rect 11317 1022 11345 1050
rect 11381 1022 11409 1050
rect 11445 1022 11473 1050
rect 11509 1022 11537 1050
rect 10933 936 10961 964
rect 10997 936 11025 964
rect 11061 936 11089 964
rect 11125 936 11153 964
rect 11189 936 11217 964
rect 11253 936 11281 964
rect 11317 936 11345 964
rect 11381 936 11409 964
rect 11445 936 11473 964
rect 11509 936 11537 964
rect 10933 850 10961 878
rect 10997 850 11025 878
rect 11061 850 11089 878
rect 11125 850 11153 878
rect 11189 850 11217 878
rect 11253 850 11281 878
rect 11317 850 11345 878
rect 11381 850 11409 878
rect 11445 850 11473 878
rect 11509 850 11537 878
rect 11575 1022 11603 1050
rect 11639 1022 11667 1050
rect 11703 1022 11731 1050
rect 11767 1022 11795 1050
rect 11831 1022 11859 1050
rect 11895 1022 11923 1050
rect 11959 1022 11987 1050
rect 12023 1022 12051 1050
rect 12087 1022 12115 1050
rect 12151 1022 12179 1050
rect 11575 936 11603 964
rect 11639 936 11667 964
rect 11703 936 11731 964
rect 11767 936 11795 964
rect 11831 936 11859 964
rect 11895 936 11923 964
rect 11959 936 11987 964
rect 12023 936 12051 964
rect 12087 936 12115 964
rect 12151 936 12179 964
rect 11575 850 11603 878
rect 11639 850 11667 878
rect 11703 850 11731 878
rect 11767 850 11795 878
rect 11831 850 11859 878
rect 11895 850 11923 878
rect 11959 850 11987 878
rect 12023 850 12051 878
rect 12087 850 12115 878
rect 12151 850 12179 878
rect 12217 1022 12245 1050
rect 12281 1022 12309 1050
rect 12345 1022 12373 1050
rect 12409 1022 12437 1050
rect 12473 1022 12501 1050
rect 12537 1022 12565 1050
rect 12601 1022 12629 1050
rect 12665 1022 12693 1050
rect 12729 1022 12757 1050
rect 12793 1022 12821 1050
rect 12217 936 12245 964
rect 12281 936 12309 964
rect 12345 936 12373 964
rect 12409 936 12437 964
rect 12473 936 12501 964
rect 12537 936 12565 964
rect 12601 936 12629 964
rect 12665 936 12693 964
rect 12729 936 12757 964
rect 12793 936 12821 964
rect 12217 850 12245 878
rect 12281 850 12309 878
rect 12345 850 12373 878
rect 12409 850 12437 878
rect 12473 850 12501 878
rect 12537 850 12565 878
rect 12601 850 12629 878
rect 12665 850 12693 878
rect 12729 850 12757 878
rect 12793 850 12821 878
rect 19 642 47 670
rect 83 642 111 670
rect 147 642 175 670
rect 211 642 239 670
rect 275 642 303 670
rect 339 642 367 670
rect 403 642 431 670
rect 467 642 495 670
rect 531 642 559 670
rect 595 642 623 670
rect 19 556 47 584
rect 83 556 111 584
rect 147 556 175 584
rect 211 556 239 584
rect 275 556 303 584
rect 339 556 367 584
rect 403 556 431 584
rect 467 556 495 584
rect 531 556 559 584
rect 595 556 623 584
rect 19 470 47 498
rect 83 470 111 498
rect 147 470 175 498
rect 211 470 239 498
rect 275 470 303 498
rect 339 470 367 498
rect 403 470 431 498
rect 467 470 495 498
rect 531 470 559 498
rect 595 470 623 498
rect 661 642 689 670
rect 725 642 753 670
rect 789 642 817 670
rect 853 642 881 670
rect 917 642 945 670
rect 981 642 1009 670
rect 1045 642 1073 670
rect 1109 642 1137 670
rect 1173 642 1201 670
rect 1237 642 1265 670
rect 661 556 689 584
rect 725 556 753 584
rect 789 556 817 584
rect 853 556 881 584
rect 917 556 945 584
rect 981 556 1009 584
rect 1045 556 1073 584
rect 1109 556 1137 584
rect 1173 556 1201 584
rect 1237 556 1265 584
rect 661 470 689 498
rect 725 470 753 498
rect 789 470 817 498
rect 853 470 881 498
rect 917 470 945 498
rect 981 470 1009 498
rect 1045 470 1073 498
rect 1109 470 1137 498
rect 1173 470 1201 498
rect 1237 470 1265 498
rect 1303 642 1331 670
rect 1367 642 1395 670
rect 1431 642 1459 670
rect 1495 642 1523 670
rect 1559 642 1587 670
rect 1623 642 1651 670
rect 1687 642 1715 670
rect 1751 642 1779 670
rect 1815 642 1843 670
rect 1879 642 1907 670
rect 1303 556 1331 584
rect 1367 556 1395 584
rect 1431 556 1459 584
rect 1495 556 1523 584
rect 1559 556 1587 584
rect 1623 556 1651 584
rect 1687 556 1715 584
rect 1751 556 1779 584
rect 1815 556 1843 584
rect 1879 556 1907 584
rect 1303 470 1331 498
rect 1367 470 1395 498
rect 1431 470 1459 498
rect 1495 470 1523 498
rect 1559 470 1587 498
rect 1623 470 1651 498
rect 1687 470 1715 498
rect 1751 470 1779 498
rect 1815 470 1843 498
rect 1879 470 1907 498
rect 1945 642 1973 670
rect 2009 642 2037 670
rect 2073 642 2101 670
rect 2137 642 2165 670
rect 2201 642 2229 670
rect 2265 642 2293 670
rect 2329 642 2357 670
rect 2393 642 2421 670
rect 2457 642 2485 670
rect 2521 642 2549 670
rect 1945 556 1973 584
rect 2009 556 2037 584
rect 2073 556 2101 584
rect 2137 556 2165 584
rect 2201 556 2229 584
rect 2265 556 2293 584
rect 2329 556 2357 584
rect 2393 556 2421 584
rect 2457 556 2485 584
rect 2521 556 2549 584
rect 1945 470 1973 498
rect 2009 470 2037 498
rect 2073 470 2101 498
rect 2137 470 2165 498
rect 2201 470 2229 498
rect 2265 470 2293 498
rect 2329 470 2357 498
rect 2393 470 2421 498
rect 2457 470 2485 498
rect 2521 470 2549 498
rect 2587 642 2615 670
rect 2651 642 2679 670
rect 2715 642 2743 670
rect 2779 642 2807 670
rect 2843 642 2871 670
rect 2907 642 2935 670
rect 2971 642 2999 670
rect 3035 642 3063 670
rect 3099 642 3127 670
rect 3163 642 3191 670
rect 2587 556 2615 584
rect 2651 556 2679 584
rect 2715 556 2743 584
rect 2779 556 2807 584
rect 2843 556 2871 584
rect 2907 556 2935 584
rect 2971 556 2999 584
rect 3035 556 3063 584
rect 3099 556 3127 584
rect 3163 556 3191 584
rect 2587 470 2615 498
rect 2651 470 2679 498
rect 2715 470 2743 498
rect 2779 470 2807 498
rect 2843 470 2871 498
rect 2907 470 2935 498
rect 2971 470 2999 498
rect 3035 470 3063 498
rect 3099 470 3127 498
rect 3163 470 3191 498
rect 3229 642 3257 670
rect 3293 642 3321 670
rect 3357 642 3385 670
rect 3421 642 3449 670
rect 3485 642 3513 670
rect 3549 642 3577 670
rect 3613 642 3641 670
rect 3677 642 3705 670
rect 3741 642 3769 670
rect 3805 642 3833 670
rect 3229 556 3257 584
rect 3293 556 3321 584
rect 3357 556 3385 584
rect 3421 556 3449 584
rect 3485 556 3513 584
rect 3549 556 3577 584
rect 3613 556 3641 584
rect 3677 556 3705 584
rect 3741 556 3769 584
rect 3805 556 3833 584
rect 3229 470 3257 498
rect 3293 470 3321 498
rect 3357 470 3385 498
rect 3421 470 3449 498
rect 3485 470 3513 498
rect 3549 470 3577 498
rect 3613 470 3641 498
rect 3677 470 3705 498
rect 3741 470 3769 498
rect 3805 470 3833 498
rect 3871 642 3899 670
rect 3935 642 3963 670
rect 3999 642 4027 670
rect 4063 642 4091 670
rect 4127 642 4155 670
rect 4191 642 4219 670
rect 4255 642 4283 670
rect 4319 642 4347 670
rect 4383 642 4411 670
rect 4447 642 4475 670
rect 3871 556 3899 584
rect 3935 556 3963 584
rect 3999 556 4027 584
rect 4063 556 4091 584
rect 4127 556 4155 584
rect 4191 556 4219 584
rect 4255 556 4283 584
rect 4319 556 4347 584
rect 4383 556 4411 584
rect 4447 556 4475 584
rect 3871 470 3899 498
rect 3935 470 3963 498
rect 3999 470 4027 498
rect 4063 470 4091 498
rect 4127 470 4155 498
rect 4191 470 4219 498
rect 4255 470 4283 498
rect 4319 470 4347 498
rect 4383 470 4411 498
rect 4447 470 4475 498
rect 4513 642 4541 670
rect 4577 642 4605 670
rect 4641 642 4669 670
rect 4705 642 4733 670
rect 4769 642 4797 670
rect 4833 642 4861 670
rect 4897 642 4925 670
rect 4961 642 4989 670
rect 5025 642 5053 670
rect 5089 642 5117 670
rect 4513 556 4541 584
rect 4577 556 4605 584
rect 4641 556 4669 584
rect 4705 556 4733 584
rect 4769 556 4797 584
rect 4833 556 4861 584
rect 4897 556 4925 584
rect 4961 556 4989 584
rect 5025 556 5053 584
rect 5089 556 5117 584
rect 4513 470 4541 498
rect 4577 470 4605 498
rect 4641 470 4669 498
rect 4705 470 4733 498
rect 4769 470 4797 498
rect 4833 470 4861 498
rect 4897 470 4925 498
rect 4961 470 4989 498
rect 5025 470 5053 498
rect 5089 470 5117 498
rect 5155 642 5183 670
rect 5219 642 5247 670
rect 5283 642 5311 670
rect 5347 642 5375 670
rect 5411 642 5439 670
rect 5475 642 5503 670
rect 5539 642 5567 670
rect 5603 642 5631 670
rect 5667 642 5695 670
rect 5731 642 5759 670
rect 5155 556 5183 584
rect 5219 556 5247 584
rect 5283 556 5311 584
rect 5347 556 5375 584
rect 5411 556 5439 584
rect 5475 556 5503 584
rect 5539 556 5567 584
rect 5603 556 5631 584
rect 5667 556 5695 584
rect 5731 556 5759 584
rect 5155 470 5183 498
rect 5219 470 5247 498
rect 5283 470 5311 498
rect 5347 470 5375 498
rect 5411 470 5439 498
rect 5475 470 5503 498
rect 5539 470 5567 498
rect 5603 470 5631 498
rect 5667 470 5695 498
rect 5731 470 5759 498
rect 5797 642 5825 670
rect 5861 642 5889 670
rect 5925 642 5953 670
rect 5989 642 6017 670
rect 6053 642 6081 670
rect 6117 642 6145 670
rect 6181 642 6209 670
rect 6245 642 6273 670
rect 6309 642 6337 670
rect 6373 642 6401 670
rect 5797 556 5825 584
rect 5861 556 5889 584
rect 5925 556 5953 584
rect 5989 556 6017 584
rect 6053 556 6081 584
rect 6117 556 6145 584
rect 6181 556 6209 584
rect 6245 556 6273 584
rect 6309 556 6337 584
rect 6373 556 6401 584
rect 5797 470 5825 498
rect 5861 470 5889 498
rect 5925 470 5953 498
rect 5989 470 6017 498
rect 6053 470 6081 498
rect 6117 470 6145 498
rect 6181 470 6209 498
rect 6245 470 6273 498
rect 6309 470 6337 498
rect 6373 470 6401 498
rect 6439 642 6467 670
rect 6503 642 6531 670
rect 6567 642 6595 670
rect 6631 642 6659 670
rect 6695 642 6723 670
rect 6759 642 6787 670
rect 6823 642 6851 670
rect 6887 642 6915 670
rect 6951 642 6979 670
rect 7015 642 7043 670
rect 6439 556 6467 584
rect 6503 556 6531 584
rect 6567 556 6595 584
rect 6631 556 6659 584
rect 6695 556 6723 584
rect 6759 556 6787 584
rect 6823 556 6851 584
rect 6887 556 6915 584
rect 6951 556 6979 584
rect 7015 556 7043 584
rect 6439 470 6467 498
rect 6503 470 6531 498
rect 6567 470 6595 498
rect 6631 470 6659 498
rect 6695 470 6723 498
rect 6759 470 6787 498
rect 6823 470 6851 498
rect 6887 470 6915 498
rect 6951 470 6979 498
rect 7015 470 7043 498
rect 7081 642 7109 670
rect 7145 642 7173 670
rect 7209 642 7237 670
rect 7273 642 7301 670
rect 7337 642 7365 670
rect 7401 642 7429 670
rect 7465 642 7493 670
rect 7529 642 7557 670
rect 7593 642 7621 670
rect 7657 642 7685 670
rect 7081 556 7109 584
rect 7145 556 7173 584
rect 7209 556 7237 584
rect 7273 556 7301 584
rect 7337 556 7365 584
rect 7401 556 7429 584
rect 7465 556 7493 584
rect 7529 556 7557 584
rect 7593 556 7621 584
rect 7657 556 7685 584
rect 7081 470 7109 498
rect 7145 470 7173 498
rect 7209 470 7237 498
rect 7273 470 7301 498
rect 7337 470 7365 498
rect 7401 470 7429 498
rect 7465 470 7493 498
rect 7529 470 7557 498
rect 7593 470 7621 498
rect 7657 470 7685 498
rect 7723 642 7751 670
rect 7787 642 7815 670
rect 7851 642 7879 670
rect 7915 642 7943 670
rect 7979 642 8007 670
rect 8043 642 8071 670
rect 8107 642 8135 670
rect 8171 642 8199 670
rect 8235 642 8263 670
rect 8299 642 8327 670
rect 7723 556 7751 584
rect 7787 556 7815 584
rect 7851 556 7879 584
rect 7915 556 7943 584
rect 7979 556 8007 584
rect 8043 556 8071 584
rect 8107 556 8135 584
rect 8171 556 8199 584
rect 8235 556 8263 584
rect 8299 556 8327 584
rect 7723 470 7751 498
rect 7787 470 7815 498
rect 7851 470 7879 498
rect 7915 470 7943 498
rect 7979 470 8007 498
rect 8043 470 8071 498
rect 8107 470 8135 498
rect 8171 470 8199 498
rect 8235 470 8263 498
rect 8299 470 8327 498
rect 8365 642 8393 670
rect 8429 642 8457 670
rect 8493 642 8521 670
rect 8557 642 8585 670
rect 8621 642 8649 670
rect 8685 642 8713 670
rect 8749 642 8777 670
rect 8813 642 8841 670
rect 8877 642 8905 670
rect 8941 642 8969 670
rect 8365 556 8393 584
rect 8429 556 8457 584
rect 8493 556 8521 584
rect 8557 556 8585 584
rect 8621 556 8649 584
rect 8685 556 8713 584
rect 8749 556 8777 584
rect 8813 556 8841 584
rect 8877 556 8905 584
rect 8941 556 8969 584
rect 8365 470 8393 498
rect 8429 470 8457 498
rect 8493 470 8521 498
rect 8557 470 8585 498
rect 8621 470 8649 498
rect 8685 470 8713 498
rect 8749 470 8777 498
rect 8813 470 8841 498
rect 8877 470 8905 498
rect 8941 470 8969 498
rect 9007 642 9035 670
rect 9071 642 9099 670
rect 9135 642 9163 670
rect 9199 642 9227 670
rect 9263 642 9291 670
rect 9327 642 9355 670
rect 9391 642 9419 670
rect 9455 642 9483 670
rect 9519 642 9547 670
rect 9583 642 9611 670
rect 9007 556 9035 584
rect 9071 556 9099 584
rect 9135 556 9163 584
rect 9199 556 9227 584
rect 9263 556 9291 584
rect 9327 556 9355 584
rect 9391 556 9419 584
rect 9455 556 9483 584
rect 9519 556 9547 584
rect 9583 556 9611 584
rect 9007 470 9035 498
rect 9071 470 9099 498
rect 9135 470 9163 498
rect 9199 470 9227 498
rect 9263 470 9291 498
rect 9327 470 9355 498
rect 9391 470 9419 498
rect 9455 470 9483 498
rect 9519 470 9547 498
rect 9583 470 9611 498
rect 9649 642 9677 670
rect 9713 642 9741 670
rect 9777 642 9805 670
rect 9841 642 9869 670
rect 9905 642 9933 670
rect 9969 642 9997 670
rect 10033 642 10061 670
rect 10097 642 10125 670
rect 10161 642 10189 670
rect 10225 642 10253 670
rect 9649 556 9677 584
rect 9713 556 9741 584
rect 9777 556 9805 584
rect 9841 556 9869 584
rect 9905 556 9933 584
rect 9969 556 9997 584
rect 10033 556 10061 584
rect 10097 556 10125 584
rect 10161 556 10189 584
rect 10225 556 10253 584
rect 9649 470 9677 498
rect 9713 470 9741 498
rect 9777 470 9805 498
rect 9841 470 9869 498
rect 9905 470 9933 498
rect 9969 470 9997 498
rect 10033 470 10061 498
rect 10097 470 10125 498
rect 10161 470 10189 498
rect 10225 470 10253 498
rect 10291 642 10319 670
rect 10355 642 10383 670
rect 10419 642 10447 670
rect 10483 642 10511 670
rect 10547 642 10575 670
rect 10611 642 10639 670
rect 10675 642 10703 670
rect 10739 642 10767 670
rect 10803 642 10831 670
rect 10867 642 10895 670
rect 10291 556 10319 584
rect 10355 556 10383 584
rect 10419 556 10447 584
rect 10483 556 10511 584
rect 10547 556 10575 584
rect 10611 556 10639 584
rect 10675 556 10703 584
rect 10739 556 10767 584
rect 10803 556 10831 584
rect 10867 556 10895 584
rect 10291 470 10319 498
rect 10355 470 10383 498
rect 10419 470 10447 498
rect 10483 470 10511 498
rect 10547 470 10575 498
rect 10611 470 10639 498
rect 10675 470 10703 498
rect 10739 470 10767 498
rect 10803 470 10831 498
rect 10867 470 10895 498
rect 10933 642 10961 670
rect 10997 642 11025 670
rect 11061 642 11089 670
rect 11125 642 11153 670
rect 11189 642 11217 670
rect 11253 642 11281 670
rect 11317 642 11345 670
rect 11381 642 11409 670
rect 11445 642 11473 670
rect 11509 642 11537 670
rect 10933 556 10961 584
rect 10997 556 11025 584
rect 11061 556 11089 584
rect 11125 556 11153 584
rect 11189 556 11217 584
rect 11253 556 11281 584
rect 11317 556 11345 584
rect 11381 556 11409 584
rect 11445 556 11473 584
rect 11509 556 11537 584
rect 10933 470 10961 498
rect 10997 470 11025 498
rect 11061 470 11089 498
rect 11125 470 11153 498
rect 11189 470 11217 498
rect 11253 470 11281 498
rect 11317 470 11345 498
rect 11381 470 11409 498
rect 11445 470 11473 498
rect 11509 470 11537 498
rect 11575 642 11603 670
rect 11639 642 11667 670
rect 11703 642 11731 670
rect 11767 642 11795 670
rect 11831 642 11859 670
rect 11895 642 11923 670
rect 11959 642 11987 670
rect 12023 642 12051 670
rect 12087 642 12115 670
rect 12151 642 12179 670
rect 11575 556 11603 584
rect 11639 556 11667 584
rect 11703 556 11731 584
rect 11767 556 11795 584
rect 11831 556 11859 584
rect 11895 556 11923 584
rect 11959 556 11987 584
rect 12023 556 12051 584
rect 12087 556 12115 584
rect 12151 556 12179 584
rect 11575 470 11603 498
rect 11639 470 11667 498
rect 11703 470 11731 498
rect 11767 470 11795 498
rect 11831 470 11859 498
rect 11895 470 11923 498
rect 11959 470 11987 498
rect 12023 470 12051 498
rect 12087 470 12115 498
rect 12151 470 12179 498
rect 12217 642 12245 670
rect 12281 642 12309 670
rect 12345 642 12373 670
rect 12409 642 12437 670
rect 12473 642 12501 670
rect 12537 642 12565 670
rect 12601 642 12629 670
rect 12665 642 12693 670
rect 12729 642 12757 670
rect 12793 642 12821 670
rect 12217 556 12245 584
rect 12281 556 12309 584
rect 12345 556 12373 584
rect 12409 556 12437 584
rect 12473 556 12501 584
rect 12537 556 12565 584
rect 12601 556 12629 584
rect 12665 556 12693 584
rect 12729 556 12757 584
rect 12793 556 12821 584
rect 12217 470 12245 498
rect 12281 470 12309 498
rect 12345 470 12373 498
rect 12409 470 12437 498
rect 12473 470 12501 498
rect 12537 470 12565 498
rect 12601 470 12629 498
rect 12665 470 12693 498
rect 12729 470 12757 498
rect 12793 470 12821 498
rect 19 262 47 290
rect 83 262 111 290
rect 147 262 175 290
rect 211 262 239 290
rect 275 262 303 290
rect 339 262 367 290
rect 403 262 431 290
rect 467 262 495 290
rect 531 262 559 290
rect 595 262 623 290
rect 19 176 47 204
rect 83 176 111 204
rect 147 176 175 204
rect 211 176 239 204
rect 275 176 303 204
rect 339 176 367 204
rect 403 176 431 204
rect 467 176 495 204
rect 531 176 559 204
rect 595 176 623 204
rect 661 262 689 290
rect 725 262 753 290
rect 789 262 817 290
rect 853 262 881 290
rect 917 262 945 290
rect 981 262 1009 290
rect 1045 262 1073 290
rect 1109 262 1137 290
rect 1173 262 1201 290
rect 1237 262 1265 290
rect 661 176 689 204
rect 725 176 753 204
rect 789 176 817 204
rect 853 176 881 204
rect 917 176 945 204
rect 981 176 1009 204
rect 1045 176 1073 204
rect 1109 176 1137 204
rect 1173 176 1201 204
rect 1237 176 1265 204
rect 1303 262 1331 290
rect 1367 262 1395 290
rect 1431 262 1459 290
rect 1495 262 1523 290
rect 1559 262 1587 290
rect 1623 262 1651 290
rect 1687 262 1715 290
rect 1751 262 1779 290
rect 1815 262 1843 290
rect 1879 262 1907 290
rect 1303 176 1331 204
rect 1367 176 1395 204
rect 1431 176 1459 204
rect 1495 176 1523 204
rect 1559 176 1587 204
rect 1623 176 1651 204
rect 1687 176 1715 204
rect 1751 176 1779 204
rect 1815 176 1843 204
rect 1879 176 1907 204
rect 1945 262 1973 290
rect 2009 262 2037 290
rect 2073 262 2101 290
rect 2137 262 2165 290
rect 2201 262 2229 290
rect 2265 262 2293 290
rect 2329 262 2357 290
rect 2393 262 2421 290
rect 2457 262 2485 290
rect 2521 262 2549 290
rect 1945 176 1973 204
rect 2009 176 2037 204
rect 2073 176 2101 204
rect 2137 176 2165 204
rect 2201 176 2229 204
rect 2265 176 2293 204
rect 2329 176 2357 204
rect 2393 176 2421 204
rect 2457 176 2485 204
rect 2521 176 2549 204
rect 2587 262 2615 290
rect 2651 262 2679 290
rect 2715 262 2743 290
rect 2779 262 2807 290
rect 2843 262 2871 290
rect 2907 262 2935 290
rect 2971 262 2999 290
rect 3035 262 3063 290
rect 3099 262 3127 290
rect 3163 262 3191 290
rect 2587 176 2615 204
rect 2651 176 2679 204
rect 2715 176 2743 204
rect 2779 176 2807 204
rect 2843 176 2871 204
rect 2907 176 2935 204
rect 2971 176 2999 204
rect 3035 176 3063 204
rect 3099 176 3127 204
rect 3163 176 3191 204
rect 3229 262 3257 290
rect 3293 262 3321 290
rect 3357 262 3385 290
rect 3421 262 3449 290
rect 3485 262 3513 290
rect 3549 262 3577 290
rect 3613 262 3641 290
rect 3677 262 3705 290
rect 3741 262 3769 290
rect 3805 262 3833 290
rect 3229 176 3257 204
rect 3293 176 3321 204
rect 3357 176 3385 204
rect 3421 176 3449 204
rect 3485 176 3513 204
rect 3549 176 3577 204
rect 3613 176 3641 204
rect 3677 176 3705 204
rect 3741 176 3769 204
rect 3805 176 3833 204
rect 3871 262 3899 290
rect 3935 262 3963 290
rect 3999 262 4027 290
rect 4063 262 4091 290
rect 4127 262 4155 290
rect 4191 262 4219 290
rect 4255 262 4283 290
rect 4319 262 4347 290
rect 4383 262 4411 290
rect 4447 262 4475 290
rect 3871 176 3899 204
rect 3935 176 3963 204
rect 3999 176 4027 204
rect 4063 176 4091 204
rect 4127 176 4155 204
rect 4191 176 4219 204
rect 4255 176 4283 204
rect 4319 176 4347 204
rect 4383 176 4411 204
rect 4447 176 4475 204
rect 19 90 47 118
rect 83 90 111 118
rect 147 90 175 118
rect 211 90 239 118
rect 275 90 303 118
rect 339 90 367 118
rect 403 90 431 118
rect 467 90 495 118
rect 531 90 559 118
rect 595 90 623 118
rect 661 90 689 118
rect 725 90 753 118
rect 789 90 817 118
rect 853 90 881 118
rect 917 90 945 118
rect 981 90 1009 118
rect 1045 90 1073 118
rect 1109 90 1137 118
rect 1173 90 1201 118
rect 1237 90 1265 118
rect 1303 90 1331 118
rect 1367 90 1395 118
rect 1431 90 1459 118
rect 1495 90 1523 118
rect 1559 90 1587 118
rect 1623 90 1651 118
rect 1687 90 1715 118
rect 1751 90 1779 118
rect 1815 90 1843 118
rect 1879 90 1907 118
rect 1945 90 1973 118
rect 2009 90 2037 118
rect 2073 90 2101 118
rect 2137 90 2165 118
rect 2201 90 2229 118
rect 2265 90 2293 118
rect 2329 90 2357 118
rect 2393 90 2421 118
rect 2457 90 2485 118
rect 2521 90 2549 118
rect 2587 90 2615 118
rect 2651 90 2679 118
rect 2715 90 2743 118
rect 2779 90 2807 118
rect 2843 90 2871 118
rect 2907 90 2935 118
rect 2971 90 2999 118
rect 3035 90 3063 118
rect 3099 90 3127 118
rect 3163 90 3191 118
rect 3229 90 3257 118
rect 3293 90 3321 118
rect 3357 90 3385 118
rect 3421 90 3449 118
rect 3485 90 3513 118
rect 3549 90 3577 118
rect 3613 90 3641 118
rect 3677 90 3705 118
rect 3741 90 3769 118
rect 3805 90 3833 118
rect 3871 90 3899 118
rect 3935 90 3963 118
rect 3999 90 4027 118
rect 4063 90 4091 118
rect 4127 90 4155 118
rect 4191 90 4219 118
rect 4255 90 4283 118
rect 4319 90 4347 118
rect 4383 90 4411 118
rect 4447 90 4475 118
rect 4513 262 4541 290
rect 4577 262 4605 290
rect 4641 262 4669 290
rect 4705 262 4733 290
rect 4769 262 4797 290
rect 4833 262 4861 290
rect 4897 262 4925 290
rect 4961 262 4989 290
rect 5025 262 5053 290
rect 5089 262 5117 290
rect 4513 176 4541 204
rect 4577 176 4605 204
rect 4641 176 4669 204
rect 4705 176 4733 204
rect 4769 176 4797 204
rect 4833 176 4861 204
rect 4897 176 4925 204
rect 4961 176 4989 204
rect 5025 176 5053 204
rect 5089 176 5117 204
rect 4513 90 4541 118
rect 4577 90 4605 118
rect 4641 90 4669 118
rect 4705 90 4733 118
rect 4769 90 4797 118
rect 4833 90 4861 118
rect 4897 90 4925 118
rect 4961 90 4989 118
rect 5025 90 5053 118
rect 5089 90 5117 118
rect 5155 262 5183 290
rect 5219 262 5247 290
rect 5283 262 5311 290
rect 5347 262 5375 290
rect 5411 262 5439 290
rect 5475 262 5503 290
rect 5539 262 5567 290
rect 5603 262 5631 290
rect 5667 262 5695 290
rect 5731 262 5759 290
rect 5155 176 5183 204
rect 5219 176 5247 204
rect 5283 176 5311 204
rect 5347 176 5375 204
rect 5411 176 5439 204
rect 5475 176 5503 204
rect 5539 176 5567 204
rect 5603 176 5631 204
rect 5667 176 5695 204
rect 5731 176 5759 204
rect 5797 262 5825 290
rect 5861 262 5889 290
rect 5925 262 5953 290
rect 5989 262 6017 290
rect 6053 262 6081 290
rect 6117 262 6145 290
rect 6181 262 6209 290
rect 6245 262 6273 290
rect 6309 262 6337 290
rect 6373 262 6401 290
rect 5797 176 5825 204
rect 5861 176 5889 204
rect 5925 176 5953 204
rect 5989 176 6017 204
rect 6053 176 6081 204
rect 6117 176 6145 204
rect 6181 176 6209 204
rect 6245 176 6273 204
rect 6309 176 6337 204
rect 6373 176 6401 204
rect 6439 262 6467 290
rect 6503 262 6531 290
rect 6567 262 6595 290
rect 6631 262 6659 290
rect 6695 262 6723 290
rect 6759 262 6787 290
rect 6823 262 6851 290
rect 6887 262 6915 290
rect 6951 262 6979 290
rect 7015 262 7043 290
rect 6439 176 6467 204
rect 6503 176 6531 204
rect 6567 176 6595 204
rect 6631 176 6659 204
rect 6695 176 6723 204
rect 6759 176 6787 204
rect 6823 176 6851 204
rect 6887 176 6915 204
rect 6951 176 6979 204
rect 7015 176 7043 204
rect 7081 262 7109 290
rect 7145 262 7173 290
rect 7209 262 7237 290
rect 7273 262 7301 290
rect 7337 262 7365 290
rect 7401 262 7429 290
rect 7465 262 7493 290
rect 7529 262 7557 290
rect 7593 262 7621 290
rect 7657 262 7685 290
rect 7081 176 7109 204
rect 7145 176 7173 204
rect 7209 176 7237 204
rect 7273 176 7301 204
rect 7337 176 7365 204
rect 7401 176 7429 204
rect 7465 176 7493 204
rect 7529 176 7557 204
rect 7593 176 7621 204
rect 7657 176 7685 204
rect 5155 90 5183 118
rect 5219 90 5247 118
rect 5283 90 5311 118
rect 5347 90 5375 118
rect 5411 90 5439 118
rect 5475 90 5503 118
rect 5539 90 5567 118
rect 5603 90 5631 118
rect 5667 90 5695 118
rect 5731 90 5759 118
rect 5797 90 5825 118
rect 5861 90 5889 118
rect 5925 90 5953 118
rect 5989 90 6017 118
rect 6053 90 6081 118
rect 6117 90 6145 118
rect 6181 90 6209 118
rect 6245 90 6273 118
rect 6309 90 6337 118
rect 6373 90 6401 118
rect 6439 90 6467 118
rect 6503 90 6531 118
rect 6567 90 6595 118
rect 6631 90 6659 118
rect 6695 90 6723 118
rect 6759 90 6787 118
rect 6823 90 6851 118
rect 6887 90 6915 118
rect 6951 90 6979 118
rect 7015 90 7043 118
rect 7081 90 7109 118
rect 7145 90 7173 118
rect 7209 90 7237 118
rect 7273 90 7301 118
rect 7337 90 7365 118
rect 7401 90 7429 118
rect 7465 90 7493 118
rect 7529 90 7557 118
rect 7593 90 7621 118
rect 7657 90 7685 118
rect 7723 262 7751 290
rect 7787 262 7815 290
rect 7851 262 7879 290
rect 7915 262 7943 290
rect 7979 262 8007 290
rect 8043 262 8071 290
rect 8107 262 8135 290
rect 8171 262 8199 290
rect 8235 262 8263 290
rect 8299 262 8327 290
rect 7723 176 7751 204
rect 7787 176 7815 204
rect 7851 176 7879 204
rect 7915 176 7943 204
rect 7979 176 8007 204
rect 8043 176 8071 204
rect 8107 176 8135 204
rect 8171 176 8199 204
rect 8235 176 8263 204
rect 8299 176 8327 204
rect 7723 90 7751 118
rect 7787 90 7815 118
rect 7851 90 7879 118
rect 7915 90 7943 118
rect 7979 90 8007 118
rect 8043 90 8071 118
rect 8107 90 8135 118
rect 8171 90 8199 118
rect 8235 90 8263 118
rect 8299 90 8327 118
rect 8365 262 8393 290
rect 8429 262 8457 290
rect 8493 262 8521 290
rect 8557 262 8585 290
rect 8621 262 8649 290
rect 8685 262 8713 290
rect 8749 262 8777 290
rect 8813 262 8841 290
rect 8877 262 8905 290
rect 8941 262 8969 290
rect 8365 176 8393 204
rect 8429 176 8457 204
rect 8493 176 8521 204
rect 8557 176 8585 204
rect 8621 176 8649 204
rect 8685 176 8713 204
rect 8749 176 8777 204
rect 8813 176 8841 204
rect 8877 176 8905 204
rect 8941 176 8969 204
rect 9007 262 9035 290
rect 9071 262 9099 290
rect 9135 262 9163 290
rect 9199 262 9227 290
rect 9263 262 9291 290
rect 9327 262 9355 290
rect 9391 262 9419 290
rect 9455 262 9483 290
rect 9519 262 9547 290
rect 9583 262 9611 290
rect 8365 90 8393 118
rect 8429 90 8457 118
rect 8493 90 8521 118
rect 8557 90 8585 118
rect 8621 90 8649 118
rect 8685 90 8713 118
rect 8749 90 8777 118
rect 8813 90 8841 118
rect 8877 90 8905 118
rect 8941 90 8969 118
rect 9007 176 9035 204
rect 9071 176 9099 204
rect 9135 176 9163 204
rect 9199 176 9227 204
rect 9263 176 9291 204
rect 9327 176 9355 204
rect 9391 176 9419 204
rect 9455 176 9483 204
rect 9519 176 9547 204
rect 9583 176 9611 204
rect 9649 262 9677 290
rect 9713 262 9741 290
rect 9777 262 9805 290
rect 9841 262 9869 290
rect 9905 262 9933 290
rect 9969 262 9997 290
rect 10033 262 10061 290
rect 10097 262 10125 290
rect 10161 262 10189 290
rect 10225 262 10253 290
rect 9007 90 9035 118
rect 9071 90 9099 118
rect 9135 90 9163 118
rect 9199 90 9227 118
rect 9263 90 9291 118
rect 9327 90 9355 118
rect 9391 90 9419 118
rect 9455 90 9483 118
rect 9519 90 9547 118
rect 9583 90 9611 118
rect 9649 176 9677 204
rect 9713 176 9741 204
rect 9777 176 9805 204
rect 9841 176 9869 204
rect 9905 176 9933 204
rect 9969 176 9997 204
rect 10033 176 10061 204
rect 10097 176 10125 204
rect 10161 176 10189 204
rect 10225 176 10253 204
rect 10291 262 10319 290
rect 10355 262 10383 290
rect 10419 262 10447 290
rect 10483 262 10511 290
rect 10547 262 10575 290
rect 10611 262 10639 290
rect 10675 262 10703 290
rect 10739 262 10767 290
rect 10803 262 10831 290
rect 10867 262 10895 290
rect 9649 90 9677 118
rect 9713 90 9741 118
rect 9777 90 9805 118
rect 9841 90 9869 118
rect 9905 90 9933 118
rect 9969 90 9997 118
rect 10033 90 10061 118
rect 10097 90 10125 118
rect 10161 90 10189 118
rect 10225 90 10253 118
rect 10291 176 10319 204
rect 10355 176 10383 204
rect 10419 176 10447 204
rect 10483 176 10511 204
rect 10547 176 10575 204
rect 10611 176 10639 204
rect 10675 176 10703 204
rect 10739 176 10767 204
rect 10803 176 10831 204
rect 10867 176 10895 204
rect 10291 90 10319 118
rect 10355 90 10383 118
rect 10419 90 10447 118
rect 10483 90 10511 118
rect 10547 90 10575 118
rect 10611 90 10639 118
rect 10675 90 10703 118
rect 10739 90 10767 118
rect 10803 90 10831 118
rect 10867 90 10895 118
rect 10933 262 10961 290
rect 10997 262 11025 290
rect 11061 262 11089 290
rect 11125 262 11153 290
rect 11189 262 11217 290
rect 11253 262 11281 290
rect 11317 262 11345 290
rect 11381 262 11409 290
rect 11445 262 11473 290
rect 11509 262 11537 290
rect 10933 176 10961 204
rect 10997 176 11025 204
rect 11061 176 11089 204
rect 11125 176 11153 204
rect 11189 176 11217 204
rect 11253 176 11281 204
rect 11317 176 11345 204
rect 11381 176 11409 204
rect 11445 176 11473 204
rect 11509 176 11537 204
rect 10933 90 10961 118
rect 10997 90 11025 118
rect 11061 90 11089 118
rect 11125 90 11153 118
rect 11189 90 11217 118
rect 11253 90 11281 118
rect 11317 90 11345 118
rect 11381 90 11409 118
rect 11445 90 11473 118
rect 11509 90 11537 118
rect 11575 262 11603 290
rect 11639 262 11667 290
rect 11703 262 11731 290
rect 11767 262 11795 290
rect 11831 262 11859 290
rect 11895 262 11923 290
rect 11959 262 11987 290
rect 12023 262 12051 290
rect 12087 262 12115 290
rect 12151 262 12179 290
rect 11575 176 11603 204
rect 11639 176 11667 204
rect 11703 176 11731 204
rect 11767 176 11795 204
rect 11831 176 11859 204
rect 11895 176 11923 204
rect 11959 176 11987 204
rect 12023 176 12051 204
rect 12087 176 12115 204
rect 12151 176 12179 204
rect 12217 262 12245 290
rect 12281 262 12309 290
rect 12345 262 12373 290
rect 12409 262 12437 290
rect 12473 262 12501 290
rect 12537 262 12565 290
rect 12601 262 12629 290
rect 12665 262 12693 290
rect 12729 262 12757 290
rect 12793 262 12821 290
rect 12217 176 12245 204
rect 12281 176 12309 204
rect 12345 176 12373 204
rect 12409 176 12437 204
rect 12473 176 12501 204
rect 12537 176 12565 204
rect 12601 176 12629 204
rect 12665 176 12693 204
rect 12729 176 12757 204
rect 12793 176 12821 204
rect 11575 90 11603 118
rect 11639 90 11667 118
rect 11703 90 11731 118
rect 11767 90 11795 118
rect 11831 90 11859 118
rect 11895 90 11923 118
rect 11959 90 11987 118
rect 12023 90 12051 118
rect 12087 90 12115 118
rect 12151 90 12179 118
rect 12217 90 12245 118
rect 12281 90 12309 118
rect 12345 90 12373 118
rect 12409 90 12437 118
rect 12473 90 12501 118
rect 12537 90 12565 118
rect 12601 90 12629 118
rect 12665 90 12693 118
rect 12729 90 12757 118
rect 12793 90 12821 118
<< metal3 >>
rect 16 1430 50 1469
rect 16 1402 19 1430
rect 47 1402 50 1430
rect 16 1344 50 1402
rect 16 1316 19 1344
rect 47 1316 50 1344
rect 16 1258 50 1316
rect 16 1230 19 1258
rect 47 1230 50 1258
rect 16 1191 50 1230
rect 80 1430 114 1469
rect 80 1402 83 1430
rect 111 1402 114 1430
rect 80 1344 114 1402
rect 80 1316 83 1344
rect 111 1316 114 1344
rect 80 1258 114 1316
rect 80 1230 83 1258
rect 111 1230 114 1258
rect 80 1191 114 1230
rect 144 1430 178 1469
rect 144 1402 147 1430
rect 175 1402 178 1430
rect 144 1344 178 1402
rect 144 1316 147 1344
rect 175 1316 178 1344
rect 144 1258 178 1316
rect 144 1230 147 1258
rect 175 1230 178 1258
rect 144 1191 178 1230
rect 208 1430 242 1469
rect 208 1402 211 1430
rect 239 1402 242 1430
rect 208 1344 242 1402
rect 208 1316 211 1344
rect 239 1316 242 1344
rect 208 1258 242 1316
rect 208 1230 211 1258
rect 239 1230 242 1258
rect 208 1191 242 1230
rect 272 1430 306 1469
rect 272 1402 275 1430
rect 303 1402 306 1430
rect 272 1344 306 1402
rect 272 1316 275 1344
rect 303 1316 306 1344
rect 272 1258 306 1316
rect 272 1230 275 1258
rect 303 1230 306 1258
rect 272 1191 306 1230
rect 336 1430 370 1469
rect 336 1402 339 1430
rect 367 1402 370 1430
rect 336 1344 370 1402
rect 336 1316 339 1344
rect 367 1316 370 1344
rect 336 1258 370 1316
rect 336 1230 339 1258
rect 367 1230 370 1258
rect 336 1191 370 1230
rect 400 1430 434 1469
rect 400 1402 403 1430
rect 431 1402 434 1430
rect 400 1344 434 1402
rect 400 1316 403 1344
rect 431 1316 434 1344
rect 400 1258 434 1316
rect 400 1230 403 1258
rect 431 1230 434 1258
rect 400 1191 434 1230
rect 464 1430 498 1469
rect 464 1402 467 1430
rect 495 1402 498 1430
rect 464 1344 498 1402
rect 464 1316 467 1344
rect 495 1316 498 1344
rect 464 1258 498 1316
rect 464 1230 467 1258
rect 495 1230 498 1258
rect 464 1191 498 1230
rect 528 1430 562 1469
rect 528 1402 531 1430
rect 559 1402 562 1430
rect 528 1344 562 1402
rect 528 1316 531 1344
rect 559 1316 562 1344
rect 528 1258 562 1316
rect 528 1230 531 1258
rect 559 1230 562 1258
rect 528 1191 562 1230
rect 592 1430 626 1469
rect 592 1402 595 1430
rect 623 1402 626 1430
rect 592 1344 626 1402
rect 592 1316 595 1344
rect 623 1316 626 1344
rect 592 1258 626 1316
rect 592 1230 595 1258
rect 623 1230 626 1258
rect 592 1191 626 1230
rect 658 1430 692 1469
rect 658 1402 661 1430
rect 689 1402 692 1430
rect 658 1344 692 1402
rect 658 1316 661 1344
rect 689 1316 692 1344
rect 658 1258 692 1316
rect 658 1230 661 1258
rect 689 1230 692 1258
rect 658 1191 692 1230
rect 722 1430 756 1469
rect 722 1402 725 1430
rect 753 1402 756 1430
rect 722 1344 756 1402
rect 722 1316 725 1344
rect 753 1316 756 1344
rect 722 1258 756 1316
rect 722 1230 725 1258
rect 753 1230 756 1258
rect 722 1191 756 1230
rect 786 1430 820 1469
rect 786 1402 789 1430
rect 817 1402 820 1430
rect 786 1344 820 1402
rect 786 1316 789 1344
rect 817 1316 820 1344
rect 786 1258 820 1316
rect 786 1230 789 1258
rect 817 1230 820 1258
rect 786 1191 820 1230
rect 850 1430 884 1469
rect 850 1402 853 1430
rect 881 1402 884 1430
rect 850 1344 884 1402
rect 850 1316 853 1344
rect 881 1316 884 1344
rect 850 1258 884 1316
rect 850 1230 853 1258
rect 881 1230 884 1258
rect 850 1191 884 1230
rect 914 1430 948 1469
rect 914 1402 917 1430
rect 945 1402 948 1430
rect 914 1344 948 1402
rect 914 1316 917 1344
rect 945 1316 948 1344
rect 914 1258 948 1316
rect 914 1230 917 1258
rect 945 1230 948 1258
rect 914 1191 948 1230
rect 978 1430 1012 1469
rect 978 1402 981 1430
rect 1009 1402 1012 1430
rect 978 1344 1012 1402
rect 978 1316 981 1344
rect 1009 1316 1012 1344
rect 978 1258 1012 1316
rect 978 1230 981 1258
rect 1009 1230 1012 1258
rect 978 1191 1012 1230
rect 1042 1430 1076 1469
rect 1042 1402 1045 1430
rect 1073 1402 1076 1430
rect 1042 1344 1076 1402
rect 1042 1316 1045 1344
rect 1073 1316 1076 1344
rect 1042 1258 1076 1316
rect 1042 1230 1045 1258
rect 1073 1230 1076 1258
rect 1042 1191 1076 1230
rect 1106 1430 1140 1469
rect 1106 1402 1109 1430
rect 1137 1402 1140 1430
rect 1106 1344 1140 1402
rect 1106 1316 1109 1344
rect 1137 1316 1140 1344
rect 1106 1258 1140 1316
rect 1106 1230 1109 1258
rect 1137 1230 1140 1258
rect 1106 1191 1140 1230
rect 1170 1430 1204 1469
rect 1170 1402 1173 1430
rect 1201 1402 1204 1430
rect 1170 1344 1204 1402
rect 1170 1316 1173 1344
rect 1201 1316 1204 1344
rect 1170 1258 1204 1316
rect 1170 1230 1173 1258
rect 1201 1230 1204 1258
rect 1170 1191 1204 1230
rect 1234 1430 1268 1469
rect 1234 1402 1237 1430
rect 1265 1402 1268 1430
rect 1234 1344 1268 1402
rect 1234 1316 1237 1344
rect 1265 1316 1268 1344
rect 1234 1258 1268 1316
rect 1234 1230 1237 1258
rect 1265 1230 1268 1258
rect 1234 1191 1268 1230
rect 1300 1430 1334 1469
rect 1300 1402 1303 1430
rect 1331 1402 1334 1430
rect 1300 1344 1334 1402
rect 1300 1316 1303 1344
rect 1331 1316 1334 1344
rect 1300 1258 1334 1316
rect 1300 1230 1303 1258
rect 1331 1230 1334 1258
rect 1300 1191 1334 1230
rect 1364 1430 1398 1469
rect 1364 1402 1367 1430
rect 1395 1402 1398 1430
rect 1364 1344 1398 1402
rect 1364 1316 1367 1344
rect 1395 1316 1398 1344
rect 1364 1258 1398 1316
rect 1364 1230 1367 1258
rect 1395 1230 1398 1258
rect 1364 1191 1398 1230
rect 1428 1430 1462 1469
rect 1428 1402 1431 1430
rect 1459 1402 1462 1430
rect 1428 1344 1462 1402
rect 1428 1316 1431 1344
rect 1459 1316 1462 1344
rect 1428 1258 1462 1316
rect 1428 1230 1431 1258
rect 1459 1230 1462 1258
rect 1428 1191 1462 1230
rect 1492 1430 1526 1469
rect 1492 1402 1495 1430
rect 1523 1402 1526 1430
rect 1492 1344 1526 1402
rect 1492 1316 1495 1344
rect 1523 1316 1526 1344
rect 1492 1258 1526 1316
rect 1492 1230 1495 1258
rect 1523 1230 1526 1258
rect 1492 1191 1526 1230
rect 1556 1430 1590 1469
rect 1556 1402 1559 1430
rect 1587 1402 1590 1430
rect 1556 1344 1590 1402
rect 1556 1316 1559 1344
rect 1587 1316 1590 1344
rect 1556 1258 1590 1316
rect 1556 1230 1559 1258
rect 1587 1230 1590 1258
rect 1556 1191 1590 1230
rect 1620 1430 1654 1469
rect 1620 1402 1623 1430
rect 1651 1402 1654 1430
rect 1620 1344 1654 1402
rect 1620 1316 1623 1344
rect 1651 1316 1654 1344
rect 1620 1258 1654 1316
rect 1620 1230 1623 1258
rect 1651 1230 1654 1258
rect 1620 1191 1654 1230
rect 1684 1430 1718 1469
rect 1684 1402 1687 1430
rect 1715 1402 1718 1430
rect 1684 1344 1718 1402
rect 1684 1316 1687 1344
rect 1715 1316 1718 1344
rect 1684 1258 1718 1316
rect 1684 1230 1687 1258
rect 1715 1230 1718 1258
rect 1684 1191 1718 1230
rect 1748 1430 1782 1469
rect 1748 1402 1751 1430
rect 1779 1402 1782 1430
rect 1748 1344 1782 1402
rect 1748 1316 1751 1344
rect 1779 1316 1782 1344
rect 1748 1258 1782 1316
rect 1748 1230 1751 1258
rect 1779 1230 1782 1258
rect 1748 1191 1782 1230
rect 1812 1430 1846 1469
rect 1812 1402 1815 1430
rect 1843 1402 1846 1430
rect 1812 1344 1846 1402
rect 1812 1316 1815 1344
rect 1843 1316 1846 1344
rect 1812 1258 1846 1316
rect 1812 1230 1815 1258
rect 1843 1230 1846 1258
rect 1812 1191 1846 1230
rect 1876 1430 1910 1469
rect 1876 1402 1879 1430
rect 1907 1402 1910 1430
rect 1876 1344 1910 1402
rect 1876 1316 1879 1344
rect 1907 1316 1910 1344
rect 1876 1258 1910 1316
rect 1876 1230 1879 1258
rect 1907 1230 1910 1258
rect 1876 1191 1910 1230
rect 1942 1430 1976 1469
rect 1942 1402 1945 1430
rect 1973 1402 1976 1430
rect 1942 1344 1976 1402
rect 1942 1316 1945 1344
rect 1973 1316 1976 1344
rect 1942 1258 1976 1316
rect 1942 1230 1945 1258
rect 1973 1230 1976 1258
rect 1942 1191 1976 1230
rect 2006 1430 2040 1469
rect 2006 1402 2009 1430
rect 2037 1402 2040 1430
rect 2006 1344 2040 1402
rect 2006 1316 2009 1344
rect 2037 1316 2040 1344
rect 2006 1258 2040 1316
rect 2006 1230 2009 1258
rect 2037 1230 2040 1258
rect 2006 1191 2040 1230
rect 2070 1430 2104 1469
rect 2070 1402 2073 1430
rect 2101 1402 2104 1430
rect 2070 1344 2104 1402
rect 2070 1316 2073 1344
rect 2101 1316 2104 1344
rect 2070 1258 2104 1316
rect 2070 1230 2073 1258
rect 2101 1230 2104 1258
rect 2070 1191 2104 1230
rect 2134 1430 2168 1469
rect 2134 1402 2137 1430
rect 2165 1402 2168 1430
rect 2134 1344 2168 1402
rect 2134 1316 2137 1344
rect 2165 1316 2168 1344
rect 2134 1258 2168 1316
rect 2134 1230 2137 1258
rect 2165 1230 2168 1258
rect 2134 1191 2168 1230
rect 2198 1430 2232 1469
rect 2198 1402 2201 1430
rect 2229 1402 2232 1430
rect 2198 1344 2232 1402
rect 2198 1316 2201 1344
rect 2229 1316 2232 1344
rect 2198 1258 2232 1316
rect 2198 1230 2201 1258
rect 2229 1230 2232 1258
rect 2198 1191 2232 1230
rect 2262 1430 2296 1469
rect 2262 1402 2265 1430
rect 2293 1402 2296 1430
rect 2262 1344 2296 1402
rect 2262 1316 2265 1344
rect 2293 1316 2296 1344
rect 2262 1258 2296 1316
rect 2262 1230 2265 1258
rect 2293 1230 2296 1258
rect 2262 1191 2296 1230
rect 2326 1430 2360 1469
rect 2326 1402 2329 1430
rect 2357 1402 2360 1430
rect 2326 1344 2360 1402
rect 2326 1316 2329 1344
rect 2357 1316 2360 1344
rect 2326 1258 2360 1316
rect 2326 1230 2329 1258
rect 2357 1230 2360 1258
rect 2326 1191 2360 1230
rect 2390 1430 2424 1469
rect 2390 1402 2393 1430
rect 2421 1402 2424 1430
rect 2390 1344 2424 1402
rect 2390 1316 2393 1344
rect 2421 1316 2424 1344
rect 2390 1258 2424 1316
rect 2390 1230 2393 1258
rect 2421 1230 2424 1258
rect 2390 1191 2424 1230
rect 2454 1430 2488 1469
rect 2454 1402 2457 1430
rect 2485 1402 2488 1430
rect 2454 1344 2488 1402
rect 2454 1316 2457 1344
rect 2485 1316 2488 1344
rect 2454 1258 2488 1316
rect 2454 1230 2457 1258
rect 2485 1230 2488 1258
rect 2454 1191 2488 1230
rect 2518 1430 2552 1469
rect 2518 1402 2521 1430
rect 2549 1402 2552 1430
rect 2518 1344 2552 1402
rect 2518 1316 2521 1344
rect 2549 1316 2552 1344
rect 2518 1258 2552 1316
rect 2518 1230 2521 1258
rect 2549 1230 2552 1258
rect 2518 1191 2552 1230
rect 2584 1430 2618 1469
rect 2584 1402 2587 1430
rect 2615 1402 2618 1430
rect 2584 1344 2618 1402
rect 2584 1316 2587 1344
rect 2615 1316 2618 1344
rect 2584 1258 2618 1316
rect 2584 1230 2587 1258
rect 2615 1230 2618 1258
rect 2584 1191 2618 1230
rect 2648 1430 2682 1469
rect 2648 1402 2651 1430
rect 2679 1402 2682 1430
rect 2648 1344 2682 1402
rect 2648 1316 2651 1344
rect 2679 1316 2682 1344
rect 2648 1258 2682 1316
rect 2648 1230 2651 1258
rect 2679 1230 2682 1258
rect 2648 1191 2682 1230
rect 2712 1430 2746 1469
rect 2712 1402 2715 1430
rect 2743 1402 2746 1430
rect 2712 1344 2746 1402
rect 2712 1316 2715 1344
rect 2743 1316 2746 1344
rect 2712 1258 2746 1316
rect 2712 1230 2715 1258
rect 2743 1230 2746 1258
rect 2712 1191 2746 1230
rect 2776 1430 2810 1469
rect 2776 1402 2779 1430
rect 2807 1402 2810 1430
rect 2776 1344 2810 1402
rect 2776 1316 2779 1344
rect 2807 1316 2810 1344
rect 2776 1258 2810 1316
rect 2776 1230 2779 1258
rect 2807 1230 2810 1258
rect 2776 1191 2810 1230
rect 2840 1430 2874 1469
rect 2840 1402 2843 1430
rect 2871 1402 2874 1430
rect 2840 1344 2874 1402
rect 2840 1316 2843 1344
rect 2871 1316 2874 1344
rect 2840 1258 2874 1316
rect 2840 1230 2843 1258
rect 2871 1230 2874 1258
rect 2840 1191 2874 1230
rect 2904 1430 2938 1469
rect 2904 1402 2907 1430
rect 2935 1402 2938 1430
rect 2904 1344 2938 1402
rect 2904 1316 2907 1344
rect 2935 1316 2938 1344
rect 2904 1258 2938 1316
rect 2904 1230 2907 1258
rect 2935 1230 2938 1258
rect 2904 1191 2938 1230
rect 2968 1430 3002 1469
rect 2968 1402 2971 1430
rect 2999 1402 3002 1430
rect 2968 1344 3002 1402
rect 2968 1316 2971 1344
rect 2999 1316 3002 1344
rect 2968 1258 3002 1316
rect 2968 1230 2971 1258
rect 2999 1230 3002 1258
rect 2968 1191 3002 1230
rect 3032 1430 3066 1469
rect 3032 1402 3035 1430
rect 3063 1402 3066 1430
rect 3032 1344 3066 1402
rect 3032 1316 3035 1344
rect 3063 1316 3066 1344
rect 3032 1258 3066 1316
rect 3032 1230 3035 1258
rect 3063 1230 3066 1258
rect 3032 1191 3066 1230
rect 3096 1430 3130 1469
rect 3096 1402 3099 1430
rect 3127 1402 3130 1430
rect 3096 1344 3130 1402
rect 3096 1316 3099 1344
rect 3127 1316 3130 1344
rect 3096 1258 3130 1316
rect 3096 1230 3099 1258
rect 3127 1230 3130 1258
rect 3096 1191 3130 1230
rect 3160 1430 3194 1469
rect 3160 1402 3163 1430
rect 3191 1402 3194 1430
rect 3160 1344 3194 1402
rect 3160 1316 3163 1344
rect 3191 1316 3194 1344
rect 3160 1258 3194 1316
rect 3160 1230 3163 1258
rect 3191 1230 3194 1258
rect 3160 1191 3194 1230
rect 3226 1430 3260 1469
rect 3226 1402 3229 1430
rect 3257 1402 3260 1430
rect 3226 1344 3260 1402
rect 3226 1316 3229 1344
rect 3257 1316 3260 1344
rect 3226 1258 3260 1316
rect 3226 1230 3229 1258
rect 3257 1230 3260 1258
rect 3226 1191 3260 1230
rect 3290 1430 3324 1469
rect 3290 1402 3293 1430
rect 3321 1402 3324 1430
rect 3290 1344 3324 1402
rect 3290 1316 3293 1344
rect 3321 1316 3324 1344
rect 3290 1258 3324 1316
rect 3290 1230 3293 1258
rect 3321 1230 3324 1258
rect 3290 1191 3324 1230
rect 3354 1430 3388 1469
rect 3354 1402 3357 1430
rect 3385 1402 3388 1430
rect 3354 1344 3388 1402
rect 3354 1316 3357 1344
rect 3385 1316 3388 1344
rect 3354 1258 3388 1316
rect 3354 1230 3357 1258
rect 3385 1230 3388 1258
rect 3354 1191 3388 1230
rect 3418 1430 3452 1469
rect 3418 1402 3421 1430
rect 3449 1402 3452 1430
rect 3418 1344 3452 1402
rect 3418 1316 3421 1344
rect 3449 1316 3452 1344
rect 3418 1258 3452 1316
rect 3418 1230 3421 1258
rect 3449 1230 3452 1258
rect 3418 1191 3452 1230
rect 3482 1430 3516 1469
rect 3482 1402 3485 1430
rect 3513 1402 3516 1430
rect 3482 1344 3516 1402
rect 3482 1316 3485 1344
rect 3513 1316 3516 1344
rect 3482 1258 3516 1316
rect 3482 1230 3485 1258
rect 3513 1230 3516 1258
rect 3482 1191 3516 1230
rect 3546 1430 3580 1469
rect 3546 1402 3549 1430
rect 3577 1402 3580 1430
rect 3546 1344 3580 1402
rect 3546 1316 3549 1344
rect 3577 1316 3580 1344
rect 3546 1258 3580 1316
rect 3546 1230 3549 1258
rect 3577 1230 3580 1258
rect 3546 1191 3580 1230
rect 3610 1430 3644 1469
rect 3610 1402 3613 1430
rect 3641 1402 3644 1430
rect 3610 1344 3644 1402
rect 3610 1316 3613 1344
rect 3641 1316 3644 1344
rect 3610 1258 3644 1316
rect 3610 1230 3613 1258
rect 3641 1230 3644 1258
rect 3610 1191 3644 1230
rect 3674 1430 3708 1469
rect 3674 1402 3677 1430
rect 3705 1402 3708 1430
rect 3674 1344 3708 1402
rect 3674 1316 3677 1344
rect 3705 1316 3708 1344
rect 3674 1258 3708 1316
rect 3674 1230 3677 1258
rect 3705 1230 3708 1258
rect 3674 1191 3708 1230
rect 3738 1430 3772 1469
rect 3738 1402 3741 1430
rect 3769 1402 3772 1430
rect 3738 1344 3772 1402
rect 3738 1316 3741 1344
rect 3769 1316 3772 1344
rect 3738 1258 3772 1316
rect 3738 1230 3741 1258
rect 3769 1230 3772 1258
rect 3738 1191 3772 1230
rect 3802 1430 3836 1469
rect 3802 1402 3805 1430
rect 3833 1402 3836 1430
rect 3802 1344 3836 1402
rect 3802 1316 3805 1344
rect 3833 1316 3836 1344
rect 3802 1258 3836 1316
rect 3802 1230 3805 1258
rect 3833 1230 3836 1258
rect 3802 1191 3836 1230
rect 3868 1430 3902 1469
rect 3868 1402 3871 1430
rect 3899 1402 3902 1430
rect 3868 1344 3902 1402
rect 3868 1316 3871 1344
rect 3899 1316 3902 1344
rect 3868 1258 3902 1316
rect 3868 1230 3871 1258
rect 3899 1230 3902 1258
rect 3868 1191 3902 1230
rect 3932 1430 3966 1469
rect 3932 1402 3935 1430
rect 3963 1402 3966 1430
rect 3932 1344 3966 1402
rect 3932 1316 3935 1344
rect 3963 1316 3966 1344
rect 3932 1258 3966 1316
rect 3932 1230 3935 1258
rect 3963 1230 3966 1258
rect 3932 1191 3966 1230
rect 3996 1430 4030 1469
rect 3996 1402 3999 1430
rect 4027 1402 4030 1430
rect 3996 1344 4030 1402
rect 3996 1316 3999 1344
rect 4027 1316 4030 1344
rect 3996 1258 4030 1316
rect 3996 1230 3999 1258
rect 4027 1230 4030 1258
rect 3996 1191 4030 1230
rect 4060 1430 4094 1469
rect 4060 1402 4063 1430
rect 4091 1402 4094 1430
rect 4060 1344 4094 1402
rect 4060 1316 4063 1344
rect 4091 1316 4094 1344
rect 4060 1258 4094 1316
rect 4060 1230 4063 1258
rect 4091 1230 4094 1258
rect 4060 1191 4094 1230
rect 4124 1430 4158 1469
rect 4124 1402 4127 1430
rect 4155 1402 4158 1430
rect 4124 1344 4158 1402
rect 4124 1316 4127 1344
rect 4155 1316 4158 1344
rect 4124 1258 4158 1316
rect 4124 1230 4127 1258
rect 4155 1230 4158 1258
rect 4124 1191 4158 1230
rect 4188 1430 4222 1469
rect 4188 1402 4191 1430
rect 4219 1402 4222 1430
rect 4188 1344 4222 1402
rect 4188 1316 4191 1344
rect 4219 1316 4222 1344
rect 4188 1258 4222 1316
rect 4188 1230 4191 1258
rect 4219 1230 4222 1258
rect 4188 1191 4222 1230
rect 4252 1430 4286 1469
rect 4252 1402 4255 1430
rect 4283 1402 4286 1430
rect 4252 1344 4286 1402
rect 4252 1316 4255 1344
rect 4283 1316 4286 1344
rect 4252 1258 4286 1316
rect 4252 1230 4255 1258
rect 4283 1230 4286 1258
rect 4252 1191 4286 1230
rect 4316 1430 4350 1469
rect 4316 1402 4319 1430
rect 4347 1402 4350 1430
rect 4316 1344 4350 1402
rect 4316 1316 4319 1344
rect 4347 1316 4350 1344
rect 4316 1258 4350 1316
rect 4316 1230 4319 1258
rect 4347 1230 4350 1258
rect 4316 1191 4350 1230
rect 4380 1430 4414 1469
rect 4380 1402 4383 1430
rect 4411 1402 4414 1430
rect 4380 1344 4414 1402
rect 4380 1316 4383 1344
rect 4411 1316 4414 1344
rect 4380 1258 4414 1316
rect 4380 1230 4383 1258
rect 4411 1230 4414 1258
rect 4380 1191 4414 1230
rect 4444 1430 4478 1469
rect 4444 1402 4447 1430
rect 4475 1402 4478 1430
rect 4444 1344 4478 1402
rect 4444 1316 4447 1344
rect 4475 1316 4478 1344
rect 4444 1258 4478 1316
rect 4444 1230 4447 1258
rect 4475 1230 4478 1258
rect 4444 1191 4478 1230
rect 4510 1430 4544 1469
rect 4510 1402 4513 1430
rect 4541 1402 4544 1430
rect 4510 1344 4544 1402
rect 4510 1316 4513 1344
rect 4541 1316 4544 1344
rect 4510 1258 4544 1316
rect 4510 1230 4513 1258
rect 4541 1230 4544 1258
rect 4510 1191 4544 1230
rect 4574 1430 4608 1469
rect 4574 1402 4577 1430
rect 4605 1402 4608 1430
rect 4574 1344 4608 1402
rect 4574 1316 4577 1344
rect 4605 1316 4608 1344
rect 4574 1258 4608 1316
rect 4574 1230 4577 1258
rect 4605 1230 4608 1258
rect 4574 1191 4608 1230
rect 4638 1430 4672 1469
rect 4638 1402 4641 1430
rect 4669 1402 4672 1430
rect 4638 1344 4672 1402
rect 4638 1316 4641 1344
rect 4669 1316 4672 1344
rect 4638 1258 4672 1316
rect 4638 1230 4641 1258
rect 4669 1230 4672 1258
rect 4638 1191 4672 1230
rect 4702 1430 4736 1469
rect 4702 1402 4705 1430
rect 4733 1402 4736 1430
rect 4702 1344 4736 1402
rect 4702 1316 4705 1344
rect 4733 1316 4736 1344
rect 4702 1258 4736 1316
rect 4702 1230 4705 1258
rect 4733 1230 4736 1258
rect 4702 1191 4736 1230
rect 4766 1430 4800 1469
rect 4766 1402 4769 1430
rect 4797 1402 4800 1430
rect 4766 1344 4800 1402
rect 4766 1316 4769 1344
rect 4797 1316 4800 1344
rect 4766 1258 4800 1316
rect 4766 1230 4769 1258
rect 4797 1230 4800 1258
rect 4766 1191 4800 1230
rect 4830 1430 4864 1469
rect 4830 1402 4833 1430
rect 4861 1402 4864 1430
rect 4830 1344 4864 1402
rect 4830 1316 4833 1344
rect 4861 1316 4864 1344
rect 4830 1258 4864 1316
rect 4830 1230 4833 1258
rect 4861 1230 4864 1258
rect 4830 1191 4864 1230
rect 4894 1430 4928 1469
rect 4894 1402 4897 1430
rect 4925 1402 4928 1430
rect 4894 1344 4928 1402
rect 4894 1316 4897 1344
rect 4925 1316 4928 1344
rect 4894 1258 4928 1316
rect 4894 1230 4897 1258
rect 4925 1230 4928 1258
rect 4894 1191 4928 1230
rect 4958 1430 4992 1469
rect 4958 1402 4961 1430
rect 4989 1402 4992 1430
rect 4958 1344 4992 1402
rect 4958 1316 4961 1344
rect 4989 1316 4992 1344
rect 4958 1258 4992 1316
rect 4958 1230 4961 1258
rect 4989 1230 4992 1258
rect 4958 1191 4992 1230
rect 5022 1430 5056 1469
rect 5022 1402 5025 1430
rect 5053 1402 5056 1430
rect 5022 1344 5056 1402
rect 5022 1316 5025 1344
rect 5053 1316 5056 1344
rect 5022 1258 5056 1316
rect 5022 1230 5025 1258
rect 5053 1230 5056 1258
rect 5022 1191 5056 1230
rect 5086 1430 5120 1469
rect 5086 1402 5089 1430
rect 5117 1402 5120 1430
rect 5086 1344 5120 1402
rect 5086 1316 5089 1344
rect 5117 1316 5120 1344
rect 5086 1258 5120 1316
rect 5086 1230 5089 1258
rect 5117 1230 5120 1258
rect 5086 1191 5120 1230
rect 5152 1430 5186 1469
rect 5152 1402 5155 1430
rect 5183 1402 5186 1430
rect 5152 1344 5186 1402
rect 5152 1316 5155 1344
rect 5183 1316 5186 1344
rect 5152 1258 5186 1316
rect 5152 1230 5155 1258
rect 5183 1230 5186 1258
rect 5152 1191 5186 1230
rect 5216 1430 5250 1469
rect 5216 1402 5219 1430
rect 5247 1402 5250 1430
rect 5216 1344 5250 1402
rect 5216 1316 5219 1344
rect 5247 1316 5250 1344
rect 5216 1258 5250 1316
rect 5216 1230 5219 1258
rect 5247 1230 5250 1258
rect 5216 1191 5250 1230
rect 5280 1430 5314 1469
rect 5280 1402 5283 1430
rect 5311 1402 5314 1430
rect 5280 1344 5314 1402
rect 5280 1316 5283 1344
rect 5311 1316 5314 1344
rect 5280 1258 5314 1316
rect 5280 1230 5283 1258
rect 5311 1230 5314 1258
rect 5280 1191 5314 1230
rect 5344 1430 5378 1469
rect 5344 1402 5347 1430
rect 5375 1402 5378 1430
rect 5344 1344 5378 1402
rect 5344 1316 5347 1344
rect 5375 1316 5378 1344
rect 5344 1258 5378 1316
rect 5344 1230 5347 1258
rect 5375 1230 5378 1258
rect 5344 1191 5378 1230
rect 5408 1430 5442 1469
rect 5408 1402 5411 1430
rect 5439 1402 5442 1430
rect 5408 1344 5442 1402
rect 5408 1316 5411 1344
rect 5439 1316 5442 1344
rect 5408 1258 5442 1316
rect 5408 1230 5411 1258
rect 5439 1230 5442 1258
rect 5408 1191 5442 1230
rect 5472 1430 5506 1469
rect 5472 1402 5475 1430
rect 5503 1402 5506 1430
rect 5472 1344 5506 1402
rect 5472 1316 5475 1344
rect 5503 1316 5506 1344
rect 5472 1258 5506 1316
rect 5472 1230 5475 1258
rect 5503 1230 5506 1258
rect 5472 1191 5506 1230
rect 5536 1430 5570 1469
rect 5536 1402 5539 1430
rect 5567 1402 5570 1430
rect 5536 1344 5570 1402
rect 5536 1316 5539 1344
rect 5567 1316 5570 1344
rect 5536 1258 5570 1316
rect 5536 1230 5539 1258
rect 5567 1230 5570 1258
rect 5536 1191 5570 1230
rect 5600 1430 5634 1469
rect 5600 1402 5603 1430
rect 5631 1402 5634 1430
rect 5600 1344 5634 1402
rect 5600 1316 5603 1344
rect 5631 1316 5634 1344
rect 5600 1258 5634 1316
rect 5600 1230 5603 1258
rect 5631 1230 5634 1258
rect 5600 1191 5634 1230
rect 5664 1430 5698 1469
rect 5664 1402 5667 1430
rect 5695 1402 5698 1430
rect 5664 1344 5698 1402
rect 5664 1316 5667 1344
rect 5695 1316 5698 1344
rect 5664 1258 5698 1316
rect 5664 1230 5667 1258
rect 5695 1230 5698 1258
rect 5664 1191 5698 1230
rect 5728 1430 5762 1469
rect 5728 1402 5731 1430
rect 5759 1402 5762 1430
rect 5728 1344 5762 1402
rect 5728 1316 5731 1344
rect 5759 1316 5762 1344
rect 5728 1258 5762 1316
rect 5728 1230 5731 1258
rect 5759 1230 5762 1258
rect 5728 1191 5762 1230
rect 5794 1430 5828 1469
rect 5794 1402 5797 1430
rect 5825 1402 5828 1430
rect 5794 1344 5828 1402
rect 5794 1316 5797 1344
rect 5825 1316 5828 1344
rect 5794 1258 5828 1316
rect 5794 1230 5797 1258
rect 5825 1230 5828 1258
rect 5794 1191 5828 1230
rect 5858 1430 5892 1469
rect 5858 1402 5861 1430
rect 5889 1402 5892 1430
rect 5858 1344 5892 1402
rect 5858 1316 5861 1344
rect 5889 1316 5892 1344
rect 5858 1258 5892 1316
rect 5858 1230 5861 1258
rect 5889 1230 5892 1258
rect 5858 1191 5892 1230
rect 5922 1430 5956 1469
rect 5922 1402 5925 1430
rect 5953 1402 5956 1430
rect 5922 1344 5956 1402
rect 5922 1316 5925 1344
rect 5953 1316 5956 1344
rect 5922 1258 5956 1316
rect 5922 1230 5925 1258
rect 5953 1230 5956 1258
rect 5922 1191 5956 1230
rect 5986 1430 6020 1469
rect 5986 1402 5989 1430
rect 6017 1402 6020 1430
rect 5986 1344 6020 1402
rect 5986 1316 5989 1344
rect 6017 1316 6020 1344
rect 5986 1258 6020 1316
rect 5986 1230 5989 1258
rect 6017 1230 6020 1258
rect 5986 1191 6020 1230
rect 6050 1430 6084 1469
rect 6050 1402 6053 1430
rect 6081 1402 6084 1430
rect 6050 1344 6084 1402
rect 6050 1316 6053 1344
rect 6081 1316 6084 1344
rect 6050 1258 6084 1316
rect 6050 1230 6053 1258
rect 6081 1230 6084 1258
rect 6050 1191 6084 1230
rect 6114 1430 6148 1469
rect 6114 1402 6117 1430
rect 6145 1402 6148 1430
rect 6114 1344 6148 1402
rect 6114 1316 6117 1344
rect 6145 1316 6148 1344
rect 6114 1258 6148 1316
rect 6114 1230 6117 1258
rect 6145 1230 6148 1258
rect 6114 1191 6148 1230
rect 6178 1430 6212 1469
rect 6178 1402 6181 1430
rect 6209 1402 6212 1430
rect 6178 1344 6212 1402
rect 6178 1316 6181 1344
rect 6209 1316 6212 1344
rect 6178 1258 6212 1316
rect 6178 1230 6181 1258
rect 6209 1230 6212 1258
rect 6178 1191 6212 1230
rect 6242 1430 6276 1469
rect 6242 1402 6245 1430
rect 6273 1402 6276 1430
rect 6242 1344 6276 1402
rect 6242 1316 6245 1344
rect 6273 1316 6276 1344
rect 6242 1258 6276 1316
rect 6242 1230 6245 1258
rect 6273 1230 6276 1258
rect 6242 1191 6276 1230
rect 6306 1430 6340 1469
rect 6306 1402 6309 1430
rect 6337 1402 6340 1430
rect 6306 1344 6340 1402
rect 6306 1316 6309 1344
rect 6337 1316 6340 1344
rect 6306 1258 6340 1316
rect 6306 1230 6309 1258
rect 6337 1230 6340 1258
rect 6306 1191 6340 1230
rect 6370 1430 6404 1469
rect 6370 1402 6373 1430
rect 6401 1402 6404 1430
rect 6370 1344 6404 1402
rect 6370 1316 6373 1344
rect 6401 1316 6404 1344
rect 6370 1258 6404 1316
rect 6370 1230 6373 1258
rect 6401 1230 6404 1258
rect 6370 1191 6404 1230
rect 6436 1430 6470 1469
rect 6436 1402 6439 1430
rect 6467 1402 6470 1430
rect 6436 1344 6470 1402
rect 6436 1316 6439 1344
rect 6467 1316 6470 1344
rect 6436 1258 6470 1316
rect 6436 1230 6439 1258
rect 6467 1230 6470 1258
rect 6436 1191 6470 1230
rect 6500 1430 6534 1469
rect 6500 1402 6503 1430
rect 6531 1402 6534 1430
rect 6500 1344 6534 1402
rect 6500 1316 6503 1344
rect 6531 1316 6534 1344
rect 6500 1258 6534 1316
rect 6500 1230 6503 1258
rect 6531 1230 6534 1258
rect 6500 1191 6534 1230
rect 6564 1430 6598 1469
rect 6564 1402 6567 1430
rect 6595 1402 6598 1430
rect 6564 1344 6598 1402
rect 6564 1316 6567 1344
rect 6595 1316 6598 1344
rect 6564 1258 6598 1316
rect 6564 1230 6567 1258
rect 6595 1230 6598 1258
rect 6564 1191 6598 1230
rect 6628 1430 6662 1469
rect 6628 1402 6631 1430
rect 6659 1402 6662 1430
rect 6628 1344 6662 1402
rect 6628 1316 6631 1344
rect 6659 1316 6662 1344
rect 6628 1258 6662 1316
rect 6628 1230 6631 1258
rect 6659 1230 6662 1258
rect 6628 1191 6662 1230
rect 6692 1430 6726 1469
rect 6692 1402 6695 1430
rect 6723 1402 6726 1430
rect 6692 1344 6726 1402
rect 6692 1316 6695 1344
rect 6723 1316 6726 1344
rect 6692 1258 6726 1316
rect 6692 1230 6695 1258
rect 6723 1230 6726 1258
rect 6692 1191 6726 1230
rect 6756 1430 6790 1469
rect 6756 1402 6759 1430
rect 6787 1402 6790 1430
rect 6756 1344 6790 1402
rect 6756 1316 6759 1344
rect 6787 1316 6790 1344
rect 6756 1258 6790 1316
rect 6756 1230 6759 1258
rect 6787 1230 6790 1258
rect 6756 1191 6790 1230
rect 6820 1430 6854 1469
rect 6820 1402 6823 1430
rect 6851 1402 6854 1430
rect 6820 1344 6854 1402
rect 6820 1316 6823 1344
rect 6851 1316 6854 1344
rect 6820 1258 6854 1316
rect 6820 1230 6823 1258
rect 6851 1230 6854 1258
rect 6820 1191 6854 1230
rect 6884 1430 6918 1469
rect 6884 1402 6887 1430
rect 6915 1402 6918 1430
rect 6884 1344 6918 1402
rect 6884 1316 6887 1344
rect 6915 1316 6918 1344
rect 6884 1258 6918 1316
rect 6884 1230 6887 1258
rect 6915 1230 6918 1258
rect 6884 1191 6918 1230
rect 6948 1430 6982 1469
rect 6948 1402 6951 1430
rect 6979 1402 6982 1430
rect 6948 1344 6982 1402
rect 6948 1316 6951 1344
rect 6979 1316 6982 1344
rect 6948 1258 6982 1316
rect 6948 1230 6951 1258
rect 6979 1230 6982 1258
rect 6948 1191 6982 1230
rect 7012 1430 7046 1469
rect 7012 1402 7015 1430
rect 7043 1402 7046 1430
rect 7012 1344 7046 1402
rect 7012 1316 7015 1344
rect 7043 1316 7046 1344
rect 7012 1258 7046 1316
rect 7012 1230 7015 1258
rect 7043 1230 7046 1258
rect 7012 1191 7046 1230
rect 7078 1430 7112 1469
rect 7078 1402 7081 1430
rect 7109 1402 7112 1430
rect 7078 1344 7112 1402
rect 7078 1316 7081 1344
rect 7109 1316 7112 1344
rect 7078 1258 7112 1316
rect 7078 1230 7081 1258
rect 7109 1230 7112 1258
rect 7078 1191 7112 1230
rect 7142 1430 7176 1469
rect 7142 1402 7145 1430
rect 7173 1402 7176 1430
rect 7142 1344 7176 1402
rect 7142 1316 7145 1344
rect 7173 1316 7176 1344
rect 7142 1258 7176 1316
rect 7142 1230 7145 1258
rect 7173 1230 7176 1258
rect 7142 1191 7176 1230
rect 7206 1430 7240 1469
rect 7206 1402 7209 1430
rect 7237 1402 7240 1430
rect 7206 1344 7240 1402
rect 7206 1316 7209 1344
rect 7237 1316 7240 1344
rect 7206 1258 7240 1316
rect 7206 1230 7209 1258
rect 7237 1230 7240 1258
rect 7206 1191 7240 1230
rect 7270 1430 7304 1469
rect 7270 1402 7273 1430
rect 7301 1402 7304 1430
rect 7270 1344 7304 1402
rect 7270 1316 7273 1344
rect 7301 1316 7304 1344
rect 7270 1258 7304 1316
rect 7270 1230 7273 1258
rect 7301 1230 7304 1258
rect 7270 1191 7304 1230
rect 7334 1430 7368 1469
rect 7334 1402 7337 1430
rect 7365 1402 7368 1430
rect 7334 1344 7368 1402
rect 7334 1316 7337 1344
rect 7365 1316 7368 1344
rect 7334 1258 7368 1316
rect 7334 1230 7337 1258
rect 7365 1230 7368 1258
rect 7334 1191 7368 1230
rect 7398 1430 7432 1469
rect 7398 1402 7401 1430
rect 7429 1402 7432 1430
rect 7398 1344 7432 1402
rect 7398 1316 7401 1344
rect 7429 1316 7432 1344
rect 7398 1258 7432 1316
rect 7398 1230 7401 1258
rect 7429 1230 7432 1258
rect 7398 1191 7432 1230
rect 7462 1430 7496 1469
rect 7462 1402 7465 1430
rect 7493 1402 7496 1430
rect 7462 1344 7496 1402
rect 7462 1316 7465 1344
rect 7493 1316 7496 1344
rect 7462 1258 7496 1316
rect 7462 1230 7465 1258
rect 7493 1230 7496 1258
rect 7462 1191 7496 1230
rect 7526 1430 7560 1469
rect 7526 1402 7529 1430
rect 7557 1402 7560 1430
rect 7526 1344 7560 1402
rect 7526 1316 7529 1344
rect 7557 1316 7560 1344
rect 7526 1258 7560 1316
rect 7526 1230 7529 1258
rect 7557 1230 7560 1258
rect 7526 1191 7560 1230
rect 7590 1430 7624 1469
rect 7590 1402 7593 1430
rect 7621 1402 7624 1430
rect 7590 1344 7624 1402
rect 7590 1316 7593 1344
rect 7621 1316 7624 1344
rect 7590 1258 7624 1316
rect 7590 1230 7593 1258
rect 7621 1230 7624 1258
rect 7590 1191 7624 1230
rect 7654 1430 7688 1469
rect 7654 1402 7657 1430
rect 7685 1402 7688 1430
rect 7654 1344 7688 1402
rect 7654 1316 7657 1344
rect 7685 1316 7688 1344
rect 7654 1258 7688 1316
rect 7654 1230 7657 1258
rect 7685 1230 7688 1258
rect 7654 1191 7688 1230
rect 7720 1430 7754 1469
rect 7720 1402 7723 1430
rect 7751 1402 7754 1430
rect 7720 1344 7754 1402
rect 7720 1316 7723 1344
rect 7751 1316 7754 1344
rect 7720 1258 7754 1316
rect 7720 1230 7723 1258
rect 7751 1230 7754 1258
rect 7720 1191 7754 1230
rect 7784 1430 7818 1469
rect 7784 1402 7787 1430
rect 7815 1402 7818 1430
rect 7784 1344 7818 1402
rect 7784 1316 7787 1344
rect 7815 1316 7818 1344
rect 7784 1258 7818 1316
rect 7784 1230 7787 1258
rect 7815 1230 7818 1258
rect 7784 1191 7818 1230
rect 7848 1430 7882 1469
rect 7848 1402 7851 1430
rect 7879 1402 7882 1430
rect 7848 1344 7882 1402
rect 7848 1316 7851 1344
rect 7879 1316 7882 1344
rect 7848 1258 7882 1316
rect 7848 1230 7851 1258
rect 7879 1230 7882 1258
rect 7848 1191 7882 1230
rect 7912 1430 7946 1469
rect 7912 1402 7915 1430
rect 7943 1402 7946 1430
rect 7912 1344 7946 1402
rect 7912 1316 7915 1344
rect 7943 1316 7946 1344
rect 7912 1258 7946 1316
rect 7912 1230 7915 1258
rect 7943 1230 7946 1258
rect 7912 1191 7946 1230
rect 7976 1430 8010 1469
rect 7976 1402 7979 1430
rect 8007 1402 8010 1430
rect 7976 1344 8010 1402
rect 7976 1316 7979 1344
rect 8007 1316 8010 1344
rect 7976 1258 8010 1316
rect 7976 1230 7979 1258
rect 8007 1230 8010 1258
rect 7976 1191 8010 1230
rect 8040 1430 8074 1469
rect 8040 1402 8043 1430
rect 8071 1402 8074 1430
rect 8040 1344 8074 1402
rect 8040 1316 8043 1344
rect 8071 1316 8074 1344
rect 8040 1258 8074 1316
rect 8040 1230 8043 1258
rect 8071 1230 8074 1258
rect 8040 1191 8074 1230
rect 8104 1430 8138 1469
rect 8104 1402 8107 1430
rect 8135 1402 8138 1430
rect 8104 1344 8138 1402
rect 8104 1316 8107 1344
rect 8135 1316 8138 1344
rect 8104 1258 8138 1316
rect 8104 1230 8107 1258
rect 8135 1230 8138 1258
rect 8104 1191 8138 1230
rect 8168 1430 8202 1469
rect 8168 1402 8171 1430
rect 8199 1402 8202 1430
rect 8168 1344 8202 1402
rect 8168 1316 8171 1344
rect 8199 1316 8202 1344
rect 8168 1258 8202 1316
rect 8168 1230 8171 1258
rect 8199 1230 8202 1258
rect 8168 1191 8202 1230
rect 8232 1430 8266 1469
rect 8232 1402 8235 1430
rect 8263 1402 8266 1430
rect 8232 1344 8266 1402
rect 8232 1316 8235 1344
rect 8263 1316 8266 1344
rect 8232 1258 8266 1316
rect 8232 1230 8235 1258
rect 8263 1230 8266 1258
rect 8232 1191 8266 1230
rect 8296 1430 8330 1469
rect 8296 1402 8299 1430
rect 8327 1402 8330 1430
rect 8296 1344 8330 1402
rect 8296 1316 8299 1344
rect 8327 1316 8330 1344
rect 8296 1258 8330 1316
rect 8296 1230 8299 1258
rect 8327 1230 8330 1258
rect 8296 1191 8330 1230
rect 8362 1430 8396 1469
rect 8362 1402 8365 1430
rect 8393 1402 8396 1430
rect 8362 1344 8396 1402
rect 8362 1316 8365 1344
rect 8393 1316 8396 1344
rect 8362 1258 8396 1316
rect 8362 1230 8365 1258
rect 8393 1230 8396 1258
rect 8362 1191 8396 1230
rect 8426 1430 8460 1469
rect 8426 1402 8429 1430
rect 8457 1402 8460 1430
rect 8426 1344 8460 1402
rect 8426 1316 8429 1344
rect 8457 1316 8460 1344
rect 8426 1258 8460 1316
rect 8426 1230 8429 1258
rect 8457 1230 8460 1258
rect 8426 1191 8460 1230
rect 8490 1430 8524 1469
rect 8490 1402 8493 1430
rect 8521 1402 8524 1430
rect 8490 1344 8524 1402
rect 8490 1316 8493 1344
rect 8521 1316 8524 1344
rect 8490 1258 8524 1316
rect 8490 1230 8493 1258
rect 8521 1230 8524 1258
rect 8490 1191 8524 1230
rect 8554 1430 8588 1469
rect 8554 1402 8557 1430
rect 8585 1402 8588 1430
rect 8554 1344 8588 1402
rect 8554 1316 8557 1344
rect 8585 1316 8588 1344
rect 8554 1258 8588 1316
rect 8554 1230 8557 1258
rect 8585 1230 8588 1258
rect 8554 1191 8588 1230
rect 8618 1430 8652 1469
rect 8618 1402 8621 1430
rect 8649 1402 8652 1430
rect 8618 1344 8652 1402
rect 8618 1316 8621 1344
rect 8649 1316 8652 1344
rect 8618 1258 8652 1316
rect 8618 1230 8621 1258
rect 8649 1230 8652 1258
rect 8618 1191 8652 1230
rect 8682 1430 8716 1469
rect 8682 1402 8685 1430
rect 8713 1402 8716 1430
rect 8682 1344 8716 1402
rect 8682 1316 8685 1344
rect 8713 1316 8716 1344
rect 8682 1258 8716 1316
rect 8682 1230 8685 1258
rect 8713 1230 8716 1258
rect 8682 1191 8716 1230
rect 8746 1430 8780 1469
rect 8746 1402 8749 1430
rect 8777 1402 8780 1430
rect 8746 1344 8780 1402
rect 8746 1316 8749 1344
rect 8777 1316 8780 1344
rect 8746 1258 8780 1316
rect 8746 1230 8749 1258
rect 8777 1230 8780 1258
rect 8746 1191 8780 1230
rect 8810 1430 8844 1469
rect 8810 1402 8813 1430
rect 8841 1402 8844 1430
rect 8810 1344 8844 1402
rect 8810 1316 8813 1344
rect 8841 1316 8844 1344
rect 8810 1258 8844 1316
rect 8810 1230 8813 1258
rect 8841 1230 8844 1258
rect 8810 1191 8844 1230
rect 8874 1430 8908 1469
rect 8874 1402 8877 1430
rect 8905 1402 8908 1430
rect 8874 1344 8908 1402
rect 8874 1316 8877 1344
rect 8905 1316 8908 1344
rect 8874 1258 8908 1316
rect 8874 1230 8877 1258
rect 8905 1230 8908 1258
rect 8874 1191 8908 1230
rect 8938 1430 8972 1469
rect 8938 1402 8941 1430
rect 8969 1402 8972 1430
rect 8938 1344 8972 1402
rect 8938 1316 8941 1344
rect 8969 1316 8972 1344
rect 8938 1258 8972 1316
rect 8938 1230 8941 1258
rect 8969 1230 8972 1258
rect 8938 1191 8972 1230
rect 9004 1430 9038 1469
rect 9004 1402 9007 1430
rect 9035 1402 9038 1430
rect 9004 1344 9038 1402
rect 9004 1316 9007 1344
rect 9035 1316 9038 1344
rect 9004 1258 9038 1316
rect 9004 1230 9007 1258
rect 9035 1230 9038 1258
rect 9004 1191 9038 1230
rect 9068 1430 9102 1469
rect 9068 1402 9071 1430
rect 9099 1402 9102 1430
rect 9068 1344 9102 1402
rect 9068 1316 9071 1344
rect 9099 1316 9102 1344
rect 9068 1258 9102 1316
rect 9068 1230 9071 1258
rect 9099 1230 9102 1258
rect 9068 1191 9102 1230
rect 9132 1430 9166 1469
rect 9132 1402 9135 1430
rect 9163 1402 9166 1430
rect 9132 1344 9166 1402
rect 9132 1316 9135 1344
rect 9163 1316 9166 1344
rect 9132 1258 9166 1316
rect 9132 1230 9135 1258
rect 9163 1230 9166 1258
rect 9132 1191 9166 1230
rect 9196 1430 9230 1469
rect 9196 1402 9199 1430
rect 9227 1402 9230 1430
rect 9196 1344 9230 1402
rect 9196 1316 9199 1344
rect 9227 1316 9230 1344
rect 9196 1258 9230 1316
rect 9196 1230 9199 1258
rect 9227 1230 9230 1258
rect 9196 1191 9230 1230
rect 9260 1430 9294 1469
rect 9260 1402 9263 1430
rect 9291 1402 9294 1430
rect 9260 1344 9294 1402
rect 9260 1316 9263 1344
rect 9291 1316 9294 1344
rect 9260 1258 9294 1316
rect 9260 1230 9263 1258
rect 9291 1230 9294 1258
rect 9260 1191 9294 1230
rect 9324 1430 9358 1469
rect 9324 1402 9327 1430
rect 9355 1402 9358 1430
rect 9324 1344 9358 1402
rect 9324 1316 9327 1344
rect 9355 1316 9358 1344
rect 9324 1258 9358 1316
rect 9324 1230 9327 1258
rect 9355 1230 9358 1258
rect 9324 1191 9358 1230
rect 9388 1430 9422 1469
rect 9388 1402 9391 1430
rect 9419 1402 9422 1430
rect 9388 1344 9422 1402
rect 9388 1316 9391 1344
rect 9419 1316 9422 1344
rect 9388 1258 9422 1316
rect 9388 1230 9391 1258
rect 9419 1230 9422 1258
rect 9388 1191 9422 1230
rect 9452 1430 9486 1469
rect 9452 1402 9455 1430
rect 9483 1402 9486 1430
rect 9452 1344 9486 1402
rect 9452 1316 9455 1344
rect 9483 1316 9486 1344
rect 9452 1258 9486 1316
rect 9452 1230 9455 1258
rect 9483 1230 9486 1258
rect 9452 1191 9486 1230
rect 9516 1430 9550 1469
rect 9516 1402 9519 1430
rect 9547 1402 9550 1430
rect 9516 1344 9550 1402
rect 9516 1316 9519 1344
rect 9547 1316 9550 1344
rect 9516 1258 9550 1316
rect 9516 1230 9519 1258
rect 9547 1230 9550 1258
rect 9516 1191 9550 1230
rect 9580 1430 9614 1469
rect 9580 1402 9583 1430
rect 9611 1402 9614 1430
rect 9580 1344 9614 1402
rect 9580 1316 9583 1344
rect 9611 1316 9614 1344
rect 9580 1258 9614 1316
rect 9580 1230 9583 1258
rect 9611 1230 9614 1258
rect 9580 1191 9614 1230
rect 9646 1430 9680 1469
rect 9646 1402 9649 1430
rect 9677 1402 9680 1430
rect 9646 1344 9680 1402
rect 9646 1316 9649 1344
rect 9677 1316 9680 1344
rect 9646 1258 9680 1316
rect 9646 1230 9649 1258
rect 9677 1230 9680 1258
rect 9646 1191 9680 1230
rect 9710 1430 9744 1469
rect 9710 1402 9713 1430
rect 9741 1402 9744 1430
rect 9710 1344 9744 1402
rect 9710 1316 9713 1344
rect 9741 1316 9744 1344
rect 9710 1258 9744 1316
rect 9710 1230 9713 1258
rect 9741 1230 9744 1258
rect 9710 1191 9744 1230
rect 9774 1430 9808 1469
rect 9774 1402 9777 1430
rect 9805 1402 9808 1430
rect 9774 1344 9808 1402
rect 9774 1316 9777 1344
rect 9805 1316 9808 1344
rect 9774 1258 9808 1316
rect 9774 1230 9777 1258
rect 9805 1230 9808 1258
rect 9774 1191 9808 1230
rect 9838 1430 9872 1469
rect 9838 1402 9841 1430
rect 9869 1402 9872 1430
rect 9838 1344 9872 1402
rect 9838 1316 9841 1344
rect 9869 1316 9872 1344
rect 9838 1258 9872 1316
rect 9838 1230 9841 1258
rect 9869 1230 9872 1258
rect 9838 1191 9872 1230
rect 9902 1430 9936 1469
rect 9902 1402 9905 1430
rect 9933 1402 9936 1430
rect 9902 1344 9936 1402
rect 9902 1316 9905 1344
rect 9933 1316 9936 1344
rect 9902 1258 9936 1316
rect 9902 1230 9905 1258
rect 9933 1230 9936 1258
rect 9902 1191 9936 1230
rect 9966 1430 10000 1469
rect 9966 1402 9969 1430
rect 9997 1402 10000 1430
rect 9966 1344 10000 1402
rect 9966 1316 9969 1344
rect 9997 1316 10000 1344
rect 9966 1258 10000 1316
rect 9966 1230 9969 1258
rect 9997 1230 10000 1258
rect 9966 1191 10000 1230
rect 10030 1430 10064 1469
rect 10030 1402 10033 1430
rect 10061 1402 10064 1430
rect 10030 1344 10064 1402
rect 10030 1316 10033 1344
rect 10061 1316 10064 1344
rect 10030 1258 10064 1316
rect 10030 1230 10033 1258
rect 10061 1230 10064 1258
rect 10030 1191 10064 1230
rect 10094 1430 10128 1469
rect 10094 1402 10097 1430
rect 10125 1402 10128 1430
rect 10094 1344 10128 1402
rect 10094 1316 10097 1344
rect 10125 1316 10128 1344
rect 10094 1258 10128 1316
rect 10094 1230 10097 1258
rect 10125 1230 10128 1258
rect 10094 1191 10128 1230
rect 10158 1430 10192 1469
rect 10158 1402 10161 1430
rect 10189 1402 10192 1430
rect 10158 1344 10192 1402
rect 10158 1316 10161 1344
rect 10189 1316 10192 1344
rect 10158 1258 10192 1316
rect 10158 1230 10161 1258
rect 10189 1230 10192 1258
rect 10158 1191 10192 1230
rect 10222 1430 10256 1469
rect 10222 1402 10225 1430
rect 10253 1402 10256 1430
rect 10222 1344 10256 1402
rect 10222 1316 10225 1344
rect 10253 1316 10256 1344
rect 10222 1258 10256 1316
rect 10222 1230 10225 1258
rect 10253 1230 10256 1258
rect 10222 1191 10256 1230
rect 10288 1430 10322 1469
rect 10288 1402 10291 1430
rect 10319 1402 10322 1430
rect 10288 1344 10322 1402
rect 10288 1316 10291 1344
rect 10319 1316 10322 1344
rect 10288 1258 10322 1316
rect 10288 1230 10291 1258
rect 10319 1230 10322 1258
rect 10288 1191 10322 1230
rect 10352 1430 10386 1469
rect 10352 1402 10355 1430
rect 10383 1402 10386 1430
rect 10352 1344 10386 1402
rect 10352 1316 10355 1344
rect 10383 1316 10386 1344
rect 10352 1258 10386 1316
rect 10352 1230 10355 1258
rect 10383 1230 10386 1258
rect 10352 1191 10386 1230
rect 10416 1430 10450 1469
rect 10416 1402 10419 1430
rect 10447 1402 10450 1430
rect 10416 1344 10450 1402
rect 10416 1316 10419 1344
rect 10447 1316 10450 1344
rect 10416 1258 10450 1316
rect 10416 1230 10419 1258
rect 10447 1230 10450 1258
rect 10416 1191 10450 1230
rect 10480 1430 10514 1469
rect 10480 1402 10483 1430
rect 10511 1402 10514 1430
rect 10480 1344 10514 1402
rect 10480 1316 10483 1344
rect 10511 1316 10514 1344
rect 10480 1258 10514 1316
rect 10480 1230 10483 1258
rect 10511 1230 10514 1258
rect 10480 1191 10514 1230
rect 10544 1430 10578 1469
rect 10544 1402 10547 1430
rect 10575 1402 10578 1430
rect 10544 1344 10578 1402
rect 10544 1316 10547 1344
rect 10575 1316 10578 1344
rect 10544 1258 10578 1316
rect 10544 1230 10547 1258
rect 10575 1230 10578 1258
rect 10544 1191 10578 1230
rect 10608 1430 10642 1469
rect 10608 1402 10611 1430
rect 10639 1402 10642 1430
rect 10608 1344 10642 1402
rect 10608 1316 10611 1344
rect 10639 1316 10642 1344
rect 10608 1258 10642 1316
rect 10608 1230 10611 1258
rect 10639 1230 10642 1258
rect 10608 1191 10642 1230
rect 10672 1430 10706 1469
rect 10672 1402 10675 1430
rect 10703 1402 10706 1430
rect 10672 1344 10706 1402
rect 10672 1316 10675 1344
rect 10703 1316 10706 1344
rect 10672 1258 10706 1316
rect 10672 1230 10675 1258
rect 10703 1230 10706 1258
rect 10672 1191 10706 1230
rect 10736 1430 10770 1469
rect 10736 1402 10739 1430
rect 10767 1402 10770 1430
rect 10736 1344 10770 1402
rect 10736 1316 10739 1344
rect 10767 1316 10770 1344
rect 10736 1258 10770 1316
rect 10736 1230 10739 1258
rect 10767 1230 10770 1258
rect 10736 1191 10770 1230
rect 10800 1430 10834 1469
rect 10800 1402 10803 1430
rect 10831 1402 10834 1430
rect 10800 1344 10834 1402
rect 10800 1316 10803 1344
rect 10831 1316 10834 1344
rect 10800 1258 10834 1316
rect 10800 1230 10803 1258
rect 10831 1230 10834 1258
rect 10800 1191 10834 1230
rect 10864 1430 10898 1469
rect 10864 1402 10867 1430
rect 10895 1402 10898 1430
rect 10864 1344 10898 1402
rect 10864 1316 10867 1344
rect 10895 1316 10898 1344
rect 10864 1258 10898 1316
rect 10864 1230 10867 1258
rect 10895 1230 10898 1258
rect 10864 1191 10898 1230
rect 10930 1430 10964 1469
rect 10930 1402 10933 1430
rect 10961 1402 10964 1430
rect 10930 1344 10964 1402
rect 10930 1316 10933 1344
rect 10961 1316 10964 1344
rect 10930 1258 10964 1316
rect 10930 1230 10933 1258
rect 10961 1230 10964 1258
rect 10930 1191 10964 1230
rect 10994 1430 11028 1469
rect 10994 1402 10997 1430
rect 11025 1402 11028 1430
rect 10994 1344 11028 1402
rect 10994 1316 10997 1344
rect 11025 1316 11028 1344
rect 10994 1258 11028 1316
rect 10994 1230 10997 1258
rect 11025 1230 11028 1258
rect 10994 1191 11028 1230
rect 11058 1430 11092 1469
rect 11058 1402 11061 1430
rect 11089 1402 11092 1430
rect 11058 1344 11092 1402
rect 11058 1316 11061 1344
rect 11089 1316 11092 1344
rect 11058 1258 11092 1316
rect 11058 1230 11061 1258
rect 11089 1230 11092 1258
rect 11058 1191 11092 1230
rect 11122 1430 11156 1469
rect 11122 1402 11125 1430
rect 11153 1402 11156 1430
rect 11122 1344 11156 1402
rect 11122 1316 11125 1344
rect 11153 1316 11156 1344
rect 11122 1258 11156 1316
rect 11122 1230 11125 1258
rect 11153 1230 11156 1258
rect 11122 1191 11156 1230
rect 11186 1430 11220 1469
rect 11186 1402 11189 1430
rect 11217 1402 11220 1430
rect 11186 1344 11220 1402
rect 11186 1316 11189 1344
rect 11217 1316 11220 1344
rect 11186 1258 11220 1316
rect 11186 1230 11189 1258
rect 11217 1230 11220 1258
rect 11186 1191 11220 1230
rect 11250 1430 11284 1469
rect 11250 1402 11253 1430
rect 11281 1402 11284 1430
rect 11250 1344 11284 1402
rect 11250 1316 11253 1344
rect 11281 1316 11284 1344
rect 11250 1258 11284 1316
rect 11250 1230 11253 1258
rect 11281 1230 11284 1258
rect 11250 1191 11284 1230
rect 11314 1430 11348 1469
rect 11314 1402 11317 1430
rect 11345 1402 11348 1430
rect 11314 1344 11348 1402
rect 11314 1316 11317 1344
rect 11345 1316 11348 1344
rect 11314 1258 11348 1316
rect 11314 1230 11317 1258
rect 11345 1230 11348 1258
rect 11314 1191 11348 1230
rect 11378 1430 11412 1469
rect 11378 1402 11381 1430
rect 11409 1402 11412 1430
rect 11378 1344 11412 1402
rect 11378 1316 11381 1344
rect 11409 1316 11412 1344
rect 11378 1258 11412 1316
rect 11378 1230 11381 1258
rect 11409 1230 11412 1258
rect 11378 1191 11412 1230
rect 11442 1430 11476 1469
rect 11442 1402 11445 1430
rect 11473 1402 11476 1430
rect 11442 1344 11476 1402
rect 11442 1316 11445 1344
rect 11473 1316 11476 1344
rect 11442 1258 11476 1316
rect 11442 1230 11445 1258
rect 11473 1230 11476 1258
rect 11442 1191 11476 1230
rect 11506 1430 11540 1469
rect 11506 1402 11509 1430
rect 11537 1402 11540 1430
rect 11506 1344 11540 1402
rect 11506 1316 11509 1344
rect 11537 1316 11540 1344
rect 11506 1258 11540 1316
rect 11506 1230 11509 1258
rect 11537 1230 11540 1258
rect 11506 1191 11540 1230
rect 11572 1430 11606 1469
rect 11572 1402 11575 1430
rect 11603 1402 11606 1430
rect 11572 1344 11606 1402
rect 11572 1316 11575 1344
rect 11603 1316 11606 1344
rect 11572 1258 11606 1316
rect 11572 1230 11575 1258
rect 11603 1230 11606 1258
rect 11572 1191 11606 1230
rect 11636 1430 11670 1469
rect 11636 1402 11639 1430
rect 11667 1402 11670 1430
rect 11636 1344 11670 1402
rect 11636 1316 11639 1344
rect 11667 1316 11670 1344
rect 11636 1258 11670 1316
rect 11636 1230 11639 1258
rect 11667 1230 11670 1258
rect 11636 1191 11670 1230
rect 11700 1430 11734 1469
rect 11700 1402 11703 1430
rect 11731 1402 11734 1430
rect 11700 1344 11734 1402
rect 11700 1316 11703 1344
rect 11731 1316 11734 1344
rect 11700 1258 11734 1316
rect 11700 1230 11703 1258
rect 11731 1230 11734 1258
rect 11700 1191 11734 1230
rect 11764 1430 11798 1469
rect 11764 1402 11767 1430
rect 11795 1402 11798 1430
rect 11764 1344 11798 1402
rect 11764 1316 11767 1344
rect 11795 1316 11798 1344
rect 11764 1258 11798 1316
rect 11764 1230 11767 1258
rect 11795 1230 11798 1258
rect 11764 1191 11798 1230
rect 11828 1430 11862 1469
rect 11828 1402 11831 1430
rect 11859 1402 11862 1430
rect 11828 1344 11862 1402
rect 11828 1316 11831 1344
rect 11859 1316 11862 1344
rect 11828 1258 11862 1316
rect 11828 1230 11831 1258
rect 11859 1230 11862 1258
rect 11828 1191 11862 1230
rect 11892 1430 11926 1469
rect 11892 1402 11895 1430
rect 11923 1402 11926 1430
rect 11892 1344 11926 1402
rect 11892 1316 11895 1344
rect 11923 1316 11926 1344
rect 11892 1258 11926 1316
rect 11892 1230 11895 1258
rect 11923 1230 11926 1258
rect 11892 1191 11926 1230
rect 11956 1430 11990 1469
rect 11956 1402 11959 1430
rect 11987 1402 11990 1430
rect 11956 1344 11990 1402
rect 11956 1316 11959 1344
rect 11987 1316 11990 1344
rect 11956 1258 11990 1316
rect 11956 1230 11959 1258
rect 11987 1230 11990 1258
rect 11956 1191 11990 1230
rect 12020 1430 12054 1469
rect 12020 1402 12023 1430
rect 12051 1402 12054 1430
rect 12020 1344 12054 1402
rect 12020 1316 12023 1344
rect 12051 1316 12054 1344
rect 12020 1258 12054 1316
rect 12020 1230 12023 1258
rect 12051 1230 12054 1258
rect 12020 1191 12054 1230
rect 12084 1430 12118 1469
rect 12084 1402 12087 1430
rect 12115 1402 12118 1430
rect 12084 1344 12118 1402
rect 12084 1316 12087 1344
rect 12115 1316 12118 1344
rect 12084 1258 12118 1316
rect 12084 1230 12087 1258
rect 12115 1230 12118 1258
rect 12084 1191 12118 1230
rect 12148 1430 12182 1469
rect 12148 1402 12151 1430
rect 12179 1402 12182 1430
rect 12148 1344 12182 1402
rect 12148 1316 12151 1344
rect 12179 1316 12182 1344
rect 12148 1258 12182 1316
rect 12148 1230 12151 1258
rect 12179 1230 12182 1258
rect 12148 1191 12182 1230
rect 12214 1430 12248 1469
rect 12214 1402 12217 1430
rect 12245 1402 12248 1430
rect 12214 1344 12248 1402
rect 12214 1316 12217 1344
rect 12245 1316 12248 1344
rect 12214 1258 12248 1316
rect 12214 1230 12217 1258
rect 12245 1230 12248 1258
rect 12214 1191 12248 1230
rect 12278 1430 12312 1469
rect 12278 1402 12281 1430
rect 12309 1402 12312 1430
rect 12278 1344 12312 1402
rect 12278 1316 12281 1344
rect 12309 1316 12312 1344
rect 12278 1258 12312 1316
rect 12278 1230 12281 1258
rect 12309 1230 12312 1258
rect 12278 1191 12312 1230
rect 12342 1430 12376 1469
rect 12342 1402 12345 1430
rect 12373 1402 12376 1430
rect 12342 1344 12376 1402
rect 12342 1316 12345 1344
rect 12373 1316 12376 1344
rect 12342 1258 12376 1316
rect 12342 1230 12345 1258
rect 12373 1230 12376 1258
rect 12342 1191 12376 1230
rect 12406 1430 12440 1469
rect 12406 1402 12409 1430
rect 12437 1402 12440 1430
rect 12406 1344 12440 1402
rect 12406 1316 12409 1344
rect 12437 1316 12440 1344
rect 12406 1258 12440 1316
rect 12406 1230 12409 1258
rect 12437 1230 12440 1258
rect 12406 1191 12440 1230
rect 12470 1430 12504 1469
rect 12470 1402 12473 1430
rect 12501 1402 12504 1430
rect 12470 1344 12504 1402
rect 12470 1316 12473 1344
rect 12501 1316 12504 1344
rect 12470 1258 12504 1316
rect 12470 1230 12473 1258
rect 12501 1230 12504 1258
rect 12470 1191 12504 1230
rect 12534 1430 12568 1469
rect 12534 1402 12537 1430
rect 12565 1402 12568 1430
rect 12534 1344 12568 1402
rect 12534 1316 12537 1344
rect 12565 1316 12568 1344
rect 12534 1258 12568 1316
rect 12534 1230 12537 1258
rect 12565 1230 12568 1258
rect 12534 1191 12568 1230
rect 12598 1430 12632 1469
rect 12598 1402 12601 1430
rect 12629 1402 12632 1430
rect 12598 1344 12632 1402
rect 12598 1316 12601 1344
rect 12629 1316 12632 1344
rect 12598 1258 12632 1316
rect 12598 1230 12601 1258
rect 12629 1230 12632 1258
rect 12598 1191 12632 1230
rect 12662 1430 12696 1469
rect 12662 1402 12665 1430
rect 12693 1402 12696 1430
rect 12662 1344 12696 1402
rect 12662 1316 12665 1344
rect 12693 1316 12696 1344
rect 12662 1258 12696 1316
rect 12662 1230 12665 1258
rect 12693 1230 12696 1258
rect 12662 1191 12696 1230
rect 12726 1430 12760 1469
rect 12726 1402 12729 1430
rect 12757 1402 12760 1430
rect 12726 1344 12760 1402
rect 12726 1316 12729 1344
rect 12757 1316 12760 1344
rect 12726 1258 12760 1316
rect 12726 1230 12729 1258
rect 12757 1230 12760 1258
rect 12726 1191 12760 1230
rect 12790 1430 12824 1469
rect 12790 1402 12793 1430
rect 12821 1402 12824 1430
rect 12790 1344 12824 1402
rect 12790 1316 12793 1344
rect 12821 1316 12824 1344
rect 12790 1258 12824 1316
rect 12790 1230 12793 1258
rect 12821 1230 12824 1258
rect 12790 1191 12824 1230
rect 16 1050 50 1089
rect 16 1022 19 1050
rect 47 1022 50 1050
rect 16 964 50 1022
rect 16 936 19 964
rect 47 936 50 964
rect 16 878 50 936
rect 16 850 19 878
rect 47 850 50 878
rect 16 811 50 850
rect 80 1050 114 1089
rect 80 1022 83 1050
rect 111 1022 114 1050
rect 80 964 114 1022
rect 80 936 83 964
rect 111 936 114 964
rect 80 878 114 936
rect 80 850 83 878
rect 111 850 114 878
rect 80 811 114 850
rect 144 1050 178 1089
rect 144 1022 147 1050
rect 175 1022 178 1050
rect 144 964 178 1022
rect 144 936 147 964
rect 175 936 178 964
rect 144 878 178 936
rect 144 850 147 878
rect 175 850 178 878
rect 144 811 178 850
rect 208 1050 242 1089
rect 208 1022 211 1050
rect 239 1022 242 1050
rect 208 964 242 1022
rect 208 936 211 964
rect 239 936 242 964
rect 208 878 242 936
rect 208 850 211 878
rect 239 850 242 878
rect 208 811 242 850
rect 272 1050 306 1089
rect 272 1022 275 1050
rect 303 1022 306 1050
rect 272 964 306 1022
rect 272 936 275 964
rect 303 936 306 964
rect 272 878 306 936
rect 272 850 275 878
rect 303 850 306 878
rect 272 811 306 850
rect 336 1050 370 1089
rect 336 1022 339 1050
rect 367 1022 370 1050
rect 336 964 370 1022
rect 336 936 339 964
rect 367 936 370 964
rect 336 878 370 936
rect 336 850 339 878
rect 367 850 370 878
rect 336 811 370 850
rect 400 1050 434 1089
rect 400 1022 403 1050
rect 431 1022 434 1050
rect 400 964 434 1022
rect 400 936 403 964
rect 431 936 434 964
rect 400 878 434 936
rect 400 850 403 878
rect 431 850 434 878
rect 400 811 434 850
rect 464 1050 498 1089
rect 464 1022 467 1050
rect 495 1022 498 1050
rect 464 964 498 1022
rect 464 936 467 964
rect 495 936 498 964
rect 464 878 498 936
rect 464 850 467 878
rect 495 850 498 878
rect 464 811 498 850
rect 528 1050 562 1089
rect 528 1022 531 1050
rect 559 1022 562 1050
rect 528 964 562 1022
rect 528 936 531 964
rect 559 936 562 964
rect 528 878 562 936
rect 528 850 531 878
rect 559 850 562 878
rect 528 811 562 850
rect 592 1050 626 1089
rect 592 1022 595 1050
rect 623 1022 626 1050
rect 592 964 626 1022
rect 592 936 595 964
rect 623 936 626 964
rect 592 878 626 936
rect 592 850 595 878
rect 623 850 626 878
rect 592 811 626 850
rect 658 1050 692 1089
rect 658 1022 661 1050
rect 689 1022 692 1050
rect 658 964 692 1022
rect 658 936 661 964
rect 689 936 692 964
rect 658 878 692 936
rect 658 850 661 878
rect 689 850 692 878
rect 658 811 692 850
rect 722 1050 756 1089
rect 722 1022 725 1050
rect 753 1022 756 1050
rect 722 964 756 1022
rect 722 936 725 964
rect 753 936 756 964
rect 722 878 756 936
rect 722 850 725 878
rect 753 850 756 878
rect 722 811 756 850
rect 786 1050 820 1089
rect 786 1022 789 1050
rect 817 1022 820 1050
rect 786 964 820 1022
rect 786 936 789 964
rect 817 936 820 964
rect 786 878 820 936
rect 786 850 789 878
rect 817 850 820 878
rect 786 811 820 850
rect 850 1050 884 1089
rect 850 1022 853 1050
rect 881 1022 884 1050
rect 850 964 884 1022
rect 850 936 853 964
rect 881 936 884 964
rect 850 878 884 936
rect 850 850 853 878
rect 881 850 884 878
rect 850 811 884 850
rect 914 1050 948 1089
rect 914 1022 917 1050
rect 945 1022 948 1050
rect 914 964 948 1022
rect 914 936 917 964
rect 945 936 948 964
rect 914 878 948 936
rect 914 850 917 878
rect 945 850 948 878
rect 914 811 948 850
rect 978 1050 1012 1089
rect 978 1022 981 1050
rect 1009 1022 1012 1050
rect 978 964 1012 1022
rect 978 936 981 964
rect 1009 936 1012 964
rect 978 878 1012 936
rect 978 850 981 878
rect 1009 850 1012 878
rect 978 811 1012 850
rect 1042 1050 1076 1089
rect 1042 1022 1045 1050
rect 1073 1022 1076 1050
rect 1042 964 1076 1022
rect 1042 936 1045 964
rect 1073 936 1076 964
rect 1042 878 1076 936
rect 1042 850 1045 878
rect 1073 850 1076 878
rect 1042 811 1076 850
rect 1106 1050 1140 1089
rect 1106 1022 1109 1050
rect 1137 1022 1140 1050
rect 1106 964 1140 1022
rect 1106 936 1109 964
rect 1137 936 1140 964
rect 1106 878 1140 936
rect 1106 850 1109 878
rect 1137 850 1140 878
rect 1106 811 1140 850
rect 1170 1050 1204 1089
rect 1170 1022 1173 1050
rect 1201 1022 1204 1050
rect 1170 964 1204 1022
rect 1170 936 1173 964
rect 1201 936 1204 964
rect 1170 878 1204 936
rect 1170 850 1173 878
rect 1201 850 1204 878
rect 1170 811 1204 850
rect 1234 1050 1268 1089
rect 1234 1022 1237 1050
rect 1265 1022 1268 1050
rect 1234 964 1268 1022
rect 1234 936 1237 964
rect 1265 936 1268 964
rect 1234 878 1268 936
rect 1234 850 1237 878
rect 1265 850 1268 878
rect 1234 811 1268 850
rect 1300 1050 1334 1089
rect 1300 1022 1303 1050
rect 1331 1022 1334 1050
rect 1300 964 1334 1022
rect 1300 936 1303 964
rect 1331 936 1334 964
rect 1300 878 1334 936
rect 1300 850 1303 878
rect 1331 850 1334 878
rect 1300 811 1334 850
rect 1364 1050 1398 1089
rect 1364 1022 1367 1050
rect 1395 1022 1398 1050
rect 1364 964 1398 1022
rect 1364 936 1367 964
rect 1395 936 1398 964
rect 1364 878 1398 936
rect 1364 850 1367 878
rect 1395 850 1398 878
rect 1364 811 1398 850
rect 1428 1050 1462 1089
rect 1428 1022 1431 1050
rect 1459 1022 1462 1050
rect 1428 964 1462 1022
rect 1428 936 1431 964
rect 1459 936 1462 964
rect 1428 878 1462 936
rect 1428 850 1431 878
rect 1459 850 1462 878
rect 1428 811 1462 850
rect 1492 1050 1526 1089
rect 1492 1022 1495 1050
rect 1523 1022 1526 1050
rect 1492 964 1526 1022
rect 1492 936 1495 964
rect 1523 936 1526 964
rect 1492 878 1526 936
rect 1492 850 1495 878
rect 1523 850 1526 878
rect 1492 811 1526 850
rect 1556 1050 1590 1089
rect 1556 1022 1559 1050
rect 1587 1022 1590 1050
rect 1556 964 1590 1022
rect 1556 936 1559 964
rect 1587 936 1590 964
rect 1556 878 1590 936
rect 1556 850 1559 878
rect 1587 850 1590 878
rect 1556 811 1590 850
rect 1620 1050 1654 1089
rect 1620 1022 1623 1050
rect 1651 1022 1654 1050
rect 1620 964 1654 1022
rect 1620 936 1623 964
rect 1651 936 1654 964
rect 1620 878 1654 936
rect 1620 850 1623 878
rect 1651 850 1654 878
rect 1620 811 1654 850
rect 1684 1050 1718 1089
rect 1684 1022 1687 1050
rect 1715 1022 1718 1050
rect 1684 964 1718 1022
rect 1684 936 1687 964
rect 1715 936 1718 964
rect 1684 878 1718 936
rect 1684 850 1687 878
rect 1715 850 1718 878
rect 1684 811 1718 850
rect 1748 1050 1782 1089
rect 1748 1022 1751 1050
rect 1779 1022 1782 1050
rect 1748 964 1782 1022
rect 1748 936 1751 964
rect 1779 936 1782 964
rect 1748 878 1782 936
rect 1748 850 1751 878
rect 1779 850 1782 878
rect 1748 811 1782 850
rect 1812 1050 1846 1089
rect 1812 1022 1815 1050
rect 1843 1022 1846 1050
rect 1812 964 1846 1022
rect 1812 936 1815 964
rect 1843 936 1846 964
rect 1812 878 1846 936
rect 1812 850 1815 878
rect 1843 850 1846 878
rect 1812 811 1846 850
rect 1876 1050 1910 1089
rect 1876 1022 1879 1050
rect 1907 1022 1910 1050
rect 1876 964 1910 1022
rect 1876 936 1879 964
rect 1907 936 1910 964
rect 1876 878 1910 936
rect 1876 850 1879 878
rect 1907 850 1910 878
rect 1876 811 1910 850
rect 1942 1050 1976 1089
rect 1942 1022 1945 1050
rect 1973 1022 1976 1050
rect 1942 964 1976 1022
rect 1942 936 1945 964
rect 1973 936 1976 964
rect 1942 878 1976 936
rect 1942 850 1945 878
rect 1973 850 1976 878
rect 1942 811 1976 850
rect 2006 1050 2040 1089
rect 2006 1022 2009 1050
rect 2037 1022 2040 1050
rect 2006 964 2040 1022
rect 2006 936 2009 964
rect 2037 936 2040 964
rect 2006 878 2040 936
rect 2006 850 2009 878
rect 2037 850 2040 878
rect 2006 811 2040 850
rect 2070 1050 2104 1089
rect 2070 1022 2073 1050
rect 2101 1022 2104 1050
rect 2070 964 2104 1022
rect 2070 936 2073 964
rect 2101 936 2104 964
rect 2070 878 2104 936
rect 2070 850 2073 878
rect 2101 850 2104 878
rect 2070 811 2104 850
rect 2134 1050 2168 1089
rect 2134 1022 2137 1050
rect 2165 1022 2168 1050
rect 2134 964 2168 1022
rect 2134 936 2137 964
rect 2165 936 2168 964
rect 2134 878 2168 936
rect 2134 850 2137 878
rect 2165 850 2168 878
rect 2134 811 2168 850
rect 2198 1050 2232 1089
rect 2198 1022 2201 1050
rect 2229 1022 2232 1050
rect 2198 964 2232 1022
rect 2198 936 2201 964
rect 2229 936 2232 964
rect 2198 878 2232 936
rect 2198 850 2201 878
rect 2229 850 2232 878
rect 2198 811 2232 850
rect 2262 1050 2296 1089
rect 2262 1022 2265 1050
rect 2293 1022 2296 1050
rect 2262 964 2296 1022
rect 2262 936 2265 964
rect 2293 936 2296 964
rect 2262 878 2296 936
rect 2262 850 2265 878
rect 2293 850 2296 878
rect 2262 811 2296 850
rect 2326 1050 2360 1089
rect 2326 1022 2329 1050
rect 2357 1022 2360 1050
rect 2326 964 2360 1022
rect 2326 936 2329 964
rect 2357 936 2360 964
rect 2326 878 2360 936
rect 2326 850 2329 878
rect 2357 850 2360 878
rect 2326 811 2360 850
rect 2390 1050 2424 1089
rect 2390 1022 2393 1050
rect 2421 1022 2424 1050
rect 2390 964 2424 1022
rect 2390 936 2393 964
rect 2421 936 2424 964
rect 2390 878 2424 936
rect 2390 850 2393 878
rect 2421 850 2424 878
rect 2390 811 2424 850
rect 2454 1050 2488 1089
rect 2454 1022 2457 1050
rect 2485 1022 2488 1050
rect 2454 964 2488 1022
rect 2454 936 2457 964
rect 2485 936 2488 964
rect 2454 878 2488 936
rect 2454 850 2457 878
rect 2485 850 2488 878
rect 2454 811 2488 850
rect 2518 1050 2552 1089
rect 2518 1022 2521 1050
rect 2549 1022 2552 1050
rect 2518 964 2552 1022
rect 2518 936 2521 964
rect 2549 936 2552 964
rect 2518 878 2552 936
rect 2518 850 2521 878
rect 2549 850 2552 878
rect 2518 811 2552 850
rect 2584 1050 2618 1089
rect 2584 1022 2587 1050
rect 2615 1022 2618 1050
rect 2584 964 2618 1022
rect 2584 936 2587 964
rect 2615 936 2618 964
rect 2584 878 2618 936
rect 2584 850 2587 878
rect 2615 850 2618 878
rect 2584 811 2618 850
rect 2648 1050 2682 1089
rect 2648 1022 2651 1050
rect 2679 1022 2682 1050
rect 2648 964 2682 1022
rect 2648 936 2651 964
rect 2679 936 2682 964
rect 2648 878 2682 936
rect 2648 850 2651 878
rect 2679 850 2682 878
rect 2648 811 2682 850
rect 2712 1050 2746 1089
rect 2712 1022 2715 1050
rect 2743 1022 2746 1050
rect 2712 964 2746 1022
rect 2712 936 2715 964
rect 2743 936 2746 964
rect 2712 878 2746 936
rect 2712 850 2715 878
rect 2743 850 2746 878
rect 2712 811 2746 850
rect 2776 1050 2810 1089
rect 2776 1022 2779 1050
rect 2807 1022 2810 1050
rect 2776 964 2810 1022
rect 2776 936 2779 964
rect 2807 936 2810 964
rect 2776 878 2810 936
rect 2776 850 2779 878
rect 2807 850 2810 878
rect 2776 811 2810 850
rect 2840 1050 2874 1089
rect 2840 1022 2843 1050
rect 2871 1022 2874 1050
rect 2840 964 2874 1022
rect 2840 936 2843 964
rect 2871 936 2874 964
rect 2840 878 2874 936
rect 2840 850 2843 878
rect 2871 850 2874 878
rect 2840 811 2874 850
rect 2904 1050 2938 1089
rect 2904 1022 2907 1050
rect 2935 1022 2938 1050
rect 2904 964 2938 1022
rect 2904 936 2907 964
rect 2935 936 2938 964
rect 2904 878 2938 936
rect 2904 850 2907 878
rect 2935 850 2938 878
rect 2904 811 2938 850
rect 2968 1050 3002 1089
rect 2968 1022 2971 1050
rect 2999 1022 3002 1050
rect 2968 964 3002 1022
rect 2968 936 2971 964
rect 2999 936 3002 964
rect 2968 878 3002 936
rect 2968 850 2971 878
rect 2999 850 3002 878
rect 2968 811 3002 850
rect 3032 1050 3066 1089
rect 3032 1022 3035 1050
rect 3063 1022 3066 1050
rect 3032 964 3066 1022
rect 3032 936 3035 964
rect 3063 936 3066 964
rect 3032 878 3066 936
rect 3032 850 3035 878
rect 3063 850 3066 878
rect 3032 811 3066 850
rect 3096 1050 3130 1089
rect 3096 1022 3099 1050
rect 3127 1022 3130 1050
rect 3096 964 3130 1022
rect 3096 936 3099 964
rect 3127 936 3130 964
rect 3096 878 3130 936
rect 3096 850 3099 878
rect 3127 850 3130 878
rect 3096 811 3130 850
rect 3160 1050 3194 1089
rect 3160 1022 3163 1050
rect 3191 1022 3194 1050
rect 3160 964 3194 1022
rect 3160 936 3163 964
rect 3191 936 3194 964
rect 3160 878 3194 936
rect 3160 850 3163 878
rect 3191 850 3194 878
rect 3160 811 3194 850
rect 3226 1050 3260 1089
rect 3226 1022 3229 1050
rect 3257 1022 3260 1050
rect 3226 964 3260 1022
rect 3226 936 3229 964
rect 3257 936 3260 964
rect 3226 878 3260 936
rect 3226 850 3229 878
rect 3257 850 3260 878
rect 3226 811 3260 850
rect 3290 1050 3324 1089
rect 3290 1022 3293 1050
rect 3321 1022 3324 1050
rect 3290 964 3324 1022
rect 3290 936 3293 964
rect 3321 936 3324 964
rect 3290 878 3324 936
rect 3290 850 3293 878
rect 3321 850 3324 878
rect 3290 811 3324 850
rect 3354 1050 3388 1089
rect 3354 1022 3357 1050
rect 3385 1022 3388 1050
rect 3354 964 3388 1022
rect 3354 936 3357 964
rect 3385 936 3388 964
rect 3354 878 3388 936
rect 3354 850 3357 878
rect 3385 850 3388 878
rect 3354 811 3388 850
rect 3418 1050 3452 1089
rect 3418 1022 3421 1050
rect 3449 1022 3452 1050
rect 3418 964 3452 1022
rect 3418 936 3421 964
rect 3449 936 3452 964
rect 3418 878 3452 936
rect 3418 850 3421 878
rect 3449 850 3452 878
rect 3418 811 3452 850
rect 3482 1050 3516 1089
rect 3482 1022 3485 1050
rect 3513 1022 3516 1050
rect 3482 964 3516 1022
rect 3482 936 3485 964
rect 3513 936 3516 964
rect 3482 878 3516 936
rect 3482 850 3485 878
rect 3513 850 3516 878
rect 3482 811 3516 850
rect 3546 1050 3580 1089
rect 3546 1022 3549 1050
rect 3577 1022 3580 1050
rect 3546 964 3580 1022
rect 3546 936 3549 964
rect 3577 936 3580 964
rect 3546 878 3580 936
rect 3546 850 3549 878
rect 3577 850 3580 878
rect 3546 811 3580 850
rect 3610 1050 3644 1089
rect 3610 1022 3613 1050
rect 3641 1022 3644 1050
rect 3610 964 3644 1022
rect 3610 936 3613 964
rect 3641 936 3644 964
rect 3610 878 3644 936
rect 3610 850 3613 878
rect 3641 850 3644 878
rect 3610 811 3644 850
rect 3674 1050 3708 1089
rect 3674 1022 3677 1050
rect 3705 1022 3708 1050
rect 3674 964 3708 1022
rect 3674 936 3677 964
rect 3705 936 3708 964
rect 3674 878 3708 936
rect 3674 850 3677 878
rect 3705 850 3708 878
rect 3674 811 3708 850
rect 3738 1050 3772 1089
rect 3738 1022 3741 1050
rect 3769 1022 3772 1050
rect 3738 964 3772 1022
rect 3738 936 3741 964
rect 3769 936 3772 964
rect 3738 878 3772 936
rect 3738 850 3741 878
rect 3769 850 3772 878
rect 3738 811 3772 850
rect 3802 1050 3836 1089
rect 3802 1022 3805 1050
rect 3833 1022 3836 1050
rect 3802 964 3836 1022
rect 3802 936 3805 964
rect 3833 936 3836 964
rect 3802 878 3836 936
rect 3802 850 3805 878
rect 3833 850 3836 878
rect 3802 811 3836 850
rect 3868 1050 3902 1089
rect 3868 1022 3871 1050
rect 3899 1022 3902 1050
rect 3868 964 3902 1022
rect 3868 936 3871 964
rect 3899 936 3902 964
rect 3868 878 3902 936
rect 3868 850 3871 878
rect 3899 850 3902 878
rect 3868 811 3902 850
rect 3932 1050 3966 1089
rect 3932 1022 3935 1050
rect 3963 1022 3966 1050
rect 3932 964 3966 1022
rect 3932 936 3935 964
rect 3963 936 3966 964
rect 3932 878 3966 936
rect 3932 850 3935 878
rect 3963 850 3966 878
rect 3932 811 3966 850
rect 3996 1050 4030 1089
rect 3996 1022 3999 1050
rect 4027 1022 4030 1050
rect 3996 964 4030 1022
rect 3996 936 3999 964
rect 4027 936 4030 964
rect 3996 878 4030 936
rect 3996 850 3999 878
rect 4027 850 4030 878
rect 3996 811 4030 850
rect 4060 1050 4094 1089
rect 4060 1022 4063 1050
rect 4091 1022 4094 1050
rect 4060 964 4094 1022
rect 4060 936 4063 964
rect 4091 936 4094 964
rect 4060 878 4094 936
rect 4060 850 4063 878
rect 4091 850 4094 878
rect 4060 811 4094 850
rect 4124 1050 4158 1089
rect 4124 1022 4127 1050
rect 4155 1022 4158 1050
rect 4124 964 4158 1022
rect 4124 936 4127 964
rect 4155 936 4158 964
rect 4124 878 4158 936
rect 4124 850 4127 878
rect 4155 850 4158 878
rect 4124 811 4158 850
rect 4188 1050 4222 1089
rect 4188 1022 4191 1050
rect 4219 1022 4222 1050
rect 4188 964 4222 1022
rect 4188 936 4191 964
rect 4219 936 4222 964
rect 4188 878 4222 936
rect 4188 850 4191 878
rect 4219 850 4222 878
rect 4188 811 4222 850
rect 4252 1050 4286 1089
rect 4252 1022 4255 1050
rect 4283 1022 4286 1050
rect 4252 964 4286 1022
rect 4252 936 4255 964
rect 4283 936 4286 964
rect 4252 878 4286 936
rect 4252 850 4255 878
rect 4283 850 4286 878
rect 4252 811 4286 850
rect 4316 1050 4350 1089
rect 4316 1022 4319 1050
rect 4347 1022 4350 1050
rect 4316 964 4350 1022
rect 4316 936 4319 964
rect 4347 936 4350 964
rect 4316 878 4350 936
rect 4316 850 4319 878
rect 4347 850 4350 878
rect 4316 811 4350 850
rect 4380 1050 4414 1089
rect 4380 1022 4383 1050
rect 4411 1022 4414 1050
rect 4380 964 4414 1022
rect 4380 936 4383 964
rect 4411 936 4414 964
rect 4380 878 4414 936
rect 4380 850 4383 878
rect 4411 850 4414 878
rect 4380 811 4414 850
rect 4444 1050 4478 1089
rect 4444 1022 4447 1050
rect 4475 1022 4478 1050
rect 4444 964 4478 1022
rect 4444 936 4447 964
rect 4475 936 4478 964
rect 4444 878 4478 936
rect 4444 850 4447 878
rect 4475 850 4478 878
rect 4444 811 4478 850
rect 4510 1050 4544 1089
rect 4510 1022 4513 1050
rect 4541 1022 4544 1050
rect 4510 964 4544 1022
rect 4510 936 4513 964
rect 4541 936 4544 964
rect 4510 878 4544 936
rect 4510 850 4513 878
rect 4541 850 4544 878
rect 4510 811 4544 850
rect 4574 1050 4608 1089
rect 4574 1022 4577 1050
rect 4605 1022 4608 1050
rect 4574 964 4608 1022
rect 4574 936 4577 964
rect 4605 936 4608 964
rect 4574 878 4608 936
rect 4574 850 4577 878
rect 4605 850 4608 878
rect 4574 811 4608 850
rect 4638 1050 4672 1089
rect 4638 1022 4641 1050
rect 4669 1022 4672 1050
rect 4638 964 4672 1022
rect 4638 936 4641 964
rect 4669 936 4672 964
rect 4638 878 4672 936
rect 4638 850 4641 878
rect 4669 850 4672 878
rect 4638 811 4672 850
rect 4702 1050 4736 1089
rect 4702 1022 4705 1050
rect 4733 1022 4736 1050
rect 4702 964 4736 1022
rect 4702 936 4705 964
rect 4733 936 4736 964
rect 4702 878 4736 936
rect 4702 850 4705 878
rect 4733 850 4736 878
rect 4702 811 4736 850
rect 4766 1050 4800 1089
rect 4766 1022 4769 1050
rect 4797 1022 4800 1050
rect 4766 964 4800 1022
rect 4766 936 4769 964
rect 4797 936 4800 964
rect 4766 878 4800 936
rect 4766 850 4769 878
rect 4797 850 4800 878
rect 4766 811 4800 850
rect 4830 1050 4864 1089
rect 4830 1022 4833 1050
rect 4861 1022 4864 1050
rect 4830 964 4864 1022
rect 4830 936 4833 964
rect 4861 936 4864 964
rect 4830 878 4864 936
rect 4830 850 4833 878
rect 4861 850 4864 878
rect 4830 811 4864 850
rect 4894 1050 4928 1089
rect 4894 1022 4897 1050
rect 4925 1022 4928 1050
rect 4894 964 4928 1022
rect 4894 936 4897 964
rect 4925 936 4928 964
rect 4894 878 4928 936
rect 4894 850 4897 878
rect 4925 850 4928 878
rect 4894 811 4928 850
rect 4958 1050 4992 1089
rect 4958 1022 4961 1050
rect 4989 1022 4992 1050
rect 4958 964 4992 1022
rect 4958 936 4961 964
rect 4989 936 4992 964
rect 4958 878 4992 936
rect 4958 850 4961 878
rect 4989 850 4992 878
rect 4958 811 4992 850
rect 5022 1050 5056 1089
rect 5022 1022 5025 1050
rect 5053 1022 5056 1050
rect 5022 964 5056 1022
rect 5022 936 5025 964
rect 5053 936 5056 964
rect 5022 878 5056 936
rect 5022 850 5025 878
rect 5053 850 5056 878
rect 5022 811 5056 850
rect 5086 1050 5120 1089
rect 5086 1022 5089 1050
rect 5117 1022 5120 1050
rect 5086 964 5120 1022
rect 5086 936 5089 964
rect 5117 936 5120 964
rect 5086 878 5120 936
rect 5086 850 5089 878
rect 5117 850 5120 878
rect 5086 811 5120 850
rect 5152 1050 5186 1089
rect 5152 1022 5155 1050
rect 5183 1022 5186 1050
rect 5152 964 5186 1022
rect 5152 936 5155 964
rect 5183 936 5186 964
rect 5152 878 5186 936
rect 5152 850 5155 878
rect 5183 850 5186 878
rect 5152 811 5186 850
rect 5216 1050 5250 1089
rect 5216 1022 5219 1050
rect 5247 1022 5250 1050
rect 5216 964 5250 1022
rect 5216 936 5219 964
rect 5247 936 5250 964
rect 5216 878 5250 936
rect 5216 850 5219 878
rect 5247 850 5250 878
rect 5216 811 5250 850
rect 5280 1050 5314 1089
rect 5280 1022 5283 1050
rect 5311 1022 5314 1050
rect 5280 964 5314 1022
rect 5280 936 5283 964
rect 5311 936 5314 964
rect 5280 878 5314 936
rect 5280 850 5283 878
rect 5311 850 5314 878
rect 5280 811 5314 850
rect 5344 1050 5378 1089
rect 5344 1022 5347 1050
rect 5375 1022 5378 1050
rect 5344 964 5378 1022
rect 5344 936 5347 964
rect 5375 936 5378 964
rect 5344 878 5378 936
rect 5344 850 5347 878
rect 5375 850 5378 878
rect 5344 811 5378 850
rect 5408 1050 5442 1089
rect 5408 1022 5411 1050
rect 5439 1022 5442 1050
rect 5408 964 5442 1022
rect 5408 936 5411 964
rect 5439 936 5442 964
rect 5408 878 5442 936
rect 5408 850 5411 878
rect 5439 850 5442 878
rect 5408 811 5442 850
rect 5472 1050 5506 1089
rect 5472 1022 5475 1050
rect 5503 1022 5506 1050
rect 5472 964 5506 1022
rect 5472 936 5475 964
rect 5503 936 5506 964
rect 5472 878 5506 936
rect 5472 850 5475 878
rect 5503 850 5506 878
rect 5472 811 5506 850
rect 5536 1050 5570 1089
rect 5536 1022 5539 1050
rect 5567 1022 5570 1050
rect 5536 964 5570 1022
rect 5536 936 5539 964
rect 5567 936 5570 964
rect 5536 878 5570 936
rect 5536 850 5539 878
rect 5567 850 5570 878
rect 5536 811 5570 850
rect 5600 1050 5634 1089
rect 5600 1022 5603 1050
rect 5631 1022 5634 1050
rect 5600 964 5634 1022
rect 5600 936 5603 964
rect 5631 936 5634 964
rect 5600 878 5634 936
rect 5600 850 5603 878
rect 5631 850 5634 878
rect 5600 811 5634 850
rect 5664 1050 5698 1089
rect 5664 1022 5667 1050
rect 5695 1022 5698 1050
rect 5664 964 5698 1022
rect 5664 936 5667 964
rect 5695 936 5698 964
rect 5664 878 5698 936
rect 5664 850 5667 878
rect 5695 850 5698 878
rect 5664 811 5698 850
rect 5728 1050 5762 1089
rect 5728 1022 5731 1050
rect 5759 1022 5762 1050
rect 5728 964 5762 1022
rect 5728 936 5731 964
rect 5759 936 5762 964
rect 5728 878 5762 936
rect 5728 850 5731 878
rect 5759 850 5762 878
rect 5728 811 5762 850
rect 5794 1050 5828 1089
rect 5794 1022 5797 1050
rect 5825 1022 5828 1050
rect 5794 964 5828 1022
rect 5794 936 5797 964
rect 5825 936 5828 964
rect 5794 878 5828 936
rect 5794 850 5797 878
rect 5825 850 5828 878
rect 5794 811 5828 850
rect 5858 1050 5892 1089
rect 5858 1022 5861 1050
rect 5889 1022 5892 1050
rect 5858 964 5892 1022
rect 5858 936 5861 964
rect 5889 936 5892 964
rect 5858 878 5892 936
rect 5858 850 5861 878
rect 5889 850 5892 878
rect 5858 811 5892 850
rect 5922 1050 5956 1089
rect 5922 1022 5925 1050
rect 5953 1022 5956 1050
rect 5922 964 5956 1022
rect 5922 936 5925 964
rect 5953 936 5956 964
rect 5922 878 5956 936
rect 5922 850 5925 878
rect 5953 850 5956 878
rect 5922 811 5956 850
rect 5986 1050 6020 1089
rect 5986 1022 5989 1050
rect 6017 1022 6020 1050
rect 5986 964 6020 1022
rect 5986 936 5989 964
rect 6017 936 6020 964
rect 5986 878 6020 936
rect 5986 850 5989 878
rect 6017 850 6020 878
rect 5986 811 6020 850
rect 6050 1050 6084 1089
rect 6050 1022 6053 1050
rect 6081 1022 6084 1050
rect 6050 964 6084 1022
rect 6050 936 6053 964
rect 6081 936 6084 964
rect 6050 878 6084 936
rect 6050 850 6053 878
rect 6081 850 6084 878
rect 6050 811 6084 850
rect 6114 1050 6148 1089
rect 6114 1022 6117 1050
rect 6145 1022 6148 1050
rect 6114 964 6148 1022
rect 6114 936 6117 964
rect 6145 936 6148 964
rect 6114 878 6148 936
rect 6114 850 6117 878
rect 6145 850 6148 878
rect 6114 811 6148 850
rect 6178 1050 6212 1089
rect 6178 1022 6181 1050
rect 6209 1022 6212 1050
rect 6178 964 6212 1022
rect 6178 936 6181 964
rect 6209 936 6212 964
rect 6178 878 6212 936
rect 6178 850 6181 878
rect 6209 850 6212 878
rect 6178 811 6212 850
rect 6242 1050 6276 1089
rect 6242 1022 6245 1050
rect 6273 1022 6276 1050
rect 6242 964 6276 1022
rect 6242 936 6245 964
rect 6273 936 6276 964
rect 6242 878 6276 936
rect 6242 850 6245 878
rect 6273 850 6276 878
rect 6242 811 6276 850
rect 6306 1050 6340 1089
rect 6306 1022 6309 1050
rect 6337 1022 6340 1050
rect 6306 964 6340 1022
rect 6306 936 6309 964
rect 6337 936 6340 964
rect 6306 878 6340 936
rect 6306 850 6309 878
rect 6337 850 6340 878
rect 6306 811 6340 850
rect 6370 1050 6404 1089
rect 6370 1022 6373 1050
rect 6401 1022 6404 1050
rect 6370 964 6404 1022
rect 6370 936 6373 964
rect 6401 936 6404 964
rect 6370 878 6404 936
rect 6370 850 6373 878
rect 6401 850 6404 878
rect 6370 811 6404 850
rect 6436 1050 6470 1089
rect 6436 1022 6439 1050
rect 6467 1022 6470 1050
rect 6436 964 6470 1022
rect 6436 936 6439 964
rect 6467 936 6470 964
rect 6436 878 6470 936
rect 6436 850 6439 878
rect 6467 850 6470 878
rect 6436 811 6470 850
rect 6500 1050 6534 1089
rect 6500 1022 6503 1050
rect 6531 1022 6534 1050
rect 6500 964 6534 1022
rect 6500 936 6503 964
rect 6531 936 6534 964
rect 6500 878 6534 936
rect 6500 850 6503 878
rect 6531 850 6534 878
rect 6500 811 6534 850
rect 6564 1050 6598 1089
rect 6564 1022 6567 1050
rect 6595 1022 6598 1050
rect 6564 964 6598 1022
rect 6564 936 6567 964
rect 6595 936 6598 964
rect 6564 878 6598 936
rect 6564 850 6567 878
rect 6595 850 6598 878
rect 6564 811 6598 850
rect 6628 1050 6662 1089
rect 6628 1022 6631 1050
rect 6659 1022 6662 1050
rect 6628 964 6662 1022
rect 6628 936 6631 964
rect 6659 936 6662 964
rect 6628 878 6662 936
rect 6628 850 6631 878
rect 6659 850 6662 878
rect 6628 811 6662 850
rect 6692 1050 6726 1089
rect 6692 1022 6695 1050
rect 6723 1022 6726 1050
rect 6692 964 6726 1022
rect 6692 936 6695 964
rect 6723 936 6726 964
rect 6692 878 6726 936
rect 6692 850 6695 878
rect 6723 850 6726 878
rect 6692 811 6726 850
rect 6756 1050 6790 1089
rect 6756 1022 6759 1050
rect 6787 1022 6790 1050
rect 6756 964 6790 1022
rect 6756 936 6759 964
rect 6787 936 6790 964
rect 6756 878 6790 936
rect 6756 850 6759 878
rect 6787 850 6790 878
rect 6756 811 6790 850
rect 6820 1050 6854 1089
rect 6820 1022 6823 1050
rect 6851 1022 6854 1050
rect 6820 964 6854 1022
rect 6820 936 6823 964
rect 6851 936 6854 964
rect 6820 878 6854 936
rect 6820 850 6823 878
rect 6851 850 6854 878
rect 6820 811 6854 850
rect 6884 1050 6918 1089
rect 6884 1022 6887 1050
rect 6915 1022 6918 1050
rect 6884 964 6918 1022
rect 6884 936 6887 964
rect 6915 936 6918 964
rect 6884 878 6918 936
rect 6884 850 6887 878
rect 6915 850 6918 878
rect 6884 811 6918 850
rect 6948 1050 6982 1089
rect 6948 1022 6951 1050
rect 6979 1022 6982 1050
rect 6948 964 6982 1022
rect 6948 936 6951 964
rect 6979 936 6982 964
rect 6948 878 6982 936
rect 6948 850 6951 878
rect 6979 850 6982 878
rect 6948 811 6982 850
rect 7012 1050 7046 1089
rect 7012 1022 7015 1050
rect 7043 1022 7046 1050
rect 7012 964 7046 1022
rect 7012 936 7015 964
rect 7043 936 7046 964
rect 7012 878 7046 936
rect 7012 850 7015 878
rect 7043 850 7046 878
rect 7012 811 7046 850
rect 7078 1050 7112 1089
rect 7078 1022 7081 1050
rect 7109 1022 7112 1050
rect 7078 964 7112 1022
rect 7078 936 7081 964
rect 7109 936 7112 964
rect 7078 878 7112 936
rect 7078 850 7081 878
rect 7109 850 7112 878
rect 7078 811 7112 850
rect 7142 1050 7176 1089
rect 7142 1022 7145 1050
rect 7173 1022 7176 1050
rect 7142 964 7176 1022
rect 7142 936 7145 964
rect 7173 936 7176 964
rect 7142 878 7176 936
rect 7142 850 7145 878
rect 7173 850 7176 878
rect 7142 811 7176 850
rect 7206 1050 7240 1089
rect 7206 1022 7209 1050
rect 7237 1022 7240 1050
rect 7206 964 7240 1022
rect 7206 936 7209 964
rect 7237 936 7240 964
rect 7206 878 7240 936
rect 7206 850 7209 878
rect 7237 850 7240 878
rect 7206 811 7240 850
rect 7270 1050 7304 1089
rect 7270 1022 7273 1050
rect 7301 1022 7304 1050
rect 7270 964 7304 1022
rect 7270 936 7273 964
rect 7301 936 7304 964
rect 7270 878 7304 936
rect 7270 850 7273 878
rect 7301 850 7304 878
rect 7270 811 7304 850
rect 7334 1050 7368 1089
rect 7334 1022 7337 1050
rect 7365 1022 7368 1050
rect 7334 964 7368 1022
rect 7334 936 7337 964
rect 7365 936 7368 964
rect 7334 878 7368 936
rect 7334 850 7337 878
rect 7365 850 7368 878
rect 7334 811 7368 850
rect 7398 1050 7432 1089
rect 7398 1022 7401 1050
rect 7429 1022 7432 1050
rect 7398 964 7432 1022
rect 7398 936 7401 964
rect 7429 936 7432 964
rect 7398 878 7432 936
rect 7398 850 7401 878
rect 7429 850 7432 878
rect 7398 811 7432 850
rect 7462 1050 7496 1089
rect 7462 1022 7465 1050
rect 7493 1022 7496 1050
rect 7462 964 7496 1022
rect 7462 936 7465 964
rect 7493 936 7496 964
rect 7462 878 7496 936
rect 7462 850 7465 878
rect 7493 850 7496 878
rect 7462 811 7496 850
rect 7526 1050 7560 1089
rect 7526 1022 7529 1050
rect 7557 1022 7560 1050
rect 7526 964 7560 1022
rect 7526 936 7529 964
rect 7557 936 7560 964
rect 7526 878 7560 936
rect 7526 850 7529 878
rect 7557 850 7560 878
rect 7526 811 7560 850
rect 7590 1050 7624 1089
rect 7590 1022 7593 1050
rect 7621 1022 7624 1050
rect 7590 964 7624 1022
rect 7590 936 7593 964
rect 7621 936 7624 964
rect 7590 878 7624 936
rect 7590 850 7593 878
rect 7621 850 7624 878
rect 7590 811 7624 850
rect 7654 1050 7688 1089
rect 7654 1022 7657 1050
rect 7685 1022 7688 1050
rect 7654 964 7688 1022
rect 7654 936 7657 964
rect 7685 936 7688 964
rect 7654 878 7688 936
rect 7654 850 7657 878
rect 7685 850 7688 878
rect 7654 811 7688 850
rect 7720 1050 7754 1089
rect 7720 1022 7723 1050
rect 7751 1022 7754 1050
rect 7720 964 7754 1022
rect 7720 936 7723 964
rect 7751 936 7754 964
rect 7720 878 7754 936
rect 7720 850 7723 878
rect 7751 850 7754 878
rect 7720 811 7754 850
rect 7784 1050 7818 1089
rect 7784 1022 7787 1050
rect 7815 1022 7818 1050
rect 7784 964 7818 1022
rect 7784 936 7787 964
rect 7815 936 7818 964
rect 7784 878 7818 936
rect 7784 850 7787 878
rect 7815 850 7818 878
rect 7784 811 7818 850
rect 7848 1050 7882 1089
rect 7848 1022 7851 1050
rect 7879 1022 7882 1050
rect 7848 964 7882 1022
rect 7848 936 7851 964
rect 7879 936 7882 964
rect 7848 878 7882 936
rect 7848 850 7851 878
rect 7879 850 7882 878
rect 7848 811 7882 850
rect 7912 1050 7946 1089
rect 7912 1022 7915 1050
rect 7943 1022 7946 1050
rect 7912 964 7946 1022
rect 7912 936 7915 964
rect 7943 936 7946 964
rect 7912 878 7946 936
rect 7912 850 7915 878
rect 7943 850 7946 878
rect 7912 811 7946 850
rect 7976 1050 8010 1089
rect 7976 1022 7979 1050
rect 8007 1022 8010 1050
rect 7976 964 8010 1022
rect 7976 936 7979 964
rect 8007 936 8010 964
rect 7976 878 8010 936
rect 7976 850 7979 878
rect 8007 850 8010 878
rect 7976 811 8010 850
rect 8040 1050 8074 1089
rect 8040 1022 8043 1050
rect 8071 1022 8074 1050
rect 8040 964 8074 1022
rect 8040 936 8043 964
rect 8071 936 8074 964
rect 8040 878 8074 936
rect 8040 850 8043 878
rect 8071 850 8074 878
rect 8040 811 8074 850
rect 8104 1050 8138 1089
rect 8104 1022 8107 1050
rect 8135 1022 8138 1050
rect 8104 964 8138 1022
rect 8104 936 8107 964
rect 8135 936 8138 964
rect 8104 878 8138 936
rect 8104 850 8107 878
rect 8135 850 8138 878
rect 8104 811 8138 850
rect 8168 1050 8202 1089
rect 8168 1022 8171 1050
rect 8199 1022 8202 1050
rect 8168 964 8202 1022
rect 8168 936 8171 964
rect 8199 936 8202 964
rect 8168 878 8202 936
rect 8168 850 8171 878
rect 8199 850 8202 878
rect 8168 811 8202 850
rect 8232 1050 8266 1089
rect 8232 1022 8235 1050
rect 8263 1022 8266 1050
rect 8232 964 8266 1022
rect 8232 936 8235 964
rect 8263 936 8266 964
rect 8232 878 8266 936
rect 8232 850 8235 878
rect 8263 850 8266 878
rect 8232 811 8266 850
rect 8296 1050 8330 1089
rect 8296 1022 8299 1050
rect 8327 1022 8330 1050
rect 8296 964 8330 1022
rect 8296 936 8299 964
rect 8327 936 8330 964
rect 8296 878 8330 936
rect 8296 850 8299 878
rect 8327 850 8330 878
rect 8296 811 8330 850
rect 8362 1050 8396 1089
rect 8362 1022 8365 1050
rect 8393 1022 8396 1050
rect 8362 964 8396 1022
rect 8362 936 8365 964
rect 8393 936 8396 964
rect 8362 878 8396 936
rect 8362 850 8365 878
rect 8393 850 8396 878
rect 8362 811 8396 850
rect 8426 1050 8460 1089
rect 8426 1022 8429 1050
rect 8457 1022 8460 1050
rect 8426 964 8460 1022
rect 8426 936 8429 964
rect 8457 936 8460 964
rect 8426 878 8460 936
rect 8426 850 8429 878
rect 8457 850 8460 878
rect 8426 811 8460 850
rect 8490 1050 8524 1089
rect 8490 1022 8493 1050
rect 8521 1022 8524 1050
rect 8490 964 8524 1022
rect 8490 936 8493 964
rect 8521 936 8524 964
rect 8490 878 8524 936
rect 8490 850 8493 878
rect 8521 850 8524 878
rect 8490 811 8524 850
rect 8554 1050 8588 1089
rect 8554 1022 8557 1050
rect 8585 1022 8588 1050
rect 8554 964 8588 1022
rect 8554 936 8557 964
rect 8585 936 8588 964
rect 8554 878 8588 936
rect 8554 850 8557 878
rect 8585 850 8588 878
rect 8554 811 8588 850
rect 8618 1050 8652 1089
rect 8618 1022 8621 1050
rect 8649 1022 8652 1050
rect 8618 964 8652 1022
rect 8618 936 8621 964
rect 8649 936 8652 964
rect 8618 878 8652 936
rect 8618 850 8621 878
rect 8649 850 8652 878
rect 8618 811 8652 850
rect 8682 1050 8716 1089
rect 8682 1022 8685 1050
rect 8713 1022 8716 1050
rect 8682 964 8716 1022
rect 8682 936 8685 964
rect 8713 936 8716 964
rect 8682 878 8716 936
rect 8682 850 8685 878
rect 8713 850 8716 878
rect 8682 811 8716 850
rect 8746 1050 8780 1089
rect 8746 1022 8749 1050
rect 8777 1022 8780 1050
rect 8746 964 8780 1022
rect 8746 936 8749 964
rect 8777 936 8780 964
rect 8746 878 8780 936
rect 8746 850 8749 878
rect 8777 850 8780 878
rect 8746 811 8780 850
rect 8810 1050 8844 1089
rect 8810 1022 8813 1050
rect 8841 1022 8844 1050
rect 8810 964 8844 1022
rect 8810 936 8813 964
rect 8841 936 8844 964
rect 8810 878 8844 936
rect 8810 850 8813 878
rect 8841 850 8844 878
rect 8810 811 8844 850
rect 8874 1050 8908 1089
rect 8874 1022 8877 1050
rect 8905 1022 8908 1050
rect 8874 964 8908 1022
rect 8874 936 8877 964
rect 8905 936 8908 964
rect 8874 878 8908 936
rect 8874 850 8877 878
rect 8905 850 8908 878
rect 8874 811 8908 850
rect 8938 1050 8972 1089
rect 8938 1022 8941 1050
rect 8969 1022 8972 1050
rect 8938 964 8972 1022
rect 8938 936 8941 964
rect 8969 936 8972 964
rect 8938 878 8972 936
rect 8938 850 8941 878
rect 8969 850 8972 878
rect 8938 811 8972 850
rect 9004 1050 9038 1089
rect 9004 1022 9007 1050
rect 9035 1022 9038 1050
rect 9004 964 9038 1022
rect 9004 936 9007 964
rect 9035 936 9038 964
rect 9004 878 9038 936
rect 9004 850 9007 878
rect 9035 850 9038 878
rect 9004 811 9038 850
rect 9068 1050 9102 1089
rect 9068 1022 9071 1050
rect 9099 1022 9102 1050
rect 9068 964 9102 1022
rect 9068 936 9071 964
rect 9099 936 9102 964
rect 9068 878 9102 936
rect 9068 850 9071 878
rect 9099 850 9102 878
rect 9068 811 9102 850
rect 9132 1050 9166 1089
rect 9132 1022 9135 1050
rect 9163 1022 9166 1050
rect 9132 964 9166 1022
rect 9132 936 9135 964
rect 9163 936 9166 964
rect 9132 878 9166 936
rect 9132 850 9135 878
rect 9163 850 9166 878
rect 9132 811 9166 850
rect 9196 1050 9230 1089
rect 9196 1022 9199 1050
rect 9227 1022 9230 1050
rect 9196 964 9230 1022
rect 9196 936 9199 964
rect 9227 936 9230 964
rect 9196 878 9230 936
rect 9196 850 9199 878
rect 9227 850 9230 878
rect 9196 811 9230 850
rect 9260 1050 9294 1089
rect 9260 1022 9263 1050
rect 9291 1022 9294 1050
rect 9260 964 9294 1022
rect 9260 936 9263 964
rect 9291 936 9294 964
rect 9260 878 9294 936
rect 9260 850 9263 878
rect 9291 850 9294 878
rect 9260 811 9294 850
rect 9324 1050 9358 1089
rect 9324 1022 9327 1050
rect 9355 1022 9358 1050
rect 9324 964 9358 1022
rect 9324 936 9327 964
rect 9355 936 9358 964
rect 9324 878 9358 936
rect 9324 850 9327 878
rect 9355 850 9358 878
rect 9324 811 9358 850
rect 9388 1050 9422 1089
rect 9388 1022 9391 1050
rect 9419 1022 9422 1050
rect 9388 964 9422 1022
rect 9388 936 9391 964
rect 9419 936 9422 964
rect 9388 878 9422 936
rect 9388 850 9391 878
rect 9419 850 9422 878
rect 9388 811 9422 850
rect 9452 1050 9486 1089
rect 9452 1022 9455 1050
rect 9483 1022 9486 1050
rect 9452 964 9486 1022
rect 9452 936 9455 964
rect 9483 936 9486 964
rect 9452 878 9486 936
rect 9452 850 9455 878
rect 9483 850 9486 878
rect 9452 811 9486 850
rect 9516 1050 9550 1089
rect 9516 1022 9519 1050
rect 9547 1022 9550 1050
rect 9516 964 9550 1022
rect 9516 936 9519 964
rect 9547 936 9550 964
rect 9516 878 9550 936
rect 9516 850 9519 878
rect 9547 850 9550 878
rect 9516 811 9550 850
rect 9580 1050 9614 1089
rect 9580 1022 9583 1050
rect 9611 1022 9614 1050
rect 9580 964 9614 1022
rect 9580 936 9583 964
rect 9611 936 9614 964
rect 9580 878 9614 936
rect 9580 850 9583 878
rect 9611 850 9614 878
rect 9580 811 9614 850
rect 9646 1050 9680 1089
rect 9646 1022 9649 1050
rect 9677 1022 9680 1050
rect 9646 964 9680 1022
rect 9646 936 9649 964
rect 9677 936 9680 964
rect 9646 878 9680 936
rect 9646 850 9649 878
rect 9677 850 9680 878
rect 9646 811 9680 850
rect 9710 1050 9744 1089
rect 9710 1022 9713 1050
rect 9741 1022 9744 1050
rect 9710 964 9744 1022
rect 9710 936 9713 964
rect 9741 936 9744 964
rect 9710 878 9744 936
rect 9710 850 9713 878
rect 9741 850 9744 878
rect 9710 811 9744 850
rect 9774 1050 9808 1089
rect 9774 1022 9777 1050
rect 9805 1022 9808 1050
rect 9774 964 9808 1022
rect 9774 936 9777 964
rect 9805 936 9808 964
rect 9774 878 9808 936
rect 9774 850 9777 878
rect 9805 850 9808 878
rect 9774 811 9808 850
rect 9838 1050 9872 1089
rect 9838 1022 9841 1050
rect 9869 1022 9872 1050
rect 9838 964 9872 1022
rect 9838 936 9841 964
rect 9869 936 9872 964
rect 9838 878 9872 936
rect 9838 850 9841 878
rect 9869 850 9872 878
rect 9838 811 9872 850
rect 9902 1050 9936 1089
rect 9902 1022 9905 1050
rect 9933 1022 9936 1050
rect 9902 964 9936 1022
rect 9902 936 9905 964
rect 9933 936 9936 964
rect 9902 878 9936 936
rect 9902 850 9905 878
rect 9933 850 9936 878
rect 9902 811 9936 850
rect 9966 1050 10000 1089
rect 9966 1022 9969 1050
rect 9997 1022 10000 1050
rect 9966 964 10000 1022
rect 9966 936 9969 964
rect 9997 936 10000 964
rect 9966 878 10000 936
rect 9966 850 9969 878
rect 9997 850 10000 878
rect 9966 811 10000 850
rect 10030 1050 10064 1089
rect 10030 1022 10033 1050
rect 10061 1022 10064 1050
rect 10030 964 10064 1022
rect 10030 936 10033 964
rect 10061 936 10064 964
rect 10030 878 10064 936
rect 10030 850 10033 878
rect 10061 850 10064 878
rect 10030 811 10064 850
rect 10094 1050 10128 1089
rect 10094 1022 10097 1050
rect 10125 1022 10128 1050
rect 10094 964 10128 1022
rect 10094 936 10097 964
rect 10125 936 10128 964
rect 10094 878 10128 936
rect 10094 850 10097 878
rect 10125 850 10128 878
rect 10094 811 10128 850
rect 10158 1050 10192 1089
rect 10158 1022 10161 1050
rect 10189 1022 10192 1050
rect 10158 964 10192 1022
rect 10158 936 10161 964
rect 10189 936 10192 964
rect 10158 878 10192 936
rect 10158 850 10161 878
rect 10189 850 10192 878
rect 10158 811 10192 850
rect 10222 1050 10256 1089
rect 10222 1022 10225 1050
rect 10253 1022 10256 1050
rect 10222 964 10256 1022
rect 10222 936 10225 964
rect 10253 936 10256 964
rect 10222 878 10256 936
rect 10222 850 10225 878
rect 10253 850 10256 878
rect 10222 811 10256 850
rect 10288 1050 10322 1089
rect 10288 1022 10291 1050
rect 10319 1022 10322 1050
rect 10288 964 10322 1022
rect 10288 936 10291 964
rect 10319 936 10322 964
rect 10288 878 10322 936
rect 10288 850 10291 878
rect 10319 850 10322 878
rect 10288 811 10322 850
rect 10352 1050 10386 1089
rect 10352 1022 10355 1050
rect 10383 1022 10386 1050
rect 10352 964 10386 1022
rect 10352 936 10355 964
rect 10383 936 10386 964
rect 10352 878 10386 936
rect 10352 850 10355 878
rect 10383 850 10386 878
rect 10352 811 10386 850
rect 10416 1050 10450 1089
rect 10416 1022 10419 1050
rect 10447 1022 10450 1050
rect 10416 964 10450 1022
rect 10416 936 10419 964
rect 10447 936 10450 964
rect 10416 878 10450 936
rect 10416 850 10419 878
rect 10447 850 10450 878
rect 10416 811 10450 850
rect 10480 1050 10514 1089
rect 10480 1022 10483 1050
rect 10511 1022 10514 1050
rect 10480 964 10514 1022
rect 10480 936 10483 964
rect 10511 936 10514 964
rect 10480 878 10514 936
rect 10480 850 10483 878
rect 10511 850 10514 878
rect 10480 811 10514 850
rect 10544 1050 10578 1089
rect 10544 1022 10547 1050
rect 10575 1022 10578 1050
rect 10544 964 10578 1022
rect 10544 936 10547 964
rect 10575 936 10578 964
rect 10544 878 10578 936
rect 10544 850 10547 878
rect 10575 850 10578 878
rect 10544 811 10578 850
rect 10608 1050 10642 1089
rect 10608 1022 10611 1050
rect 10639 1022 10642 1050
rect 10608 964 10642 1022
rect 10608 936 10611 964
rect 10639 936 10642 964
rect 10608 878 10642 936
rect 10608 850 10611 878
rect 10639 850 10642 878
rect 10608 811 10642 850
rect 10672 1050 10706 1089
rect 10672 1022 10675 1050
rect 10703 1022 10706 1050
rect 10672 964 10706 1022
rect 10672 936 10675 964
rect 10703 936 10706 964
rect 10672 878 10706 936
rect 10672 850 10675 878
rect 10703 850 10706 878
rect 10672 811 10706 850
rect 10736 1050 10770 1089
rect 10736 1022 10739 1050
rect 10767 1022 10770 1050
rect 10736 964 10770 1022
rect 10736 936 10739 964
rect 10767 936 10770 964
rect 10736 878 10770 936
rect 10736 850 10739 878
rect 10767 850 10770 878
rect 10736 811 10770 850
rect 10800 1050 10834 1089
rect 10800 1022 10803 1050
rect 10831 1022 10834 1050
rect 10800 964 10834 1022
rect 10800 936 10803 964
rect 10831 936 10834 964
rect 10800 878 10834 936
rect 10800 850 10803 878
rect 10831 850 10834 878
rect 10800 811 10834 850
rect 10864 1050 10898 1089
rect 10864 1022 10867 1050
rect 10895 1022 10898 1050
rect 10864 964 10898 1022
rect 10864 936 10867 964
rect 10895 936 10898 964
rect 10864 878 10898 936
rect 10864 850 10867 878
rect 10895 850 10898 878
rect 10864 811 10898 850
rect 10930 1050 10964 1089
rect 10930 1022 10933 1050
rect 10961 1022 10964 1050
rect 10930 964 10964 1022
rect 10930 936 10933 964
rect 10961 936 10964 964
rect 10930 878 10964 936
rect 10930 850 10933 878
rect 10961 850 10964 878
rect 10930 811 10964 850
rect 10994 1050 11028 1089
rect 10994 1022 10997 1050
rect 11025 1022 11028 1050
rect 10994 964 11028 1022
rect 10994 936 10997 964
rect 11025 936 11028 964
rect 10994 878 11028 936
rect 10994 850 10997 878
rect 11025 850 11028 878
rect 10994 811 11028 850
rect 11058 1050 11092 1089
rect 11058 1022 11061 1050
rect 11089 1022 11092 1050
rect 11058 964 11092 1022
rect 11058 936 11061 964
rect 11089 936 11092 964
rect 11058 878 11092 936
rect 11058 850 11061 878
rect 11089 850 11092 878
rect 11058 811 11092 850
rect 11122 1050 11156 1089
rect 11122 1022 11125 1050
rect 11153 1022 11156 1050
rect 11122 964 11156 1022
rect 11122 936 11125 964
rect 11153 936 11156 964
rect 11122 878 11156 936
rect 11122 850 11125 878
rect 11153 850 11156 878
rect 11122 811 11156 850
rect 11186 1050 11220 1089
rect 11186 1022 11189 1050
rect 11217 1022 11220 1050
rect 11186 964 11220 1022
rect 11186 936 11189 964
rect 11217 936 11220 964
rect 11186 878 11220 936
rect 11186 850 11189 878
rect 11217 850 11220 878
rect 11186 811 11220 850
rect 11250 1050 11284 1089
rect 11250 1022 11253 1050
rect 11281 1022 11284 1050
rect 11250 964 11284 1022
rect 11250 936 11253 964
rect 11281 936 11284 964
rect 11250 878 11284 936
rect 11250 850 11253 878
rect 11281 850 11284 878
rect 11250 811 11284 850
rect 11314 1050 11348 1089
rect 11314 1022 11317 1050
rect 11345 1022 11348 1050
rect 11314 964 11348 1022
rect 11314 936 11317 964
rect 11345 936 11348 964
rect 11314 878 11348 936
rect 11314 850 11317 878
rect 11345 850 11348 878
rect 11314 811 11348 850
rect 11378 1050 11412 1089
rect 11378 1022 11381 1050
rect 11409 1022 11412 1050
rect 11378 964 11412 1022
rect 11378 936 11381 964
rect 11409 936 11412 964
rect 11378 878 11412 936
rect 11378 850 11381 878
rect 11409 850 11412 878
rect 11378 811 11412 850
rect 11442 1050 11476 1089
rect 11442 1022 11445 1050
rect 11473 1022 11476 1050
rect 11442 964 11476 1022
rect 11442 936 11445 964
rect 11473 936 11476 964
rect 11442 878 11476 936
rect 11442 850 11445 878
rect 11473 850 11476 878
rect 11442 811 11476 850
rect 11506 1050 11540 1089
rect 11506 1022 11509 1050
rect 11537 1022 11540 1050
rect 11506 964 11540 1022
rect 11506 936 11509 964
rect 11537 936 11540 964
rect 11506 878 11540 936
rect 11506 850 11509 878
rect 11537 850 11540 878
rect 11506 811 11540 850
rect 11572 1050 11606 1089
rect 11572 1022 11575 1050
rect 11603 1022 11606 1050
rect 11572 964 11606 1022
rect 11572 936 11575 964
rect 11603 936 11606 964
rect 11572 878 11606 936
rect 11572 850 11575 878
rect 11603 850 11606 878
rect 11572 811 11606 850
rect 11636 1050 11670 1089
rect 11636 1022 11639 1050
rect 11667 1022 11670 1050
rect 11636 964 11670 1022
rect 11636 936 11639 964
rect 11667 936 11670 964
rect 11636 878 11670 936
rect 11636 850 11639 878
rect 11667 850 11670 878
rect 11636 811 11670 850
rect 11700 1050 11734 1089
rect 11700 1022 11703 1050
rect 11731 1022 11734 1050
rect 11700 964 11734 1022
rect 11700 936 11703 964
rect 11731 936 11734 964
rect 11700 878 11734 936
rect 11700 850 11703 878
rect 11731 850 11734 878
rect 11700 811 11734 850
rect 11764 1050 11798 1089
rect 11764 1022 11767 1050
rect 11795 1022 11798 1050
rect 11764 964 11798 1022
rect 11764 936 11767 964
rect 11795 936 11798 964
rect 11764 878 11798 936
rect 11764 850 11767 878
rect 11795 850 11798 878
rect 11764 811 11798 850
rect 11828 1050 11862 1089
rect 11828 1022 11831 1050
rect 11859 1022 11862 1050
rect 11828 964 11862 1022
rect 11828 936 11831 964
rect 11859 936 11862 964
rect 11828 878 11862 936
rect 11828 850 11831 878
rect 11859 850 11862 878
rect 11828 811 11862 850
rect 11892 1050 11926 1089
rect 11892 1022 11895 1050
rect 11923 1022 11926 1050
rect 11892 964 11926 1022
rect 11892 936 11895 964
rect 11923 936 11926 964
rect 11892 878 11926 936
rect 11892 850 11895 878
rect 11923 850 11926 878
rect 11892 811 11926 850
rect 11956 1050 11990 1089
rect 11956 1022 11959 1050
rect 11987 1022 11990 1050
rect 11956 964 11990 1022
rect 11956 936 11959 964
rect 11987 936 11990 964
rect 11956 878 11990 936
rect 11956 850 11959 878
rect 11987 850 11990 878
rect 11956 811 11990 850
rect 12020 1050 12054 1089
rect 12020 1022 12023 1050
rect 12051 1022 12054 1050
rect 12020 964 12054 1022
rect 12020 936 12023 964
rect 12051 936 12054 964
rect 12020 878 12054 936
rect 12020 850 12023 878
rect 12051 850 12054 878
rect 12020 811 12054 850
rect 12084 1050 12118 1089
rect 12084 1022 12087 1050
rect 12115 1022 12118 1050
rect 12084 964 12118 1022
rect 12084 936 12087 964
rect 12115 936 12118 964
rect 12084 878 12118 936
rect 12084 850 12087 878
rect 12115 850 12118 878
rect 12084 811 12118 850
rect 12148 1050 12182 1089
rect 12148 1022 12151 1050
rect 12179 1022 12182 1050
rect 12148 964 12182 1022
rect 12148 936 12151 964
rect 12179 936 12182 964
rect 12148 878 12182 936
rect 12148 850 12151 878
rect 12179 850 12182 878
rect 12148 811 12182 850
rect 12214 1050 12248 1089
rect 12214 1022 12217 1050
rect 12245 1022 12248 1050
rect 12214 964 12248 1022
rect 12214 936 12217 964
rect 12245 936 12248 964
rect 12214 878 12248 936
rect 12214 850 12217 878
rect 12245 850 12248 878
rect 12214 811 12248 850
rect 12278 1050 12312 1089
rect 12278 1022 12281 1050
rect 12309 1022 12312 1050
rect 12278 964 12312 1022
rect 12278 936 12281 964
rect 12309 936 12312 964
rect 12278 878 12312 936
rect 12278 850 12281 878
rect 12309 850 12312 878
rect 12278 811 12312 850
rect 12342 1050 12376 1089
rect 12342 1022 12345 1050
rect 12373 1022 12376 1050
rect 12342 964 12376 1022
rect 12342 936 12345 964
rect 12373 936 12376 964
rect 12342 878 12376 936
rect 12342 850 12345 878
rect 12373 850 12376 878
rect 12342 811 12376 850
rect 12406 1050 12440 1089
rect 12406 1022 12409 1050
rect 12437 1022 12440 1050
rect 12406 964 12440 1022
rect 12406 936 12409 964
rect 12437 936 12440 964
rect 12406 878 12440 936
rect 12406 850 12409 878
rect 12437 850 12440 878
rect 12406 811 12440 850
rect 12470 1050 12504 1089
rect 12470 1022 12473 1050
rect 12501 1022 12504 1050
rect 12470 964 12504 1022
rect 12470 936 12473 964
rect 12501 936 12504 964
rect 12470 878 12504 936
rect 12470 850 12473 878
rect 12501 850 12504 878
rect 12470 811 12504 850
rect 12534 1050 12568 1089
rect 12534 1022 12537 1050
rect 12565 1022 12568 1050
rect 12534 964 12568 1022
rect 12534 936 12537 964
rect 12565 936 12568 964
rect 12534 878 12568 936
rect 12534 850 12537 878
rect 12565 850 12568 878
rect 12534 811 12568 850
rect 12598 1050 12632 1089
rect 12598 1022 12601 1050
rect 12629 1022 12632 1050
rect 12598 964 12632 1022
rect 12598 936 12601 964
rect 12629 936 12632 964
rect 12598 878 12632 936
rect 12598 850 12601 878
rect 12629 850 12632 878
rect 12598 811 12632 850
rect 12662 1050 12696 1089
rect 12662 1022 12665 1050
rect 12693 1022 12696 1050
rect 12662 964 12696 1022
rect 12662 936 12665 964
rect 12693 936 12696 964
rect 12662 878 12696 936
rect 12662 850 12665 878
rect 12693 850 12696 878
rect 12662 811 12696 850
rect 12726 1050 12760 1089
rect 12726 1022 12729 1050
rect 12757 1022 12760 1050
rect 12726 964 12760 1022
rect 12726 936 12729 964
rect 12757 936 12760 964
rect 12726 878 12760 936
rect 12726 850 12729 878
rect 12757 850 12760 878
rect 12726 811 12760 850
rect 12790 1050 12824 1089
rect 12790 1022 12793 1050
rect 12821 1022 12824 1050
rect 12790 964 12824 1022
rect 12790 936 12793 964
rect 12821 936 12824 964
rect 12790 878 12824 936
rect 12790 850 12793 878
rect 12821 850 12824 878
rect 12790 811 12824 850
rect 16 670 50 709
rect 16 642 19 670
rect 47 642 50 670
rect 16 584 50 642
rect 16 556 19 584
rect 47 556 50 584
rect 16 498 50 556
rect 16 470 19 498
rect 47 470 50 498
rect 16 431 50 470
rect 80 670 114 709
rect 80 642 83 670
rect 111 642 114 670
rect 80 584 114 642
rect 80 556 83 584
rect 111 556 114 584
rect 80 498 114 556
rect 80 470 83 498
rect 111 470 114 498
rect 80 431 114 470
rect 144 670 178 709
rect 144 642 147 670
rect 175 642 178 670
rect 144 584 178 642
rect 144 556 147 584
rect 175 556 178 584
rect 144 498 178 556
rect 144 470 147 498
rect 175 470 178 498
rect 144 431 178 470
rect 208 670 242 709
rect 208 642 211 670
rect 239 642 242 670
rect 208 584 242 642
rect 208 556 211 584
rect 239 556 242 584
rect 208 498 242 556
rect 208 470 211 498
rect 239 470 242 498
rect 208 431 242 470
rect 272 670 306 709
rect 272 642 275 670
rect 303 642 306 670
rect 272 584 306 642
rect 272 556 275 584
rect 303 556 306 584
rect 272 498 306 556
rect 272 470 275 498
rect 303 470 306 498
rect 272 431 306 470
rect 336 670 370 709
rect 336 642 339 670
rect 367 642 370 670
rect 336 584 370 642
rect 336 556 339 584
rect 367 556 370 584
rect 336 498 370 556
rect 336 470 339 498
rect 367 470 370 498
rect 336 431 370 470
rect 400 670 434 709
rect 400 642 403 670
rect 431 642 434 670
rect 400 584 434 642
rect 400 556 403 584
rect 431 556 434 584
rect 400 498 434 556
rect 400 470 403 498
rect 431 470 434 498
rect 400 431 434 470
rect 464 670 498 709
rect 464 642 467 670
rect 495 642 498 670
rect 464 584 498 642
rect 464 556 467 584
rect 495 556 498 584
rect 464 498 498 556
rect 464 470 467 498
rect 495 470 498 498
rect 464 431 498 470
rect 528 670 562 709
rect 528 642 531 670
rect 559 642 562 670
rect 528 584 562 642
rect 528 556 531 584
rect 559 556 562 584
rect 528 498 562 556
rect 528 470 531 498
rect 559 470 562 498
rect 528 431 562 470
rect 592 670 626 709
rect 592 642 595 670
rect 623 642 626 670
rect 592 584 626 642
rect 592 556 595 584
rect 623 556 626 584
rect 592 498 626 556
rect 592 470 595 498
rect 623 470 626 498
rect 592 431 626 470
rect 658 670 692 709
rect 658 642 661 670
rect 689 642 692 670
rect 658 584 692 642
rect 658 556 661 584
rect 689 556 692 584
rect 658 498 692 556
rect 658 470 661 498
rect 689 470 692 498
rect 658 431 692 470
rect 722 670 756 709
rect 722 642 725 670
rect 753 642 756 670
rect 722 584 756 642
rect 722 556 725 584
rect 753 556 756 584
rect 722 498 756 556
rect 722 470 725 498
rect 753 470 756 498
rect 722 431 756 470
rect 786 670 820 709
rect 786 642 789 670
rect 817 642 820 670
rect 786 584 820 642
rect 786 556 789 584
rect 817 556 820 584
rect 786 498 820 556
rect 786 470 789 498
rect 817 470 820 498
rect 786 431 820 470
rect 850 670 884 709
rect 850 642 853 670
rect 881 642 884 670
rect 850 584 884 642
rect 850 556 853 584
rect 881 556 884 584
rect 850 498 884 556
rect 850 470 853 498
rect 881 470 884 498
rect 850 431 884 470
rect 914 670 948 709
rect 914 642 917 670
rect 945 642 948 670
rect 914 584 948 642
rect 914 556 917 584
rect 945 556 948 584
rect 914 498 948 556
rect 914 470 917 498
rect 945 470 948 498
rect 914 431 948 470
rect 978 670 1012 709
rect 978 642 981 670
rect 1009 642 1012 670
rect 978 584 1012 642
rect 978 556 981 584
rect 1009 556 1012 584
rect 978 498 1012 556
rect 978 470 981 498
rect 1009 470 1012 498
rect 978 431 1012 470
rect 1042 670 1076 709
rect 1042 642 1045 670
rect 1073 642 1076 670
rect 1042 584 1076 642
rect 1042 556 1045 584
rect 1073 556 1076 584
rect 1042 498 1076 556
rect 1042 470 1045 498
rect 1073 470 1076 498
rect 1042 431 1076 470
rect 1106 670 1140 709
rect 1106 642 1109 670
rect 1137 642 1140 670
rect 1106 584 1140 642
rect 1106 556 1109 584
rect 1137 556 1140 584
rect 1106 498 1140 556
rect 1106 470 1109 498
rect 1137 470 1140 498
rect 1106 431 1140 470
rect 1170 670 1204 709
rect 1170 642 1173 670
rect 1201 642 1204 670
rect 1170 584 1204 642
rect 1170 556 1173 584
rect 1201 556 1204 584
rect 1170 498 1204 556
rect 1170 470 1173 498
rect 1201 470 1204 498
rect 1170 431 1204 470
rect 1234 670 1268 709
rect 1234 642 1237 670
rect 1265 642 1268 670
rect 1234 584 1268 642
rect 1234 556 1237 584
rect 1265 556 1268 584
rect 1234 498 1268 556
rect 1234 470 1237 498
rect 1265 470 1268 498
rect 1234 431 1268 470
rect 1300 670 1334 709
rect 1300 642 1303 670
rect 1331 642 1334 670
rect 1300 584 1334 642
rect 1300 556 1303 584
rect 1331 556 1334 584
rect 1300 498 1334 556
rect 1300 470 1303 498
rect 1331 470 1334 498
rect 1300 431 1334 470
rect 1364 670 1398 709
rect 1364 642 1367 670
rect 1395 642 1398 670
rect 1364 584 1398 642
rect 1364 556 1367 584
rect 1395 556 1398 584
rect 1364 498 1398 556
rect 1364 470 1367 498
rect 1395 470 1398 498
rect 1364 431 1398 470
rect 1428 670 1462 709
rect 1428 642 1431 670
rect 1459 642 1462 670
rect 1428 584 1462 642
rect 1428 556 1431 584
rect 1459 556 1462 584
rect 1428 498 1462 556
rect 1428 470 1431 498
rect 1459 470 1462 498
rect 1428 431 1462 470
rect 1492 670 1526 709
rect 1492 642 1495 670
rect 1523 642 1526 670
rect 1492 584 1526 642
rect 1492 556 1495 584
rect 1523 556 1526 584
rect 1492 498 1526 556
rect 1492 470 1495 498
rect 1523 470 1526 498
rect 1492 431 1526 470
rect 1556 670 1590 709
rect 1556 642 1559 670
rect 1587 642 1590 670
rect 1556 584 1590 642
rect 1556 556 1559 584
rect 1587 556 1590 584
rect 1556 498 1590 556
rect 1556 470 1559 498
rect 1587 470 1590 498
rect 1556 431 1590 470
rect 1620 670 1654 709
rect 1620 642 1623 670
rect 1651 642 1654 670
rect 1620 584 1654 642
rect 1620 556 1623 584
rect 1651 556 1654 584
rect 1620 498 1654 556
rect 1620 470 1623 498
rect 1651 470 1654 498
rect 1620 431 1654 470
rect 1684 670 1718 709
rect 1684 642 1687 670
rect 1715 642 1718 670
rect 1684 584 1718 642
rect 1684 556 1687 584
rect 1715 556 1718 584
rect 1684 498 1718 556
rect 1684 470 1687 498
rect 1715 470 1718 498
rect 1684 431 1718 470
rect 1748 670 1782 709
rect 1748 642 1751 670
rect 1779 642 1782 670
rect 1748 584 1782 642
rect 1748 556 1751 584
rect 1779 556 1782 584
rect 1748 498 1782 556
rect 1748 470 1751 498
rect 1779 470 1782 498
rect 1748 431 1782 470
rect 1812 670 1846 709
rect 1812 642 1815 670
rect 1843 642 1846 670
rect 1812 584 1846 642
rect 1812 556 1815 584
rect 1843 556 1846 584
rect 1812 498 1846 556
rect 1812 470 1815 498
rect 1843 470 1846 498
rect 1812 431 1846 470
rect 1876 670 1910 709
rect 1876 642 1879 670
rect 1907 642 1910 670
rect 1876 584 1910 642
rect 1876 556 1879 584
rect 1907 556 1910 584
rect 1876 498 1910 556
rect 1876 470 1879 498
rect 1907 470 1910 498
rect 1876 431 1910 470
rect 1942 670 1976 709
rect 1942 642 1945 670
rect 1973 642 1976 670
rect 1942 584 1976 642
rect 1942 556 1945 584
rect 1973 556 1976 584
rect 1942 498 1976 556
rect 1942 470 1945 498
rect 1973 470 1976 498
rect 1942 431 1976 470
rect 2006 670 2040 709
rect 2006 642 2009 670
rect 2037 642 2040 670
rect 2006 584 2040 642
rect 2006 556 2009 584
rect 2037 556 2040 584
rect 2006 498 2040 556
rect 2006 470 2009 498
rect 2037 470 2040 498
rect 2006 431 2040 470
rect 2070 670 2104 709
rect 2070 642 2073 670
rect 2101 642 2104 670
rect 2070 584 2104 642
rect 2070 556 2073 584
rect 2101 556 2104 584
rect 2070 498 2104 556
rect 2070 470 2073 498
rect 2101 470 2104 498
rect 2070 431 2104 470
rect 2134 670 2168 709
rect 2134 642 2137 670
rect 2165 642 2168 670
rect 2134 584 2168 642
rect 2134 556 2137 584
rect 2165 556 2168 584
rect 2134 498 2168 556
rect 2134 470 2137 498
rect 2165 470 2168 498
rect 2134 431 2168 470
rect 2198 670 2232 709
rect 2198 642 2201 670
rect 2229 642 2232 670
rect 2198 584 2232 642
rect 2198 556 2201 584
rect 2229 556 2232 584
rect 2198 498 2232 556
rect 2198 470 2201 498
rect 2229 470 2232 498
rect 2198 431 2232 470
rect 2262 670 2296 709
rect 2262 642 2265 670
rect 2293 642 2296 670
rect 2262 584 2296 642
rect 2262 556 2265 584
rect 2293 556 2296 584
rect 2262 498 2296 556
rect 2262 470 2265 498
rect 2293 470 2296 498
rect 2262 431 2296 470
rect 2326 670 2360 709
rect 2326 642 2329 670
rect 2357 642 2360 670
rect 2326 584 2360 642
rect 2326 556 2329 584
rect 2357 556 2360 584
rect 2326 498 2360 556
rect 2326 470 2329 498
rect 2357 470 2360 498
rect 2326 431 2360 470
rect 2390 670 2424 709
rect 2390 642 2393 670
rect 2421 642 2424 670
rect 2390 584 2424 642
rect 2390 556 2393 584
rect 2421 556 2424 584
rect 2390 498 2424 556
rect 2390 470 2393 498
rect 2421 470 2424 498
rect 2390 431 2424 470
rect 2454 670 2488 709
rect 2454 642 2457 670
rect 2485 642 2488 670
rect 2454 584 2488 642
rect 2454 556 2457 584
rect 2485 556 2488 584
rect 2454 498 2488 556
rect 2454 470 2457 498
rect 2485 470 2488 498
rect 2454 431 2488 470
rect 2518 670 2552 709
rect 2518 642 2521 670
rect 2549 642 2552 670
rect 2518 584 2552 642
rect 2518 556 2521 584
rect 2549 556 2552 584
rect 2518 498 2552 556
rect 2518 470 2521 498
rect 2549 470 2552 498
rect 2518 431 2552 470
rect 2584 670 2618 709
rect 2584 642 2587 670
rect 2615 642 2618 670
rect 2584 584 2618 642
rect 2584 556 2587 584
rect 2615 556 2618 584
rect 2584 498 2618 556
rect 2584 470 2587 498
rect 2615 470 2618 498
rect 2584 431 2618 470
rect 2648 670 2682 709
rect 2648 642 2651 670
rect 2679 642 2682 670
rect 2648 584 2682 642
rect 2648 556 2651 584
rect 2679 556 2682 584
rect 2648 498 2682 556
rect 2648 470 2651 498
rect 2679 470 2682 498
rect 2648 431 2682 470
rect 2712 670 2746 709
rect 2712 642 2715 670
rect 2743 642 2746 670
rect 2712 584 2746 642
rect 2712 556 2715 584
rect 2743 556 2746 584
rect 2712 498 2746 556
rect 2712 470 2715 498
rect 2743 470 2746 498
rect 2712 431 2746 470
rect 2776 670 2810 709
rect 2776 642 2779 670
rect 2807 642 2810 670
rect 2776 584 2810 642
rect 2776 556 2779 584
rect 2807 556 2810 584
rect 2776 498 2810 556
rect 2776 470 2779 498
rect 2807 470 2810 498
rect 2776 431 2810 470
rect 2840 670 2874 709
rect 2840 642 2843 670
rect 2871 642 2874 670
rect 2840 584 2874 642
rect 2840 556 2843 584
rect 2871 556 2874 584
rect 2840 498 2874 556
rect 2840 470 2843 498
rect 2871 470 2874 498
rect 2840 431 2874 470
rect 2904 670 2938 709
rect 2904 642 2907 670
rect 2935 642 2938 670
rect 2904 584 2938 642
rect 2904 556 2907 584
rect 2935 556 2938 584
rect 2904 498 2938 556
rect 2904 470 2907 498
rect 2935 470 2938 498
rect 2904 431 2938 470
rect 2968 670 3002 709
rect 2968 642 2971 670
rect 2999 642 3002 670
rect 2968 584 3002 642
rect 2968 556 2971 584
rect 2999 556 3002 584
rect 2968 498 3002 556
rect 2968 470 2971 498
rect 2999 470 3002 498
rect 2968 431 3002 470
rect 3032 670 3066 709
rect 3032 642 3035 670
rect 3063 642 3066 670
rect 3032 584 3066 642
rect 3032 556 3035 584
rect 3063 556 3066 584
rect 3032 498 3066 556
rect 3032 470 3035 498
rect 3063 470 3066 498
rect 3032 431 3066 470
rect 3096 670 3130 709
rect 3096 642 3099 670
rect 3127 642 3130 670
rect 3096 584 3130 642
rect 3096 556 3099 584
rect 3127 556 3130 584
rect 3096 498 3130 556
rect 3096 470 3099 498
rect 3127 470 3130 498
rect 3096 431 3130 470
rect 3160 670 3194 709
rect 3160 642 3163 670
rect 3191 642 3194 670
rect 3160 584 3194 642
rect 3160 556 3163 584
rect 3191 556 3194 584
rect 3160 498 3194 556
rect 3160 470 3163 498
rect 3191 470 3194 498
rect 3160 431 3194 470
rect 3226 670 3260 709
rect 3226 642 3229 670
rect 3257 642 3260 670
rect 3226 584 3260 642
rect 3226 556 3229 584
rect 3257 556 3260 584
rect 3226 498 3260 556
rect 3226 470 3229 498
rect 3257 470 3260 498
rect 3226 431 3260 470
rect 3290 670 3324 709
rect 3290 642 3293 670
rect 3321 642 3324 670
rect 3290 584 3324 642
rect 3290 556 3293 584
rect 3321 556 3324 584
rect 3290 498 3324 556
rect 3290 470 3293 498
rect 3321 470 3324 498
rect 3290 431 3324 470
rect 3354 670 3388 709
rect 3354 642 3357 670
rect 3385 642 3388 670
rect 3354 584 3388 642
rect 3354 556 3357 584
rect 3385 556 3388 584
rect 3354 498 3388 556
rect 3354 470 3357 498
rect 3385 470 3388 498
rect 3354 431 3388 470
rect 3418 670 3452 709
rect 3418 642 3421 670
rect 3449 642 3452 670
rect 3418 584 3452 642
rect 3418 556 3421 584
rect 3449 556 3452 584
rect 3418 498 3452 556
rect 3418 470 3421 498
rect 3449 470 3452 498
rect 3418 431 3452 470
rect 3482 670 3516 709
rect 3482 642 3485 670
rect 3513 642 3516 670
rect 3482 584 3516 642
rect 3482 556 3485 584
rect 3513 556 3516 584
rect 3482 498 3516 556
rect 3482 470 3485 498
rect 3513 470 3516 498
rect 3482 431 3516 470
rect 3546 670 3580 709
rect 3546 642 3549 670
rect 3577 642 3580 670
rect 3546 584 3580 642
rect 3546 556 3549 584
rect 3577 556 3580 584
rect 3546 498 3580 556
rect 3546 470 3549 498
rect 3577 470 3580 498
rect 3546 431 3580 470
rect 3610 670 3644 709
rect 3610 642 3613 670
rect 3641 642 3644 670
rect 3610 584 3644 642
rect 3610 556 3613 584
rect 3641 556 3644 584
rect 3610 498 3644 556
rect 3610 470 3613 498
rect 3641 470 3644 498
rect 3610 431 3644 470
rect 3674 670 3708 709
rect 3674 642 3677 670
rect 3705 642 3708 670
rect 3674 584 3708 642
rect 3674 556 3677 584
rect 3705 556 3708 584
rect 3674 498 3708 556
rect 3674 470 3677 498
rect 3705 470 3708 498
rect 3674 431 3708 470
rect 3738 670 3772 709
rect 3738 642 3741 670
rect 3769 642 3772 670
rect 3738 584 3772 642
rect 3738 556 3741 584
rect 3769 556 3772 584
rect 3738 498 3772 556
rect 3738 470 3741 498
rect 3769 470 3772 498
rect 3738 431 3772 470
rect 3802 670 3836 709
rect 3802 642 3805 670
rect 3833 642 3836 670
rect 3802 584 3836 642
rect 3802 556 3805 584
rect 3833 556 3836 584
rect 3802 498 3836 556
rect 3802 470 3805 498
rect 3833 470 3836 498
rect 3802 431 3836 470
rect 3868 670 3902 709
rect 3868 642 3871 670
rect 3899 642 3902 670
rect 3868 584 3902 642
rect 3868 556 3871 584
rect 3899 556 3902 584
rect 3868 498 3902 556
rect 3868 470 3871 498
rect 3899 470 3902 498
rect 3868 431 3902 470
rect 3932 670 3966 709
rect 3932 642 3935 670
rect 3963 642 3966 670
rect 3932 584 3966 642
rect 3932 556 3935 584
rect 3963 556 3966 584
rect 3932 498 3966 556
rect 3932 470 3935 498
rect 3963 470 3966 498
rect 3932 431 3966 470
rect 3996 670 4030 709
rect 3996 642 3999 670
rect 4027 642 4030 670
rect 3996 584 4030 642
rect 3996 556 3999 584
rect 4027 556 4030 584
rect 3996 498 4030 556
rect 3996 470 3999 498
rect 4027 470 4030 498
rect 3996 431 4030 470
rect 4060 670 4094 709
rect 4060 642 4063 670
rect 4091 642 4094 670
rect 4060 584 4094 642
rect 4060 556 4063 584
rect 4091 556 4094 584
rect 4060 498 4094 556
rect 4060 470 4063 498
rect 4091 470 4094 498
rect 4060 431 4094 470
rect 4124 670 4158 709
rect 4124 642 4127 670
rect 4155 642 4158 670
rect 4124 584 4158 642
rect 4124 556 4127 584
rect 4155 556 4158 584
rect 4124 498 4158 556
rect 4124 470 4127 498
rect 4155 470 4158 498
rect 4124 431 4158 470
rect 4188 670 4222 709
rect 4188 642 4191 670
rect 4219 642 4222 670
rect 4188 584 4222 642
rect 4188 556 4191 584
rect 4219 556 4222 584
rect 4188 498 4222 556
rect 4188 470 4191 498
rect 4219 470 4222 498
rect 4188 431 4222 470
rect 4252 670 4286 709
rect 4252 642 4255 670
rect 4283 642 4286 670
rect 4252 584 4286 642
rect 4252 556 4255 584
rect 4283 556 4286 584
rect 4252 498 4286 556
rect 4252 470 4255 498
rect 4283 470 4286 498
rect 4252 431 4286 470
rect 4316 670 4350 709
rect 4316 642 4319 670
rect 4347 642 4350 670
rect 4316 584 4350 642
rect 4316 556 4319 584
rect 4347 556 4350 584
rect 4316 498 4350 556
rect 4316 470 4319 498
rect 4347 470 4350 498
rect 4316 431 4350 470
rect 4380 670 4414 709
rect 4380 642 4383 670
rect 4411 642 4414 670
rect 4380 584 4414 642
rect 4380 556 4383 584
rect 4411 556 4414 584
rect 4380 498 4414 556
rect 4380 470 4383 498
rect 4411 470 4414 498
rect 4380 431 4414 470
rect 4444 670 4478 709
rect 4444 642 4447 670
rect 4475 642 4478 670
rect 4444 584 4478 642
rect 4444 556 4447 584
rect 4475 556 4478 584
rect 4444 498 4478 556
rect 4444 470 4447 498
rect 4475 470 4478 498
rect 4444 431 4478 470
rect 4510 670 4544 709
rect 4510 642 4513 670
rect 4541 642 4544 670
rect 4510 584 4544 642
rect 4510 556 4513 584
rect 4541 556 4544 584
rect 4510 498 4544 556
rect 4510 470 4513 498
rect 4541 470 4544 498
rect 4510 431 4544 470
rect 4574 670 4608 709
rect 4574 642 4577 670
rect 4605 642 4608 670
rect 4574 584 4608 642
rect 4574 556 4577 584
rect 4605 556 4608 584
rect 4574 498 4608 556
rect 4574 470 4577 498
rect 4605 470 4608 498
rect 4574 431 4608 470
rect 4638 670 4672 709
rect 4638 642 4641 670
rect 4669 642 4672 670
rect 4638 584 4672 642
rect 4638 556 4641 584
rect 4669 556 4672 584
rect 4638 498 4672 556
rect 4638 470 4641 498
rect 4669 470 4672 498
rect 4638 431 4672 470
rect 4702 670 4736 709
rect 4702 642 4705 670
rect 4733 642 4736 670
rect 4702 584 4736 642
rect 4702 556 4705 584
rect 4733 556 4736 584
rect 4702 498 4736 556
rect 4702 470 4705 498
rect 4733 470 4736 498
rect 4702 431 4736 470
rect 4766 670 4800 709
rect 4766 642 4769 670
rect 4797 642 4800 670
rect 4766 584 4800 642
rect 4766 556 4769 584
rect 4797 556 4800 584
rect 4766 498 4800 556
rect 4766 470 4769 498
rect 4797 470 4800 498
rect 4766 431 4800 470
rect 4830 670 4864 709
rect 4830 642 4833 670
rect 4861 642 4864 670
rect 4830 584 4864 642
rect 4830 556 4833 584
rect 4861 556 4864 584
rect 4830 498 4864 556
rect 4830 470 4833 498
rect 4861 470 4864 498
rect 4830 431 4864 470
rect 4894 670 4928 709
rect 4894 642 4897 670
rect 4925 642 4928 670
rect 4894 584 4928 642
rect 4894 556 4897 584
rect 4925 556 4928 584
rect 4894 498 4928 556
rect 4894 470 4897 498
rect 4925 470 4928 498
rect 4894 431 4928 470
rect 4958 670 4992 709
rect 4958 642 4961 670
rect 4989 642 4992 670
rect 4958 584 4992 642
rect 4958 556 4961 584
rect 4989 556 4992 584
rect 4958 498 4992 556
rect 4958 470 4961 498
rect 4989 470 4992 498
rect 4958 431 4992 470
rect 5022 670 5056 709
rect 5022 642 5025 670
rect 5053 642 5056 670
rect 5022 584 5056 642
rect 5022 556 5025 584
rect 5053 556 5056 584
rect 5022 498 5056 556
rect 5022 470 5025 498
rect 5053 470 5056 498
rect 5022 431 5056 470
rect 5086 670 5120 709
rect 5086 642 5089 670
rect 5117 642 5120 670
rect 5086 584 5120 642
rect 5086 556 5089 584
rect 5117 556 5120 584
rect 5086 498 5120 556
rect 5086 470 5089 498
rect 5117 470 5120 498
rect 5086 431 5120 470
rect 5152 670 5186 709
rect 5152 642 5155 670
rect 5183 642 5186 670
rect 5152 584 5186 642
rect 5152 556 5155 584
rect 5183 556 5186 584
rect 5152 498 5186 556
rect 5152 470 5155 498
rect 5183 470 5186 498
rect 5152 431 5186 470
rect 5216 670 5250 709
rect 5216 642 5219 670
rect 5247 642 5250 670
rect 5216 584 5250 642
rect 5216 556 5219 584
rect 5247 556 5250 584
rect 5216 498 5250 556
rect 5216 470 5219 498
rect 5247 470 5250 498
rect 5216 431 5250 470
rect 5280 670 5314 709
rect 5280 642 5283 670
rect 5311 642 5314 670
rect 5280 584 5314 642
rect 5280 556 5283 584
rect 5311 556 5314 584
rect 5280 498 5314 556
rect 5280 470 5283 498
rect 5311 470 5314 498
rect 5280 431 5314 470
rect 5344 670 5378 709
rect 5344 642 5347 670
rect 5375 642 5378 670
rect 5344 584 5378 642
rect 5344 556 5347 584
rect 5375 556 5378 584
rect 5344 498 5378 556
rect 5344 470 5347 498
rect 5375 470 5378 498
rect 5344 431 5378 470
rect 5408 670 5442 709
rect 5408 642 5411 670
rect 5439 642 5442 670
rect 5408 584 5442 642
rect 5408 556 5411 584
rect 5439 556 5442 584
rect 5408 498 5442 556
rect 5408 470 5411 498
rect 5439 470 5442 498
rect 5408 431 5442 470
rect 5472 670 5506 709
rect 5472 642 5475 670
rect 5503 642 5506 670
rect 5472 584 5506 642
rect 5472 556 5475 584
rect 5503 556 5506 584
rect 5472 498 5506 556
rect 5472 470 5475 498
rect 5503 470 5506 498
rect 5472 431 5506 470
rect 5536 670 5570 709
rect 5536 642 5539 670
rect 5567 642 5570 670
rect 5536 584 5570 642
rect 5536 556 5539 584
rect 5567 556 5570 584
rect 5536 498 5570 556
rect 5536 470 5539 498
rect 5567 470 5570 498
rect 5536 431 5570 470
rect 5600 670 5634 709
rect 5600 642 5603 670
rect 5631 642 5634 670
rect 5600 584 5634 642
rect 5600 556 5603 584
rect 5631 556 5634 584
rect 5600 498 5634 556
rect 5600 470 5603 498
rect 5631 470 5634 498
rect 5600 431 5634 470
rect 5664 670 5698 709
rect 5664 642 5667 670
rect 5695 642 5698 670
rect 5664 584 5698 642
rect 5664 556 5667 584
rect 5695 556 5698 584
rect 5664 498 5698 556
rect 5664 470 5667 498
rect 5695 470 5698 498
rect 5664 431 5698 470
rect 5728 670 5762 709
rect 5728 642 5731 670
rect 5759 642 5762 670
rect 5728 584 5762 642
rect 5728 556 5731 584
rect 5759 556 5762 584
rect 5728 498 5762 556
rect 5728 470 5731 498
rect 5759 470 5762 498
rect 5728 431 5762 470
rect 5794 670 5828 709
rect 5794 642 5797 670
rect 5825 642 5828 670
rect 5794 584 5828 642
rect 5794 556 5797 584
rect 5825 556 5828 584
rect 5794 498 5828 556
rect 5794 470 5797 498
rect 5825 470 5828 498
rect 5794 431 5828 470
rect 5858 670 5892 709
rect 5858 642 5861 670
rect 5889 642 5892 670
rect 5858 584 5892 642
rect 5858 556 5861 584
rect 5889 556 5892 584
rect 5858 498 5892 556
rect 5858 470 5861 498
rect 5889 470 5892 498
rect 5858 431 5892 470
rect 5922 670 5956 709
rect 5922 642 5925 670
rect 5953 642 5956 670
rect 5922 584 5956 642
rect 5922 556 5925 584
rect 5953 556 5956 584
rect 5922 498 5956 556
rect 5922 470 5925 498
rect 5953 470 5956 498
rect 5922 431 5956 470
rect 5986 670 6020 709
rect 5986 642 5989 670
rect 6017 642 6020 670
rect 5986 584 6020 642
rect 5986 556 5989 584
rect 6017 556 6020 584
rect 5986 498 6020 556
rect 5986 470 5989 498
rect 6017 470 6020 498
rect 5986 431 6020 470
rect 6050 670 6084 709
rect 6050 642 6053 670
rect 6081 642 6084 670
rect 6050 584 6084 642
rect 6050 556 6053 584
rect 6081 556 6084 584
rect 6050 498 6084 556
rect 6050 470 6053 498
rect 6081 470 6084 498
rect 6050 431 6084 470
rect 6114 670 6148 709
rect 6114 642 6117 670
rect 6145 642 6148 670
rect 6114 584 6148 642
rect 6114 556 6117 584
rect 6145 556 6148 584
rect 6114 498 6148 556
rect 6114 470 6117 498
rect 6145 470 6148 498
rect 6114 431 6148 470
rect 6178 670 6212 709
rect 6178 642 6181 670
rect 6209 642 6212 670
rect 6178 584 6212 642
rect 6178 556 6181 584
rect 6209 556 6212 584
rect 6178 498 6212 556
rect 6178 470 6181 498
rect 6209 470 6212 498
rect 6178 431 6212 470
rect 6242 670 6276 709
rect 6242 642 6245 670
rect 6273 642 6276 670
rect 6242 584 6276 642
rect 6242 556 6245 584
rect 6273 556 6276 584
rect 6242 498 6276 556
rect 6242 470 6245 498
rect 6273 470 6276 498
rect 6242 431 6276 470
rect 6306 670 6340 709
rect 6306 642 6309 670
rect 6337 642 6340 670
rect 6306 584 6340 642
rect 6306 556 6309 584
rect 6337 556 6340 584
rect 6306 498 6340 556
rect 6306 470 6309 498
rect 6337 470 6340 498
rect 6306 431 6340 470
rect 6370 670 6404 709
rect 6370 642 6373 670
rect 6401 642 6404 670
rect 6370 584 6404 642
rect 6370 556 6373 584
rect 6401 556 6404 584
rect 6370 498 6404 556
rect 6370 470 6373 498
rect 6401 470 6404 498
rect 6370 431 6404 470
rect 6436 670 6470 709
rect 6436 642 6439 670
rect 6467 642 6470 670
rect 6436 584 6470 642
rect 6436 556 6439 584
rect 6467 556 6470 584
rect 6436 498 6470 556
rect 6436 470 6439 498
rect 6467 470 6470 498
rect 6436 431 6470 470
rect 6500 670 6534 709
rect 6500 642 6503 670
rect 6531 642 6534 670
rect 6500 584 6534 642
rect 6500 556 6503 584
rect 6531 556 6534 584
rect 6500 498 6534 556
rect 6500 470 6503 498
rect 6531 470 6534 498
rect 6500 431 6534 470
rect 6564 670 6598 709
rect 6564 642 6567 670
rect 6595 642 6598 670
rect 6564 584 6598 642
rect 6564 556 6567 584
rect 6595 556 6598 584
rect 6564 498 6598 556
rect 6564 470 6567 498
rect 6595 470 6598 498
rect 6564 431 6598 470
rect 6628 670 6662 709
rect 6628 642 6631 670
rect 6659 642 6662 670
rect 6628 584 6662 642
rect 6628 556 6631 584
rect 6659 556 6662 584
rect 6628 498 6662 556
rect 6628 470 6631 498
rect 6659 470 6662 498
rect 6628 431 6662 470
rect 6692 670 6726 709
rect 6692 642 6695 670
rect 6723 642 6726 670
rect 6692 584 6726 642
rect 6692 556 6695 584
rect 6723 556 6726 584
rect 6692 498 6726 556
rect 6692 470 6695 498
rect 6723 470 6726 498
rect 6692 431 6726 470
rect 6756 670 6790 709
rect 6756 642 6759 670
rect 6787 642 6790 670
rect 6756 584 6790 642
rect 6756 556 6759 584
rect 6787 556 6790 584
rect 6756 498 6790 556
rect 6756 470 6759 498
rect 6787 470 6790 498
rect 6756 431 6790 470
rect 6820 670 6854 709
rect 6820 642 6823 670
rect 6851 642 6854 670
rect 6820 584 6854 642
rect 6820 556 6823 584
rect 6851 556 6854 584
rect 6820 498 6854 556
rect 6820 470 6823 498
rect 6851 470 6854 498
rect 6820 431 6854 470
rect 6884 670 6918 709
rect 6884 642 6887 670
rect 6915 642 6918 670
rect 6884 584 6918 642
rect 6884 556 6887 584
rect 6915 556 6918 584
rect 6884 498 6918 556
rect 6884 470 6887 498
rect 6915 470 6918 498
rect 6884 431 6918 470
rect 6948 670 6982 709
rect 6948 642 6951 670
rect 6979 642 6982 670
rect 6948 584 6982 642
rect 6948 556 6951 584
rect 6979 556 6982 584
rect 6948 498 6982 556
rect 6948 470 6951 498
rect 6979 470 6982 498
rect 6948 431 6982 470
rect 7012 670 7046 709
rect 7012 642 7015 670
rect 7043 642 7046 670
rect 7012 584 7046 642
rect 7012 556 7015 584
rect 7043 556 7046 584
rect 7012 498 7046 556
rect 7012 470 7015 498
rect 7043 470 7046 498
rect 7012 431 7046 470
rect 7078 670 7112 709
rect 7078 642 7081 670
rect 7109 642 7112 670
rect 7078 584 7112 642
rect 7078 556 7081 584
rect 7109 556 7112 584
rect 7078 498 7112 556
rect 7078 470 7081 498
rect 7109 470 7112 498
rect 7078 431 7112 470
rect 7142 670 7176 709
rect 7142 642 7145 670
rect 7173 642 7176 670
rect 7142 584 7176 642
rect 7142 556 7145 584
rect 7173 556 7176 584
rect 7142 498 7176 556
rect 7142 470 7145 498
rect 7173 470 7176 498
rect 7142 431 7176 470
rect 7206 670 7240 709
rect 7206 642 7209 670
rect 7237 642 7240 670
rect 7206 584 7240 642
rect 7206 556 7209 584
rect 7237 556 7240 584
rect 7206 498 7240 556
rect 7206 470 7209 498
rect 7237 470 7240 498
rect 7206 431 7240 470
rect 7270 670 7304 709
rect 7270 642 7273 670
rect 7301 642 7304 670
rect 7270 584 7304 642
rect 7270 556 7273 584
rect 7301 556 7304 584
rect 7270 498 7304 556
rect 7270 470 7273 498
rect 7301 470 7304 498
rect 7270 431 7304 470
rect 7334 670 7368 709
rect 7334 642 7337 670
rect 7365 642 7368 670
rect 7334 584 7368 642
rect 7334 556 7337 584
rect 7365 556 7368 584
rect 7334 498 7368 556
rect 7334 470 7337 498
rect 7365 470 7368 498
rect 7334 431 7368 470
rect 7398 670 7432 709
rect 7398 642 7401 670
rect 7429 642 7432 670
rect 7398 584 7432 642
rect 7398 556 7401 584
rect 7429 556 7432 584
rect 7398 498 7432 556
rect 7398 470 7401 498
rect 7429 470 7432 498
rect 7398 431 7432 470
rect 7462 670 7496 709
rect 7462 642 7465 670
rect 7493 642 7496 670
rect 7462 584 7496 642
rect 7462 556 7465 584
rect 7493 556 7496 584
rect 7462 498 7496 556
rect 7462 470 7465 498
rect 7493 470 7496 498
rect 7462 431 7496 470
rect 7526 670 7560 709
rect 7526 642 7529 670
rect 7557 642 7560 670
rect 7526 584 7560 642
rect 7526 556 7529 584
rect 7557 556 7560 584
rect 7526 498 7560 556
rect 7526 470 7529 498
rect 7557 470 7560 498
rect 7526 431 7560 470
rect 7590 670 7624 709
rect 7590 642 7593 670
rect 7621 642 7624 670
rect 7590 584 7624 642
rect 7590 556 7593 584
rect 7621 556 7624 584
rect 7590 498 7624 556
rect 7590 470 7593 498
rect 7621 470 7624 498
rect 7590 431 7624 470
rect 7654 670 7688 709
rect 7654 642 7657 670
rect 7685 642 7688 670
rect 7654 584 7688 642
rect 7654 556 7657 584
rect 7685 556 7688 584
rect 7654 498 7688 556
rect 7654 470 7657 498
rect 7685 470 7688 498
rect 7654 431 7688 470
rect 7720 670 7754 709
rect 7720 642 7723 670
rect 7751 642 7754 670
rect 7720 584 7754 642
rect 7720 556 7723 584
rect 7751 556 7754 584
rect 7720 498 7754 556
rect 7720 470 7723 498
rect 7751 470 7754 498
rect 7720 431 7754 470
rect 7784 670 7818 709
rect 7784 642 7787 670
rect 7815 642 7818 670
rect 7784 584 7818 642
rect 7784 556 7787 584
rect 7815 556 7818 584
rect 7784 498 7818 556
rect 7784 470 7787 498
rect 7815 470 7818 498
rect 7784 431 7818 470
rect 7848 670 7882 709
rect 7848 642 7851 670
rect 7879 642 7882 670
rect 7848 584 7882 642
rect 7848 556 7851 584
rect 7879 556 7882 584
rect 7848 498 7882 556
rect 7848 470 7851 498
rect 7879 470 7882 498
rect 7848 431 7882 470
rect 7912 670 7946 709
rect 7912 642 7915 670
rect 7943 642 7946 670
rect 7912 584 7946 642
rect 7912 556 7915 584
rect 7943 556 7946 584
rect 7912 498 7946 556
rect 7912 470 7915 498
rect 7943 470 7946 498
rect 7912 431 7946 470
rect 7976 670 8010 709
rect 7976 642 7979 670
rect 8007 642 8010 670
rect 7976 584 8010 642
rect 7976 556 7979 584
rect 8007 556 8010 584
rect 7976 498 8010 556
rect 7976 470 7979 498
rect 8007 470 8010 498
rect 7976 431 8010 470
rect 8040 670 8074 709
rect 8040 642 8043 670
rect 8071 642 8074 670
rect 8040 584 8074 642
rect 8040 556 8043 584
rect 8071 556 8074 584
rect 8040 498 8074 556
rect 8040 470 8043 498
rect 8071 470 8074 498
rect 8040 431 8074 470
rect 8104 670 8138 709
rect 8104 642 8107 670
rect 8135 642 8138 670
rect 8104 584 8138 642
rect 8104 556 8107 584
rect 8135 556 8138 584
rect 8104 498 8138 556
rect 8104 470 8107 498
rect 8135 470 8138 498
rect 8104 431 8138 470
rect 8168 670 8202 709
rect 8168 642 8171 670
rect 8199 642 8202 670
rect 8168 584 8202 642
rect 8168 556 8171 584
rect 8199 556 8202 584
rect 8168 498 8202 556
rect 8168 470 8171 498
rect 8199 470 8202 498
rect 8168 431 8202 470
rect 8232 670 8266 709
rect 8232 642 8235 670
rect 8263 642 8266 670
rect 8232 584 8266 642
rect 8232 556 8235 584
rect 8263 556 8266 584
rect 8232 498 8266 556
rect 8232 470 8235 498
rect 8263 470 8266 498
rect 8232 431 8266 470
rect 8296 670 8330 709
rect 8296 642 8299 670
rect 8327 642 8330 670
rect 8296 584 8330 642
rect 8296 556 8299 584
rect 8327 556 8330 584
rect 8296 498 8330 556
rect 8296 470 8299 498
rect 8327 470 8330 498
rect 8296 431 8330 470
rect 8362 670 8396 709
rect 8362 642 8365 670
rect 8393 642 8396 670
rect 8362 584 8396 642
rect 8362 556 8365 584
rect 8393 556 8396 584
rect 8362 498 8396 556
rect 8362 470 8365 498
rect 8393 470 8396 498
rect 8362 431 8396 470
rect 8426 670 8460 709
rect 8426 642 8429 670
rect 8457 642 8460 670
rect 8426 584 8460 642
rect 8426 556 8429 584
rect 8457 556 8460 584
rect 8426 498 8460 556
rect 8426 470 8429 498
rect 8457 470 8460 498
rect 8426 431 8460 470
rect 8490 670 8524 709
rect 8490 642 8493 670
rect 8521 642 8524 670
rect 8490 584 8524 642
rect 8490 556 8493 584
rect 8521 556 8524 584
rect 8490 498 8524 556
rect 8490 470 8493 498
rect 8521 470 8524 498
rect 8490 431 8524 470
rect 8554 670 8588 709
rect 8554 642 8557 670
rect 8585 642 8588 670
rect 8554 584 8588 642
rect 8554 556 8557 584
rect 8585 556 8588 584
rect 8554 498 8588 556
rect 8554 470 8557 498
rect 8585 470 8588 498
rect 8554 431 8588 470
rect 8618 670 8652 709
rect 8618 642 8621 670
rect 8649 642 8652 670
rect 8618 584 8652 642
rect 8618 556 8621 584
rect 8649 556 8652 584
rect 8618 498 8652 556
rect 8618 470 8621 498
rect 8649 470 8652 498
rect 8618 431 8652 470
rect 8682 670 8716 709
rect 8682 642 8685 670
rect 8713 642 8716 670
rect 8682 584 8716 642
rect 8682 556 8685 584
rect 8713 556 8716 584
rect 8682 498 8716 556
rect 8682 470 8685 498
rect 8713 470 8716 498
rect 8682 431 8716 470
rect 8746 670 8780 709
rect 8746 642 8749 670
rect 8777 642 8780 670
rect 8746 584 8780 642
rect 8746 556 8749 584
rect 8777 556 8780 584
rect 8746 498 8780 556
rect 8746 470 8749 498
rect 8777 470 8780 498
rect 8746 431 8780 470
rect 8810 670 8844 709
rect 8810 642 8813 670
rect 8841 642 8844 670
rect 8810 584 8844 642
rect 8810 556 8813 584
rect 8841 556 8844 584
rect 8810 498 8844 556
rect 8810 470 8813 498
rect 8841 470 8844 498
rect 8810 431 8844 470
rect 8874 670 8908 709
rect 8874 642 8877 670
rect 8905 642 8908 670
rect 8874 584 8908 642
rect 8874 556 8877 584
rect 8905 556 8908 584
rect 8874 498 8908 556
rect 8874 470 8877 498
rect 8905 470 8908 498
rect 8874 431 8908 470
rect 8938 670 8972 709
rect 8938 642 8941 670
rect 8969 642 8972 670
rect 8938 584 8972 642
rect 8938 556 8941 584
rect 8969 556 8972 584
rect 8938 498 8972 556
rect 8938 470 8941 498
rect 8969 470 8972 498
rect 8938 431 8972 470
rect 9004 670 9038 709
rect 9004 642 9007 670
rect 9035 642 9038 670
rect 9004 584 9038 642
rect 9004 556 9007 584
rect 9035 556 9038 584
rect 9004 498 9038 556
rect 9004 470 9007 498
rect 9035 470 9038 498
rect 9004 431 9038 470
rect 9068 670 9102 709
rect 9068 642 9071 670
rect 9099 642 9102 670
rect 9068 584 9102 642
rect 9068 556 9071 584
rect 9099 556 9102 584
rect 9068 498 9102 556
rect 9068 470 9071 498
rect 9099 470 9102 498
rect 9068 431 9102 470
rect 9132 670 9166 709
rect 9132 642 9135 670
rect 9163 642 9166 670
rect 9132 584 9166 642
rect 9132 556 9135 584
rect 9163 556 9166 584
rect 9132 498 9166 556
rect 9132 470 9135 498
rect 9163 470 9166 498
rect 9132 431 9166 470
rect 9196 670 9230 709
rect 9196 642 9199 670
rect 9227 642 9230 670
rect 9196 584 9230 642
rect 9196 556 9199 584
rect 9227 556 9230 584
rect 9196 498 9230 556
rect 9196 470 9199 498
rect 9227 470 9230 498
rect 9196 431 9230 470
rect 9260 670 9294 709
rect 9260 642 9263 670
rect 9291 642 9294 670
rect 9260 584 9294 642
rect 9260 556 9263 584
rect 9291 556 9294 584
rect 9260 498 9294 556
rect 9260 470 9263 498
rect 9291 470 9294 498
rect 9260 431 9294 470
rect 9324 670 9358 709
rect 9324 642 9327 670
rect 9355 642 9358 670
rect 9324 584 9358 642
rect 9324 556 9327 584
rect 9355 556 9358 584
rect 9324 498 9358 556
rect 9324 470 9327 498
rect 9355 470 9358 498
rect 9324 431 9358 470
rect 9388 670 9422 709
rect 9388 642 9391 670
rect 9419 642 9422 670
rect 9388 584 9422 642
rect 9388 556 9391 584
rect 9419 556 9422 584
rect 9388 498 9422 556
rect 9388 470 9391 498
rect 9419 470 9422 498
rect 9388 431 9422 470
rect 9452 670 9486 709
rect 9452 642 9455 670
rect 9483 642 9486 670
rect 9452 584 9486 642
rect 9452 556 9455 584
rect 9483 556 9486 584
rect 9452 498 9486 556
rect 9452 470 9455 498
rect 9483 470 9486 498
rect 9452 431 9486 470
rect 9516 670 9550 709
rect 9516 642 9519 670
rect 9547 642 9550 670
rect 9516 584 9550 642
rect 9516 556 9519 584
rect 9547 556 9550 584
rect 9516 498 9550 556
rect 9516 470 9519 498
rect 9547 470 9550 498
rect 9516 431 9550 470
rect 9580 670 9614 709
rect 9580 642 9583 670
rect 9611 642 9614 670
rect 9580 584 9614 642
rect 9580 556 9583 584
rect 9611 556 9614 584
rect 9580 498 9614 556
rect 9580 470 9583 498
rect 9611 470 9614 498
rect 9580 431 9614 470
rect 9646 670 9680 709
rect 9646 642 9649 670
rect 9677 642 9680 670
rect 9646 584 9680 642
rect 9646 556 9649 584
rect 9677 556 9680 584
rect 9646 498 9680 556
rect 9646 470 9649 498
rect 9677 470 9680 498
rect 9646 431 9680 470
rect 9710 670 9744 709
rect 9710 642 9713 670
rect 9741 642 9744 670
rect 9710 584 9744 642
rect 9710 556 9713 584
rect 9741 556 9744 584
rect 9710 498 9744 556
rect 9710 470 9713 498
rect 9741 470 9744 498
rect 9710 431 9744 470
rect 9774 670 9808 709
rect 9774 642 9777 670
rect 9805 642 9808 670
rect 9774 584 9808 642
rect 9774 556 9777 584
rect 9805 556 9808 584
rect 9774 498 9808 556
rect 9774 470 9777 498
rect 9805 470 9808 498
rect 9774 431 9808 470
rect 9838 670 9872 709
rect 9838 642 9841 670
rect 9869 642 9872 670
rect 9838 584 9872 642
rect 9838 556 9841 584
rect 9869 556 9872 584
rect 9838 498 9872 556
rect 9838 470 9841 498
rect 9869 470 9872 498
rect 9838 431 9872 470
rect 9902 670 9936 709
rect 9902 642 9905 670
rect 9933 642 9936 670
rect 9902 584 9936 642
rect 9902 556 9905 584
rect 9933 556 9936 584
rect 9902 498 9936 556
rect 9902 470 9905 498
rect 9933 470 9936 498
rect 9902 431 9936 470
rect 9966 670 10000 709
rect 9966 642 9969 670
rect 9997 642 10000 670
rect 9966 584 10000 642
rect 9966 556 9969 584
rect 9997 556 10000 584
rect 9966 498 10000 556
rect 9966 470 9969 498
rect 9997 470 10000 498
rect 9966 431 10000 470
rect 10030 670 10064 709
rect 10030 642 10033 670
rect 10061 642 10064 670
rect 10030 584 10064 642
rect 10030 556 10033 584
rect 10061 556 10064 584
rect 10030 498 10064 556
rect 10030 470 10033 498
rect 10061 470 10064 498
rect 10030 431 10064 470
rect 10094 670 10128 709
rect 10094 642 10097 670
rect 10125 642 10128 670
rect 10094 584 10128 642
rect 10094 556 10097 584
rect 10125 556 10128 584
rect 10094 498 10128 556
rect 10094 470 10097 498
rect 10125 470 10128 498
rect 10094 431 10128 470
rect 10158 670 10192 709
rect 10158 642 10161 670
rect 10189 642 10192 670
rect 10158 584 10192 642
rect 10158 556 10161 584
rect 10189 556 10192 584
rect 10158 498 10192 556
rect 10158 470 10161 498
rect 10189 470 10192 498
rect 10158 431 10192 470
rect 10222 670 10256 709
rect 10222 642 10225 670
rect 10253 642 10256 670
rect 10222 584 10256 642
rect 10222 556 10225 584
rect 10253 556 10256 584
rect 10222 498 10256 556
rect 10222 470 10225 498
rect 10253 470 10256 498
rect 10222 431 10256 470
rect 10288 670 10322 709
rect 10288 642 10291 670
rect 10319 642 10322 670
rect 10288 584 10322 642
rect 10288 556 10291 584
rect 10319 556 10322 584
rect 10288 498 10322 556
rect 10288 470 10291 498
rect 10319 470 10322 498
rect 10288 431 10322 470
rect 10352 670 10386 709
rect 10352 642 10355 670
rect 10383 642 10386 670
rect 10352 584 10386 642
rect 10352 556 10355 584
rect 10383 556 10386 584
rect 10352 498 10386 556
rect 10352 470 10355 498
rect 10383 470 10386 498
rect 10352 431 10386 470
rect 10416 670 10450 709
rect 10416 642 10419 670
rect 10447 642 10450 670
rect 10416 584 10450 642
rect 10416 556 10419 584
rect 10447 556 10450 584
rect 10416 498 10450 556
rect 10416 470 10419 498
rect 10447 470 10450 498
rect 10416 431 10450 470
rect 10480 670 10514 709
rect 10480 642 10483 670
rect 10511 642 10514 670
rect 10480 584 10514 642
rect 10480 556 10483 584
rect 10511 556 10514 584
rect 10480 498 10514 556
rect 10480 470 10483 498
rect 10511 470 10514 498
rect 10480 431 10514 470
rect 10544 670 10578 709
rect 10544 642 10547 670
rect 10575 642 10578 670
rect 10544 584 10578 642
rect 10544 556 10547 584
rect 10575 556 10578 584
rect 10544 498 10578 556
rect 10544 470 10547 498
rect 10575 470 10578 498
rect 10544 431 10578 470
rect 10608 670 10642 709
rect 10608 642 10611 670
rect 10639 642 10642 670
rect 10608 584 10642 642
rect 10608 556 10611 584
rect 10639 556 10642 584
rect 10608 498 10642 556
rect 10608 470 10611 498
rect 10639 470 10642 498
rect 10608 431 10642 470
rect 10672 670 10706 709
rect 10672 642 10675 670
rect 10703 642 10706 670
rect 10672 584 10706 642
rect 10672 556 10675 584
rect 10703 556 10706 584
rect 10672 498 10706 556
rect 10672 470 10675 498
rect 10703 470 10706 498
rect 10672 431 10706 470
rect 10736 670 10770 709
rect 10736 642 10739 670
rect 10767 642 10770 670
rect 10736 584 10770 642
rect 10736 556 10739 584
rect 10767 556 10770 584
rect 10736 498 10770 556
rect 10736 470 10739 498
rect 10767 470 10770 498
rect 10736 431 10770 470
rect 10800 670 10834 709
rect 10800 642 10803 670
rect 10831 642 10834 670
rect 10800 584 10834 642
rect 10800 556 10803 584
rect 10831 556 10834 584
rect 10800 498 10834 556
rect 10800 470 10803 498
rect 10831 470 10834 498
rect 10800 431 10834 470
rect 10864 670 10898 709
rect 10864 642 10867 670
rect 10895 642 10898 670
rect 10864 584 10898 642
rect 10864 556 10867 584
rect 10895 556 10898 584
rect 10864 498 10898 556
rect 10864 470 10867 498
rect 10895 470 10898 498
rect 10864 431 10898 470
rect 10930 670 10964 709
rect 10930 642 10933 670
rect 10961 642 10964 670
rect 10930 584 10964 642
rect 10930 556 10933 584
rect 10961 556 10964 584
rect 10930 498 10964 556
rect 10930 470 10933 498
rect 10961 470 10964 498
rect 10930 431 10964 470
rect 10994 670 11028 709
rect 10994 642 10997 670
rect 11025 642 11028 670
rect 10994 584 11028 642
rect 10994 556 10997 584
rect 11025 556 11028 584
rect 10994 498 11028 556
rect 10994 470 10997 498
rect 11025 470 11028 498
rect 10994 431 11028 470
rect 11058 670 11092 709
rect 11058 642 11061 670
rect 11089 642 11092 670
rect 11058 584 11092 642
rect 11058 556 11061 584
rect 11089 556 11092 584
rect 11058 498 11092 556
rect 11058 470 11061 498
rect 11089 470 11092 498
rect 11058 431 11092 470
rect 11122 670 11156 709
rect 11122 642 11125 670
rect 11153 642 11156 670
rect 11122 584 11156 642
rect 11122 556 11125 584
rect 11153 556 11156 584
rect 11122 498 11156 556
rect 11122 470 11125 498
rect 11153 470 11156 498
rect 11122 431 11156 470
rect 11186 670 11220 709
rect 11186 642 11189 670
rect 11217 642 11220 670
rect 11186 584 11220 642
rect 11186 556 11189 584
rect 11217 556 11220 584
rect 11186 498 11220 556
rect 11186 470 11189 498
rect 11217 470 11220 498
rect 11186 431 11220 470
rect 11250 670 11284 709
rect 11250 642 11253 670
rect 11281 642 11284 670
rect 11250 584 11284 642
rect 11250 556 11253 584
rect 11281 556 11284 584
rect 11250 498 11284 556
rect 11250 470 11253 498
rect 11281 470 11284 498
rect 11250 431 11284 470
rect 11314 670 11348 709
rect 11314 642 11317 670
rect 11345 642 11348 670
rect 11314 584 11348 642
rect 11314 556 11317 584
rect 11345 556 11348 584
rect 11314 498 11348 556
rect 11314 470 11317 498
rect 11345 470 11348 498
rect 11314 431 11348 470
rect 11378 670 11412 709
rect 11378 642 11381 670
rect 11409 642 11412 670
rect 11378 584 11412 642
rect 11378 556 11381 584
rect 11409 556 11412 584
rect 11378 498 11412 556
rect 11378 470 11381 498
rect 11409 470 11412 498
rect 11378 431 11412 470
rect 11442 670 11476 709
rect 11442 642 11445 670
rect 11473 642 11476 670
rect 11442 584 11476 642
rect 11442 556 11445 584
rect 11473 556 11476 584
rect 11442 498 11476 556
rect 11442 470 11445 498
rect 11473 470 11476 498
rect 11442 431 11476 470
rect 11506 670 11540 709
rect 11506 642 11509 670
rect 11537 642 11540 670
rect 11506 584 11540 642
rect 11506 556 11509 584
rect 11537 556 11540 584
rect 11506 498 11540 556
rect 11506 470 11509 498
rect 11537 470 11540 498
rect 11506 431 11540 470
rect 11572 670 11606 709
rect 11572 642 11575 670
rect 11603 642 11606 670
rect 11572 584 11606 642
rect 11572 556 11575 584
rect 11603 556 11606 584
rect 11572 498 11606 556
rect 11572 470 11575 498
rect 11603 470 11606 498
rect 11572 431 11606 470
rect 11636 670 11670 709
rect 11636 642 11639 670
rect 11667 642 11670 670
rect 11636 584 11670 642
rect 11636 556 11639 584
rect 11667 556 11670 584
rect 11636 498 11670 556
rect 11636 470 11639 498
rect 11667 470 11670 498
rect 11636 431 11670 470
rect 11700 670 11734 709
rect 11700 642 11703 670
rect 11731 642 11734 670
rect 11700 584 11734 642
rect 11700 556 11703 584
rect 11731 556 11734 584
rect 11700 498 11734 556
rect 11700 470 11703 498
rect 11731 470 11734 498
rect 11700 431 11734 470
rect 11764 670 11798 709
rect 11764 642 11767 670
rect 11795 642 11798 670
rect 11764 584 11798 642
rect 11764 556 11767 584
rect 11795 556 11798 584
rect 11764 498 11798 556
rect 11764 470 11767 498
rect 11795 470 11798 498
rect 11764 431 11798 470
rect 11828 670 11862 709
rect 11828 642 11831 670
rect 11859 642 11862 670
rect 11828 584 11862 642
rect 11828 556 11831 584
rect 11859 556 11862 584
rect 11828 498 11862 556
rect 11828 470 11831 498
rect 11859 470 11862 498
rect 11828 431 11862 470
rect 11892 670 11926 709
rect 11892 642 11895 670
rect 11923 642 11926 670
rect 11892 584 11926 642
rect 11892 556 11895 584
rect 11923 556 11926 584
rect 11892 498 11926 556
rect 11892 470 11895 498
rect 11923 470 11926 498
rect 11892 431 11926 470
rect 11956 670 11990 709
rect 11956 642 11959 670
rect 11987 642 11990 670
rect 11956 584 11990 642
rect 11956 556 11959 584
rect 11987 556 11990 584
rect 11956 498 11990 556
rect 11956 470 11959 498
rect 11987 470 11990 498
rect 11956 431 11990 470
rect 12020 670 12054 709
rect 12020 642 12023 670
rect 12051 642 12054 670
rect 12020 584 12054 642
rect 12020 556 12023 584
rect 12051 556 12054 584
rect 12020 498 12054 556
rect 12020 470 12023 498
rect 12051 470 12054 498
rect 12020 431 12054 470
rect 12084 670 12118 709
rect 12084 642 12087 670
rect 12115 642 12118 670
rect 12084 584 12118 642
rect 12084 556 12087 584
rect 12115 556 12118 584
rect 12084 498 12118 556
rect 12084 470 12087 498
rect 12115 470 12118 498
rect 12084 431 12118 470
rect 12148 670 12182 709
rect 12148 642 12151 670
rect 12179 642 12182 670
rect 12148 584 12182 642
rect 12148 556 12151 584
rect 12179 556 12182 584
rect 12148 498 12182 556
rect 12148 470 12151 498
rect 12179 470 12182 498
rect 12148 431 12182 470
rect 12214 670 12248 709
rect 12214 642 12217 670
rect 12245 642 12248 670
rect 12214 584 12248 642
rect 12214 556 12217 584
rect 12245 556 12248 584
rect 12214 498 12248 556
rect 12214 470 12217 498
rect 12245 470 12248 498
rect 12214 431 12248 470
rect 12278 670 12312 709
rect 12278 642 12281 670
rect 12309 642 12312 670
rect 12278 584 12312 642
rect 12278 556 12281 584
rect 12309 556 12312 584
rect 12278 498 12312 556
rect 12278 470 12281 498
rect 12309 470 12312 498
rect 12278 431 12312 470
rect 12342 670 12376 709
rect 12342 642 12345 670
rect 12373 642 12376 670
rect 12342 584 12376 642
rect 12342 556 12345 584
rect 12373 556 12376 584
rect 12342 498 12376 556
rect 12342 470 12345 498
rect 12373 470 12376 498
rect 12342 431 12376 470
rect 12406 670 12440 709
rect 12406 642 12409 670
rect 12437 642 12440 670
rect 12406 584 12440 642
rect 12406 556 12409 584
rect 12437 556 12440 584
rect 12406 498 12440 556
rect 12406 470 12409 498
rect 12437 470 12440 498
rect 12406 431 12440 470
rect 12470 670 12504 709
rect 12470 642 12473 670
rect 12501 642 12504 670
rect 12470 584 12504 642
rect 12470 556 12473 584
rect 12501 556 12504 584
rect 12470 498 12504 556
rect 12470 470 12473 498
rect 12501 470 12504 498
rect 12470 431 12504 470
rect 12534 670 12568 709
rect 12534 642 12537 670
rect 12565 642 12568 670
rect 12534 584 12568 642
rect 12534 556 12537 584
rect 12565 556 12568 584
rect 12534 498 12568 556
rect 12534 470 12537 498
rect 12565 470 12568 498
rect 12534 431 12568 470
rect 12598 670 12632 709
rect 12598 642 12601 670
rect 12629 642 12632 670
rect 12598 584 12632 642
rect 12598 556 12601 584
rect 12629 556 12632 584
rect 12598 498 12632 556
rect 12598 470 12601 498
rect 12629 470 12632 498
rect 12598 431 12632 470
rect 12662 670 12696 709
rect 12662 642 12665 670
rect 12693 642 12696 670
rect 12662 584 12696 642
rect 12662 556 12665 584
rect 12693 556 12696 584
rect 12662 498 12696 556
rect 12662 470 12665 498
rect 12693 470 12696 498
rect 12662 431 12696 470
rect 12726 670 12760 709
rect 12726 642 12729 670
rect 12757 642 12760 670
rect 12726 584 12760 642
rect 12726 556 12729 584
rect 12757 556 12760 584
rect 12726 498 12760 556
rect 12726 470 12729 498
rect 12757 470 12760 498
rect 12726 431 12760 470
rect 12790 670 12824 709
rect 12790 642 12793 670
rect 12821 642 12824 670
rect 12790 584 12824 642
rect 12790 556 12793 584
rect 12821 556 12824 584
rect 12790 498 12824 556
rect 12790 470 12793 498
rect 12821 470 12824 498
rect 12790 431 12824 470
rect 16 290 50 329
rect 16 262 19 290
rect 47 262 50 290
rect 16 204 50 262
rect 16 176 19 204
rect 47 176 50 204
rect 16 118 50 176
rect 16 90 19 118
rect 47 90 50 118
rect 16 51 50 90
rect 80 290 114 329
rect 80 262 83 290
rect 111 262 114 290
rect 80 204 114 262
rect 80 176 83 204
rect 111 176 114 204
rect 80 118 114 176
rect 80 90 83 118
rect 111 90 114 118
rect 80 51 114 90
rect 144 290 178 329
rect 144 262 147 290
rect 175 262 178 290
rect 144 204 178 262
rect 144 176 147 204
rect 175 176 178 204
rect 144 118 178 176
rect 144 90 147 118
rect 175 90 178 118
rect 144 51 178 90
rect 208 290 242 329
rect 208 262 211 290
rect 239 262 242 290
rect 208 204 242 262
rect 208 176 211 204
rect 239 176 242 204
rect 208 118 242 176
rect 208 90 211 118
rect 239 90 242 118
rect 208 51 242 90
rect 272 290 306 329
rect 272 262 275 290
rect 303 262 306 290
rect 272 204 306 262
rect 272 176 275 204
rect 303 176 306 204
rect 272 118 306 176
rect 272 90 275 118
rect 303 90 306 118
rect 272 51 306 90
rect 336 290 370 329
rect 336 262 339 290
rect 367 262 370 290
rect 336 204 370 262
rect 336 176 339 204
rect 367 176 370 204
rect 336 118 370 176
rect 336 90 339 118
rect 367 90 370 118
rect 336 51 370 90
rect 400 290 434 329
rect 400 262 403 290
rect 431 262 434 290
rect 400 204 434 262
rect 400 176 403 204
rect 431 176 434 204
rect 400 118 434 176
rect 400 90 403 118
rect 431 90 434 118
rect 400 51 434 90
rect 464 290 498 329
rect 464 262 467 290
rect 495 262 498 290
rect 464 204 498 262
rect 464 176 467 204
rect 495 176 498 204
rect 464 118 498 176
rect 464 90 467 118
rect 495 90 498 118
rect 464 51 498 90
rect 528 290 562 329
rect 528 262 531 290
rect 559 262 562 290
rect 528 204 562 262
rect 528 176 531 204
rect 559 176 562 204
rect 528 118 562 176
rect 528 90 531 118
rect 559 90 562 118
rect 528 51 562 90
rect 592 290 626 329
rect 592 262 595 290
rect 623 262 626 290
rect 592 204 626 262
rect 592 176 595 204
rect 623 176 626 204
rect 592 118 626 176
rect 592 90 595 118
rect 623 90 626 118
rect 592 51 626 90
rect 658 290 692 329
rect 658 262 661 290
rect 689 262 692 290
rect 658 204 692 262
rect 658 176 661 204
rect 689 176 692 204
rect 658 118 692 176
rect 658 90 661 118
rect 689 90 692 118
rect 658 51 692 90
rect 722 290 756 329
rect 722 262 725 290
rect 753 262 756 290
rect 722 204 756 262
rect 722 176 725 204
rect 753 176 756 204
rect 722 118 756 176
rect 722 90 725 118
rect 753 90 756 118
rect 722 51 756 90
rect 786 290 820 329
rect 786 262 789 290
rect 817 262 820 290
rect 786 204 820 262
rect 786 176 789 204
rect 817 176 820 204
rect 786 118 820 176
rect 786 90 789 118
rect 817 90 820 118
rect 786 51 820 90
rect 850 290 884 329
rect 850 262 853 290
rect 881 262 884 290
rect 850 204 884 262
rect 850 176 853 204
rect 881 176 884 204
rect 850 118 884 176
rect 850 90 853 118
rect 881 90 884 118
rect 850 51 884 90
rect 914 290 948 329
rect 914 262 917 290
rect 945 262 948 290
rect 914 204 948 262
rect 914 176 917 204
rect 945 176 948 204
rect 914 118 948 176
rect 914 90 917 118
rect 945 90 948 118
rect 914 51 948 90
rect 978 290 1012 329
rect 978 262 981 290
rect 1009 262 1012 290
rect 978 204 1012 262
rect 978 176 981 204
rect 1009 176 1012 204
rect 978 118 1012 176
rect 978 90 981 118
rect 1009 90 1012 118
rect 978 51 1012 90
rect 1042 290 1076 329
rect 1042 262 1045 290
rect 1073 262 1076 290
rect 1042 204 1076 262
rect 1042 176 1045 204
rect 1073 176 1076 204
rect 1042 118 1076 176
rect 1042 90 1045 118
rect 1073 90 1076 118
rect 1042 51 1076 90
rect 1106 290 1140 329
rect 1106 262 1109 290
rect 1137 262 1140 290
rect 1106 204 1140 262
rect 1106 176 1109 204
rect 1137 176 1140 204
rect 1106 118 1140 176
rect 1106 90 1109 118
rect 1137 90 1140 118
rect 1106 51 1140 90
rect 1170 290 1204 329
rect 1170 262 1173 290
rect 1201 262 1204 290
rect 1170 204 1204 262
rect 1170 176 1173 204
rect 1201 176 1204 204
rect 1170 118 1204 176
rect 1170 90 1173 118
rect 1201 90 1204 118
rect 1170 51 1204 90
rect 1234 290 1268 329
rect 1234 262 1237 290
rect 1265 262 1268 290
rect 1234 204 1268 262
rect 1234 176 1237 204
rect 1265 176 1268 204
rect 1234 118 1268 176
rect 1234 90 1237 118
rect 1265 90 1268 118
rect 1234 51 1268 90
rect 1300 290 1334 329
rect 1300 262 1303 290
rect 1331 262 1334 290
rect 1300 204 1334 262
rect 1300 176 1303 204
rect 1331 176 1334 204
rect 1300 118 1334 176
rect 1300 90 1303 118
rect 1331 90 1334 118
rect 1300 51 1334 90
rect 1364 290 1398 329
rect 1364 262 1367 290
rect 1395 262 1398 290
rect 1364 204 1398 262
rect 1364 176 1367 204
rect 1395 176 1398 204
rect 1364 118 1398 176
rect 1364 90 1367 118
rect 1395 90 1398 118
rect 1364 51 1398 90
rect 1428 290 1462 329
rect 1428 262 1431 290
rect 1459 262 1462 290
rect 1428 204 1462 262
rect 1428 176 1431 204
rect 1459 176 1462 204
rect 1428 118 1462 176
rect 1428 90 1431 118
rect 1459 90 1462 118
rect 1428 51 1462 90
rect 1492 290 1526 329
rect 1492 262 1495 290
rect 1523 262 1526 290
rect 1492 204 1526 262
rect 1492 176 1495 204
rect 1523 176 1526 204
rect 1492 118 1526 176
rect 1492 90 1495 118
rect 1523 90 1526 118
rect 1492 51 1526 90
rect 1556 290 1590 329
rect 1556 262 1559 290
rect 1587 262 1590 290
rect 1556 204 1590 262
rect 1556 176 1559 204
rect 1587 176 1590 204
rect 1556 118 1590 176
rect 1556 90 1559 118
rect 1587 90 1590 118
rect 1556 51 1590 90
rect 1620 290 1654 329
rect 1620 262 1623 290
rect 1651 262 1654 290
rect 1620 204 1654 262
rect 1620 176 1623 204
rect 1651 176 1654 204
rect 1620 118 1654 176
rect 1620 90 1623 118
rect 1651 90 1654 118
rect 1620 51 1654 90
rect 1684 290 1718 329
rect 1684 262 1687 290
rect 1715 262 1718 290
rect 1684 204 1718 262
rect 1684 176 1687 204
rect 1715 176 1718 204
rect 1684 118 1718 176
rect 1684 90 1687 118
rect 1715 90 1718 118
rect 1684 51 1718 90
rect 1748 290 1782 329
rect 1748 262 1751 290
rect 1779 262 1782 290
rect 1748 204 1782 262
rect 1748 176 1751 204
rect 1779 176 1782 204
rect 1748 118 1782 176
rect 1748 90 1751 118
rect 1779 90 1782 118
rect 1748 51 1782 90
rect 1812 290 1846 329
rect 1812 262 1815 290
rect 1843 262 1846 290
rect 1812 204 1846 262
rect 1812 176 1815 204
rect 1843 176 1846 204
rect 1812 118 1846 176
rect 1812 90 1815 118
rect 1843 90 1846 118
rect 1812 51 1846 90
rect 1876 290 1910 329
rect 1876 262 1879 290
rect 1907 262 1910 290
rect 1876 204 1910 262
rect 1876 176 1879 204
rect 1907 176 1910 204
rect 1876 118 1910 176
rect 1876 90 1879 118
rect 1907 90 1910 118
rect 1876 51 1910 90
rect 1942 290 1976 329
rect 1942 262 1945 290
rect 1973 262 1976 290
rect 1942 204 1976 262
rect 1942 176 1945 204
rect 1973 176 1976 204
rect 1942 118 1976 176
rect 1942 90 1945 118
rect 1973 90 1976 118
rect 1942 51 1976 90
rect 2006 290 2040 329
rect 2006 262 2009 290
rect 2037 262 2040 290
rect 2006 204 2040 262
rect 2006 176 2009 204
rect 2037 176 2040 204
rect 2006 118 2040 176
rect 2006 90 2009 118
rect 2037 90 2040 118
rect 2006 51 2040 90
rect 2070 290 2104 329
rect 2070 262 2073 290
rect 2101 262 2104 290
rect 2070 204 2104 262
rect 2070 176 2073 204
rect 2101 176 2104 204
rect 2070 118 2104 176
rect 2070 90 2073 118
rect 2101 90 2104 118
rect 2070 51 2104 90
rect 2134 290 2168 329
rect 2134 262 2137 290
rect 2165 262 2168 290
rect 2134 204 2168 262
rect 2134 176 2137 204
rect 2165 176 2168 204
rect 2134 118 2168 176
rect 2134 90 2137 118
rect 2165 90 2168 118
rect 2134 51 2168 90
rect 2198 290 2232 329
rect 2198 262 2201 290
rect 2229 262 2232 290
rect 2198 204 2232 262
rect 2198 176 2201 204
rect 2229 176 2232 204
rect 2198 118 2232 176
rect 2198 90 2201 118
rect 2229 90 2232 118
rect 2198 51 2232 90
rect 2262 290 2296 329
rect 2262 262 2265 290
rect 2293 262 2296 290
rect 2262 204 2296 262
rect 2262 176 2265 204
rect 2293 176 2296 204
rect 2262 118 2296 176
rect 2262 90 2265 118
rect 2293 90 2296 118
rect 2262 51 2296 90
rect 2326 290 2360 329
rect 2326 262 2329 290
rect 2357 262 2360 290
rect 2326 204 2360 262
rect 2326 176 2329 204
rect 2357 176 2360 204
rect 2326 118 2360 176
rect 2326 90 2329 118
rect 2357 90 2360 118
rect 2326 51 2360 90
rect 2390 290 2424 329
rect 2390 262 2393 290
rect 2421 262 2424 290
rect 2390 204 2424 262
rect 2390 176 2393 204
rect 2421 176 2424 204
rect 2390 118 2424 176
rect 2390 90 2393 118
rect 2421 90 2424 118
rect 2390 51 2424 90
rect 2454 290 2488 329
rect 2454 262 2457 290
rect 2485 262 2488 290
rect 2454 204 2488 262
rect 2454 176 2457 204
rect 2485 176 2488 204
rect 2454 118 2488 176
rect 2454 90 2457 118
rect 2485 90 2488 118
rect 2454 51 2488 90
rect 2518 290 2552 329
rect 2518 262 2521 290
rect 2549 262 2552 290
rect 2518 204 2552 262
rect 2518 176 2521 204
rect 2549 176 2552 204
rect 2518 118 2552 176
rect 2518 90 2521 118
rect 2549 90 2552 118
rect 2518 51 2552 90
rect 2584 290 2618 329
rect 2584 262 2587 290
rect 2615 262 2618 290
rect 2584 204 2618 262
rect 2584 176 2587 204
rect 2615 176 2618 204
rect 2584 118 2618 176
rect 2584 90 2587 118
rect 2615 90 2618 118
rect 2584 51 2618 90
rect 2648 290 2682 329
rect 2648 262 2651 290
rect 2679 262 2682 290
rect 2648 204 2682 262
rect 2648 176 2651 204
rect 2679 176 2682 204
rect 2648 118 2682 176
rect 2648 90 2651 118
rect 2679 90 2682 118
rect 2648 51 2682 90
rect 2712 290 2746 329
rect 2712 262 2715 290
rect 2743 262 2746 290
rect 2712 204 2746 262
rect 2712 176 2715 204
rect 2743 176 2746 204
rect 2712 118 2746 176
rect 2712 90 2715 118
rect 2743 90 2746 118
rect 2712 51 2746 90
rect 2776 290 2810 329
rect 2776 262 2779 290
rect 2807 262 2810 290
rect 2776 204 2810 262
rect 2776 176 2779 204
rect 2807 176 2810 204
rect 2776 118 2810 176
rect 2776 90 2779 118
rect 2807 90 2810 118
rect 2776 51 2810 90
rect 2840 290 2874 329
rect 2840 262 2843 290
rect 2871 262 2874 290
rect 2840 204 2874 262
rect 2840 176 2843 204
rect 2871 176 2874 204
rect 2840 118 2874 176
rect 2840 90 2843 118
rect 2871 90 2874 118
rect 2840 51 2874 90
rect 2904 290 2938 329
rect 2904 262 2907 290
rect 2935 262 2938 290
rect 2904 204 2938 262
rect 2904 176 2907 204
rect 2935 176 2938 204
rect 2904 118 2938 176
rect 2904 90 2907 118
rect 2935 90 2938 118
rect 2904 51 2938 90
rect 2968 290 3002 329
rect 2968 262 2971 290
rect 2999 262 3002 290
rect 2968 204 3002 262
rect 2968 176 2971 204
rect 2999 176 3002 204
rect 2968 118 3002 176
rect 2968 90 2971 118
rect 2999 90 3002 118
rect 2968 51 3002 90
rect 3032 290 3066 329
rect 3032 262 3035 290
rect 3063 262 3066 290
rect 3032 204 3066 262
rect 3032 176 3035 204
rect 3063 176 3066 204
rect 3032 118 3066 176
rect 3032 90 3035 118
rect 3063 90 3066 118
rect 3032 51 3066 90
rect 3096 290 3130 329
rect 3096 262 3099 290
rect 3127 262 3130 290
rect 3096 204 3130 262
rect 3096 176 3099 204
rect 3127 176 3130 204
rect 3096 118 3130 176
rect 3096 90 3099 118
rect 3127 90 3130 118
rect 3096 51 3130 90
rect 3160 290 3194 329
rect 3160 262 3163 290
rect 3191 262 3194 290
rect 3160 204 3194 262
rect 3160 176 3163 204
rect 3191 176 3194 204
rect 3160 118 3194 176
rect 3160 90 3163 118
rect 3191 90 3194 118
rect 3160 51 3194 90
rect 3226 290 3260 329
rect 3226 262 3229 290
rect 3257 262 3260 290
rect 3226 204 3260 262
rect 3226 176 3229 204
rect 3257 176 3260 204
rect 3226 118 3260 176
rect 3226 90 3229 118
rect 3257 90 3260 118
rect 3226 51 3260 90
rect 3290 290 3324 329
rect 3290 262 3293 290
rect 3321 262 3324 290
rect 3290 204 3324 262
rect 3290 176 3293 204
rect 3321 176 3324 204
rect 3290 118 3324 176
rect 3290 90 3293 118
rect 3321 90 3324 118
rect 3290 51 3324 90
rect 3354 290 3388 329
rect 3354 262 3357 290
rect 3385 262 3388 290
rect 3354 204 3388 262
rect 3354 176 3357 204
rect 3385 176 3388 204
rect 3354 118 3388 176
rect 3354 90 3357 118
rect 3385 90 3388 118
rect 3354 51 3388 90
rect 3418 290 3452 329
rect 3418 262 3421 290
rect 3449 262 3452 290
rect 3418 204 3452 262
rect 3418 176 3421 204
rect 3449 176 3452 204
rect 3418 118 3452 176
rect 3418 90 3421 118
rect 3449 90 3452 118
rect 3418 51 3452 90
rect 3482 290 3516 329
rect 3482 262 3485 290
rect 3513 262 3516 290
rect 3482 204 3516 262
rect 3482 176 3485 204
rect 3513 176 3516 204
rect 3482 118 3516 176
rect 3482 90 3485 118
rect 3513 90 3516 118
rect 3482 51 3516 90
rect 3546 290 3580 329
rect 3546 262 3549 290
rect 3577 262 3580 290
rect 3546 204 3580 262
rect 3546 176 3549 204
rect 3577 176 3580 204
rect 3546 118 3580 176
rect 3546 90 3549 118
rect 3577 90 3580 118
rect 3546 51 3580 90
rect 3610 290 3644 329
rect 3610 262 3613 290
rect 3641 262 3644 290
rect 3610 204 3644 262
rect 3610 176 3613 204
rect 3641 176 3644 204
rect 3610 118 3644 176
rect 3610 90 3613 118
rect 3641 90 3644 118
rect 3610 51 3644 90
rect 3674 290 3708 329
rect 3674 262 3677 290
rect 3705 262 3708 290
rect 3674 204 3708 262
rect 3674 176 3677 204
rect 3705 176 3708 204
rect 3674 118 3708 176
rect 3674 90 3677 118
rect 3705 90 3708 118
rect 3674 51 3708 90
rect 3738 290 3772 329
rect 3738 262 3741 290
rect 3769 262 3772 290
rect 3738 204 3772 262
rect 3738 176 3741 204
rect 3769 176 3772 204
rect 3738 118 3772 176
rect 3738 90 3741 118
rect 3769 90 3772 118
rect 3738 51 3772 90
rect 3802 290 3836 329
rect 3802 262 3805 290
rect 3833 262 3836 290
rect 3802 204 3836 262
rect 3802 176 3805 204
rect 3833 176 3836 204
rect 3802 118 3836 176
rect 3802 90 3805 118
rect 3833 90 3836 118
rect 3802 51 3836 90
rect 3868 290 3902 329
rect 3868 262 3871 290
rect 3899 262 3902 290
rect 3868 204 3902 262
rect 3868 176 3871 204
rect 3899 176 3902 204
rect 3868 118 3902 176
rect 3868 90 3871 118
rect 3899 90 3902 118
rect 3868 51 3902 90
rect 3932 290 3966 329
rect 3932 262 3935 290
rect 3963 262 3966 290
rect 3932 204 3966 262
rect 3932 176 3935 204
rect 3963 176 3966 204
rect 3932 118 3966 176
rect 3932 90 3935 118
rect 3963 90 3966 118
rect 3932 51 3966 90
rect 3996 290 4030 329
rect 3996 262 3999 290
rect 4027 262 4030 290
rect 3996 204 4030 262
rect 3996 176 3999 204
rect 4027 176 4030 204
rect 3996 118 4030 176
rect 3996 90 3999 118
rect 4027 90 4030 118
rect 3996 51 4030 90
rect 4060 290 4094 329
rect 4060 262 4063 290
rect 4091 262 4094 290
rect 4060 204 4094 262
rect 4060 176 4063 204
rect 4091 176 4094 204
rect 4060 118 4094 176
rect 4060 90 4063 118
rect 4091 90 4094 118
rect 4060 51 4094 90
rect 4124 290 4158 329
rect 4124 262 4127 290
rect 4155 262 4158 290
rect 4124 204 4158 262
rect 4124 176 4127 204
rect 4155 176 4158 204
rect 4124 118 4158 176
rect 4124 90 4127 118
rect 4155 90 4158 118
rect 4124 51 4158 90
rect 4188 290 4222 329
rect 4188 262 4191 290
rect 4219 262 4222 290
rect 4188 204 4222 262
rect 4188 176 4191 204
rect 4219 176 4222 204
rect 4188 118 4222 176
rect 4188 90 4191 118
rect 4219 90 4222 118
rect 4188 51 4222 90
rect 4252 290 4286 329
rect 4252 262 4255 290
rect 4283 262 4286 290
rect 4252 204 4286 262
rect 4252 176 4255 204
rect 4283 176 4286 204
rect 4252 118 4286 176
rect 4252 90 4255 118
rect 4283 90 4286 118
rect 4252 51 4286 90
rect 4316 290 4350 329
rect 4316 262 4319 290
rect 4347 262 4350 290
rect 4316 204 4350 262
rect 4316 176 4319 204
rect 4347 176 4350 204
rect 4316 118 4350 176
rect 4316 90 4319 118
rect 4347 90 4350 118
rect 4316 51 4350 90
rect 4380 290 4414 329
rect 4380 262 4383 290
rect 4411 262 4414 290
rect 4380 204 4414 262
rect 4380 176 4383 204
rect 4411 176 4414 204
rect 4380 118 4414 176
rect 4380 90 4383 118
rect 4411 90 4414 118
rect 4380 51 4414 90
rect 4444 290 4478 329
rect 4444 262 4447 290
rect 4475 262 4478 290
rect 4444 204 4478 262
rect 4444 176 4447 204
rect 4475 176 4478 204
rect 4444 118 4478 176
rect 4444 90 4447 118
rect 4475 90 4478 118
rect 4444 51 4478 90
rect 4510 290 4544 329
rect 4510 262 4513 290
rect 4541 262 4544 290
rect 4510 204 4544 262
rect 4510 176 4513 204
rect 4541 176 4544 204
rect 4510 118 4544 176
rect 4510 90 4513 118
rect 4541 90 4544 118
rect 4510 51 4544 90
rect 4574 290 4608 329
rect 4574 262 4577 290
rect 4605 262 4608 290
rect 4574 204 4608 262
rect 4574 176 4577 204
rect 4605 176 4608 204
rect 4574 118 4608 176
rect 4574 90 4577 118
rect 4605 90 4608 118
rect 4574 51 4608 90
rect 4638 290 4672 329
rect 4638 262 4641 290
rect 4669 262 4672 290
rect 4638 204 4672 262
rect 4638 176 4641 204
rect 4669 176 4672 204
rect 4638 118 4672 176
rect 4638 90 4641 118
rect 4669 90 4672 118
rect 4638 51 4672 90
rect 4702 290 4736 329
rect 4702 262 4705 290
rect 4733 262 4736 290
rect 4702 204 4736 262
rect 4702 176 4705 204
rect 4733 176 4736 204
rect 4702 118 4736 176
rect 4702 90 4705 118
rect 4733 90 4736 118
rect 4702 51 4736 90
rect 4766 290 4800 329
rect 4766 262 4769 290
rect 4797 262 4800 290
rect 4766 204 4800 262
rect 4766 176 4769 204
rect 4797 176 4800 204
rect 4766 118 4800 176
rect 4766 90 4769 118
rect 4797 90 4800 118
rect 4766 51 4800 90
rect 4830 290 4864 329
rect 4830 262 4833 290
rect 4861 262 4864 290
rect 4830 204 4864 262
rect 4830 176 4833 204
rect 4861 176 4864 204
rect 4830 118 4864 176
rect 4830 90 4833 118
rect 4861 90 4864 118
rect 4830 51 4864 90
rect 4894 290 4928 329
rect 4894 262 4897 290
rect 4925 262 4928 290
rect 4894 204 4928 262
rect 4894 176 4897 204
rect 4925 176 4928 204
rect 4894 118 4928 176
rect 4894 90 4897 118
rect 4925 90 4928 118
rect 4894 51 4928 90
rect 4958 290 4992 329
rect 4958 262 4961 290
rect 4989 262 4992 290
rect 4958 204 4992 262
rect 4958 176 4961 204
rect 4989 176 4992 204
rect 4958 118 4992 176
rect 4958 90 4961 118
rect 4989 90 4992 118
rect 4958 51 4992 90
rect 5022 290 5056 329
rect 5022 262 5025 290
rect 5053 262 5056 290
rect 5022 204 5056 262
rect 5022 176 5025 204
rect 5053 176 5056 204
rect 5022 118 5056 176
rect 5022 90 5025 118
rect 5053 90 5056 118
rect 5022 51 5056 90
rect 5086 290 5120 329
rect 5086 262 5089 290
rect 5117 262 5120 290
rect 5086 204 5120 262
rect 5086 176 5089 204
rect 5117 176 5120 204
rect 5086 118 5120 176
rect 5086 90 5089 118
rect 5117 90 5120 118
rect 5086 51 5120 90
rect 5152 290 5186 329
rect 5152 262 5155 290
rect 5183 262 5186 290
rect 5152 204 5186 262
rect 5152 176 5155 204
rect 5183 176 5186 204
rect 5152 118 5186 176
rect 5152 90 5155 118
rect 5183 90 5186 118
rect 5152 51 5186 90
rect 5216 290 5250 329
rect 5216 262 5219 290
rect 5247 262 5250 290
rect 5216 204 5250 262
rect 5216 176 5219 204
rect 5247 176 5250 204
rect 5216 118 5250 176
rect 5216 90 5219 118
rect 5247 90 5250 118
rect 5216 51 5250 90
rect 5280 290 5314 329
rect 5280 262 5283 290
rect 5311 262 5314 290
rect 5280 204 5314 262
rect 5280 176 5283 204
rect 5311 176 5314 204
rect 5280 118 5314 176
rect 5280 90 5283 118
rect 5311 90 5314 118
rect 5280 51 5314 90
rect 5344 290 5378 329
rect 5344 262 5347 290
rect 5375 262 5378 290
rect 5344 204 5378 262
rect 5344 176 5347 204
rect 5375 176 5378 204
rect 5344 118 5378 176
rect 5344 90 5347 118
rect 5375 90 5378 118
rect 5344 51 5378 90
rect 5408 290 5442 329
rect 5408 262 5411 290
rect 5439 262 5442 290
rect 5408 204 5442 262
rect 5408 176 5411 204
rect 5439 176 5442 204
rect 5408 118 5442 176
rect 5408 90 5411 118
rect 5439 90 5442 118
rect 5408 51 5442 90
rect 5472 290 5506 329
rect 5472 262 5475 290
rect 5503 262 5506 290
rect 5472 204 5506 262
rect 5472 176 5475 204
rect 5503 176 5506 204
rect 5472 118 5506 176
rect 5472 90 5475 118
rect 5503 90 5506 118
rect 5472 51 5506 90
rect 5536 290 5570 329
rect 5536 262 5539 290
rect 5567 262 5570 290
rect 5536 204 5570 262
rect 5536 176 5539 204
rect 5567 176 5570 204
rect 5536 118 5570 176
rect 5536 90 5539 118
rect 5567 90 5570 118
rect 5536 51 5570 90
rect 5600 290 5634 329
rect 5600 262 5603 290
rect 5631 262 5634 290
rect 5600 204 5634 262
rect 5600 176 5603 204
rect 5631 176 5634 204
rect 5600 118 5634 176
rect 5600 90 5603 118
rect 5631 90 5634 118
rect 5600 51 5634 90
rect 5664 290 5698 329
rect 5664 262 5667 290
rect 5695 262 5698 290
rect 5664 204 5698 262
rect 5664 176 5667 204
rect 5695 176 5698 204
rect 5664 118 5698 176
rect 5664 90 5667 118
rect 5695 90 5698 118
rect 5664 51 5698 90
rect 5728 290 5762 329
rect 5728 262 5731 290
rect 5759 262 5762 290
rect 5728 204 5762 262
rect 5728 176 5731 204
rect 5759 176 5762 204
rect 5728 118 5762 176
rect 5728 90 5731 118
rect 5759 90 5762 118
rect 5728 51 5762 90
rect 5794 290 5828 329
rect 5794 262 5797 290
rect 5825 262 5828 290
rect 5794 204 5828 262
rect 5794 176 5797 204
rect 5825 176 5828 204
rect 5794 118 5828 176
rect 5794 90 5797 118
rect 5825 90 5828 118
rect 5794 51 5828 90
rect 5858 290 5892 329
rect 5858 262 5861 290
rect 5889 262 5892 290
rect 5858 204 5892 262
rect 5858 176 5861 204
rect 5889 176 5892 204
rect 5858 118 5892 176
rect 5858 90 5861 118
rect 5889 90 5892 118
rect 5858 51 5892 90
rect 5922 290 5956 329
rect 5922 262 5925 290
rect 5953 262 5956 290
rect 5922 204 5956 262
rect 5922 176 5925 204
rect 5953 176 5956 204
rect 5922 118 5956 176
rect 5922 90 5925 118
rect 5953 90 5956 118
rect 5922 51 5956 90
rect 5986 290 6020 329
rect 5986 262 5989 290
rect 6017 262 6020 290
rect 5986 204 6020 262
rect 5986 176 5989 204
rect 6017 176 6020 204
rect 5986 118 6020 176
rect 5986 90 5989 118
rect 6017 90 6020 118
rect 5986 51 6020 90
rect 6050 290 6084 329
rect 6050 262 6053 290
rect 6081 262 6084 290
rect 6050 204 6084 262
rect 6050 176 6053 204
rect 6081 176 6084 204
rect 6050 118 6084 176
rect 6050 90 6053 118
rect 6081 90 6084 118
rect 6050 51 6084 90
rect 6114 290 6148 329
rect 6114 262 6117 290
rect 6145 262 6148 290
rect 6114 204 6148 262
rect 6114 176 6117 204
rect 6145 176 6148 204
rect 6114 118 6148 176
rect 6114 90 6117 118
rect 6145 90 6148 118
rect 6114 51 6148 90
rect 6178 290 6212 329
rect 6178 262 6181 290
rect 6209 262 6212 290
rect 6178 204 6212 262
rect 6178 176 6181 204
rect 6209 176 6212 204
rect 6178 118 6212 176
rect 6178 90 6181 118
rect 6209 90 6212 118
rect 6178 51 6212 90
rect 6242 290 6276 329
rect 6242 262 6245 290
rect 6273 262 6276 290
rect 6242 204 6276 262
rect 6242 176 6245 204
rect 6273 176 6276 204
rect 6242 118 6276 176
rect 6242 90 6245 118
rect 6273 90 6276 118
rect 6242 51 6276 90
rect 6306 290 6340 329
rect 6306 262 6309 290
rect 6337 262 6340 290
rect 6306 204 6340 262
rect 6306 176 6309 204
rect 6337 176 6340 204
rect 6306 118 6340 176
rect 6306 90 6309 118
rect 6337 90 6340 118
rect 6306 51 6340 90
rect 6370 290 6404 329
rect 6370 262 6373 290
rect 6401 262 6404 290
rect 6370 204 6404 262
rect 6370 176 6373 204
rect 6401 176 6404 204
rect 6370 118 6404 176
rect 6370 90 6373 118
rect 6401 90 6404 118
rect 6370 51 6404 90
rect 6436 290 6470 329
rect 6436 262 6439 290
rect 6467 262 6470 290
rect 6436 204 6470 262
rect 6436 176 6439 204
rect 6467 176 6470 204
rect 6436 118 6470 176
rect 6436 90 6439 118
rect 6467 90 6470 118
rect 6436 51 6470 90
rect 6500 290 6534 329
rect 6500 262 6503 290
rect 6531 262 6534 290
rect 6500 204 6534 262
rect 6500 176 6503 204
rect 6531 176 6534 204
rect 6500 118 6534 176
rect 6500 90 6503 118
rect 6531 90 6534 118
rect 6500 51 6534 90
rect 6564 290 6598 329
rect 6564 262 6567 290
rect 6595 262 6598 290
rect 6564 204 6598 262
rect 6564 176 6567 204
rect 6595 176 6598 204
rect 6564 118 6598 176
rect 6564 90 6567 118
rect 6595 90 6598 118
rect 6564 51 6598 90
rect 6628 290 6662 329
rect 6628 262 6631 290
rect 6659 262 6662 290
rect 6628 204 6662 262
rect 6628 176 6631 204
rect 6659 176 6662 204
rect 6628 118 6662 176
rect 6628 90 6631 118
rect 6659 90 6662 118
rect 6628 51 6662 90
rect 6692 290 6726 329
rect 6692 262 6695 290
rect 6723 262 6726 290
rect 6692 204 6726 262
rect 6692 176 6695 204
rect 6723 176 6726 204
rect 6692 118 6726 176
rect 6692 90 6695 118
rect 6723 90 6726 118
rect 6692 51 6726 90
rect 6756 290 6790 329
rect 6756 262 6759 290
rect 6787 262 6790 290
rect 6756 204 6790 262
rect 6756 176 6759 204
rect 6787 176 6790 204
rect 6756 118 6790 176
rect 6756 90 6759 118
rect 6787 90 6790 118
rect 6756 51 6790 90
rect 6820 290 6854 329
rect 6820 262 6823 290
rect 6851 262 6854 290
rect 6820 204 6854 262
rect 6820 176 6823 204
rect 6851 176 6854 204
rect 6820 118 6854 176
rect 6820 90 6823 118
rect 6851 90 6854 118
rect 6820 51 6854 90
rect 6884 290 6918 329
rect 6884 262 6887 290
rect 6915 262 6918 290
rect 6884 204 6918 262
rect 6884 176 6887 204
rect 6915 176 6918 204
rect 6884 118 6918 176
rect 6884 90 6887 118
rect 6915 90 6918 118
rect 6884 51 6918 90
rect 6948 290 6982 329
rect 6948 262 6951 290
rect 6979 262 6982 290
rect 6948 204 6982 262
rect 6948 176 6951 204
rect 6979 176 6982 204
rect 6948 118 6982 176
rect 6948 90 6951 118
rect 6979 90 6982 118
rect 6948 51 6982 90
rect 7012 290 7046 329
rect 7012 262 7015 290
rect 7043 262 7046 290
rect 7012 204 7046 262
rect 7012 176 7015 204
rect 7043 176 7046 204
rect 7012 118 7046 176
rect 7012 90 7015 118
rect 7043 90 7046 118
rect 7012 51 7046 90
rect 7078 290 7112 329
rect 7078 262 7081 290
rect 7109 262 7112 290
rect 7078 204 7112 262
rect 7078 176 7081 204
rect 7109 176 7112 204
rect 7078 118 7112 176
rect 7078 90 7081 118
rect 7109 90 7112 118
rect 7078 51 7112 90
rect 7142 290 7176 329
rect 7142 262 7145 290
rect 7173 262 7176 290
rect 7142 204 7176 262
rect 7142 176 7145 204
rect 7173 176 7176 204
rect 7142 118 7176 176
rect 7142 90 7145 118
rect 7173 90 7176 118
rect 7142 51 7176 90
rect 7206 290 7240 329
rect 7206 262 7209 290
rect 7237 262 7240 290
rect 7206 204 7240 262
rect 7206 176 7209 204
rect 7237 176 7240 204
rect 7206 118 7240 176
rect 7206 90 7209 118
rect 7237 90 7240 118
rect 7206 51 7240 90
rect 7270 290 7304 329
rect 7270 262 7273 290
rect 7301 262 7304 290
rect 7270 204 7304 262
rect 7270 176 7273 204
rect 7301 176 7304 204
rect 7270 118 7304 176
rect 7270 90 7273 118
rect 7301 90 7304 118
rect 7270 51 7304 90
rect 7334 290 7368 329
rect 7334 262 7337 290
rect 7365 262 7368 290
rect 7334 204 7368 262
rect 7334 176 7337 204
rect 7365 176 7368 204
rect 7334 118 7368 176
rect 7334 90 7337 118
rect 7365 90 7368 118
rect 7334 51 7368 90
rect 7398 290 7432 329
rect 7398 262 7401 290
rect 7429 262 7432 290
rect 7398 204 7432 262
rect 7398 176 7401 204
rect 7429 176 7432 204
rect 7398 118 7432 176
rect 7398 90 7401 118
rect 7429 90 7432 118
rect 7398 51 7432 90
rect 7462 290 7496 329
rect 7462 262 7465 290
rect 7493 262 7496 290
rect 7462 204 7496 262
rect 7462 176 7465 204
rect 7493 176 7496 204
rect 7462 118 7496 176
rect 7462 90 7465 118
rect 7493 90 7496 118
rect 7462 51 7496 90
rect 7526 290 7560 329
rect 7526 262 7529 290
rect 7557 262 7560 290
rect 7526 204 7560 262
rect 7526 176 7529 204
rect 7557 176 7560 204
rect 7526 118 7560 176
rect 7526 90 7529 118
rect 7557 90 7560 118
rect 7526 51 7560 90
rect 7590 290 7624 329
rect 7590 262 7593 290
rect 7621 262 7624 290
rect 7590 204 7624 262
rect 7590 176 7593 204
rect 7621 176 7624 204
rect 7590 118 7624 176
rect 7590 90 7593 118
rect 7621 90 7624 118
rect 7590 51 7624 90
rect 7654 290 7688 329
rect 7654 262 7657 290
rect 7685 262 7688 290
rect 7654 204 7688 262
rect 7654 176 7657 204
rect 7685 176 7688 204
rect 7654 118 7688 176
rect 7654 90 7657 118
rect 7685 90 7688 118
rect 7654 51 7688 90
rect 7720 290 7754 329
rect 7720 262 7723 290
rect 7751 262 7754 290
rect 7720 204 7754 262
rect 7720 176 7723 204
rect 7751 176 7754 204
rect 7720 118 7754 176
rect 7720 90 7723 118
rect 7751 90 7754 118
rect 7720 51 7754 90
rect 7784 290 7818 329
rect 7784 262 7787 290
rect 7815 262 7818 290
rect 7784 204 7818 262
rect 7784 176 7787 204
rect 7815 176 7818 204
rect 7784 118 7818 176
rect 7784 90 7787 118
rect 7815 90 7818 118
rect 7784 51 7818 90
rect 7848 290 7882 329
rect 7848 262 7851 290
rect 7879 262 7882 290
rect 7848 204 7882 262
rect 7848 176 7851 204
rect 7879 176 7882 204
rect 7848 118 7882 176
rect 7848 90 7851 118
rect 7879 90 7882 118
rect 7848 51 7882 90
rect 7912 290 7946 329
rect 7912 262 7915 290
rect 7943 262 7946 290
rect 7912 204 7946 262
rect 7912 176 7915 204
rect 7943 176 7946 204
rect 7912 118 7946 176
rect 7912 90 7915 118
rect 7943 90 7946 118
rect 7912 51 7946 90
rect 7976 290 8010 329
rect 7976 262 7979 290
rect 8007 262 8010 290
rect 7976 204 8010 262
rect 7976 176 7979 204
rect 8007 176 8010 204
rect 7976 118 8010 176
rect 7976 90 7979 118
rect 8007 90 8010 118
rect 7976 51 8010 90
rect 8040 290 8074 329
rect 8040 262 8043 290
rect 8071 262 8074 290
rect 8040 204 8074 262
rect 8040 176 8043 204
rect 8071 176 8074 204
rect 8040 118 8074 176
rect 8040 90 8043 118
rect 8071 90 8074 118
rect 8040 51 8074 90
rect 8104 290 8138 329
rect 8104 262 8107 290
rect 8135 262 8138 290
rect 8104 204 8138 262
rect 8104 176 8107 204
rect 8135 176 8138 204
rect 8104 118 8138 176
rect 8104 90 8107 118
rect 8135 90 8138 118
rect 8104 51 8138 90
rect 8168 290 8202 329
rect 8168 262 8171 290
rect 8199 262 8202 290
rect 8168 204 8202 262
rect 8168 176 8171 204
rect 8199 176 8202 204
rect 8168 118 8202 176
rect 8168 90 8171 118
rect 8199 90 8202 118
rect 8168 51 8202 90
rect 8232 290 8266 329
rect 8232 262 8235 290
rect 8263 262 8266 290
rect 8232 204 8266 262
rect 8232 176 8235 204
rect 8263 176 8266 204
rect 8232 118 8266 176
rect 8232 90 8235 118
rect 8263 90 8266 118
rect 8232 51 8266 90
rect 8296 290 8330 329
rect 8296 262 8299 290
rect 8327 262 8330 290
rect 8296 204 8330 262
rect 8296 176 8299 204
rect 8327 176 8330 204
rect 8296 118 8330 176
rect 8296 90 8299 118
rect 8327 90 8330 118
rect 8296 51 8330 90
rect 8362 290 8396 329
rect 8362 262 8365 290
rect 8393 262 8396 290
rect 8362 204 8396 262
rect 8362 176 8365 204
rect 8393 176 8396 204
rect 8362 118 8396 176
rect 8362 90 8365 118
rect 8393 90 8396 118
rect 8362 51 8396 90
rect 8426 290 8460 329
rect 8426 262 8429 290
rect 8457 262 8460 290
rect 8426 204 8460 262
rect 8426 176 8429 204
rect 8457 176 8460 204
rect 8426 118 8460 176
rect 8426 90 8429 118
rect 8457 90 8460 118
rect 8426 51 8460 90
rect 8490 290 8524 329
rect 8490 262 8493 290
rect 8521 262 8524 290
rect 8490 204 8524 262
rect 8490 176 8493 204
rect 8521 176 8524 204
rect 8490 118 8524 176
rect 8490 90 8493 118
rect 8521 90 8524 118
rect 8490 51 8524 90
rect 8554 290 8588 329
rect 8554 262 8557 290
rect 8585 262 8588 290
rect 8554 204 8588 262
rect 8554 176 8557 204
rect 8585 176 8588 204
rect 8554 118 8588 176
rect 8554 90 8557 118
rect 8585 90 8588 118
rect 8554 51 8588 90
rect 8618 290 8652 329
rect 8618 262 8621 290
rect 8649 262 8652 290
rect 8618 204 8652 262
rect 8618 176 8621 204
rect 8649 176 8652 204
rect 8618 118 8652 176
rect 8618 90 8621 118
rect 8649 90 8652 118
rect 8618 51 8652 90
rect 8682 290 8716 329
rect 8682 262 8685 290
rect 8713 262 8716 290
rect 8682 204 8716 262
rect 8682 176 8685 204
rect 8713 176 8716 204
rect 8682 118 8716 176
rect 8682 90 8685 118
rect 8713 90 8716 118
rect 8682 51 8716 90
rect 8746 290 8780 329
rect 8746 262 8749 290
rect 8777 262 8780 290
rect 8746 204 8780 262
rect 8746 176 8749 204
rect 8777 176 8780 204
rect 8746 118 8780 176
rect 8746 90 8749 118
rect 8777 90 8780 118
rect 8746 51 8780 90
rect 8810 290 8844 329
rect 8810 262 8813 290
rect 8841 262 8844 290
rect 8810 204 8844 262
rect 8810 176 8813 204
rect 8841 176 8844 204
rect 8810 118 8844 176
rect 8810 90 8813 118
rect 8841 90 8844 118
rect 8810 51 8844 90
rect 8874 290 8908 329
rect 8874 262 8877 290
rect 8905 262 8908 290
rect 8874 204 8908 262
rect 8874 176 8877 204
rect 8905 176 8908 204
rect 8874 118 8908 176
rect 8874 90 8877 118
rect 8905 90 8908 118
rect 8874 51 8908 90
rect 8938 290 8972 329
rect 8938 262 8941 290
rect 8969 262 8972 290
rect 8938 204 8972 262
rect 8938 176 8941 204
rect 8969 176 8972 204
rect 8938 118 8972 176
rect 8938 90 8941 118
rect 8969 90 8972 118
rect 8938 51 8972 90
rect 9004 290 9038 329
rect 9004 262 9007 290
rect 9035 262 9038 290
rect 9004 204 9038 262
rect 9004 176 9007 204
rect 9035 176 9038 204
rect 9004 118 9038 176
rect 9004 90 9007 118
rect 9035 90 9038 118
rect 9004 51 9038 90
rect 9068 290 9102 329
rect 9068 262 9071 290
rect 9099 262 9102 290
rect 9068 204 9102 262
rect 9068 176 9071 204
rect 9099 176 9102 204
rect 9068 118 9102 176
rect 9068 90 9071 118
rect 9099 90 9102 118
rect 9068 51 9102 90
rect 9132 290 9166 329
rect 9132 262 9135 290
rect 9163 262 9166 290
rect 9132 204 9166 262
rect 9132 176 9135 204
rect 9163 176 9166 204
rect 9132 118 9166 176
rect 9132 90 9135 118
rect 9163 90 9166 118
rect 9132 51 9166 90
rect 9196 290 9230 329
rect 9196 262 9199 290
rect 9227 262 9230 290
rect 9196 204 9230 262
rect 9196 176 9199 204
rect 9227 176 9230 204
rect 9196 118 9230 176
rect 9196 90 9199 118
rect 9227 90 9230 118
rect 9196 51 9230 90
rect 9260 290 9294 329
rect 9260 262 9263 290
rect 9291 262 9294 290
rect 9260 204 9294 262
rect 9260 176 9263 204
rect 9291 176 9294 204
rect 9260 118 9294 176
rect 9260 90 9263 118
rect 9291 90 9294 118
rect 9260 51 9294 90
rect 9324 290 9358 329
rect 9324 262 9327 290
rect 9355 262 9358 290
rect 9324 204 9358 262
rect 9324 176 9327 204
rect 9355 176 9358 204
rect 9324 118 9358 176
rect 9324 90 9327 118
rect 9355 90 9358 118
rect 9324 51 9358 90
rect 9388 290 9422 329
rect 9388 262 9391 290
rect 9419 262 9422 290
rect 9388 204 9422 262
rect 9388 176 9391 204
rect 9419 176 9422 204
rect 9388 118 9422 176
rect 9388 90 9391 118
rect 9419 90 9422 118
rect 9388 51 9422 90
rect 9452 290 9486 329
rect 9452 262 9455 290
rect 9483 262 9486 290
rect 9452 204 9486 262
rect 9452 176 9455 204
rect 9483 176 9486 204
rect 9452 118 9486 176
rect 9452 90 9455 118
rect 9483 90 9486 118
rect 9452 51 9486 90
rect 9516 290 9550 329
rect 9516 262 9519 290
rect 9547 262 9550 290
rect 9516 204 9550 262
rect 9516 176 9519 204
rect 9547 176 9550 204
rect 9516 118 9550 176
rect 9516 90 9519 118
rect 9547 90 9550 118
rect 9516 51 9550 90
rect 9580 290 9614 329
rect 9580 262 9583 290
rect 9611 262 9614 290
rect 9580 204 9614 262
rect 9580 176 9583 204
rect 9611 176 9614 204
rect 9580 118 9614 176
rect 9580 90 9583 118
rect 9611 90 9614 118
rect 9580 51 9614 90
rect 9646 290 9680 329
rect 9646 262 9649 290
rect 9677 262 9680 290
rect 9646 204 9680 262
rect 9646 176 9649 204
rect 9677 176 9680 204
rect 9646 118 9680 176
rect 9646 90 9649 118
rect 9677 90 9680 118
rect 9646 51 9680 90
rect 9710 290 9744 329
rect 9710 262 9713 290
rect 9741 262 9744 290
rect 9710 204 9744 262
rect 9710 176 9713 204
rect 9741 176 9744 204
rect 9710 118 9744 176
rect 9710 90 9713 118
rect 9741 90 9744 118
rect 9710 51 9744 90
rect 9774 290 9808 329
rect 9774 262 9777 290
rect 9805 262 9808 290
rect 9774 204 9808 262
rect 9774 176 9777 204
rect 9805 176 9808 204
rect 9774 118 9808 176
rect 9774 90 9777 118
rect 9805 90 9808 118
rect 9774 51 9808 90
rect 9838 290 9872 329
rect 9838 262 9841 290
rect 9869 262 9872 290
rect 9838 204 9872 262
rect 9838 176 9841 204
rect 9869 176 9872 204
rect 9838 118 9872 176
rect 9838 90 9841 118
rect 9869 90 9872 118
rect 9838 51 9872 90
rect 9902 290 9936 329
rect 9902 262 9905 290
rect 9933 262 9936 290
rect 9902 204 9936 262
rect 9902 176 9905 204
rect 9933 176 9936 204
rect 9902 118 9936 176
rect 9902 90 9905 118
rect 9933 90 9936 118
rect 9902 51 9936 90
rect 9966 290 10000 329
rect 9966 262 9969 290
rect 9997 262 10000 290
rect 9966 204 10000 262
rect 9966 176 9969 204
rect 9997 176 10000 204
rect 9966 118 10000 176
rect 9966 90 9969 118
rect 9997 90 10000 118
rect 9966 51 10000 90
rect 10030 290 10064 329
rect 10030 262 10033 290
rect 10061 262 10064 290
rect 10030 204 10064 262
rect 10030 176 10033 204
rect 10061 176 10064 204
rect 10030 118 10064 176
rect 10030 90 10033 118
rect 10061 90 10064 118
rect 10030 51 10064 90
rect 10094 290 10128 329
rect 10094 262 10097 290
rect 10125 262 10128 290
rect 10094 204 10128 262
rect 10094 176 10097 204
rect 10125 176 10128 204
rect 10094 118 10128 176
rect 10094 90 10097 118
rect 10125 90 10128 118
rect 10094 51 10128 90
rect 10158 290 10192 329
rect 10158 262 10161 290
rect 10189 262 10192 290
rect 10158 204 10192 262
rect 10158 176 10161 204
rect 10189 176 10192 204
rect 10158 118 10192 176
rect 10158 90 10161 118
rect 10189 90 10192 118
rect 10158 51 10192 90
rect 10222 290 10256 329
rect 10222 262 10225 290
rect 10253 262 10256 290
rect 10222 204 10256 262
rect 10222 176 10225 204
rect 10253 176 10256 204
rect 10222 118 10256 176
rect 10222 90 10225 118
rect 10253 90 10256 118
rect 10222 51 10256 90
rect 10288 290 10322 329
rect 10288 262 10291 290
rect 10319 262 10322 290
rect 10288 204 10322 262
rect 10288 176 10291 204
rect 10319 176 10322 204
rect 10288 118 10322 176
rect 10288 90 10291 118
rect 10319 90 10322 118
rect 10288 51 10322 90
rect 10352 290 10386 329
rect 10352 262 10355 290
rect 10383 262 10386 290
rect 10352 204 10386 262
rect 10352 176 10355 204
rect 10383 176 10386 204
rect 10352 118 10386 176
rect 10352 90 10355 118
rect 10383 90 10386 118
rect 10352 51 10386 90
rect 10416 290 10450 329
rect 10416 262 10419 290
rect 10447 262 10450 290
rect 10416 204 10450 262
rect 10416 176 10419 204
rect 10447 176 10450 204
rect 10416 118 10450 176
rect 10416 90 10419 118
rect 10447 90 10450 118
rect 10416 51 10450 90
rect 10480 290 10514 329
rect 10480 262 10483 290
rect 10511 262 10514 290
rect 10480 204 10514 262
rect 10480 176 10483 204
rect 10511 176 10514 204
rect 10480 118 10514 176
rect 10480 90 10483 118
rect 10511 90 10514 118
rect 10480 51 10514 90
rect 10544 290 10578 329
rect 10544 262 10547 290
rect 10575 262 10578 290
rect 10544 204 10578 262
rect 10544 176 10547 204
rect 10575 176 10578 204
rect 10544 118 10578 176
rect 10544 90 10547 118
rect 10575 90 10578 118
rect 10544 51 10578 90
rect 10608 290 10642 329
rect 10608 262 10611 290
rect 10639 262 10642 290
rect 10608 204 10642 262
rect 10608 176 10611 204
rect 10639 176 10642 204
rect 10608 118 10642 176
rect 10608 90 10611 118
rect 10639 90 10642 118
rect 10608 51 10642 90
rect 10672 290 10706 329
rect 10672 262 10675 290
rect 10703 262 10706 290
rect 10672 204 10706 262
rect 10672 176 10675 204
rect 10703 176 10706 204
rect 10672 118 10706 176
rect 10672 90 10675 118
rect 10703 90 10706 118
rect 10672 51 10706 90
rect 10736 290 10770 329
rect 10736 262 10739 290
rect 10767 262 10770 290
rect 10736 204 10770 262
rect 10736 176 10739 204
rect 10767 176 10770 204
rect 10736 118 10770 176
rect 10736 90 10739 118
rect 10767 90 10770 118
rect 10736 51 10770 90
rect 10800 290 10834 329
rect 10800 262 10803 290
rect 10831 262 10834 290
rect 10800 204 10834 262
rect 10800 176 10803 204
rect 10831 176 10834 204
rect 10800 118 10834 176
rect 10800 90 10803 118
rect 10831 90 10834 118
rect 10800 51 10834 90
rect 10864 290 10898 329
rect 10864 262 10867 290
rect 10895 262 10898 290
rect 10864 204 10898 262
rect 10864 176 10867 204
rect 10895 176 10898 204
rect 10864 118 10898 176
rect 10864 90 10867 118
rect 10895 90 10898 118
rect 10864 51 10898 90
rect 10930 290 10964 329
rect 10930 262 10933 290
rect 10961 262 10964 290
rect 10930 204 10964 262
rect 10930 176 10933 204
rect 10961 176 10964 204
rect 10930 118 10964 176
rect 10930 90 10933 118
rect 10961 90 10964 118
rect 10930 51 10964 90
rect 10994 290 11028 329
rect 10994 262 10997 290
rect 11025 262 11028 290
rect 10994 204 11028 262
rect 10994 176 10997 204
rect 11025 176 11028 204
rect 10994 118 11028 176
rect 10994 90 10997 118
rect 11025 90 11028 118
rect 10994 51 11028 90
rect 11058 290 11092 329
rect 11058 262 11061 290
rect 11089 262 11092 290
rect 11058 204 11092 262
rect 11058 176 11061 204
rect 11089 176 11092 204
rect 11058 118 11092 176
rect 11058 90 11061 118
rect 11089 90 11092 118
rect 11058 51 11092 90
rect 11122 290 11156 329
rect 11122 262 11125 290
rect 11153 262 11156 290
rect 11122 204 11156 262
rect 11122 176 11125 204
rect 11153 176 11156 204
rect 11122 118 11156 176
rect 11122 90 11125 118
rect 11153 90 11156 118
rect 11122 51 11156 90
rect 11186 290 11220 329
rect 11186 262 11189 290
rect 11217 262 11220 290
rect 11186 204 11220 262
rect 11186 176 11189 204
rect 11217 176 11220 204
rect 11186 118 11220 176
rect 11186 90 11189 118
rect 11217 90 11220 118
rect 11186 51 11220 90
rect 11250 290 11284 329
rect 11250 262 11253 290
rect 11281 262 11284 290
rect 11250 204 11284 262
rect 11250 176 11253 204
rect 11281 176 11284 204
rect 11250 118 11284 176
rect 11250 90 11253 118
rect 11281 90 11284 118
rect 11250 51 11284 90
rect 11314 290 11348 329
rect 11314 262 11317 290
rect 11345 262 11348 290
rect 11314 204 11348 262
rect 11314 176 11317 204
rect 11345 176 11348 204
rect 11314 118 11348 176
rect 11314 90 11317 118
rect 11345 90 11348 118
rect 11314 51 11348 90
rect 11378 290 11412 329
rect 11378 262 11381 290
rect 11409 262 11412 290
rect 11378 204 11412 262
rect 11378 176 11381 204
rect 11409 176 11412 204
rect 11378 118 11412 176
rect 11378 90 11381 118
rect 11409 90 11412 118
rect 11378 51 11412 90
rect 11442 290 11476 329
rect 11442 262 11445 290
rect 11473 262 11476 290
rect 11442 204 11476 262
rect 11442 176 11445 204
rect 11473 176 11476 204
rect 11442 118 11476 176
rect 11442 90 11445 118
rect 11473 90 11476 118
rect 11442 51 11476 90
rect 11506 290 11540 329
rect 11506 262 11509 290
rect 11537 262 11540 290
rect 11506 204 11540 262
rect 11506 176 11509 204
rect 11537 176 11540 204
rect 11506 118 11540 176
rect 11506 90 11509 118
rect 11537 90 11540 118
rect 11506 51 11540 90
rect 11572 290 11606 329
rect 11572 262 11575 290
rect 11603 262 11606 290
rect 11572 204 11606 262
rect 11572 176 11575 204
rect 11603 176 11606 204
rect 11572 118 11606 176
rect 11572 90 11575 118
rect 11603 90 11606 118
rect 11572 51 11606 90
rect 11636 290 11670 329
rect 11636 262 11639 290
rect 11667 262 11670 290
rect 11636 204 11670 262
rect 11636 176 11639 204
rect 11667 176 11670 204
rect 11636 118 11670 176
rect 11636 90 11639 118
rect 11667 90 11670 118
rect 11636 51 11670 90
rect 11700 290 11734 329
rect 11700 262 11703 290
rect 11731 262 11734 290
rect 11700 204 11734 262
rect 11700 176 11703 204
rect 11731 176 11734 204
rect 11700 118 11734 176
rect 11700 90 11703 118
rect 11731 90 11734 118
rect 11700 51 11734 90
rect 11764 290 11798 329
rect 11764 262 11767 290
rect 11795 262 11798 290
rect 11764 204 11798 262
rect 11764 176 11767 204
rect 11795 176 11798 204
rect 11764 118 11798 176
rect 11764 90 11767 118
rect 11795 90 11798 118
rect 11764 51 11798 90
rect 11828 290 11862 329
rect 11828 262 11831 290
rect 11859 262 11862 290
rect 11828 204 11862 262
rect 11828 176 11831 204
rect 11859 176 11862 204
rect 11828 118 11862 176
rect 11828 90 11831 118
rect 11859 90 11862 118
rect 11828 51 11862 90
rect 11892 290 11926 329
rect 11892 262 11895 290
rect 11923 262 11926 290
rect 11892 204 11926 262
rect 11892 176 11895 204
rect 11923 176 11926 204
rect 11892 118 11926 176
rect 11892 90 11895 118
rect 11923 90 11926 118
rect 11892 51 11926 90
rect 11956 290 11990 329
rect 11956 262 11959 290
rect 11987 262 11990 290
rect 11956 204 11990 262
rect 11956 176 11959 204
rect 11987 176 11990 204
rect 11956 118 11990 176
rect 11956 90 11959 118
rect 11987 90 11990 118
rect 11956 51 11990 90
rect 12020 290 12054 329
rect 12020 262 12023 290
rect 12051 262 12054 290
rect 12020 204 12054 262
rect 12020 176 12023 204
rect 12051 176 12054 204
rect 12020 118 12054 176
rect 12020 90 12023 118
rect 12051 90 12054 118
rect 12020 51 12054 90
rect 12084 290 12118 329
rect 12084 262 12087 290
rect 12115 262 12118 290
rect 12084 204 12118 262
rect 12084 176 12087 204
rect 12115 176 12118 204
rect 12084 118 12118 176
rect 12084 90 12087 118
rect 12115 90 12118 118
rect 12084 51 12118 90
rect 12148 290 12182 329
rect 12148 262 12151 290
rect 12179 262 12182 290
rect 12148 204 12182 262
rect 12148 176 12151 204
rect 12179 176 12182 204
rect 12148 118 12182 176
rect 12148 90 12151 118
rect 12179 90 12182 118
rect 12148 51 12182 90
rect 12214 290 12248 329
rect 12214 262 12217 290
rect 12245 262 12248 290
rect 12214 204 12248 262
rect 12214 176 12217 204
rect 12245 176 12248 204
rect 12214 118 12248 176
rect 12214 90 12217 118
rect 12245 90 12248 118
rect 12214 51 12248 90
rect 12278 290 12312 329
rect 12278 262 12281 290
rect 12309 262 12312 290
rect 12278 204 12312 262
rect 12278 176 12281 204
rect 12309 176 12312 204
rect 12278 118 12312 176
rect 12278 90 12281 118
rect 12309 90 12312 118
rect 12278 51 12312 90
rect 12342 290 12376 329
rect 12342 262 12345 290
rect 12373 262 12376 290
rect 12342 204 12376 262
rect 12342 176 12345 204
rect 12373 176 12376 204
rect 12342 118 12376 176
rect 12342 90 12345 118
rect 12373 90 12376 118
rect 12342 51 12376 90
rect 12406 290 12440 329
rect 12406 262 12409 290
rect 12437 262 12440 290
rect 12406 204 12440 262
rect 12406 176 12409 204
rect 12437 176 12440 204
rect 12406 118 12440 176
rect 12406 90 12409 118
rect 12437 90 12440 118
rect 12406 51 12440 90
rect 12470 290 12504 329
rect 12470 262 12473 290
rect 12501 262 12504 290
rect 12470 204 12504 262
rect 12470 176 12473 204
rect 12501 176 12504 204
rect 12470 118 12504 176
rect 12470 90 12473 118
rect 12501 90 12504 118
rect 12470 51 12504 90
rect 12534 290 12568 329
rect 12534 262 12537 290
rect 12565 262 12568 290
rect 12534 204 12568 262
rect 12534 176 12537 204
rect 12565 176 12568 204
rect 12534 118 12568 176
rect 12534 90 12537 118
rect 12565 90 12568 118
rect 12534 51 12568 90
rect 12598 290 12632 329
rect 12598 262 12601 290
rect 12629 262 12632 290
rect 12598 204 12632 262
rect 12598 176 12601 204
rect 12629 176 12632 204
rect 12598 118 12632 176
rect 12598 90 12601 118
rect 12629 90 12632 118
rect 12598 51 12632 90
rect 12662 290 12696 329
rect 12662 262 12665 290
rect 12693 262 12696 290
rect 12662 204 12696 262
rect 12662 176 12665 204
rect 12693 176 12696 204
rect 12662 118 12696 176
rect 12662 90 12665 118
rect 12693 90 12696 118
rect 12662 51 12696 90
rect 12726 290 12760 329
rect 12726 262 12729 290
rect 12757 262 12760 290
rect 12726 204 12760 262
rect 12726 176 12729 204
rect 12757 176 12760 204
rect 12726 118 12760 176
rect 12726 90 12729 118
rect 12757 90 12760 118
rect 12726 51 12760 90
rect 12790 290 12824 329
rect 12790 262 12793 290
rect 12821 262 12824 290
rect 12790 204 12824 262
rect 12790 176 12793 204
rect 12821 176 12824 204
rect 12790 118 12824 176
rect 12790 90 12793 118
rect 12821 90 12824 118
rect 12790 51 12824 90
<< metal4 >>
rect 0 1505 12840 1535
rect 18 1185 48 1475
rect 82 1155 112 1505
rect 146 1155 176 1505
rect 210 1155 240 1505
rect 274 1155 304 1505
rect 338 1155 368 1505
rect 402 1155 432 1505
rect 466 1155 496 1505
rect 530 1155 560 1505
rect 594 1185 624 1475
rect 660 1185 690 1475
rect 724 1185 754 1505
rect 788 1185 818 1505
rect 852 1185 882 1505
rect 916 1185 946 1505
rect 980 1185 1010 1505
rect 1044 1185 1074 1505
rect 1108 1185 1138 1505
rect 1172 1185 1202 1505
rect 1236 1185 1266 1475
rect 1302 1185 1332 1475
rect 1366 1185 1396 1505
rect 1430 1185 1460 1505
rect 1494 1185 1524 1505
rect 1558 1185 1588 1505
rect 1622 1185 1652 1505
rect 1686 1185 1716 1505
rect 1750 1185 1780 1505
rect 1814 1185 1844 1505
rect 1878 1185 1908 1475
rect 1944 1185 1974 1475
rect 2008 1185 2038 1505
rect 2072 1185 2102 1505
rect 2136 1185 2166 1505
rect 2200 1185 2230 1505
rect 2264 1185 2294 1505
rect 2328 1185 2358 1505
rect 2392 1185 2422 1505
rect 2456 1185 2486 1505
rect 2520 1185 2550 1475
rect 2586 1185 2616 1475
rect 2650 1155 2680 1505
rect 2714 1155 2744 1505
rect 2778 1155 2808 1505
rect 2842 1155 2872 1505
rect 2906 1155 2936 1505
rect 2970 1155 3000 1505
rect 3034 1155 3064 1505
rect 3098 1155 3128 1505
rect 3162 1185 3192 1475
rect 3228 1185 3258 1475
rect 3292 1155 3322 1505
rect 3356 1155 3386 1505
rect 3420 1155 3450 1505
rect 3484 1155 3514 1505
rect 3548 1155 3578 1505
rect 3612 1155 3642 1505
rect 3676 1155 3706 1505
rect 3740 1155 3770 1505
rect 3804 1185 3834 1475
rect 3870 1185 3900 1475
rect 3934 1186 3964 1505
rect 3998 1186 4028 1505
rect 4062 1186 4092 1505
rect 4126 1186 4156 1505
rect 4190 1186 4220 1505
rect 4254 1186 4284 1505
rect 4318 1186 4348 1505
rect 4382 1186 4412 1505
rect 4446 1186 4476 1475
rect 4512 1186 4542 1475
rect 4576 1186 4606 1505
rect 4640 1186 4670 1505
rect 4704 1186 4734 1505
rect 4768 1186 4798 1505
rect 4832 1186 4862 1505
rect 4896 1186 4926 1505
rect 4960 1186 4990 1505
rect 5024 1186 5054 1505
rect 5088 1186 5118 1475
rect 5154 1186 5184 1475
rect 5218 1186 5248 1505
rect 5282 1186 5312 1505
rect 5346 1186 5376 1505
rect 5410 1186 5440 1505
rect 5474 1186 5504 1505
rect 5538 1186 5568 1505
rect 5602 1186 5632 1505
rect 5666 1186 5696 1505
rect 5730 1185 5760 1475
rect 5796 1185 5826 1475
rect 3934 1155 3964 1156
rect 3998 1155 4028 1156
rect 4062 1155 4092 1156
rect 4126 1155 4156 1156
rect 4190 1155 4220 1156
rect 4254 1155 4284 1156
rect 4318 1155 4348 1156
rect 4382 1155 4412 1156
rect 4576 1155 4606 1156
rect 4640 1155 4670 1156
rect 4704 1155 4734 1156
rect 4768 1155 4798 1156
rect 4832 1155 4862 1156
rect 4896 1155 4926 1156
rect 4960 1155 4990 1156
rect 5024 1155 5054 1156
rect 5218 1155 5248 1156
rect 5282 1155 5312 1156
rect 5346 1155 5376 1156
rect 5410 1155 5440 1156
rect 5474 1155 5504 1156
rect 5538 1155 5568 1156
rect 5602 1155 5632 1156
rect 5666 1155 5696 1156
rect 5860 1155 5890 1505
rect 5924 1155 5954 1505
rect 5988 1155 6018 1505
rect 6052 1155 6082 1505
rect 6116 1155 6146 1505
rect 6180 1155 6210 1505
rect 6244 1155 6274 1505
rect 6308 1155 6338 1505
rect 6372 1185 6402 1475
rect 6438 1185 6468 1475
rect 6502 1155 6532 1505
rect 6566 1155 6596 1505
rect 6630 1155 6660 1505
rect 6694 1155 6724 1505
rect 6758 1155 6788 1505
rect 6822 1155 6852 1505
rect 6886 1155 6916 1505
rect 6950 1155 6980 1505
rect 7014 1185 7044 1475
rect 7080 1185 7110 1475
rect 7144 1185 7174 1505
rect 7208 1185 7238 1505
rect 7272 1185 7302 1505
rect 7336 1185 7366 1505
rect 7400 1185 7430 1505
rect 7464 1185 7494 1505
rect 7528 1185 7558 1505
rect 7592 1185 7622 1505
rect 7656 1185 7686 1475
rect 7722 1185 7752 1475
rect 7786 1185 7816 1505
rect 7850 1185 7880 1505
rect 7914 1185 7944 1505
rect 7978 1185 8008 1505
rect 8042 1185 8072 1505
rect 8106 1185 8136 1505
rect 8170 1185 8200 1505
rect 8234 1185 8264 1505
rect 8298 1185 8328 1475
rect 8364 1185 8394 1475
rect 8428 1185 8458 1505
rect 8492 1185 8522 1505
rect 8556 1185 8586 1505
rect 8620 1185 8650 1505
rect 8684 1185 8714 1505
rect 8748 1185 8778 1505
rect 8812 1185 8842 1505
rect 8876 1185 8906 1505
rect 8940 1185 8970 1475
rect 9006 1185 9036 1475
rect 9070 1155 9100 1505
rect 9134 1155 9164 1505
rect 9198 1155 9228 1505
rect 9262 1155 9292 1505
rect 9326 1155 9356 1505
rect 9390 1155 9420 1505
rect 9454 1155 9484 1505
rect 9518 1155 9548 1505
rect 9582 1185 9612 1475
rect 9648 1185 9678 1475
rect 9712 1155 9742 1505
rect 9776 1155 9806 1505
rect 9840 1155 9870 1505
rect 9904 1155 9934 1505
rect 9968 1155 9998 1505
rect 10032 1155 10062 1505
rect 10096 1155 10126 1505
rect 10160 1155 10190 1505
rect 10224 1185 10254 1475
rect 10290 1185 10320 1475
rect 10354 1185 10384 1505
rect 10418 1185 10448 1505
rect 10482 1185 10512 1505
rect 10546 1185 10576 1505
rect 10610 1185 10640 1505
rect 10674 1185 10704 1505
rect 10738 1185 10768 1505
rect 10802 1185 10832 1505
rect 10866 1185 10896 1475
rect 10932 1185 10962 1475
rect 10996 1185 11026 1505
rect 11060 1185 11090 1505
rect 11124 1185 11154 1505
rect 11188 1185 11218 1505
rect 11252 1185 11282 1505
rect 11316 1185 11346 1505
rect 11380 1185 11410 1505
rect 11444 1185 11474 1505
rect 11508 1185 11538 1475
rect 11574 1185 11604 1475
rect 11638 1185 11668 1505
rect 11702 1185 11732 1505
rect 11766 1185 11796 1505
rect 11830 1185 11860 1505
rect 11894 1185 11924 1505
rect 11958 1185 11988 1505
rect 12022 1185 12052 1505
rect 12086 1185 12116 1505
rect 12150 1185 12180 1475
rect 12216 1185 12246 1475
rect 12280 1155 12310 1505
rect 12344 1155 12374 1505
rect 12408 1155 12438 1505
rect 12472 1155 12502 1505
rect 12536 1155 12566 1505
rect 12600 1155 12630 1505
rect 12664 1155 12694 1505
rect 12728 1155 12758 1505
rect 12792 1185 12822 1475
rect 0 1125 625 1155
rect 659 1125 2551 1155
rect 2585 1125 3835 1155
rect 3869 1125 5761 1155
rect 5795 1125 7045 1155
rect 7079 1125 8971 1155
rect 9005 1125 10255 1155
rect 10289 1125 12181 1155
rect 12215 1125 12840 1155
rect 18 805 48 1095
rect 82 775 112 1125
rect 146 775 176 1125
rect 210 775 240 1125
rect 274 775 304 1125
rect 338 775 368 1125
rect 402 775 432 1125
rect 466 775 496 1125
rect 530 775 560 1125
rect 594 805 624 1095
rect 660 805 690 1095
rect 724 775 754 1125
rect 788 775 818 1125
rect 852 775 882 1125
rect 916 775 946 1125
rect 980 775 1010 1125
rect 1044 775 1074 1125
rect 1108 775 1138 1125
rect 1172 775 1202 1125
rect 1236 805 1266 1095
rect 1302 805 1332 1095
rect 1366 775 1396 1125
rect 1430 775 1460 1125
rect 1494 775 1524 1125
rect 1558 775 1588 1125
rect 1622 775 1652 1125
rect 1686 775 1716 1125
rect 1750 775 1780 1125
rect 1814 775 1844 1125
rect 1878 805 1908 1095
rect 1944 805 1974 1095
rect 2008 775 2038 1125
rect 2072 775 2102 1125
rect 2136 775 2166 1125
rect 2200 775 2230 1125
rect 2264 775 2294 1125
rect 2328 775 2358 1125
rect 2392 775 2422 1125
rect 2456 775 2486 1125
rect 2520 805 2550 1095
rect 2586 805 2616 1095
rect 2650 775 2680 1125
rect 2714 775 2744 1125
rect 2778 775 2808 1125
rect 2842 775 2872 1125
rect 2906 775 2936 1125
rect 2970 775 3000 1125
rect 3034 775 3064 1125
rect 3098 775 3128 1125
rect 3162 805 3192 1095
rect 3228 805 3258 1095
rect 3292 775 3322 1125
rect 3356 775 3386 1125
rect 3420 775 3450 1125
rect 3484 775 3514 1125
rect 3548 775 3578 1125
rect 3612 775 3642 1125
rect 3676 775 3706 1125
rect 3740 775 3770 1125
rect 3804 805 3834 1095
rect 3870 805 3900 1095
rect 3934 775 3964 1125
rect 3998 775 4028 1125
rect 4062 775 4092 1125
rect 4126 775 4156 1125
rect 4190 775 4220 1125
rect 4254 775 4284 1125
rect 4318 775 4348 1125
rect 4382 775 4412 1125
rect 4446 805 4476 1095
rect 4512 805 4542 1095
rect 4576 775 4606 1125
rect 4640 775 4670 1125
rect 4704 775 4734 1125
rect 4768 775 4798 1125
rect 4832 775 4862 1125
rect 4896 775 4926 1125
rect 4960 775 4990 1125
rect 5024 775 5054 1125
rect 5088 805 5118 1095
rect 5154 805 5184 1095
rect 5218 775 5248 1125
rect 5282 775 5312 1125
rect 5346 775 5376 1125
rect 5410 775 5440 1125
rect 5474 775 5504 1125
rect 5538 775 5568 1125
rect 5602 775 5632 1125
rect 5666 775 5696 1125
rect 5730 805 5760 1095
rect 5796 805 5826 1095
rect 5860 775 5890 1125
rect 5924 775 5954 1125
rect 5988 775 6018 1125
rect 6052 775 6082 1125
rect 6116 775 6146 1125
rect 6180 775 6210 1125
rect 6244 775 6274 1125
rect 6308 775 6338 1125
rect 6372 805 6402 1095
rect 6438 805 6468 1095
rect 6502 775 6532 1125
rect 6566 775 6596 1125
rect 6630 775 6660 1125
rect 6694 775 6724 1125
rect 6758 775 6788 1125
rect 6822 775 6852 1125
rect 6886 775 6916 1125
rect 6950 775 6980 1125
rect 7014 805 7044 1095
rect 7080 805 7110 1095
rect 7144 775 7174 1125
rect 7208 775 7238 1125
rect 7272 775 7302 1125
rect 7336 775 7366 1125
rect 7400 775 7430 1125
rect 7464 775 7494 1125
rect 7528 775 7558 1125
rect 7592 775 7622 1125
rect 7656 805 7686 1095
rect 7722 805 7752 1095
rect 7786 775 7816 1125
rect 7850 775 7880 1125
rect 7914 775 7944 1125
rect 7978 775 8008 1125
rect 8042 775 8072 1125
rect 8106 775 8136 1125
rect 8170 775 8200 1125
rect 8234 775 8264 1125
rect 8298 805 8328 1095
rect 8364 805 8394 1095
rect 8428 775 8458 1125
rect 8492 775 8522 1125
rect 8556 775 8586 1125
rect 8620 775 8650 1125
rect 8684 775 8714 1125
rect 8748 775 8778 1125
rect 8812 775 8842 1125
rect 8876 775 8906 1125
rect 8940 805 8970 1095
rect 9006 805 9036 1095
rect 9070 775 9100 1125
rect 9134 775 9164 1125
rect 9198 775 9228 1125
rect 9262 775 9292 1125
rect 9326 775 9356 1125
rect 9390 775 9420 1125
rect 9454 775 9484 1125
rect 9518 775 9548 1125
rect 9582 805 9612 1095
rect 9648 805 9678 1095
rect 9712 775 9742 1125
rect 9776 775 9806 1125
rect 9840 775 9870 1125
rect 9904 775 9934 1125
rect 9968 775 9998 1125
rect 10032 775 10062 1125
rect 10096 775 10126 1125
rect 10160 775 10190 1125
rect 10224 805 10254 1095
rect 10290 805 10320 1095
rect 10354 775 10384 1125
rect 10418 775 10448 1125
rect 10482 775 10512 1125
rect 10546 775 10576 1125
rect 10610 775 10640 1125
rect 10674 775 10704 1125
rect 10738 775 10768 1125
rect 10802 775 10832 1125
rect 10866 805 10896 1095
rect 10932 805 10962 1095
rect 10996 775 11026 1125
rect 11060 775 11090 1125
rect 11124 775 11154 1125
rect 11188 775 11218 1125
rect 11252 775 11282 1125
rect 11316 775 11346 1125
rect 11380 775 11410 1125
rect 11444 775 11474 1125
rect 11508 805 11538 1095
rect 11574 805 11604 1095
rect 11638 775 11668 1125
rect 11702 775 11732 1125
rect 11766 775 11796 1125
rect 11830 775 11860 1125
rect 11894 775 11924 1125
rect 11958 775 11988 1125
rect 12022 775 12052 1125
rect 12086 775 12116 1125
rect 12150 805 12180 1095
rect 12216 805 12246 1095
rect 12280 775 12310 1125
rect 12344 775 12374 1125
rect 12408 775 12438 1125
rect 12472 775 12502 1125
rect 12536 775 12566 1125
rect 12600 775 12630 1125
rect 12664 775 12694 1125
rect 12728 775 12758 1125
rect 12792 805 12822 1095
rect 0 745 625 775
rect 659 745 2551 775
rect 2585 745 3835 775
rect 3869 745 5761 775
rect 5795 745 7045 775
rect 7079 745 8971 775
rect 9005 745 10255 775
rect 10289 745 12181 775
rect 12215 745 12840 775
rect 18 425 48 715
rect 82 395 112 745
rect 146 395 176 745
rect 210 395 240 745
rect 274 395 304 745
rect 338 395 368 745
rect 402 395 432 745
rect 466 395 496 745
rect 530 395 560 745
rect 594 425 624 715
rect 660 425 690 715
rect 724 395 754 745
rect 788 395 818 745
rect 852 395 882 745
rect 916 395 946 745
rect 980 395 1010 745
rect 1044 395 1074 745
rect 1108 395 1138 745
rect 1172 395 1202 745
rect 1236 425 1266 715
rect 1302 425 1332 715
rect 1366 395 1396 745
rect 1430 395 1460 745
rect 1494 395 1524 745
rect 1558 395 1588 745
rect 1622 395 1652 745
rect 1686 395 1716 745
rect 1750 395 1780 745
rect 1814 395 1844 745
rect 1878 425 1908 715
rect 1944 425 1974 715
rect 2008 395 2038 745
rect 2072 395 2102 745
rect 2136 395 2166 745
rect 2200 395 2230 745
rect 2264 395 2294 745
rect 2328 395 2358 745
rect 2392 395 2422 745
rect 2456 395 2486 745
rect 2520 425 2550 715
rect 2586 425 2616 715
rect 2650 395 2680 745
rect 2714 395 2744 745
rect 2778 395 2808 745
rect 2842 395 2872 745
rect 2906 395 2936 745
rect 2970 395 3000 745
rect 3034 395 3064 745
rect 3098 395 3128 745
rect 3162 425 3192 715
rect 3228 425 3258 715
rect 3292 395 3322 745
rect 3356 395 3386 745
rect 3420 395 3450 745
rect 3484 395 3514 745
rect 3548 395 3578 745
rect 3612 395 3642 745
rect 3676 395 3706 745
rect 3740 395 3770 745
rect 3804 425 3834 715
rect 3870 425 3900 715
rect 3934 395 3964 745
rect 3998 395 4028 745
rect 4062 395 4092 745
rect 4126 395 4156 745
rect 4190 395 4220 745
rect 4254 395 4284 745
rect 4318 395 4348 745
rect 4382 395 4412 745
rect 4446 425 4476 715
rect 4512 425 4542 715
rect 4576 395 4606 745
rect 4640 395 4670 745
rect 4704 395 4734 745
rect 4768 395 4798 745
rect 4832 395 4862 745
rect 4896 395 4926 745
rect 4960 395 4990 745
rect 5024 395 5054 745
rect 5088 425 5118 715
rect 5154 425 5184 715
rect 5218 395 5248 745
rect 5282 395 5312 745
rect 5346 395 5376 745
rect 5410 395 5440 745
rect 5474 395 5504 745
rect 5538 395 5568 745
rect 5602 395 5632 745
rect 5666 395 5696 745
rect 5730 425 5760 715
rect 5796 425 5826 715
rect 5860 395 5890 745
rect 5924 395 5954 745
rect 5988 395 6018 745
rect 6052 395 6082 745
rect 6116 395 6146 745
rect 6180 395 6210 745
rect 6244 395 6274 745
rect 6308 395 6338 745
rect 6372 425 6402 715
rect 6438 425 6468 715
rect 6502 395 6532 745
rect 6566 395 6596 745
rect 6630 395 6660 745
rect 6694 395 6724 745
rect 6758 395 6788 745
rect 6822 395 6852 745
rect 6886 395 6916 745
rect 6950 395 6980 745
rect 7014 425 7044 715
rect 7080 425 7110 715
rect 7144 395 7174 745
rect 7208 395 7238 745
rect 7272 395 7302 745
rect 7336 395 7366 745
rect 7400 395 7430 745
rect 7464 395 7494 745
rect 7528 395 7558 745
rect 7592 395 7622 745
rect 7656 425 7686 715
rect 7722 425 7752 715
rect 7786 395 7816 745
rect 7850 395 7880 745
rect 7914 395 7944 745
rect 7978 395 8008 745
rect 8042 395 8072 745
rect 8106 395 8136 745
rect 8170 395 8200 745
rect 8234 395 8264 745
rect 8298 425 8328 715
rect 8364 425 8394 715
rect 8428 395 8458 745
rect 8492 395 8522 745
rect 8556 395 8586 745
rect 8620 395 8650 745
rect 8684 395 8714 745
rect 8748 395 8778 745
rect 8812 395 8842 745
rect 8876 395 8906 745
rect 8940 425 8970 715
rect 9006 425 9036 715
rect 9070 395 9100 745
rect 9134 395 9164 745
rect 9198 395 9228 745
rect 9262 395 9292 745
rect 9326 395 9356 745
rect 9390 395 9420 745
rect 9454 395 9484 745
rect 9518 395 9548 745
rect 9582 425 9612 715
rect 9648 425 9678 715
rect 9712 395 9742 745
rect 9776 395 9806 745
rect 9840 395 9870 745
rect 9904 395 9934 745
rect 9968 395 9998 745
rect 10032 395 10062 745
rect 10096 395 10126 745
rect 10160 395 10190 745
rect 10224 425 10254 715
rect 10290 425 10320 715
rect 10354 395 10384 745
rect 10418 395 10448 745
rect 10482 395 10512 745
rect 10546 395 10576 745
rect 10610 395 10640 745
rect 10674 395 10704 745
rect 10738 395 10768 745
rect 10802 395 10832 745
rect 10866 425 10896 715
rect 10932 425 10962 715
rect 10996 395 11026 745
rect 11060 395 11090 745
rect 11124 395 11154 745
rect 11188 395 11218 745
rect 11252 395 11282 745
rect 11316 395 11346 745
rect 11380 395 11410 745
rect 11444 395 11474 745
rect 11508 425 11538 715
rect 11574 425 11604 715
rect 11638 395 11668 745
rect 11702 395 11732 745
rect 11766 395 11796 745
rect 11830 395 11860 745
rect 11894 395 11924 745
rect 11958 395 11988 745
rect 12022 395 12052 745
rect 12086 395 12116 745
rect 12150 425 12180 715
rect 12216 425 12246 715
rect 12280 395 12310 745
rect 12344 395 12374 745
rect 12408 395 12438 745
rect 12472 395 12502 745
rect 12536 395 12566 745
rect 12600 395 12630 745
rect 12664 395 12694 745
rect 12728 395 12758 745
rect 12792 425 12822 715
rect 0 365 625 395
rect 659 365 2551 395
rect 2585 365 3835 395
rect 3869 365 5761 395
rect 5795 365 7045 395
rect 7079 365 8971 395
rect 9005 365 10255 395
rect 10289 365 12181 395
rect 12215 365 12840 395
rect 18 45 48 335
rect 82 15 112 365
rect 146 15 176 365
rect 210 15 240 365
rect 274 15 304 365
rect 338 15 368 365
rect 402 15 432 365
rect 466 15 496 365
rect 530 15 560 365
rect 594 45 624 335
rect 660 45 690 335
rect 724 15 754 335
rect 788 15 818 335
rect 852 15 882 335
rect 916 15 946 335
rect 980 15 1010 335
rect 1044 15 1074 335
rect 1108 15 1138 335
rect 1172 15 1202 335
rect 1236 45 1266 335
rect 1302 45 1332 335
rect 1366 15 1396 335
rect 1430 15 1460 335
rect 1494 15 1524 335
rect 1558 15 1588 335
rect 1622 15 1652 335
rect 1686 15 1716 335
rect 1750 15 1780 335
rect 1814 15 1844 335
rect 1878 45 1908 335
rect 1944 45 1974 335
rect 2008 15 2038 335
rect 2072 15 2102 335
rect 2136 15 2166 335
rect 2200 15 2230 335
rect 2264 15 2294 335
rect 2328 15 2358 335
rect 2392 15 2422 335
rect 2456 15 2486 335
rect 2520 45 2550 335
rect 2586 45 2616 335
rect 2650 15 2680 365
rect 2714 15 2744 365
rect 2778 15 2808 365
rect 2842 15 2872 365
rect 2906 15 2936 365
rect 2970 15 3000 365
rect 3034 15 3064 365
rect 3098 15 3128 365
rect 3162 45 3192 335
rect 3228 45 3258 335
rect 3292 15 3322 365
rect 3356 15 3386 365
rect 3420 15 3450 365
rect 3484 15 3514 365
rect 3548 15 3578 365
rect 3612 15 3642 365
rect 3676 15 3706 365
rect 3740 15 3770 365
rect 3804 45 3834 335
rect 3870 45 3900 335
rect 3934 15 3964 335
rect 3998 15 4028 335
rect 4062 15 4092 335
rect 4126 15 4156 335
rect 4190 15 4220 335
rect 4254 15 4284 335
rect 4318 15 4348 335
rect 4382 15 4412 335
rect 4446 45 4476 335
rect 4512 45 4542 335
rect 4576 15 4606 335
rect 4640 15 4670 335
rect 4704 15 4734 335
rect 4768 15 4798 335
rect 4832 15 4862 365
rect 4896 15 4926 365
rect 4960 15 4990 365
rect 5024 15 5054 365
rect 5088 45 5118 335
rect 5154 45 5184 335
rect 5218 15 5248 335
rect 5282 15 5312 335
rect 5346 15 5376 335
rect 5410 15 5440 335
rect 5474 15 5504 335
rect 5538 15 5568 335
rect 5602 15 5632 335
rect 5666 15 5696 335
rect 5730 45 5760 335
rect 5796 45 5826 335
rect 5860 15 5890 365
rect 5924 15 5954 365
rect 5988 15 6018 365
rect 6052 15 6082 365
rect 6116 15 6146 365
rect 6180 15 6210 365
rect 6244 15 6274 365
rect 6308 15 6338 365
rect 6372 45 6402 335
rect 6438 45 6468 335
rect 6502 15 6532 365
rect 6566 15 6596 365
rect 6630 15 6660 365
rect 6694 15 6724 365
rect 6758 15 6788 365
rect 6822 15 6852 365
rect 6886 15 6916 365
rect 6950 15 6980 365
rect 7014 45 7044 335
rect 7080 45 7110 335
rect 7144 15 7174 335
rect 7208 15 7238 335
rect 7272 15 7302 335
rect 7336 15 7366 335
rect 7400 15 7430 335
rect 7464 15 7494 335
rect 7528 15 7558 335
rect 7592 15 7622 335
rect 7656 45 7686 335
rect 7722 45 7752 335
rect 7786 15 7816 335
rect 7850 15 7880 335
rect 7914 15 7944 335
rect 7978 15 8008 335
rect 8042 15 8072 335
rect 8106 15 8136 335
rect 8170 15 8200 365
rect 8234 15 8264 365
rect 8298 45 8328 335
rect 8364 45 8394 335
rect 8428 15 8458 335
rect 8492 15 8522 335
rect 8556 15 8586 335
rect 8620 15 8650 335
rect 8684 15 8714 335
rect 8748 15 8778 335
rect 8812 15 8842 335
rect 8876 15 8906 335
rect 8940 45 8970 335
rect 9006 45 9036 335
rect 9070 15 9100 365
rect 9134 15 9164 365
rect 9198 15 9228 365
rect 9262 15 9292 365
rect 9326 15 9356 365
rect 9390 15 9420 365
rect 9454 15 9484 365
rect 9518 15 9548 365
rect 9582 45 9612 335
rect 9648 45 9678 335
rect 9712 15 9742 365
rect 9776 15 9806 365
rect 9840 15 9870 365
rect 9904 15 9934 365
rect 9968 15 9998 365
rect 10032 15 10062 365
rect 10096 15 10126 365
rect 10160 15 10190 365
rect 10224 45 10254 335
rect 10290 45 10320 335
rect 10354 15 10384 335
rect 10418 15 10448 335
rect 10482 15 10512 335
rect 10546 15 10576 335
rect 10610 15 10640 335
rect 10674 15 10704 335
rect 10738 15 10768 335
rect 10802 15 10832 335
rect 10866 45 10896 335
rect 10932 45 10962 335
rect 10996 15 11026 335
rect 11060 15 11090 335
rect 11124 15 11154 335
rect 11188 15 11218 335
rect 11252 15 11282 335
rect 11316 15 11346 335
rect 11380 15 11410 335
rect 11444 15 11474 365
rect 11508 45 11538 335
rect 11574 45 11604 335
rect 11638 15 11668 335
rect 11702 15 11732 335
rect 11766 15 11796 335
rect 11830 15 11860 335
rect 11894 15 11924 335
rect 11958 15 11988 335
rect 12022 15 12052 335
rect 12086 15 12116 335
rect 12150 45 12180 335
rect 12216 45 12246 335
rect 12280 15 12310 365
rect 12344 15 12374 365
rect 12408 15 12438 365
rect 12472 15 12502 365
rect 12536 15 12566 365
rect 12600 15 12630 365
rect 12664 15 12694 365
rect 12728 15 12758 365
rect 12792 45 12822 335
rect 0 -15 4478 15
rect 4510 -15 4798 15
rect 4828 -15 5120 15
rect 5152 -15 7688 15
rect 7720 -15 8136 15
rect 8166 -15 8299 15
rect 8362 -15 10898 15
rect 10930 -15 11410 15
rect 11440 -15 11478 15
rect 11572 -15 12840 15
<< labels >>
rlabel metal4 0 745 0 775 7 dummy_top
rlabel metal2 14 790 14 820 7 dummy_bot
rlabel metal4 659 365 659 395 7 top_8
rlabel metal2 656 410 656 440 7 bot_8
rlabel metal4 3869 365 3869 395 7 top_4
rlabel metal2 3866 410 3866 440 7 bot_4
rlabel metal4 7079 365 7079 395 7 top_2
rlabel metal2 7076 410 7076 440 7 bot_2
rlabel metal4 10289 365 10289 395 7 top_1
rlabel metal2 10286 410 10286 440 7 bot_1
<< end >>
