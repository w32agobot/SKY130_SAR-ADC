* SPICE3 file created from adc_array_fingercap_8(1)x700aF_23um2.ext - technology: sky130A

C0 cbot floatingmetal 2.60fF
C1 cbot ctop 0.70fF
C2 floatingmetal VSUBS 0.33fF
C3 ctop VSUBS 0.22fF
C4 cbot VSUBS 1.90fF
