magic
tech sky130A
magscale 1 2
timestamp 1662655812
<< nwell >>
rect -38 247 1878 582
<< pwell >>
rect 1 -17 1839 214
<< nmos >>
rect 160 95 959 179
rect 1154 80 1184 164
rect 1250 80 1280 164
rect 1454 80 1484 164
rect 1550 80 1580 164
<< pmos >>
rect 1132 296 1162 456
rect 1228 296 1258 456
rect 1548 296 1578 456
rect 1644 296 1674 456
<< pmoslvt >>
rect 160 283 959 443
<< ndiff >>
rect 102 167 160 179
rect 102 107 114 167
rect 148 107 160 167
rect 102 95 160 107
rect 959 167 1017 179
rect 959 107 971 167
rect 1005 107 1017 167
rect 959 95 1017 107
rect 1094 152 1154 164
rect 1094 92 1104 152
rect 1138 92 1154 152
rect 1094 80 1154 92
rect 1184 152 1250 164
rect 1184 92 1200 152
rect 1234 92 1250 152
rect 1184 80 1250 92
rect 1280 152 1338 164
rect 1280 92 1296 152
rect 1330 92 1338 152
rect 1280 80 1338 92
rect 1392 152 1454 164
rect 1392 92 1404 152
rect 1438 92 1454 152
rect 1392 80 1454 92
rect 1484 152 1550 164
rect 1484 92 1500 152
rect 1534 92 1550 152
rect 1484 80 1550 92
rect 1580 152 1642 164
rect 1580 92 1596 152
rect 1630 92 1642 152
rect 1580 80 1642 92
<< pdiff >>
rect 1072 444 1132 456
rect 102 431 160 443
rect 102 295 114 431
rect 148 295 160 431
rect 102 283 160 295
rect 959 431 1017 443
rect 959 295 971 431
rect 1005 295 1017 431
rect 1072 308 1082 444
rect 1116 308 1132 444
rect 1072 296 1132 308
rect 1162 444 1228 456
rect 1162 308 1178 444
rect 1212 308 1228 444
rect 1162 296 1228 308
rect 1258 444 1318 456
rect 1258 308 1274 444
rect 1308 308 1318 444
rect 1258 296 1318 308
rect 1486 444 1548 456
rect 1486 308 1498 444
rect 1532 308 1548 444
rect 1486 296 1548 308
rect 1578 444 1644 456
rect 1578 308 1594 444
rect 1628 308 1644 444
rect 1578 296 1644 308
rect 1674 444 1734 456
rect 1674 308 1690 444
rect 1724 308 1734 444
rect 1674 296 1734 308
rect 959 283 1017 295
<< ndiffc >>
rect 114 107 148 167
rect 971 107 1005 167
rect 1104 92 1138 152
rect 1200 92 1234 152
rect 1296 92 1330 152
rect 1404 92 1438 152
rect 1500 92 1534 152
rect 1596 92 1630 152
<< pdiffc >>
rect 114 295 148 431
rect 971 295 1005 431
rect 1082 308 1116 444
rect 1178 308 1212 444
rect 1274 308 1308 444
rect 1498 308 1532 444
rect 1594 308 1628 444
rect 1690 308 1724 444
<< poly >>
rect 160 443 959 479
rect 1132 456 1162 490
rect 1228 456 1258 490
rect 1548 456 1578 490
rect 1644 456 1674 490
rect 160 264 959 283
rect 25 248 959 264
rect 1132 280 1162 296
rect 1228 280 1258 296
rect 1132 258 1280 280
rect 25 214 35 248
rect 70 214 959 248
rect 25 198 959 214
rect 1074 250 1280 258
rect 1074 248 1184 250
rect 1074 214 1112 248
rect 1146 214 1184 248
rect 1074 202 1184 214
rect 160 179 959 198
rect 1154 164 1184 202
rect 1250 164 1280 250
rect 1340 252 1406 262
rect 1340 218 1356 252
rect 1390 220 1406 252
rect 1548 220 1578 296
rect 1644 220 1674 296
rect 1390 218 1674 220
rect 1340 190 1674 218
rect 1454 164 1484 190
rect 1550 164 1580 190
rect 160 69 959 95
rect 1154 54 1184 80
rect 1250 54 1280 80
rect 1454 54 1484 80
rect 1550 54 1580 80
<< polycont >>
rect 35 214 70 248
rect 1112 214 1146 248
rect 1356 218 1390 252
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1840 561
rect 114 431 148 447
rect 114 279 148 295
rect 971 431 1005 447
rect 25 248 73 264
rect 25 214 35 248
rect 70 214 73 248
rect 25 198 73 214
rect 971 258 1005 295
rect 1082 444 1116 527
rect 1082 292 1116 308
rect 1178 444 1212 460
rect 1178 292 1212 308
rect 1274 444 1308 460
rect 1274 292 1308 308
rect 971 248 1162 258
rect 971 214 1112 248
rect 1146 214 1162 248
rect 971 202 1162 214
rect 1356 252 1390 268
rect 1424 258 1458 527
rect 1492 444 1532 460
rect 1492 308 1498 444
rect 1492 292 1532 308
rect 1594 444 1628 460
rect 1424 224 1534 258
rect 1356 202 1390 218
rect 114 167 148 183
rect 114 91 148 107
rect 971 167 1005 202
rect 971 73 1005 107
rect 1104 152 1138 168
rect 405 17 439 48
rect 913 17 947 48
rect 1104 17 1138 92
rect 1200 152 1234 168
rect 1200 76 1234 92
rect 1296 76 1330 92
rect 1404 152 1438 168
rect 1404 76 1438 92
rect 1500 152 1534 224
rect 1594 236 1628 308
rect 1690 444 1730 460
rect 1724 308 1730 444
rect 1690 292 1730 308
rect 1732 254 1778 258
rect 1594 202 1698 236
rect 1500 76 1534 92
rect 1596 152 1630 168
rect 1596 76 1630 92
rect 1664 17 1698 202
rect 1732 220 1738 254
rect 1772 220 1778 254
rect 1732 196 1778 220
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1840 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 114 295 148 431
rect 1178 308 1212 444
rect 1274 308 1308 364
rect 1356 218 1390 252
rect 1498 328 1532 444
rect 114 107 148 167
rect 1200 92 1234 152
rect 1296 152 1330 178
rect 1296 144 1330 152
rect 1404 92 1438 132
rect 1690 328 1724 444
rect 1596 92 1630 132
rect 1738 220 1772 254
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
<< metal1 >>
rect 0 561 1840 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1840 561
rect 0 496 1840 527
rect 108 431 154 496
rect 108 295 114 431
rect 148 295 154 431
rect 1172 444 1730 456
rect 1172 308 1178 444
rect 1212 422 1498 444
rect 1212 308 1218 422
rect 1172 296 1218 308
rect 1268 364 1314 394
rect 1268 308 1274 364
rect 1308 308 1314 364
rect 1492 328 1498 422
rect 1532 422 1690 444
rect 1532 328 1538 422
rect 1492 316 1538 328
rect 1684 328 1690 422
rect 1724 328 1730 444
rect 1684 316 1730 328
rect 108 283 154 295
rect 1268 248 1314 308
rect 1350 252 1396 264
rect 1350 248 1356 252
rect 1268 220 1356 248
rect 1290 218 1356 220
rect 1390 248 1396 252
rect 1726 254 1784 260
rect 1726 248 1738 254
rect 1390 220 1738 248
rect 1772 220 1784 254
rect 1390 218 1396 220
rect 1290 206 1396 218
rect 1726 214 1784 220
rect 108 167 154 182
rect 108 107 114 167
rect 148 107 154 167
rect 1290 178 1336 206
rect 108 48 154 107
rect 1194 152 1240 164
rect 1194 92 1200 152
rect 1234 104 1240 152
rect 1290 144 1296 178
rect 1330 144 1336 178
rect 1290 132 1336 144
rect 1398 132 1444 144
rect 1398 104 1404 132
rect 1234 92 1404 104
rect 1438 104 1444 132
rect 1590 132 1636 144
rect 1590 104 1596 132
rect 1438 92 1596 104
rect 1630 92 1636 132
rect 1194 76 1636 92
rect 0 17 1840 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1840 17
rect 0 -48 1840 -17
<< labels >>
flabel metal1 s 0 496 1840 592 0 FreeSans 160 0 0 0 VPWR
port 3 nsew power bidirectional abutment
flabel metal1 s 213 527 247 561 0 FreeSans 160 0 0 0 VPWR
port 3 nsew power bidirectional abutment
flabel metal1 s 213 -17 247 17 0 FreeSans 160 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 0 -48 1840 48 0 FreeSans 160 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel nwell s 213 527 247 561 0 FreeSans 160 0 0 0 VPB
port 5 nsew power bidirectional
flabel pwell s 213 -17 247 17 0 FreeSans 160 0 0 0 VNB
port 6 nsew ground bidirectional
flabel metal1 s 1738 220 1772 254 0 FreeSans 160 0 0 0 out
port 2 nsew signal output
flabel locali s 38 221 72 255 7 FreeSans 160 0 0 0 in
port 1 nsew signal input
rlabel locali 971 169 1005 169 1 cap_top
<< properties >>
string FIXED_BBOX 0 0 1840 544
string LEFclass CORE
string LEForigin 0 0
string LEFsite unithd
string LEFsource USER
<< end >>
