* SPICE3 file created from adc_array_wafflecap_8(1)x560aF_25um2.ext - technology: sky130A

.subckt adc_array_wafflecap_8(1)x560aF_25um2 cbot ctop
C0 ctop cbot 0.57fF
C1 cbot nc 3.78fF
C2 cbot VSUBS 2.01fF
C3 nc VSUBS 0.46fF
.ends
