* SPICE3 file created from adc_noise_decoup_cell1.ext - technology: sky130A

.subckt adc_noise_decoup_cell1 nmoscap_top nmoscap_bot mimcap_top mimcap_bot pwell
X0 mimcap_top mimcap_bot sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X1 nmoscap_bot nmoscap_top nmoscap_bot pwell sky130_fd_pr__nfet_01v8 ad=2.296e+13p pd=6.84e+07u as=0p ps=0u w=1.64e+07u l=1.6e+07u
C0 nmoscap_top mimcap_bot 15.25fF
C1 nmoscap_top nmoscap_bot 510.69fF
C2 mimcap_bot nmoscap_bot 16.58fF
C3 nmoscap_top mimcap_top 2.89fF
C4 mimcap_top mimcap_bot 33.25fF
C5 nmoscap_top pwell 13.14fF
C6 mimcap_top pwell 2.10fF
C7 mimcap_bot pwell 2.60fF
C8 nmoscap_bot pwell 8.64fF
.ends
