magic
tech sky130A
magscale 1 2
timestamp 1661178173
<< metal3 >>
rect -750 4522 749 4550
rect -750 2378 665 4522
rect 729 2378 749 4522
rect -750 2350 749 2378
rect -750 2222 749 2250
rect -750 78 665 2222
rect 729 78 749 2222
rect -750 50 749 78
rect -750 -78 749 -50
rect -750 -2222 665 -78
rect 729 -2222 749 -78
rect -750 -2250 749 -2222
rect -750 -2378 749 -2350
rect -750 -4522 665 -2378
rect 729 -4522 749 -2378
rect -750 -4550 749 -4522
<< via3 >>
rect 665 2378 729 4522
rect 665 78 729 2222
rect 665 -2222 729 -78
rect 665 -4522 729 -2378
<< mimcap >>
rect -650 4410 550 4450
rect -650 2490 -610 4410
rect 510 2490 550 4410
rect -650 2450 550 2490
rect -650 2110 550 2150
rect -650 190 -610 2110
rect 510 190 550 2110
rect -650 150 550 190
rect -650 -190 550 -150
rect -650 -2110 -610 -190
rect 510 -2110 550 -190
rect -650 -2150 550 -2110
rect -650 -2490 550 -2450
rect -650 -4410 -610 -2490
rect 510 -4410 550 -2490
rect -650 -4450 550 -4410
<< mimcapcontact >>
rect -610 2490 510 4410
rect -610 190 510 2110
rect -610 -2110 510 -190
rect -610 -4410 510 -2490
<< metal4 >>
rect -102 4411 2 4600
rect 618 4538 722 4600
rect 618 4522 745 4538
rect -611 4410 511 4411
rect -611 2490 -610 4410
rect 510 2490 511 4410
rect -611 2489 511 2490
rect -102 2111 2 2489
rect 618 2378 665 4522
rect 729 2378 745 4522
rect 618 2362 745 2378
rect 618 2238 722 2362
rect 618 2222 745 2238
rect -611 2110 511 2111
rect -611 190 -610 2110
rect 510 190 511 2110
rect -611 189 511 190
rect -102 -189 2 189
rect 618 78 665 2222
rect 729 78 745 2222
rect 618 62 745 78
rect 618 -62 722 62
rect 618 -78 745 -62
rect -611 -190 511 -189
rect -611 -2110 -610 -190
rect 510 -2110 511 -190
rect -611 -2111 511 -2110
rect -102 -2489 2 -2111
rect 618 -2222 665 -78
rect 729 -2222 745 -78
rect 618 -2238 745 -2222
rect 618 -2362 722 -2238
rect 618 -2378 745 -2362
rect -611 -2490 511 -2489
rect -611 -4410 -610 -2490
rect 510 -4410 511 -2490
rect -611 -4411 511 -4410
rect -102 -4600 2 -4411
rect 618 -4522 665 -2378
rect 729 -4522 745 -2378
rect 618 -4538 745 -4522
rect 618 -4600 722 -4538
<< properties >>
string FIXED_BBOX -750 2350 650 4550
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 6 l 10 val 126.08 carea 2.00 cperi 0.19 nx 1 ny 4 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
