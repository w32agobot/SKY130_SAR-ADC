* NGSPICE file created from adc_vcm_generator.ext - technology: sky130A

.subckt sky130_fd_sc_hd__inv_1 A VGND VPWR Y VNB VPB
X0 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
.ends

.subckt pfet_01v8_w500_l500_nf2 a_n29_0# a_129_0# a_n129_n26# w_n224_n36# a_n187_0#
+ a_29_n26#
X0 a_129_0# a_29_n26# a_n29_0# w_n224_n36# sky130_fd_pr__pfet_01v8 ad=1.45e+11p pd=1.58e+06u as=1.45e+11p ps=1.58e+06u w=500000u l=500000u
X1 a_n29_0# a_n129_n26# a_n187_0# w_n224_n36# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.45e+11p ps=1.58e+06u w=500000u l=500000u
.ends

.subckt sky130_fd_sc_hd__buf_4 A VGND VPWR X VNB VPB
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=8e+11p pd=7.6e+06u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=5.2e+11p ps=5.5e+06u w=650000u l=150000u
X5 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X9 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__dlymetal6s6s_1 A VGND VPWR X VNB VPB
X0 X a_629_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=5.82e+11p ps=5.85e+06u w=650000u l=150000u
X1 a_523_47# a_346_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X2 VGND a_240_47# a_346_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X3 a_240_47# a_63_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X4 VPWR a_240_47# a_346_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=8.445e+11p pd=7.95e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X5 VGND A a_63_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X6 VPWR A a_63_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X7 VPWR a_523_47# a_629_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X8 VGND a_523_47# a_629_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X9 a_523_47# a_346_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X10 a_240_47# a_63_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X11 X a_629_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt adc_noise_decoup_cell1 nmoscap_top nmoscap_bot mimcap_top mimcap_bot pwell
X0 mimcap_top mimcap_bot sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X1 nmoscap_bot nmoscap_top nmoscap_bot pwell sky130_fd_pr__nfet_01v8 ad=2.296e+13p pd=6.84e+07u as=0p ps=0u w=1.64e+07u l=1.6e+07u
.ends

.subckt nfet_01v8_w500_l500_nf2 a_n129_n76# a_n29_n50# a_n187_n50# a_29_n76# a_129_n50#
+ VSUBS
X0 a_129_n50# a_29_n76# a_n29_n50# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45e+11p pd=1.58e+06u as=1.45e+11p ps=1.58e+06u w=500000u l=500000u
X1 a_n29_n50# a_n129_n76# a_n187_n50# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.45e+11p ps=1.58e+06u w=500000u l=500000u
.ends

.subckt sky130_fd_sc_hd__nand2_1 A B VGND VPWR Y VNB VPB
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=5.2e+11p pd=5.04e+06u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1 Y A a_113_47# VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X2 a_113_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X3 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt adc_vcm_generator VPWR VGND clk vcm
Xsky130_fd_sc_hd__inv_1_4 clk VGND VPWR sky130_fd_sc_hd__inv_1_4/Y VGND VPWR sky130_fd_sc_hd__inv_1
Xpfet_01v8_w500_l500_nf2_0 mimtop2 vcm phi1_n VPWR vcm phi1_n pfet_01v8_w500_l500_nf2
Xpfet_01v8_w500_l500_nf2_1 mimtop1 vcm phi1_n VPWR vcm phi1_n pfet_01v8_w500_l500_nf2
Xsky130_fd_sc_hd__buf_4_0 sky130_fd_sc_hd__inv_1_2/A VGND VPWR phi1 VGND VPWR sky130_fd_sc_hd__buf_4
Xpfet_01v8_w500_l500_nf2_2 mimtop2 mimbot1 phi2_n VPWR mimbot1 phi2_n pfet_01v8_w500_l500_nf2
Xsky130_fd_sc_hd__buf_4_1 sky130_fd_sc_hd__inv_1_2/Y VGND VPWR phi1_n VGND VPWR sky130_fd_sc_hd__buf_4
Xpfet_01v8_w500_l500_nf2_3 VPWR mimtop1 phi2_n VPWR mimtop1 phi2_n pfet_01v8_w500_l500_nf2
Xpfet_01v8_w500_l500_nf2_4 mimbot1 VGND phi1_n VPWR VGND phi1_n pfet_01v8_w500_l500_nf2
Xsky130_fd_sc_hd__buf_4_2 sky130_fd_sc_hd__inv_1_3/A VGND VPWR phi2 VGND VPWR sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_3 sky130_fd_sc_hd__inv_1_3/Y VGND VPWR phi2_n VGND VPWR sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__dlymetal6s6s_1_0 sky130_fd_sc_hd__nand2_1_0/Y VGND VPWR sky130_fd_sc_hd__dlymetal6s6s_1_2/A
+ VGND VPWR sky130_fd_sc_hd__dlymetal6s6s_1
Xsky130_fd_sc_hd__dlymetal6s6s_1_1 sky130_fd_sc_hd__nand2_1_1/Y VGND VPWR sky130_fd_sc_hd__dlymetal6s6s_1_4/A
+ VGND VPWR sky130_fd_sc_hd__dlymetal6s6s_1
Xsky130_fd_sc_hd__dlymetal6s6s_1_2 sky130_fd_sc_hd__dlymetal6s6s_1_2/A VGND VPWR sky130_fd_sc_hd__dlymetal6s6s_1_3/A
+ VGND VPWR sky130_fd_sc_hd__dlymetal6s6s_1
Xsky130_fd_sc_hd__dlymetal6s6s_1_3 sky130_fd_sc_hd__dlymetal6s6s_1_3/A VGND VPWR sky130_fd_sc_hd__inv_1_0/A
+ VGND VPWR sky130_fd_sc_hd__dlymetal6s6s_1
Xsky130_fd_sc_hd__dlymetal6s6s_1_4 sky130_fd_sc_hd__dlymetal6s6s_1_4/A VGND VPWR sky130_fd_sc_hd__dlymetal6s6s_1_5/A
+ VGND VPWR sky130_fd_sc_hd__dlymetal6s6s_1
Xsky130_fd_sc_hd__dlymetal6s6s_1_5 sky130_fd_sc_hd__dlymetal6s6s_1_5/A VGND VPWR sky130_fd_sc_hd__inv_1_1/A
+ VGND VPWR sky130_fd_sc_hd__dlymetal6s6s_1
Xadc_noise_decoup_cell1_0[0] VPWR VGND VPWR VGND VGND adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_0[1] VPWR VGND VPWR VGND VGND adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_0[2] VPWR VGND VPWR VGND VGND adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[0|0] vcm VGND mimtop2 VGND VGND adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[1|0] vcm VGND mimtop2 VGND VGND adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[2|0] vcm VGND mimtop2 VGND VGND adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[3|0] vcm VGND mimtop2 VGND VGND adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[4|0] vcm VGND mimtop2 VGND VGND adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[5|0] vcm VGND mimtop2 VGND VGND adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[6|0] vcm VGND mimtop2 VGND VGND adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[7|0] vcm VGND mimtop2 VGND VGND adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[0|1] vcm VGND mimtop2 VGND VGND adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[1|1] vcm VGND mimtop2 VGND VGND adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[2|1] vcm VGND mimtop2 VGND VGND adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[3|1] vcm VGND mimtop2 VGND VGND adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[4|1] vcm VGND mimtop2 VGND VGND adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[5|1] vcm VGND mimtop2 VGND VGND adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[6|1] vcm VGND mimtop2 VGND VGND adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[7|1] vcm VGND mimtop2 VGND VGND adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[0|2] vcm VGND mimtop2 VGND VGND adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[1|2] vcm VGND mimtop2 VGND VGND adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[2|2] vcm VGND mimtop2 VGND VGND adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[3|2] vcm VGND mimtop2 VGND VGND adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[4|2] vcm VGND mimtop2 VGND VGND adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[5|2] vcm VGND mimtop2 VGND VGND adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[6|2] vcm VGND mimtop2 VGND VGND adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[7|2] vcm VGND mimtop2 VGND VGND adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[0|3] vcm VGND mimtop2 VGND VGND adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[1|3] vcm VGND mimtop2 VGND VGND adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[2|3] vcm VGND mimtop2 VGND VGND adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[3|3] vcm VGND mimtop2 VGND VGND adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[4|3] vcm VGND mimtop2 VGND VGND adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[5|3] vcm VGND mimtop2 VGND VGND adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[6|3] vcm VGND mimtop2 VGND VGND adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[7|3] vcm VGND mimtop2 VGND VGND adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[0|4] vcm VGND mimtop2 VGND VGND adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[1|4] vcm VGND mimtop2 VGND VGND adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[2|4] vcm VGND mimtop2 VGND VGND adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[3|4] vcm VGND mimtop2 VGND VGND adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[4|4] vcm VGND mimtop2 VGND VGND adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[5|4] vcm VGND mimtop2 VGND VGND adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[6|4] vcm VGND mimtop2 VGND VGND adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[7|4] vcm VGND mimtop2 VGND VGND adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[0|0] vcm VGND mimtop1 mimbot1 VGND adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[1|0] vcm VGND mimtop1 mimbot1 VGND adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[2|0] vcm VGND mimtop1 mimbot1 VGND adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[3|0] vcm VGND mimtop1 mimbot1 VGND adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[4|0] vcm VGND mimtop1 mimbot1 VGND adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[5|0] vcm VGND mimtop1 mimbot1 VGND adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[6|0] vcm VGND mimtop1 mimbot1 VGND adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[7|0] vcm VGND mimtop1 mimbot1 VGND adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[0|1] vcm VGND mimtop1 mimbot1 VGND adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[1|1] vcm VGND mimtop1 mimbot1 VGND adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[2|1] vcm VGND mimtop1 mimbot1 VGND adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[3|1] vcm VGND mimtop1 mimbot1 VGND adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[4|1] vcm VGND mimtop1 mimbot1 VGND adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[5|1] vcm VGND mimtop1 mimbot1 VGND adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[6|1] vcm VGND mimtop1 mimbot1 VGND adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[7|1] vcm VGND mimtop1 mimbot1 VGND adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[0|2] vcm VGND mimtop1 mimbot1 VGND adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[1|2] vcm VGND mimtop1 mimbot1 VGND adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[2|2] vcm VGND mimtop1 mimbot1 VGND adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[3|2] vcm VGND mimtop1 mimbot1 VGND adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[4|2] vcm VGND mimtop1 mimbot1 VGND adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[5|2] vcm VGND mimtop1 mimbot1 VGND adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[6|2] vcm VGND mimtop1 mimbot1 VGND adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[7|2] vcm VGND mimtop1 mimbot1 VGND adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[0|3] vcm VGND mimtop1 mimbot1 VGND adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[1|3] vcm VGND mimtop1 mimbot1 VGND adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[2|3] vcm VGND mimtop1 mimbot1 VGND adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[3|3] vcm VGND mimtop1 mimbot1 VGND adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[4|3] vcm VGND mimtop1 mimbot1 VGND adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[5|3] vcm VGND mimtop1 mimbot1 VGND adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[6|3] vcm VGND mimtop1 mimbot1 VGND adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[7|3] vcm VGND mimtop1 mimbot1 VGND adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[0|4] vcm VGND mimtop1 mimbot1 VGND adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[1|4] vcm VGND mimtop1 mimbot1 VGND adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[2|4] vcm VGND mimtop1 mimbot1 VGND adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[3|4] vcm VGND mimtop1 mimbot1 VGND adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[4|4] vcm VGND mimtop1 mimbot1 VGND adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[5|4] vcm VGND mimtop1 mimbot1 VGND adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[6|4] vcm VGND mimtop1 mimbot1 VGND adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[7|4] vcm VGND mimtop1 mimbot1 VGND adc_noise_decoup_cell1
Xnfet_01v8_w500_l500_nf2_0 phi1 mimtop2 vcm phi1 vcm VGND nfet_01v8_w500_l500_nf2
Xnfet_01v8_w500_l500_nf2_1 phi1 mimtop1 vcm phi1 vcm VGND nfet_01v8_w500_l500_nf2
Xsky130_fd_sc_hd__nand2_1_0 clk sky130_fd_sc_hd__inv_1_3/Y VGND VPWR sky130_fd_sc_hd__nand2_1_0/Y
+ VGND VPWR sky130_fd_sc_hd__nand2_1
Xnfet_01v8_w500_l500_nf2_2 phi2 mimtop2 mimbot1 phi2 mimbot1 VGND nfet_01v8_w500_l500_nf2
Xnfet_01v8_w500_l500_nf2_3 phi2 VPWR mimtop1 phi2 mimtop1 VGND nfet_01v8_w500_l500_nf2
Xsky130_fd_sc_hd__nand2_1_1 sky130_fd_sc_hd__inv_1_2/Y sky130_fd_sc_hd__inv_1_4/Y
+ VGND VPWR sky130_fd_sc_hd__nand2_1_1/Y VGND VPWR sky130_fd_sc_hd__nand2_1
Xnfet_01v8_w500_l500_nf2_4 phi1 mimbot1 VGND phi1 VGND VGND nfet_01v8_w500_l500_nf2
Xsky130_fd_sc_hd__inv_1_0 sky130_fd_sc_hd__inv_1_0/A VGND VPWR sky130_fd_sc_hd__inv_1_2/A
+ VGND VPWR sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_1 sky130_fd_sc_hd__inv_1_1/A VGND VPWR sky130_fd_sc_hd__inv_1_3/A
+ VGND VPWR sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_2 sky130_fd_sc_hd__inv_1_2/A VGND VPWR sky130_fd_sc_hd__inv_1_2/Y
+ VGND VPWR sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_3 sky130_fd_sc_hd__inv_1_3/A VGND VPWR sky130_fd_sc_hd__inv_1_3/Y
+ VGND VPWR sky130_fd_sc_hd__inv_1
.ends

