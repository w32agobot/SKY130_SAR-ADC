magic
tech sky130A
timestamp 1661327437
<< metal2 >>
rect 14 545 334 550
rect 14 513 19 545
rect 51 513 297 545
rect 329 513 334 545
rect 14 421 334 513
rect 14 389 19 421
rect 51 389 297 421
rect 329 389 334 421
rect 14 297 334 389
rect 14 265 19 297
rect 51 265 297 297
rect 329 265 334 297
rect 14 173 334 265
rect 14 141 19 173
rect 51 141 297 173
rect 329 141 334 173
rect 14 49 334 141
rect 14 17 19 49
rect 51 17 297 49
rect 329 17 334 49
rect 14 12 334 17
<< via2 >>
rect 19 513 51 545
rect 297 513 329 545
rect 19 389 51 421
rect 297 389 329 421
rect 19 265 51 297
rect 297 265 329 297
rect 19 141 51 173
rect 297 141 329 173
rect 19 17 51 49
rect 297 17 329 49
<< metal3 >>
rect 16 546 54 548
rect 294 546 332 548
rect 16 545 83 546
rect 16 513 19 545
rect 51 513 83 545
rect 16 512 83 513
rect 265 545 332 546
rect 265 513 297 545
rect 329 513 332 545
rect 265 512 332 513
rect 16 510 54 512
rect 294 510 332 512
rect 16 422 54 424
rect 294 422 332 424
rect 16 421 83 422
rect 16 389 19 421
rect 51 389 83 421
rect 16 388 83 389
rect 265 421 332 422
rect 265 389 297 421
rect 329 389 332 421
rect 265 388 332 389
rect 16 386 54 388
rect 294 386 332 388
rect 16 298 54 300
rect 294 298 332 300
rect 16 297 83 298
rect 16 265 19 297
rect 51 265 83 297
rect 16 264 83 265
rect 265 297 332 298
rect 265 265 297 297
rect 329 265 332 297
rect 265 264 332 265
rect 16 262 54 264
rect 294 262 332 264
rect 16 174 54 176
rect 294 174 332 176
rect 16 173 83 174
rect 16 141 19 173
rect 51 141 83 173
rect 16 140 83 141
rect 265 173 332 174
rect 265 141 297 173
rect 329 141 332 173
rect 265 140 332 141
rect 16 138 54 140
rect 294 138 332 140
rect 16 50 54 52
rect 294 50 332 52
rect 16 49 83 50
rect 16 17 19 49
rect 51 17 83 49
rect 16 16 83 17
rect 265 49 332 50
rect 265 17 297 49
rect 329 17 332 49
rect 265 16 332 17
rect 16 14 54 16
rect 294 14 332 16
<< via3 >>
rect 19 513 51 545
rect 297 513 329 545
rect 19 389 51 421
rect 297 389 329 421
rect 19 265 51 297
rect 297 265 329 297
rect 19 141 51 173
rect 297 141 329 173
rect 19 17 51 49
rect 297 17 329 49
<< metal4 >>
rect 18 545 52 546
rect 18 544 19 545
rect 16 514 19 544
rect 18 513 19 514
rect 51 544 52 545
rect 51 514 130 544
rect 51 513 52 514
rect 18 512 52 513
rect 160 482 190 564
rect 296 545 330 546
rect 296 544 297 545
rect 220 514 297 544
rect 296 513 297 514
rect 329 544 330 545
rect 329 514 332 544
rect 329 513 330 514
rect 296 512 330 513
rect 0 452 348 482
rect 18 421 52 422
rect 18 420 19 421
rect 16 390 19 420
rect 18 389 19 390
rect 51 420 52 421
rect 51 390 130 420
rect 51 389 52 390
rect 18 388 52 389
rect 160 358 190 452
rect 296 421 330 422
rect 296 420 297 421
rect 220 390 297 420
rect 296 389 297 390
rect 329 420 330 421
rect 329 390 332 420
rect 329 389 330 390
rect 296 388 330 389
rect 0 328 348 358
rect 18 297 52 298
rect 18 296 19 297
rect 16 266 19 296
rect 18 265 19 266
rect 51 296 52 297
rect 51 266 130 296
rect 51 265 52 266
rect 18 264 52 265
rect 160 234 190 328
rect 296 297 330 298
rect 296 296 297 297
rect 220 266 297 296
rect 296 265 297 266
rect 329 296 330 297
rect 329 266 332 296
rect 329 265 330 266
rect 296 264 330 265
rect 0 204 348 234
rect 18 173 52 174
rect 18 172 19 173
rect 16 142 19 172
rect 18 141 19 142
rect 51 172 52 173
rect 51 142 130 172
rect 51 141 52 142
rect 18 140 52 141
rect 160 110 190 204
rect 296 173 330 174
rect 296 172 297 173
rect 220 142 297 172
rect 296 141 297 142
rect 329 172 330 173
rect 329 142 332 172
rect 329 141 330 142
rect 296 140 330 141
rect 0 80 348 110
rect 18 49 52 50
rect 18 48 19 49
rect 16 18 19 48
rect 18 17 19 18
rect 51 48 52 49
rect 51 18 130 48
rect 51 17 52 18
rect 18 16 52 17
rect 160 -2 190 80
rect 296 49 330 50
rect 296 48 297 49
rect 220 18 297 48
rect 296 17 297 18
rect 329 48 330 49
rect 329 18 332 48
rect 329 17 330 18
rect 296 16 330 17
<< comment >>
rect 0 550 14 564
rect 334 550 348 564
rect 0 -2 14 12
rect 334 -2 348 12
<< end >>
