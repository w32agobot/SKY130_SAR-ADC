VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO adc_vcm_generator
  CLASS BLOCK ;
  FOREIGN adc_vcm_generator ;
  ORIGIN 0.000 0.000 ;
  SIZE 111.850 BY 380.000 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 6.750 194.150 7.590 194.155 ;
        RECT 12.155 194.150 14.705 194.155 ;
        RECT 6.395 192.925 23.795 194.150 ;
        RECT 6.395 191.320 24.255 192.925 ;
        RECT 6.395 187.105 24.255 188.710 ;
        RECT 7.315 185.885 23.795 187.105 ;
        RECT 7.315 185.880 9.625 185.885 ;
        RECT 14.675 185.880 23.795 185.885 ;
      LAYER li1 ;
        RECT 7.025 192.825 7.315 193.990 ;
        RECT 6.940 192.655 7.400 192.825 ;
        RECT 14.950 192.820 15.240 193.985 ;
        RECT 15.560 192.820 15.890 193.970 ;
        RECT 16.400 192.820 16.730 193.620 ;
        RECT 17.250 192.820 17.490 193.620 ;
        RECT 18.320 192.820 18.650 193.970 ;
        RECT 19.160 192.820 19.490 193.620 ;
        RECT 20.010 192.820 20.250 193.620 ;
        RECT 21.675 192.820 21.885 193.960 ;
        RECT 23.055 192.820 23.265 193.960 ;
        RECT 7.965 192.650 24.065 192.820 ;
        RECT 8.050 191.485 8.340 192.650 ;
        RECT 8.510 191.510 8.770 192.650 ;
        RECT 9.440 191.510 9.720 192.650 ;
        RECT 10.500 192.225 10.885 192.650 ;
        RECT 11.915 192.225 12.300 192.650 ;
        RECT 13.330 192.225 13.715 192.650 ;
        RECT 15.100 192.225 15.485 192.650 ;
        RECT 16.515 192.225 16.900 192.650 ;
        RECT 17.930 192.225 18.315 192.650 ;
        RECT 19.700 192.225 20.085 192.650 ;
        RECT 21.115 192.225 21.500 192.650 ;
        RECT 22.530 192.225 22.915 192.650 ;
        RECT 23.690 191.485 23.980 192.650 ;
        RECT 6.670 187.380 6.960 188.545 ;
        RECT 7.385 187.380 7.595 188.520 ;
        RECT 8.510 187.380 8.790 188.520 ;
        RECT 9.460 187.380 9.720 188.520 ;
        RECT 10.500 187.380 10.885 187.805 ;
        RECT 11.915 187.380 12.300 187.805 ;
        RECT 13.330 187.380 13.715 187.805 ;
        RECT 15.100 187.380 15.485 187.805 ;
        RECT 16.515 187.380 16.900 187.805 ;
        RECT 17.930 187.380 18.315 187.805 ;
        RECT 19.700 187.380 20.085 187.805 ;
        RECT 21.115 187.380 21.500 187.805 ;
        RECT 22.530 187.380 22.915 187.805 ;
        RECT 23.690 187.380 23.980 188.545 ;
        RECT 6.585 187.210 24.065 187.380 ;
        RECT 7.590 186.045 7.880 187.210 ;
        RECT 10.570 186.560 10.745 187.210 ;
        RECT 10.575 184.605 10.745 186.560 ;
        RECT 14.950 186.045 15.240 187.210 ;
        RECT 15.560 186.060 15.890 187.210 ;
        RECT 16.400 186.410 16.730 187.210 ;
        RECT 17.250 186.410 17.490 187.210 ;
        RECT 18.320 186.060 18.650 187.210 ;
        RECT 19.160 186.410 19.490 187.210 ;
        RECT 20.010 186.410 20.250 187.210 ;
        RECT 21.675 186.070 21.885 187.210 ;
        RECT 23.055 186.070 23.265 187.210 ;
        RECT 43.835 180.260 47.835 180.460 ;
        RECT 43.835 179.660 44.235 180.260 ;
        RECT 43.835 179.460 47.835 179.660 ;
        RECT 43.835 178.860 44.235 179.460 ;
        RECT 43.835 178.660 47.835 178.860 ;
        RECT 43.835 178.060 44.235 178.660 ;
        RECT 43.835 177.860 47.835 178.060 ;
        RECT 43.835 177.260 44.235 177.860 ;
        RECT 43.835 177.060 47.835 177.260 ;
        RECT 43.835 176.460 44.235 177.060 ;
        RECT 43.835 176.260 47.835 176.460 ;
        RECT 43.835 175.660 44.235 176.260 ;
        RECT 43.835 175.460 47.835 175.660 ;
        RECT 43.835 174.860 44.235 175.460 ;
        RECT 43.835 174.660 47.835 174.860 ;
        RECT 43.835 174.060 44.235 174.660 ;
        RECT 43.835 173.860 47.835 174.060 ;
        RECT 43.835 173.260 44.235 173.860 ;
        RECT 43.835 173.060 47.835 173.260 ;
        RECT 43.835 172.860 44.235 173.060 ;
        RECT 48.585 172.860 48.785 180.460 ;
        RECT 49.385 172.860 49.585 180.460 ;
        RECT 50.185 172.860 50.385 180.460 ;
        RECT 50.985 172.860 51.185 180.460 ;
        RECT 51.785 172.860 51.985 180.460 ;
        RECT 43.835 172.460 51.985 172.860 ;
        RECT 43.835 172.260 44.235 172.460 ;
        RECT 43.835 172.060 47.835 172.260 ;
        RECT 43.835 171.460 44.235 172.060 ;
        RECT 43.835 171.260 47.835 171.460 ;
        RECT 43.835 170.660 44.235 171.260 ;
        RECT 43.835 170.460 47.835 170.660 ;
        RECT 43.835 169.860 44.235 170.460 ;
        RECT 43.835 169.660 47.835 169.860 ;
        RECT 43.835 169.060 44.235 169.660 ;
        RECT 43.835 168.860 47.835 169.060 ;
        RECT 43.835 168.260 44.235 168.860 ;
        RECT 43.835 168.060 47.835 168.260 ;
        RECT 43.835 167.460 44.235 168.060 ;
        RECT 43.835 167.260 47.835 167.460 ;
        RECT 43.835 166.660 44.235 167.260 ;
        RECT 43.835 166.460 47.835 166.660 ;
        RECT 43.835 165.860 44.235 166.460 ;
        RECT 43.835 165.660 47.835 165.860 ;
        RECT 43.835 165.060 44.235 165.660 ;
        RECT 43.835 164.860 47.835 165.060 ;
        RECT 48.585 164.860 48.785 172.460 ;
        RECT 49.385 164.860 49.585 172.460 ;
        RECT 50.185 164.860 50.385 172.460 ;
        RECT 50.985 164.860 51.185 172.460 ;
        RECT 51.785 164.860 51.985 172.460 ;
        RECT 53.285 172.860 53.485 180.460 ;
        RECT 54.085 172.860 54.285 180.460 ;
        RECT 54.885 172.860 55.085 180.460 ;
        RECT 55.685 172.860 55.885 180.460 ;
        RECT 56.485 172.860 56.685 180.460 ;
        RECT 57.435 180.260 61.435 180.460 ;
        RECT 61.035 179.660 61.435 180.260 ;
        RECT 57.435 179.460 61.435 179.660 ;
        RECT 61.035 178.860 61.435 179.460 ;
        RECT 57.435 178.660 61.435 178.860 ;
        RECT 61.035 178.060 61.435 178.660 ;
        RECT 57.435 177.860 61.435 178.060 ;
        RECT 61.035 177.260 61.435 177.860 ;
        RECT 57.435 177.060 61.435 177.260 ;
        RECT 61.035 176.460 61.435 177.060 ;
        RECT 57.435 176.260 61.435 176.460 ;
        RECT 61.035 175.660 61.435 176.260 ;
        RECT 57.435 175.460 61.435 175.660 ;
        RECT 61.035 174.860 61.435 175.460 ;
        RECT 57.435 174.660 61.435 174.860 ;
        RECT 61.035 174.060 61.435 174.660 ;
        RECT 57.435 173.860 61.435 174.060 ;
        RECT 61.035 173.260 61.435 173.860 ;
        RECT 57.435 173.060 61.435 173.260 ;
        RECT 61.035 172.860 61.435 173.060 ;
        RECT 53.285 172.460 61.435 172.860 ;
        RECT 53.285 164.860 53.485 172.460 ;
        RECT 54.085 164.860 54.285 172.460 ;
        RECT 54.885 164.860 55.085 172.460 ;
        RECT 55.685 164.860 55.885 172.460 ;
        RECT 56.485 164.860 56.685 172.460 ;
        RECT 61.035 172.260 61.435 172.460 ;
        RECT 57.435 172.060 61.435 172.260 ;
        RECT 61.035 171.460 61.435 172.060 ;
        RECT 57.435 171.260 61.435 171.460 ;
        RECT 61.035 170.660 61.435 171.260 ;
        RECT 57.435 170.460 61.435 170.660 ;
        RECT 61.035 169.860 61.435 170.460 ;
        RECT 57.435 169.660 61.435 169.860 ;
        RECT 61.035 169.060 61.435 169.660 ;
        RECT 57.435 168.860 61.435 169.060 ;
        RECT 61.035 168.260 61.435 168.860 ;
        RECT 57.435 168.060 61.435 168.260 ;
        RECT 61.035 167.460 61.435 168.060 ;
        RECT 57.435 167.260 61.435 167.460 ;
        RECT 61.035 166.660 61.435 167.260 ;
        RECT 57.435 166.460 61.435 166.660 ;
        RECT 61.035 165.860 61.435 166.460 ;
        RECT 57.435 165.660 61.435 165.860 ;
        RECT 61.035 165.060 61.435 165.660 ;
        RECT 57.435 164.860 61.435 165.060 ;
        RECT 63.835 180.260 67.835 180.460 ;
        RECT 63.835 179.660 64.235 180.260 ;
        RECT 63.835 179.460 67.835 179.660 ;
        RECT 63.835 178.860 64.235 179.460 ;
        RECT 63.835 178.660 67.835 178.860 ;
        RECT 63.835 178.060 64.235 178.660 ;
        RECT 63.835 177.860 67.835 178.060 ;
        RECT 63.835 177.260 64.235 177.860 ;
        RECT 63.835 177.060 67.835 177.260 ;
        RECT 63.835 176.460 64.235 177.060 ;
        RECT 63.835 176.260 67.835 176.460 ;
        RECT 63.835 175.660 64.235 176.260 ;
        RECT 63.835 175.460 67.835 175.660 ;
        RECT 63.835 174.860 64.235 175.460 ;
        RECT 63.835 174.660 67.835 174.860 ;
        RECT 63.835 174.060 64.235 174.660 ;
        RECT 63.835 173.860 67.835 174.060 ;
        RECT 63.835 173.260 64.235 173.860 ;
        RECT 63.835 173.060 67.835 173.260 ;
        RECT 63.835 172.860 64.235 173.060 ;
        RECT 68.585 172.860 68.785 180.460 ;
        RECT 69.385 172.860 69.585 180.460 ;
        RECT 70.185 172.860 70.385 180.460 ;
        RECT 70.985 172.860 71.185 180.460 ;
        RECT 71.785 172.860 71.985 180.460 ;
        RECT 63.835 172.460 71.985 172.860 ;
        RECT 63.835 172.260 64.235 172.460 ;
        RECT 63.835 172.060 67.835 172.260 ;
        RECT 63.835 171.460 64.235 172.060 ;
        RECT 63.835 171.260 67.835 171.460 ;
        RECT 63.835 170.660 64.235 171.260 ;
        RECT 63.835 170.460 67.835 170.660 ;
        RECT 63.835 169.860 64.235 170.460 ;
        RECT 63.835 169.660 67.835 169.860 ;
        RECT 63.835 169.060 64.235 169.660 ;
        RECT 63.835 168.860 67.835 169.060 ;
        RECT 63.835 168.260 64.235 168.860 ;
        RECT 63.835 168.060 67.835 168.260 ;
        RECT 63.835 167.460 64.235 168.060 ;
        RECT 63.835 167.260 67.835 167.460 ;
        RECT 63.835 166.660 64.235 167.260 ;
        RECT 63.835 166.460 67.835 166.660 ;
        RECT 63.835 165.860 64.235 166.460 ;
        RECT 63.835 165.660 67.835 165.860 ;
        RECT 63.835 165.060 64.235 165.660 ;
        RECT 63.835 164.860 67.835 165.060 ;
        RECT 68.585 164.860 68.785 172.460 ;
        RECT 69.385 164.860 69.585 172.460 ;
        RECT 70.185 164.860 70.385 172.460 ;
        RECT 70.985 164.860 71.185 172.460 ;
        RECT 71.785 164.860 71.985 172.460 ;
        RECT 73.285 172.860 73.485 180.460 ;
        RECT 74.085 172.860 74.285 180.460 ;
        RECT 74.885 172.860 75.085 180.460 ;
        RECT 75.685 172.860 75.885 180.460 ;
        RECT 76.485 172.860 76.685 180.460 ;
        RECT 77.435 180.260 81.435 180.460 ;
        RECT 81.035 179.660 81.435 180.260 ;
        RECT 77.435 179.460 81.435 179.660 ;
        RECT 81.035 178.860 81.435 179.460 ;
        RECT 77.435 178.660 81.435 178.860 ;
        RECT 81.035 178.060 81.435 178.660 ;
        RECT 77.435 177.860 81.435 178.060 ;
        RECT 81.035 177.260 81.435 177.860 ;
        RECT 77.435 177.060 81.435 177.260 ;
        RECT 81.035 176.460 81.435 177.060 ;
        RECT 77.435 176.260 81.435 176.460 ;
        RECT 81.035 175.660 81.435 176.260 ;
        RECT 77.435 175.460 81.435 175.660 ;
        RECT 81.035 174.860 81.435 175.460 ;
        RECT 77.435 174.660 81.435 174.860 ;
        RECT 81.035 174.060 81.435 174.660 ;
        RECT 77.435 173.860 81.435 174.060 ;
        RECT 81.035 173.260 81.435 173.860 ;
        RECT 77.435 173.060 81.435 173.260 ;
        RECT 81.035 172.860 81.435 173.060 ;
        RECT 73.285 172.460 81.435 172.860 ;
        RECT 73.285 164.860 73.485 172.460 ;
        RECT 74.085 164.860 74.285 172.460 ;
        RECT 74.885 164.860 75.085 172.460 ;
        RECT 75.685 164.860 75.885 172.460 ;
        RECT 76.485 164.860 76.685 172.460 ;
        RECT 81.035 172.260 81.435 172.460 ;
        RECT 77.435 172.060 81.435 172.260 ;
        RECT 81.035 171.460 81.435 172.060 ;
        RECT 77.435 171.260 81.435 171.460 ;
        RECT 81.035 170.660 81.435 171.260 ;
        RECT 77.435 170.460 81.435 170.660 ;
        RECT 81.035 169.860 81.435 170.460 ;
        RECT 77.435 169.660 81.435 169.860 ;
        RECT 81.035 169.060 81.435 169.660 ;
        RECT 77.435 168.860 81.435 169.060 ;
        RECT 81.035 168.260 81.435 168.860 ;
        RECT 77.435 168.060 81.435 168.260 ;
        RECT 81.035 167.460 81.435 168.060 ;
        RECT 77.435 167.260 81.435 167.460 ;
        RECT 81.035 166.660 81.435 167.260 ;
        RECT 77.435 166.460 81.435 166.660 ;
        RECT 81.035 165.860 81.435 166.460 ;
        RECT 77.435 165.660 81.435 165.860 ;
        RECT 81.035 165.060 81.435 165.660 ;
        RECT 77.435 164.860 81.435 165.060 ;
        RECT 83.835 180.260 87.835 180.460 ;
        RECT 83.835 179.660 84.235 180.260 ;
        RECT 83.835 179.460 87.835 179.660 ;
        RECT 83.835 178.860 84.235 179.460 ;
        RECT 83.835 178.660 87.835 178.860 ;
        RECT 83.835 178.060 84.235 178.660 ;
        RECT 83.835 177.860 87.835 178.060 ;
        RECT 83.835 177.260 84.235 177.860 ;
        RECT 83.835 177.060 87.835 177.260 ;
        RECT 83.835 176.460 84.235 177.060 ;
        RECT 83.835 176.260 87.835 176.460 ;
        RECT 83.835 175.660 84.235 176.260 ;
        RECT 83.835 175.460 87.835 175.660 ;
        RECT 83.835 174.860 84.235 175.460 ;
        RECT 83.835 174.660 87.835 174.860 ;
        RECT 83.835 174.060 84.235 174.660 ;
        RECT 83.835 173.860 87.835 174.060 ;
        RECT 83.835 173.260 84.235 173.860 ;
        RECT 83.835 173.060 87.835 173.260 ;
        RECT 83.835 172.860 84.235 173.060 ;
        RECT 88.585 172.860 88.785 180.460 ;
        RECT 89.385 172.860 89.585 180.460 ;
        RECT 90.185 172.860 90.385 180.460 ;
        RECT 90.985 172.860 91.185 180.460 ;
        RECT 91.785 172.860 91.985 180.460 ;
        RECT 83.835 172.460 91.985 172.860 ;
        RECT 83.835 172.260 84.235 172.460 ;
        RECT 83.835 172.060 87.835 172.260 ;
        RECT 83.835 171.460 84.235 172.060 ;
        RECT 83.835 171.260 87.835 171.460 ;
        RECT 83.835 170.660 84.235 171.260 ;
        RECT 83.835 170.460 87.835 170.660 ;
        RECT 83.835 169.860 84.235 170.460 ;
        RECT 83.835 169.660 87.835 169.860 ;
        RECT 83.835 169.060 84.235 169.660 ;
        RECT 83.835 168.860 87.835 169.060 ;
        RECT 83.835 168.260 84.235 168.860 ;
        RECT 83.835 168.060 87.835 168.260 ;
        RECT 83.835 167.460 84.235 168.060 ;
        RECT 83.835 167.260 87.835 167.460 ;
        RECT 83.835 166.660 84.235 167.260 ;
        RECT 83.835 166.460 87.835 166.660 ;
        RECT 83.835 165.860 84.235 166.460 ;
        RECT 83.835 165.660 87.835 165.860 ;
        RECT 83.835 165.060 84.235 165.660 ;
        RECT 83.835 164.860 87.835 165.060 ;
        RECT 88.585 164.860 88.785 172.460 ;
        RECT 89.385 164.860 89.585 172.460 ;
        RECT 90.185 164.860 90.385 172.460 ;
        RECT 90.985 164.860 91.185 172.460 ;
        RECT 91.785 164.860 91.985 172.460 ;
        RECT 93.285 172.860 93.485 180.460 ;
        RECT 94.085 172.860 94.285 180.460 ;
        RECT 94.885 172.860 95.085 180.460 ;
        RECT 95.685 172.860 95.885 180.460 ;
        RECT 96.485 172.860 96.685 180.460 ;
        RECT 97.435 180.260 101.435 180.460 ;
        RECT 101.035 179.660 101.435 180.260 ;
        RECT 97.435 179.460 101.435 179.660 ;
        RECT 101.035 178.860 101.435 179.460 ;
        RECT 97.435 178.660 101.435 178.860 ;
        RECT 101.035 178.060 101.435 178.660 ;
        RECT 97.435 177.860 101.435 178.060 ;
        RECT 101.035 177.260 101.435 177.860 ;
        RECT 97.435 177.060 101.435 177.260 ;
        RECT 101.035 176.460 101.435 177.060 ;
        RECT 97.435 176.260 101.435 176.460 ;
        RECT 101.035 175.660 101.435 176.260 ;
        RECT 97.435 175.460 101.435 175.660 ;
        RECT 101.035 174.860 101.435 175.460 ;
        RECT 97.435 174.660 101.435 174.860 ;
        RECT 101.035 174.060 101.435 174.660 ;
        RECT 97.435 173.860 101.435 174.060 ;
        RECT 101.035 173.260 101.435 173.860 ;
        RECT 97.435 173.060 101.435 173.260 ;
        RECT 101.035 172.860 101.435 173.060 ;
        RECT 93.285 172.460 101.435 172.860 ;
        RECT 93.285 164.860 93.485 172.460 ;
        RECT 94.085 164.860 94.285 172.460 ;
        RECT 94.885 164.860 95.085 172.460 ;
        RECT 95.685 164.860 95.885 172.460 ;
        RECT 96.485 164.860 96.685 172.460 ;
        RECT 101.035 172.260 101.435 172.460 ;
        RECT 97.435 172.060 101.435 172.260 ;
        RECT 101.035 171.460 101.435 172.060 ;
        RECT 97.435 171.260 101.435 171.460 ;
        RECT 101.035 170.660 101.435 171.260 ;
        RECT 97.435 170.460 101.435 170.660 ;
        RECT 101.035 169.860 101.435 170.460 ;
        RECT 97.435 169.660 101.435 169.860 ;
        RECT 101.035 169.060 101.435 169.660 ;
        RECT 97.435 168.860 101.435 169.060 ;
        RECT 101.035 168.260 101.435 168.860 ;
        RECT 97.435 168.060 101.435 168.260 ;
        RECT 101.035 167.460 101.435 168.060 ;
        RECT 97.435 167.260 101.435 167.460 ;
        RECT 101.035 166.660 101.435 167.260 ;
        RECT 97.435 166.460 101.435 166.660 ;
        RECT 101.035 165.860 101.435 166.460 ;
        RECT 97.435 165.660 101.435 165.860 ;
        RECT 101.035 165.060 101.435 165.660 ;
        RECT 97.435 164.860 101.435 165.060 ;
      LAYER mcon ;
        RECT 7.085 192.655 7.255 192.825 ;
        RECT 8.110 192.650 8.280 192.820 ;
        RECT 8.570 192.650 8.740 192.820 ;
        RECT 9.030 192.650 9.200 192.820 ;
        RECT 9.490 192.650 9.660 192.820 ;
        RECT 9.950 192.650 10.120 192.820 ;
        RECT 10.410 192.650 10.580 192.820 ;
        RECT 10.870 192.650 11.040 192.820 ;
        RECT 11.330 192.650 11.500 192.820 ;
        RECT 11.790 192.650 11.960 192.820 ;
        RECT 12.250 192.650 12.420 192.820 ;
        RECT 12.710 192.650 12.880 192.820 ;
        RECT 13.170 192.650 13.340 192.820 ;
        RECT 13.630 192.650 13.800 192.820 ;
        RECT 14.090 192.650 14.260 192.820 ;
        RECT 14.550 192.650 14.720 192.820 ;
        RECT 15.010 192.650 15.180 192.820 ;
        RECT 15.470 192.650 15.640 192.820 ;
        RECT 15.930 192.650 16.100 192.820 ;
        RECT 16.390 192.650 16.560 192.820 ;
        RECT 16.850 192.650 17.020 192.820 ;
        RECT 17.310 192.650 17.480 192.820 ;
        RECT 17.770 192.650 17.940 192.820 ;
        RECT 18.230 192.650 18.400 192.820 ;
        RECT 18.690 192.650 18.860 192.820 ;
        RECT 19.150 192.650 19.320 192.820 ;
        RECT 19.610 192.650 19.780 192.820 ;
        RECT 20.070 192.650 20.240 192.820 ;
        RECT 20.530 192.650 20.700 192.820 ;
        RECT 20.990 192.650 21.160 192.820 ;
        RECT 21.450 192.650 21.620 192.820 ;
        RECT 21.910 192.650 22.080 192.820 ;
        RECT 22.370 192.650 22.540 192.820 ;
        RECT 22.830 192.650 23.000 192.820 ;
        RECT 23.290 192.650 23.460 192.820 ;
        RECT 23.750 192.650 23.920 192.820 ;
        RECT 6.730 187.210 6.900 187.380 ;
        RECT 7.190 187.210 7.360 187.380 ;
        RECT 7.650 187.210 7.820 187.380 ;
        RECT 8.110 187.210 8.280 187.380 ;
        RECT 8.570 187.210 8.740 187.380 ;
        RECT 9.030 187.210 9.200 187.380 ;
        RECT 9.490 187.210 9.660 187.380 ;
        RECT 9.950 187.210 10.120 187.380 ;
        RECT 10.410 187.210 10.580 187.380 ;
        RECT 10.870 187.210 11.040 187.380 ;
        RECT 11.330 187.210 11.500 187.380 ;
        RECT 11.790 187.210 11.960 187.380 ;
        RECT 12.250 187.210 12.420 187.380 ;
        RECT 12.710 187.210 12.880 187.380 ;
        RECT 13.170 187.210 13.340 187.380 ;
        RECT 13.630 187.210 13.800 187.380 ;
        RECT 14.090 187.210 14.260 187.380 ;
        RECT 14.550 187.210 14.720 187.380 ;
        RECT 15.010 187.210 15.180 187.380 ;
        RECT 15.470 187.210 15.640 187.380 ;
        RECT 15.930 187.210 16.100 187.380 ;
        RECT 16.390 187.210 16.560 187.380 ;
        RECT 16.850 187.210 17.020 187.380 ;
        RECT 17.310 187.210 17.480 187.380 ;
        RECT 17.770 187.210 17.940 187.380 ;
        RECT 18.230 187.210 18.400 187.380 ;
        RECT 18.690 187.210 18.860 187.380 ;
        RECT 19.150 187.210 19.320 187.380 ;
        RECT 19.610 187.210 19.780 187.380 ;
        RECT 20.070 187.210 20.240 187.380 ;
        RECT 20.530 187.210 20.700 187.380 ;
        RECT 20.990 187.210 21.160 187.380 ;
        RECT 21.450 187.210 21.620 187.380 ;
        RECT 21.910 187.210 22.080 187.380 ;
        RECT 22.370 187.210 22.540 187.380 ;
        RECT 22.830 187.210 23.000 187.380 ;
        RECT 23.290 187.210 23.460 187.380 ;
        RECT 23.750 187.210 23.920 187.380 ;
        RECT 43.885 176.960 44.185 177.410 ;
        RECT 43.885 176.210 44.185 176.660 ;
        RECT 43.885 175.460 44.185 175.910 ;
        RECT 43.885 174.710 44.185 175.160 ;
        RECT 43.885 173.960 44.185 174.410 ;
        RECT 43.885 173.210 44.185 173.660 ;
        RECT 43.885 172.460 44.185 172.910 ;
        RECT 43.885 171.710 44.185 172.160 ;
        RECT 43.885 170.960 44.185 171.410 ;
        RECT 43.885 170.210 44.185 170.660 ;
        RECT 43.885 169.460 44.185 169.910 ;
        RECT 43.885 168.710 44.185 169.160 ;
        RECT 43.885 167.960 44.185 168.410 ;
        RECT 61.085 176.960 61.385 177.410 ;
        RECT 61.085 176.210 61.385 176.660 ;
        RECT 61.085 175.460 61.385 175.910 ;
        RECT 61.085 174.710 61.385 175.160 ;
        RECT 61.085 173.960 61.385 174.410 ;
        RECT 61.085 173.210 61.385 173.660 ;
        RECT 61.085 172.460 61.385 172.910 ;
        RECT 61.085 171.710 61.385 172.160 ;
        RECT 61.085 170.960 61.385 171.410 ;
        RECT 61.085 170.210 61.385 170.660 ;
        RECT 61.085 169.460 61.385 169.910 ;
        RECT 61.085 168.710 61.385 169.160 ;
        RECT 61.085 167.960 61.385 168.410 ;
        RECT 63.885 176.960 64.185 177.410 ;
        RECT 63.885 176.210 64.185 176.660 ;
        RECT 63.885 175.460 64.185 175.910 ;
        RECT 63.885 174.710 64.185 175.160 ;
        RECT 63.885 173.960 64.185 174.410 ;
        RECT 63.885 173.210 64.185 173.660 ;
        RECT 63.885 172.460 64.185 172.910 ;
        RECT 63.885 171.710 64.185 172.160 ;
        RECT 63.885 170.960 64.185 171.410 ;
        RECT 63.885 170.210 64.185 170.660 ;
        RECT 63.885 169.460 64.185 169.910 ;
        RECT 63.885 168.710 64.185 169.160 ;
        RECT 63.885 167.960 64.185 168.410 ;
        RECT 81.085 176.960 81.385 177.410 ;
        RECT 81.085 176.210 81.385 176.660 ;
        RECT 81.085 175.460 81.385 175.910 ;
        RECT 81.085 174.710 81.385 175.160 ;
        RECT 81.085 173.960 81.385 174.410 ;
        RECT 81.085 173.210 81.385 173.660 ;
        RECT 81.085 172.460 81.385 172.910 ;
        RECT 81.085 171.710 81.385 172.160 ;
        RECT 81.085 170.960 81.385 171.410 ;
        RECT 81.085 170.210 81.385 170.660 ;
        RECT 81.085 169.460 81.385 169.910 ;
        RECT 81.085 168.710 81.385 169.160 ;
        RECT 81.085 167.960 81.385 168.410 ;
        RECT 83.885 176.960 84.185 177.410 ;
        RECT 83.885 176.210 84.185 176.660 ;
        RECT 83.885 175.460 84.185 175.910 ;
        RECT 83.885 174.710 84.185 175.160 ;
        RECT 83.885 173.960 84.185 174.410 ;
        RECT 83.885 173.210 84.185 173.660 ;
        RECT 83.885 172.460 84.185 172.910 ;
        RECT 83.885 171.710 84.185 172.160 ;
        RECT 83.885 170.960 84.185 171.410 ;
        RECT 83.885 170.210 84.185 170.660 ;
        RECT 83.885 169.460 84.185 169.910 ;
        RECT 83.885 168.710 84.185 169.160 ;
        RECT 83.885 167.960 84.185 168.410 ;
        RECT 101.085 176.960 101.385 177.410 ;
        RECT 101.085 176.210 101.385 176.660 ;
        RECT 101.085 175.460 101.385 175.910 ;
        RECT 101.085 174.710 101.385 175.160 ;
        RECT 101.085 173.960 101.385 174.410 ;
        RECT 101.085 173.210 101.385 173.660 ;
        RECT 101.085 172.460 101.385 172.910 ;
        RECT 101.085 171.710 101.385 172.160 ;
        RECT 101.085 170.960 101.385 171.410 ;
        RECT 101.085 170.210 101.385 170.660 ;
        RECT 101.085 169.460 101.385 169.910 ;
        RECT 101.085 168.710 101.385 169.160 ;
        RECT 101.085 167.960 101.385 168.410 ;
      LAYER met1 ;
        RECT 16.435 198.760 22.105 198.765 ;
        RECT 0.000 197.485 109.510 198.760 ;
        RECT 6.940 192.975 7.400 192.980 ;
        RECT 0.000 192.495 24.065 192.975 ;
        RECT 0.000 187.055 24.065 187.535 ;
        RECT 49.435 181.460 55.835 182.660 ;
        RECT 69.435 181.460 75.835 182.660 ;
        RECT 89.435 181.460 95.835 182.660 ;
        RECT 52.135 180.810 53.135 181.460 ;
        RECT 72.135 180.810 73.135 181.460 ;
        RECT 92.135 180.810 93.135 181.460 ;
        RECT 48.785 180.660 56.485 180.810 ;
        RECT 68.785 180.660 76.485 180.810 ;
        RECT 88.785 180.660 96.485 180.810 ;
        RECT 43.835 175.860 44.585 177.660 ;
        RECT 42.635 173.110 44.585 175.860 ;
        RECT 42.635 172.210 42.785 173.110 ;
        RECT 43.435 172.960 44.585 173.110 ;
        RECT 44.735 172.960 44.885 180.510 ;
        RECT 45.335 172.960 45.485 180.510 ;
        RECT 45.935 172.960 46.085 180.510 ;
        RECT 46.535 172.960 46.685 180.510 ;
        RECT 47.135 172.960 47.285 180.510 ;
        RECT 47.735 172.960 47.885 180.510 ;
        RECT 52.135 180.210 53.135 180.660 ;
        RECT 48.785 180.060 56.485 180.210 ;
        RECT 52.135 179.610 53.135 180.060 ;
        RECT 48.785 179.460 56.485 179.610 ;
        RECT 52.135 179.010 53.135 179.460 ;
        RECT 48.785 178.860 56.485 179.010 ;
        RECT 52.135 178.410 53.135 178.860 ;
        RECT 48.785 178.260 56.485 178.410 ;
        RECT 52.135 177.810 53.135 178.260 ;
        RECT 48.785 177.660 56.485 177.810 ;
        RECT 52.135 177.210 53.135 177.660 ;
        RECT 48.785 177.060 56.485 177.210 ;
        RECT 52.135 176.610 53.135 177.060 ;
        RECT 48.785 176.460 56.485 176.610 ;
        RECT 52.135 176.010 53.135 176.460 ;
        RECT 48.785 175.860 56.485 176.010 ;
        RECT 52.135 175.410 53.135 175.860 ;
        RECT 48.785 175.260 56.485 175.410 ;
        RECT 52.135 174.810 53.135 175.260 ;
        RECT 48.785 174.660 56.485 174.810 ;
        RECT 52.135 174.210 53.135 174.660 ;
        RECT 48.785 174.060 56.485 174.210 ;
        RECT 52.135 173.610 53.135 174.060 ;
        RECT 48.785 173.460 56.485 173.610 ;
        RECT 52.135 172.960 53.135 173.460 ;
        RECT 57.385 172.960 57.535 180.510 ;
        RECT 57.985 172.960 58.135 180.510 ;
        RECT 58.585 172.960 58.735 180.510 ;
        RECT 59.185 172.960 59.335 180.510 ;
        RECT 59.785 172.960 59.935 180.510 ;
        RECT 60.385 172.960 60.535 180.510 ;
        RECT 60.685 175.860 61.435 177.660 ;
        RECT 63.835 175.860 64.585 177.660 ;
        RECT 60.685 173.110 64.585 175.860 ;
        RECT 60.685 172.960 61.835 173.110 ;
        RECT 43.435 172.360 61.835 172.960 ;
        RECT 43.435 172.210 44.585 172.360 ;
        RECT 42.635 169.460 44.585 172.210 ;
        RECT 43.835 167.710 44.585 169.460 ;
        RECT 44.735 164.810 44.885 172.360 ;
        RECT 45.335 164.810 45.485 172.360 ;
        RECT 45.935 164.810 46.085 172.360 ;
        RECT 46.535 164.810 46.685 172.360 ;
        RECT 47.135 164.810 47.285 172.360 ;
        RECT 47.735 164.810 47.885 172.360 ;
        RECT 52.135 171.860 53.135 172.360 ;
        RECT 48.785 171.710 56.485 171.860 ;
        RECT 52.135 171.260 53.135 171.710 ;
        RECT 48.785 171.110 56.485 171.260 ;
        RECT 52.135 170.660 53.135 171.110 ;
        RECT 48.785 170.510 56.485 170.660 ;
        RECT 52.135 170.060 53.135 170.510 ;
        RECT 48.785 169.910 56.485 170.060 ;
        RECT 52.135 169.460 53.135 169.910 ;
        RECT 48.785 169.310 56.485 169.460 ;
        RECT 52.135 168.860 53.135 169.310 ;
        RECT 48.785 168.710 56.485 168.860 ;
        RECT 52.135 168.260 53.135 168.710 ;
        RECT 48.785 168.110 56.485 168.260 ;
        RECT 52.135 167.660 53.135 168.110 ;
        RECT 48.785 167.510 56.485 167.660 ;
        RECT 52.135 167.060 53.135 167.510 ;
        RECT 48.785 166.910 56.485 167.060 ;
        RECT 52.135 166.460 53.135 166.910 ;
        RECT 48.785 166.310 56.485 166.460 ;
        RECT 52.135 165.860 53.135 166.310 ;
        RECT 48.785 165.710 56.485 165.860 ;
        RECT 52.135 165.260 53.135 165.710 ;
        RECT 48.785 165.110 56.485 165.260 ;
        RECT 52.135 164.660 53.135 165.110 ;
        RECT 57.385 164.810 57.535 172.360 ;
        RECT 57.985 164.810 58.135 172.360 ;
        RECT 58.585 164.810 58.735 172.360 ;
        RECT 59.185 164.810 59.335 172.360 ;
        RECT 59.785 164.810 59.935 172.360 ;
        RECT 60.385 164.810 60.535 172.360 ;
        RECT 60.685 172.210 61.835 172.360 ;
        RECT 62.485 172.210 62.785 173.110 ;
        RECT 63.435 172.960 64.585 173.110 ;
        RECT 64.735 172.960 64.885 180.510 ;
        RECT 65.335 172.960 65.485 180.510 ;
        RECT 65.935 172.960 66.085 180.510 ;
        RECT 66.535 172.960 66.685 180.510 ;
        RECT 67.135 172.960 67.285 180.510 ;
        RECT 67.735 172.960 67.885 180.510 ;
        RECT 72.135 180.210 73.135 180.660 ;
        RECT 68.785 180.060 76.485 180.210 ;
        RECT 72.135 179.610 73.135 180.060 ;
        RECT 68.785 179.460 76.485 179.610 ;
        RECT 72.135 179.010 73.135 179.460 ;
        RECT 68.785 178.860 76.485 179.010 ;
        RECT 72.135 178.410 73.135 178.860 ;
        RECT 68.785 178.260 76.485 178.410 ;
        RECT 72.135 177.810 73.135 178.260 ;
        RECT 68.785 177.660 76.485 177.810 ;
        RECT 72.135 177.210 73.135 177.660 ;
        RECT 68.785 177.060 76.485 177.210 ;
        RECT 72.135 176.610 73.135 177.060 ;
        RECT 68.785 176.460 76.485 176.610 ;
        RECT 72.135 176.010 73.135 176.460 ;
        RECT 68.785 175.860 76.485 176.010 ;
        RECT 72.135 175.410 73.135 175.860 ;
        RECT 68.785 175.260 76.485 175.410 ;
        RECT 72.135 174.810 73.135 175.260 ;
        RECT 68.785 174.660 76.485 174.810 ;
        RECT 72.135 174.210 73.135 174.660 ;
        RECT 68.785 174.060 76.485 174.210 ;
        RECT 72.135 173.610 73.135 174.060 ;
        RECT 68.785 173.460 76.485 173.610 ;
        RECT 72.135 172.960 73.135 173.460 ;
        RECT 77.385 172.960 77.535 180.510 ;
        RECT 77.985 172.960 78.135 180.510 ;
        RECT 78.585 172.960 78.735 180.510 ;
        RECT 79.185 172.960 79.335 180.510 ;
        RECT 79.785 172.960 79.935 180.510 ;
        RECT 80.385 172.960 80.535 180.510 ;
        RECT 80.685 175.860 81.435 177.660 ;
        RECT 83.835 175.860 84.585 177.660 ;
        RECT 80.685 173.110 84.585 175.860 ;
        RECT 80.685 172.960 81.835 173.110 ;
        RECT 63.435 172.360 81.835 172.960 ;
        RECT 63.435 172.210 64.585 172.360 ;
        RECT 60.685 169.460 64.585 172.210 ;
        RECT 60.685 167.710 61.435 169.460 ;
        RECT 63.835 167.710 64.585 169.460 ;
        RECT 64.735 164.810 64.885 172.360 ;
        RECT 65.335 164.810 65.485 172.360 ;
        RECT 65.935 164.810 66.085 172.360 ;
        RECT 66.535 164.810 66.685 172.360 ;
        RECT 67.135 164.810 67.285 172.360 ;
        RECT 67.735 164.810 67.885 172.360 ;
        RECT 72.135 171.860 73.135 172.360 ;
        RECT 68.785 171.710 76.485 171.860 ;
        RECT 72.135 171.260 73.135 171.710 ;
        RECT 68.785 171.110 76.485 171.260 ;
        RECT 72.135 170.660 73.135 171.110 ;
        RECT 68.785 170.510 76.485 170.660 ;
        RECT 72.135 170.060 73.135 170.510 ;
        RECT 68.785 169.910 76.485 170.060 ;
        RECT 72.135 169.460 73.135 169.910 ;
        RECT 68.785 169.310 76.485 169.460 ;
        RECT 72.135 168.860 73.135 169.310 ;
        RECT 68.785 168.710 76.485 168.860 ;
        RECT 72.135 168.260 73.135 168.710 ;
        RECT 68.785 168.110 76.485 168.260 ;
        RECT 72.135 167.660 73.135 168.110 ;
        RECT 68.785 167.510 76.485 167.660 ;
        RECT 72.135 167.060 73.135 167.510 ;
        RECT 68.785 166.910 76.485 167.060 ;
        RECT 72.135 166.460 73.135 166.910 ;
        RECT 68.785 166.310 76.485 166.460 ;
        RECT 72.135 165.860 73.135 166.310 ;
        RECT 68.785 165.710 76.485 165.860 ;
        RECT 72.135 165.260 73.135 165.710 ;
        RECT 68.785 165.110 76.485 165.260 ;
        RECT 72.135 164.660 73.135 165.110 ;
        RECT 77.385 164.810 77.535 172.360 ;
        RECT 77.985 164.810 78.135 172.360 ;
        RECT 78.585 164.810 78.735 172.360 ;
        RECT 79.185 164.810 79.335 172.360 ;
        RECT 79.785 164.810 79.935 172.360 ;
        RECT 80.385 164.810 80.535 172.360 ;
        RECT 80.685 172.210 81.835 172.360 ;
        RECT 82.485 172.210 82.785 173.110 ;
        RECT 83.435 172.960 84.585 173.110 ;
        RECT 84.735 172.960 84.885 180.510 ;
        RECT 85.335 172.960 85.485 180.510 ;
        RECT 85.935 172.960 86.085 180.510 ;
        RECT 86.535 172.960 86.685 180.510 ;
        RECT 87.135 172.960 87.285 180.510 ;
        RECT 87.735 172.960 87.885 180.510 ;
        RECT 92.135 180.210 93.135 180.660 ;
        RECT 88.785 180.060 96.485 180.210 ;
        RECT 92.135 179.610 93.135 180.060 ;
        RECT 88.785 179.460 96.485 179.610 ;
        RECT 92.135 179.010 93.135 179.460 ;
        RECT 88.785 178.860 96.485 179.010 ;
        RECT 92.135 178.410 93.135 178.860 ;
        RECT 88.785 178.260 96.485 178.410 ;
        RECT 92.135 177.810 93.135 178.260 ;
        RECT 88.785 177.660 96.485 177.810 ;
        RECT 92.135 177.210 93.135 177.660 ;
        RECT 88.785 177.060 96.485 177.210 ;
        RECT 92.135 176.610 93.135 177.060 ;
        RECT 88.785 176.460 96.485 176.610 ;
        RECT 92.135 176.010 93.135 176.460 ;
        RECT 88.785 175.860 96.485 176.010 ;
        RECT 92.135 175.410 93.135 175.860 ;
        RECT 88.785 175.260 96.485 175.410 ;
        RECT 92.135 174.810 93.135 175.260 ;
        RECT 88.785 174.660 96.485 174.810 ;
        RECT 92.135 174.210 93.135 174.660 ;
        RECT 88.785 174.060 96.485 174.210 ;
        RECT 92.135 173.610 93.135 174.060 ;
        RECT 88.785 173.460 96.485 173.610 ;
        RECT 92.135 172.960 93.135 173.460 ;
        RECT 97.385 172.960 97.535 180.510 ;
        RECT 97.985 172.960 98.135 180.510 ;
        RECT 98.585 172.960 98.735 180.510 ;
        RECT 99.185 172.960 99.335 180.510 ;
        RECT 99.785 172.960 99.935 180.510 ;
        RECT 100.385 172.960 100.535 180.510 ;
        RECT 100.685 175.860 101.435 177.660 ;
        RECT 100.685 173.510 102.635 175.860 ;
        RECT 100.685 173.110 109.510 173.510 ;
        RECT 100.685 172.960 101.835 173.110 ;
        RECT 83.435 172.360 101.835 172.960 ;
        RECT 83.435 172.210 84.585 172.360 ;
        RECT 80.685 169.460 84.585 172.210 ;
        RECT 80.685 167.710 81.435 169.460 ;
        RECT 83.835 167.710 84.585 169.460 ;
        RECT 84.735 164.810 84.885 172.360 ;
        RECT 85.335 164.810 85.485 172.360 ;
        RECT 85.935 164.810 86.085 172.360 ;
        RECT 86.535 164.810 86.685 172.360 ;
        RECT 87.135 164.810 87.285 172.360 ;
        RECT 87.735 164.810 87.885 172.360 ;
        RECT 92.135 171.860 93.135 172.360 ;
        RECT 88.785 171.710 96.485 171.860 ;
        RECT 92.135 171.260 93.135 171.710 ;
        RECT 88.785 171.110 96.485 171.260 ;
        RECT 92.135 170.660 93.135 171.110 ;
        RECT 88.785 170.510 96.485 170.660 ;
        RECT 92.135 170.060 93.135 170.510 ;
        RECT 88.785 169.910 96.485 170.060 ;
        RECT 92.135 169.460 93.135 169.910 ;
        RECT 88.785 169.310 96.485 169.460 ;
        RECT 92.135 168.860 93.135 169.310 ;
        RECT 88.785 168.710 96.485 168.860 ;
        RECT 92.135 168.260 93.135 168.710 ;
        RECT 88.785 168.110 96.485 168.260 ;
        RECT 92.135 167.660 93.135 168.110 ;
        RECT 88.785 167.510 96.485 167.660 ;
        RECT 92.135 167.060 93.135 167.510 ;
        RECT 88.785 166.910 96.485 167.060 ;
        RECT 92.135 166.460 93.135 166.910 ;
        RECT 88.785 166.310 96.485 166.460 ;
        RECT 92.135 165.860 93.135 166.310 ;
        RECT 88.785 165.710 96.485 165.860 ;
        RECT 92.135 165.260 93.135 165.710 ;
        RECT 88.785 165.110 96.485 165.260 ;
        RECT 92.135 164.660 93.135 165.110 ;
        RECT 97.385 164.810 97.535 172.360 ;
        RECT 97.985 164.810 98.135 172.360 ;
        RECT 98.585 164.810 98.735 172.360 ;
        RECT 99.185 164.810 99.335 172.360 ;
        RECT 99.785 164.810 99.935 172.360 ;
        RECT 100.385 164.810 100.535 172.360 ;
        RECT 100.685 172.210 101.835 172.360 ;
        RECT 102.485 172.235 109.510 173.110 ;
        RECT 102.485 172.210 102.635 172.235 ;
        RECT 100.685 169.460 102.635 172.210 ;
        RECT 100.685 167.710 101.435 169.460 ;
        RECT 48.785 164.510 56.485 164.660 ;
        RECT 68.785 164.510 76.485 164.660 ;
        RECT 88.785 164.510 96.485 164.660 ;
        RECT 52.135 163.860 53.135 164.510 ;
        RECT 72.135 163.860 73.135 164.510 ;
        RECT 92.135 163.860 93.135 164.510 ;
        RECT 49.435 162.660 55.835 163.860 ;
        RECT 69.435 162.660 75.835 163.860 ;
        RECT 89.435 162.660 95.835 163.860 ;
      LAYER via ;
        RECT 0.160 198.305 0.560 198.705 ;
        RECT 0.785 198.305 1.185 198.705 ;
        RECT 1.410 198.305 1.810 198.705 ;
        RECT 107.675 198.230 108.075 198.630 ;
        RECT 108.300 198.230 108.700 198.630 ;
        RECT 108.925 198.230 109.325 198.630 ;
        RECT 0.160 197.775 0.560 198.175 ;
        RECT 0.785 197.775 1.185 198.175 ;
        RECT 1.410 197.775 1.810 198.175 ;
        RECT 107.670 197.630 108.070 198.030 ;
        RECT 108.295 197.630 108.695 198.030 ;
        RECT 108.920 197.630 109.320 198.030 ;
        RECT 0.080 192.540 0.490 192.930 ;
        RECT 0.650 192.540 1.060 192.930 ;
        RECT 1.220 192.540 1.630 192.930 ;
        RECT 0.080 187.100 0.490 187.490 ;
        RECT 0.650 187.100 1.060 187.490 ;
        RECT 1.220 187.100 1.630 187.490 ;
        RECT 49.535 181.560 50.535 182.560 ;
        RECT 50.685 181.560 51.685 182.560 ;
        RECT 51.835 181.560 53.435 182.560 ;
        RECT 53.585 181.560 54.585 182.560 ;
        RECT 54.735 181.560 55.735 182.560 ;
        RECT 69.535 181.560 70.535 182.560 ;
        RECT 70.685 181.560 71.685 182.560 ;
        RECT 71.835 181.560 73.435 182.560 ;
        RECT 73.585 181.560 74.585 182.560 ;
        RECT 74.735 181.560 75.735 182.560 ;
        RECT 89.535 181.560 90.535 182.560 ;
        RECT 90.685 181.560 91.685 182.560 ;
        RECT 91.835 181.560 93.435 182.560 ;
        RECT 93.585 181.560 94.585 182.560 ;
        RECT 94.735 181.560 95.735 182.560 ;
        RECT 42.735 175.060 43.435 175.760 ;
        RECT 42.735 174.210 43.435 174.910 ;
        RECT 42.735 173.360 43.435 174.060 ;
        RECT 61.835 175.060 62.535 175.760 ;
        RECT 62.735 175.060 63.435 175.760 ;
        RECT 61.835 174.210 62.535 174.910 ;
        RECT 62.735 174.210 63.435 174.910 ;
        RECT 61.835 173.360 62.535 174.060 ;
        RECT 62.735 173.360 63.435 174.060 ;
        RECT 42.735 171.260 43.435 171.960 ;
        RECT 42.735 170.410 43.435 171.110 ;
        RECT 42.735 169.560 43.435 170.260 ;
        RECT 81.835 175.060 82.535 175.760 ;
        RECT 82.735 175.060 83.435 175.760 ;
        RECT 81.835 174.210 82.535 174.910 ;
        RECT 82.735 174.210 83.435 174.910 ;
        RECT 81.835 173.360 82.535 174.060 ;
        RECT 82.735 173.360 83.435 174.060 ;
        RECT 61.835 171.260 62.535 171.960 ;
        RECT 62.735 171.260 63.435 171.960 ;
        RECT 61.835 170.410 62.535 171.110 ;
        RECT 62.735 170.410 63.435 171.110 ;
        RECT 61.835 169.560 62.535 170.260 ;
        RECT 62.735 169.560 63.435 170.260 ;
        RECT 101.835 175.060 102.535 175.760 ;
        RECT 101.835 174.210 102.535 174.910 ;
        RECT 101.835 173.360 102.535 174.060 ;
        RECT 81.835 171.260 82.535 171.960 ;
        RECT 82.735 171.260 83.435 171.960 ;
        RECT 81.835 170.410 82.535 171.110 ;
        RECT 82.735 170.410 83.435 171.110 ;
        RECT 81.835 169.560 82.535 170.260 ;
        RECT 82.735 169.560 83.435 170.260 ;
        RECT 102.800 172.980 103.200 173.380 ;
        RECT 103.425 172.980 103.825 173.380 ;
        RECT 104.050 172.980 104.450 173.380 ;
        RECT 107.675 172.980 108.075 173.380 ;
        RECT 108.300 172.980 108.700 173.380 ;
        RECT 108.925 172.980 109.325 173.380 ;
        RECT 102.795 172.380 103.195 172.780 ;
        RECT 103.420 172.380 103.820 172.780 ;
        RECT 104.045 172.380 104.445 172.780 ;
        RECT 107.670 172.380 108.070 172.780 ;
        RECT 108.295 172.380 108.695 172.780 ;
        RECT 108.920 172.380 109.320 172.780 ;
        RECT 101.835 171.260 102.535 171.960 ;
        RECT 101.835 170.410 102.535 171.110 ;
        RECT 101.835 169.560 102.535 170.260 ;
        RECT 49.535 162.760 50.535 163.760 ;
        RECT 50.635 162.760 51.635 163.760 ;
        RECT 51.785 162.760 53.385 163.760 ;
        RECT 53.585 162.760 54.585 163.760 ;
        RECT 54.735 162.760 55.735 163.760 ;
        RECT 69.535 162.760 70.535 163.760 ;
        RECT 70.635 162.760 71.635 163.760 ;
        RECT 71.785 162.760 73.385 163.760 ;
        RECT 73.585 162.760 74.585 163.760 ;
        RECT 74.735 162.760 75.735 163.760 ;
        RECT 89.535 162.760 90.535 163.760 ;
        RECT 90.635 162.760 91.635 163.760 ;
        RECT 91.785 162.760 93.385 163.760 ;
        RECT 93.585 162.760 94.585 163.760 ;
        RECT 94.735 162.760 95.735 163.760 ;
      LAYER met2 ;
        RECT 0.000 197.640 2.000 198.760 ;
        RECT 107.510 197.485 109.510 198.760 ;
        RECT 0.000 192.495 1.710 192.975 ;
        RECT 0.000 187.055 1.710 187.535 ;
        RECT 49.435 181.760 55.835 182.660 ;
        RECT 69.435 181.760 75.835 182.660 ;
        RECT 89.435 181.760 95.835 182.660 ;
        RECT 47.535 181.260 57.735 181.760 ;
        RECT 67.535 181.260 77.735 181.760 ;
        RECT 87.535 181.260 97.735 181.760 ;
        RECT 44.435 181.210 60.835 181.260 ;
        RECT 44.435 180.660 48.235 181.210 ;
        RECT 47.935 180.210 48.235 180.660 ;
        RECT 44.385 180.060 48.235 180.210 ;
        RECT 47.935 179.610 48.235 180.060 ;
        RECT 44.385 179.460 48.235 179.610 ;
        RECT 47.935 179.010 48.235 179.460 ;
        RECT 44.385 178.860 48.235 179.010 ;
        RECT 47.935 178.410 48.235 178.860 ;
        RECT 44.385 178.260 48.235 178.410 ;
        RECT 47.935 177.810 48.235 178.260 ;
        RECT 44.385 177.660 48.235 177.810 ;
        RECT 47.935 177.210 48.235 177.660 ;
        RECT 44.385 177.060 48.235 177.210 ;
        RECT 47.935 176.610 48.235 177.060 ;
        RECT 44.385 176.460 48.235 176.610 ;
        RECT 47.935 176.010 48.235 176.460 ;
        RECT 44.385 175.860 48.235 176.010 ;
        RECT 42.635 169.460 43.535 175.860 ;
        RECT 47.935 175.410 48.235 175.860 ;
        RECT 44.385 175.260 48.235 175.410 ;
        RECT 47.935 174.810 48.235 175.260 ;
        RECT 44.385 174.660 48.235 174.810 ;
        RECT 47.935 174.210 48.235 174.660 ;
        RECT 44.385 174.060 48.235 174.210 ;
        RECT 47.935 173.610 48.235 174.060 ;
        RECT 44.385 173.460 48.235 173.610 ;
        RECT 47.935 173.010 48.235 173.460 ;
        RECT 48.685 173.010 48.835 181.210 ;
        RECT 49.285 173.010 49.435 181.210 ;
        RECT 49.885 173.010 50.035 181.210 ;
        RECT 50.485 173.010 50.635 181.210 ;
        RECT 51.085 173.010 51.235 181.210 ;
        RECT 51.685 173.010 51.835 181.210 ;
        RECT 47.935 171.860 48.235 172.310 ;
        RECT 44.385 171.710 48.235 171.860 ;
        RECT 47.935 171.260 48.235 171.710 ;
        RECT 44.385 171.110 48.235 171.260 ;
        RECT 47.935 170.660 48.235 171.110 ;
        RECT 44.385 170.510 48.235 170.660 ;
        RECT 47.935 170.060 48.235 170.510 ;
        RECT 44.385 169.910 48.235 170.060 ;
        RECT 47.935 169.460 48.235 169.910 ;
        RECT 44.385 169.310 48.235 169.460 ;
        RECT 47.935 168.860 48.235 169.310 ;
        RECT 44.385 168.710 48.235 168.860 ;
        RECT 47.935 168.260 48.235 168.710 ;
        RECT 44.385 168.110 48.235 168.260 ;
        RECT 47.935 167.660 48.235 168.110 ;
        RECT 44.385 167.510 48.235 167.660 ;
        RECT 47.935 167.060 48.235 167.510 ;
        RECT 44.385 166.910 48.235 167.060 ;
        RECT 47.935 166.460 48.235 166.910 ;
        RECT 44.385 166.310 48.235 166.460 ;
        RECT 47.935 165.860 48.235 166.310 ;
        RECT 44.385 165.710 48.235 165.860 ;
        RECT 47.935 165.260 48.235 165.710 ;
        RECT 44.385 165.110 48.235 165.260 ;
        RECT 47.935 164.660 48.235 165.110 ;
        RECT 44.435 164.110 48.235 164.660 ;
        RECT 48.685 164.110 48.835 172.310 ;
        RECT 49.285 164.110 49.435 172.310 ;
        RECT 49.885 164.110 50.035 172.310 ;
        RECT 50.485 164.110 50.635 172.310 ;
        RECT 51.085 164.110 51.235 172.310 ;
        RECT 51.685 164.110 51.835 172.310 ;
        RECT 52.285 164.110 52.985 181.210 ;
        RECT 53.435 173.010 53.585 181.210 ;
        RECT 54.035 173.010 54.185 181.210 ;
        RECT 54.635 173.010 54.785 181.210 ;
        RECT 55.235 173.010 55.385 181.210 ;
        RECT 55.835 173.010 55.985 181.210 ;
        RECT 56.435 173.010 56.585 181.210 ;
        RECT 57.035 180.660 60.835 181.210 ;
        RECT 64.435 181.210 80.835 181.260 ;
        RECT 64.435 180.660 68.235 181.210 ;
        RECT 57.035 180.210 57.335 180.660 ;
        RECT 67.935 180.210 68.235 180.660 ;
        RECT 57.035 180.060 60.885 180.210 ;
        RECT 64.385 180.060 68.235 180.210 ;
        RECT 57.035 179.610 57.335 180.060 ;
        RECT 67.935 179.610 68.235 180.060 ;
        RECT 57.035 179.460 60.885 179.610 ;
        RECT 64.385 179.460 68.235 179.610 ;
        RECT 57.035 179.010 57.335 179.460 ;
        RECT 67.935 179.010 68.235 179.460 ;
        RECT 57.035 178.860 60.885 179.010 ;
        RECT 64.385 178.860 68.235 179.010 ;
        RECT 57.035 178.410 57.335 178.860 ;
        RECT 67.935 178.410 68.235 178.860 ;
        RECT 57.035 178.260 60.885 178.410 ;
        RECT 64.385 178.260 68.235 178.410 ;
        RECT 57.035 177.810 57.335 178.260 ;
        RECT 67.935 177.810 68.235 178.260 ;
        RECT 57.035 177.660 60.885 177.810 ;
        RECT 64.385 177.660 68.235 177.810 ;
        RECT 57.035 177.210 57.335 177.660 ;
        RECT 67.935 177.210 68.235 177.660 ;
        RECT 57.035 177.060 60.885 177.210 ;
        RECT 64.385 177.060 68.235 177.210 ;
        RECT 57.035 176.610 57.335 177.060 ;
        RECT 67.935 176.610 68.235 177.060 ;
        RECT 57.035 176.460 60.885 176.610 ;
        RECT 64.385 176.460 68.235 176.610 ;
        RECT 57.035 176.010 57.335 176.460 ;
        RECT 67.935 176.010 68.235 176.460 ;
        RECT 57.035 175.860 60.885 176.010 ;
        RECT 64.385 175.860 68.235 176.010 ;
        RECT 57.035 175.410 57.335 175.860 ;
        RECT 57.035 175.260 60.885 175.410 ;
        RECT 57.035 174.810 57.335 175.260 ;
        RECT 57.035 174.660 60.885 174.810 ;
        RECT 57.035 174.210 57.335 174.660 ;
        RECT 57.035 174.060 60.885 174.210 ;
        RECT 57.035 173.610 57.335 174.060 ;
        RECT 57.035 173.460 60.885 173.610 ;
        RECT 57.035 173.010 57.335 173.460 ;
        RECT 53.435 164.110 53.585 172.310 ;
        RECT 54.035 164.110 54.185 172.310 ;
        RECT 54.635 164.110 54.785 172.310 ;
        RECT 55.235 164.110 55.385 172.310 ;
        RECT 55.835 164.110 55.985 172.310 ;
        RECT 56.435 164.110 56.585 172.310 ;
        RECT 57.035 171.860 57.335 172.310 ;
        RECT 57.035 171.710 60.885 171.860 ;
        RECT 57.035 171.260 57.335 171.710 ;
        RECT 57.035 171.110 60.885 171.260 ;
        RECT 57.035 170.660 57.335 171.110 ;
        RECT 57.035 170.510 60.885 170.660 ;
        RECT 57.035 170.060 57.335 170.510 ;
        RECT 57.035 169.910 60.885 170.060 ;
        RECT 57.035 169.460 57.335 169.910 ;
        RECT 61.735 169.460 63.535 175.860 ;
        RECT 67.935 175.410 68.235 175.860 ;
        RECT 64.385 175.260 68.235 175.410 ;
        RECT 67.935 174.810 68.235 175.260 ;
        RECT 64.385 174.660 68.235 174.810 ;
        RECT 67.935 174.210 68.235 174.660 ;
        RECT 64.385 174.060 68.235 174.210 ;
        RECT 67.935 173.610 68.235 174.060 ;
        RECT 64.385 173.460 68.235 173.610 ;
        RECT 67.935 173.010 68.235 173.460 ;
        RECT 68.685 173.010 68.835 181.210 ;
        RECT 69.285 173.010 69.435 181.210 ;
        RECT 69.885 173.010 70.035 181.210 ;
        RECT 70.485 173.010 70.635 181.210 ;
        RECT 71.085 173.010 71.235 181.210 ;
        RECT 71.685 173.010 71.835 181.210 ;
        RECT 67.935 171.860 68.235 172.310 ;
        RECT 64.385 171.710 68.235 171.860 ;
        RECT 67.935 171.260 68.235 171.710 ;
        RECT 64.385 171.110 68.235 171.260 ;
        RECT 67.935 170.660 68.235 171.110 ;
        RECT 64.385 170.510 68.235 170.660 ;
        RECT 67.935 170.060 68.235 170.510 ;
        RECT 64.385 169.910 68.235 170.060 ;
        RECT 67.935 169.460 68.235 169.910 ;
        RECT 57.035 169.310 60.885 169.460 ;
        RECT 64.385 169.310 68.235 169.460 ;
        RECT 57.035 168.860 57.335 169.310 ;
        RECT 67.935 168.860 68.235 169.310 ;
        RECT 57.035 168.710 60.885 168.860 ;
        RECT 64.385 168.710 68.235 168.860 ;
        RECT 57.035 168.260 57.335 168.710 ;
        RECT 67.935 168.260 68.235 168.710 ;
        RECT 57.035 168.110 60.885 168.260 ;
        RECT 64.385 168.110 68.235 168.260 ;
        RECT 57.035 167.660 57.335 168.110 ;
        RECT 67.935 167.660 68.235 168.110 ;
        RECT 57.035 167.510 60.885 167.660 ;
        RECT 64.385 167.510 68.235 167.660 ;
        RECT 57.035 167.060 57.335 167.510 ;
        RECT 67.935 167.060 68.235 167.510 ;
        RECT 57.035 166.910 60.885 167.060 ;
        RECT 64.385 166.910 68.235 167.060 ;
        RECT 57.035 166.460 57.335 166.910 ;
        RECT 67.935 166.460 68.235 166.910 ;
        RECT 57.035 166.310 60.885 166.460 ;
        RECT 64.385 166.310 68.235 166.460 ;
        RECT 57.035 165.860 57.335 166.310 ;
        RECT 67.935 165.860 68.235 166.310 ;
        RECT 57.035 165.710 60.885 165.860 ;
        RECT 64.385 165.710 68.235 165.860 ;
        RECT 57.035 165.260 57.335 165.710 ;
        RECT 67.935 165.260 68.235 165.710 ;
        RECT 57.035 165.110 60.885 165.260 ;
        RECT 64.385 165.110 68.235 165.260 ;
        RECT 57.035 164.660 57.335 165.110 ;
        RECT 67.935 164.660 68.235 165.110 ;
        RECT 57.035 164.110 60.835 164.660 ;
        RECT 44.435 164.060 60.835 164.110 ;
        RECT 64.435 164.110 68.235 164.660 ;
        RECT 68.685 164.110 68.835 172.310 ;
        RECT 69.285 164.110 69.435 172.310 ;
        RECT 69.885 164.110 70.035 172.310 ;
        RECT 70.485 164.110 70.635 172.310 ;
        RECT 71.085 164.110 71.235 172.310 ;
        RECT 71.685 164.110 71.835 172.310 ;
        RECT 72.285 164.110 72.985 181.210 ;
        RECT 73.435 173.010 73.585 181.210 ;
        RECT 74.035 173.010 74.185 181.210 ;
        RECT 74.635 173.010 74.785 181.210 ;
        RECT 75.235 173.010 75.385 181.210 ;
        RECT 75.835 173.010 75.985 181.210 ;
        RECT 76.435 173.010 76.585 181.210 ;
        RECT 77.035 180.660 80.835 181.210 ;
        RECT 84.435 181.210 100.835 181.260 ;
        RECT 84.435 180.660 88.235 181.210 ;
        RECT 77.035 180.210 77.335 180.660 ;
        RECT 87.935 180.210 88.235 180.660 ;
        RECT 77.035 180.060 80.885 180.210 ;
        RECT 84.385 180.060 88.235 180.210 ;
        RECT 77.035 179.610 77.335 180.060 ;
        RECT 87.935 179.610 88.235 180.060 ;
        RECT 77.035 179.460 80.885 179.610 ;
        RECT 84.385 179.460 88.235 179.610 ;
        RECT 77.035 179.010 77.335 179.460 ;
        RECT 87.935 179.010 88.235 179.460 ;
        RECT 77.035 178.860 80.885 179.010 ;
        RECT 84.385 178.860 88.235 179.010 ;
        RECT 77.035 178.410 77.335 178.860 ;
        RECT 87.935 178.410 88.235 178.860 ;
        RECT 77.035 178.260 80.885 178.410 ;
        RECT 84.385 178.260 88.235 178.410 ;
        RECT 77.035 177.810 77.335 178.260 ;
        RECT 87.935 177.810 88.235 178.260 ;
        RECT 77.035 177.660 80.885 177.810 ;
        RECT 84.385 177.660 88.235 177.810 ;
        RECT 77.035 177.210 77.335 177.660 ;
        RECT 87.935 177.210 88.235 177.660 ;
        RECT 77.035 177.060 80.885 177.210 ;
        RECT 84.385 177.060 88.235 177.210 ;
        RECT 77.035 176.610 77.335 177.060 ;
        RECT 87.935 176.610 88.235 177.060 ;
        RECT 77.035 176.460 80.885 176.610 ;
        RECT 84.385 176.460 88.235 176.610 ;
        RECT 77.035 176.010 77.335 176.460 ;
        RECT 87.935 176.010 88.235 176.460 ;
        RECT 77.035 175.860 80.885 176.010 ;
        RECT 84.385 175.860 88.235 176.010 ;
        RECT 77.035 175.410 77.335 175.860 ;
        RECT 77.035 175.260 80.885 175.410 ;
        RECT 77.035 174.810 77.335 175.260 ;
        RECT 77.035 174.660 80.885 174.810 ;
        RECT 77.035 174.210 77.335 174.660 ;
        RECT 77.035 174.060 80.885 174.210 ;
        RECT 77.035 173.610 77.335 174.060 ;
        RECT 77.035 173.460 80.885 173.610 ;
        RECT 77.035 173.010 77.335 173.460 ;
        RECT 73.435 164.110 73.585 172.310 ;
        RECT 74.035 164.110 74.185 172.310 ;
        RECT 74.635 164.110 74.785 172.310 ;
        RECT 75.235 164.110 75.385 172.310 ;
        RECT 75.835 164.110 75.985 172.310 ;
        RECT 76.435 164.110 76.585 172.310 ;
        RECT 77.035 171.860 77.335 172.310 ;
        RECT 77.035 171.710 80.885 171.860 ;
        RECT 77.035 171.260 77.335 171.710 ;
        RECT 77.035 171.110 80.885 171.260 ;
        RECT 77.035 170.660 77.335 171.110 ;
        RECT 77.035 170.510 80.885 170.660 ;
        RECT 77.035 170.060 77.335 170.510 ;
        RECT 77.035 169.910 80.885 170.060 ;
        RECT 77.035 169.460 77.335 169.910 ;
        RECT 81.735 169.460 83.535 175.860 ;
        RECT 87.935 175.410 88.235 175.860 ;
        RECT 84.385 175.260 88.235 175.410 ;
        RECT 87.935 174.810 88.235 175.260 ;
        RECT 84.385 174.660 88.235 174.810 ;
        RECT 87.935 174.210 88.235 174.660 ;
        RECT 84.385 174.060 88.235 174.210 ;
        RECT 87.935 173.610 88.235 174.060 ;
        RECT 84.385 173.460 88.235 173.610 ;
        RECT 87.935 173.010 88.235 173.460 ;
        RECT 88.685 173.010 88.835 181.210 ;
        RECT 89.285 173.010 89.435 181.210 ;
        RECT 89.885 173.010 90.035 181.210 ;
        RECT 90.485 173.010 90.635 181.210 ;
        RECT 91.085 173.010 91.235 181.210 ;
        RECT 91.685 173.010 91.835 181.210 ;
        RECT 87.935 171.860 88.235 172.310 ;
        RECT 84.385 171.710 88.235 171.860 ;
        RECT 87.935 171.260 88.235 171.710 ;
        RECT 84.385 171.110 88.235 171.260 ;
        RECT 87.935 170.660 88.235 171.110 ;
        RECT 84.385 170.510 88.235 170.660 ;
        RECT 87.935 170.060 88.235 170.510 ;
        RECT 84.385 169.910 88.235 170.060 ;
        RECT 87.935 169.460 88.235 169.910 ;
        RECT 77.035 169.310 80.885 169.460 ;
        RECT 84.385 169.310 88.235 169.460 ;
        RECT 77.035 168.860 77.335 169.310 ;
        RECT 87.935 168.860 88.235 169.310 ;
        RECT 77.035 168.710 80.885 168.860 ;
        RECT 84.385 168.710 88.235 168.860 ;
        RECT 77.035 168.260 77.335 168.710 ;
        RECT 87.935 168.260 88.235 168.710 ;
        RECT 77.035 168.110 80.885 168.260 ;
        RECT 84.385 168.110 88.235 168.260 ;
        RECT 77.035 167.660 77.335 168.110 ;
        RECT 87.935 167.660 88.235 168.110 ;
        RECT 77.035 167.510 80.885 167.660 ;
        RECT 84.385 167.510 88.235 167.660 ;
        RECT 77.035 167.060 77.335 167.510 ;
        RECT 87.935 167.060 88.235 167.510 ;
        RECT 77.035 166.910 80.885 167.060 ;
        RECT 84.385 166.910 88.235 167.060 ;
        RECT 77.035 166.460 77.335 166.910 ;
        RECT 87.935 166.460 88.235 166.910 ;
        RECT 77.035 166.310 80.885 166.460 ;
        RECT 84.385 166.310 88.235 166.460 ;
        RECT 77.035 165.860 77.335 166.310 ;
        RECT 87.935 165.860 88.235 166.310 ;
        RECT 77.035 165.710 80.885 165.860 ;
        RECT 84.385 165.710 88.235 165.860 ;
        RECT 77.035 165.260 77.335 165.710 ;
        RECT 87.935 165.260 88.235 165.710 ;
        RECT 77.035 165.110 80.885 165.260 ;
        RECT 84.385 165.110 88.235 165.260 ;
        RECT 77.035 164.660 77.335 165.110 ;
        RECT 87.935 164.660 88.235 165.110 ;
        RECT 77.035 164.110 80.835 164.660 ;
        RECT 64.435 164.060 80.835 164.110 ;
        RECT 84.435 164.110 88.235 164.660 ;
        RECT 88.685 164.110 88.835 172.310 ;
        RECT 89.285 164.110 89.435 172.310 ;
        RECT 89.885 164.110 90.035 172.310 ;
        RECT 90.485 164.110 90.635 172.310 ;
        RECT 91.085 164.110 91.235 172.310 ;
        RECT 91.685 164.110 91.835 172.310 ;
        RECT 92.285 164.110 92.985 181.210 ;
        RECT 93.435 173.010 93.585 181.210 ;
        RECT 94.035 173.010 94.185 181.210 ;
        RECT 94.635 173.010 94.785 181.210 ;
        RECT 95.235 173.010 95.385 181.210 ;
        RECT 95.835 173.010 95.985 181.210 ;
        RECT 96.435 173.010 96.585 181.210 ;
        RECT 97.035 180.660 100.835 181.210 ;
        RECT 97.035 180.210 97.335 180.660 ;
        RECT 97.035 180.060 100.885 180.210 ;
        RECT 97.035 179.610 97.335 180.060 ;
        RECT 97.035 179.460 100.885 179.610 ;
        RECT 97.035 179.010 97.335 179.460 ;
        RECT 97.035 178.860 100.885 179.010 ;
        RECT 97.035 178.410 97.335 178.860 ;
        RECT 97.035 178.260 100.885 178.410 ;
        RECT 97.035 177.810 97.335 178.260 ;
        RECT 97.035 177.660 100.885 177.810 ;
        RECT 97.035 177.210 97.335 177.660 ;
        RECT 97.035 177.060 100.885 177.210 ;
        RECT 97.035 176.610 97.335 177.060 ;
        RECT 97.035 176.460 100.885 176.610 ;
        RECT 97.035 176.010 97.335 176.460 ;
        RECT 97.035 175.860 100.885 176.010 ;
        RECT 97.035 175.410 97.335 175.860 ;
        RECT 97.035 175.260 100.885 175.410 ;
        RECT 97.035 174.810 97.335 175.260 ;
        RECT 97.035 174.660 100.885 174.810 ;
        RECT 97.035 174.210 97.335 174.660 ;
        RECT 97.035 174.060 100.885 174.210 ;
        RECT 97.035 173.610 97.335 174.060 ;
        RECT 97.035 173.460 100.885 173.610 ;
        RECT 101.735 173.510 102.635 175.860 ;
        RECT 97.035 173.010 97.335 173.460 ;
        RECT 93.435 164.110 93.585 172.310 ;
        RECT 94.035 164.110 94.185 172.310 ;
        RECT 94.635 164.110 94.785 172.310 ;
        RECT 95.235 164.110 95.385 172.310 ;
        RECT 95.835 164.110 95.985 172.310 ;
        RECT 96.435 164.110 96.585 172.310 ;
        RECT 97.035 171.860 97.335 172.310 ;
        RECT 101.735 172.235 104.635 173.510 ;
        RECT 107.510 172.235 109.510 173.510 ;
        RECT 97.035 171.710 100.885 171.860 ;
        RECT 97.035 171.260 97.335 171.710 ;
        RECT 97.035 171.110 100.885 171.260 ;
        RECT 97.035 170.660 97.335 171.110 ;
        RECT 97.035 170.510 100.885 170.660 ;
        RECT 97.035 170.060 97.335 170.510 ;
        RECT 97.035 169.910 100.885 170.060 ;
        RECT 97.035 169.460 97.335 169.910 ;
        RECT 101.735 169.460 102.635 172.235 ;
        RECT 97.035 169.310 100.885 169.460 ;
        RECT 97.035 168.860 97.335 169.310 ;
        RECT 97.035 168.710 100.885 168.860 ;
        RECT 97.035 168.260 97.335 168.710 ;
        RECT 97.035 168.110 100.885 168.260 ;
        RECT 97.035 167.660 97.335 168.110 ;
        RECT 97.035 167.510 100.885 167.660 ;
        RECT 97.035 167.060 97.335 167.510 ;
        RECT 97.035 166.910 100.885 167.060 ;
        RECT 97.035 166.460 97.335 166.910 ;
        RECT 97.035 166.310 100.885 166.460 ;
        RECT 97.035 165.860 97.335 166.310 ;
        RECT 97.035 165.710 100.885 165.860 ;
        RECT 97.035 165.260 97.335 165.710 ;
        RECT 97.035 165.110 100.885 165.260 ;
        RECT 97.035 164.660 97.335 165.110 ;
        RECT 97.035 164.110 100.835 164.660 ;
        RECT 84.435 164.060 100.835 164.110 ;
        RECT 47.535 163.560 57.735 164.060 ;
        RECT 67.535 163.560 77.735 164.060 ;
        RECT 87.535 163.560 97.735 164.060 ;
        RECT 49.435 162.660 55.835 163.560 ;
        RECT 69.435 162.660 75.835 163.560 ;
        RECT 89.435 162.660 95.835 163.560 ;
      LAYER via2 ;
        RECT 0.160 198.305 0.560 198.705 ;
        RECT 0.785 198.305 1.185 198.705 ;
        RECT 1.410 198.305 1.810 198.705 ;
        RECT 0.160 197.775 0.560 198.175 ;
        RECT 0.785 197.775 1.185 198.175 ;
        RECT 1.410 197.775 1.810 198.175 ;
        RECT 107.675 198.230 108.075 198.630 ;
        RECT 108.300 198.230 108.700 198.630 ;
        RECT 108.925 198.230 109.325 198.630 ;
        RECT 107.670 197.630 108.070 198.030 ;
        RECT 108.295 197.630 108.695 198.030 ;
        RECT 108.920 197.630 109.320 198.030 ;
        RECT 0.080 192.540 0.490 192.930 ;
        RECT 0.650 192.540 1.060 192.930 ;
        RECT 1.220 192.540 1.630 192.930 ;
        RECT 0.080 187.100 0.490 187.490 ;
        RECT 0.650 187.100 1.060 187.490 ;
        RECT 1.220 187.100 1.630 187.490 ;
        RECT 102.800 172.980 103.200 173.380 ;
        RECT 103.425 172.980 103.825 173.380 ;
        RECT 104.050 172.980 104.450 173.380 ;
        RECT 102.795 172.380 103.195 172.780 ;
        RECT 103.420 172.380 103.820 172.780 ;
        RECT 104.045 172.380 104.445 172.780 ;
        RECT 107.675 172.980 108.075 173.380 ;
        RECT 108.300 172.980 108.700 173.380 ;
        RECT 108.925 172.980 109.325 173.380 ;
        RECT 107.670 172.380 108.070 172.780 ;
        RECT 108.295 172.380 108.695 172.780 ;
        RECT 108.920 172.380 109.320 172.780 ;
      LAYER met3 ;
        RECT 0.000 197.640 2.000 198.760 ;
        RECT 107.510 197.485 109.510 198.760 ;
        RECT 0.000 192.495 1.710 192.975 ;
        RECT 0.000 187.055 1.710 187.535 ;
        RECT 49.435 181.810 55.835 182.660 ;
        RECT 69.435 181.810 75.835 182.660 ;
        RECT 89.435 181.810 95.835 182.660 ;
        RECT 42.635 169.460 43.485 175.860 ;
        RECT 61.785 169.460 63.485 175.860 ;
        RECT 81.785 169.460 83.485 175.860 ;
        RECT 101.785 173.510 102.635 175.860 ;
        RECT 101.785 172.235 104.635 173.510 ;
        RECT 107.510 172.235 109.510 173.510 ;
        RECT 101.785 169.460 102.635 172.235 ;
        RECT 49.435 162.660 55.835 163.510 ;
        RECT 69.435 162.660 75.835 163.510 ;
        RECT 89.435 162.660 95.835 163.510 ;
      LAYER via3 ;
        RECT 0.160 198.305 0.555 198.705 ;
        RECT 0.780 198.305 1.180 198.705 ;
        RECT 1.410 198.305 1.810 198.705 ;
        RECT 0.160 197.775 0.555 198.175 ;
        RECT 0.780 197.775 1.180 198.175 ;
        RECT 1.410 197.775 1.810 198.175 ;
        RECT 107.675 198.230 108.075 198.630 ;
        RECT 108.300 198.230 108.700 198.630 ;
        RECT 108.925 198.230 109.325 198.630 ;
        RECT 107.670 197.630 108.070 198.030 ;
        RECT 108.295 197.630 108.695 198.030 ;
        RECT 108.920 197.630 109.320 198.030 ;
        RECT 0.075 192.535 0.495 192.935 ;
        RECT 0.645 192.535 1.065 192.935 ;
        RECT 1.215 192.535 1.635 192.935 ;
        RECT 0.075 187.095 0.495 187.495 ;
        RECT 0.645 187.095 1.065 187.495 ;
        RECT 1.215 187.095 1.635 187.495 ;
        RECT 49.535 181.910 50.185 182.560 ;
        RECT 50.335 181.910 50.985 182.560 ;
        RECT 51.135 181.910 51.785 182.560 ;
        RECT 53.485 181.910 54.135 182.560 ;
        RECT 54.285 181.910 54.935 182.560 ;
        RECT 55.085 181.910 55.735 182.560 ;
        RECT 69.535 181.910 70.185 182.560 ;
        RECT 70.335 181.910 70.985 182.560 ;
        RECT 71.135 181.910 71.785 182.560 ;
        RECT 73.485 181.910 74.135 182.560 ;
        RECT 74.285 181.910 74.935 182.560 ;
        RECT 75.085 181.910 75.735 182.560 ;
        RECT 89.535 181.910 90.185 182.560 ;
        RECT 90.335 181.910 90.985 182.560 ;
        RECT 91.135 181.910 91.785 182.560 ;
        RECT 93.485 181.910 94.135 182.560 ;
        RECT 94.285 181.910 94.935 182.560 ;
        RECT 95.085 181.910 95.735 182.560 ;
        RECT 42.735 175.110 43.385 175.760 ;
        RECT 42.735 174.310 43.385 174.960 ;
        RECT 42.735 173.510 43.385 174.160 ;
        RECT 42.735 171.160 43.385 171.810 ;
        RECT 42.735 170.360 43.385 171.010 ;
        RECT 42.735 169.560 43.385 170.210 ;
        RECT 61.885 175.110 62.535 175.760 ;
        RECT 62.735 175.110 63.385 175.760 ;
        RECT 61.885 174.310 62.535 174.960 ;
        RECT 62.735 174.310 63.385 174.960 ;
        RECT 61.885 173.510 62.535 174.160 ;
        RECT 62.735 173.510 63.385 174.160 ;
        RECT 61.885 171.160 62.535 171.810 ;
        RECT 62.735 171.160 63.385 171.810 ;
        RECT 61.885 170.360 62.535 171.010 ;
        RECT 62.735 170.360 63.385 171.010 ;
        RECT 61.885 169.560 62.535 170.210 ;
        RECT 62.735 169.560 63.385 170.210 ;
        RECT 81.885 175.110 82.535 175.760 ;
        RECT 82.735 175.110 83.385 175.760 ;
        RECT 81.885 174.310 82.535 174.960 ;
        RECT 82.735 174.310 83.385 174.960 ;
        RECT 81.885 173.510 82.535 174.160 ;
        RECT 82.735 173.510 83.385 174.160 ;
        RECT 81.885 171.160 82.535 171.810 ;
        RECT 82.735 171.160 83.385 171.810 ;
        RECT 81.885 170.360 82.535 171.010 ;
        RECT 82.735 170.360 83.385 171.010 ;
        RECT 81.885 169.560 82.535 170.210 ;
        RECT 82.735 169.560 83.385 170.210 ;
        RECT 101.885 175.110 102.535 175.760 ;
        RECT 101.885 174.310 102.535 174.960 ;
        RECT 101.885 173.510 102.535 174.160 ;
        RECT 102.800 172.980 103.200 173.380 ;
        RECT 103.425 172.980 103.825 173.380 ;
        RECT 104.050 172.980 104.450 173.380 ;
        RECT 102.795 172.380 103.195 172.780 ;
        RECT 103.420 172.380 103.820 172.780 ;
        RECT 104.045 172.380 104.445 172.780 ;
        RECT 107.675 172.980 108.075 173.380 ;
        RECT 108.300 172.980 108.700 173.380 ;
        RECT 108.925 172.980 109.325 173.380 ;
        RECT 107.670 172.380 108.070 172.780 ;
        RECT 108.295 172.380 108.695 172.780 ;
        RECT 108.920 172.380 109.320 172.780 ;
        RECT 101.885 171.160 102.535 171.810 ;
        RECT 101.885 170.360 102.535 171.010 ;
        RECT 101.885 169.560 102.535 170.210 ;
        RECT 49.535 162.760 50.185 163.410 ;
        RECT 50.335 162.760 50.985 163.410 ;
        RECT 51.135 162.760 51.785 163.410 ;
        RECT 53.485 162.760 54.135 163.410 ;
        RECT 54.285 162.760 54.935 163.410 ;
        RECT 55.085 162.760 55.735 163.410 ;
        RECT 69.535 162.760 70.185 163.410 ;
        RECT 70.335 162.760 70.985 163.410 ;
        RECT 71.135 162.760 71.785 163.410 ;
        RECT 73.485 162.760 74.135 163.410 ;
        RECT 74.285 162.760 74.935 163.410 ;
        RECT 75.085 162.760 75.735 163.410 ;
        RECT 89.535 162.760 90.185 163.410 ;
        RECT 90.335 162.760 90.985 163.410 ;
        RECT 91.135 162.760 91.785 163.410 ;
        RECT 93.485 162.760 94.135 163.410 ;
        RECT 94.285 162.760 94.935 163.410 ;
        RECT 95.085 162.760 95.735 163.410 ;
      LAYER met4 ;
        RECT 0.000 0.000 2.000 380.000 ;
        RECT 49.435 181.210 55.835 182.660 ;
        RECT 69.435 181.210 75.835 182.660 ;
        RECT 89.435 181.210 95.835 182.660 ;
        RECT 44.085 175.860 61.185 181.210 ;
        RECT 64.085 175.860 81.185 181.210 ;
        RECT 84.085 175.860 101.185 181.210 ;
        RECT 42.635 173.510 102.635 175.860 ;
        RECT 42.635 172.235 104.635 173.510 ;
        RECT 42.635 169.460 102.635 172.235 ;
        RECT 44.085 164.110 61.185 169.460 ;
        RECT 64.085 164.110 81.185 169.460 ;
        RECT 84.085 164.110 101.185 169.460 ;
        RECT 49.435 162.660 55.835 164.110 ;
        RECT 69.435 162.660 75.835 164.110 ;
        RECT 89.435 162.660 95.835 164.110 ;
        RECT 107.510 0.000 109.510 380.000 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 9.130 379.100 11.530 380.000 ;
        RECT 17.930 379.100 20.330 380.000 ;
        RECT 29.130 379.100 31.530 380.000 ;
        RECT 37.930 379.100 40.330 380.000 ;
        RECT 49.130 379.100 51.530 380.000 ;
        RECT 57.930 379.100 60.330 380.000 ;
        RECT 69.130 379.100 71.530 380.000 ;
        RECT 77.930 379.100 80.330 380.000 ;
        RECT 89.130 379.100 91.530 380.000 ;
        RECT 97.930 379.100 100.330 380.000 ;
        RECT 5.880 378.900 23.830 379.100 ;
        RECT 25.880 378.900 43.830 379.100 ;
        RECT 45.880 378.900 63.830 379.100 ;
        RECT 65.880 378.900 83.830 379.100 ;
        RECT 85.880 378.900 103.830 379.100 ;
        RECT 5.830 378.800 23.830 378.900 ;
        RECT 25.830 378.800 43.830 378.900 ;
        RECT 45.830 378.800 63.830 378.900 ;
        RECT 65.830 378.800 83.830 378.900 ;
        RECT 85.830 378.800 103.830 378.900 ;
        RECT 5.680 375.600 23.830 378.800 ;
        RECT 25.680 375.600 43.830 378.800 ;
        RECT 45.680 375.600 63.830 378.800 ;
        RECT 65.680 375.600 83.830 378.800 ;
        RECT 85.680 375.600 103.830 378.800 ;
        RECT 4.730 373.200 104.730 375.600 ;
        RECT 5.630 366.800 23.830 373.200 ;
        RECT 25.630 366.800 43.830 373.200 ;
        RECT 45.630 366.800 63.830 373.200 ;
        RECT 65.630 366.800 83.830 373.200 ;
        RECT 85.630 366.800 103.830 373.200 ;
        RECT 4.730 364.400 104.730 366.800 ;
        RECT 5.630 360.900 23.830 364.400 ;
        RECT 25.630 360.900 43.830 364.400 ;
        RECT 45.630 360.900 63.830 364.400 ;
        RECT 65.630 360.900 83.830 364.400 ;
        RECT 85.630 360.900 103.830 364.400 ;
        RECT 9.130 359.100 11.530 360.900 ;
        RECT 17.930 359.100 20.330 360.900 ;
        RECT 29.130 359.100 31.530 360.900 ;
        RECT 37.930 359.100 40.330 360.900 ;
        RECT 49.130 359.100 51.530 360.900 ;
        RECT 57.930 359.100 60.330 360.900 ;
        RECT 69.130 359.100 71.530 360.900 ;
        RECT 77.930 359.100 80.330 360.900 ;
        RECT 89.130 359.100 91.530 360.900 ;
        RECT 97.930 359.100 100.330 360.900 ;
        RECT 5.880 358.900 23.830 359.100 ;
        RECT 25.880 358.900 43.830 359.100 ;
        RECT 45.880 358.900 63.830 359.100 ;
        RECT 65.880 358.900 83.830 359.100 ;
        RECT 85.880 358.900 103.830 359.100 ;
        RECT 5.830 358.800 23.830 358.900 ;
        RECT 25.830 358.800 43.830 358.900 ;
        RECT 45.830 358.800 63.830 358.900 ;
        RECT 65.830 358.800 83.830 358.900 ;
        RECT 85.830 358.800 103.830 358.900 ;
        RECT 5.680 355.600 23.830 358.800 ;
        RECT 25.680 355.600 43.830 358.800 ;
        RECT 45.680 355.600 63.830 358.800 ;
        RECT 65.680 355.600 83.830 358.800 ;
        RECT 85.680 355.600 103.830 358.800 ;
        RECT 4.730 353.200 104.730 355.600 ;
        RECT 5.630 346.800 23.830 353.200 ;
        RECT 25.630 346.800 43.830 353.200 ;
        RECT 45.630 346.800 63.830 353.200 ;
        RECT 65.630 346.800 83.830 353.200 ;
        RECT 85.630 346.800 103.830 353.200 ;
        RECT 4.730 344.400 104.730 346.800 ;
        RECT 5.630 340.900 23.830 344.400 ;
        RECT 25.630 340.900 43.830 344.400 ;
        RECT 45.630 340.900 63.830 344.400 ;
        RECT 65.630 340.900 83.830 344.400 ;
        RECT 85.630 340.900 103.830 344.400 ;
        RECT 9.130 339.100 11.530 340.900 ;
        RECT 17.930 339.100 20.330 340.900 ;
        RECT 29.130 339.100 31.530 340.900 ;
        RECT 37.930 339.100 40.330 340.900 ;
        RECT 49.130 339.100 51.530 340.900 ;
        RECT 57.930 339.100 60.330 340.900 ;
        RECT 69.130 339.100 71.530 340.900 ;
        RECT 77.930 339.100 80.330 340.900 ;
        RECT 89.130 339.100 91.530 340.900 ;
        RECT 97.930 339.100 100.330 340.900 ;
        RECT 5.880 338.900 23.830 339.100 ;
        RECT 25.880 338.900 43.830 339.100 ;
        RECT 45.880 338.900 63.830 339.100 ;
        RECT 65.880 338.900 83.830 339.100 ;
        RECT 85.880 338.900 103.830 339.100 ;
        RECT 5.830 338.800 23.830 338.900 ;
        RECT 25.830 338.800 43.830 338.900 ;
        RECT 45.830 338.800 63.830 338.900 ;
        RECT 65.830 338.800 83.830 338.900 ;
        RECT 85.830 338.800 103.830 338.900 ;
        RECT 5.680 335.600 23.830 338.800 ;
        RECT 25.680 335.600 43.830 338.800 ;
        RECT 45.680 335.600 63.830 338.800 ;
        RECT 65.680 335.600 83.830 338.800 ;
        RECT 85.680 335.600 103.830 338.800 ;
        RECT 4.730 333.200 104.730 335.600 ;
        RECT 5.630 326.800 23.830 333.200 ;
        RECT 25.630 326.800 43.830 333.200 ;
        RECT 45.630 326.800 63.830 333.200 ;
        RECT 65.630 326.800 83.830 333.200 ;
        RECT 85.630 326.800 103.830 333.200 ;
        RECT 4.730 324.400 104.730 326.800 ;
        RECT 5.630 320.900 23.830 324.400 ;
        RECT 25.630 320.900 43.830 324.400 ;
        RECT 45.630 320.900 63.830 324.400 ;
        RECT 65.630 320.900 83.830 324.400 ;
        RECT 85.630 320.900 103.830 324.400 ;
        RECT 9.130 319.100 11.530 320.900 ;
        RECT 17.930 319.100 20.330 320.900 ;
        RECT 29.130 319.100 31.530 320.900 ;
        RECT 37.930 319.100 40.330 320.900 ;
        RECT 49.130 319.100 51.530 320.900 ;
        RECT 57.930 319.100 60.330 320.900 ;
        RECT 69.130 319.100 71.530 320.900 ;
        RECT 77.930 319.100 80.330 320.900 ;
        RECT 89.130 319.100 91.530 320.900 ;
        RECT 97.930 319.100 100.330 320.900 ;
        RECT 5.880 318.900 23.830 319.100 ;
        RECT 25.880 318.900 43.830 319.100 ;
        RECT 45.880 318.900 63.830 319.100 ;
        RECT 65.880 318.900 83.830 319.100 ;
        RECT 85.880 318.900 103.830 319.100 ;
        RECT 5.830 318.800 23.830 318.900 ;
        RECT 25.830 318.800 43.830 318.900 ;
        RECT 45.830 318.800 63.830 318.900 ;
        RECT 65.830 318.800 83.830 318.900 ;
        RECT 85.830 318.800 103.830 318.900 ;
        RECT 5.680 315.600 23.830 318.800 ;
        RECT 25.680 315.600 43.830 318.800 ;
        RECT 45.680 315.600 63.830 318.800 ;
        RECT 65.680 315.600 83.830 318.800 ;
        RECT 85.680 315.600 103.830 318.800 ;
        RECT 4.730 313.200 104.730 315.600 ;
        RECT 5.630 306.800 23.830 313.200 ;
        RECT 25.630 306.800 43.830 313.200 ;
        RECT 45.630 306.800 63.830 313.200 ;
        RECT 65.630 306.800 83.830 313.200 ;
        RECT 85.630 306.800 103.830 313.200 ;
        RECT 4.730 304.400 104.730 306.800 ;
        RECT 5.630 300.900 23.830 304.400 ;
        RECT 25.630 300.900 43.830 304.400 ;
        RECT 45.630 300.900 63.830 304.400 ;
        RECT 65.630 300.900 83.830 304.400 ;
        RECT 85.630 300.900 103.830 304.400 ;
        RECT 9.130 299.100 11.530 300.900 ;
        RECT 17.930 299.100 20.330 300.900 ;
        RECT 29.130 299.100 31.530 300.900 ;
        RECT 37.930 299.100 40.330 300.900 ;
        RECT 49.130 299.100 51.530 300.900 ;
        RECT 57.930 299.100 60.330 300.900 ;
        RECT 69.130 299.100 71.530 300.900 ;
        RECT 77.930 299.100 80.330 300.900 ;
        RECT 89.130 299.100 91.530 300.900 ;
        RECT 97.930 299.100 100.330 300.900 ;
        RECT 5.880 298.900 23.830 299.100 ;
        RECT 25.880 298.900 43.830 299.100 ;
        RECT 45.880 298.900 63.830 299.100 ;
        RECT 65.880 298.900 83.830 299.100 ;
        RECT 85.880 298.900 103.830 299.100 ;
        RECT 5.830 298.800 23.830 298.900 ;
        RECT 25.830 298.800 43.830 298.900 ;
        RECT 45.830 298.800 63.830 298.900 ;
        RECT 65.830 298.800 83.830 298.900 ;
        RECT 85.830 298.800 103.830 298.900 ;
        RECT 5.680 295.600 23.830 298.800 ;
        RECT 25.680 295.600 43.830 298.800 ;
        RECT 45.680 295.600 63.830 298.800 ;
        RECT 65.680 295.600 83.830 298.800 ;
        RECT 85.680 295.600 103.830 298.800 ;
        RECT 4.730 293.200 104.730 295.600 ;
        RECT 5.630 286.800 23.830 293.200 ;
        RECT 25.630 286.800 43.830 293.200 ;
        RECT 45.630 286.800 63.830 293.200 ;
        RECT 65.630 286.800 83.830 293.200 ;
        RECT 85.630 286.800 103.830 293.200 ;
        RECT 4.730 284.400 104.730 286.800 ;
        RECT 5.630 280.900 23.830 284.400 ;
        RECT 25.630 280.900 43.830 284.400 ;
        RECT 45.630 280.900 63.830 284.400 ;
        RECT 65.630 280.900 83.830 284.400 ;
        RECT 85.630 280.900 103.830 284.400 ;
        RECT 9.130 279.100 11.530 280.900 ;
        RECT 17.930 279.100 20.330 280.900 ;
        RECT 29.130 279.100 31.530 280.900 ;
        RECT 37.930 279.100 40.330 280.900 ;
        RECT 49.130 279.100 51.530 280.900 ;
        RECT 57.930 279.100 60.330 280.900 ;
        RECT 69.130 279.100 71.530 280.900 ;
        RECT 77.930 279.100 80.330 280.900 ;
        RECT 89.130 279.100 91.530 280.900 ;
        RECT 97.930 279.100 100.330 280.900 ;
        RECT 5.880 278.900 23.830 279.100 ;
        RECT 25.880 278.900 43.830 279.100 ;
        RECT 45.880 278.900 63.830 279.100 ;
        RECT 65.880 278.900 83.830 279.100 ;
        RECT 85.880 278.900 103.830 279.100 ;
        RECT 5.830 278.800 23.830 278.900 ;
        RECT 25.830 278.800 43.830 278.900 ;
        RECT 45.830 278.800 63.830 278.900 ;
        RECT 65.830 278.800 83.830 278.900 ;
        RECT 85.830 278.800 103.830 278.900 ;
        RECT 5.680 275.600 23.830 278.800 ;
        RECT 25.680 275.600 43.830 278.800 ;
        RECT 45.680 275.600 63.830 278.800 ;
        RECT 65.680 275.600 83.830 278.800 ;
        RECT 85.680 275.600 103.830 278.800 ;
        RECT 4.730 273.200 104.730 275.600 ;
        RECT 5.630 266.800 23.830 273.200 ;
        RECT 25.630 266.800 43.830 273.200 ;
        RECT 45.630 266.800 63.830 273.200 ;
        RECT 65.630 266.800 83.830 273.200 ;
        RECT 85.630 266.800 103.830 273.200 ;
        RECT 4.730 264.400 104.730 266.800 ;
        RECT 5.630 260.900 23.830 264.400 ;
        RECT 25.630 260.900 43.830 264.400 ;
        RECT 45.630 260.900 63.830 264.400 ;
        RECT 65.630 260.900 83.830 264.400 ;
        RECT 85.630 260.900 103.830 264.400 ;
        RECT 9.130 259.100 11.530 260.900 ;
        RECT 17.930 259.100 20.330 260.900 ;
        RECT 29.130 259.100 31.530 260.900 ;
        RECT 37.930 259.100 40.330 260.900 ;
        RECT 49.130 259.100 51.530 260.900 ;
        RECT 57.930 259.100 60.330 260.900 ;
        RECT 69.130 259.100 71.530 260.900 ;
        RECT 77.930 259.100 80.330 260.900 ;
        RECT 89.130 259.100 91.530 260.900 ;
        RECT 97.930 259.100 100.330 260.900 ;
        RECT 5.880 258.900 23.830 259.100 ;
        RECT 25.880 258.900 43.830 259.100 ;
        RECT 45.880 258.900 63.830 259.100 ;
        RECT 65.880 258.900 83.830 259.100 ;
        RECT 85.880 258.900 103.830 259.100 ;
        RECT 5.830 258.800 23.830 258.900 ;
        RECT 25.830 258.800 43.830 258.900 ;
        RECT 45.830 258.800 63.830 258.900 ;
        RECT 65.830 258.800 83.830 258.900 ;
        RECT 85.830 258.800 103.830 258.900 ;
        RECT 5.680 255.600 23.830 258.800 ;
        RECT 25.680 255.600 43.830 258.800 ;
        RECT 45.680 255.600 63.830 258.800 ;
        RECT 65.680 255.600 83.830 258.800 ;
        RECT 85.680 255.600 103.830 258.800 ;
        RECT 4.730 253.200 104.730 255.600 ;
        RECT 5.630 246.800 23.830 253.200 ;
        RECT 25.630 246.800 43.830 253.200 ;
        RECT 45.630 246.800 63.830 253.200 ;
        RECT 65.630 246.800 83.830 253.200 ;
        RECT 85.630 246.800 103.830 253.200 ;
        RECT 4.730 244.400 104.730 246.800 ;
        RECT 5.630 240.900 23.830 244.400 ;
        RECT 25.630 240.900 43.830 244.400 ;
        RECT 45.630 240.900 63.830 244.400 ;
        RECT 65.630 240.900 83.830 244.400 ;
        RECT 85.630 240.900 103.830 244.400 ;
        RECT 9.130 239.100 11.530 240.900 ;
        RECT 17.930 239.100 20.330 240.900 ;
        RECT 29.130 239.100 31.530 240.900 ;
        RECT 37.930 239.100 40.330 240.900 ;
        RECT 49.130 239.100 51.530 240.900 ;
        RECT 57.930 239.100 60.330 240.900 ;
        RECT 69.130 239.100 71.530 240.900 ;
        RECT 77.930 239.100 80.330 240.900 ;
        RECT 89.130 239.100 91.530 240.900 ;
        RECT 97.930 239.100 100.330 240.900 ;
        RECT 5.880 238.900 23.830 239.100 ;
        RECT 25.880 238.900 43.830 239.100 ;
        RECT 45.880 238.900 63.830 239.100 ;
        RECT 65.880 238.900 83.830 239.100 ;
        RECT 85.880 238.900 103.830 239.100 ;
        RECT 5.830 238.800 23.830 238.900 ;
        RECT 25.830 238.800 43.830 238.900 ;
        RECT 45.830 238.800 63.830 238.900 ;
        RECT 65.830 238.800 83.830 238.900 ;
        RECT 85.830 238.800 103.830 238.900 ;
        RECT 5.680 235.600 23.830 238.800 ;
        RECT 25.680 235.600 43.830 238.800 ;
        RECT 45.680 235.600 63.830 238.800 ;
        RECT 65.680 235.600 83.830 238.800 ;
        RECT 85.680 235.600 103.830 238.800 ;
        RECT 4.730 233.200 104.730 235.600 ;
        RECT 5.630 226.800 23.830 233.200 ;
        RECT 25.630 226.800 43.830 233.200 ;
        RECT 45.630 226.800 63.830 233.200 ;
        RECT 65.630 226.800 83.830 233.200 ;
        RECT 85.630 226.800 103.830 233.200 ;
        RECT 4.730 224.400 104.730 226.800 ;
        RECT 5.630 220.900 23.830 224.400 ;
        RECT 25.630 220.900 43.830 224.400 ;
        RECT 45.630 220.900 63.830 224.400 ;
        RECT 65.630 220.900 83.830 224.400 ;
        RECT 85.630 220.900 103.830 224.400 ;
        RECT 9.130 220.000 11.530 220.900 ;
        RECT 17.930 220.000 20.330 220.900 ;
        RECT 29.130 220.000 31.530 220.900 ;
        RECT 37.930 220.000 40.330 220.900 ;
        RECT 49.130 220.000 51.530 220.900 ;
        RECT 57.930 220.000 60.330 220.900 ;
        RECT 69.130 220.000 71.530 220.900 ;
        RECT 77.930 220.000 80.330 220.900 ;
        RECT 89.130 220.000 91.530 220.900 ;
        RECT 97.930 220.000 100.330 220.900 ;
        RECT 6.955 194.485 7.385 195.270 ;
        RECT 14.880 194.480 15.310 195.265 ;
        RECT 7.980 190.205 8.410 190.990 ;
        RECT 23.620 190.205 24.050 190.990 ;
        RECT 6.600 189.040 7.030 189.825 ;
        RECT 23.620 189.040 24.050 189.825 ;
        RECT 7.520 184.765 7.950 185.550 ;
        RECT 14.880 184.765 15.310 185.550 ;
        RECT 47.035 181.760 49.435 182.660 ;
        RECT 55.835 181.760 58.235 182.660 ;
        RECT 67.035 181.760 69.435 182.660 ;
        RECT 75.835 181.760 78.235 182.660 ;
        RECT 87.035 181.760 89.435 182.660 ;
        RECT 95.835 181.760 98.235 182.660 ;
        RECT 43.785 181.560 61.735 181.760 ;
        RECT 63.785 181.560 81.735 181.760 ;
        RECT 83.785 181.560 101.735 181.760 ;
        RECT 43.735 181.460 61.735 181.560 ;
        RECT 63.735 181.460 81.735 181.560 ;
        RECT 83.735 181.460 101.735 181.560 ;
        RECT 43.585 178.260 61.735 181.460 ;
        RECT 63.585 178.260 81.735 181.460 ;
        RECT 83.585 178.260 101.735 181.460 ;
        RECT 42.635 175.860 102.635 178.260 ;
        RECT 43.535 169.460 61.735 175.860 ;
        RECT 63.535 169.460 81.735 175.860 ;
        RECT 83.535 169.460 101.735 175.860 ;
        RECT 42.635 167.060 102.635 169.460 ;
        RECT 43.535 163.560 61.735 167.060 ;
        RECT 63.535 163.560 81.735 167.060 ;
        RECT 83.535 163.560 101.735 167.060 ;
        RECT 47.035 162.660 49.435 163.560 ;
        RECT 55.835 162.660 58.235 163.560 ;
        RECT 67.035 162.660 69.435 163.560 ;
        RECT 75.835 162.660 78.235 163.560 ;
        RECT 87.035 162.660 89.435 163.560 ;
        RECT 95.835 162.660 98.235 163.560 ;
        RECT 9.130 159.100 11.530 160.000 ;
        RECT 17.930 159.100 20.330 160.000 ;
        RECT 29.130 159.100 31.530 160.000 ;
        RECT 37.930 159.100 40.330 160.000 ;
        RECT 49.130 159.100 51.530 160.000 ;
        RECT 57.930 159.100 60.330 160.000 ;
        RECT 69.130 159.100 71.530 160.000 ;
        RECT 77.930 159.100 80.330 160.000 ;
        RECT 89.130 159.100 91.530 160.000 ;
        RECT 97.930 159.100 100.330 160.000 ;
        RECT 5.880 158.900 23.830 159.100 ;
        RECT 25.880 158.900 43.830 159.100 ;
        RECT 45.880 158.900 63.830 159.100 ;
        RECT 65.880 158.900 83.830 159.100 ;
        RECT 85.880 158.900 103.830 159.100 ;
        RECT 5.830 158.800 23.830 158.900 ;
        RECT 25.830 158.800 43.830 158.900 ;
        RECT 45.830 158.800 63.830 158.900 ;
        RECT 65.830 158.800 83.830 158.900 ;
        RECT 85.830 158.800 103.830 158.900 ;
        RECT 5.680 155.600 23.830 158.800 ;
        RECT 25.680 155.600 43.830 158.800 ;
        RECT 45.680 155.600 63.830 158.800 ;
        RECT 65.680 155.600 83.830 158.800 ;
        RECT 85.680 155.600 103.830 158.800 ;
        RECT 4.730 153.200 104.730 155.600 ;
        RECT 5.630 146.800 23.830 153.200 ;
        RECT 25.630 146.800 43.830 153.200 ;
        RECT 45.630 146.800 63.830 153.200 ;
        RECT 65.630 146.800 83.830 153.200 ;
        RECT 85.630 146.800 103.830 153.200 ;
        RECT 4.730 144.400 104.730 146.800 ;
        RECT 5.630 140.900 23.830 144.400 ;
        RECT 25.630 140.900 43.830 144.400 ;
        RECT 45.630 140.900 63.830 144.400 ;
        RECT 65.630 140.900 83.830 144.400 ;
        RECT 85.630 140.900 103.830 144.400 ;
        RECT 9.130 139.100 11.530 140.900 ;
        RECT 17.930 139.100 20.330 140.900 ;
        RECT 29.130 139.100 31.530 140.900 ;
        RECT 37.930 139.100 40.330 140.900 ;
        RECT 49.130 139.100 51.530 140.900 ;
        RECT 57.930 139.100 60.330 140.900 ;
        RECT 69.130 139.100 71.530 140.900 ;
        RECT 77.930 139.100 80.330 140.900 ;
        RECT 89.130 139.100 91.530 140.900 ;
        RECT 97.930 139.100 100.330 140.900 ;
        RECT 5.880 138.900 23.830 139.100 ;
        RECT 25.880 138.900 43.830 139.100 ;
        RECT 45.880 138.900 63.830 139.100 ;
        RECT 65.880 138.900 83.830 139.100 ;
        RECT 85.880 138.900 103.830 139.100 ;
        RECT 5.830 138.800 23.830 138.900 ;
        RECT 25.830 138.800 43.830 138.900 ;
        RECT 45.830 138.800 63.830 138.900 ;
        RECT 65.830 138.800 83.830 138.900 ;
        RECT 85.830 138.800 103.830 138.900 ;
        RECT 5.680 135.600 23.830 138.800 ;
        RECT 25.680 135.600 43.830 138.800 ;
        RECT 45.680 135.600 63.830 138.800 ;
        RECT 65.680 135.600 83.830 138.800 ;
        RECT 85.680 135.600 103.830 138.800 ;
        RECT 4.730 133.200 104.730 135.600 ;
        RECT 5.630 126.800 23.830 133.200 ;
        RECT 25.630 126.800 43.830 133.200 ;
        RECT 45.630 126.800 63.830 133.200 ;
        RECT 65.630 126.800 83.830 133.200 ;
        RECT 85.630 126.800 103.830 133.200 ;
        RECT 4.730 124.400 104.730 126.800 ;
        RECT 5.630 120.900 23.830 124.400 ;
        RECT 25.630 120.900 43.830 124.400 ;
        RECT 45.630 120.900 63.830 124.400 ;
        RECT 65.630 120.900 83.830 124.400 ;
        RECT 85.630 120.900 103.830 124.400 ;
        RECT 9.130 119.100 11.530 120.900 ;
        RECT 17.930 119.100 20.330 120.900 ;
        RECT 29.130 119.100 31.530 120.900 ;
        RECT 37.930 119.100 40.330 120.900 ;
        RECT 49.130 119.100 51.530 120.900 ;
        RECT 57.930 119.100 60.330 120.900 ;
        RECT 69.130 119.100 71.530 120.900 ;
        RECT 77.930 119.100 80.330 120.900 ;
        RECT 89.130 119.100 91.530 120.900 ;
        RECT 97.930 119.100 100.330 120.900 ;
        RECT 5.880 118.900 23.830 119.100 ;
        RECT 25.880 118.900 43.830 119.100 ;
        RECT 45.880 118.900 63.830 119.100 ;
        RECT 65.880 118.900 83.830 119.100 ;
        RECT 85.880 118.900 103.830 119.100 ;
        RECT 5.830 118.800 23.830 118.900 ;
        RECT 25.830 118.800 43.830 118.900 ;
        RECT 45.830 118.800 63.830 118.900 ;
        RECT 65.830 118.800 83.830 118.900 ;
        RECT 85.830 118.800 103.830 118.900 ;
        RECT 5.680 115.600 23.830 118.800 ;
        RECT 25.680 115.600 43.830 118.800 ;
        RECT 45.680 115.600 63.830 118.800 ;
        RECT 65.680 115.600 83.830 118.800 ;
        RECT 85.680 115.600 103.830 118.800 ;
        RECT 4.730 113.200 104.730 115.600 ;
        RECT 5.630 106.800 23.830 113.200 ;
        RECT 25.630 106.800 43.830 113.200 ;
        RECT 45.630 106.800 63.830 113.200 ;
        RECT 65.630 106.800 83.830 113.200 ;
        RECT 85.630 106.800 103.830 113.200 ;
        RECT 4.730 104.400 104.730 106.800 ;
        RECT 5.630 100.900 23.830 104.400 ;
        RECT 25.630 100.900 43.830 104.400 ;
        RECT 45.630 100.900 63.830 104.400 ;
        RECT 65.630 100.900 83.830 104.400 ;
        RECT 85.630 100.900 103.830 104.400 ;
        RECT 9.130 99.100 11.530 100.900 ;
        RECT 17.930 99.100 20.330 100.900 ;
        RECT 29.130 99.100 31.530 100.900 ;
        RECT 37.930 99.100 40.330 100.900 ;
        RECT 49.130 99.100 51.530 100.900 ;
        RECT 57.930 99.100 60.330 100.900 ;
        RECT 69.130 99.100 71.530 100.900 ;
        RECT 77.930 99.100 80.330 100.900 ;
        RECT 89.130 99.100 91.530 100.900 ;
        RECT 97.930 99.100 100.330 100.900 ;
        RECT 5.880 98.900 23.830 99.100 ;
        RECT 25.880 98.900 43.830 99.100 ;
        RECT 45.880 98.900 63.830 99.100 ;
        RECT 65.880 98.900 83.830 99.100 ;
        RECT 85.880 98.900 103.830 99.100 ;
        RECT 5.830 98.800 23.830 98.900 ;
        RECT 25.830 98.800 43.830 98.900 ;
        RECT 45.830 98.800 63.830 98.900 ;
        RECT 65.830 98.800 83.830 98.900 ;
        RECT 85.830 98.800 103.830 98.900 ;
        RECT 5.680 95.600 23.830 98.800 ;
        RECT 25.680 95.600 43.830 98.800 ;
        RECT 45.680 95.600 63.830 98.800 ;
        RECT 65.680 95.600 83.830 98.800 ;
        RECT 85.680 95.600 103.830 98.800 ;
        RECT 4.730 93.200 104.730 95.600 ;
        RECT 5.630 86.800 23.830 93.200 ;
        RECT 25.630 86.800 43.830 93.200 ;
        RECT 45.630 86.800 63.830 93.200 ;
        RECT 65.630 86.800 83.830 93.200 ;
        RECT 85.630 86.800 103.830 93.200 ;
        RECT 4.730 84.400 104.730 86.800 ;
        RECT 5.630 80.900 23.830 84.400 ;
        RECT 25.630 80.900 43.830 84.400 ;
        RECT 45.630 80.900 63.830 84.400 ;
        RECT 65.630 80.900 83.830 84.400 ;
        RECT 85.630 80.900 103.830 84.400 ;
        RECT 9.130 79.100 11.530 80.900 ;
        RECT 17.930 79.100 20.330 80.900 ;
        RECT 29.130 79.100 31.530 80.900 ;
        RECT 37.930 79.100 40.330 80.900 ;
        RECT 49.130 79.100 51.530 80.900 ;
        RECT 57.930 79.100 60.330 80.900 ;
        RECT 69.130 79.100 71.530 80.900 ;
        RECT 77.930 79.100 80.330 80.900 ;
        RECT 89.130 79.100 91.530 80.900 ;
        RECT 97.930 79.100 100.330 80.900 ;
        RECT 5.880 78.900 23.830 79.100 ;
        RECT 25.880 78.900 43.830 79.100 ;
        RECT 45.880 78.900 63.830 79.100 ;
        RECT 65.880 78.900 83.830 79.100 ;
        RECT 85.880 78.900 103.830 79.100 ;
        RECT 5.830 78.800 23.830 78.900 ;
        RECT 25.830 78.800 43.830 78.900 ;
        RECT 45.830 78.800 63.830 78.900 ;
        RECT 65.830 78.800 83.830 78.900 ;
        RECT 85.830 78.800 103.830 78.900 ;
        RECT 5.680 75.600 23.830 78.800 ;
        RECT 25.680 75.600 43.830 78.800 ;
        RECT 45.680 75.600 63.830 78.800 ;
        RECT 65.680 75.600 83.830 78.800 ;
        RECT 85.680 75.600 103.830 78.800 ;
        RECT 4.730 73.200 104.730 75.600 ;
        RECT 5.630 66.800 23.830 73.200 ;
        RECT 25.630 66.800 43.830 73.200 ;
        RECT 45.630 66.800 63.830 73.200 ;
        RECT 65.630 66.800 83.830 73.200 ;
        RECT 85.630 66.800 103.830 73.200 ;
        RECT 4.730 64.400 104.730 66.800 ;
        RECT 5.630 60.900 23.830 64.400 ;
        RECT 25.630 60.900 43.830 64.400 ;
        RECT 45.630 60.900 63.830 64.400 ;
        RECT 65.630 60.900 83.830 64.400 ;
        RECT 85.630 60.900 103.830 64.400 ;
        RECT 9.130 59.100 11.530 60.900 ;
        RECT 17.930 59.100 20.330 60.900 ;
        RECT 29.130 59.100 31.530 60.900 ;
        RECT 37.930 59.100 40.330 60.900 ;
        RECT 49.130 59.100 51.530 60.900 ;
        RECT 57.930 59.100 60.330 60.900 ;
        RECT 69.130 59.100 71.530 60.900 ;
        RECT 77.930 59.100 80.330 60.900 ;
        RECT 89.130 59.100 91.530 60.900 ;
        RECT 97.930 59.100 100.330 60.900 ;
        RECT 5.880 58.900 23.830 59.100 ;
        RECT 25.880 58.900 43.830 59.100 ;
        RECT 45.880 58.900 63.830 59.100 ;
        RECT 65.880 58.900 83.830 59.100 ;
        RECT 85.880 58.900 103.830 59.100 ;
        RECT 5.830 58.800 23.830 58.900 ;
        RECT 25.830 58.800 43.830 58.900 ;
        RECT 45.830 58.800 63.830 58.900 ;
        RECT 65.830 58.800 83.830 58.900 ;
        RECT 85.830 58.800 103.830 58.900 ;
        RECT 5.680 55.600 23.830 58.800 ;
        RECT 25.680 55.600 43.830 58.800 ;
        RECT 45.680 55.600 63.830 58.800 ;
        RECT 65.680 55.600 83.830 58.800 ;
        RECT 85.680 55.600 103.830 58.800 ;
        RECT 4.730 53.200 104.730 55.600 ;
        RECT 5.630 46.800 23.830 53.200 ;
        RECT 25.630 46.800 43.830 53.200 ;
        RECT 45.630 46.800 63.830 53.200 ;
        RECT 65.630 46.800 83.830 53.200 ;
        RECT 85.630 46.800 103.830 53.200 ;
        RECT 4.730 44.400 104.730 46.800 ;
        RECT 5.630 40.900 23.830 44.400 ;
        RECT 25.630 40.900 43.830 44.400 ;
        RECT 45.630 40.900 63.830 44.400 ;
        RECT 65.630 40.900 83.830 44.400 ;
        RECT 85.630 40.900 103.830 44.400 ;
        RECT 9.130 39.100 11.530 40.900 ;
        RECT 17.930 39.100 20.330 40.900 ;
        RECT 29.130 39.100 31.530 40.900 ;
        RECT 37.930 39.100 40.330 40.900 ;
        RECT 49.130 39.100 51.530 40.900 ;
        RECT 57.930 39.100 60.330 40.900 ;
        RECT 69.130 39.100 71.530 40.900 ;
        RECT 77.930 39.100 80.330 40.900 ;
        RECT 89.130 39.100 91.530 40.900 ;
        RECT 97.930 39.100 100.330 40.900 ;
        RECT 5.880 38.900 23.830 39.100 ;
        RECT 25.880 38.900 43.830 39.100 ;
        RECT 45.880 38.900 63.830 39.100 ;
        RECT 65.880 38.900 83.830 39.100 ;
        RECT 85.880 38.900 103.830 39.100 ;
        RECT 5.830 38.800 23.830 38.900 ;
        RECT 25.830 38.800 43.830 38.900 ;
        RECT 45.830 38.800 63.830 38.900 ;
        RECT 65.830 38.800 83.830 38.900 ;
        RECT 85.830 38.800 103.830 38.900 ;
        RECT 5.680 35.600 23.830 38.800 ;
        RECT 25.680 35.600 43.830 38.800 ;
        RECT 45.680 35.600 63.830 38.800 ;
        RECT 65.680 35.600 83.830 38.800 ;
        RECT 85.680 35.600 103.830 38.800 ;
        RECT 4.730 33.200 104.730 35.600 ;
        RECT 5.630 26.800 23.830 33.200 ;
        RECT 25.630 26.800 43.830 33.200 ;
        RECT 45.630 26.800 63.830 33.200 ;
        RECT 65.630 26.800 83.830 33.200 ;
        RECT 85.630 26.800 103.830 33.200 ;
        RECT 4.730 24.400 104.730 26.800 ;
        RECT 5.630 20.900 23.830 24.400 ;
        RECT 25.630 20.900 43.830 24.400 ;
        RECT 45.630 20.900 63.830 24.400 ;
        RECT 65.630 20.900 83.830 24.400 ;
        RECT 85.630 20.900 103.830 24.400 ;
        RECT 9.130 19.100 11.530 20.900 ;
        RECT 17.930 19.100 20.330 20.900 ;
        RECT 29.130 19.100 31.530 20.900 ;
        RECT 37.930 19.100 40.330 20.900 ;
        RECT 49.130 19.100 51.530 20.900 ;
        RECT 57.930 19.100 60.330 20.900 ;
        RECT 69.130 19.100 71.530 20.900 ;
        RECT 77.930 19.100 80.330 20.900 ;
        RECT 89.130 19.100 91.530 20.900 ;
        RECT 97.930 19.100 100.330 20.900 ;
        RECT 5.880 18.900 23.830 19.100 ;
        RECT 25.880 18.900 43.830 19.100 ;
        RECT 45.880 18.900 63.830 19.100 ;
        RECT 65.880 18.900 83.830 19.100 ;
        RECT 85.880 18.900 103.830 19.100 ;
        RECT 5.830 18.800 23.830 18.900 ;
        RECT 25.830 18.800 43.830 18.900 ;
        RECT 45.830 18.800 63.830 18.900 ;
        RECT 65.830 18.800 83.830 18.900 ;
        RECT 85.830 18.800 103.830 18.900 ;
        RECT 5.680 15.600 23.830 18.800 ;
        RECT 25.680 15.600 43.830 18.800 ;
        RECT 45.680 15.600 63.830 18.800 ;
        RECT 65.680 15.600 83.830 18.800 ;
        RECT 85.680 15.600 103.830 18.800 ;
        RECT 4.730 13.200 104.730 15.600 ;
        RECT 5.630 6.800 23.830 13.200 ;
        RECT 25.630 6.800 43.830 13.200 ;
        RECT 45.630 6.800 63.830 13.200 ;
        RECT 65.630 6.800 83.830 13.200 ;
        RECT 85.630 6.800 103.830 13.200 ;
        RECT 4.730 4.400 104.730 6.800 ;
        RECT 5.630 0.900 23.830 4.400 ;
        RECT 25.630 0.900 43.830 4.400 ;
        RECT 45.630 0.900 63.830 4.400 ;
        RECT 65.630 0.900 83.830 4.400 ;
        RECT 85.630 0.900 103.830 4.400 ;
        RECT 9.130 0.000 11.530 0.900 ;
        RECT 17.930 0.000 20.330 0.900 ;
        RECT 29.130 0.000 31.530 0.900 ;
        RECT 37.930 0.000 40.330 0.900 ;
        RECT 49.130 0.000 51.530 0.900 ;
        RECT 57.930 0.000 60.330 0.900 ;
        RECT 69.130 0.000 71.530 0.900 ;
        RECT 77.930 0.000 80.330 0.900 ;
        RECT 89.130 0.000 91.530 0.900 ;
        RECT 97.930 0.000 100.330 0.900 ;
      LAYER li1 ;
        RECT 9.180 379.600 11.480 380.000 ;
        RECT 17.980 379.600 20.280 380.000 ;
        RECT 29.180 379.600 31.480 380.000 ;
        RECT 37.980 379.600 40.280 380.000 ;
        RECT 49.180 379.600 51.480 380.000 ;
        RECT 57.980 379.600 60.280 380.000 ;
        RECT 69.180 379.600 71.480 380.000 ;
        RECT 77.980 379.600 80.280 380.000 ;
        RECT 89.180 379.600 91.480 380.000 ;
        RECT 97.980 379.600 100.280 380.000 ;
        RECT 5.130 379.200 24.330 379.600 ;
        RECT 2.515 376.880 2.875 377.260 ;
        RECT 3.145 376.880 3.505 377.260 ;
        RECT 3.745 376.880 4.105 377.260 ;
        RECT 2.515 376.290 2.875 376.670 ;
        RECT 3.145 376.290 3.505 376.670 ;
        RECT 3.745 376.290 4.105 376.670 ;
        RECT 5.130 375.550 5.530 379.200 ;
        RECT 9.180 379.150 11.480 379.200 ;
        RECT 17.980 379.150 20.280 379.200 ;
        RECT 6.530 378.000 22.930 378.600 ;
        RECT 10.130 377.400 10.480 378.000 ;
        RECT 6.530 377.200 10.480 377.400 ;
        RECT 10.130 376.600 10.480 377.200 ;
        RECT 6.530 376.400 10.480 376.600 ;
        RECT 10.130 375.800 10.480 376.400 ;
        RECT 6.530 375.600 10.480 375.800 ;
        RECT 4.730 375.545 5.580 375.550 ;
        RECT 2.315 373.250 5.580 375.545 ;
        RECT 10.130 375.000 10.480 375.600 ;
        RECT 6.530 374.800 10.480 375.000 ;
        RECT 10.130 374.200 10.480 374.800 ;
        RECT 6.530 374.000 10.480 374.200 ;
        RECT 10.130 373.400 10.480 374.000 ;
        RECT 5.130 366.750 5.530 373.250 ;
        RECT 6.530 373.200 10.480 373.400 ;
        RECT 10.130 372.600 10.480 373.200 ;
        RECT 6.530 372.400 10.480 372.600 ;
        RECT 10.130 371.800 10.480 372.400 ;
        RECT 6.530 371.600 10.480 371.800 ;
        RECT 10.130 371.000 10.480 371.600 ;
        RECT 6.530 370.800 10.480 371.000 ;
        RECT 10.130 370.400 10.480 370.800 ;
        RECT 11.080 370.400 11.280 378.000 ;
        RECT 11.880 370.400 12.080 378.000 ;
        RECT 12.680 370.400 12.880 378.000 ;
        RECT 13.480 370.400 13.680 378.000 ;
        RECT 10.130 369.200 10.480 369.600 ;
        RECT 6.530 369.000 10.480 369.200 ;
        RECT 10.130 368.400 10.480 369.000 ;
        RECT 6.530 368.200 10.480 368.400 ;
        RECT 10.130 367.600 10.480 368.200 ;
        RECT 6.530 367.400 10.480 367.600 ;
        RECT 10.130 366.800 10.480 367.400 ;
        RECT 4.730 366.745 5.580 366.750 ;
        RECT 2.315 364.450 5.580 366.745 ;
        RECT 6.530 366.600 10.480 366.800 ;
        RECT 10.130 366.000 10.480 366.600 ;
        RECT 6.530 365.800 10.480 366.000 ;
        RECT 10.130 365.200 10.480 365.800 ;
        RECT 6.530 365.000 10.480 365.200 ;
        RECT 2.515 363.515 2.875 363.895 ;
        RECT 3.145 363.515 3.505 363.895 ;
        RECT 3.745 363.515 4.105 363.895 ;
        RECT 2.515 362.925 2.875 363.305 ;
        RECT 3.145 362.925 3.505 363.305 ;
        RECT 3.745 362.925 4.105 363.305 ;
        RECT 5.130 360.800 5.530 364.450 ;
        RECT 10.130 364.400 10.480 365.000 ;
        RECT 6.530 364.200 10.480 364.400 ;
        RECT 10.130 363.600 10.480 364.200 ;
        RECT 6.530 363.400 10.480 363.600 ;
        RECT 10.130 362.800 10.480 363.400 ;
        RECT 6.530 362.600 10.480 362.800 ;
        RECT 10.130 362.000 10.480 362.600 ;
        RECT 11.080 362.000 11.280 369.600 ;
        RECT 11.880 362.000 12.080 369.600 ;
        RECT 12.680 362.000 12.880 369.600 ;
        RECT 13.480 362.000 13.680 369.600 ;
        RECT 14.280 362.000 15.180 378.000 ;
        RECT 15.780 370.400 15.980 378.000 ;
        RECT 16.580 370.400 16.780 378.000 ;
        RECT 17.380 370.400 17.580 378.000 ;
        RECT 18.180 370.400 18.380 378.000 ;
        RECT 18.980 377.400 19.330 378.000 ;
        RECT 18.980 377.200 22.930 377.400 ;
        RECT 18.980 376.600 19.330 377.200 ;
        RECT 18.980 376.400 22.930 376.600 ;
        RECT 18.980 375.800 19.330 376.400 ;
        RECT 18.980 375.600 22.930 375.800 ;
        RECT 18.980 375.000 19.330 375.600 ;
        RECT 23.930 375.550 24.330 379.200 ;
        RECT 25.130 379.200 44.330 379.600 ;
        RECT 25.130 375.550 25.530 379.200 ;
        RECT 29.180 379.150 31.480 379.200 ;
        RECT 37.980 379.150 40.280 379.200 ;
        RECT 26.530 378.000 42.930 378.600 ;
        RECT 30.130 377.400 30.480 378.000 ;
        RECT 26.530 377.200 30.480 377.400 ;
        RECT 30.130 376.600 30.480 377.200 ;
        RECT 26.530 376.400 30.480 376.600 ;
        RECT 30.130 375.800 30.480 376.400 ;
        RECT 26.530 375.600 30.480 375.800 ;
        RECT 18.980 374.800 22.930 375.000 ;
        RECT 18.980 374.200 19.330 374.800 ;
        RECT 18.980 374.000 22.930 374.200 ;
        RECT 18.980 373.400 19.330 374.000 ;
        RECT 18.980 373.200 22.930 373.400 ;
        RECT 23.880 373.250 25.580 375.550 ;
        RECT 30.130 375.000 30.480 375.600 ;
        RECT 26.530 374.800 30.480 375.000 ;
        RECT 30.130 374.200 30.480 374.800 ;
        RECT 26.530 374.000 30.480 374.200 ;
        RECT 30.130 373.400 30.480 374.000 ;
        RECT 18.980 372.600 19.330 373.200 ;
        RECT 18.980 372.400 22.930 372.600 ;
        RECT 18.980 371.800 19.330 372.400 ;
        RECT 18.980 371.600 22.930 371.800 ;
        RECT 18.980 371.000 19.330 371.600 ;
        RECT 18.980 370.800 22.930 371.000 ;
        RECT 18.980 370.400 19.330 370.800 ;
        RECT 15.780 362.000 15.980 369.600 ;
        RECT 16.580 362.000 16.780 369.600 ;
        RECT 17.380 362.000 17.580 369.600 ;
        RECT 18.180 362.000 18.380 369.600 ;
        RECT 18.980 369.200 19.330 369.600 ;
        RECT 18.980 369.000 22.930 369.200 ;
        RECT 18.980 368.400 19.330 369.000 ;
        RECT 18.980 368.200 22.930 368.400 ;
        RECT 18.980 367.600 19.330 368.200 ;
        RECT 18.980 367.400 22.930 367.600 ;
        RECT 18.980 366.800 19.330 367.400 ;
        RECT 18.980 366.600 22.930 366.800 ;
        RECT 23.930 366.750 24.330 373.250 ;
        RECT 25.130 366.750 25.530 373.250 ;
        RECT 26.530 373.200 30.480 373.400 ;
        RECT 30.130 372.600 30.480 373.200 ;
        RECT 26.530 372.400 30.480 372.600 ;
        RECT 30.130 371.800 30.480 372.400 ;
        RECT 26.530 371.600 30.480 371.800 ;
        RECT 30.130 371.000 30.480 371.600 ;
        RECT 26.530 370.800 30.480 371.000 ;
        RECT 30.130 370.400 30.480 370.800 ;
        RECT 31.080 370.400 31.280 378.000 ;
        RECT 31.880 370.400 32.080 378.000 ;
        RECT 32.680 370.400 32.880 378.000 ;
        RECT 33.480 370.400 33.680 378.000 ;
        RECT 30.130 369.200 30.480 369.600 ;
        RECT 26.530 369.000 30.480 369.200 ;
        RECT 30.130 368.400 30.480 369.000 ;
        RECT 26.530 368.200 30.480 368.400 ;
        RECT 30.130 367.600 30.480 368.200 ;
        RECT 26.530 367.400 30.480 367.600 ;
        RECT 30.130 366.800 30.480 367.400 ;
        RECT 18.980 366.000 19.330 366.600 ;
        RECT 18.980 365.800 22.930 366.000 ;
        RECT 18.980 365.200 19.330 365.800 ;
        RECT 18.980 365.000 22.930 365.200 ;
        RECT 18.980 364.400 19.330 365.000 ;
        RECT 23.880 364.450 25.580 366.750 ;
        RECT 26.530 366.600 30.480 366.800 ;
        RECT 30.130 366.000 30.480 366.600 ;
        RECT 26.530 365.800 30.480 366.000 ;
        RECT 30.130 365.200 30.480 365.800 ;
        RECT 26.530 365.000 30.480 365.200 ;
        RECT 18.980 364.200 22.930 364.400 ;
        RECT 18.980 363.600 19.330 364.200 ;
        RECT 18.980 363.400 22.930 363.600 ;
        RECT 18.980 362.800 19.330 363.400 ;
        RECT 18.980 362.600 22.930 362.800 ;
        RECT 18.980 362.000 19.330 362.600 ;
        RECT 6.530 361.400 22.930 362.000 ;
        RECT 9.180 360.800 11.480 360.850 ;
        RECT 17.980 360.800 20.280 360.850 ;
        RECT 23.930 360.800 24.330 364.450 ;
        RECT 5.130 360.400 24.330 360.800 ;
        RECT 25.130 360.800 25.530 364.450 ;
        RECT 30.130 364.400 30.480 365.000 ;
        RECT 26.530 364.200 30.480 364.400 ;
        RECT 30.130 363.600 30.480 364.200 ;
        RECT 26.530 363.400 30.480 363.600 ;
        RECT 30.130 362.800 30.480 363.400 ;
        RECT 26.530 362.600 30.480 362.800 ;
        RECT 30.130 362.000 30.480 362.600 ;
        RECT 31.080 362.000 31.280 369.600 ;
        RECT 31.880 362.000 32.080 369.600 ;
        RECT 32.680 362.000 32.880 369.600 ;
        RECT 33.480 362.000 33.680 369.600 ;
        RECT 34.280 362.000 35.180 378.000 ;
        RECT 35.780 370.400 35.980 378.000 ;
        RECT 36.580 370.400 36.780 378.000 ;
        RECT 37.380 370.400 37.580 378.000 ;
        RECT 38.180 370.400 38.380 378.000 ;
        RECT 38.980 377.400 39.330 378.000 ;
        RECT 38.980 377.200 42.930 377.400 ;
        RECT 38.980 376.600 39.330 377.200 ;
        RECT 38.980 376.400 42.930 376.600 ;
        RECT 38.980 375.800 39.330 376.400 ;
        RECT 38.980 375.600 42.930 375.800 ;
        RECT 38.980 375.000 39.330 375.600 ;
        RECT 43.930 375.550 44.330 379.200 ;
        RECT 45.130 379.200 64.330 379.600 ;
        RECT 45.130 375.550 45.530 379.200 ;
        RECT 49.180 379.150 51.480 379.200 ;
        RECT 57.980 379.150 60.280 379.200 ;
        RECT 46.530 378.000 62.930 378.600 ;
        RECT 50.130 377.400 50.480 378.000 ;
        RECT 46.530 377.200 50.480 377.400 ;
        RECT 50.130 376.600 50.480 377.200 ;
        RECT 46.530 376.400 50.480 376.600 ;
        RECT 50.130 375.800 50.480 376.400 ;
        RECT 46.530 375.600 50.480 375.800 ;
        RECT 38.980 374.800 42.930 375.000 ;
        RECT 38.980 374.200 39.330 374.800 ;
        RECT 38.980 374.000 42.930 374.200 ;
        RECT 38.980 373.400 39.330 374.000 ;
        RECT 38.980 373.200 42.930 373.400 ;
        RECT 43.880 373.250 45.580 375.550 ;
        RECT 50.130 375.000 50.480 375.600 ;
        RECT 46.530 374.800 50.480 375.000 ;
        RECT 50.130 374.200 50.480 374.800 ;
        RECT 46.530 374.000 50.480 374.200 ;
        RECT 50.130 373.400 50.480 374.000 ;
        RECT 38.980 372.600 39.330 373.200 ;
        RECT 38.980 372.400 42.930 372.600 ;
        RECT 38.980 371.800 39.330 372.400 ;
        RECT 38.980 371.600 42.930 371.800 ;
        RECT 38.980 371.000 39.330 371.600 ;
        RECT 38.980 370.800 42.930 371.000 ;
        RECT 38.980 370.400 39.330 370.800 ;
        RECT 35.780 362.000 35.980 369.600 ;
        RECT 36.580 362.000 36.780 369.600 ;
        RECT 37.380 362.000 37.580 369.600 ;
        RECT 38.180 362.000 38.380 369.600 ;
        RECT 38.980 369.200 39.330 369.600 ;
        RECT 38.980 369.000 42.930 369.200 ;
        RECT 38.980 368.400 39.330 369.000 ;
        RECT 38.980 368.200 42.930 368.400 ;
        RECT 38.980 367.600 39.330 368.200 ;
        RECT 38.980 367.400 42.930 367.600 ;
        RECT 38.980 366.800 39.330 367.400 ;
        RECT 38.980 366.600 42.930 366.800 ;
        RECT 43.930 366.750 44.330 373.250 ;
        RECT 45.130 366.750 45.530 373.250 ;
        RECT 46.530 373.200 50.480 373.400 ;
        RECT 50.130 372.600 50.480 373.200 ;
        RECT 46.530 372.400 50.480 372.600 ;
        RECT 50.130 371.800 50.480 372.400 ;
        RECT 46.530 371.600 50.480 371.800 ;
        RECT 50.130 371.000 50.480 371.600 ;
        RECT 46.530 370.800 50.480 371.000 ;
        RECT 50.130 370.400 50.480 370.800 ;
        RECT 51.080 370.400 51.280 378.000 ;
        RECT 51.880 370.400 52.080 378.000 ;
        RECT 52.680 370.400 52.880 378.000 ;
        RECT 53.480 370.400 53.680 378.000 ;
        RECT 50.130 369.200 50.480 369.600 ;
        RECT 46.530 369.000 50.480 369.200 ;
        RECT 50.130 368.400 50.480 369.000 ;
        RECT 46.530 368.200 50.480 368.400 ;
        RECT 50.130 367.600 50.480 368.200 ;
        RECT 46.530 367.400 50.480 367.600 ;
        RECT 50.130 366.800 50.480 367.400 ;
        RECT 38.980 366.000 39.330 366.600 ;
        RECT 38.980 365.800 42.930 366.000 ;
        RECT 38.980 365.200 39.330 365.800 ;
        RECT 38.980 365.000 42.930 365.200 ;
        RECT 38.980 364.400 39.330 365.000 ;
        RECT 43.880 364.450 45.580 366.750 ;
        RECT 46.530 366.600 50.480 366.800 ;
        RECT 50.130 366.000 50.480 366.600 ;
        RECT 46.530 365.800 50.480 366.000 ;
        RECT 50.130 365.200 50.480 365.800 ;
        RECT 46.530 365.000 50.480 365.200 ;
        RECT 38.980 364.200 42.930 364.400 ;
        RECT 38.980 363.600 39.330 364.200 ;
        RECT 38.980 363.400 42.930 363.600 ;
        RECT 38.980 362.800 39.330 363.400 ;
        RECT 38.980 362.600 42.930 362.800 ;
        RECT 38.980 362.000 39.330 362.600 ;
        RECT 26.530 361.400 42.930 362.000 ;
        RECT 29.180 360.800 31.480 360.850 ;
        RECT 37.980 360.800 40.280 360.850 ;
        RECT 43.930 360.800 44.330 364.450 ;
        RECT 25.130 360.400 44.330 360.800 ;
        RECT 45.130 360.800 45.530 364.450 ;
        RECT 50.130 364.400 50.480 365.000 ;
        RECT 46.530 364.200 50.480 364.400 ;
        RECT 50.130 363.600 50.480 364.200 ;
        RECT 46.530 363.400 50.480 363.600 ;
        RECT 50.130 362.800 50.480 363.400 ;
        RECT 46.530 362.600 50.480 362.800 ;
        RECT 50.130 362.000 50.480 362.600 ;
        RECT 51.080 362.000 51.280 369.600 ;
        RECT 51.880 362.000 52.080 369.600 ;
        RECT 52.680 362.000 52.880 369.600 ;
        RECT 53.480 362.000 53.680 369.600 ;
        RECT 54.280 362.000 55.180 378.000 ;
        RECT 55.780 370.400 55.980 378.000 ;
        RECT 56.580 370.400 56.780 378.000 ;
        RECT 57.380 370.400 57.580 378.000 ;
        RECT 58.180 370.400 58.380 378.000 ;
        RECT 58.980 377.400 59.330 378.000 ;
        RECT 58.980 377.200 62.930 377.400 ;
        RECT 58.980 376.600 59.330 377.200 ;
        RECT 58.980 376.400 62.930 376.600 ;
        RECT 58.980 375.800 59.330 376.400 ;
        RECT 58.980 375.600 62.930 375.800 ;
        RECT 58.980 375.000 59.330 375.600 ;
        RECT 63.930 375.550 64.330 379.200 ;
        RECT 65.130 379.200 84.330 379.600 ;
        RECT 65.130 375.550 65.530 379.200 ;
        RECT 69.180 379.150 71.480 379.200 ;
        RECT 77.980 379.150 80.280 379.200 ;
        RECT 66.530 378.000 82.930 378.600 ;
        RECT 70.130 377.400 70.480 378.000 ;
        RECT 66.530 377.200 70.480 377.400 ;
        RECT 70.130 376.600 70.480 377.200 ;
        RECT 66.530 376.400 70.480 376.600 ;
        RECT 70.130 375.800 70.480 376.400 ;
        RECT 66.530 375.600 70.480 375.800 ;
        RECT 58.980 374.800 62.930 375.000 ;
        RECT 58.980 374.200 59.330 374.800 ;
        RECT 58.980 374.000 62.930 374.200 ;
        RECT 58.980 373.400 59.330 374.000 ;
        RECT 58.980 373.200 62.930 373.400 ;
        RECT 63.880 373.250 65.580 375.550 ;
        RECT 70.130 375.000 70.480 375.600 ;
        RECT 66.530 374.800 70.480 375.000 ;
        RECT 70.130 374.200 70.480 374.800 ;
        RECT 66.530 374.000 70.480 374.200 ;
        RECT 70.130 373.400 70.480 374.000 ;
        RECT 58.980 372.600 59.330 373.200 ;
        RECT 58.980 372.400 62.930 372.600 ;
        RECT 58.980 371.800 59.330 372.400 ;
        RECT 58.980 371.600 62.930 371.800 ;
        RECT 58.980 371.000 59.330 371.600 ;
        RECT 58.980 370.800 62.930 371.000 ;
        RECT 58.980 370.400 59.330 370.800 ;
        RECT 55.780 362.000 55.980 369.600 ;
        RECT 56.580 362.000 56.780 369.600 ;
        RECT 57.380 362.000 57.580 369.600 ;
        RECT 58.180 362.000 58.380 369.600 ;
        RECT 58.980 369.200 59.330 369.600 ;
        RECT 58.980 369.000 62.930 369.200 ;
        RECT 58.980 368.400 59.330 369.000 ;
        RECT 58.980 368.200 62.930 368.400 ;
        RECT 58.980 367.600 59.330 368.200 ;
        RECT 58.980 367.400 62.930 367.600 ;
        RECT 58.980 366.800 59.330 367.400 ;
        RECT 58.980 366.600 62.930 366.800 ;
        RECT 63.930 366.750 64.330 373.250 ;
        RECT 65.130 366.750 65.530 373.250 ;
        RECT 66.530 373.200 70.480 373.400 ;
        RECT 70.130 372.600 70.480 373.200 ;
        RECT 66.530 372.400 70.480 372.600 ;
        RECT 70.130 371.800 70.480 372.400 ;
        RECT 66.530 371.600 70.480 371.800 ;
        RECT 70.130 371.000 70.480 371.600 ;
        RECT 66.530 370.800 70.480 371.000 ;
        RECT 70.130 370.400 70.480 370.800 ;
        RECT 71.080 370.400 71.280 378.000 ;
        RECT 71.880 370.400 72.080 378.000 ;
        RECT 72.680 370.400 72.880 378.000 ;
        RECT 73.480 370.400 73.680 378.000 ;
        RECT 70.130 369.200 70.480 369.600 ;
        RECT 66.530 369.000 70.480 369.200 ;
        RECT 70.130 368.400 70.480 369.000 ;
        RECT 66.530 368.200 70.480 368.400 ;
        RECT 70.130 367.600 70.480 368.200 ;
        RECT 66.530 367.400 70.480 367.600 ;
        RECT 70.130 366.800 70.480 367.400 ;
        RECT 58.980 366.000 59.330 366.600 ;
        RECT 58.980 365.800 62.930 366.000 ;
        RECT 58.980 365.200 59.330 365.800 ;
        RECT 58.980 365.000 62.930 365.200 ;
        RECT 58.980 364.400 59.330 365.000 ;
        RECT 63.880 364.450 65.580 366.750 ;
        RECT 66.530 366.600 70.480 366.800 ;
        RECT 70.130 366.000 70.480 366.600 ;
        RECT 66.530 365.800 70.480 366.000 ;
        RECT 70.130 365.200 70.480 365.800 ;
        RECT 66.530 365.000 70.480 365.200 ;
        RECT 58.980 364.200 62.930 364.400 ;
        RECT 58.980 363.600 59.330 364.200 ;
        RECT 58.980 363.400 62.930 363.600 ;
        RECT 58.980 362.800 59.330 363.400 ;
        RECT 58.980 362.600 62.930 362.800 ;
        RECT 58.980 362.000 59.330 362.600 ;
        RECT 46.530 361.400 62.930 362.000 ;
        RECT 49.180 360.800 51.480 360.850 ;
        RECT 57.980 360.800 60.280 360.850 ;
        RECT 63.930 360.800 64.330 364.450 ;
        RECT 45.130 360.400 64.330 360.800 ;
        RECT 65.130 360.800 65.530 364.450 ;
        RECT 70.130 364.400 70.480 365.000 ;
        RECT 66.530 364.200 70.480 364.400 ;
        RECT 70.130 363.600 70.480 364.200 ;
        RECT 66.530 363.400 70.480 363.600 ;
        RECT 70.130 362.800 70.480 363.400 ;
        RECT 66.530 362.600 70.480 362.800 ;
        RECT 70.130 362.000 70.480 362.600 ;
        RECT 71.080 362.000 71.280 369.600 ;
        RECT 71.880 362.000 72.080 369.600 ;
        RECT 72.680 362.000 72.880 369.600 ;
        RECT 73.480 362.000 73.680 369.600 ;
        RECT 74.280 362.000 75.180 378.000 ;
        RECT 75.780 370.400 75.980 378.000 ;
        RECT 76.580 370.400 76.780 378.000 ;
        RECT 77.380 370.400 77.580 378.000 ;
        RECT 78.180 370.400 78.380 378.000 ;
        RECT 78.980 377.400 79.330 378.000 ;
        RECT 78.980 377.200 82.930 377.400 ;
        RECT 78.980 376.600 79.330 377.200 ;
        RECT 78.980 376.400 82.930 376.600 ;
        RECT 78.980 375.800 79.330 376.400 ;
        RECT 78.980 375.600 82.930 375.800 ;
        RECT 78.980 375.000 79.330 375.600 ;
        RECT 83.930 375.550 84.330 379.200 ;
        RECT 85.130 379.200 104.330 379.600 ;
        RECT 85.130 375.550 85.530 379.200 ;
        RECT 89.180 379.150 91.480 379.200 ;
        RECT 97.980 379.150 100.280 379.200 ;
        RECT 86.530 378.000 102.930 378.600 ;
        RECT 90.130 377.400 90.480 378.000 ;
        RECT 86.530 377.200 90.480 377.400 ;
        RECT 90.130 376.600 90.480 377.200 ;
        RECT 86.530 376.400 90.480 376.600 ;
        RECT 90.130 375.800 90.480 376.400 ;
        RECT 86.530 375.600 90.480 375.800 ;
        RECT 78.980 374.800 82.930 375.000 ;
        RECT 78.980 374.200 79.330 374.800 ;
        RECT 78.980 374.000 82.930 374.200 ;
        RECT 78.980 373.400 79.330 374.000 ;
        RECT 78.980 373.200 82.930 373.400 ;
        RECT 83.880 373.250 85.580 375.550 ;
        RECT 90.130 375.000 90.480 375.600 ;
        RECT 86.530 374.800 90.480 375.000 ;
        RECT 90.130 374.200 90.480 374.800 ;
        RECT 86.530 374.000 90.480 374.200 ;
        RECT 90.130 373.400 90.480 374.000 ;
        RECT 78.980 372.600 79.330 373.200 ;
        RECT 78.980 372.400 82.930 372.600 ;
        RECT 78.980 371.800 79.330 372.400 ;
        RECT 78.980 371.600 82.930 371.800 ;
        RECT 78.980 371.000 79.330 371.600 ;
        RECT 78.980 370.800 82.930 371.000 ;
        RECT 78.980 370.400 79.330 370.800 ;
        RECT 75.780 362.000 75.980 369.600 ;
        RECT 76.580 362.000 76.780 369.600 ;
        RECT 77.380 362.000 77.580 369.600 ;
        RECT 78.180 362.000 78.380 369.600 ;
        RECT 78.980 369.200 79.330 369.600 ;
        RECT 78.980 369.000 82.930 369.200 ;
        RECT 78.980 368.400 79.330 369.000 ;
        RECT 78.980 368.200 82.930 368.400 ;
        RECT 78.980 367.600 79.330 368.200 ;
        RECT 78.980 367.400 82.930 367.600 ;
        RECT 78.980 366.800 79.330 367.400 ;
        RECT 78.980 366.600 82.930 366.800 ;
        RECT 83.930 366.750 84.330 373.250 ;
        RECT 85.130 366.750 85.530 373.250 ;
        RECT 86.530 373.200 90.480 373.400 ;
        RECT 90.130 372.600 90.480 373.200 ;
        RECT 86.530 372.400 90.480 372.600 ;
        RECT 90.130 371.800 90.480 372.400 ;
        RECT 86.530 371.600 90.480 371.800 ;
        RECT 90.130 371.000 90.480 371.600 ;
        RECT 86.530 370.800 90.480 371.000 ;
        RECT 90.130 370.400 90.480 370.800 ;
        RECT 91.080 370.400 91.280 378.000 ;
        RECT 91.880 370.400 92.080 378.000 ;
        RECT 92.680 370.400 92.880 378.000 ;
        RECT 93.480 370.400 93.680 378.000 ;
        RECT 90.130 369.200 90.480 369.600 ;
        RECT 86.530 369.000 90.480 369.200 ;
        RECT 90.130 368.400 90.480 369.000 ;
        RECT 86.530 368.200 90.480 368.400 ;
        RECT 90.130 367.600 90.480 368.200 ;
        RECT 86.530 367.400 90.480 367.600 ;
        RECT 90.130 366.800 90.480 367.400 ;
        RECT 78.980 366.000 79.330 366.600 ;
        RECT 78.980 365.800 82.930 366.000 ;
        RECT 78.980 365.200 79.330 365.800 ;
        RECT 78.980 365.000 82.930 365.200 ;
        RECT 78.980 364.400 79.330 365.000 ;
        RECT 83.880 364.450 85.580 366.750 ;
        RECT 86.530 366.600 90.480 366.800 ;
        RECT 90.130 366.000 90.480 366.600 ;
        RECT 86.530 365.800 90.480 366.000 ;
        RECT 90.130 365.200 90.480 365.800 ;
        RECT 86.530 365.000 90.480 365.200 ;
        RECT 78.980 364.200 82.930 364.400 ;
        RECT 78.980 363.600 79.330 364.200 ;
        RECT 78.980 363.400 82.930 363.600 ;
        RECT 78.980 362.800 79.330 363.400 ;
        RECT 78.980 362.600 82.930 362.800 ;
        RECT 78.980 362.000 79.330 362.600 ;
        RECT 66.530 361.400 82.930 362.000 ;
        RECT 69.180 360.800 71.480 360.850 ;
        RECT 77.980 360.800 80.280 360.850 ;
        RECT 83.930 360.800 84.330 364.450 ;
        RECT 65.130 360.400 84.330 360.800 ;
        RECT 85.130 360.800 85.530 364.450 ;
        RECT 90.130 364.400 90.480 365.000 ;
        RECT 86.530 364.200 90.480 364.400 ;
        RECT 90.130 363.600 90.480 364.200 ;
        RECT 86.530 363.400 90.480 363.600 ;
        RECT 90.130 362.800 90.480 363.400 ;
        RECT 86.530 362.600 90.480 362.800 ;
        RECT 90.130 362.000 90.480 362.600 ;
        RECT 91.080 362.000 91.280 369.600 ;
        RECT 91.880 362.000 92.080 369.600 ;
        RECT 92.680 362.000 92.880 369.600 ;
        RECT 93.480 362.000 93.680 369.600 ;
        RECT 94.280 362.000 95.180 378.000 ;
        RECT 95.780 370.400 95.980 378.000 ;
        RECT 96.580 370.400 96.780 378.000 ;
        RECT 97.380 370.400 97.580 378.000 ;
        RECT 98.180 370.400 98.380 378.000 ;
        RECT 98.980 377.400 99.330 378.000 ;
        RECT 98.980 377.200 102.930 377.400 ;
        RECT 98.980 376.600 99.330 377.200 ;
        RECT 98.980 376.400 102.930 376.600 ;
        RECT 98.980 375.800 99.330 376.400 ;
        RECT 98.980 375.600 102.930 375.800 ;
        RECT 98.980 375.000 99.330 375.600 ;
        RECT 103.930 375.550 104.330 379.200 ;
        RECT 105.340 377.080 105.700 377.460 ;
        RECT 105.970 377.080 106.330 377.460 ;
        RECT 106.570 377.080 106.930 377.460 ;
        RECT 105.340 376.490 105.700 376.870 ;
        RECT 105.970 376.490 106.330 376.870 ;
        RECT 106.570 376.490 106.930 376.870 ;
        RECT 98.980 374.800 102.930 375.000 ;
        RECT 98.980 374.200 99.330 374.800 ;
        RECT 98.980 374.000 102.930 374.200 ;
        RECT 98.980 373.400 99.330 374.000 ;
        RECT 98.980 373.200 102.930 373.400 ;
        RECT 103.880 373.250 104.730 375.550 ;
        RECT 98.980 372.600 99.330 373.200 ;
        RECT 98.980 372.400 102.930 372.600 ;
        RECT 98.980 371.800 99.330 372.400 ;
        RECT 98.980 371.600 102.930 371.800 ;
        RECT 98.980 371.000 99.330 371.600 ;
        RECT 98.980 370.800 102.930 371.000 ;
        RECT 98.980 370.400 99.330 370.800 ;
        RECT 95.780 362.000 95.980 369.600 ;
        RECT 96.580 362.000 96.780 369.600 ;
        RECT 97.380 362.000 97.580 369.600 ;
        RECT 98.180 362.000 98.380 369.600 ;
        RECT 98.980 369.200 99.330 369.600 ;
        RECT 98.980 369.000 102.930 369.200 ;
        RECT 98.980 368.400 99.330 369.000 ;
        RECT 98.980 368.200 102.930 368.400 ;
        RECT 98.980 367.600 99.330 368.200 ;
        RECT 98.980 367.400 102.930 367.600 ;
        RECT 98.980 366.800 99.330 367.400 ;
        RECT 98.980 366.600 102.930 366.800 ;
        RECT 103.930 366.750 104.330 373.250 ;
        RECT 98.980 366.000 99.330 366.600 ;
        RECT 98.980 365.800 102.930 366.000 ;
        RECT 98.980 365.200 99.330 365.800 ;
        RECT 98.980 365.000 102.930 365.200 ;
        RECT 98.980 364.400 99.330 365.000 ;
        RECT 103.880 364.450 104.730 366.750 ;
        RECT 98.980 364.200 102.930 364.400 ;
        RECT 98.980 363.600 99.330 364.200 ;
        RECT 98.980 363.400 102.930 363.600 ;
        RECT 98.980 362.800 99.330 363.400 ;
        RECT 98.980 362.600 102.930 362.800 ;
        RECT 98.980 362.000 99.330 362.600 ;
        RECT 86.530 361.400 102.930 362.000 ;
        RECT 89.180 360.800 91.480 360.850 ;
        RECT 97.980 360.800 100.280 360.850 ;
        RECT 103.930 360.800 104.330 364.450 ;
        RECT 105.340 363.095 105.700 363.475 ;
        RECT 105.970 363.095 106.330 363.475 ;
        RECT 106.570 363.095 106.930 363.475 ;
        RECT 105.340 362.505 105.700 362.885 ;
        RECT 105.970 362.505 106.330 362.885 ;
        RECT 106.570 362.505 106.930 362.885 ;
        RECT 85.130 360.400 104.330 360.800 ;
        RECT 9.180 359.600 11.480 360.400 ;
        RECT 17.980 359.600 20.280 360.400 ;
        RECT 29.180 359.600 31.480 360.400 ;
        RECT 37.980 359.600 40.280 360.400 ;
        RECT 49.180 359.600 51.480 360.400 ;
        RECT 57.980 359.600 60.280 360.400 ;
        RECT 69.180 359.600 71.480 360.400 ;
        RECT 77.980 359.600 80.280 360.400 ;
        RECT 89.180 359.600 91.480 360.400 ;
        RECT 97.980 359.600 100.280 360.400 ;
        RECT 5.130 359.200 24.330 359.600 ;
        RECT 2.515 356.880 2.875 357.260 ;
        RECT 3.145 356.880 3.505 357.260 ;
        RECT 3.745 356.880 4.105 357.260 ;
        RECT 2.515 356.290 2.875 356.670 ;
        RECT 3.145 356.290 3.505 356.670 ;
        RECT 3.745 356.290 4.105 356.670 ;
        RECT 5.130 355.550 5.530 359.200 ;
        RECT 9.180 359.150 11.480 359.200 ;
        RECT 17.980 359.150 20.280 359.200 ;
        RECT 6.530 358.000 22.930 358.600 ;
        RECT 10.130 357.400 10.480 358.000 ;
        RECT 6.530 357.200 10.480 357.400 ;
        RECT 10.130 356.600 10.480 357.200 ;
        RECT 6.530 356.400 10.480 356.600 ;
        RECT 10.130 355.800 10.480 356.400 ;
        RECT 6.530 355.600 10.480 355.800 ;
        RECT 4.730 355.545 5.580 355.550 ;
        RECT 2.315 353.250 5.580 355.545 ;
        RECT 10.130 355.000 10.480 355.600 ;
        RECT 6.530 354.800 10.480 355.000 ;
        RECT 10.130 354.200 10.480 354.800 ;
        RECT 6.530 354.000 10.480 354.200 ;
        RECT 10.130 353.400 10.480 354.000 ;
        RECT 5.130 346.750 5.530 353.250 ;
        RECT 6.530 353.200 10.480 353.400 ;
        RECT 10.130 352.600 10.480 353.200 ;
        RECT 6.530 352.400 10.480 352.600 ;
        RECT 10.130 351.800 10.480 352.400 ;
        RECT 6.530 351.600 10.480 351.800 ;
        RECT 10.130 351.000 10.480 351.600 ;
        RECT 6.530 350.800 10.480 351.000 ;
        RECT 10.130 350.400 10.480 350.800 ;
        RECT 11.080 350.400 11.280 358.000 ;
        RECT 11.880 350.400 12.080 358.000 ;
        RECT 12.680 350.400 12.880 358.000 ;
        RECT 13.480 350.400 13.680 358.000 ;
        RECT 10.130 349.200 10.480 349.600 ;
        RECT 6.530 349.000 10.480 349.200 ;
        RECT 10.130 348.400 10.480 349.000 ;
        RECT 6.530 348.200 10.480 348.400 ;
        RECT 10.130 347.600 10.480 348.200 ;
        RECT 6.530 347.400 10.480 347.600 ;
        RECT 10.130 346.800 10.480 347.400 ;
        RECT 4.730 346.745 5.580 346.750 ;
        RECT 2.315 344.450 5.580 346.745 ;
        RECT 6.530 346.600 10.480 346.800 ;
        RECT 10.130 346.000 10.480 346.600 ;
        RECT 6.530 345.800 10.480 346.000 ;
        RECT 10.130 345.200 10.480 345.800 ;
        RECT 6.530 345.000 10.480 345.200 ;
        RECT 2.515 343.515 2.875 343.895 ;
        RECT 3.145 343.515 3.505 343.895 ;
        RECT 3.745 343.515 4.105 343.895 ;
        RECT 2.515 342.925 2.875 343.305 ;
        RECT 3.145 342.925 3.505 343.305 ;
        RECT 3.745 342.925 4.105 343.305 ;
        RECT 5.130 340.800 5.530 344.450 ;
        RECT 10.130 344.400 10.480 345.000 ;
        RECT 6.530 344.200 10.480 344.400 ;
        RECT 10.130 343.600 10.480 344.200 ;
        RECT 6.530 343.400 10.480 343.600 ;
        RECT 10.130 342.800 10.480 343.400 ;
        RECT 6.530 342.600 10.480 342.800 ;
        RECT 10.130 342.000 10.480 342.600 ;
        RECT 11.080 342.000 11.280 349.600 ;
        RECT 11.880 342.000 12.080 349.600 ;
        RECT 12.680 342.000 12.880 349.600 ;
        RECT 13.480 342.000 13.680 349.600 ;
        RECT 14.280 342.000 15.180 358.000 ;
        RECT 15.780 350.400 15.980 358.000 ;
        RECT 16.580 350.400 16.780 358.000 ;
        RECT 17.380 350.400 17.580 358.000 ;
        RECT 18.180 350.400 18.380 358.000 ;
        RECT 18.980 357.400 19.330 358.000 ;
        RECT 18.980 357.200 22.930 357.400 ;
        RECT 18.980 356.600 19.330 357.200 ;
        RECT 18.980 356.400 22.930 356.600 ;
        RECT 18.980 355.800 19.330 356.400 ;
        RECT 18.980 355.600 22.930 355.800 ;
        RECT 18.980 355.000 19.330 355.600 ;
        RECT 23.930 355.550 24.330 359.200 ;
        RECT 25.130 359.200 44.330 359.600 ;
        RECT 25.130 355.550 25.530 359.200 ;
        RECT 29.180 359.150 31.480 359.200 ;
        RECT 37.980 359.150 40.280 359.200 ;
        RECT 26.530 358.000 42.930 358.600 ;
        RECT 30.130 357.400 30.480 358.000 ;
        RECT 26.530 357.200 30.480 357.400 ;
        RECT 30.130 356.600 30.480 357.200 ;
        RECT 26.530 356.400 30.480 356.600 ;
        RECT 30.130 355.800 30.480 356.400 ;
        RECT 26.530 355.600 30.480 355.800 ;
        RECT 18.980 354.800 22.930 355.000 ;
        RECT 18.980 354.200 19.330 354.800 ;
        RECT 18.980 354.000 22.930 354.200 ;
        RECT 18.980 353.400 19.330 354.000 ;
        RECT 18.980 353.200 22.930 353.400 ;
        RECT 23.880 353.250 25.580 355.550 ;
        RECT 30.130 355.000 30.480 355.600 ;
        RECT 26.530 354.800 30.480 355.000 ;
        RECT 30.130 354.200 30.480 354.800 ;
        RECT 26.530 354.000 30.480 354.200 ;
        RECT 30.130 353.400 30.480 354.000 ;
        RECT 18.980 352.600 19.330 353.200 ;
        RECT 18.980 352.400 22.930 352.600 ;
        RECT 18.980 351.800 19.330 352.400 ;
        RECT 18.980 351.600 22.930 351.800 ;
        RECT 18.980 351.000 19.330 351.600 ;
        RECT 18.980 350.800 22.930 351.000 ;
        RECT 18.980 350.400 19.330 350.800 ;
        RECT 15.780 342.000 15.980 349.600 ;
        RECT 16.580 342.000 16.780 349.600 ;
        RECT 17.380 342.000 17.580 349.600 ;
        RECT 18.180 342.000 18.380 349.600 ;
        RECT 18.980 349.200 19.330 349.600 ;
        RECT 18.980 349.000 22.930 349.200 ;
        RECT 18.980 348.400 19.330 349.000 ;
        RECT 18.980 348.200 22.930 348.400 ;
        RECT 18.980 347.600 19.330 348.200 ;
        RECT 18.980 347.400 22.930 347.600 ;
        RECT 18.980 346.800 19.330 347.400 ;
        RECT 18.980 346.600 22.930 346.800 ;
        RECT 23.930 346.750 24.330 353.250 ;
        RECT 25.130 346.750 25.530 353.250 ;
        RECT 26.530 353.200 30.480 353.400 ;
        RECT 30.130 352.600 30.480 353.200 ;
        RECT 26.530 352.400 30.480 352.600 ;
        RECT 30.130 351.800 30.480 352.400 ;
        RECT 26.530 351.600 30.480 351.800 ;
        RECT 30.130 351.000 30.480 351.600 ;
        RECT 26.530 350.800 30.480 351.000 ;
        RECT 30.130 350.400 30.480 350.800 ;
        RECT 31.080 350.400 31.280 358.000 ;
        RECT 31.880 350.400 32.080 358.000 ;
        RECT 32.680 350.400 32.880 358.000 ;
        RECT 33.480 350.400 33.680 358.000 ;
        RECT 30.130 349.200 30.480 349.600 ;
        RECT 26.530 349.000 30.480 349.200 ;
        RECT 30.130 348.400 30.480 349.000 ;
        RECT 26.530 348.200 30.480 348.400 ;
        RECT 30.130 347.600 30.480 348.200 ;
        RECT 26.530 347.400 30.480 347.600 ;
        RECT 30.130 346.800 30.480 347.400 ;
        RECT 18.980 346.000 19.330 346.600 ;
        RECT 18.980 345.800 22.930 346.000 ;
        RECT 18.980 345.200 19.330 345.800 ;
        RECT 18.980 345.000 22.930 345.200 ;
        RECT 18.980 344.400 19.330 345.000 ;
        RECT 23.880 344.450 25.580 346.750 ;
        RECT 26.530 346.600 30.480 346.800 ;
        RECT 30.130 346.000 30.480 346.600 ;
        RECT 26.530 345.800 30.480 346.000 ;
        RECT 30.130 345.200 30.480 345.800 ;
        RECT 26.530 345.000 30.480 345.200 ;
        RECT 18.980 344.200 22.930 344.400 ;
        RECT 18.980 343.600 19.330 344.200 ;
        RECT 18.980 343.400 22.930 343.600 ;
        RECT 18.980 342.800 19.330 343.400 ;
        RECT 18.980 342.600 22.930 342.800 ;
        RECT 18.980 342.000 19.330 342.600 ;
        RECT 6.530 341.400 22.930 342.000 ;
        RECT 9.180 340.800 11.480 340.850 ;
        RECT 17.980 340.800 20.280 340.850 ;
        RECT 23.930 340.800 24.330 344.450 ;
        RECT 5.130 340.400 24.330 340.800 ;
        RECT 25.130 340.800 25.530 344.450 ;
        RECT 30.130 344.400 30.480 345.000 ;
        RECT 26.530 344.200 30.480 344.400 ;
        RECT 30.130 343.600 30.480 344.200 ;
        RECT 26.530 343.400 30.480 343.600 ;
        RECT 30.130 342.800 30.480 343.400 ;
        RECT 26.530 342.600 30.480 342.800 ;
        RECT 30.130 342.000 30.480 342.600 ;
        RECT 31.080 342.000 31.280 349.600 ;
        RECT 31.880 342.000 32.080 349.600 ;
        RECT 32.680 342.000 32.880 349.600 ;
        RECT 33.480 342.000 33.680 349.600 ;
        RECT 34.280 342.000 35.180 358.000 ;
        RECT 35.780 350.400 35.980 358.000 ;
        RECT 36.580 350.400 36.780 358.000 ;
        RECT 37.380 350.400 37.580 358.000 ;
        RECT 38.180 350.400 38.380 358.000 ;
        RECT 38.980 357.400 39.330 358.000 ;
        RECT 38.980 357.200 42.930 357.400 ;
        RECT 38.980 356.600 39.330 357.200 ;
        RECT 38.980 356.400 42.930 356.600 ;
        RECT 38.980 355.800 39.330 356.400 ;
        RECT 38.980 355.600 42.930 355.800 ;
        RECT 38.980 355.000 39.330 355.600 ;
        RECT 43.930 355.550 44.330 359.200 ;
        RECT 45.130 359.200 64.330 359.600 ;
        RECT 45.130 355.550 45.530 359.200 ;
        RECT 49.180 359.150 51.480 359.200 ;
        RECT 57.980 359.150 60.280 359.200 ;
        RECT 46.530 358.000 62.930 358.600 ;
        RECT 50.130 357.400 50.480 358.000 ;
        RECT 46.530 357.200 50.480 357.400 ;
        RECT 50.130 356.600 50.480 357.200 ;
        RECT 46.530 356.400 50.480 356.600 ;
        RECT 50.130 355.800 50.480 356.400 ;
        RECT 46.530 355.600 50.480 355.800 ;
        RECT 38.980 354.800 42.930 355.000 ;
        RECT 38.980 354.200 39.330 354.800 ;
        RECT 38.980 354.000 42.930 354.200 ;
        RECT 38.980 353.400 39.330 354.000 ;
        RECT 38.980 353.200 42.930 353.400 ;
        RECT 43.880 353.250 45.580 355.550 ;
        RECT 50.130 355.000 50.480 355.600 ;
        RECT 46.530 354.800 50.480 355.000 ;
        RECT 50.130 354.200 50.480 354.800 ;
        RECT 46.530 354.000 50.480 354.200 ;
        RECT 50.130 353.400 50.480 354.000 ;
        RECT 38.980 352.600 39.330 353.200 ;
        RECT 38.980 352.400 42.930 352.600 ;
        RECT 38.980 351.800 39.330 352.400 ;
        RECT 38.980 351.600 42.930 351.800 ;
        RECT 38.980 351.000 39.330 351.600 ;
        RECT 38.980 350.800 42.930 351.000 ;
        RECT 38.980 350.400 39.330 350.800 ;
        RECT 35.780 342.000 35.980 349.600 ;
        RECT 36.580 342.000 36.780 349.600 ;
        RECT 37.380 342.000 37.580 349.600 ;
        RECT 38.180 342.000 38.380 349.600 ;
        RECT 38.980 349.200 39.330 349.600 ;
        RECT 38.980 349.000 42.930 349.200 ;
        RECT 38.980 348.400 39.330 349.000 ;
        RECT 38.980 348.200 42.930 348.400 ;
        RECT 38.980 347.600 39.330 348.200 ;
        RECT 38.980 347.400 42.930 347.600 ;
        RECT 38.980 346.800 39.330 347.400 ;
        RECT 38.980 346.600 42.930 346.800 ;
        RECT 43.930 346.750 44.330 353.250 ;
        RECT 45.130 346.750 45.530 353.250 ;
        RECT 46.530 353.200 50.480 353.400 ;
        RECT 50.130 352.600 50.480 353.200 ;
        RECT 46.530 352.400 50.480 352.600 ;
        RECT 50.130 351.800 50.480 352.400 ;
        RECT 46.530 351.600 50.480 351.800 ;
        RECT 50.130 351.000 50.480 351.600 ;
        RECT 46.530 350.800 50.480 351.000 ;
        RECT 50.130 350.400 50.480 350.800 ;
        RECT 51.080 350.400 51.280 358.000 ;
        RECT 51.880 350.400 52.080 358.000 ;
        RECT 52.680 350.400 52.880 358.000 ;
        RECT 53.480 350.400 53.680 358.000 ;
        RECT 50.130 349.200 50.480 349.600 ;
        RECT 46.530 349.000 50.480 349.200 ;
        RECT 50.130 348.400 50.480 349.000 ;
        RECT 46.530 348.200 50.480 348.400 ;
        RECT 50.130 347.600 50.480 348.200 ;
        RECT 46.530 347.400 50.480 347.600 ;
        RECT 50.130 346.800 50.480 347.400 ;
        RECT 38.980 346.000 39.330 346.600 ;
        RECT 38.980 345.800 42.930 346.000 ;
        RECT 38.980 345.200 39.330 345.800 ;
        RECT 38.980 345.000 42.930 345.200 ;
        RECT 38.980 344.400 39.330 345.000 ;
        RECT 43.880 344.450 45.580 346.750 ;
        RECT 46.530 346.600 50.480 346.800 ;
        RECT 50.130 346.000 50.480 346.600 ;
        RECT 46.530 345.800 50.480 346.000 ;
        RECT 50.130 345.200 50.480 345.800 ;
        RECT 46.530 345.000 50.480 345.200 ;
        RECT 38.980 344.200 42.930 344.400 ;
        RECT 38.980 343.600 39.330 344.200 ;
        RECT 38.980 343.400 42.930 343.600 ;
        RECT 38.980 342.800 39.330 343.400 ;
        RECT 38.980 342.600 42.930 342.800 ;
        RECT 38.980 342.000 39.330 342.600 ;
        RECT 26.530 341.400 42.930 342.000 ;
        RECT 29.180 340.800 31.480 340.850 ;
        RECT 37.980 340.800 40.280 340.850 ;
        RECT 43.930 340.800 44.330 344.450 ;
        RECT 25.130 340.400 44.330 340.800 ;
        RECT 45.130 340.800 45.530 344.450 ;
        RECT 50.130 344.400 50.480 345.000 ;
        RECT 46.530 344.200 50.480 344.400 ;
        RECT 50.130 343.600 50.480 344.200 ;
        RECT 46.530 343.400 50.480 343.600 ;
        RECT 50.130 342.800 50.480 343.400 ;
        RECT 46.530 342.600 50.480 342.800 ;
        RECT 50.130 342.000 50.480 342.600 ;
        RECT 51.080 342.000 51.280 349.600 ;
        RECT 51.880 342.000 52.080 349.600 ;
        RECT 52.680 342.000 52.880 349.600 ;
        RECT 53.480 342.000 53.680 349.600 ;
        RECT 54.280 342.000 55.180 358.000 ;
        RECT 55.780 350.400 55.980 358.000 ;
        RECT 56.580 350.400 56.780 358.000 ;
        RECT 57.380 350.400 57.580 358.000 ;
        RECT 58.180 350.400 58.380 358.000 ;
        RECT 58.980 357.400 59.330 358.000 ;
        RECT 58.980 357.200 62.930 357.400 ;
        RECT 58.980 356.600 59.330 357.200 ;
        RECT 58.980 356.400 62.930 356.600 ;
        RECT 58.980 355.800 59.330 356.400 ;
        RECT 58.980 355.600 62.930 355.800 ;
        RECT 58.980 355.000 59.330 355.600 ;
        RECT 63.930 355.550 64.330 359.200 ;
        RECT 65.130 359.200 84.330 359.600 ;
        RECT 65.130 355.550 65.530 359.200 ;
        RECT 69.180 359.150 71.480 359.200 ;
        RECT 77.980 359.150 80.280 359.200 ;
        RECT 66.530 358.000 82.930 358.600 ;
        RECT 70.130 357.400 70.480 358.000 ;
        RECT 66.530 357.200 70.480 357.400 ;
        RECT 70.130 356.600 70.480 357.200 ;
        RECT 66.530 356.400 70.480 356.600 ;
        RECT 70.130 355.800 70.480 356.400 ;
        RECT 66.530 355.600 70.480 355.800 ;
        RECT 58.980 354.800 62.930 355.000 ;
        RECT 58.980 354.200 59.330 354.800 ;
        RECT 58.980 354.000 62.930 354.200 ;
        RECT 58.980 353.400 59.330 354.000 ;
        RECT 58.980 353.200 62.930 353.400 ;
        RECT 63.880 353.250 65.580 355.550 ;
        RECT 70.130 355.000 70.480 355.600 ;
        RECT 66.530 354.800 70.480 355.000 ;
        RECT 70.130 354.200 70.480 354.800 ;
        RECT 66.530 354.000 70.480 354.200 ;
        RECT 70.130 353.400 70.480 354.000 ;
        RECT 58.980 352.600 59.330 353.200 ;
        RECT 58.980 352.400 62.930 352.600 ;
        RECT 58.980 351.800 59.330 352.400 ;
        RECT 58.980 351.600 62.930 351.800 ;
        RECT 58.980 351.000 59.330 351.600 ;
        RECT 58.980 350.800 62.930 351.000 ;
        RECT 58.980 350.400 59.330 350.800 ;
        RECT 55.780 342.000 55.980 349.600 ;
        RECT 56.580 342.000 56.780 349.600 ;
        RECT 57.380 342.000 57.580 349.600 ;
        RECT 58.180 342.000 58.380 349.600 ;
        RECT 58.980 349.200 59.330 349.600 ;
        RECT 58.980 349.000 62.930 349.200 ;
        RECT 58.980 348.400 59.330 349.000 ;
        RECT 58.980 348.200 62.930 348.400 ;
        RECT 58.980 347.600 59.330 348.200 ;
        RECT 58.980 347.400 62.930 347.600 ;
        RECT 58.980 346.800 59.330 347.400 ;
        RECT 58.980 346.600 62.930 346.800 ;
        RECT 63.930 346.750 64.330 353.250 ;
        RECT 65.130 346.750 65.530 353.250 ;
        RECT 66.530 353.200 70.480 353.400 ;
        RECT 70.130 352.600 70.480 353.200 ;
        RECT 66.530 352.400 70.480 352.600 ;
        RECT 70.130 351.800 70.480 352.400 ;
        RECT 66.530 351.600 70.480 351.800 ;
        RECT 70.130 351.000 70.480 351.600 ;
        RECT 66.530 350.800 70.480 351.000 ;
        RECT 70.130 350.400 70.480 350.800 ;
        RECT 71.080 350.400 71.280 358.000 ;
        RECT 71.880 350.400 72.080 358.000 ;
        RECT 72.680 350.400 72.880 358.000 ;
        RECT 73.480 350.400 73.680 358.000 ;
        RECT 70.130 349.200 70.480 349.600 ;
        RECT 66.530 349.000 70.480 349.200 ;
        RECT 70.130 348.400 70.480 349.000 ;
        RECT 66.530 348.200 70.480 348.400 ;
        RECT 70.130 347.600 70.480 348.200 ;
        RECT 66.530 347.400 70.480 347.600 ;
        RECT 70.130 346.800 70.480 347.400 ;
        RECT 58.980 346.000 59.330 346.600 ;
        RECT 58.980 345.800 62.930 346.000 ;
        RECT 58.980 345.200 59.330 345.800 ;
        RECT 58.980 345.000 62.930 345.200 ;
        RECT 58.980 344.400 59.330 345.000 ;
        RECT 63.880 344.450 65.580 346.750 ;
        RECT 66.530 346.600 70.480 346.800 ;
        RECT 70.130 346.000 70.480 346.600 ;
        RECT 66.530 345.800 70.480 346.000 ;
        RECT 70.130 345.200 70.480 345.800 ;
        RECT 66.530 345.000 70.480 345.200 ;
        RECT 58.980 344.200 62.930 344.400 ;
        RECT 58.980 343.600 59.330 344.200 ;
        RECT 58.980 343.400 62.930 343.600 ;
        RECT 58.980 342.800 59.330 343.400 ;
        RECT 58.980 342.600 62.930 342.800 ;
        RECT 58.980 342.000 59.330 342.600 ;
        RECT 46.530 341.400 62.930 342.000 ;
        RECT 49.180 340.800 51.480 340.850 ;
        RECT 57.980 340.800 60.280 340.850 ;
        RECT 63.930 340.800 64.330 344.450 ;
        RECT 45.130 340.400 64.330 340.800 ;
        RECT 65.130 340.800 65.530 344.450 ;
        RECT 70.130 344.400 70.480 345.000 ;
        RECT 66.530 344.200 70.480 344.400 ;
        RECT 70.130 343.600 70.480 344.200 ;
        RECT 66.530 343.400 70.480 343.600 ;
        RECT 70.130 342.800 70.480 343.400 ;
        RECT 66.530 342.600 70.480 342.800 ;
        RECT 70.130 342.000 70.480 342.600 ;
        RECT 71.080 342.000 71.280 349.600 ;
        RECT 71.880 342.000 72.080 349.600 ;
        RECT 72.680 342.000 72.880 349.600 ;
        RECT 73.480 342.000 73.680 349.600 ;
        RECT 74.280 342.000 75.180 358.000 ;
        RECT 75.780 350.400 75.980 358.000 ;
        RECT 76.580 350.400 76.780 358.000 ;
        RECT 77.380 350.400 77.580 358.000 ;
        RECT 78.180 350.400 78.380 358.000 ;
        RECT 78.980 357.400 79.330 358.000 ;
        RECT 78.980 357.200 82.930 357.400 ;
        RECT 78.980 356.600 79.330 357.200 ;
        RECT 78.980 356.400 82.930 356.600 ;
        RECT 78.980 355.800 79.330 356.400 ;
        RECT 78.980 355.600 82.930 355.800 ;
        RECT 78.980 355.000 79.330 355.600 ;
        RECT 83.930 355.550 84.330 359.200 ;
        RECT 85.130 359.200 104.330 359.600 ;
        RECT 85.130 355.550 85.530 359.200 ;
        RECT 89.180 359.150 91.480 359.200 ;
        RECT 97.980 359.150 100.280 359.200 ;
        RECT 86.530 358.000 102.930 358.600 ;
        RECT 90.130 357.400 90.480 358.000 ;
        RECT 86.530 357.200 90.480 357.400 ;
        RECT 90.130 356.600 90.480 357.200 ;
        RECT 86.530 356.400 90.480 356.600 ;
        RECT 90.130 355.800 90.480 356.400 ;
        RECT 86.530 355.600 90.480 355.800 ;
        RECT 78.980 354.800 82.930 355.000 ;
        RECT 78.980 354.200 79.330 354.800 ;
        RECT 78.980 354.000 82.930 354.200 ;
        RECT 78.980 353.400 79.330 354.000 ;
        RECT 78.980 353.200 82.930 353.400 ;
        RECT 83.880 353.250 85.580 355.550 ;
        RECT 90.130 355.000 90.480 355.600 ;
        RECT 86.530 354.800 90.480 355.000 ;
        RECT 90.130 354.200 90.480 354.800 ;
        RECT 86.530 354.000 90.480 354.200 ;
        RECT 90.130 353.400 90.480 354.000 ;
        RECT 78.980 352.600 79.330 353.200 ;
        RECT 78.980 352.400 82.930 352.600 ;
        RECT 78.980 351.800 79.330 352.400 ;
        RECT 78.980 351.600 82.930 351.800 ;
        RECT 78.980 351.000 79.330 351.600 ;
        RECT 78.980 350.800 82.930 351.000 ;
        RECT 78.980 350.400 79.330 350.800 ;
        RECT 75.780 342.000 75.980 349.600 ;
        RECT 76.580 342.000 76.780 349.600 ;
        RECT 77.380 342.000 77.580 349.600 ;
        RECT 78.180 342.000 78.380 349.600 ;
        RECT 78.980 349.200 79.330 349.600 ;
        RECT 78.980 349.000 82.930 349.200 ;
        RECT 78.980 348.400 79.330 349.000 ;
        RECT 78.980 348.200 82.930 348.400 ;
        RECT 78.980 347.600 79.330 348.200 ;
        RECT 78.980 347.400 82.930 347.600 ;
        RECT 78.980 346.800 79.330 347.400 ;
        RECT 78.980 346.600 82.930 346.800 ;
        RECT 83.930 346.750 84.330 353.250 ;
        RECT 85.130 346.750 85.530 353.250 ;
        RECT 86.530 353.200 90.480 353.400 ;
        RECT 90.130 352.600 90.480 353.200 ;
        RECT 86.530 352.400 90.480 352.600 ;
        RECT 90.130 351.800 90.480 352.400 ;
        RECT 86.530 351.600 90.480 351.800 ;
        RECT 90.130 351.000 90.480 351.600 ;
        RECT 86.530 350.800 90.480 351.000 ;
        RECT 90.130 350.400 90.480 350.800 ;
        RECT 91.080 350.400 91.280 358.000 ;
        RECT 91.880 350.400 92.080 358.000 ;
        RECT 92.680 350.400 92.880 358.000 ;
        RECT 93.480 350.400 93.680 358.000 ;
        RECT 90.130 349.200 90.480 349.600 ;
        RECT 86.530 349.000 90.480 349.200 ;
        RECT 90.130 348.400 90.480 349.000 ;
        RECT 86.530 348.200 90.480 348.400 ;
        RECT 90.130 347.600 90.480 348.200 ;
        RECT 86.530 347.400 90.480 347.600 ;
        RECT 90.130 346.800 90.480 347.400 ;
        RECT 78.980 346.000 79.330 346.600 ;
        RECT 78.980 345.800 82.930 346.000 ;
        RECT 78.980 345.200 79.330 345.800 ;
        RECT 78.980 345.000 82.930 345.200 ;
        RECT 78.980 344.400 79.330 345.000 ;
        RECT 83.880 344.450 85.580 346.750 ;
        RECT 86.530 346.600 90.480 346.800 ;
        RECT 90.130 346.000 90.480 346.600 ;
        RECT 86.530 345.800 90.480 346.000 ;
        RECT 90.130 345.200 90.480 345.800 ;
        RECT 86.530 345.000 90.480 345.200 ;
        RECT 78.980 344.200 82.930 344.400 ;
        RECT 78.980 343.600 79.330 344.200 ;
        RECT 78.980 343.400 82.930 343.600 ;
        RECT 78.980 342.800 79.330 343.400 ;
        RECT 78.980 342.600 82.930 342.800 ;
        RECT 78.980 342.000 79.330 342.600 ;
        RECT 66.530 341.400 82.930 342.000 ;
        RECT 69.180 340.800 71.480 340.850 ;
        RECT 77.980 340.800 80.280 340.850 ;
        RECT 83.930 340.800 84.330 344.450 ;
        RECT 65.130 340.400 84.330 340.800 ;
        RECT 85.130 340.800 85.530 344.450 ;
        RECT 90.130 344.400 90.480 345.000 ;
        RECT 86.530 344.200 90.480 344.400 ;
        RECT 90.130 343.600 90.480 344.200 ;
        RECT 86.530 343.400 90.480 343.600 ;
        RECT 90.130 342.800 90.480 343.400 ;
        RECT 86.530 342.600 90.480 342.800 ;
        RECT 90.130 342.000 90.480 342.600 ;
        RECT 91.080 342.000 91.280 349.600 ;
        RECT 91.880 342.000 92.080 349.600 ;
        RECT 92.680 342.000 92.880 349.600 ;
        RECT 93.480 342.000 93.680 349.600 ;
        RECT 94.280 342.000 95.180 358.000 ;
        RECT 95.780 350.400 95.980 358.000 ;
        RECT 96.580 350.400 96.780 358.000 ;
        RECT 97.380 350.400 97.580 358.000 ;
        RECT 98.180 350.400 98.380 358.000 ;
        RECT 98.980 357.400 99.330 358.000 ;
        RECT 98.980 357.200 102.930 357.400 ;
        RECT 98.980 356.600 99.330 357.200 ;
        RECT 98.980 356.400 102.930 356.600 ;
        RECT 98.980 355.800 99.330 356.400 ;
        RECT 98.980 355.600 102.930 355.800 ;
        RECT 98.980 355.000 99.330 355.600 ;
        RECT 103.930 355.550 104.330 359.200 ;
        RECT 105.340 357.080 105.700 357.460 ;
        RECT 105.970 357.080 106.330 357.460 ;
        RECT 106.570 357.080 106.930 357.460 ;
        RECT 105.340 356.490 105.700 356.870 ;
        RECT 105.970 356.490 106.330 356.870 ;
        RECT 106.570 356.490 106.930 356.870 ;
        RECT 98.980 354.800 102.930 355.000 ;
        RECT 98.980 354.200 99.330 354.800 ;
        RECT 98.980 354.000 102.930 354.200 ;
        RECT 98.980 353.400 99.330 354.000 ;
        RECT 98.980 353.200 102.930 353.400 ;
        RECT 103.880 353.250 104.730 355.550 ;
        RECT 98.980 352.600 99.330 353.200 ;
        RECT 98.980 352.400 102.930 352.600 ;
        RECT 98.980 351.800 99.330 352.400 ;
        RECT 98.980 351.600 102.930 351.800 ;
        RECT 98.980 351.000 99.330 351.600 ;
        RECT 98.980 350.800 102.930 351.000 ;
        RECT 98.980 350.400 99.330 350.800 ;
        RECT 95.780 342.000 95.980 349.600 ;
        RECT 96.580 342.000 96.780 349.600 ;
        RECT 97.380 342.000 97.580 349.600 ;
        RECT 98.180 342.000 98.380 349.600 ;
        RECT 98.980 349.200 99.330 349.600 ;
        RECT 98.980 349.000 102.930 349.200 ;
        RECT 98.980 348.400 99.330 349.000 ;
        RECT 98.980 348.200 102.930 348.400 ;
        RECT 98.980 347.600 99.330 348.200 ;
        RECT 98.980 347.400 102.930 347.600 ;
        RECT 98.980 346.800 99.330 347.400 ;
        RECT 98.980 346.600 102.930 346.800 ;
        RECT 103.930 346.750 104.330 353.250 ;
        RECT 98.980 346.000 99.330 346.600 ;
        RECT 98.980 345.800 102.930 346.000 ;
        RECT 98.980 345.200 99.330 345.800 ;
        RECT 98.980 345.000 102.930 345.200 ;
        RECT 98.980 344.400 99.330 345.000 ;
        RECT 103.880 344.450 104.730 346.750 ;
        RECT 98.980 344.200 102.930 344.400 ;
        RECT 98.980 343.600 99.330 344.200 ;
        RECT 98.980 343.400 102.930 343.600 ;
        RECT 98.980 342.800 99.330 343.400 ;
        RECT 98.980 342.600 102.930 342.800 ;
        RECT 98.980 342.000 99.330 342.600 ;
        RECT 86.530 341.400 102.930 342.000 ;
        RECT 89.180 340.800 91.480 340.850 ;
        RECT 97.980 340.800 100.280 340.850 ;
        RECT 103.930 340.800 104.330 344.450 ;
        RECT 105.340 343.095 105.700 343.475 ;
        RECT 105.970 343.095 106.330 343.475 ;
        RECT 106.570 343.095 106.930 343.475 ;
        RECT 105.340 342.505 105.700 342.885 ;
        RECT 105.970 342.505 106.330 342.885 ;
        RECT 106.570 342.505 106.930 342.885 ;
        RECT 85.130 340.400 104.330 340.800 ;
        RECT 9.180 339.600 11.480 340.400 ;
        RECT 17.980 339.600 20.280 340.400 ;
        RECT 29.180 339.600 31.480 340.400 ;
        RECT 37.980 339.600 40.280 340.400 ;
        RECT 49.180 339.600 51.480 340.400 ;
        RECT 57.980 339.600 60.280 340.400 ;
        RECT 69.180 339.600 71.480 340.400 ;
        RECT 77.980 339.600 80.280 340.400 ;
        RECT 89.180 339.600 91.480 340.400 ;
        RECT 97.980 339.600 100.280 340.400 ;
        RECT 5.130 339.200 24.330 339.600 ;
        RECT 2.515 336.870 2.875 337.250 ;
        RECT 3.145 336.870 3.505 337.250 ;
        RECT 3.745 336.870 4.105 337.250 ;
        RECT 2.515 336.280 2.875 336.660 ;
        RECT 3.145 336.280 3.505 336.660 ;
        RECT 3.745 336.280 4.105 336.660 ;
        RECT 5.130 335.550 5.530 339.200 ;
        RECT 9.180 339.150 11.480 339.200 ;
        RECT 17.980 339.150 20.280 339.200 ;
        RECT 6.530 338.000 22.930 338.600 ;
        RECT 10.130 337.400 10.480 338.000 ;
        RECT 6.530 337.200 10.480 337.400 ;
        RECT 10.130 336.600 10.480 337.200 ;
        RECT 6.530 336.400 10.480 336.600 ;
        RECT 10.130 335.800 10.480 336.400 ;
        RECT 6.530 335.600 10.480 335.800 ;
        RECT 4.730 335.545 5.580 335.550 ;
        RECT 2.315 333.250 5.580 335.545 ;
        RECT 10.130 335.000 10.480 335.600 ;
        RECT 6.530 334.800 10.480 335.000 ;
        RECT 10.130 334.200 10.480 334.800 ;
        RECT 6.530 334.000 10.480 334.200 ;
        RECT 10.130 333.400 10.480 334.000 ;
        RECT 5.130 326.750 5.530 333.250 ;
        RECT 6.530 333.200 10.480 333.400 ;
        RECT 10.130 332.600 10.480 333.200 ;
        RECT 6.530 332.400 10.480 332.600 ;
        RECT 10.130 331.800 10.480 332.400 ;
        RECT 6.530 331.600 10.480 331.800 ;
        RECT 10.130 331.000 10.480 331.600 ;
        RECT 6.530 330.800 10.480 331.000 ;
        RECT 10.130 330.400 10.480 330.800 ;
        RECT 11.080 330.400 11.280 338.000 ;
        RECT 11.880 330.400 12.080 338.000 ;
        RECT 12.680 330.400 12.880 338.000 ;
        RECT 13.480 330.400 13.680 338.000 ;
        RECT 10.130 329.200 10.480 329.600 ;
        RECT 6.530 329.000 10.480 329.200 ;
        RECT 10.130 328.400 10.480 329.000 ;
        RECT 6.530 328.200 10.480 328.400 ;
        RECT 10.130 327.600 10.480 328.200 ;
        RECT 6.530 327.400 10.480 327.600 ;
        RECT 10.130 326.800 10.480 327.400 ;
        RECT 2.315 324.455 5.580 326.750 ;
        RECT 6.530 326.600 10.480 326.800 ;
        RECT 10.130 326.000 10.480 326.600 ;
        RECT 6.530 325.800 10.480 326.000 ;
        RECT 10.130 325.200 10.480 325.800 ;
        RECT 6.530 325.000 10.480 325.200 ;
        RECT 4.730 324.450 5.580 324.455 ;
        RECT 2.515 323.170 2.875 323.550 ;
        RECT 3.145 323.170 3.505 323.550 ;
        RECT 3.745 323.170 4.105 323.550 ;
        RECT 2.515 322.580 2.875 322.960 ;
        RECT 3.145 322.580 3.505 322.960 ;
        RECT 3.745 322.580 4.105 322.960 ;
        RECT 5.130 320.800 5.530 324.450 ;
        RECT 10.130 324.400 10.480 325.000 ;
        RECT 6.530 324.200 10.480 324.400 ;
        RECT 10.130 323.600 10.480 324.200 ;
        RECT 6.530 323.400 10.480 323.600 ;
        RECT 10.130 322.800 10.480 323.400 ;
        RECT 6.530 322.600 10.480 322.800 ;
        RECT 10.130 322.000 10.480 322.600 ;
        RECT 11.080 322.000 11.280 329.600 ;
        RECT 11.880 322.000 12.080 329.600 ;
        RECT 12.680 322.000 12.880 329.600 ;
        RECT 13.480 322.000 13.680 329.600 ;
        RECT 14.280 322.000 15.180 338.000 ;
        RECT 15.780 330.400 15.980 338.000 ;
        RECT 16.580 330.400 16.780 338.000 ;
        RECT 17.380 330.400 17.580 338.000 ;
        RECT 18.180 330.400 18.380 338.000 ;
        RECT 18.980 337.400 19.330 338.000 ;
        RECT 18.980 337.200 22.930 337.400 ;
        RECT 18.980 336.600 19.330 337.200 ;
        RECT 18.980 336.400 22.930 336.600 ;
        RECT 18.980 335.800 19.330 336.400 ;
        RECT 18.980 335.600 22.930 335.800 ;
        RECT 18.980 335.000 19.330 335.600 ;
        RECT 23.930 335.550 24.330 339.200 ;
        RECT 25.130 339.200 44.330 339.600 ;
        RECT 25.130 335.550 25.530 339.200 ;
        RECT 29.180 339.150 31.480 339.200 ;
        RECT 37.980 339.150 40.280 339.200 ;
        RECT 26.530 338.000 42.930 338.600 ;
        RECT 30.130 337.400 30.480 338.000 ;
        RECT 26.530 337.200 30.480 337.400 ;
        RECT 30.130 336.600 30.480 337.200 ;
        RECT 26.530 336.400 30.480 336.600 ;
        RECT 30.130 335.800 30.480 336.400 ;
        RECT 26.530 335.600 30.480 335.800 ;
        RECT 18.980 334.800 22.930 335.000 ;
        RECT 18.980 334.200 19.330 334.800 ;
        RECT 18.980 334.000 22.930 334.200 ;
        RECT 18.980 333.400 19.330 334.000 ;
        RECT 18.980 333.200 22.930 333.400 ;
        RECT 23.880 333.250 25.580 335.550 ;
        RECT 30.130 335.000 30.480 335.600 ;
        RECT 26.530 334.800 30.480 335.000 ;
        RECT 30.130 334.200 30.480 334.800 ;
        RECT 26.530 334.000 30.480 334.200 ;
        RECT 30.130 333.400 30.480 334.000 ;
        RECT 18.980 332.600 19.330 333.200 ;
        RECT 18.980 332.400 22.930 332.600 ;
        RECT 18.980 331.800 19.330 332.400 ;
        RECT 18.980 331.600 22.930 331.800 ;
        RECT 18.980 331.000 19.330 331.600 ;
        RECT 18.980 330.800 22.930 331.000 ;
        RECT 18.980 330.400 19.330 330.800 ;
        RECT 15.780 322.000 15.980 329.600 ;
        RECT 16.580 322.000 16.780 329.600 ;
        RECT 17.380 322.000 17.580 329.600 ;
        RECT 18.180 322.000 18.380 329.600 ;
        RECT 18.980 329.200 19.330 329.600 ;
        RECT 18.980 329.000 22.930 329.200 ;
        RECT 18.980 328.400 19.330 329.000 ;
        RECT 18.980 328.200 22.930 328.400 ;
        RECT 18.980 327.600 19.330 328.200 ;
        RECT 18.980 327.400 22.930 327.600 ;
        RECT 18.980 326.800 19.330 327.400 ;
        RECT 18.980 326.600 22.930 326.800 ;
        RECT 23.930 326.750 24.330 333.250 ;
        RECT 25.130 326.750 25.530 333.250 ;
        RECT 26.530 333.200 30.480 333.400 ;
        RECT 30.130 332.600 30.480 333.200 ;
        RECT 26.530 332.400 30.480 332.600 ;
        RECT 30.130 331.800 30.480 332.400 ;
        RECT 26.530 331.600 30.480 331.800 ;
        RECT 30.130 331.000 30.480 331.600 ;
        RECT 26.530 330.800 30.480 331.000 ;
        RECT 30.130 330.400 30.480 330.800 ;
        RECT 31.080 330.400 31.280 338.000 ;
        RECT 31.880 330.400 32.080 338.000 ;
        RECT 32.680 330.400 32.880 338.000 ;
        RECT 33.480 330.400 33.680 338.000 ;
        RECT 30.130 329.200 30.480 329.600 ;
        RECT 26.530 329.000 30.480 329.200 ;
        RECT 30.130 328.400 30.480 329.000 ;
        RECT 26.530 328.200 30.480 328.400 ;
        RECT 30.130 327.600 30.480 328.200 ;
        RECT 26.530 327.400 30.480 327.600 ;
        RECT 30.130 326.800 30.480 327.400 ;
        RECT 18.980 326.000 19.330 326.600 ;
        RECT 18.980 325.800 22.930 326.000 ;
        RECT 18.980 325.200 19.330 325.800 ;
        RECT 18.980 325.000 22.930 325.200 ;
        RECT 18.980 324.400 19.330 325.000 ;
        RECT 23.880 324.450 25.580 326.750 ;
        RECT 26.530 326.600 30.480 326.800 ;
        RECT 30.130 326.000 30.480 326.600 ;
        RECT 26.530 325.800 30.480 326.000 ;
        RECT 30.130 325.200 30.480 325.800 ;
        RECT 26.530 325.000 30.480 325.200 ;
        RECT 18.980 324.200 22.930 324.400 ;
        RECT 18.980 323.600 19.330 324.200 ;
        RECT 18.980 323.400 22.930 323.600 ;
        RECT 18.980 322.800 19.330 323.400 ;
        RECT 18.980 322.600 22.930 322.800 ;
        RECT 18.980 322.000 19.330 322.600 ;
        RECT 6.530 321.400 22.930 322.000 ;
        RECT 9.180 320.800 11.480 320.850 ;
        RECT 17.980 320.800 20.280 320.850 ;
        RECT 23.930 320.800 24.330 324.450 ;
        RECT 5.130 320.400 24.330 320.800 ;
        RECT 25.130 320.800 25.530 324.450 ;
        RECT 30.130 324.400 30.480 325.000 ;
        RECT 26.530 324.200 30.480 324.400 ;
        RECT 30.130 323.600 30.480 324.200 ;
        RECT 26.530 323.400 30.480 323.600 ;
        RECT 30.130 322.800 30.480 323.400 ;
        RECT 26.530 322.600 30.480 322.800 ;
        RECT 30.130 322.000 30.480 322.600 ;
        RECT 31.080 322.000 31.280 329.600 ;
        RECT 31.880 322.000 32.080 329.600 ;
        RECT 32.680 322.000 32.880 329.600 ;
        RECT 33.480 322.000 33.680 329.600 ;
        RECT 34.280 322.000 35.180 338.000 ;
        RECT 35.780 330.400 35.980 338.000 ;
        RECT 36.580 330.400 36.780 338.000 ;
        RECT 37.380 330.400 37.580 338.000 ;
        RECT 38.180 330.400 38.380 338.000 ;
        RECT 38.980 337.400 39.330 338.000 ;
        RECT 38.980 337.200 42.930 337.400 ;
        RECT 38.980 336.600 39.330 337.200 ;
        RECT 38.980 336.400 42.930 336.600 ;
        RECT 38.980 335.800 39.330 336.400 ;
        RECT 38.980 335.600 42.930 335.800 ;
        RECT 38.980 335.000 39.330 335.600 ;
        RECT 43.930 335.550 44.330 339.200 ;
        RECT 45.130 339.200 64.330 339.600 ;
        RECT 45.130 335.550 45.530 339.200 ;
        RECT 49.180 339.150 51.480 339.200 ;
        RECT 57.980 339.150 60.280 339.200 ;
        RECT 46.530 338.000 62.930 338.600 ;
        RECT 50.130 337.400 50.480 338.000 ;
        RECT 46.530 337.200 50.480 337.400 ;
        RECT 50.130 336.600 50.480 337.200 ;
        RECT 46.530 336.400 50.480 336.600 ;
        RECT 50.130 335.800 50.480 336.400 ;
        RECT 46.530 335.600 50.480 335.800 ;
        RECT 38.980 334.800 42.930 335.000 ;
        RECT 38.980 334.200 39.330 334.800 ;
        RECT 38.980 334.000 42.930 334.200 ;
        RECT 38.980 333.400 39.330 334.000 ;
        RECT 38.980 333.200 42.930 333.400 ;
        RECT 43.880 333.250 45.580 335.550 ;
        RECT 50.130 335.000 50.480 335.600 ;
        RECT 46.530 334.800 50.480 335.000 ;
        RECT 50.130 334.200 50.480 334.800 ;
        RECT 46.530 334.000 50.480 334.200 ;
        RECT 50.130 333.400 50.480 334.000 ;
        RECT 38.980 332.600 39.330 333.200 ;
        RECT 38.980 332.400 42.930 332.600 ;
        RECT 38.980 331.800 39.330 332.400 ;
        RECT 38.980 331.600 42.930 331.800 ;
        RECT 38.980 331.000 39.330 331.600 ;
        RECT 38.980 330.800 42.930 331.000 ;
        RECT 38.980 330.400 39.330 330.800 ;
        RECT 35.780 322.000 35.980 329.600 ;
        RECT 36.580 322.000 36.780 329.600 ;
        RECT 37.380 322.000 37.580 329.600 ;
        RECT 38.180 322.000 38.380 329.600 ;
        RECT 38.980 329.200 39.330 329.600 ;
        RECT 38.980 329.000 42.930 329.200 ;
        RECT 38.980 328.400 39.330 329.000 ;
        RECT 38.980 328.200 42.930 328.400 ;
        RECT 38.980 327.600 39.330 328.200 ;
        RECT 38.980 327.400 42.930 327.600 ;
        RECT 38.980 326.800 39.330 327.400 ;
        RECT 38.980 326.600 42.930 326.800 ;
        RECT 43.930 326.750 44.330 333.250 ;
        RECT 45.130 326.750 45.530 333.250 ;
        RECT 46.530 333.200 50.480 333.400 ;
        RECT 50.130 332.600 50.480 333.200 ;
        RECT 46.530 332.400 50.480 332.600 ;
        RECT 50.130 331.800 50.480 332.400 ;
        RECT 46.530 331.600 50.480 331.800 ;
        RECT 50.130 331.000 50.480 331.600 ;
        RECT 46.530 330.800 50.480 331.000 ;
        RECT 50.130 330.400 50.480 330.800 ;
        RECT 51.080 330.400 51.280 338.000 ;
        RECT 51.880 330.400 52.080 338.000 ;
        RECT 52.680 330.400 52.880 338.000 ;
        RECT 53.480 330.400 53.680 338.000 ;
        RECT 50.130 329.200 50.480 329.600 ;
        RECT 46.530 329.000 50.480 329.200 ;
        RECT 50.130 328.400 50.480 329.000 ;
        RECT 46.530 328.200 50.480 328.400 ;
        RECT 50.130 327.600 50.480 328.200 ;
        RECT 46.530 327.400 50.480 327.600 ;
        RECT 50.130 326.800 50.480 327.400 ;
        RECT 38.980 326.000 39.330 326.600 ;
        RECT 38.980 325.800 42.930 326.000 ;
        RECT 38.980 325.200 39.330 325.800 ;
        RECT 38.980 325.000 42.930 325.200 ;
        RECT 38.980 324.400 39.330 325.000 ;
        RECT 43.880 324.450 45.580 326.750 ;
        RECT 46.530 326.600 50.480 326.800 ;
        RECT 50.130 326.000 50.480 326.600 ;
        RECT 46.530 325.800 50.480 326.000 ;
        RECT 50.130 325.200 50.480 325.800 ;
        RECT 46.530 325.000 50.480 325.200 ;
        RECT 38.980 324.200 42.930 324.400 ;
        RECT 38.980 323.600 39.330 324.200 ;
        RECT 38.980 323.400 42.930 323.600 ;
        RECT 38.980 322.800 39.330 323.400 ;
        RECT 38.980 322.600 42.930 322.800 ;
        RECT 38.980 322.000 39.330 322.600 ;
        RECT 26.530 321.400 42.930 322.000 ;
        RECT 29.180 320.800 31.480 320.850 ;
        RECT 37.980 320.800 40.280 320.850 ;
        RECT 43.930 320.800 44.330 324.450 ;
        RECT 25.130 320.400 44.330 320.800 ;
        RECT 45.130 320.800 45.530 324.450 ;
        RECT 50.130 324.400 50.480 325.000 ;
        RECT 46.530 324.200 50.480 324.400 ;
        RECT 50.130 323.600 50.480 324.200 ;
        RECT 46.530 323.400 50.480 323.600 ;
        RECT 50.130 322.800 50.480 323.400 ;
        RECT 46.530 322.600 50.480 322.800 ;
        RECT 50.130 322.000 50.480 322.600 ;
        RECT 51.080 322.000 51.280 329.600 ;
        RECT 51.880 322.000 52.080 329.600 ;
        RECT 52.680 322.000 52.880 329.600 ;
        RECT 53.480 322.000 53.680 329.600 ;
        RECT 54.280 322.000 55.180 338.000 ;
        RECT 55.780 330.400 55.980 338.000 ;
        RECT 56.580 330.400 56.780 338.000 ;
        RECT 57.380 330.400 57.580 338.000 ;
        RECT 58.180 330.400 58.380 338.000 ;
        RECT 58.980 337.400 59.330 338.000 ;
        RECT 58.980 337.200 62.930 337.400 ;
        RECT 58.980 336.600 59.330 337.200 ;
        RECT 58.980 336.400 62.930 336.600 ;
        RECT 58.980 335.800 59.330 336.400 ;
        RECT 58.980 335.600 62.930 335.800 ;
        RECT 58.980 335.000 59.330 335.600 ;
        RECT 63.930 335.550 64.330 339.200 ;
        RECT 65.130 339.200 84.330 339.600 ;
        RECT 65.130 335.550 65.530 339.200 ;
        RECT 69.180 339.150 71.480 339.200 ;
        RECT 77.980 339.150 80.280 339.200 ;
        RECT 66.530 338.000 82.930 338.600 ;
        RECT 70.130 337.400 70.480 338.000 ;
        RECT 66.530 337.200 70.480 337.400 ;
        RECT 70.130 336.600 70.480 337.200 ;
        RECT 66.530 336.400 70.480 336.600 ;
        RECT 70.130 335.800 70.480 336.400 ;
        RECT 66.530 335.600 70.480 335.800 ;
        RECT 58.980 334.800 62.930 335.000 ;
        RECT 58.980 334.200 59.330 334.800 ;
        RECT 58.980 334.000 62.930 334.200 ;
        RECT 58.980 333.400 59.330 334.000 ;
        RECT 58.980 333.200 62.930 333.400 ;
        RECT 63.880 333.250 65.580 335.550 ;
        RECT 70.130 335.000 70.480 335.600 ;
        RECT 66.530 334.800 70.480 335.000 ;
        RECT 70.130 334.200 70.480 334.800 ;
        RECT 66.530 334.000 70.480 334.200 ;
        RECT 70.130 333.400 70.480 334.000 ;
        RECT 58.980 332.600 59.330 333.200 ;
        RECT 58.980 332.400 62.930 332.600 ;
        RECT 58.980 331.800 59.330 332.400 ;
        RECT 58.980 331.600 62.930 331.800 ;
        RECT 58.980 331.000 59.330 331.600 ;
        RECT 58.980 330.800 62.930 331.000 ;
        RECT 58.980 330.400 59.330 330.800 ;
        RECT 55.780 322.000 55.980 329.600 ;
        RECT 56.580 322.000 56.780 329.600 ;
        RECT 57.380 322.000 57.580 329.600 ;
        RECT 58.180 322.000 58.380 329.600 ;
        RECT 58.980 329.200 59.330 329.600 ;
        RECT 58.980 329.000 62.930 329.200 ;
        RECT 58.980 328.400 59.330 329.000 ;
        RECT 58.980 328.200 62.930 328.400 ;
        RECT 58.980 327.600 59.330 328.200 ;
        RECT 58.980 327.400 62.930 327.600 ;
        RECT 58.980 326.800 59.330 327.400 ;
        RECT 58.980 326.600 62.930 326.800 ;
        RECT 63.930 326.750 64.330 333.250 ;
        RECT 65.130 326.750 65.530 333.250 ;
        RECT 66.530 333.200 70.480 333.400 ;
        RECT 70.130 332.600 70.480 333.200 ;
        RECT 66.530 332.400 70.480 332.600 ;
        RECT 70.130 331.800 70.480 332.400 ;
        RECT 66.530 331.600 70.480 331.800 ;
        RECT 70.130 331.000 70.480 331.600 ;
        RECT 66.530 330.800 70.480 331.000 ;
        RECT 70.130 330.400 70.480 330.800 ;
        RECT 71.080 330.400 71.280 338.000 ;
        RECT 71.880 330.400 72.080 338.000 ;
        RECT 72.680 330.400 72.880 338.000 ;
        RECT 73.480 330.400 73.680 338.000 ;
        RECT 70.130 329.200 70.480 329.600 ;
        RECT 66.530 329.000 70.480 329.200 ;
        RECT 70.130 328.400 70.480 329.000 ;
        RECT 66.530 328.200 70.480 328.400 ;
        RECT 70.130 327.600 70.480 328.200 ;
        RECT 66.530 327.400 70.480 327.600 ;
        RECT 70.130 326.800 70.480 327.400 ;
        RECT 58.980 326.000 59.330 326.600 ;
        RECT 58.980 325.800 62.930 326.000 ;
        RECT 58.980 325.200 59.330 325.800 ;
        RECT 58.980 325.000 62.930 325.200 ;
        RECT 58.980 324.400 59.330 325.000 ;
        RECT 63.880 324.450 65.580 326.750 ;
        RECT 66.530 326.600 70.480 326.800 ;
        RECT 70.130 326.000 70.480 326.600 ;
        RECT 66.530 325.800 70.480 326.000 ;
        RECT 70.130 325.200 70.480 325.800 ;
        RECT 66.530 325.000 70.480 325.200 ;
        RECT 58.980 324.200 62.930 324.400 ;
        RECT 58.980 323.600 59.330 324.200 ;
        RECT 58.980 323.400 62.930 323.600 ;
        RECT 58.980 322.800 59.330 323.400 ;
        RECT 58.980 322.600 62.930 322.800 ;
        RECT 58.980 322.000 59.330 322.600 ;
        RECT 46.530 321.400 62.930 322.000 ;
        RECT 49.180 320.800 51.480 320.850 ;
        RECT 57.980 320.800 60.280 320.850 ;
        RECT 63.930 320.800 64.330 324.450 ;
        RECT 45.130 320.400 64.330 320.800 ;
        RECT 65.130 320.800 65.530 324.450 ;
        RECT 70.130 324.400 70.480 325.000 ;
        RECT 66.530 324.200 70.480 324.400 ;
        RECT 70.130 323.600 70.480 324.200 ;
        RECT 66.530 323.400 70.480 323.600 ;
        RECT 70.130 322.800 70.480 323.400 ;
        RECT 66.530 322.600 70.480 322.800 ;
        RECT 70.130 322.000 70.480 322.600 ;
        RECT 71.080 322.000 71.280 329.600 ;
        RECT 71.880 322.000 72.080 329.600 ;
        RECT 72.680 322.000 72.880 329.600 ;
        RECT 73.480 322.000 73.680 329.600 ;
        RECT 74.280 322.000 75.180 338.000 ;
        RECT 75.780 330.400 75.980 338.000 ;
        RECT 76.580 330.400 76.780 338.000 ;
        RECT 77.380 330.400 77.580 338.000 ;
        RECT 78.180 330.400 78.380 338.000 ;
        RECT 78.980 337.400 79.330 338.000 ;
        RECT 78.980 337.200 82.930 337.400 ;
        RECT 78.980 336.600 79.330 337.200 ;
        RECT 78.980 336.400 82.930 336.600 ;
        RECT 78.980 335.800 79.330 336.400 ;
        RECT 78.980 335.600 82.930 335.800 ;
        RECT 78.980 335.000 79.330 335.600 ;
        RECT 83.930 335.550 84.330 339.200 ;
        RECT 85.130 339.200 104.330 339.600 ;
        RECT 85.130 335.550 85.530 339.200 ;
        RECT 89.180 339.150 91.480 339.200 ;
        RECT 97.980 339.150 100.280 339.200 ;
        RECT 86.530 338.000 102.930 338.600 ;
        RECT 90.130 337.400 90.480 338.000 ;
        RECT 86.530 337.200 90.480 337.400 ;
        RECT 90.130 336.600 90.480 337.200 ;
        RECT 86.530 336.400 90.480 336.600 ;
        RECT 90.130 335.800 90.480 336.400 ;
        RECT 86.530 335.600 90.480 335.800 ;
        RECT 78.980 334.800 82.930 335.000 ;
        RECT 78.980 334.200 79.330 334.800 ;
        RECT 78.980 334.000 82.930 334.200 ;
        RECT 78.980 333.400 79.330 334.000 ;
        RECT 78.980 333.200 82.930 333.400 ;
        RECT 83.880 333.250 85.580 335.550 ;
        RECT 90.130 335.000 90.480 335.600 ;
        RECT 86.530 334.800 90.480 335.000 ;
        RECT 90.130 334.200 90.480 334.800 ;
        RECT 86.530 334.000 90.480 334.200 ;
        RECT 90.130 333.400 90.480 334.000 ;
        RECT 78.980 332.600 79.330 333.200 ;
        RECT 78.980 332.400 82.930 332.600 ;
        RECT 78.980 331.800 79.330 332.400 ;
        RECT 78.980 331.600 82.930 331.800 ;
        RECT 78.980 331.000 79.330 331.600 ;
        RECT 78.980 330.800 82.930 331.000 ;
        RECT 78.980 330.400 79.330 330.800 ;
        RECT 75.780 322.000 75.980 329.600 ;
        RECT 76.580 322.000 76.780 329.600 ;
        RECT 77.380 322.000 77.580 329.600 ;
        RECT 78.180 322.000 78.380 329.600 ;
        RECT 78.980 329.200 79.330 329.600 ;
        RECT 78.980 329.000 82.930 329.200 ;
        RECT 78.980 328.400 79.330 329.000 ;
        RECT 78.980 328.200 82.930 328.400 ;
        RECT 78.980 327.600 79.330 328.200 ;
        RECT 78.980 327.400 82.930 327.600 ;
        RECT 78.980 326.800 79.330 327.400 ;
        RECT 78.980 326.600 82.930 326.800 ;
        RECT 83.930 326.750 84.330 333.250 ;
        RECT 85.130 326.750 85.530 333.250 ;
        RECT 86.530 333.200 90.480 333.400 ;
        RECT 90.130 332.600 90.480 333.200 ;
        RECT 86.530 332.400 90.480 332.600 ;
        RECT 90.130 331.800 90.480 332.400 ;
        RECT 86.530 331.600 90.480 331.800 ;
        RECT 90.130 331.000 90.480 331.600 ;
        RECT 86.530 330.800 90.480 331.000 ;
        RECT 90.130 330.400 90.480 330.800 ;
        RECT 91.080 330.400 91.280 338.000 ;
        RECT 91.880 330.400 92.080 338.000 ;
        RECT 92.680 330.400 92.880 338.000 ;
        RECT 93.480 330.400 93.680 338.000 ;
        RECT 90.130 329.200 90.480 329.600 ;
        RECT 86.530 329.000 90.480 329.200 ;
        RECT 90.130 328.400 90.480 329.000 ;
        RECT 86.530 328.200 90.480 328.400 ;
        RECT 90.130 327.600 90.480 328.200 ;
        RECT 86.530 327.400 90.480 327.600 ;
        RECT 90.130 326.800 90.480 327.400 ;
        RECT 78.980 326.000 79.330 326.600 ;
        RECT 78.980 325.800 82.930 326.000 ;
        RECT 78.980 325.200 79.330 325.800 ;
        RECT 78.980 325.000 82.930 325.200 ;
        RECT 78.980 324.400 79.330 325.000 ;
        RECT 83.880 324.450 85.580 326.750 ;
        RECT 86.530 326.600 90.480 326.800 ;
        RECT 90.130 326.000 90.480 326.600 ;
        RECT 86.530 325.800 90.480 326.000 ;
        RECT 90.130 325.200 90.480 325.800 ;
        RECT 86.530 325.000 90.480 325.200 ;
        RECT 78.980 324.200 82.930 324.400 ;
        RECT 78.980 323.600 79.330 324.200 ;
        RECT 78.980 323.400 82.930 323.600 ;
        RECT 78.980 322.800 79.330 323.400 ;
        RECT 78.980 322.600 82.930 322.800 ;
        RECT 78.980 322.000 79.330 322.600 ;
        RECT 66.530 321.400 82.930 322.000 ;
        RECT 69.180 320.800 71.480 320.850 ;
        RECT 77.980 320.800 80.280 320.850 ;
        RECT 83.930 320.800 84.330 324.450 ;
        RECT 65.130 320.400 84.330 320.800 ;
        RECT 85.130 320.800 85.530 324.450 ;
        RECT 90.130 324.400 90.480 325.000 ;
        RECT 86.530 324.200 90.480 324.400 ;
        RECT 90.130 323.600 90.480 324.200 ;
        RECT 86.530 323.400 90.480 323.600 ;
        RECT 90.130 322.800 90.480 323.400 ;
        RECT 86.530 322.600 90.480 322.800 ;
        RECT 90.130 322.000 90.480 322.600 ;
        RECT 91.080 322.000 91.280 329.600 ;
        RECT 91.880 322.000 92.080 329.600 ;
        RECT 92.680 322.000 92.880 329.600 ;
        RECT 93.480 322.000 93.680 329.600 ;
        RECT 94.280 322.000 95.180 338.000 ;
        RECT 95.780 330.400 95.980 338.000 ;
        RECT 96.580 330.400 96.780 338.000 ;
        RECT 97.380 330.400 97.580 338.000 ;
        RECT 98.180 330.400 98.380 338.000 ;
        RECT 98.980 337.400 99.330 338.000 ;
        RECT 98.980 337.200 102.930 337.400 ;
        RECT 98.980 336.600 99.330 337.200 ;
        RECT 98.980 336.400 102.930 336.600 ;
        RECT 98.980 335.800 99.330 336.400 ;
        RECT 98.980 335.600 102.930 335.800 ;
        RECT 98.980 335.000 99.330 335.600 ;
        RECT 103.930 335.550 104.330 339.200 ;
        RECT 105.340 337.080 105.700 337.460 ;
        RECT 105.970 337.080 106.330 337.460 ;
        RECT 106.570 337.080 106.930 337.460 ;
        RECT 105.340 336.490 105.700 336.870 ;
        RECT 105.970 336.490 106.330 336.870 ;
        RECT 106.570 336.490 106.930 336.870 ;
        RECT 98.980 334.800 102.930 335.000 ;
        RECT 98.980 334.200 99.330 334.800 ;
        RECT 98.980 334.000 102.930 334.200 ;
        RECT 98.980 333.400 99.330 334.000 ;
        RECT 98.980 333.200 102.930 333.400 ;
        RECT 103.880 333.250 104.730 335.550 ;
        RECT 98.980 332.600 99.330 333.200 ;
        RECT 98.980 332.400 102.930 332.600 ;
        RECT 98.980 331.800 99.330 332.400 ;
        RECT 98.980 331.600 102.930 331.800 ;
        RECT 98.980 331.000 99.330 331.600 ;
        RECT 98.980 330.800 102.930 331.000 ;
        RECT 98.980 330.400 99.330 330.800 ;
        RECT 95.780 322.000 95.980 329.600 ;
        RECT 96.580 322.000 96.780 329.600 ;
        RECT 97.380 322.000 97.580 329.600 ;
        RECT 98.180 322.000 98.380 329.600 ;
        RECT 98.980 329.200 99.330 329.600 ;
        RECT 98.980 329.000 102.930 329.200 ;
        RECT 98.980 328.400 99.330 329.000 ;
        RECT 98.980 328.200 102.930 328.400 ;
        RECT 98.980 327.600 99.330 328.200 ;
        RECT 98.980 327.400 102.930 327.600 ;
        RECT 98.980 326.800 99.330 327.400 ;
        RECT 98.980 326.600 102.930 326.800 ;
        RECT 103.930 326.750 104.330 333.250 ;
        RECT 98.980 326.000 99.330 326.600 ;
        RECT 98.980 325.800 102.930 326.000 ;
        RECT 98.980 325.200 99.330 325.800 ;
        RECT 98.980 325.000 102.930 325.200 ;
        RECT 98.980 324.400 99.330 325.000 ;
        RECT 103.880 324.450 104.730 326.750 ;
        RECT 98.980 324.200 102.930 324.400 ;
        RECT 98.980 323.600 99.330 324.200 ;
        RECT 98.980 323.400 102.930 323.600 ;
        RECT 98.980 322.800 99.330 323.400 ;
        RECT 98.980 322.600 102.930 322.800 ;
        RECT 98.980 322.000 99.330 322.600 ;
        RECT 86.530 321.400 102.930 322.000 ;
        RECT 89.180 320.800 91.480 320.850 ;
        RECT 97.980 320.800 100.280 320.850 ;
        RECT 103.930 320.800 104.330 324.450 ;
        RECT 105.340 323.095 105.700 323.475 ;
        RECT 105.970 323.095 106.330 323.475 ;
        RECT 106.570 323.095 106.930 323.475 ;
        RECT 105.340 322.505 105.700 322.885 ;
        RECT 105.970 322.505 106.330 322.885 ;
        RECT 106.570 322.505 106.930 322.885 ;
        RECT 85.130 320.400 104.330 320.800 ;
        RECT 9.180 319.600 11.480 320.400 ;
        RECT 17.980 319.600 20.280 320.400 ;
        RECT 29.180 319.600 31.480 320.400 ;
        RECT 37.980 319.600 40.280 320.400 ;
        RECT 49.180 319.600 51.480 320.400 ;
        RECT 57.980 319.600 60.280 320.400 ;
        RECT 69.180 319.600 71.480 320.400 ;
        RECT 77.980 319.600 80.280 320.400 ;
        RECT 89.180 319.600 91.480 320.400 ;
        RECT 97.980 319.600 100.280 320.400 ;
        RECT 5.130 319.200 24.330 319.600 ;
        RECT 2.515 317.280 2.875 317.660 ;
        RECT 3.145 317.280 3.505 317.660 ;
        RECT 3.745 317.280 4.105 317.660 ;
        RECT 2.515 316.690 2.875 317.070 ;
        RECT 3.145 316.690 3.505 317.070 ;
        RECT 3.745 316.690 4.105 317.070 ;
        RECT 5.130 315.550 5.530 319.200 ;
        RECT 9.180 319.150 11.480 319.200 ;
        RECT 17.980 319.150 20.280 319.200 ;
        RECT 6.530 318.000 22.930 318.600 ;
        RECT 10.130 317.400 10.480 318.000 ;
        RECT 6.530 317.200 10.480 317.400 ;
        RECT 10.130 316.600 10.480 317.200 ;
        RECT 6.530 316.400 10.480 316.600 ;
        RECT 10.130 315.800 10.480 316.400 ;
        RECT 6.530 315.600 10.480 315.800 ;
        RECT 4.730 315.545 5.580 315.550 ;
        RECT 2.320 315.340 5.580 315.545 ;
        RECT 2.315 313.250 5.580 315.340 ;
        RECT 10.130 315.000 10.480 315.600 ;
        RECT 6.530 314.800 10.480 315.000 ;
        RECT 10.130 314.200 10.480 314.800 ;
        RECT 6.530 314.000 10.480 314.200 ;
        RECT 10.130 313.400 10.480 314.000 ;
        RECT 5.130 306.750 5.530 313.250 ;
        RECT 6.530 313.200 10.480 313.400 ;
        RECT 10.130 312.600 10.480 313.200 ;
        RECT 6.530 312.400 10.480 312.600 ;
        RECT 10.130 311.800 10.480 312.400 ;
        RECT 6.530 311.600 10.480 311.800 ;
        RECT 10.130 311.000 10.480 311.600 ;
        RECT 6.530 310.800 10.480 311.000 ;
        RECT 10.130 310.400 10.480 310.800 ;
        RECT 11.080 310.400 11.280 318.000 ;
        RECT 11.880 310.400 12.080 318.000 ;
        RECT 12.680 310.400 12.880 318.000 ;
        RECT 13.480 310.400 13.680 318.000 ;
        RECT 10.130 309.200 10.480 309.600 ;
        RECT 6.530 309.000 10.480 309.200 ;
        RECT 10.130 308.400 10.480 309.000 ;
        RECT 6.530 308.200 10.480 308.400 ;
        RECT 10.130 307.600 10.480 308.200 ;
        RECT 6.530 307.400 10.480 307.600 ;
        RECT 10.130 306.800 10.480 307.400 ;
        RECT 2.315 304.455 5.580 306.750 ;
        RECT 6.530 306.600 10.480 306.800 ;
        RECT 10.130 306.000 10.480 306.600 ;
        RECT 6.530 305.800 10.480 306.000 ;
        RECT 10.130 305.200 10.480 305.800 ;
        RECT 6.530 305.000 10.480 305.200 ;
        RECT 4.730 304.450 5.580 304.455 ;
        RECT 2.515 303.040 2.875 303.420 ;
        RECT 3.145 303.040 3.505 303.420 ;
        RECT 3.745 303.040 4.105 303.420 ;
        RECT 2.515 302.450 2.875 302.830 ;
        RECT 3.145 302.450 3.505 302.830 ;
        RECT 3.745 302.450 4.105 302.830 ;
        RECT 5.130 300.800 5.530 304.450 ;
        RECT 10.130 304.400 10.480 305.000 ;
        RECT 6.530 304.200 10.480 304.400 ;
        RECT 10.130 303.600 10.480 304.200 ;
        RECT 6.530 303.400 10.480 303.600 ;
        RECT 10.130 302.800 10.480 303.400 ;
        RECT 6.530 302.600 10.480 302.800 ;
        RECT 10.130 302.000 10.480 302.600 ;
        RECT 11.080 302.000 11.280 309.600 ;
        RECT 11.880 302.000 12.080 309.600 ;
        RECT 12.680 302.000 12.880 309.600 ;
        RECT 13.480 302.000 13.680 309.600 ;
        RECT 14.280 302.000 15.180 318.000 ;
        RECT 15.780 310.400 15.980 318.000 ;
        RECT 16.580 310.400 16.780 318.000 ;
        RECT 17.380 310.400 17.580 318.000 ;
        RECT 18.180 310.400 18.380 318.000 ;
        RECT 18.980 317.400 19.330 318.000 ;
        RECT 18.980 317.200 22.930 317.400 ;
        RECT 18.980 316.600 19.330 317.200 ;
        RECT 18.980 316.400 22.930 316.600 ;
        RECT 18.980 315.800 19.330 316.400 ;
        RECT 18.980 315.600 22.930 315.800 ;
        RECT 18.980 315.000 19.330 315.600 ;
        RECT 23.930 315.550 24.330 319.200 ;
        RECT 25.130 319.200 44.330 319.600 ;
        RECT 25.130 315.550 25.530 319.200 ;
        RECT 29.180 319.150 31.480 319.200 ;
        RECT 37.980 319.150 40.280 319.200 ;
        RECT 26.530 318.000 42.930 318.600 ;
        RECT 30.130 317.400 30.480 318.000 ;
        RECT 26.530 317.200 30.480 317.400 ;
        RECT 30.130 316.600 30.480 317.200 ;
        RECT 26.530 316.400 30.480 316.600 ;
        RECT 30.130 315.800 30.480 316.400 ;
        RECT 26.530 315.600 30.480 315.800 ;
        RECT 18.980 314.800 22.930 315.000 ;
        RECT 18.980 314.200 19.330 314.800 ;
        RECT 18.980 314.000 22.930 314.200 ;
        RECT 18.980 313.400 19.330 314.000 ;
        RECT 18.980 313.200 22.930 313.400 ;
        RECT 23.880 313.250 25.580 315.550 ;
        RECT 30.130 315.000 30.480 315.600 ;
        RECT 26.530 314.800 30.480 315.000 ;
        RECT 30.130 314.200 30.480 314.800 ;
        RECT 26.530 314.000 30.480 314.200 ;
        RECT 30.130 313.400 30.480 314.000 ;
        RECT 18.980 312.600 19.330 313.200 ;
        RECT 18.980 312.400 22.930 312.600 ;
        RECT 18.980 311.800 19.330 312.400 ;
        RECT 18.980 311.600 22.930 311.800 ;
        RECT 18.980 311.000 19.330 311.600 ;
        RECT 18.980 310.800 22.930 311.000 ;
        RECT 18.980 310.400 19.330 310.800 ;
        RECT 15.780 302.000 15.980 309.600 ;
        RECT 16.580 302.000 16.780 309.600 ;
        RECT 17.380 302.000 17.580 309.600 ;
        RECT 18.180 302.000 18.380 309.600 ;
        RECT 18.980 309.200 19.330 309.600 ;
        RECT 18.980 309.000 22.930 309.200 ;
        RECT 18.980 308.400 19.330 309.000 ;
        RECT 18.980 308.200 22.930 308.400 ;
        RECT 18.980 307.600 19.330 308.200 ;
        RECT 18.980 307.400 22.930 307.600 ;
        RECT 18.980 306.800 19.330 307.400 ;
        RECT 18.980 306.600 22.930 306.800 ;
        RECT 23.930 306.750 24.330 313.250 ;
        RECT 25.130 306.750 25.530 313.250 ;
        RECT 26.530 313.200 30.480 313.400 ;
        RECT 30.130 312.600 30.480 313.200 ;
        RECT 26.530 312.400 30.480 312.600 ;
        RECT 30.130 311.800 30.480 312.400 ;
        RECT 26.530 311.600 30.480 311.800 ;
        RECT 30.130 311.000 30.480 311.600 ;
        RECT 26.530 310.800 30.480 311.000 ;
        RECT 30.130 310.400 30.480 310.800 ;
        RECT 31.080 310.400 31.280 318.000 ;
        RECT 31.880 310.400 32.080 318.000 ;
        RECT 32.680 310.400 32.880 318.000 ;
        RECT 33.480 310.400 33.680 318.000 ;
        RECT 30.130 309.200 30.480 309.600 ;
        RECT 26.530 309.000 30.480 309.200 ;
        RECT 30.130 308.400 30.480 309.000 ;
        RECT 26.530 308.200 30.480 308.400 ;
        RECT 30.130 307.600 30.480 308.200 ;
        RECT 26.530 307.400 30.480 307.600 ;
        RECT 30.130 306.800 30.480 307.400 ;
        RECT 18.980 306.000 19.330 306.600 ;
        RECT 18.980 305.800 22.930 306.000 ;
        RECT 18.980 305.200 19.330 305.800 ;
        RECT 18.980 305.000 22.930 305.200 ;
        RECT 18.980 304.400 19.330 305.000 ;
        RECT 23.880 304.450 25.580 306.750 ;
        RECT 26.530 306.600 30.480 306.800 ;
        RECT 30.130 306.000 30.480 306.600 ;
        RECT 26.530 305.800 30.480 306.000 ;
        RECT 30.130 305.200 30.480 305.800 ;
        RECT 26.530 305.000 30.480 305.200 ;
        RECT 18.980 304.200 22.930 304.400 ;
        RECT 18.980 303.600 19.330 304.200 ;
        RECT 18.980 303.400 22.930 303.600 ;
        RECT 18.980 302.800 19.330 303.400 ;
        RECT 18.980 302.600 22.930 302.800 ;
        RECT 18.980 302.000 19.330 302.600 ;
        RECT 6.530 301.400 22.930 302.000 ;
        RECT 9.180 300.800 11.480 300.850 ;
        RECT 17.980 300.800 20.280 300.850 ;
        RECT 23.930 300.800 24.330 304.450 ;
        RECT 5.130 300.400 24.330 300.800 ;
        RECT 25.130 300.800 25.530 304.450 ;
        RECT 30.130 304.400 30.480 305.000 ;
        RECT 26.530 304.200 30.480 304.400 ;
        RECT 30.130 303.600 30.480 304.200 ;
        RECT 26.530 303.400 30.480 303.600 ;
        RECT 30.130 302.800 30.480 303.400 ;
        RECT 26.530 302.600 30.480 302.800 ;
        RECT 30.130 302.000 30.480 302.600 ;
        RECT 31.080 302.000 31.280 309.600 ;
        RECT 31.880 302.000 32.080 309.600 ;
        RECT 32.680 302.000 32.880 309.600 ;
        RECT 33.480 302.000 33.680 309.600 ;
        RECT 34.280 302.000 35.180 318.000 ;
        RECT 35.780 310.400 35.980 318.000 ;
        RECT 36.580 310.400 36.780 318.000 ;
        RECT 37.380 310.400 37.580 318.000 ;
        RECT 38.180 310.400 38.380 318.000 ;
        RECT 38.980 317.400 39.330 318.000 ;
        RECT 38.980 317.200 42.930 317.400 ;
        RECT 38.980 316.600 39.330 317.200 ;
        RECT 38.980 316.400 42.930 316.600 ;
        RECT 38.980 315.800 39.330 316.400 ;
        RECT 38.980 315.600 42.930 315.800 ;
        RECT 38.980 315.000 39.330 315.600 ;
        RECT 43.930 315.550 44.330 319.200 ;
        RECT 45.130 319.200 64.330 319.600 ;
        RECT 45.130 315.550 45.530 319.200 ;
        RECT 49.180 319.150 51.480 319.200 ;
        RECT 57.980 319.150 60.280 319.200 ;
        RECT 46.530 318.000 62.930 318.600 ;
        RECT 50.130 317.400 50.480 318.000 ;
        RECT 46.530 317.200 50.480 317.400 ;
        RECT 50.130 316.600 50.480 317.200 ;
        RECT 46.530 316.400 50.480 316.600 ;
        RECT 50.130 315.800 50.480 316.400 ;
        RECT 46.530 315.600 50.480 315.800 ;
        RECT 38.980 314.800 42.930 315.000 ;
        RECT 38.980 314.200 39.330 314.800 ;
        RECT 38.980 314.000 42.930 314.200 ;
        RECT 38.980 313.400 39.330 314.000 ;
        RECT 38.980 313.200 42.930 313.400 ;
        RECT 43.880 313.250 45.580 315.550 ;
        RECT 50.130 315.000 50.480 315.600 ;
        RECT 46.530 314.800 50.480 315.000 ;
        RECT 50.130 314.200 50.480 314.800 ;
        RECT 46.530 314.000 50.480 314.200 ;
        RECT 50.130 313.400 50.480 314.000 ;
        RECT 38.980 312.600 39.330 313.200 ;
        RECT 38.980 312.400 42.930 312.600 ;
        RECT 38.980 311.800 39.330 312.400 ;
        RECT 38.980 311.600 42.930 311.800 ;
        RECT 38.980 311.000 39.330 311.600 ;
        RECT 38.980 310.800 42.930 311.000 ;
        RECT 38.980 310.400 39.330 310.800 ;
        RECT 35.780 302.000 35.980 309.600 ;
        RECT 36.580 302.000 36.780 309.600 ;
        RECT 37.380 302.000 37.580 309.600 ;
        RECT 38.180 302.000 38.380 309.600 ;
        RECT 38.980 309.200 39.330 309.600 ;
        RECT 38.980 309.000 42.930 309.200 ;
        RECT 38.980 308.400 39.330 309.000 ;
        RECT 38.980 308.200 42.930 308.400 ;
        RECT 38.980 307.600 39.330 308.200 ;
        RECT 38.980 307.400 42.930 307.600 ;
        RECT 38.980 306.800 39.330 307.400 ;
        RECT 38.980 306.600 42.930 306.800 ;
        RECT 43.930 306.750 44.330 313.250 ;
        RECT 45.130 306.750 45.530 313.250 ;
        RECT 46.530 313.200 50.480 313.400 ;
        RECT 50.130 312.600 50.480 313.200 ;
        RECT 46.530 312.400 50.480 312.600 ;
        RECT 50.130 311.800 50.480 312.400 ;
        RECT 46.530 311.600 50.480 311.800 ;
        RECT 50.130 311.000 50.480 311.600 ;
        RECT 46.530 310.800 50.480 311.000 ;
        RECT 50.130 310.400 50.480 310.800 ;
        RECT 51.080 310.400 51.280 318.000 ;
        RECT 51.880 310.400 52.080 318.000 ;
        RECT 52.680 310.400 52.880 318.000 ;
        RECT 53.480 310.400 53.680 318.000 ;
        RECT 50.130 309.200 50.480 309.600 ;
        RECT 46.530 309.000 50.480 309.200 ;
        RECT 50.130 308.400 50.480 309.000 ;
        RECT 46.530 308.200 50.480 308.400 ;
        RECT 50.130 307.600 50.480 308.200 ;
        RECT 46.530 307.400 50.480 307.600 ;
        RECT 50.130 306.800 50.480 307.400 ;
        RECT 38.980 306.000 39.330 306.600 ;
        RECT 38.980 305.800 42.930 306.000 ;
        RECT 38.980 305.200 39.330 305.800 ;
        RECT 38.980 305.000 42.930 305.200 ;
        RECT 38.980 304.400 39.330 305.000 ;
        RECT 43.880 304.450 45.580 306.750 ;
        RECT 46.530 306.600 50.480 306.800 ;
        RECT 50.130 306.000 50.480 306.600 ;
        RECT 46.530 305.800 50.480 306.000 ;
        RECT 50.130 305.200 50.480 305.800 ;
        RECT 46.530 305.000 50.480 305.200 ;
        RECT 38.980 304.200 42.930 304.400 ;
        RECT 38.980 303.600 39.330 304.200 ;
        RECT 38.980 303.400 42.930 303.600 ;
        RECT 38.980 302.800 39.330 303.400 ;
        RECT 38.980 302.600 42.930 302.800 ;
        RECT 38.980 302.000 39.330 302.600 ;
        RECT 26.530 301.400 42.930 302.000 ;
        RECT 29.180 300.800 31.480 300.850 ;
        RECT 37.980 300.800 40.280 300.850 ;
        RECT 43.930 300.800 44.330 304.450 ;
        RECT 25.130 300.400 44.330 300.800 ;
        RECT 45.130 300.800 45.530 304.450 ;
        RECT 50.130 304.400 50.480 305.000 ;
        RECT 46.530 304.200 50.480 304.400 ;
        RECT 50.130 303.600 50.480 304.200 ;
        RECT 46.530 303.400 50.480 303.600 ;
        RECT 50.130 302.800 50.480 303.400 ;
        RECT 46.530 302.600 50.480 302.800 ;
        RECT 50.130 302.000 50.480 302.600 ;
        RECT 51.080 302.000 51.280 309.600 ;
        RECT 51.880 302.000 52.080 309.600 ;
        RECT 52.680 302.000 52.880 309.600 ;
        RECT 53.480 302.000 53.680 309.600 ;
        RECT 54.280 302.000 55.180 318.000 ;
        RECT 55.780 310.400 55.980 318.000 ;
        RECT 56.580 310.400 56.780 318.000 ;
        RECT 57.380 310.400 57.580 318.000 ;
        RECT 58.180 310.400 58.380 318.000 ;
        RECT 58.980 317.400 59.330 318.000 ;
        RECT 58.980 317.200 62.930 317.400 ;
        RECT 58.980 316.600 59.330 317.200 ;
        RECT 58.980 316.400 62.930 316.600 ;
        RECT 58.980 315.800 59.330 316.400 ;
        RECT 58.980 315.600 62.930 315.800 ;
        RECT 58.980 315.000 59.330 315.600 ;
        RECT 63.930 315.550 64.330 319.200 ;
        RECT 65.130 319.200 84.330 319.600 ;
        RECT 65.130 315.550 65.530 319.200 ;
        RECT 69.180 319.150 71.480 319.200 ;
        RECT 77.980 319.150 80.280 319.200 ;
        RECT 66.530 318.000 82.930 318.600 ;
        RECT 70.130 317.400 70.480 318.000 ;
        RECT 66.530 317.200 70.480 317.400 ;
        RECT 70.130 316.600 70.480 317.200 ;
        RECT 66.530 316.400 70.480 316.600 ;
        RECT 70.130 315.800 70.480 316.400 ;
        RECT 66.530 315.600 70.480 315.800 ;
        RECT 58.980 314.800 62.930 315.000 ;
        RECT 58.980 314.200 59.330 314.800 ;
        RECT 58.980 314.000 62.930 314.200 ;
        RECT 58.980 313.400 59.330 314.000 ;
        RECT 58.980 313.200 62.930 313.400 ;
        RECT 63.880 313.250 65.580 315.550 ;
        RECT 70.130 315.000 70.480 315.600 ;
        RECT 66.530 314.800 70.480 315.000 ;
        RECT 70.130 314.200 70.480 314.800 ;
        RECT 66.530 314.000 70.480 314.200 ;
        RECT 70.130 313.400 70.480 314.000 ;
        RECT 58.980 312.600 59.330 313.200 ;
        RECT 58.980 312.400 62.930 312.600 ;
        RECT 58.980 311.800 59.330 312.400 ;
        RECT 58.980 311.600 62.930 311.800 ;
        RECT 58.980 311.000 59.330 311.600 ;
        RECT 58.980 310.800 62.930 311.000 ;
        RECT 58.980 310.400 59.330 310.800 ;
        RECT 55.780 302.000 55.980 309.600 ;
        RECT 56.580 302.000 56.780 309.600 ;
        RECT 57.380 302.000 57.580 309.600 ;
        RECT 58.180 302.000 58.380 309.600 ;
        RECT 58.980 309.200 59.330 309.600 ;
        RECT 58.980 309.000 62.930 309.200 ;
        RECT 58.980 308.400 59.330 309.000 ;
        RECT 58.980 308.200 62.930 308.400 ;
        RECT 58.980 307.600 59.330 308.200 ;
        RECT 58.980 307.400 62.930 307.600 ;
        RECT 58.980 306.800 59.330 307.400 ;
        RECT 58.980 306.600 62.930 306.800 ;
        RECT 63.930 306.750 64.330 313.250 ;
        RECT 65.130 306.750 65.530 313.250 ;
        RECT 66.530 313.200 70.480 313.400 ;
        RECT 70.130 312.600 70.480 313.200 ;
        RECT 66.530 312.400 70.480 312.600 ;
        RECT 70.130 311.800 70.480 312.400 ;
        RECT 66.530 311.600 70.480 311.800 ;
        RECT 70.130 311.000 70.480 311.600 ;
        RECT 66.530 310.800 70.480 311.000 ;
        RECT 70.130 310.400 70.480 310.800 ;
        RECT 71.080 310.400 71.280 318.000 ;
        RECT 71.880 310.400 72.080 318.000 ;
        RECT 72.680 310.400 72.880 318.000 ;
        RECT 73.480 310.400 73.680 318.000 ;
        RECT 70.130 309.200 70.480 309.600 ;
        RECT 66.530 309.000 70.480 309.200 ;
        RECT 70.130 308.400 70.480 309.000 ;
        RECT 66.530 308.200 70.480 308.400 ;
        RECT 70.130 307.600 70.480 308.200 ;
        RECT 66.530 307.400 70.480 307.600 ;
        RECT 70.130 306.800 70.480 307.400 ;
        RECT 58.980 306.000 59.330 306.600 ;
        RECT 58.980 305.800 62.930 306.000 ;
        RECT 58.980 305.200 59.330 305.800 ;
        RECT 58.980 305.000 62.930 305.200 ;
        RECT 58.980 304.400 59.330 305.000 ;
        RECT 63.880 304.450 65.580 306.750 ;
        RECT 66.530 306.600 70.480 306.800 ;
        RECT 70.130 306.000 70.480 306.600 ;
        RECT 66.530 305.800 70.480 306.000 ;
        RECT 70.130 305.200 70.480 305.800 ;
        RECT 66.530 305.000 70.480 305.200 ;
        RECT 58.980 304.200 62.930 304.400 ;
        RECT 58.980 303.600 59.330 304.200 ;
        RECT 58.980 303.400 62.930 303.600 ;
        RECT 58.980 302.800 59.330 303.400 ;
        RECT 58.980 302.600 62.930 302.800 ;
        RECT 58.980 302.000 59.330 302.600 ;
        RECT 46.530 301.400 62.930 302.000 ;
        RECT 49.180 300.800 51.480 300.850 ;
        RECT 57.980 300.800 60.280 300.850 ;
        RECT 63.930 300.800 64.330 304.450 ;
        RECT 45.130 300.400 64.330 300.800 ;
        RECT 65.130 300.800 65.530 304.450 ;
        RECT 70.130 304.400 70.480 305.000 ;
        RECT 66.530 304.200 70.480 304.400 ;
        RECT 70.130 303.600 70.480 304.200 ;
        RECT 66.530 303.400 70.480 303.600 ;
        RECT 70.130 302.800 70.480 303.400 ;
        RECT 66.530 302.600 70.480 302.800 ;
        RECT 70.130 302.000 70.480 302.600 ;
        RECT 71.080 302.000 71.280 309.600 ;
        RECT 71.880 302.000 72.080 309.600 ;
        RECT 72.680 302.000 72.880 309.600 ;
        RECT 73.480 302.000 73.680 309.600 ;
        RECT 74.280 302.000 75.180 318.000 ;
        RECT 75.780 310.400 75.980 318.000 ;
        RECT 76.580 310.400 76.780 318.000 ;
        RECT 77.380 310.400 77.580 318.000 ;
        RECT 78.180 310.400 78.380 318.000 ;
        RECT 78.980 317.400 79.330 318.000 ;
        RECT 78.980 317.200 82.930 317.400 ;
        RECT 78.980 316.600 79.330 317.200 ;
        RECT 78.980 316.400 82.930 316.600 ;
        RECT 78.980 315.800 79.330 316.400 ;
        RECT 78.980 315.600 82.930 315.800 ;
        RECT 78.980 315.000 79.330 315.600 ;
        RECT 83.930 315.550 84.330 319.200 ;
        RECT 85.130 319.200 104.330 319.600 ;
        RECT 85.130 315.550 85.530 319.200 ;
        RECT 89.180 319.150 91.480 319.200 ;
        RECT 97.980 319.150 100.280 319.200 ;
        RECT 86.530 318.000 102.930 318.600 ;
        RECT 90.130 317.400 90.480 318.000 ;
        RECT 86.530 317.200 90.480 317.400 ;
        RECT 90.130 316.600 90.480 317.200 ;
        RECT 86.530 316.400 90.480 316.600 ;
        RECT 90.130 315.800 90.480 316.400 ;
        RECT 86.530 315.600 90.480 315.800 ;
        RECT 78.980 314.800 82.930 315.000 ;
        RECT 78.980 314.200 79.330 314.800 ;
        RECT 78.980 314.000 82.930 314.200 ;
        RECT 78.980 313.400 79.330 314.000 ;
        RECT 78.980 313.200 82.930 313.400 ;
        RECT 83.880 313.250 85.580 315.550 ;
        RECT 90.130 315.000 90.480 315.600 ;
        RECT 86.530 314.800 90.480 315.000 ;
        RECT 90.130 314.200 90.480 314.800 ;
        RECT 86.530 314.000 90.480 314.200 ;
        RECT 90.130 313.400 90.480 314.000 ;
        RECT 78.980 312.600 79.330 313.200 ;
        RECT 78.980 312.400 82.930 312.600 ;
        RECT 78.980 311.800 79.330 312.400 ;
        RECT 78.980 311.600 82.930 311.800 ;
        RECT 78.980 311.000 79.330 311.600 ;
        RECT 78.980 310.800 82.930 311.000 ;
        RECT 78.980 310.400 79.330 310.800 ;
        RECT 75.780 302.000 75.980 309.600 ;
        RECT 76.580 302.000 76.780 309.600 ;
        RECT 77.380 302.000 77.580 309.600 ;
        RECT 78.180 302.000 78.380 309.600 ;
        RECT 78.980 309.200 79.330 309.600 ;
        RECT 78.980 309.000 82.930 309.200 ;
        RECT 78.980 308.400 79.330 309.000 ;
        RECT 78.980 308.200 82.930 308.400 ;
        RECT 78.980 307.600 79.330 308.200 ;
        RECT 78.980 307.400 82.930 307.600 ;
        RECT 78.980 306.800 79.330 307.400 ;
        RECT 78.980 306.600 82.930 306.800 ;
        RECT 83.930 306.750 84.330 313.250 ;
        RECT 85.130 306.750 85.530 313.250 ;
        RECT 86.530 313.200 90.480 313.400 ;
        RECT 90.130 312.600 90.480 313.200 ;
        RECT 86.530 312.400 90.480 312.600 ;
        RECT 90.130 311.800 90.480 312.400 ;
        RECT 86.530 311.600 90.480 311.800 ;
        RECT 90.130 311.000 90.480 311.600 ;
        RECT 86.530 310.800 90.480 311.000 ;
        RECT 90.130 310.400 90.480 310.800 ;
        RECT 91.080 310.400 91.280 318.000 ;
        RECT 91.880 310.400 92.080 318.000 ;
        RECT 92.680 310.400 92.880 318.000 ;
        RECT 93.480 310.400 93.680 318.000 ;
        RECT 90.130 309.200 90.480 309.600 ;
        RECT 86.530 309.000 90.480 309.200 ;
        RECT 90.130 308.400 90.480 309.000 ;
        RECT 86.530 308.200 90.480 308.400 ;
        RECT 90.130 307.600 90.480 308.200 ;
        RECT 86.530 307.400 90.480 307.600 ;
        RECT 90.130 306.800 90.480 307.400 ;
        RECT 78.980 306.000 79.330 306.600 ;
        RECT 78.980 305.800 82.930 306.000 ;
        RECT 78.980 305.200 79.330 305.800 ;
        RECT 78.980 305.000 82.930 305.200 ;
        RECT 78.980 304.400 79.330 305.000 ;
        RECT 83.880 304.450 85.580 306.750 ;
        RECT 86.530 306.600 90.480 306.800 ;
        RECT 90.130 306.000 90.480 306.600 ;
        RECT 86.530 305.800 90.480 306.000 ;
        RECT 90.130 305.200 90.480 305.800 ;
        RECT 86.530 305.000 90.480 305.200 ;
        RECT 78.980 304.200 82.930 304.400 ;
        RECT 78.980 303.600 79.330 304.200 ;
        RECT 78.980 303.400 82.930 303.600 ;
        RECT 78.980 302.800 79.330 303.400 ;
        RECT 78.980 302.600 82.930 302.800 ;
        RECT 78.980 302.000 79.330 302.600 ;
        RECT 66.530 301.400 82.930 302.000 ;
        RECT 69.180 300.800 71.480 300.850 ;
        RECT 77.980 300.800 80.280 300.850 ;
        RECT 83.930 300.800 84.330 304.450 ;
        RECT 65.130 300.400 84.330 300.800 ;
        RECT 85.130 300.800 85.530 304.450 ;
        RECT 90.130 304.400 90.480 305.000 ;
        RECT 86.530 304.200 90.480 304.400 ;
        RECT 90.130 303.600 90.480 304.200 ;
        RECT 86.530 303.400 90.480 303.600 ;
        RECT 90.130 302.800 90.480 303.400 ;
        RECT 86.530 302.600 90.480 302.800 ;
        RECT 90.130 302.000 90.480 302.600 ;
        RECT 91.080 302.000 91.280 309.600 ;
        RECT 91.880 302.000 92.080 309.600 ;
        RECT 92.680 302.000 92.880 309.600 ;
        RECT 93.480 302.000 93.680 309.600 ;
        RECT 94.280 302.000 95.180 318.000 ;
        RECT 95.780 310.400 95.980 318.000 ;
        RECT 96.580 310.400 96.780 318.000 ;
        RECT 97.380 310.400 97.580 318.000 ;
        RECT 98.180 310.400 98.380 318.000 ;
        RECT 98.980 317.400 99.330 318.000 ;
        RECT 98.980 317.200 102.930 317.400 ;
        RECT 98.980 316.600 99.330 317.200 ;
        RECT 98.980 316.400 102.930 316.600 ;
        RECT 98.980 315.800 99.330 316.400 ;
        RECT 98.980 315.600 102.930 315.800 ;
        RECT 98.980 315.000 99.330 315.600 ;
        RECT 103.930 315.550 104.330 319.200 ;
        RECT 105.340 317.080 105.700 317.460 ;
        RECT 105.970 317.080 106.330 317.460 ;
        RECT 106.570 317.080 106.930 317.460 ;
        RECT 105.340 316.490 105.700 316.870 ;
        RECT 105.970 316.490 106.330 316.870 ;
        RECT 106.570 316.490 106.930 316.870 ;
        RECT 98.980 314.800 102.930 315.000 ;
        RECT 98.980 314.200 99.330 314.800 ;
        RECT 98.980 314.000 102.930 314.200 ;
        RECT 98.980 313.400 99.330 314.000 ;
        RECT 98.980 313.200 102.930 313.400 ;
        RECT 103.880 313.250 104.730 315.550 ;
        RECT 98.980 312.600 99.330 313.200 ;
        RECT 98.980 312.400 102.930 312.600 ;
        RECT 98.980 311.800 99.330 312.400 ;
        RECT 98.980 311.600 102.930 311.800 ;
        RECT 98.980 311.000 99.330 311.600 ;
        RECT 98.980 310.800 102.930 311.000 ;
        RECT 98.980 310.400 99.330 310.800 ;
        RECT 95.780 302.000 95.980 309.600 ;
        RECT 96.580 302.000 96.780 309.600 ;
        RECT 97.380 302.000 97.580 309.600 ;
        RECT 98.180 302.000 98.380 309.600 ;
        RECT 98.980 309.200 99.330 309.600 ;
        RECT 98.980 309.000 102.930 309.200 ;
        RECT 98.980 308.400 99.330 309.000 ;
        RECT 98.980 308.200 102.930 308.400 ;
        RECT 98.980 307.600 99.330 308.200 ;
        RECT 98.980 307.400 102.930 307.600 ;
        RECT 98.980 306.800 99.330 307.400 ;
        RECT 98.980 306.600 102.930 306.800 ;
        RECT 103.930 306.750 104.330 313.250 ;
        RECT 98.980 306.000 99.330 306.600 ;
        RECT 98.980 305.800 102.930 306.000 ;
        RECT 98.980 305.200 99.330 305.800 ;
        RECT 98.980 305.000 102.930 305.200 ;
        RECT 98.980 304.400 99.330 305.000 ;
        RECT 103.880 304.450 104.730 306.750 ;
        RECT 98.980 304.200 102.930 304.400 ;
        RECT 98.980 303.600 99.330 304.200 ;
        RECT 98.980 303.400 102.930 303.600 ;
        RECT 98.980 302.800 99.330 303.400 ;
        RECT 98.980 302.600 102.930 302.800 ;
        RECT 98.980 302.000 99.330 302.600 ;
        RECT 86.530 301.400 102.930 302.000 ;
        RECT 89.180 300.800 91.480 300.850 ;
        RECT 97.980 300.800 100.280 300.850 ;
        RECT 103.930 300.800 104.330 304.450 ;
        RECT 105.340 303.095 105.700 303.475 ;
        RECT 105.970 303.095 106.330 303.475 ;
        RECT 106.570 303.095 106.930 303.475 ;
        RECT 105.340 302.505 105.700 302.885 ;
        RECT 105.970 302.505 106.330 302.885 ;
        RECT 106.570 302.505 106.930 302.885 ;
        RECT 85.130 300.400 104.330 300.800 ;
        RECT 9.180 299.600 11.480 300.400 ;
        RECT 17.980 299.600 20.280 300.400 ;
        RECT 29.180 299.600 31.480 300.400 ;
        RECT 37.980 299.600 40.280 300.400 ;
        RECT 49.180 299.600 51.480 300.400 ;
        RECT 57.980 299.600 60.280 300.400 ;
        RECT 69.180 299.600 71.480 300.400 ;
        RECT 77.980 299.600 80.280 300.400 ;
        RECT 89.180 299.600 91.480 300.400 ;
        RECT 97.980 299.600 100.280 300.400 ;
        RECT 5.130 299.200 24.330 299.600 ;
        RECT 2.515 297.025 2.875 297.405 ;
        RECT 3.145 297.025 3.505 297.405 ;
        RECT 3.745 297.025 4.105 297.405 ;
        RECT 2.515 296.435 2.875 296.815 ;
        RECT 3.145 296.435 3.505 296.815 ;
        RECT 3.745 296.435 4.105 296.815 ;
        RECT 5.130 295.550 5.530 299.200 ;
        RECT 9.180 299.150 11.480 299.200 ;
        RECT 17.980 299.150 20.280 299.200 ;
        RECT 6.530 298.000 22.930 298.600 ;
        RECT 10.130 297.400 10.480 298.000 ;
        RECT 6.530 297.200 10.480 297.400 ;
        RECT 10.130 296.600 10.480 297.200 ;
        RECT 6.530 296.400 10.480 296.600 ;
        RECT 10.130 295.800 10.480 296.400 ;
        RECT 6.530 295.600 10.480 295.800 ;
        RECT 4.730 295.545 5.580 295.550 ;
        RECT 2.320 295.340 5.580 295.545 ;
        RECT 2.315 293.250 5.580 295.340 ;
        RECT 10.130 295.000 10.480 295.600 ;
        RECT 6.530 294.800 10.480 295.000 ;
        RECT 10.130 294.200 10.480 294.800 ;
        RECT 6.530 294.000 10.480 294.200 ;
        RECT 10.130 293.400 10.480 294.000 ;
        RECT 5.130 286.750 5.530 293.250 ;
        RECT 6.530 293.200 10.480 293.400 ;
        RECT 10.130 292.600 10.480 293.200 ;
        RECT 6.530 292.400 10.480 292.600 ;
        RECT 10.130 291.800 10.480 292.400 ;
        RECT 6.530 291.600 10.480 291.800 ;
        RECT 10.130 291.000 10.480 291.600 ;
        RECT 6.530 290.800 10.480 291.000 ;
        RECT 10.130 290.400 10.480 290.800 ;
        RECT 11.080 290.400 11.280 298.000 ;
        RECT 11.880 290.400 12.080 298.000 ;
        RECT 12.680 290.400 12.880 298.000 ;
        RECT 13.480 290.400 13.680 298.000 ;
        RECT 10.130 289.200 10.480 289.600 ;
        RECT 6.530 289.000 10.480 289.200 ;
        RECT 10.130 288.400 10.480 289.000 ;
        RECT 6.530 288.200 10.480 288.400 ;
        RECT 10.130 287.600 10.480 288.200 ;
        RECT 6.530 287.400 10.480 287.600 ;
        RECT 10.130 286.800 10.480 287.400 ;
        RECT 4.730 286.740 5.580 286.750 ;
        RECT 2.315 284.450 5.580 286.740 ;
        RECT 6.530 286.600 10.480 286.800 ;
        RECT 10.130 286.000 10.480 286.600 ;
        RECT 6.530 285.800 10.480 286.000 ;
        RECT 10.130 285.200 10.480 285.800 ;
        RECT 6.530 285.000 10.480 285.200 ;
        RECT 2.315 284.445 4.730 284.450 ;
        RECT 2.515 283.140 2.875 283.520 ;
        RECT 3.145 283.140 3.505 283.520 ;
        RECT 3.745 283.140 4.105 283.520 ;
        RECT 2.515 282.550 2.875 282.930 ;
        RECT 3.145 282.550 3.505 282.930 ;
        RECT 3.745 282.550 4.105 282.930 ;
        RECT 5.130 280.800 5.530 284.450 ;
        RECT 10.130 284.400 10.480 285.000 ;
        RECT 6.530 284.200 10.480 284.400 ;
        RECT 10.130 283.600 10.480 284.200 ;
        RECT 6.530 283.400 10.480 283.600 ;
        RECT 10.130 282.800 10.480 283.400 ;
        RECT 6.530 282.600 10.480 282.800 ;
        RECT 10.130 282.000 10.480 282.600 ;
        RECT 11.080 282.000 11.280 289.600 ;
        RECT 11.880 282.000 12.080 289.600 ;
        RECT 12.680 282.000 12.880 289.600 ;
        RECT 13.480 282.000 13.680 289.600 ;
        RECT 14.280 282.000 15.180 298.000 ;
        RECT 15.780 290.400 15.980 298.000 ;
        RECT 16.580 290.400 16.780 298.000 ;
        RECT 17.380 290.400 17.580 298.000 ;
        RECT 18.180 290.400 18.380 298.000 ;
        RECT 18.980 297.400 19.330 298.000 ;
        RECT 18.980 297.200 22.930 297.400 ;
        RECT 18.980 296.600 19.330 297.200 ;
        RECT 18.980 296.400 22.930 296.600 ;
        RECT 18.980 295.800 19.330 296.400 ;
        RECT 18.980 295.600 22.930 295.800 ;
        RECT 18.980 295.000 19.330 295.600 ;
        RECT 23.930 295.550 24.330 299.200 ;
        RECT 25.130 299.200 44.330 299.600 ;
        RECT 25.130 295.550 25.530 299.200 ;
        RECT 29.180 299.150 31.480 299.200 ;
        RECT 37.980 299.150 40.280 299.200 ;
        RECT 26.530 298.000 42.930 298.600 ;
        RECT 30.130 297.400 30.480 298.000 ;
        RECT 26.530 297.200 30.480 297.400 ;
        RECT 30.130 296.600 30.480 297.200 ;
        RECT 26.530 296.400 30.480 296.600 ;
        RECT 30.130 295.800 30.480 296.400 ;
        RECT 26.530 295.600 30.480 295.800 ;
        RECT 18.980 294.800 22.930 295.000 ;
        RECT 18.980 294.200 19.330 294.800 ;
        RECT 18.980 294.000 22.930 294.200 ;
        RECT 18.980 293.400 19.330 294.000 ;
        RECT 18.980 293.200 22.930 293.400 ;
        RECT 23.880 293.250 25.580 295.550 ;
        RECT 30.130 295.000 30.480 295.600 ;
        RECT 26.530 294.800 30.480 295.000 ;
        RECT 30.130 294.200 30.480 294.800 ;
        RECT 26.530 294.000 30.480 294.200 ;
        RECT 30.130 293.400 30.480 294.000 ;
        RECT 18.980 292.600 19.330 293.200 ;
        RECT 18.980 292.400 22.930 292.600 ;
        RECT 18.980 291.800 19.330 292.400 ;
        RECT 18.980 291.600 22.930 291.800 ;
        RECT 18.980 291.000 19.330 291.600 ;
        RECT 18.980 290.800 22.930 291.000 ;
        RECT 18.980 290.400 19.330 290.800 ;
        RECT 15.780 282.000 15.980 289.600 ;
        RECT 16.580 282.000 16.780 289.600 ;
        RECT 17.380 282.000 17.580 289.600 ;
        RECT 18.180 282.000 18.380 289.600 ;
        RECT 18.980 289.200 19.330 289.600 ;
        RECT 18.980 289.000 22.930 289.200 ;
        RECT 18.980 288.400 19.330 289.000 ;
        RECT 18.980 288.200 22.930 288.400 ;
        RECT 18.980 287.600 19.330 288.200 ;
        RECT 18.980 287.400 22.930 287.600 ;
        RECT 18.980 286.800 19.330 287.400 ;
        RECT 18.980 286.600 22.930 286.800 ;
        RECT 23.930 286.750 24.330 293.250 ;
        RECT 25.130 286.750 25.530 293.250 ;
        RECT 26.530 293.200 30.480 293.400 ;
        RECT 30.130 292.600 30.480 293.200 ;
        RECT 26.530 292.400 30.480 292.600 ;
        RECT 30.130 291.800 30.480 292.400 ;
        RECT 26.530 291.600 30.480 291.800 ;
        RECT 30.130 291.000 30.480 291.600 ;
        RECT 26.530 290.800 30.480 291.000 ;
        RECT 30.130 290.400 30.480 290.800 ;
        RECT 31.080 290.400 31.280 298.000 ;
        RECT 31.880 290.400 32.080 298.000 ;
        RECT 32.680 290.400 32.880 298.000 ;
        RECT 33.480 290.400 33.680 298.000 ;
        RECT 30.130 289.200 30.480 289.600 ;
        RECT 26.530 289.000 30.480 289.200 ;
        RECT 30.130 288.400 30.480 289.000 ;
        RECT 26.530 288.200 30.480 288.400 ;
        RECT 30.130 287.600 30.480 288.200 ;
        RECT 26.530 287.400 30.480 287.600 ;
        RECT 30.130 286.800 30.480 287.400 ;
        RECT 18.980 286.000 19.330 286.600 ;
        RECT 18.980 285.800 22.930 286.000 ;
        RECT 18.980 285.200 19.330 285.800 ;
        RECT 18.980 285.000 22.930 285.200 ;
        RECT 18.980 284.400 19.330 285.000 ;
        RECT 23.880 284.450 25.580 286.750 ;
        RECT 26.530 286.600 30.480 286.800 ;
        RECT 30.130 286.000 30.480 286.600 ;
        RECT 26.530 285.800 30.480 286.000 ;
        RECT 30.130 285.200 30.480 285.800 ;
        RECT 26.530 285.000 30.480 285.200 ;
        RECT 18.980 284.200 22.930 284.400 ;
        RECT 18.980 283.600 19.330 284.200 ;
        RECT 18.980 283.400 22.930 283.600 ;
        RECT 18.980 282.800 19.330 283.400 ;
        RECT 18.980 282.600 22.930 282.800 ;
        RECT 18.980 282.000 19.330 282.600 ;
        RECT 6.530 281.400 22.930 282.000 ;
        RECT 9.180 280.800 11.480 280.850 ;
        RECT 17.980 280.800 20.280 280.850 ;
        RECT 23.930 280.800 24.330 284.450 ;
        RECT 5.130 280.400 24.330 280.800 ;
        RECT 25.130 280.800 25.530 284.450 ;
        RECT 30.130 284.400 30.480 285.000 ;
        RECT 26.530 284.200 30.480 284.400 ;
        RECT 30.130 283.600 30.480 284.200 ;
        RECT 26.530 283.400 30.480 283.600 ;
        RECT 30.130 282.800 30.480 283.400 ;
        RECT 26.530 282.600 30.480 282.800 ;
        RECT 30.130 282.000 30.480 282.600 ;
        RECT 31.080 282.000 31.280 289.600 ;
        RECT 31.880 282.000 32.080 289.600 ;
        RECT 32.680 282.000 32.880 289.600 ;
        RECT 33.480 282.000 33.680 289.600 ;
        RECT 34.280 282.000 35.180 298.000 ;
        RECT 35.780 290.400 35.980 298.000 ;
        RECT 36.580 290.400 36.780 298.000 ;
        RECT 37.380 290.400 37.580 298.000 ;
        RECT 38.180 290.400 38.380 298.000 ;
        RECT 38.980 297.400 39.330 298.000 ;
        RECT 38.980 297.200 42.930 297.400 ;
        RECT 38.980 296.600 39.330 297.200 ;
        RECT 38.980 296.400 42.930 296.600 ;
        RECT 38.980 295.800 39.330 296.400 ;
        RECT 38.980 295.600 42.930 295.800 ;
        RECT 38.980 295.000 39.330 295.600 ;
        RECT 43.930 295.550 44.330 299.200 ;
        RECT 45.130 299.200 64.330 299.600 ;
        RECT 45.130 295.550 45.530 299.200 ;
        RECT 49.180 299.150 51.480 299.200 ;
        RECT 57.980 299.150 60.280 299.200 ;
        RECT 46.530 298.000 62.930 298.600 ;
        RECT 50.130 297.400 50.480 298.000 ;
        RECT 46.530 297.200 50.480 297.400 ;
        RECT 50.130 296.600 50.480 297.200 ;
        RECT 46.530 296.400 50.480 296.600 ;
        RECT 50.130 295.800 50.480 296.400 ;
        RECT 46.530 295.600 50.480 295.800 ;
        RECT 38.980 294.800 42.930 295.000 ;
        RECT 38.980 294.200 39.330 294.800 ;
        RECT 38.980 294.000 42.930 294.200 ;
        RECT 38.980 293.400 39.330 294.000 ;
        RECT 38.980 293.200 42.930 293.400 ;
        RECT 43.880 293.250 45.580 295.550 ;
        RECT 50.130 295.000 50.480 295.600 ;
        RECT 46.530 294.800 50.480 295.000 ;
        RECT 50.130 294.200 50.480 294.800 ;
        RECT 46.530 294.000 50.480 294.200 ;
        RECT 50.130 293.400 50.480 294.000 ;
        RECT 38.980 292.600 39.330 293.200 ;
        RECT 38.980 292.400 42.930 292.600 ;
        RECT 38.980 291.800 39.330 292.400 ;
        RECT 38.980 291.600 42.930 291.800 ;
        RECT 38.980 291.000 39.330 291.600 ;
        RECT 38.980 290.800 42.930 291.000 ;
        RECT 38.980 290.400 39.330 290.800 ;
        RECT 35.780 282.000 35.980 289.600 ;
        RECT 36.580 282.000 36.780 289.600 ;
        RECT 37.380 282.000 37.580 289.600 ;
        RECT 38.180 282.000 38.380 289.600 ;
        RECT 38.980 289.200 39.330 289.600 ;
        RECT 38.980 289.000 42.930 289.200 ;
        RECT 38.980 288.400 39.330 289.000 ;
        RECT 38.980 288.200 42.930 288.400 ;
        RECT 38.980 287.600 39.330 288.200 ;
        RECT 38.980 287.400 42.930 287.600 ;
        RECT 38.980 286.800 39.330 287.400 ;
        RECT 38.980 286.600 42.930 286.800 ;
        RECT 43.930 286.750 44.330 293.250 ;
        RECT 45.130 286.750 45.530 293.250 ;
        RECT 46.530 293.200 50.480 293.400 ;
        RECT 50.130 292.600 50.480 293.200 ;
        RECT 46.530 292.400 50.480 292.600 ;
        RECT 50.130 291.800 50.480 292.400 ;
        RECT 46.530 291.600 50.480 291.800 ;
        RECT 50.130 291.000 50.480 291.600 ;
        RECT 46.530 290.800 50.480 291.000 ;
        RECT 50.130 290.400 50.480 290.800 ;
        RECT 51.080 290.400 51.280 298.000 ;
        RECT 51.880 290.400 52.080 298.000 ;
        RECT 52.680 290.400 52.880 298.000 ;
        RECT 53.480 290.400 53.680 298.000 ;
        RECT 50.130 289.200 50.480 289.600 ;
        RECT 46.530 289.000 50.480 289.200 ;
        RECT 50.130 288.400 50.480 289.000 ;
        RECT 46.530 288.200 50.480 288.400 ;
        RECT 50.130 287.600 50.480 288.200 ;
        RECT 46.530 287.400 50.480 287.600 ;
        RECT 50.130 286.800 50.480 287.400 ;
        RECT 38.980 286.000 39.330 286.600 ;
        RECT 38.980 285.800 42.930 286.000 ;
        RECT 38.980 285.200 39.330 285.800 ;
        RECT 38.980 285.000 42.930 285.200 ;
        RECT 38.980 284.400 39.330 285.000 ;
        RECT 43.880 284.450 45.580 286.750 ;
        RECT 46.530 286.600 50.480 286.800 ;
        RECT 50.130 286.000 50.480 286.600 ;
        RECT 46.530 285.800 50.480 286.000 ;
        RECT 50.130 285.200 50.480 285.800 ;
        RECT 46.530 285.000 50.480 285.200 ;
        RECT 38.980 284.200 42.930 284.400 ;
        RECT 38.980 283.600 39.330 284.200 ;
        RECT 38.980 283.400 42.930 283.600 ;
        RECT 38.980 282.800 39.330 283.400 ;
        RECT 38.980 282.600 42.930 282.800 ;
        RECT 38.980 282.000 39.330 282.600 ;
        RECT 26.530 281.400 42.930 282.000 ;
        RECT 29.180 280.800 31.480 280.850 ;
        RECT 37.980 280.800 40.280 280.850 ;
        RECT 43.930 280.800 44.330 284.450 ;
        RECT 25.130 280.400 44.330 280.800 ;
        RECT 45.130 280.800 45.530 284.450 ;
        RECT 50.130 284.400 50.480 285.000 ;
        RECT 46.530 284.200 50.480 284.400 ;
        RECT 50.130 283.600 50.480 284.200 ;
        RECT 46.530 283.400 50.480 283.600 ;
        RECT 50.130 282.800 50.480 283.400 ;
        RECT 46.530 282.600 50.480 282.800 ;
        RECT 50.130 282.000 50.480 282.600 ;
        RECT 51.080 282.000 51.280 289.600 ;
        RECT 51.880 282.000 52.080 289.600 ;
        RECT 52.680 282.000 52.880 289.600 ;
        RECT 53.480 282.000 53.680 289.600 ;
        RECT 54.280 282.000 55.180 298.000 ;
        RECT 55.780 290.400 55.980 298.000 ;
        RECT 56.580 290.400 56.780 298.000 ;
        RECT 57.380 290.400 57.580 298.000 ;
        RECT 58.180 290.400 58.380 298.000 ;
        RECT 58.980 297.400 59.330 298.000 ;
        RECT 58.980 297.200 62.930 297.400 ;
        RECT 58.980 296.600 59.330 297.200 ;
        RECT 58.980 296.400 62.930 296.600 ;
        RECT 58.980 295.800 59.330 296.400 ;
        RECT 58.980 295.600 62.930 295.800 ;
        RECT 58.980 295.000 59.330 295.600 ;
        RECT 63.930 295.550 64.330 299.200 ;
        RECT 65.130 299.200 84.330 299.600 ;
        RECT 65.130 295.550 65.530 299.200 ;
        RECT 69.180 299.150 71.480 299.200 ;
        RECT 77.980 299.150 80.280 299.200 ;
        RECT 66.530 298.000 82.930 298.600 ;
        RECT 70.130 297.400 70.480 298.000 ;
        RECT 66.530 297.200 70.480 297.400 ;
        RECT 70.130 296.600 70.480 297.200 ;
        RECT 66.530 296.400 70.480 296.600 ;
        RECT 70.130 295.800 70.480 296.400 ;
        RECT 66.530 295.600 70.480 295.800 ;
        RECT 58.980 294.800 62.930 295.000 ;
        RECT 58.980 294.200 59.330 294.800 ;
        RECT 58.980 294.000 62.930 294.200 ;
        RECT 58.980 293.400 59.330 294.000 ;
        RECT 58.980 293.200 62.930 293.400 ;
        RECT 63.880 293.250 65.580 295.550 ;
        RECT 70.130 295.000 70.480 295.600 ;
        RECT 66.530 294.800 70.480 295.000 ;
        RECT 70.130 294.200 70.480 294.800 ;
        RECT 66.530 294.000 70.480 294.200 ;
        RECT 70.130 293.400 70.480 294.000 ;
        RECT 58.980 292.600 59.330 293.200 ;
        RECT 58.980 292.400 62.930 292.600 ;
        RECT 58.980 291.800 59.330 292.400 ;
        RECT 58.980 291.600 62.930 291.800 ;
        RECT 58.980 291.000 59.330 291.600 ;
        RECT 58.980 290.800 62.930 291.000 ;
        RECT 58.980 290.400 59.330 290.800 ;
        RECT 55.780 282.000 55.980 289.600 ;
        RECT 56.580 282.000 56.780 289.600 ;
        RECT 57.380 282.000 57.580 289.600 ;
        RECT 58.180 282.000 58.380 289.600 ;
        RECT 58.980 289.200 59.330 289.600 ;
        RECT 58.980 289.000 62.930 289.200 ;
        RECT 58.980 288.400 59.330 289.000 ;
        RECT 58.980 288.200 62.930 288.400 ;
        RECT 58.980 287.600 59.330 288.200 ;
        RECT 58.980 287.400 62.930 287.600 ;
        RECT 58.980 286.800 59.330 287.400 ;
        RECT 58.980 286.600 62.930 286.800 ;
        RECT 63.930 286.750 64.330 293.250 ;
        RECT 65.130 286.750 65.530 293.250 ;
        RECT 66.530 293.200 70.480 293.400 ;
        RECT 70.130 292.600 70.480 293.200 ;
        RECT 66.530 292.400 70.480 292.600 ;
        RECT 70.130 291.800 70.480 292.400 ;
        RECT 66.530 291.600 70.480 291.800 ;
        RECT 70.130 291.000 70.480 291.600 ;
        RECT 66.530 290.800 70.480 291.000 ;
        RECT 70.130 290.400 70.480 290.800 ;
        RECT 71.080 290.400 71.280 298.000 ;
        RECT 71.880 290.400 72.080 298.000 ;
        RECT 72.680 290.400 72.880 298.000 ;
        RECT 73.480 290.400 73.680 298.000 ;
        RECT 70.130 289.200 70.480 289.600 ;
        RECT 66.530 289.000 70.480 289.200 ;
        RECT 70.130 288.400 70.480 289.000 ;
        RECT 66.530 288.200 70.480 288.400 ;
        RECT 70.130 287.600 70.480 288.200 ;
        RECT 66.530 287.400 70.480 287.600 ;
        RECT 70.130 286.800 70.480 287.400 ;
        RECT 58.980 286.000 59.330 286.600 ;
        RECT 58.980 285.800 62.930 286.000 ;
        RECT 58.980 285.200 59.330 285.800 ;
        RECT 58.980 285.000 62.930 285.200 ;
        RECT 58.980 284.400 59.330 285.000 ;
        RECT 63.880 284.450 65.580 286.750 ;
        RECT 66.530 286.600 70.480 286.800 ;
        RECT 70.130 286.000 70.480 286.600 ;
        RECT 66.530 285.800 70.480 286.000 ;
        RECT 70.130 285.200 70.480 285.800 ;
        RECT 66.530 285.000 70.480 285.200 ;
        RECT 58.980 284.200 62.930 284.400 ;
        RECT 58.980 283.600 59.330 284.200 ;
        RECT 58.980 283.400 62.930 283.600 ;
        RECT 58.980 282.800 59.330 283.400 ;
        RECT 58.980 282.600 62.930 282.800 ;
        RECT 58.980 282.000 59.330 282.600 ;
        RECT 46.530 281.400 62.930 282.000 ;
        RECT 49.180 280.800 51.480 280.850 ;
        RECT 57.980 280.800 60.280 280.850 ;
        RECT 63.930 280.800 64.330 284.450 ;
        RECT 45.130 280.400 64.330 280.800 ;
        RECT 65.130 280.800 65.530 284.450 ;
        RECT 70.130 284.400 70.480 285.000 ;
        RECT 66.530 284.200 70.480 284.400 ;
        RECT 70.130 283.600 70.480 284.200 ;
        RECT 66.530 283.400 70.480 283.600 ;
        RECT 70.130 282.800 70.480 283.400 ;
        RECT 66.530 282.600 70.480 282.800 ;
        RECT 70.130 282.000 70.480 282.600 ;
        RECT 71.080 282.000 71.280 289.600 ;
        RECT 71.880 282.000 72.080 289.600 ;
        RECT 72.680 282.000 72.880 289.600 ;
        RECT 73.480 282.000 73.680 289.600 ;
        RECT 74.280 282.000 75.180 298.000 ;
        RECT 75.780 290.400 75.980 298.000 ;
        RECT 76.580 290.400 76.780 298.000 ;
        RECT 77.380 290.400 77.580 298.000 ;
        RECT 78.180 290.400 78.380 298.000 ;
        RECT 78.980 297.400 79.330 298.000 ;
        RECT 78.980 297.200 82.930 297.400 ;
        RECT 78.980 296.600 79.330 297.200 ;
        RECT 78.980 296.400 82.930 296.600 ;
        RECT 78.980 295.800 79.330 296.400 ;
        RECT 78.980 295.600 82.930 295.800 ;
        RECT 78.980 295.000 79.330 295.600 ;
        RECT 83.930 295.550 84.330 299.200 ;
        RECT 85.130 299.200 104.330 299.600 ;
        RECT 85.130 295.550 85.530 299.200 ;
        RECT 89.180 299.150 91.480 299.200 ;
        RECT 97.980 299.150 100.280 299.200 ;
        RECT 86.530 298.000 102.930 298.600 ;
        RECT 90.130 297.400 90.480 298.000 ;
        RECT 86.530 297.200 90.480 297.400 ;
        RECT 90.130 296.600 90.480 297.200 ;
        RECT 86.530 296.400 90.480 296.600 ;
        RECT 90.130 295.800 90.480 296.400 ;
        RECT 86.530 295.600 90.480 295.800 ;
        RECT 78.980 294.800 82.930 295.000 ;
        RECT 78.980 294.200 79.330 294.800 ;
        RECT 78.980 294.000 82.930 294.200 ;
        RECT 78.980 293.400 79.330 294.000 ;
        RECT 78.980 293.200 82.930 293.400 ;
        RECT 83.880 293.250 85.580 295.550 ;
        RECT 90.130 295.000 90.480 295.600 ;
        RECT 86.530 294.800 90.480 295.000 ;
        RECT 90.130 294.200 90.480 294.800 ;
        RECT 86.530 294.000 90.480 294.200 ;
        RECT 90.130 293.400 90.480 294.000 ;
        RECT 78.980 292.600 79.330 293.200 ;
        RECT 78.980 292.400 82.930 292.600 ;
        RECT 78.980 291.800 79.330 292.400 ;
        RECT 78.980 291.600 82.930 291.800 ;
        RECT 78.980 291.000 79.330 291.600 ;
        RECT 78.980 290.800 82.930 291.000 ;
        RECT 78.980 290.400 79.330 290.800 ;
        RECT 75.780 282.000 75.980 289.600 ;
        RECT 76.580 282.000 76.780 289.600 ;
        RECT 77.380 282.000 77.580 289.600 ;
        RECT 78.180 282.000 78.380 289.600 ;
        RECT 78.980 289.200 79.330 289.600 ;
        RECT 78.980 289.000 82.930 289.200 ;
        RECT 78.980 288.400 79.330 289.000 ;
        RECT 78.980 288.200 82.930 288.400 ;
        RECT 78.980 287.600 79.330 288.200 ;
        RECT 78.980 287.400 82.930 287.600 ;
        RECT 78.980 286.800 79.330 287.400 ;
        RECT 78.980 286.600 82.930 286.800 ;
        RECT 83.930 286.750 84.330 293.250 ;
        RECT 85.130 286.750 85.530 293.250 ;
        RECT 86.530 293.200 90.480 293.400 ;
        RECT 90.130 292.600 90.480 293.200 ;
        RECT 86.530 292.400 90.480 292.600 ;
        RECT 90.130 291.800 90.480 292.400 ;
        RECT 86.530 291.600 90.480 291.800 ;
        RECT 90.130 291.000 90.480 291.600 ;
        RECT 86.530 290.800 90.480 291.000 ;
        RECT 90.130 290.400 90.480 290.800 ;
        RECT 91.080 290.400 91.280 298.000 ;
        RECT 91.880 290.400 92.080 298.000 ;
        RECT 92.680 290.400 92.880 298.000 ;
        RECT 93.480 290.400 93.680 298.000 ;
        RECT 90.130 289.200 90.480 289.600 ;
        RECT 86.530 289.000 90.480 289.200 ;
        RECT 90.130 288.400 90.480 289.000 ;
        RECT 86.530 288.200 90.480 288.400 ;
        RECT 90.130 287.600 90.480 288.200 ;
        RECT 86.530 287.400 90.480 287.600 ;
        RECT 90.130 286.800 90.480 287.400 ;
        RECT 78.980 286.000 79.330 286.600 ;
        RECT 78.980 285.800 82.930 286.000 ;
        RECT 78.980 285.200 79.330 285.800 ;
        RECT 78.980 285.000 82.930 285.200 ;
        RECT 78.980 284.400 79.330 285.000 ;
        RECT 83.880 284.450 85.580 286.750 ;
        RECT 86.530 286.600 90.480 286.800 ;
        RECT 90.130 286.000 90.480 286.600 ;
        RECT 86.530 285.800 90.480 286.000 ;
        RECT 90.130 285.200 90.480 285.800 ;
        RECT 86.530 285.000 90.480 285.200 ;
        RECT 78.980 284.200 82.930 284.400 ;
        RECT 78.980 283.600 79.330 284.200 ;
        RECT 78.980 283.400 82.930 283.600 ;
        RECT 78.980 282.800 79.330 283.400 ;
        RECT 78.980 282.600 82.930 282.800 ;
        RECT 78.980 282.000 79.330 282.600 ;
        RECT 66.530 281.400 82.930 282.000 ;
        RECT 69.180 280.800 71.480 280.850 ;
        RECT 77.980 280.800 80.280 280.850 ;
        RECT 83.930 280.800 84.330 284.450 ;
        RECT 65.130 280.400 84.330 280.800 ;
        RECT 85.130 280.800 85.530 284.450 ;
        RECT 90.130 284.400 90.480 285.000 ;
        RECT 86.530 284.200 90.480 284.400 ;
        RECT 90.130 283.600 90.480 284.200 ;
        RECT 86.530 283.400 90.480 283.600 ;
        RECT 90.130 282.800 90.480 283.400 ;
        RECT 86.530 282.600 90.480 282.800 ;
        RECT 90.130 282.000 90.480 282.600 ;
        RECT 91.080 282.000 91.280 289.600 ;
        RECT 91.880 282.000 92.080 289.600 ;
        RECT 92.680 282.000 92.880 289.600 ;
        RECT 93.480 282.000 93.680 289.600 ;
        RECT 94.280 282.000 95.180 298.000 ;
        RECT 95.780 290.400 95.980 298.000 ;
        RECT 96.580 290.400 96.780 298.000 ;
        RECT 97.380 290.400 97.580 298.000 ;
        RECT 98.180 290.400 98.380 298.000 ;
        RECT 98.980 297.400 99.330 298.000 ;
        RECT 98.980 297.200 102.930 297.400 ;
        RECT 98.980 296.600 99.330 297.200 ;
        RECT 98.980 296.400 102.930 296.600 ;
        RECT 98.980 295.800 99.330 296.400 ;
        RECT 98.980 295.600 102.930 295.800 ;
        RECT 98.980 295.000 99.330 295.600 ;
        RECT 103.930 295.550 104.330 299.200 ;
        RECT 105.340 297.350 105.700 297.730 ;
        RECT 105.970 297.350 106.330 297.730 ;
        RECT 106.570 297.350 106.930 297.730 ;
        RECT 105.340 296.760 105.700 297.140 ;
        RECT 105.970 296.760 106.330 297.140 ;
        RECT 106.570 296.760 106.930 297.140 ;
        RECT 98.980 294.800 102.930 295.000 ;
        RECT 98.980 294.200 99.330 294.800 ;
        RECT 98.980 294.000 102.930 294.200 ;
        RECT 98.980 293.400 99.330 294.000 ;
        RECT 98.980 293.200 102.930 293.400 ;
        RECT 103.880 293.250 104.730 295.550 ;
        RECT 98.980 292.600 99.330 293.200 ;
        RECT 98.980 292.400 102.930 292.600 ;
        RECT 98.980 291.800 99.330 292.400 ;
        RECT 98.980 291.600 102.930 291.800 ;
        RECT 98.980 291.000 99.330 291.600 ;
        RECT 98.980 290.800 102.930 291.000 ;
        RECT 98.980 290.400 99.330 290.800 ;
        RECT 95.780 282.000 95.980 289.600 ;
        RECT 96.580 282.000 96.780 289.600 ;
        RECT 97.380 282.000 97.580 289.600 ;
        RECT 98.180 282.000 98.380 289.600 ;
        RECT 98.980 289.200 99.330 289.600 ;
        RECT 98.980 289.000 102.930 289.200 ;
        RECT 98.980 288.400 99.330 289.000 ;
        RECT 98.980 288.200 102.930 288.400 ;
        RECT 98.980 287.600 99.330 288.200 ;
        RECT 98.980 287.400 102.930 287.600 ;
        RECT 98.980 286.800 99.330 287.400 ;
        RECT 98.980 286.600 102.930 286.800 ;
        RECT 103.930 286.750 104.330 293.250 ;
        RECT 98.980 286.000 99.330 286.600 ;
        RECT 98.980 285.800 102.930 286.000 ;
        RECT 98.980 285.200 99.330 285.800 ;
        RECT 98.980 285.000 102.930 285.200 ;
        RECT 98.980 284.400 99.330 285.000 ;
        RECT 103.880 284.450 104.730 286.750 ;
        RECT 98.980 284.200 102.930 284.400 ;
        RECT 98.980 283.600 99.330 284.200 ;
        RECT 98.980 283.400 102.930 283.600 ;
        RECT 98.980 282.800 99.330 283.400 ;
        RECT 98.980 282.600 102.930 282.800 ;
        RECT 98.980 282.000 99.330 282.600 ;
        RECT 86.530 281.400 102.930 282.000 ;
        RECT 89.180 280.800 91.480 280.850 ;
        RECT 97.980 280.800 100.280 280.850 ;
        RECT 103.930 280.800 104.330 284.450 ;
        RECT 105.340 282.770 105.700 283.150 ;
        RECT 105.970 282.770 106.330 283.150 ;
        RECT 106.570 282.770 106.930 283.150 ;
        RECT 105.340 282.180 105.700 282.560 ;
        RECT 105.970 282.180 106.330 282.560 ;
        RECT 106.570 282.180 106.930 282.560 ;
        RECT 85.130 280.400 104.330 280.800 ;
        RECT 9.180 279.600 11.480 280.400 ;
        RECT 17.980 279.600 20.280 280.400 ;
        RECT 29.180 279.600 31.480 280.400 ;
        RECT 37.980 279.600 40.280 280.400 ;
        RECT 49.180 279.600 51.480 280.400 ;
        RECT 57.980 279.600 60.280 280.400 ;
        RECT 69.180 279.600 71.480 280.400 ;
        RECT 77.980 279.600 80.280 280.400 ;
        RECT 89.180 279.600 91.480 280.400 ;
        RECT 97.980 279.600 100.280 280.400 ;
        RECT 5.130 279.200 24.330 279.600 ;
        RECT 2.515 277.105 2.875 277.485 ;
        RECT 3.145 277.105 3.505 277.485 ;
        RECT 3.745 277.105 4.105 277.485 ;
        RECT 2.515 276.515 2.875 276.895 ;
        RECT 3.145 276.515 3.505 276.895 ;
        RECT 3.745 276.515 4.105 276.895 ;
        RECT 5.130 275.550 5.530 279.200 ;
        RECT 9.180 279.150 11.480 279.200 ;
        RECT 17.980 279.150 20.280 279.200 ;
        RECT 6.530 278.000 22.930 278.600 ;
        RECT 10.130 277.400 10.480 278.000 ;
        RECT 6.530 277.200 10.480 277.400 ;
        RECT 10.130 276.600 10.480 277.200 ;
        RECT 6.530 276.400 10.480 276.600 ;
        RECT 10.130 275.800 10.480 276.400 ;
        RECT 6.530 275.600 10.480 275.800 ;
        RECT 4.730 275.545 5.580 275.550 ;
        RECT 2.315 273.250 5.580 275.545 ;
        RECT 10.130 275.000 10.480 275.600 ;
        RECT 6.530 274.800 10.480 275.000 ;
        RECT 10.130 274.200 10.480 274.800 ;
        RECT 6.530 274.000 10.480 274.200 ;
        RECT 10.130 273.400 10.480 274.000 ;
        RECT 5.130 266.750 5.530 273.250 ;
        RECT 6.530 273.200 10.480 273.400 ;
        RECT 10.130 272.600 10.480 273.200 ;
        RECT 6.530 272.400 10.480 272.600 ;
        RECT 10.130 271.800 10.480 272.400 ;
        RECT 6.530 271.600 10.480 271.800 ;
        RECT 10.130 271.000 10.480 271.600 ;
        RECT 6.530 270.800 10.480 271.000 ;
        RECT 10.130 270.400 10.480 270.800 ;
        RECT 11.080 270.400 11.280 278.000 ;
        RECT 11.880 270.400 12.080 278.000 ;
        RECT 12.680 270.400 12.880 278.000 ;
        RECT 13.480 270.400 13.680 278.000 ;
        RECT 10.130 269.200 10.480 269.600 ;
        RECT 6.530 269.000 10.480 269.200 ;
        RECT 10.130 268.400 10.480 269.000 ;
        RECT 6.530 268.200 10.480 268.400 ;
        RECT 10.130 267.600 10.480 268.200 ;
        RECT 6.530 267.400 10.480 267.600 ;
        RECT 10.130 266.800 10.480 267.400 ;
        RECT 2.315 264.455 5.580 266.750 ;
        RECT 6.530 266.600 10.480 266.800 ;
        RECT 10.130 266.000 10.480 266.600 ;
        RECT 6.530 265.800 10.480 266.000 ;
        RECT 10.130 265.200 10.480 265.800 ;
        RECT 6.530 265.000 10.480 265.200 ;
        RECT 4.730 264.450 5.580 264.455 ;
        RECT 2.515 263.275 2.875 263.655 ;
        RECT 3.145 263.275 3.505 263.655 ;
        RECT 3.745 263.275 4.105 263.655 ;
        RECT 2.515 262.685 2.875 263.065 ;
        RECT 3.145 262.685 3.505 263.065 ;
        RECT 3.745 262.685 4.105 263.065 ;
        RECT 5.130 260.800 5.530 264.450 ;
        RECT 10.130 264.400 10.480 265.000 ;
        RECT 6.530 264.200 10.480 264.400 ;
        RECT 10.130 263.600 10.480 264.200 ;
        RECT 6.530 263.400 10.480 263.600 ;
        RECT 10.130 262.800 10.480 263.400 ;
        RECT 6.530 262.600 10.480 262.800 ;
        RECT 10.130 262.000 10.480 262.600 ;
        RECT 11.080 262.000 11.280 269.600 ;
        RECT 11.880 262.000 12.080 269.600 ;
        RECT 12.680 262.000 12.880 269.600 ;
        RECT 13.480 262.000 13.680 269.600 ;
        RECT 14.280 262.000 15.180 278.000 ;
        RECT 15.780 270.400 15.980 278.000 ;
        RECT 16.580 270.400 16.780 278.000 ;
        RECT 17.380 270.400 17.580 278.000 ;
        RECT 18.180 270.400 18.380 278.000 ;
        RECT 18.980 277.400 19.330 278.000 ;
        RECT 18.980 277.200 22.930 277.400 ;
        RECT 18.980 276.600 19.330 277.200 ;
        RECT 18.980 276.400 22.930 276.600 ;
        RECT 18.980 275.800 19.330 276.400 ;
        RECT 18.980 275.600 22.930 275.800 ;
        RECT 18.980 275.000 19.330 275.600 ;
        RECT 23.930 275.550 24.330 279.200 ;
        RECT 25.130 279.200 44.330 279.600 ;
        RECT 25.130 275.550 25.530 279.200 ;
        RECT 29.180 279.150 31.480 279.200 ;
        RECT 37.980 279.150 40.280 279.200 ;
        RECT 26.530 278.000 42.930 278.600 ;
        RECT 30.130 277.400 30.480 278.000 ;
        RECT 26.530 277.200 30.480 277.400 ;
        RECT 30.130 276.600 30.480 277.200 ;
        RECT 26.530 276.400 30.480 276.600 ;
        RECT 30.130 275.800 30.480 276.400 ;
        RECT 26.530 275.600 30.480 275.800 ;
        RECT 18.980 274.800 22.930 275.000 ;
        RECT 18.980 274.200 19.330 274.800 ;
        RECT 18.980 274.000 22.930 274.200 ;
        RECT 18.980 273.400 19.330 274.000 ;
        RECT 18.980 273.200 22.930 273.400 ;
        RECT 23.880 273.250 25.580 275.550 ;
        RECT 30.130 275.000 30.480 275.600 ;
        RECT 26.530 274.800 30.480 275.000 ;
        RECT 30.130 274.200 30.480 274.800 ;
        RECT 26.530 274.000 30.480 274.200 ;
        RECT 30.130 273.400 30.480 274.000 ;
        RECT 18.980 272.600 19.330 273.200 ;
        RECT 18.980 272.400 22.930 272.600 ;
        RECT 18.980 271.800 19.330 272.400 ;
        RECT 18.980 271.600 22.930 271.800 ;
        RECT 18.980 271.000 19.330 271.600 ;
        RECT 18.980 270.800 22.930 271.000 ;
        RECT 18.980 270.400 19.330 270.800 ;
        RECT 15.780 262.000 15.980 269.600 ;
        RECT 16.580 262.000 16.780 269.600 ;
        RECT 17.380 262.000 17.580 269.600 ;
        RECT 18.180 262.000 18.380 269.600 ;
        RECT 18.980 269.200 19.330 269.600 ;
        RECT 18.980 269.000 22.930 269.200 ;
        RECT 18.980 268.400 19.330 269.000 ;
        RECT 18.980 268.200 22.930 268.400 ;
        RECT 18.980 267.600 19.330 268.200 ;
        RECT 18.980 267.400 22.930 267.600 ;
        RECT 18.980 266.800 19.330 267.400 ;
        RECT 18.980 266.600 22.930 266.800 ;
        RECT 23.930 266.750 24.330 273.250 ;
        RECT 25.130 266.750 25.530 273.250 ;
        RECT 26.530 273.200 30.480 273.400 ;
        RECT 30.130 272.600 30.480 273.200 ;
        RECT 26.530 272.400 30.480 272.600 ;
        RECT 30.130 271.800 30.480 272.400 ;
        RECT 26.530 271.600 30.480 271.800 ;
        RECT 30.130 271.000 30.480 271.600 ;
        RECT 26.530 270.800 30.480 271.000 ;
        RECT 30.130 270.400 30.480 270.800 ;
        RECT 31.080 270.400 31.280 278.000 ;
        RECT 31.880 270.400 32.080 278.000 ;
        RECT 32.680 270.400 32.880 278.000 ;
        RECT 33.480 270.400 33.680 278.000 ;
        RECT 30.130 269.200 30.480 269.600 ;
        RECT 26.530 269.000 30.480 269.200 ;
        RECT 30.130 268.400 30.480 269.000 ;
        RECT 26.530 268.200 30.480 268.400 ;
        RECT 30.130 267.600 30.480 268.200 ;
        RECT 26.530 267.400 30.480 267.600 ;
        RECT 30.130 266.800 30.480 267.400 ;
        RECT 18.980 266.000 19.330 266.600 ;
        RECT 18.980 265.800 22.930 266.000 ;
        RECT 18.980 265.200 19.330 265.800 ;
        RECT 18.980 265.000 22.930 265.200 ;
        RECT 18.980 264.400 19.330 265.000 ;
        RECT 23.880 264.450 25.580 266.750 ;
        RECT 26.530 266.600 30.480 266.800 ;
        RECT 30.130 266.000 30.480 266.600 ;
        RECT 26.530 265.800 30.480 266.000 ;
        RECT 30.130 265.200 30.480 265.800 ;
        RECT 26.530 265.000 30.480 265.200 ;
        RECT 18.980 264.200 22.930 264.400 ;
        RECT 18.980 263.600 19.330 264.200 ;
        RECT 18.980 263.400 22.930 263.600 ;
        RECT 18.980 262.800 19.330 263.400 ;
        RECT 18.980 262.600 22.930 262.800 ;
        RECT 18.980 262.000 19.330 262.600 ;
        RECT 6.530 261.400 22.930 262.000 ;
        RECT 9.180 260.800 11.480 260.850 ;
        RECT 17.980 260.800 20.280 260.850 ;
        RECT 23.930 260.800 24.330 264.450 ;
        RECT 5.130 260.400 24.330 260.800 ;
        RECT 25.130 260.800 25.530 264.450 ;
        RECT 30.130 264.400 30.480 265.000 ;
        RECT 26.530 264.200 30.480 264.400 ;
        RECT 30.130 263.600 30.480 264.200 ;
        RECT 26.530 263.400 30.480 263.600 ;
        RECT 30.130 262.800 30.480 263.400 ;
        RECT 26.530 262.600 30.480 262.800 ;
        RECT 30.130 262.000 30.480 262.600 ;
        RECT 31.080 262.000 31.280 269.600 ;
        RECT 31.880 262.000 32.080 269.600 ;
        RECT 32.680 262.000 32.880 269.600 ;
        RECT 33.480 262.000 33.680 269.600 ;
        RECT 34.280 262.000 35.180 278.000 ;
        RECT 35.780 270.400 35.980 278.000 ;
        RECT 36.580 270.400 36.780 278.000 ;
        RECT 37.380 270.400 37.580 278.000 ;
        RECT 38.180 270.400 38.380 278.000 ;
        RECT 38.980 277.400 39.330 278.000 ;
        RECT 38.980 277.200 42.930 277.400 ;
        RECT 38.980 276.600 39.330 277.200 ;
        RECT 38.980 276.400 42.930 276.600 ;
        RECT 38.980 275.800 39.330 276.400 ;
        RECT 38.980 275.600 42.930 275.800 ;
        RECT 38.980 275.000 39.330 275.600 ;
        RECT 43.930 275.550 44.330 279.200 ;
        RECT 45.130 279.200 64.330 279.600 ;
        RECT 45.130 275.550 45.530 279.200 ;
        RECT 49.180 279.150 51.480 279.200 ;
        RECT 57.980 279.150 60.280 279.200 ;
        RECT 46.530 278.000 62.930 278.600 ;
        RECT 50.130 277.400 50.480 278.000 ;
        RECT 46.530 277.200 50.480 277.400 ;
        RECT 50.130 276.600 50.480 277.200 ;
        RECT 46.530 276.400 50.480 276.600 ;
        RECT 50.130 275.800 50.480 276.400 ;
        RECT 46.530 275.600 50.480 275.800 ;
        RECT 38.980 274.800 42.930 275.000 ;
        RECT 38.980 274.200 39.330 274.800 ;
        RECT 38.980 274.000 42.930 274.200 ;
        RECT 38.980 273.400 39.330 274.000 ;
        RECT 38.980 273.200 42.930 273.400 ;
        RECT 43.880 273.250 45.580 275.550 ;
        RECT 50.130 275.000 50.480 275.600 ;
        RECT 46.530 274.800 50.480 275.000 ;
        RECT 50.130 274.200 50.480 274.800 ;
        RECT 46.530 274.000 50.480 274.200 ;
        RECT 50.130 273.400 50.480 274.000 ;
        RECT 38.980 272.600 39.330 273.200 ;
        RECT 38.980 272.400 42.930 272.600 ;
        RECT 38.980 271.800 39.330 272.400 ;
        RECT 38.980 271.600 42.930 271.800 ;
        RECT 38.980 271.000 39.330 271.600 ;
        RECT 38.980 270.800 42.930 271.000 ;
        RECT 38.980 270.400 39.330 270.800 ;
        RECT 35.780 262.000 35.980 269.600 ;
        RECT 36.580 262.000 36.780 269.600 ;
        RECT 37.380 262.000 37.580 269.600 ;
        RECT 38.180 262.000 38.380 269.600 ;
        RECT 38.980 269.200 39.330 269.600 ;
        RECT 38.980 269.000 42.930 269.200 ;
        RECT 38.980 268.400 39.330 269.000 ;
        RECT 38.980 268.200 42.930 268.400 ;
        RECT 38.980 267.600 39.330 268.200 ;
        RECT 38.980 267.400 42.930 267.600 ;
        RECT 38.980 266.800 39.330 267.400 ;
        RECT 38.980 266.600 42.930 266.800 ;
        RECT 43.930 266.750 44.330 273.250 ;
        RECT 45.130 266.750 45.530 273.250 ;
        RECT 46.530 273.200 50.480 273.400 ;
        RECT 50.130 272.600 50.480 273.200 ;
        RECT 46.530 272.400 50.480 272.600 ;
        RECT 50.130 271.800 50.480 272.400 ;
        RECT 46.530 271.600 50.480 271.800 ;
        RECT 50.130 271.000 50.480 271.600 ;
        RECT 46.530 270.800 50.480 271.000 ;
        RECT 50.130 270.400 50.480 270.800 ;
        RECT 51.080 270.400 51.280 278.000 ;
        RECT 51.880 270.400 52.080 278.000 ;
        RECT 52.680 270.400 52.880 278.000 ;
        RECT 53.480 270.400 53.680 278.000 ;
        RECT 50.130 269.200 50.480 269.600 ;
        RECT 46.530 269.000 50.480 269.200 ;
        RECT 50.130 268.400 50.480 269.000 ;
        RECT 46.530 268.200 50.480 268.400 ;
        RECT 50.130 267.600 50.480 268.200 ;
        RECT 46.530 267.400 50.480 267.600 ;
        RECT 50.130 266.800 50.480 267.400 ;
        RECT 38.980 266.000 39.330 266.600 ;
        RECT 38.980 265.800 42.930 266.000 ;
        RECT 38.980 265.200 39.330 265.800 ;
        RECT 38.980 265.000 42.930 265.200 ;
        RECT 38.980 264.400 39.330 265.000 ;
        RECT 43.880 264.450 45.580 266.750 ;
        RECT 46.530 266.600 50.480 266.800 ;
        RECT 50.130 266.000 50.480 266.600 ;
        RECT 46.530 265.800 50.480 266.000 ;
        RECT 50.130 265.200 50.480 265.800 ;
        RECT 46.530 265.000 50.480 265.200 ;
        RECT 38.980 264.200 42.930 264.400 ;
        RECT 38.980 263.600 39.330 264.200 ;
        RECT 38.980 263.400 42.930 263.600 ;
        RECT 38.980 262.800 39.330 263.400 ;
        RECT 38.980 262.600 42.930 262.800 ;
        RECT 38.980 262.000 39.330 262.600 ;
        RECT 26.530 261.400 42.930 262.000 ;
        RECT 29.180 260.800 31.480 260.850 ;
        RECT 37.980 260.800 40.280 260.850 ;
        RECT 43.930 260.800 44.330 264.450 ;
        RECT 25.130 260.400 44.330 260.800 ;
        RECT 45.130 260.800 45.530 264.450 ;
        RECT 50.130 264.400 50.480 265.000 ;
        RECT 46.530 264.200 50.480 264.400 ;
        RECT 50.130 263.600 50.480 264.200 ;
        RECT 46.530 263.400 50.480 263.600 ;
        RECT 50.130 262.800 50.480 263.400 ;
        RECT 46.530 262.600 50.480 262.800 ;
        RECT 50.130 262.000 50.480 262.600 ;
        RECT 51.080 262.000 51.280 269.600 ;
        RECT 51.880 262.000 52.080 269.600 ;
        RECT 52.680 262.000 52.880 269.600 ;
        RECT 53.480 262.000 53.680 269.600 ;
        RECT 54.280 262.000 55.180 278.000 ;
        RECT 55.780 270.400 55.980 278.000 ;
        RECT 56.580 270.400 56.780 278.000 ;
        RECT 57.380 270.400 57.580 278.000 ;
        RECT 58.180 270.400 58.380 278.000 ;
        RECT 58.980 277.400 59.330 278.000 ;
        RECT 58.980 277.200 62.930 277.400 ;
        RECT 58.980 276.600 59.330 277.200 ;
        RECT 58.980 276.400 62.930 276.600 ;
        RECT 58.980 275.800 59.330 276.400 ;
        RECT 58.980 275.600 62.930 275.800 ;
        RECT 58.980 275.000 59.330 275.600 ;
        RECT 63.930 275.550 64.330 279.200 ;
        RECT 65.130 279.200 84.330 279.600 ;
        RECT 65.130 275.550 65.530 279.200 ;
        RECT 69.180 279.150 71.480 279.200 ;
        RECT 77.980 279.150 80.280 279.200 ;
        RECT 66.530 278.000 82.930 278.600 ;
        RECT 70.130 277.400 70.480 278.000 ;
        RECT 66.530 277.200 70.480 277.400 ;
        RECT 70.130 276.600 70.480 277.200 ;
        RECT 66.530 276.400 70.480 276.600 ;
        RECT 70.130 275.800 70.480 276.400 ;
        RECT 66.530 275.600 70.480 275.800 ;
        RECT 58.980 274.800 62.930 275.000 ;
        RECT 58.980 274.200 59.330 274.800 ;
        RECT 58.980 274.000 62.930 274.200 ;
        RECT 58.980 273.400 59.330 274.000 ;
        RECT 58.980 273.200 62.930 273.400 ;
        RECT 63.880 273.250 65.580 275.550 ;
        RECT 70.130 275.000 70.480 275.600 ;
        RECT 66.530 274.800 70.480 275.000 ;
        RECT 70.130 274.200 70.480 274.800 ;
        RECT 66.530 274.000 70.480 274.200 ;
        RECT 70.130 273.400 70.480 274.000 ;
        RECT 58.980 272.600 59.330 273.200 ;
        RECT 58.980 272.400 62.930 272.600 ;
        RECT 58.980 271.800 59.330 272.400 ;
        RECT 58.980 271.600 62.930 271.800 ;
        RECT 58.980 271.000 59.330 271.600 ;
        RECT 58.980 270.800 62.930 271.000 ;
        RECT 58.980 270.400 59.330 270.800 ;
        RECT 55.780 262.000 55.980 269.600 ;
        RECT 56.580 262.000 56.780 269.600 ;
        RECT 57.380 262.000 57.580 269.600 ;
        RECT 58.180 262.000 58.380 269.600 ;
        RECT 58.980 269.200 59.330 269.600 ;
        RECT 58.980 269.000 62.930 269.200 ;
        RECT 58.980 268.400 59.330 269.000 ;
        RECT 58.980 268.200 62.930 268.400 ;
        RECT 58.980 267.600 59.330 268.200 ;
        RECT 58.980 267.400 62.930 267.600 ;
        RECT 58.980 266.800 59.330 267.400 ;
        RECT 58.980 266.600 62.930 266.800 ;
        RECT 63.930 266.750 64.330 273.250 ;
        RECT 65.130 266.750 65.530 273.250 ;
        RECT 66.530 273.200 70.480 273.400 ;
        RECT 70.130 272.600 70.480 273.200 ;
        RECT 66.530 272.400 70.480 272.600 ;
        RECT 70.130 271.800 70.480 272.400 ;
        RECT 66.530 271.600 70.480 271.800 ;
        RECT 70.130 271.000 70.480 271.600 ;
        RECT 66.530 270.800 70.480 271.000 ;
        RECT 70.130 270.400 70.480 270.800 ;
        RECT 71.080 270.400 71.280 278.000 ;
        RECT 71.880 270.400 72.080 278.000 ;
        RECT 72.680 270.400 72.880 278.000 ;
        RECT 73.480 270.400 73.680 278.000 ;
        RECT 70.130 269.200 70.480 269.600 ;
        RECT 66.530 269.000 70.480 269.200 ;
        RECT 70.130 268.400 70.480 269.000 ;
        RECT 66.530 268.200 70.480 268.400 ;
        RECT 70.130 267.600 70.480 268.200 ;
        RECT 66.530 267.400 70.480 267.600 ;
        RECT 70.130 266.800 70.480 267.400 ;
        RECT 58.980 266.000 59.330 266.600 ;
        RECT 58.980 265.800 62.930 266.000 ;
        RECT 58.980 265.200 59.330 265.800 ;
        RECT 58.980 265.000 62.930 265.200 ;
        RECT 58.980 264.400 59.330 265.000 ;
        RECT 63.880 264.450 65.580 266.750 ;
        RECT 66.530 266.600 70.480 266.800 ;
        RECT 70.130 266.000 70.480 266.600 ;
        RECT 66.530 265.800 70.480 266.000 ;
        RECT 70.130 265.200 70.480 265.800 ;
        RECT 66.530 265.000 70.480 265.200 ;
        RECT 58.980 264.200 62.930 264.400 ;
        RECT 58.980 263.600 59.330 264.200 ;
        RECT 58.980 263.400 62.930 263.600 ;
        RECT 58.980 262.800 59.330 263.400 ;
        RECT 58.980 262.600 62.930 262.800 ;
        RECT 58.980 262.000 59.330 262.600 ;
        RECT 46.530 261.400 62.930 262.000 ;
        RECT 49.180 260.800 51.480 260.850 ;
        RECT 57.980 260.800 60.280 260.850 ;
        RECT 63.930 260.800 64.330 264.450 ;
        RECT 45.130 260.400 64.330 260.800 ;
        RECT 65.130 260.800 65.530 264.450 ;
        RECT 70.130 264.400 70.480 265.000 ;
        RECT 66.530 264.200 70.480 264.400 ;
        RECT 70.130 263.600 70.480 264.200 ;
        RECT 66.530 263.400 70.480 263.600 ;
        RECT 70.130 262.800 70.480 263.400 ;
        RECT 66.530 262.600 70.480 262.800 ;
        RECT 70.130 262.000 70.480 262.600 ;
        RECT 71.080 262.000 71.280 269.600 ;
        RECT 71.880 262.000 72.080 269.600 ;
        RECT 72.680 262.000 72.880 269.600 ;
        RECT 73.480 262.000 73.680 269.600 ;
        RECT 74.280 262.000 75.180 278.000 ;
        RECT 75.780 270.400 75.980 278.000 ;
        RECT 76.580 270.400 76.780 278.000 ;
        RECT 77.380 270.400 77.580 278.000 ;
        RECT 78.180 270.400 78.380 278.000 ;
        RECT 78.980 277.400 79.330 278.000 ;
        RECT 78.980 277.200 82.930 277.400 ;
        RECT 78.980 276.600 79.330 277.200 ;
        RECT 78.980 276.400 82.930 276.600 ;
        RECT 78.980 275.800 79.330 276.400 ;
        RECT 78.980 275.600 82.930 275.800 ;
        RECT 78.980 275.000 79.330 275.600 ;
        RECT 83.930 275.550 84.330 279.200 ;
        RECT 85.130 279.200 104.330 279.600 ;
        RECT 85.130 275.550 85.530 279.200 ;
        RECT 89.180 279.150 91.480 279.200 ;
        RECT 97.980 279.150 100.280 279.200 ;
        RECT 86.530 278.000 102.930 278.600 ;
        RECT 90.130 277.400 90.480 278.000 ;
        RECT 86.530 277.200 90.480 277.400 ;
        RECT 90.130 276.600 90.480 277.200 ;
        RECT 86.530 276.400 90.480 276.600 ;
        RECT 90.130 275.800 90.480 276.400 ;
        RECT 86.530 275.600 90.480 275.800 ;
        RECT 78.980 274.800 82.930 275.000 ;
        RECT 78.980 274.200 79.330 274.800 ;
        RECT 78.980 274.000 82.930 274.200 ;
        RECT 78.980 273.400 79.330 274.000 ;
        RECT 78.980 273.200 82.930 273.400 ;
        RECT 83.880 273.250 85.580 275.550 ;
        RECT 90.130 275.000 90.480 275.600 ;
        RECT 86.530 274.800 90.480 275.000 ;
        RECT 90.130 274.200 90.480 274.800 ;
        RECT 86.530 274.000 90.480 274.200 ;
        RECT 90.130 273.400 90.480 274.000 ;
        RECT 78.980 272.600 79.330 273.200 ;
        RECT 78.980 272.400 82.930 272.600 ;
        RECT 78.980 271.800 79.330 272.400 ;
        RECT 78.980 271.600 82.930 271.800 ;
        RECT 78.980 271.000 79.330 271.600 ;
        RECT 78.980 270.800 82.930 271.000 ;
        RECT 78.980 270.400 79.330 270.800 ;
        RECT 75.780 262.000 75.980 269.600 ;
        RECT 76.580 262.000 76.780 269.600 ;
        RECT 77.380 262.000 77.580 269.600 ;
        RECT 78.180 262.000 78.380 269.600 ;
        RECT 78.980 269.200 79.330 269.600 ;
        RECT 78.980 269.000 82.930 269.200 ;
        RECT 78.980 268.400 79.330 269.000 ;
        RECT 78.980 268.200 82.930 268.400 ;
        RECT 78.980 267.600 79.330 268.200 ;
        RECT 78.980 267.400 82.930 267.600 ;
        RECT 78.980 266.800 79.330 267.400 ;
        RECT 78.980 266.600 82.930 266.800 ;
        RECT 83.930 266.750 84.330 273.250 ;
        RECT 85.130 266.750 85.530 273.250 ;
        RECT 86.530 273.200 90.480 273.400 ;
        RECT 90.130 272.600 90.480 273.200 ;
        RECT 86.530 272.400 90.480 272.600 ;
        RECT 90.130 271.800 90.480 272.400 ;
        RECT 86.530 271.600 90.480 271.800 ;
        RECT 90.130 271.000 90.480 271.600 ;
        RECT 86.530 270.800 90.480 271.000 ;
        RECT 90.130 270.400 90.480 270.800 ;
        RECT 91.080 270.400 91.280 278.000 ;
        RECT 91.880 270.400 92.080 278.000 ;
        RECT 92.680 270.400 92.880 278.000 ;
        RECT 93.480 270.400 93.680 278.000 ;
        RECT 90.130 269.200 90.480 269.600 ;
        RECT 86.530 269.000 90.480 269.200 ;
        RECT 90.130 268.400 90.480 269.000 ;
        RECT 86.530 268.200 90.480 268.400 ;
        RECT 90.130 267.600 90.480 268.200 ;
        RECT 86.530 267.400 90.480 267.600 ;
        RECT 90.130 266.800 90.480 267.400 ;
        RECT 78.980 266.000 79.330 266.600 ;
        RECT 78.980 265.800 82.930 266.000 ;
        RECT 78.980 265.200 79.330 265.800 ;
        RECT 78.980 265.000 82.930 265.200 ;
        RECT 78.980 264.400 79.330 265.000 ;
        RECT 83.880 264.450 85.580 266.750 ;
        RECT 86.530 266.600 90.480 266.800 ;
        RECT 90.130 266.000 90.480 266.600 ;
        RECT 86.530 265.800 90.480 266.000 ;
        RECT 90.130 265.200 90.480 265.800 ;
        RECT 86.530 265.000 90.480 265.200 ;
        RECT 78.980 264.200 82.930 264.400 ;
        RECT 78.980 263.600 79.330 264.200 ;
        RECT 78.980 263.400 82.930 263.600 ;
        RECT 78.980 262.800 79.330 263.400 ;
        RECT 78.980 262.600 82.930 262.800 ;
        RECT 78.980 262.000 79.330 262.600 ;
        RECT 66.530 261.400 82.930 262.000 ;
        RECT 69.180 260.800 71.480 260.850 ;
        RECT 77.980 260.800 80.280 260.850 ;
        RECT 83.930 260.800 84.330 264.450 ;
        RECT 65.130 260.400 84.330 260.800 ;
        RECT 85.130 260.800 85.530 264.450 ;
        RECT 90.130 264.400 90.480 265.000 ;
        RECT 86.530 264.200 90.480 264.400 ;
        RECT 90.130 263.600 90.480 264.200 ;
        RECT 86.530 263.400 90.480 263.600 ;
        RECT 90.130 262.800 90.480 263.400 ;
        RECT 86.530 262.600 90.480 262.800 ;
        RECT 90.130 262.000 90.480 262.600 ;
        RECT 91.080 262.000 91.280 269.600 ;
        RECT 91.880 262.000 92.080 269.600 ;
        RECT 92.680 262.000 92.880 269.600 ;
        RECT 93.480 262.000 93.680 269.600 ;
        RECT 94.280 262.000 95.180 278.000 ;
        RECT 95.780 270.400 95.980 278.000 ;
        RECT 96.580 270.400 96.780 278.000 ;
        RECT 97.380 270.400 97.580 278.000 ;
        RECT 98.180 270.400 98.380 278.000 ;
        RECT 98.980 277.400 99.330 278.000 ;
        RECT 98.980 277.200 102.930 277.400 ;
        RECT 98.980 276.600 99.330 277.200 ;
        RECT 98.980 276.400 102.930 276.600 ;
        RECT 98.980 275.800 99.330 276.400 ;
        RECT 98.980 275.600 102.930 275.800 ;
        RECT 98.980 275.000 99.330 275.600 ;
        RECT 103.930 275.550 104.330 279.200 ;
        RECT 105.340 276.855 105.700 277.235 ;
        RECT 105.970 276.855 106.330 277.235 ;
        RECT 106.570 276.855 106.930 277.235 ;
        RECT 105.340 276.265 105.700 276.645 ;
        RECT 105.970 276.265 106.330 276.645 ;
        RECT 106.570 276.265 106.930 276.645 ;
        RECT 98.980 274.800 102.930 275.000 ;
        RECT 98.980 274.200 99.330 274.800 ;
        RECT 98.980 274.000 102.930 274.200 ;
        RECT 98.980 273.400 99.330 274.000 ;
        RECT 98.980 273.200 102.930 273.400 ;
        RECT 103.880 273.250 104.730 275.550 ;
        RECT 98.980 272.600 99.330 273.200 ;
        RECT 98.980 272.400 102.930 272.600 ;
        RECT 98.980 271.800 99.330 272.400 ;
        RECT 98.980 271.600 102.930 271.800 ;
        RECT 98.980 271.000 99.330 271.600 ;
        RECT 98.980 270.800 102.930 271.000 ;
        RECT 98.980 270.400 99.330 270.800 ;
        RECT 95.780 262.000 95.980 269.600 ;
        RECT 96.580 262.000 96.780 269.600 ;
        RECT 97.380 262.000 97.580 269.600 ;
        RECT 98.180 262.000 98.380 269.600 ;
        RECT 98.980 269.200 99.330 269.600 ;
        RECT 98.980 269.000 102.930 269.200 ;
        RECT 98.980 268.400 99.330 269.000 ;
        RECT 98.980 268.200 102.930 268.400 ;
        RECT 98.980 267.600 99.330 268.200 ;
        RECT 98.980 267.400 102.930 267.600 ;
        RECT 98.980 266.800 99.330 267.400 ;
        RECT 98.980 266.600 102.930 266.800 ;
        RECT 103.930 266.750 104.330 273.250 ;
        RECT 98.980 266.000 99.330 266.600 ;
        RECT 98.980 265.800 102.930 266.000 ;
        RECT 98.980 265.200 99.330 265.800 ;
        RECT 98.980 265.000 102.930 265.200 ;
        RECT 98.980 264.400 99.330 265.000 ;
        RECT 103.880 264.450 104.730 266.750 ;
        RECT 98.980 264.200 102.930 264.400 ;
        RECT 98.980 263.600 99.330 264.200 ;
        RECT 98.980 263.400 102.930 263.600 ;
        RECT 98.980 262.800 99.330 263.400 ;
        RECT 98.980 262.600 102.930 262.800 ;
        RECT 98.980 262.000 99.330 262.600 ;
        RECT 86.530 261.400 102.930 262.000 ;
        RECT 89.180 260.800 91.480 260.850 ;
        RECT 97.980 260.800 100.280 260.850 ;
        RECT 103.930 260.800 104.330 264.450 ;
        RECT 105.340 262.495 105.700 262.875 ;
        RECT 105.970 262.495 106.330 262.875 ;
        RECT 106.570 262.495 106.930 262.875 ;
        RECT 105.340 261.905 105.700 262.285 ;
        RECT 105.970 261.905 106.330 262.285 ;
        RECT 106.570 261.905 106.930 262.285 ;
        RECT 85.130 260.400 104.330 260.800 ;
        RECT 9.180 259.600 11.480 260.400 ;
        RECT 17.980 259.600 20.280 260.400 ;
        RECT 29.180 259.600 31.480 260.400 ;
        RECT 37.980 259.600 40.280 260.400 ;
        RECT 49.180 259.600 51.480 260.400 ;
        RECT 57.980 259.600 60.280 260.400 ;
        RECT 69.180 259.600 71.480 260.400 ;
        RECT 77.980 259.600 80.280 260.400 ;
        RECT 89.180 259.600 91.480 260.400 ;
        RECT 97.980 259.600 100.280 260.400 ;
        RECT 5.130 259.200 24.330 259.600 ;
        RECT 2.515 257.340 2.875 257.720 ;
        RECT 3.145 257.340 3.505 257.720 ;
        RECT 3.745 257.340 4.105 257.720 ;
        RECT 2.515 256.750 2.875 257.130 ;
        RECT 3.145 256.750 3.505 257.130 ;
        RECT 3.745 256.750 4.105 257.130 ;
        RECT 5.130 255.550 5.530 259.200 ;
        RECT 9.180 259.150 11.480 259.200 ;
        RECT 17.980 259.150 20.280 259.200 ;
        RECT 6.530 258.000 22.930 258.600 ;
        RECT 10.130 257.400 10.480 258.000 ;
        RECT 6.530 257.200 10.480 257.400 ;
        RECT 10.130 256.600 10.480 257.200 ;
        RECT 6.530 256.400 10.480 256.600 ;
        RECT 10.130 255.800 10.480 256.400 ;
        RECT 6.530 255.600 10.480 255.800 ;
        RECT 4.730 255.545 5.580 255.550 ;
        RECT 2.315 253.250 5.580 255.545 ;
        RECT 10.130 255.000 10.480 255.600 ;
        RECT 6.530 254.800 10.480 255.000 ;
        RECT 10.130 254.200 10.480 254.800 ;
        RECT 6.530 254.000 10.480 254.200 ;
        RECT 10.130 253.400 10.480 254.000 ;
        RECT 5.130 246.750 5.530 253.250 ;
        RECT 6.530 253.200 10.480 253.400 ;
        RECT 10.130 252.600 10.480 253.200 ;
        RECT 6.530 252.400 10.480 252.600 ;
        RECT 10.130 251.800 10.480 252.400 ;
        RECT 6.530 251.600 10.480 251.800 ;
        RECT 10.130 251.000 10.480 251.600 ;
        RECT 6.530 250.800 10.480 251.000 ;
        RECT 10.130 250.400 10.480 250.800 ;
        RECT 11.080 250.400 11.280 258.000 ;
        RECT 11.880 250.400 12.080 258.000 ;
        RECT 12.680 250.400 12.880 258.000 ;
        RECT 13.480 250.400 13.680 258.000 ;
        RECT 10.130 249.200 10.480 249.600 ;
        RECT 6.530 249.000 10.480 249.200 ;
        RECT 10.130 248.400 10.480 249.000 ;
        RECT 6.530 248.200 10.480 248.400 ;
        RECT 10.130 247.600 10.480 248.200 ;
        RECT 6.530 247.400 10.480 247.600 ;
        RECT 10.130 246.800 10.480 247.400 ;
        RECT 2.315 244.455 5.580 246.750 ;
        RECT 6.530 246.600 10.480 246.800 ;
        RECT 10.130 246.000 10.480 246.600 ;
        RECT 6.530 245.800 10.480 246.000 ;
        RECT 10.130 245.200 10.480 245.800 ;
        RECT 6.530 245.000 10.480 245.200 ;
        RECT 4.730 244.450 5.580 244.455 ;
        RECT 2.515 243.230 2.875 243.610 ;
        RECT 3.145 243.230 3.505 243.610 ;
        RECT 3.745 243.230 4.105 243.610 ;
        RECT 2.515 242.640 2.875 243.020 ;
        RECT 3.145 242.640 3.505 243.020 ;
        RECT 3.745 242.640 4.105 243.020 ;
        RECT 5.130 240.800 5.530 244.450 ;
        RECT 10.130 244.400 10.480 245.000 ;
        RECT 6.530 244.200 10.480 244.400 ;
        RECT 10.130 243.600 10.480 244.200 ;
        RECT 6.530 243.400 10.480 243.600 ;
        RECT 10.130 242.800 10.480 243.400 ;
        RECT 6.530 242.600 10.480 242.800 ;
        RECT 10.130 242.000 10.480 242.600 ;
        RECT 11.080 242.000 11.280 249.600 ;
        RECT 11.880 242.000 12.080 249.600 ;
        RECT 12.680 242.000 12.880 249.600 ;
        RECT 13.480 242.000 13.680 249.600 ;
        RECT 14.280 242.000 15.180 258.000 ;
        RECT 15.780 250.400 15.980 258.000 ;
        RECT 16.580 250.400 16.780 258.000 ;
        RECT 17.380 250.400 17.580 258.000 ;
        RECT 18.180 250.400 18.380 258.000 ;
        RECT 18.980 257.400 19.330 258.000 ;
        RECT 18.980 257.200 22.930 257.400 ;
        RECT 18.980 256.600 19.330 257.200 ;
        RECT 18.980 256.400 22.930 256.600 ;
        RECT 18.980 255.800 19.330 256.400 ;
        RECT 18.980 255.600 22.930 255.800 ;
        RECT 18.980 255.000 19.330 255.600 ;
        RECT 23.930 255.550 24.330 259.200 ;
        RECT 25.130 259.200 44.330 259.600 ;
        RECT 25.130 255.550 25.530 259.200 ;
        RECT 29.180 259.150 31.480 259.200 ;
        RECT 37.980 259.150 40.280 259.200 ;
        RECT 26.530 258.000 42.930 258.600 ;
        RECT 30.130 257.400 30.480 258.000 ;
        RECT 26.530 257.200 30.480 257.400 ;
        RECT 30.130 256.600 30.480 257.200 ;
        RECT 26.530 256.400 30.480 256.600 ;
        RECT 30.130 255.800 30.480 256.400 ;
        RECT 26.530 255.600 30.480 255.800 ;
        RECT 18.980 254.800 22.930 255.000 ;
        RECT 18.980 254.200 19.330 254.800 ;
        RECT 18.980 254.000 22.930 254.200 ;
        RECT 18.980 253.400 19.330 254.000 ;
        RECT 18.980 253.200 22.930 253.400 ;
        RECT 23.880 253.250 25.580 255.550 ;
        RECT 30.130 255.000 30.480 255.600 ;
        RECT 26.530 254.800 30.480 255.000 ;
        RECT 30.130 254.200 30.480 254.800 ;
        RECT 26.530 254.000 30.480 254.200 ;
        RECT 30.130 253.400 30.480 254.000 ;
        RECT 18.980 252.600 19.330 253.200 ;
        RECT 18.980 252.400 22.930 252.600 ;
        RECT 18.980 251.800 19.330 252.400 ;
        RECT 18.980 251.600 22.930 251.800 ;
        RECT 18.980 251.000 19.330 251.600 ;
        RECT 18.980 250.800 22.930 251.000 ;
        RECT 18.980 250.400 19.330 250.800 ;
        RECT 15.780 242.000 15.980 249.600 ;
        RECT 16.580 242.000 16.780 249.600 ;
        RECT 17.380 242.000 17.580 249.600 ;
        RECT 18.180 242.000 18.380 249.600 ;
        RECT 18.980 249.200 19.330 249.600 ;
        RECT 18.980 249.000 22.930 249.200 ;
        RECT 18.980 248.400 19.330 249.000 ;
        RECT 18.980 248.200 22.930 248.400 ;
        RECT 18.980 247.600 19.330 248.200 ;
        RECT 18.980 247.400 22.930 247.600 ;
        RECT 18.980 246.800 19.330 247.400 ;
        RECT 18.980 246.600 22.930 246.800 ;
        RECT 23.930 246.750 24.330 253.250 ;
        RECT 25.130 246.750 25.530 253.250 ;
        RECT 26.530 253.200 30.480 253.400 ;
        RECT 30.130 252.600 30.480 253.200 ;
        RECT 26.530 252.400 30.480 252.600 ;
        RECT 30.130 251.800 30.480 252.400 ;
        RECT 26.530 251.600 30.480 251.800 ;
        RECT 30.130 251.000 30.480 251.600 ;
        RECT 26.530 250.800 30.480 251.000 ;
        RECT 30.130 250.400 30.480 250.800 ;
        RECT 31.080 250.400 31.280 258.000 ;
        RECT 31.880 250.400 32.080 258.000 ;
        RECT 32.680 250.400 32.880 258.000 ;
        RECT 33.480 250.400 33.680 258.000 ;
        RECT 30.130 249.200 30.480 249.600 ;
        RECT 26.530 249.000 30.480 249.200 ;
        RECT 30.130 248.400 30.480 249.000 ;
        RECT 26.530 248.200 30.480 248.400 ;
        RECT 30.130 247.600 30.480 248.200 ;
        RECT 26.530 247.400 30.480 247.600 ;
        RECT 30.130 246.800 30.480 247.400 ;
        RECT 18.980 246.000 19.330 246.600 ;
        RECT 18.980 245.800 22.930 246.000 ;
        RECT 18.980 245.200 19.330 245.800 ;
        RECT 18.980 245.000 22.930 245.200 ;
        RECT 18.980 244.400 19.330 245.000 ;
        RECT 23.880 244.450 25.580 246.750 ;
        RECT 26.530 246.600 30.480 246.800 ;
        RECT 30.130 246.000 30.480 246.600 ;
        RECT 26.530 245.800 30.480 246.000 ;
        RECT 30.130 245.200 30.480 245.800 ;
        RECT 26.530 245.000 30.480 245.200 ;
        RECT 18.980 244.200 22.930 244.400 ;
        RECT 18.980 243.600 19.330 244.200 ;
        RECT 18.980 243.400 22.930 243.600 ;
        RECT 18.980 242.800 19.330 243.400 ;
        RECT 18.980 242.600 22.930 242.800 ;
        RECT 18.980 242.000 19.330 242.600 ;
        RECT 6.530 241.400 22.930 242.000 ;
        RECT 9.180 240.800 11.480 240.850 ;
        RECT 17.980 240.800 20.280 240.850 ;
        RECT 23.930 240.800 24.330 244.450 ;
        RECT 5.130 240.400 24.330 240.800 ;
        RECT 25.130 240.800 25.530 244.450 ;
        RECT 30.130 244.400 30.480 245.000 ;
        RECT 26.530 244.200 30.480 244.400 ;
        RECT 30.130 243.600 30.480 244.200 ;
        RECT 26.530 243.400 30.480 243.600 ;
        RECT 30.130 242.800 30.480 243.400 ;
        RECT 26.530 242.600 30.480 242.800 ;
        RECT 30.130 242.000 30.480 242.600 ;
        RECT 31.080 242.000 31.280 249.600 ;
        RECT 31.880 242.000 32.080 249.600 ;
        RECT 32.680 242.000 32.880 249.600 ;
        RECT 33.480 242.000 33.680 249.600 ;
        RECT 34.280 242.000 35.180 258.000 ;
        RECT 35.780 250.400 35.980 258.000 ;
        RECT 36.580 250.400 36.780 258.000 ;
        RECT 37.380 250.400 37.580 258.000 ;
        RECT 38.180 250.400 38.380 258.000 ;
        RECT 38.980 257.400 39.330 258.000 ;
        RECT 38.980 257.200 42.930 257.400 ;
        RECT 38.980 256.600 39.330 257.200 ;
        RECT 38.980 256.400 42.930 256.600 ;
        RECT 38.980 255.800 39.330 256.400 ;
        RECT 38.980 255.600 42.930 255.800 ;
        RECT 38.980 255.000 39.330 255.600 ;
        RECT 43.930 255.550 44.330 259.200 ;
        RECT 45.130 259.200 64.330 259.600 ;
        RECT 45.130 255.550 45.530 259.200 ;
        RECT 49.180 259.150 51.480 259.200 ;
        RECT 57.980 259.150 60.280 259.200 ;
        RECT 46.530 258.000 62.930 258.600 ;
        RECT 50.130 257.400 50.480 258.000 ;
        RECT 46.530 257.200 50.480 257.400 ;
        RECT 50.130 256.600 50.480 257.200 ;
        RECT 46.530 256.400 50.480 256.600 ;
        RECT 50.130 255.800 50.480 256.400 ;
        RECT 46.530 255.600 50.480 255.800 ;
        RECT 38.980 254.800 42.930 255.000 ;
        RECT 38.980 254.200 39.330 254.800 ;
        RECT 38.980 254.000 42.930 254.200 ;
        RECT 38.980 253.400 39.330 254.000 ;
        RECT 38.980 253.200 42.930 253.400 ;
        RECT 43.880 253.250 45.580 255.550 ;
        RECT 50.130 255.000 50.480 255.600 ;
        RECT 46.530 254.800 50.480 255.000 ;
        RECT 50.130 254.200 50.480 254.800 ;
        RECT 46.530 254.000 50.480 254.200 ;
        RECT 50.130 253.400 50.480 254.000 ;
        RECT 38.980 252.600 39.330 253.200 ;
        RECT 38.980 252.400 42.930 252.600 ;
        RECT 38.980 251.800 39.330 252.400 ;
        RECT 38.980 251.600 42.930 251.800 ;
        RECT 38.980 251.000 39.330 251.600 ;
        RECT 38.980 250.800 42.930 251.000 ;
        RECT 38.980 250.400 39.330 250.800 ;
        RECT 35.780 242.000 35.980 249.600 ;
        RECT 36.580 242.000 36.780 249.600 ;
        RECT 37.380 242.000 37.580 249.600 ;
        RECT 38.180 242.000 38.380 249.600 ;
        RECT 38.980 249.200 39.330 249.600 ;
        RECT 38.980 249.000 42.930 249.200 ;
        RECT 38.980 248.400 39.330 249.000 ;
        RECT 38.980 248.200 42.930 248.400 ;
        RECT 38.980 247.600 39.330 248.200 ;
        RECT 38.980 247.400 42.930 247.600 ;
        RECT 38.980 246.800 39.330 247.400 ;
        RECT 38.980 246.600 42.930 246.800 ;
        RECT 43.930 246.750 44.330 253.250 ;
        RECT 45.130 246.750 45.530 253.250 ;
        RECT 46.530 253.200 50.480 253.400 ;
        RECT 50.130 252.600 50.480 253.200 ;
        RECT 46.530 252.400 50.480 252.600 ;
        RECT 50.130 251.800 50.480 252.400 ;
        RECT 46.530 251.600 50.480 251.800 ;
        RECT 50.130 251.000 50.480 251.600 ;
        RECT 46.530 250.800 50.480 251.000 ;
        RECT 50.130 250.400 50.480 250.800 ;
        RECT 51.080 250.400 51.280 258.000 ;
        RECT 51.880 250.400 52.080 258.000 ;
        RECT 52.680 250.400 52.880 258.000 ;
        RECT 53.480 250.400 53.680 258.000 ;
        RECT 50.130 249.200 50.480 249.600 ;
        RECT 46.530 249.000 50.480 249.200 ;
        RECT 50.130 248.400 50.480 249.000 ;
        RECT 46.530 248.200 50.480 248.400 ;
        RECT 50.130 247.600 50.480 248.200 ;
        RECT 46.530 247.400 50.480 247.600 ;
        RECT 50.130 246.800 50.480 247.400 ;
        RECT 38.980 246.000 39.330 246.600 ;
        RECT 38.980 245.800 42.930 246.000 ;
        RECT 38.980 245.200 39.330 245.800 ;
        RECT 38.980 245.000 42.930 245.200 ;
        RECT 38.980 244.400 39.330 245.000 ;
        RECT 43.880 244.450 45.580 246.750 ;
        RECT 46.530 246.600 50.480 246.800 ;
        RECT 50.130 246.000 50.480 246.600 ;
        RECT 46.530 245.800 50.480 246.000 ;
        RECT 50.130 245.200 50.480 245.800 ;
        RECT 46.530 245.000 50.480 245.200 ;
        RECT 38.980 244.200 42.930 244.400 ;
        RECT 38.980 243.600 39.330 244.200 ;
        RECT 38.980 243.400 42.930 243.600 ;
        RECT 38.980 242.800 39.330 243.400 ;
        RECT 38.980 242.600 42.930 242.800 ;
        RECT 38.980 242.000 39.330 242.600 ;
        RECT 26.530 241.400 42.930 242.000 ;
        RECT 29.180 240.800 31.480 240.850 ;
        RECT 37.980 240.800 40.280 240.850 ;
        RECT 43.930 240.800 44.330 244.450 ;
        RECT 25.130 240.400 44.330 240.800 ;
        RECT 45.130 240.800 45.530 244.450 ;
        RECT 50.130 244.400 50.480 245.000 ;
        RECT 46.530 244.200 50.480 244.400 ;
        RECT 50.130 243.600 50.480 244.200 ;
        RECT 46.530 243.400 50.480 243.600 ;
        RECT 50.130 242.800 50.480 243.400 ;
        RECT 46.530 242.600 50.480 242.800 ;
        RECT 50.130 242.000 50.480 242.600 ;
        RECT 51.080 242.000 51.280 249.600 ;
        RECT 51.880 242.000 52.080 249.600 ;
        RECT 52.680 242.000 52.880 249.600 ;
        RECT 53.480 242.000 53.680 249.600 ;
        RECT 54.280 242.000 55.180 258.000 ;
        RECT 55.780 250.400 55.980 258.000 ;
        RECT 56.580 250.400 56.780 258.000 ;
        RECT 57.380 250.400 57.580 258.000 ;
        RECT 58.180 250.400 58.380 258.000 ;
        RECT 58.980 257.400 59.330 258.000 ;
        RECT 58.980 257.200 62.930 257.400 ;
        RECT 58.980 256.600 59.330 257.200 ;
        RECT 58.980 256.400 62.930 256.600 ;
        RECT 58.980 255.800 59.330 256.400 ;
        RECT 58.980 255.600 62.930 255.800 ;
        RECT 58.980 255.000 59.330 255.600 ;
        RECT 63.930 255.550 64.330 259.200 ;
        RECT 65.130 259.200 84.330 259.600 ;
        RECT 65.130 255.550 65.530 259.200 ;
        RECT 69.180 259.150 71.480 259.200 ;
        RECT 77.980 259.150 80.280 259.200 ;
        RECT 66.530 258.000 82.930 258.600 ;
        RECT 70.130 257.400 70.480 258.000 ;
        RECT 66.530 257.200 70.480 257.400 ;
        RECT 70.130 256.600 70.480 257.200 ;
        RECT 66.530 256.400 70.480 256.600 ;
        RECT 70.130 255.800 70.480 256.400 ;
        RECT 66.530 255.600 70.480 255.800 ;
        RECT 58.980 254.800 62.930 255.000 ;
        RECT 58.980 254.200 59.330 254.800 ;
        RECT 58.980 254.000 62.930 254.200 ;
        RECT 58.980 253.400 59.330 254.000 ;
        RECT 58.980 253.200 62.930 253.400 ;
        RECT 63.880 253.250 65.580 255.550 ;
        RECT 70.130 255.000 70.480 255.600 ;
        RECT 66.530 254.800 70.480 255.000 ;
        RECT 70.130 254.200 70.480 254.800 ;
        RECT 66.530 254.000 70.480 254.200 ;
        RECT 70.130 253.400 70.480 254.000 ;
        RECT 58.980 252.600 59.330 253.200 ;
        RECT 58.980 252.400 62.930 252.600 ;
        RECT 58.980 251.800 59.330 252.400 ;
        RECT 58.980 251.600 62.930 251.800 ;
        RECT 58.980 251.000 59.330 251.600 ;
        RECT 58.980 250.800 62.930 251.000 ;
        RECT 58.980 250.400 59.330 250.800 ;
        RECT 55.780 242.000 55.980 249.600 ;
        RECT 56.580 242.000 56.780 249.600 ;
        RECT 57.380 242.000 57.580 249.600 ;
        RECT 58.180 242.000 58.380 249.600 ;
        RECT 58.980 249.200 59.330 249.600 ;
        RECT 58.980 249.000 62.930 249.200 ;
        RECT 58.980 248.400 59.330 249.000 ;
        RECT 58.980 248.200 62.930 248.400 ;
        RECT 58.980 247.600 59.330 248.200 ;
        RECT 58.980 247.400 62.930 247.600 ;
        RECT 58.980 246.800 59.330 247.400 ;
        RECT 58.980 246.600 62.930 246.800 ;
        RECT 63.930 246.750 64.330 253.250 ;
        RECT 65.130 246.750 65.530 253.250 ;
        RECT 66.530 253.200 70.480 253.400 ;
        RECT 70.130 252.600 70.480 253.200 ;
        RECT 66.530 252.400 70.480 252.600 ;
        RECT 70.130 251.800 70.480 252.400 ;
        RECT 66.530 251.600 70.480 251.800 ;
        RECT 70.130 251.000 70.480 251.600 ;
        RECT 66.530 250.800 70.480 251.000 ;
        RECT 70.130 250.400 70.480 250.800 ;
        RECT 71.080 250.400 71.280 258.000 ;
        RECT 71.880 250.400 72.080 258.000 ;
        RECT 72.680 250.400 72.880 258.000 ;
        RECT 73.480 250.400 73.680 258.000 ;
        RECT 70.130 249.200 70.480 249.600 ;
        RECT 66.530 249.000 70.480 249.200 ;
        RECT 70.130 248.400 70.480 249.000 ;
        RECT 66.530 248.200 70.480 248.400 ;
        RECT 70.130 247.600 70.480 248.200 ;
        RECT 66.530 247.400 70.480 247.600 ;
        RECT 70.130 246.800 70.480 247.400 ;
        RECT 58.980 246.000 59.330 246.600 ;
        RECT 58.980 245.800 62.930 246.000 ;
        RECT 58.980 245.200 59.330 245.800 ;
        RECT 58.980 245.000 62.930 245.200 ;
        RECT 58.980 244.400 59.330 245.000 ;
        RECT 63.880 244.450 65.580 246.750 ;
        RECT 66.530 246.600 70.480 246.800 ;
        RECT 70.130 246.000 70.480 246.600 ;
        RECT 66.530 245.800 70.480 246.000 ;
        RECT 70.130 245.200 70.480 245.800 ;
        RECT 66.530 245.000 70.480 245.200 ;
        RECT 58.980 244.200 62.930 244.400 ;
        RECT 58.980 243.600 59.330 244.200 ;
        RECT 58.980 243.400 62.930 243.600 ;
        RECT 58.980 242.800 59.330 243.400 ;
        RECT 58.980 242.600 62.930 242.800 ;
        RECT 58.980 242.000 59.330 242.600 ;
        RECT 46.530 241.400 62.930 242.000 ;
        RECT 49.180 240.800 51.480 240.850 ;
        RECT 57.980 240.800 60.280 240.850 ;
        RECT 63.930 240.800 64.330 244.450 ;
        RECT 45.130 240.400 64.330 240.800 ;
        RECT 65.130 240.800 65.530 244.450 ;
        RECT 70.130 244.400 70.480 245.000 ;
        RECT 66.530 244.200 70.480 244.400 ;
        RECT 70.130 243.600 70.480 244.200 ;
        RECT 66.530 243.400 70.480 243.600 ;
        RECT 70.130 242.800 70.480 243.400 ;
        RECT 66.530 242.600 70.480 242.800 ;
        RECT 70.130 242.000 70.480 242.600 ;
        RECT 71.080 242.000 71.280 249.600 ;
        RECT 71.880 242.000 72.080 249.600 ;
        RECT 72.680 242.000 72.880 249.600 ;
        RECT 73.480 242.000 73.680 249.600 ;
        RECT 74.280 242.000 75.180 258.000 ;
        RECT 75.780 250.400 75.980 258.000 ;
        RECT 76.580 250.400 76.780 258.000 ;
        RECT 77.380 250.400 77.580 258.000 ;
        RECT 78.180 250.400 78.380 258.000 ;
        RECT 78.980 257.400 79.330 258.000 ;
        RECT 78.980 257.200 82.930 257.400 ;
        RECT 78.980 256.600 79.330 257.200 ;
        RECT 78.980 256.400 82.930 256.600 ;
        RECT 78.980 255.800 79.330 256.400 ;
        RECT 78.980 255.600 82.930 255.800 ;
        RECT 78.980 255.000 79.330 255.600 ;
        RECT 83.930 255.550 84.330 259.200 ;
        RECT 85.130 259.200 104.330 259.600 ;
        RECT 85.130 255.550 85.530 259.200 ;
        RECT 89.180 259.150 91.480 259.200 ;
        RECT 97.980 259.150 100.280 259.200 ;
        RECT 86.530 258.000 102.930 258.600 ;
        RECT 90.130 257.400 90.480 258.000 ;
        RECT 86.530 257.200 90.480 257.400 ;
        RECT 90.130 256.600 90.480 257.200 ;
        RECT 86.530 256.400 90.480 256.600 ;
        RECT 90.130 255.800 90.480 256.400 ;
        RECT 86.530 255.600 90.480 255.800 ;
        RECT 78.980 254.800 82.930 255.000 ;
        RECT 78.980 254.200 79.330 254.800 ;
        RECT 78.980 254.000 82.930 254.200 ;
        RECT 78.980 253.400 79.330 254.000 ;
        RECT 78.980 253.200 82.930 253.400 ;
        RECT 83.880 253.250 85.580 255.550 ;
        RECT 90.130 255.000 90.480 255.600 ;
        RECT 86.530 254.800 90.480 255.000 ;
        RECT 90.130 254.200 90.480 254.800 ;
        RECT 86.530 254.000 90.480 254.200 ;
        RECT 90.130 253.400 90.480 254.000 ;
        RECT 78.980 252.600 79.330 253.200 ;
        RECT 78.980 252.400 82.930 252.600 ;
        RECT 78.980 251.800 79.330 252.400 ;
        RECT 78.980 251.600 82.930 251.800 ;
        RECT 78.980 251.000 79.330 251.600 ;
        RECT 78.980 250.800 82.930 251.000 ;
        RECT 78.980 250.400 79.330 250.800 ;
        RECT 75.780 242.000 75.980 249.600 ;
        RECT 76.580 242.000 76.780 249.600 ;
        RECT 77.380 242.000 77.580 249.600 ;
        RECT 78.180 242.000 78.380 249.600 ;
        RECT 78.980 249.200 79.330 249.600 ;
        RECT 78.980 249.000 82.930 249.200 ;
        RECT 78.980 248.400 79.330 249.000 ;
        RECT 78.980 248.200 82.930 248.400 ;
        RECT 78.980 247.600 79.330 248.200 ;
        RECT 78.980 247.400 82.930 247.600 ;
        RECT 78.980 246.800 79.330 247.400 ;
        RECT 78.980 246.600 82.930 246.800 ;
        RECT 83.930 246.750 84.330 253.250 ;
        RECT 85.130 246.750 85.530 253.250 ;
        RECT 86.530 253.200 90.480 253.400 ;
        RECT 90.130 252.600 90.480 253.200 ;
        RECT 86.530 252.400 90.480 252.600 ;
        RECT 90.130 251.800 90.480 252.400 ;
        RECT 86.530 251.600 90.480 251.800 ;
        RECT 90.130 251.000 90.480 251.600 ;
        RECT 86.530 250.800 90.480 251.000 ;
        RECT 90.130 250.400 90.480 250.800 ;
        RECT 91.080 250.400 91.280 258.000 ;
        RECT 91.880 250.400 92.080 258.000 ;
        RECT 92.680 250.400 92.880 258.000 ;
        RECT 93.480 250.400 93.680 258.000 ;
        RECT 90.130 249.200 90.480 249.600 ;
        RECT 86.530 249.000 90.480 249.200 ;
        RECT 90.130 248.400 90.480 249.000 ;
        RECT 86.530 248.200 90.480 248.400 ;
        RECT 90.130 247.600 90.480 248.200 ;
        RECT 86.530 247.400 90.480 247.600 ;
        RECT 90.130 246.800 90.480 247.400 ;
        RECT 78.980 246.000 79.330 246.600 ;
        RECT 78.980 245.800 82.930 246.000 ;
        RECT 78.980 245.200 79.330 245.800 ;
        RECT 78.980 245.000 82.930 245.200 ;
        RECT 78.980 244.400 79.330 245.000 ;
        RECT 83.880 244.450 85.580 246.750 ;
        RECT 86.530 246.600 90.480 246.800 ;
        RECT 90.130 246.000 90.480 246.600 ;
        RECT 86.530 245.800 90.480 246.000 ;
        RECT 90.130 245.200 90.480 245.800 ;
        RECT 86.530 245.000 90.480 245.200 ;
        RECT 78.980 244.200 82.930 244.400 ;
        RECT 78.980 243.600 79.330 244.200 ;
        RECT 78.980 243.400 82.930 243.600 ;
        RECT 78.980 242.800 79.330 243.400 ;
        RECT 78.980 242.600 82.930 242.800 ;
        RECT 78.980 242.000 79.330 242.600 ;
        RECT 66.530 241.400 82.930 242.000 ;
        RECT 69.180 240.800 71.480 240.850 ;
        RECT 77.980 240.800 80.280 240.850 ;
        RECT 83.930 240.800 84.330 244.450 ;
        RECT 65.130 240.400 84.330 240.800 ;
        RECT 85.130 240.800 85.530 244.450 ;
        RECT 90.130 244.400 90.480 245.000 ;
        RECT 86.530 244.200 90.480 244.400 ;
        RECT 90.130 243.600 90.480 244.200 ;
        RECT 86.530 243.400 90.480 243.600 ;
        RECT 90.130 242.800 90.480 243.400 ;
        RECT 86.530 242.600 90.480 242.800 ;
        RECT 90.130 242.000 90.480 242.600 ;
        RECT 91.080 242.000 91.280 249.600 ;
        RECT 91.880 242.000 92.080 249.600 ;
        RECT 92.680 242.000 92.880 249.600 ;
        RECT 93.480 242.000 93.680 249.600 ;
        RECT 94.280 242.000 95.180 258.000 ;
        RECT 95.780 250.400 95.980 258.000 ;
        RECT 96.580 250.400 96.780 258.000 ;
        RECT 97.380 250.400 97.580 258.000 ;
        RECT 98.180 250.400 98.380 258.000 ;
        RECT 98.980 257.400 99.330 258.000 ;
        RECT 98.980 257.200 102.930 257.400 ;
        RECT 98.980 256.600 99.330 257.200 ;
        RECT 98.980 256.400 102.930 256.600 ;
        RECT 98.980 255.800 99.330 256.400 ;
        RECT 98.980 255.600 102.930 255.800 ;
        RECT 98.980 255.000 99.330 255.600 ;
        RECT 103.930 255.550 104.330 259.200 ;
        RECT 105.340 256.820 105.700 257.200 ;
        RECT 105.970 256.820 106.330 257.200 ;
        RECT 106.570 256.820 106.930 257.200 ;
        RECT 105.340 256.230 105.700 256.610 ;
        RECT 105.970 256.230 106.330 256.610 ;
        RECT 106.570 256.230 106.930 256.610 ;
        RECT 98.980 254.800 102.930 255.000 ;
        RECT 98.980 254.200 99.330 254.800 ;
        RECT 98.980 254.000 102.930 254.200 ;
        RECT 98.980 253.400 99.330 254.000 ;
        RECT 98.980 253.200 102.930 253.400 ;
        RECT 103.880 253.250 104.730 255.550 ;
        RECT 98.980 252.600 99.330 253.200 ;
        RECT 98.980 252.400 102.930 252.600 ;
        RECT 98.980 251.800 99.330 252.400 ;
        RECT 98.980 251.600 102.930 251.800 ;
        RECT 98.980 251.000 99.330 251.600 ;
        RECT 98.980 250.800 102.930 251.000 ;
        RECT 98.980 250.400 99.330 250.800 ;
        RECT 95.780 242.000 95.980 249.600 ;
        RECT 96.580 242.000 96.780 249.600 ;
        RECT 97.380 242.000 97.580 249.600 ;
        RECT 98.180 242.000 98.380 249.600 ;
        RECT 98.980 249.200 99.330 249.600 ;
        RECT 98.980 249.000 102.930 249.200 ;
        RECT 98.980 248.400 99.330 249.000 ;
        RECT 98.980 248.200 102.930 248.400 ;
        RECT 98.980 247.600 99.330 248.200 ;
        RECT 98.980 247.400 102.930 247.600 ;
        RECT 98.980 246.800 99.330 247.400 ;
        RECT 98.980 246.600 102.930 246.800 ;
        RECT 103.930 246.750 104.330 253.250 ;
        RECT 98.980 246.000 99.330 246.600 ;
        RECT 98.980 245.800 102.930 246.000 ;
        RECT 98.980 245.200 99.330 245.800 ;
        RECT 98.980 245.000 102.930 245.200 ;
        RECT 98.980 244.400 99.330 245.000 ;
        RECT 103.880 244.450 104.730 246.750 ;
        RECT 98.980 244.200 102.930 244.400 ;
        RECT 98.980 243.600 99.330 244.200 ;
        RECT 98.980 243.400 102.930 243.600 ;
        RECT 98.980 242.800 99.330 243.400 ;
        RECT 98.980 242.600 102.930 242.800 ;
        RECT 98.980 242.000 99.330 242.600 ;
        RECT 86.530 241.400 102.930 242.000 ;
        RECT 89.180 240.800 91.480 240.850 ;
        RECT 97.980 240.800 100.280 240.850 ;
        RECT 103.930 240.800 104.330 244.450 ;
        RECT 105.340 243.025 105.700 243.405 ;
        RECT 105.970 243.025 106.330 243.405 ;
        RECT 106.570 243.025 106.930 243.405 ;
        RECT 105.340 242.435 105.700 242.815 ;
        RECT 105.970 242.435 106.330 242.815 ;
        RECT 106.570 242.435 106.930 242.815 ;
        RECT 85.130 240.400 104.330 240.800 ;
        RECT 9.180 239.600 11.480 240.400 ;
        RECT 17.980 239.600 20.280 240.400 ;
        RECT 29.180 239.600 31.480 240.400 ;
        RECT 37.980 239.600 40.280 240.400 ;
        RECT 49.180 239.600 51.480 240.400 ;
        RECT 57.980 239.600 60.280 240.400 ;
        RECT 69.180 239.600 71.480 240.400 ;
        RECT 77.980 239.600 80.280 240.400 ;
        RECT 89.180 239.600 91.480 240.400 ;
        RECT 97.980 239.600 100.280 240.400 ;
        RECT 5.130 239.200 24.330 239.600 ;
        RECT 2.515 237.465 2.875 237.845 ;
        RECT 3.145 237.465 3.505 237.845 ;
        RECT 3.745 237.465 4.105 237.845 ;
        RECT 2.515 236.875 2.875 237.255 ;
        RECT 3.145 236.875 3.505 237.255 ;
        RECT 3.745 236.875 4.105 237.255 ;
        RECT 5.130 235.550 5.530 239.200 ;
        RECT 9.180 239.150 11.480 239.200 ;
        RECT 17.980 239.150 20.280 239.200 ;
        RECT 6.530 238.000 22.930 238.600 ;
        RECT 10.130 237.400 10.480 238.000 ;
        RECT 6.530 237.200 10.480 237.400 ;
        RECT 10.130 236.600 10.480 237.200 ;
        RECT 6.530 236.400 10.480 236.600 ;
        RECT 10.130 235.800 10.480 236.400 ;
        RECT 6.530 235.600 10.480 235.800 ;
        RECT 4.730 235.545 5.580 235.550 ;
        RECT 2.315 233.250 5.580 235.545 ;
        RECT 10.130 235.000 10.480 235.600 ;
        RECT 6.530 234.800 10.480 235.000 ;
        RECT 10.130 234.200 10.480 234.800 ;
        RECT 6.530 234.000 10.480 234.200 ;
        RECT 10.130 233.400 10.480 234.000 ;
        RECT 5.130 226.750 5.530 233.250 ;
        RECT 6.530 233.200 10.480 233.400 ;
        RECT 10.130 232.600 10.480 233.200 ;
        RECT 6.530 232.400 10.480 232.600 ;
        RECT 10.130 231.800 10.480 232.400 ;
        RECT 6.530 231.600 10.480 231.800 ;
        RECT 10.130 231.000 10.480 231.600 ;
        RECT 6.530 230.800 10.480 231.000 ;
        RECT 10.130 230.400 10.480 230.800 ;
        RECT 11.080 230.400 11.280 238.000 ;
        RECT 11.880 230.400 12.080 238.000 ;
        RECT 12.680 230.400 12.880 238.000 ;
        RECT 13.480 230.400 13.680 238.000 ;
        RECT 10.130 229.200 10.480 229.600 ;
        RECT 6.530 229.000 10.480 229.200 ;
        RECT 10.130 228.400 10.480 229.000 ;
        RECT 6.530 228.200 10.480 228.400 ;
        RECT 10.130 227.600 10.480 228.200 ;
        RECT 6.530 227.400 10.480 227.600 ;
        RECT 10.130 226.800 10.480 227.400 ;
        RECT 2.315 224.455 5.580 226.750 ;
        RECT 6.530 226.600 10.480 226.800 ;
        RECT 10.130 226.000 10.480 226.600 ;
        RECT 6.530 225.800 10.480 226.000 ;
        RECT 10.130 225.200 10.480 225.800 ;
        RECT 6.530 225.000 10.480 225.200 ;
        RECT 2.315 224.450 4.180 224.455 ;
        RECT 4.730 224.450 5.580 224.455 ;
        RECT 2.515 222.165 2.875 222.545 ;
        RECT 3.145 222.165 3.505 222.545 ;
        RECT 3.745 222.165 4.105 222.545 ;
        RECT 2.515 221.575 2.875 221.955 ;
        RECT 3.145 221.575 3.505 221.955 ;
        RECT 3.745 221.575 4.105 221.955 ;
        RECT 5.130 220.800 5.530 224.450 ;
        RECT 10.130 224.400 10.480 225.000 ;
        RECT 6.530 224.200 10.480 224.400 ;
        RECT 10.130 223.600 10.480 224.200 ;
        RECT 6.530 223.400 10.480 223.600 ;
        RECT 10.130 222.800 10.480 223.400 ;
        RECT 6.530 222.600 10.480 222.800 ;
        RECT 10.130 222.000 10.480 222.600 ;
        RECT 11.080 222.000 11.280 229.600 ;
        RECT 11.880 222.000 12.080 229.600 ;
        RECT 12.680 222.000 12.880 229.600 ;
        RECT 13.480 222.000 13.680 229.600 ;
        RECT 14.280 222.000 15.180 238.000 ;
        RECT 15.780 230.400 15.980 238.000 ;
        RECT 16.580 230.400 16.780 238.000 ;
        RECT 17.380 230.400 17.580 238.000 ;
        RECT 18.180 230.400 18.380 238.000 ;
        RECT 18.980 237.400 19.330 238.000 ;
        RECT 18.980 237.200 22.930 237.400 ;
        RECT 18.980 236.600 19.330 237.200 ;
        RECT 18.980 236.400 22.930 236.600 ;
        RECT 18.980 235.800 19.330 236.400 ;
        RECT 18.980 235.600 22.930 235.800 ;
        RECT 18.980 235.000 19.330 235.600 ;
        RECT 23.930 235.550 24.330 239.200 ;
        RECT 25.130 239.200 44.330 239.600 ;
        RECT 25.130 235.550 25.530 239.200 ;
        RECT 29.180 239.150 31.480 239.200 ;
        RECT 37.980 239.150 40.280 239.200 ;
        RECT 26.530 238.000 42.930 238.600 ;
        RECT 30.130 237.400 30.480 238.000 ;
        RECT 26.530 237.200 30.480 237.400 ;
        RECT 30.130 236.600 30.480 237.200 ;
        RECT 26.530 236.400 30.480 236.600 ;
        RECT 30.130 235.800 30.480 236.400 ;
        RECT 26.530 235.600 30.480 235.800 ;
        RECT 18.980 234.800 22.930 235.000 ;
        RECT 18.980 234.200 19.330 234.800 ;
        RECT 18.980 234.000 22.930 234.200 ;
        RECT 18.980 233.400 19.330 234.000 ;
        RECT 18.980 233.200 22.930 233.400 ;
        RECT 23.880 233.250 25.580 235.550 ;
        RECT 30.130 235.000 30.480 235.600 ;
        RECT 26.530 234.800 30.480 235.000 ;
        RECT 30.130 234.200 30.480 234.800 ;
        RECT 26.530 234.000 30.480 234.200 ;
        RECT 30.130 233.400 30.480 234.000 ;
        RECT 18.980 232.600 19.330 233.200 ;
        RECT 18.980 232.400 22.930 232.600 ;
        RECT 18.980 231.800 19.330 232.400 ;
        RECT 18.980 231.600 22.930 231.800 ;
        RECT 18.980 231.000 19.330 231.600 ;
        RECT 18.980 230.800 22.930 231.000 ;
        RECT 18.980 230.400 19.330 230.800 ;
        RECT 15.780 222.000 15.980 229.600 ;
        RECT 16.580 222.000 16.780 229.600 ;
        RECT 17.380 222.000 17.580 229.600 ;
        RECT 18.180 222.000 18.380 229.600 ;
        RECT 18.980 229.200 19.330 229.600 ;
        RECT 18.980 229.000 22.930 229.200 ;
        RECT 18.980 228.400 19.330 229.000 ;
        RECT 18.980 228.200 22.930 228.400 ;
        RECT 18.980 227.600 19.330 228.200 ;
        RECT 18.980 227.400 22.930 227.600 ;
        RECT 18.980 226.800 19.330 227.400 ;
        RECT 18.980 226.600 22.930 226.800 ;
        RECT 23.930 226.750 24.330 233.250 ;
        RECT 25.130 226.750 25.530 233.250 ;
        RECT 26.530 233.200 30.480 233.400 ;
        RECT 30.130 232.600 30.480 233.200 ;
        RECT 26.530 232.400 30.480 232.600 ;
        RECT 30.130 231.800 30.480 232.400 ;
        RECT 26.530 231.600 30.480 231.800 ;
        RECT 30.130 231.000 30.480 231.600 ;
        RECT 26.530 230.800 30.480 231.000 ;
        RECT 30.130 230.400 30.480 230.800 ;
        RECT 31.080 230.400 31.280 238.000 ;
        RECT 31.880 230.400 32.080 238.000 ;
        RECT 32.680 230.400 32.880 238.000 ;
        RECT 33.480 230.400 33.680 238.000 ;
        RECT 30.130 229.200 30.480 229.600 ;
        RECT 26.530 229.000 30.480 229.200 ;
        RECT 30.130 228.400 30.480 229.000 ;
        RECT 26.530 228.200 30.480 228.400 ;
        RECT 30.130 227.600 30.480 228.200 ;
        RECT 26.530 227.400 30.480 227.600 ;
        RECT 30.130 226.800 30.480 227.400 ;
        RECT 18.980 226.000 19.330 226.600 ;
        RECT 18.980 225.800 22.930 226.000 ;
        RECT 18.980 225.200 19.330 225.800 ;
        RECT 18.980 225.000 22.930 225.200 ;
        RECT 18.980 224.400 19.330 225.000 ;
        RECT 23.880 224.450 25.580 226.750 ;
        RECT 26.530 226.600 30.480 226.800 ;
        RECT 30.130 226.000 30.480 226.600 ;
        RECT 26.530 225.800 30.480 226.000 ;
        RECT 30.130 225.200 30.480 225.800 ;
        RECT 26.530 225.000 30.480 225.200 ;
        RECT 18.980 224.200 22.930 224.400 ;
        RECT 18.980 223.600 19.330 224.200 ;
        RECT 18.980 223.400 22.930 223.600 ;
        RECT 18.980 222.800 19.330 223.400 ;
        RECT 18.980 222.600 22.930 222.800 ;
        RECT 18.980 222.000 19.330 222.600 ;
        RECT 6.530 221.400 22.930 222.000 ;
        RECT 9.180 220.800 11.480 220.850 ;
        RECT 17.980 220.800 20.280 220.850 ;
        RECT 23.930 220.800 24.330 224.450 ;
        RECT 5.130 220.400 24.330 220.800 ;
        RECT 25.130 220.800 25.530 224.450 ;
        RECT 30.130 224.400 30.480 225.000 ;
        RECT 26.530 224.200 30.480 224.400 ;
        RECT 30.130 223.600 30.480 224.200 ;
        RECT 26.530 223.400 30.480 223.600 ;
        RECT 30.130 222.800 30.480 223.400 ;
        RECT 26.530 222.600 30.480 222.800 ;
        RECT 30.130 222.000 30.480 222.600 ;
        RECT 31.080 222.000 31.280 229.600 ;
        RECT 31.880 222.000 32.080 229.600 ;
        RECT 32.680 222.000 32.880 229.600 ;
        RECT 33.480 222.000 33.680 229.600 ;
        RECT 34.280 222.000 35.180 238.000 ;
        RECT 35.780 230.400 35.980 238.000 ;
        RECT 36.580 230.400 36.780 238.000 ;
        RECT 37.380 230.400 37.580 238.000 ;
        RECT 38.180 230.400 38.380 238.000 ;
        RECT 38.980 237.400 39.330 238.000 ;
        RECT 38.980 237.200 42.930 237.400 ;
        RECT 38.980 236.600 39.330 237.200 ;
        RECT 38.980 236.400 42.930 236.600 ;
        RECT 38.980 235.800 39.330 236.400 ;
        RECT 38.980 235.600 42.930 235.800 ;
        RECT 38.980 235.000 39.330 235.600 ;
        RECT 43.930 235.550 44.330 239.200 ;
        RECT 45.130 239.200 64.330 239.600 ;
        RECT 45.130 235.550 45.530 239.200 ;
        RECT 49.180 239.150 51.480 239.200 ;
        RECT 57.980 239.150 60.280 239.200 ;
        RECT 46.530 238.000 62.930 238.600 ;
        RECT 50.130 237.400 50.480 238.000 ;
        RECT 46.530 237.200 50.480 237.400 ;
        RECT 50.130 236.600 50.480 237.200 ;
        RECT 46.530 236.400 50.480 236.600 ;
        RECT 50.130 235.800 50.480 236.400 ;
        RECT 46.530 235.600 50.480 235.800 ;
        RECT 38.980 234.800 42.930 235.000 ;
        RECT 38.980 234.200 39.330 234.800 ;
        RECT 38.980 234.000 42.930 234.200 ;
        RECT 38.980 233.400 39.330 234.000 ;
        RECT 38.980 233.200 42.930 233.400 ;
        RECT 43.880 233.250 45.580 235.550 ;
        RECT 50.130 235.000 50.480 235.600 ;
        RECT 46.530 234.800 50.480 235.000 ;
        RECT 50.130 234.200 50.480 234.800 ;
        RECT 46.530 234.000 50.480 234.200 ;
        RECT 50.130 233.400 50.480 234.000 ;
        RECT 38.980 232.600 39.330 233.200 ;
        RECT 38.980 232.400 42.930 232.600 ;
        RECT 38.980 231.800 39.330 232.400 ;
        RECT 38.980 231.600 42.930 231.800 ;
        RECT 38.980 231.000 39.330 231.600 ;
        RECT 38.980 230.800 42.930 231.000 ;
        RECT 38.980 230.400 39.330 230.800 ;
        RECT 35.780 222.000 35.980 229.600 ;
        RECT 36.580 222.000 36.780 229.600 ;
        RECT 37.380 222.000 37.580 229.600 ;
        RECT 38.180 222.000 38.380 229.600 ;
        RECT 38.980 229.200 39.330 229.600 ;
        RECT 38.980 229.000 42.930 229.200 ;
        RECT 38.980 228.400 39.330 229.000 ;
        RECT 38.980 228.200 42.930 228.400 ;
        RECT 38.980 227.600 39.330 228.200 ;
        RECT 38.980 227.400 42.930 227.600 ;
        RECT 38.980 226.800 39.330 227.400 ;
        RECT 38.980 226.600 42.930 226.800 ;
        RECT 43.930 226.750 44.330 233.250 ;
        RECT 45.130 226.750 45.530 233.250 ;
        RECT 46.530 233.200 50.480 233.400 ;
        RECT 50.130 232.600 50.480 233.200 ;
        RECT 46.530 232.400 50.480 232.600 ;
        RECT 50.130 231.800 50.480 232.400 ;
        RECT 46.530 231.600 50.480 231.800 ;
        RECT 50.130 231.000 50.480 231.600 ;
        RECT 46.530 230.800 50.480 231.000 ;
        RECT 50.130 230.400 50.480 230.800 ;
        RECT 51.080 230.400 51.280 238.000 ;
        RECT 51.880 230.400 52.080 238.000 ;
        RECT 52.680 230.400 52.880 238.000 ;
        RECT 53.480 230.400 53.680 238.000 ;
        RECT 50.130 229.200 50.480 229.600 ;
        RECT 46.530 229.000 50.480 229.200 ;
        RECT 50.130 228.400 50.480 229.000 ;
        RECT 46.530 228.200 50.480 228.400 ;
        RECT 50.130 227.600 50.480 228.200 ;
        RECT 46.530 227.400 50.480 227.600 ;
        RECT 50.130 226.800 50.480 227.400 ;
        RECT 38.980 226.000 39.330 226.600 ;
        RECT 38.980 225.800 42.930 226.000 ;
        RECT 38.980 225.200 39.330 225.800 ;
        RECT 38.980 225.000 42.930 225.200 ;
        RECT 38.980 224.400 39.330 225.000 ;
        RECT 43.880 224.450 45.580 226.750 ;
        RECT 46.530 226.600 50.480 226.800 ;
        RECT 50.130 226.000 50.480 226.600 ;
        RECT 46.530 225.800 50.480 226.000 ;
        RECT 50.130 225.200 50.480 225.800 ;
        RECT 46.530 225.000 50.480 225.200 ;
        RECT 38.980 224.200 42.930 224.400 ;
        RECT 38.980 223.600 39.330 224.200 ;
        RECT 38.980 223.400 42.930 223.600 ;
        RECT 38.980 222.800 39.330 223.400 ;
        RECT 38.980 222.600 42.930 222.800 ;
        RECT 38.980 222.000 39.330 222.600 ;
        RECT 26.530 221.400 42.930 222.000 ;
        RECT 29.180 220.800 31.480 220.850 ;
        RECT 37.980 220.800 40.280 220.850 ;
        RECT 43.930 220.800 44.330 224.450 ;
        RECT 25.130 220.400 44.330 220.800 ;
        RECT 45.130 220.800 45.530 224.450 ;
        RECT 50.130 224.400 50.480 225.000 ;
        RECT 46.530 224.200 50.480 224.400 ;
        RECT 50.130 223.600 50.480 224.200 ;
        RECT 46.530 223.400 50.480 223.600 ;
        RECT 50.130 222.800 50.480 223.400 ;
        RECT 46.530 222.600 50.480 222.800 ;
        RECT 50.130 222.000 50.480 222.600 ;
        RECT 51.080 222.000 51.280 229.600 ;
        RECT 51.880 222.000 52.080 229.600 ;
        RECT 52.680 222.000 52.880 229.600 ;
        RECT 53.480 222.000 53.680 229.600 ;
        RECT 54.280 222.000 55.180 238.000 ;
        RECT 55.780 230.400 55.980 238.000 ;
        RECT 56.580 230.400 56.780 238.000 ;
        RECT 57.380 230.400 57.580 238.000 ;
        RECT 58.180 230.400 58.380 238.000 ;
        RECT 58.980 237.400 59.330 238.000 ;
        RECT 58.980 237.200 62.930 237.400 ;
        RECT 58.980 236.600 59.330 237.200 ;
        RECT 58.980 236.400 62.930 236.600 ;
        RECT 58.980 235.800 59.330 236.400 ;
        RECT 58.980 235.600 62.930 235.800 ;
        RECT 58.980 235.000 59.330 235.600 ;
        RECT 63.930 235.550 64.330 239.200 ;
        RECT 65.130 239.200 84.330 239.600 ;
        RECT 65.130 235.550 65.530 239.200 ;
        RECT 69.180 239.150 71.480 239.200 ;
        RECT 77.980 239.150 80.280 239.200 ;
        RECT 66.530 238.000 82.930 238.600 ;
        RECT 70.130 237.400 70.480 238.000 ;
        RECT 66.530 237.200 70.480 237.400 ;
        RECT 70.130 236.600 70.480 237.200 ;
        RECT 66.530 236.400 70.480 236.600 ;
        RECT 70.130 235.800 70.480 236.400 ;
        RECT 66.530 235.600 70.480 235.800 ;
        RECT 58.980 234.800 62.930 235.000 ;
        RECT 58.980 234.200 59.330 234.800 ;
        RECT 58.980 234.000 62.930 234.200 ;
        RECT 58.980 233.400 59.330 234.000 ;
        RECT 58.980 233.200 62.930 233.400 ;
        RECT 63.880 233.250 65.580 235.550 ;
        RECT 70.130 235.000 70.480 235.600 ;
        RECT 66.530 234.800 70.480 235.000 ;
        RECT 70.130 234.200 70.480 234.800 ;
        RECT 66.530 234.000 70.480 234.200 ;
        RECT 70.130 233.400 70.480 234.000 ;
        RECT 58.980 232.600 59.330 233.200 ;
        RECT 58.980 232.400 62.930 232.600 ;
        RECT 58.980 231.800 59.330 232.400 ;
        RECT 58.980 231.600 62.930 231.800 ;
        RECT 58.980 231.000 59.330 231.600 ;
        RECT 58.980 230.800 62.930 231.000 ;
        RECT 58.980 230.400 59.330 230.800 ;
        RECT 55.780 222.000 55.980 229.600 ;
        RECT 56.580 222.000 56.780 229.600 ;
        RECT 57.380 222.000 57.580 229.600 ;
        RECT 58.180 222.000 58.380 229.600 ;
        RECT 58.980 229.200 59.330 229.600 ;
        RECT 58.980 229.000 62.930 229.200 ;
        RECT 58.980 228.400 59.330 229.000 ;
        RECT 58.980 228.200 62.930 228.400 ;
        RECT 58.980 227.600 59.330 228.200 ;
        RECT 58.980 227.400 62.930 227.600 ;
        RECT 58.980 226.800 59.330 227.400 ;
        RECT 58.980 226.600 62.930 226.800 ;
        RECT 63.930 226.750 64.330 233.250 ;
        RECT 65.130 226.750 65.530 233.250 ;
        RECT 66.530 233.200 70.480 233.400 ;
        RECT 70.130 232.600 70.480 233.200 ;
        RECT 66.530 232.400 70.480 232.600 ;
        RECT 70.130 231.800 70.480 232.400 ;
        RECT 66.530 231.600 70.480 231.800 ;
        RECT 70.130 231.000 70.480 231.600 ;
        RECT 66.530 230.800 70.480 231.000 ;
        RECT 70.130 230.400 70.480 230.800 ;
        RECT 71.080 230.400 71.280 238.000 ;
        RECT 71.880 230.400 72.080 238.000 ;
        RECT 72.680 230.400 72.880 238.000 ;
        RECT 73.480 230.400 73.680 238.000 ;
        RECT 70.130 229.200 70.480 229.600 ;
        RECT 66.530 229.000 70.480 229.200 ;
        RECT 70.130 228.400 70.480 229.000 ;
        RECT 66.530 228.200 70.480 228.400 ;
        RECT 70.130 227.600 70.480 228.200 ;
        RECT 66.530 227.400 70.480 227.600 ;
        RECT 70.130 226.800 70.480 227.400 ;
        RECT 58.980 226.000 59.330 226.600 ;
        RECT 58.980 225.800 62.930 226.000 ;
        RECT 58.980 225.200 59.330 225.800 ;
        RECT 58.980 225.000 62.930 225.200 ;
        RECT 58.980 224.400 59.330 225.000 ;
        RECT 63.880 224.450 65.580 226.750 ;
        RECT 66.530 226.600 70.480 226.800 ;
        RECT 70.130 226.000 70.480 226.600 ;
        RECT 66.530 225.800 70.480 226.000 ;
        RECT 70.130 225.200 70.480 225.800 ;
        RECT 66.530 225.000 70.480 225.200 ;
        RECT 58.980 224.200 62.930 224.400 ;
        RECT 58.980 223.600 59.330 224.200 ;
        RECT 58.980 223.400 62.930 223.600 ;
        RECT 58.980 222.800 59.330 223.400 ;
        RECT 58.980 222.600 62.930 222.800 ;
        RECT 58.980 222.000 59.330 222.600 ;
        RECT 46.530 221.400 62.930 222.000 ;
        RECT 49.180 220.800 51.480 220.850 ;
        RECT 57.980 220.800 60.280 220.850 ;
        RECT 63.930 220.800 64.330 224.450 ;
        RECT 45.130 220.400 64.330 220.800 ;
        RECT 65.130 220.800 65.530 224.450 ;
        RECT 70.130 224.400 70.480 225.000 ;
        RECT 66.530 224.200 70.480 224.400 ;
        RECT 70.130 223.600 70.480 224.200 ;
        RECT 66.530 223.400 70.480 223.600 ;
        RECT 70.130 222.800 70.480 223.400 ;
        RECT 66.530 222.600 70.480 222.800 ;
        RECT 70.130 222.000 70.480 222.600 ;
        RECT 71.080 222.000 71.280 229.600 ;
        RECT 71.880 222.000 72.080 229.600 ;
        RECT 72.680 222.000 72.880 229.600 ;
        RECT 73.480 222.000 73.680 229.600 ;
        RECT 74.280 222.000 75.180 238.000 ;
        RECT 75.780 230.400 75.980 238.000 ;
        RECT 76.580 230.400 76.780 238.000 ;
        RECT 77.380 230.400 77.580 238.000 ;
        RECT 78.180 230.400 78.380 238.000 ;
        RECT 78.980 237.400 79.330 238.000 ;
        RECT 78.980 237.200 82.930 237.400 ;
        RECT 78.980 236.600 79.330 237.200 ;
        RECT 78.980 236.400 82.930 236.600 ;
        RECT 78.980 235.800 79.330 236.400 ;
        RECT 78.980 235.600 82.930 235.800 ;
        RECT 78.980 235.000 79.330 235.600 ;
        RECT 83.930 235.550 84.330 239.200 ;
        RECT 85.130 239.200 104.330 239.600 ;
        RECT 85.130 235.550 85.530 239.200 ;
        RECT 89.180 239.150 91.480 239.200 ;
        RECT 97.980 239.150 100.280 239.200 ;
        RECT 86.530 238.000 102.930 238.600 ;
        RECT 90.130 237.400 90.480 238.000 ;
        RECT 86.530 237.200 90.480 237.400 ;
        RECT 90.130 236.600 90.480 237.200 ;
        RECT 86.530 236.400 90.480 236.600 ;
        RECT 90.130 235.800 90.480 236.400 ;
        RECT 86.530 235.600 90.480 235.800 ;
        RECT 78.980 234.800 82.930 235.000 ;
        RECT 78.980 234.200 79.330 234.800 ;
        RECT 78.980 234.000 82.930 234.200 ;
        RECT 78.980 233.400 79.330 234.000 ;
        RECT 78.980 233.200 82.930 233.400 ;
        RECT 83.880 233.250 85.580 235.550 ;
        RECT 90.130 235.000 90.480 235.600 ;
        RECT 86.530 234.800 90.480 235.000 ;
        RECT 90.130 234.200 90.480 234.800 ;
        RECT 86.530 234.000 90.480 234.200 ;
        RECT 90.130 233.400 90.480 234.000 ;
        RECT 78.980 232.600 79.330 233.200 ;
        RECT 78.980 232.400 82.930 232.600 ;
        RECT 78.980 231.800 79.330 232.400 ;
        RECT 78.980 231.600 82.930 231.800 ;
        RECT 78.980 231.000 79.330 231.600 ;
        RECT 78.980 230.800 82.930 231.000 ;
        RECT 78.980 230.400 79.330 230.800 ;
        RECT 75.780 222.000 75.980 229.600 ;
        RECT 76.580 222.000 76.780 229.600 ;
        RECT 77.380 222.000 77.580 229.600 ;
        RECT 78.180 222.000 78.380 229.600 ;
        RECT 78.980 229.200 79.330 229.600 ;
        RECT 78.980 229.000 82.930 229.200 ;
        RECT 78.980 228.400 79.330 229.000 ;
        RECT 78.980 228.200 82.930 228.400 ;
        RECT 78.980 227.600 79.330 228.200 ;
        RECT 78.980 227.400 82.930 227.600 ;
        RECT 78.980 226.800 79.330 227.400 ;
        RECT 78.980 226.600 82.930 226.800 ;
        RECT 83.930 226.750 84.330 233.250 ;
        RECT 85.130 226.750 85.530 233.250 ;
        RECT 86.530 233.200 90.480 233.400 ;
        RECT 90.130 232.600 90.480 233.200 ;
        RECT 86.530 232.400 90.480 232.600 ;
        RECT 90.130 231.800 90.480 232.400 ;
        RECT 86.530 231.600 90.480 231.800 ;
        RECT 90.130 231.000 90.480 231.600 ;
        RECT 86.530 230.800 90.480 231.000 ;
        RECT 90.130 230.400 90.480 230.800 ;
        RECT 91.080 230.400 91.280 238.000 ;
        RECT 91.880 230.400 92.080 238.000 ;
        RECT 92.680 230.400 92.880 238.000 ;
        RECT 93.480 230.400 93.680 238.000 ;
        RECT 90.130 229.200 90.480 229.600 ;
        RECT 86.530 229.000 90.480 229.200 ;
        RECT 90.130 228.400 90.480 229.000 ;
        RECT 86.530 228.200 90.480 228.400 ;
        RECT 90.130 227.600 90.480 228.200 ;
        RECT 86.530 227.400 90.480 227.600 ;
        RECT 90.130 226.800 90.480 227.400 ;
        RECT 78.980 226.000 79.330 226.600 ;
        RECT 78.980 225.800 82.930 226.000 ;
        RECT 78.980 225.200 79.330 225.800 ;
        RECT 78.980 225.000 82.930 225.200 ;
        RECT 78.980 224.400 79.330 225.000 ;
        RECT 83.880 224.450 85.580 226.750 ;
        RECT 86.530 226.600 90.480 226.800 ;
        RECT 90.130 226.000 90.480 226.600 ;
        RECT 86.530 225.800 90.480 226.000 ;
        RECT 90.130 225.200 90.480 225.800 ;
        RECT 86.530 225.000 90.480 225.200 ;
        RECT 78.980 224.200 82.930 224.400 ;
        RECT 78.980 223.600 79.330 224.200 ;
        RECT 78.980 223.400 82.930 223.600 ;
        RECT 78.980 222.800 79.330 223.400 ;
        RECT 78.980 222.600 82.930 222.800 ;
        RECT 78.980 222.000 79.330 222.600 ;
        RECT 66.530 221.400 82.930 222.000 ;
        RECT 69.180 220.800 71.480 220.850 ;
        RECT 77.980 220.800 80.280 220.850 ;
        RECT 83.930 220.800 84.330 224.450 ;
        RECT 65.130 220.400 84.330 220.800 ;
        RECT 85.130 220.800 85.530 224.450 ;
        RECT 90.130 224.400 90.480 225.000 ;
        RECT 86.530 224.200 90.480 224.400 ;
        RECT 90.130 223.600 90.480 224.200 ;
        RECT 86.530 223.400 90.480 223.600 ;
        RECT 90.130 222.800 90.480 223.400 ;
        RECT 86.530 222.600 90.480 222.800 ;
        RECT 90.130 222.000 90.480 222.600 ;
        RECT 91.080 222.000 91.280 229.600 ;
        RECT 91.880 222.000 92.080 229.600 ;
        RECT 92.680 222.000 92.880 229.600 ;
        RECT 93.480 222.000 93.680 229.600 ;
        RECT 94.280 222.000 95.180 238.000 ;
        RECT 95.780 230.400 95.980 238.000 ;
        RECT 96.580 230.400 96.780 238.000 ;
        RECT 97.380 230.400 97.580 238.000 ;
        RECT 98.180 230.400 98.380 238.000 ;
        RECT 98.980 237.400 99.330 238.000 ;
        RECT 98.980 237.200 102.930 237.400 ;
        RECT 98.980 236.600 99.330 237.200 ;
        RECT 98.980 236.400 102.930 236.600 ;
        RECT 98.980 235.800 99.330 236.400 ;
        RECT 98.980 235.600 102.930 235.800 ;
        RECT 98.980 235.000 99.330 235.600 ;
        RECT 103.930 235.550 104.330 239.200 ;
        RECT 105.340 237.260 105.700 237.640 ;
        RECT 105.970 237.260 106.330 237.640 ;
        RECT 106.570 237.260 106.930 237.640 ;
        RECT 105.340 236.670 105.700 237.050 ;
        RECT 105.970 236.670 106.330 237.050 ;
        RECT 106.570 236.670 106.930 237.050 ;
        RECT 98.980 234.800 102.930 235.000 ;
        RECT 98.980 234.200 99.330 234.800 ;
        RECT 98.980 234.000 102.930 234.200 ;
        RECT 98.980 233.400 99.330 234.000 ;
        RECT 98.980 233.200 102.930 233.400 ;
        RECT 103.880 233.250 104.730 235.550 ;
        RECT 98.980 232.600 99.330 233.200 ;
        RECT 98.980 232.400 102.930 232.600 ;
        RECT 98.980 231.800 99.330 232.400 ;
        RECT 98.980 231.600 102.930 231.800 ;
        RECT 98.980 231.000 99.330 231.600 ;
        RECT 98.980 230.800 102.930 231.000 ;
        RECT 98.980 230.400 99.330 230.800 ;
        RECT 95.780 222.000 95.980 229.600 ;
        RECT 96.580 222.000 96.780 229.600 ;
        RECT 97.380 222.000 97.580 229.600 ;
        RECT 98.180 222.000 98.380 229.600 ;
        RECT 98.980 229.200 99.330 229.600 ;
        RECT 98.980 229.000 102.930 229.200 ;
        RECT 98.980 228.400 99.330 229.000 ;
        RECT 98.980 228.200 102.930 228.400 ;
        RECT 98.980 227.600 99.330 228.200 ;
        RECT 98.980 227.400 102.930 227.600 ;
        RECT 98.980 226.800 99.330 227.400 ;
        RECT 98.980 226.600 102.930 226.800 ;
        RECT 103.930 226.750 104.330 233.250 ;
        RECT 98.980 226.000 99.330 226.600 ;
        RECT 98.980 225.800 102.930 226.000 ;
        RECT 98.980 225.200 99.330 225.800 ;
        RECT 98.980 225.000 102.930 225.200 ;
        RECT 98.980 224.400 99.330 225.000 ;
        RECT 103.880 224.450 104.730 226.750 ;
        RECT 98.980 224.200 102.930 224.400 ;
        RECT 98.980 223.600 99.330 224.200 ;
        RECT 98.980 223.400 102.930 223.600 ;
        RECT 98.980 222.800 99.330 223.400 ;
        RECT 98.980 222.600 102.930 222.800 ;
        RECT 98.980 222.000 99.330 222.600 ;
        RECT 86.530 221.400 102.930 222.000 ;
        RECT 89.180 220.800 91.480 220.850 ;
        RECT 97.980 220.800 100.280 220.850 ;
        RECT 103.930 220.800 104.330 224.450 ;
        RECT 105.340 221.680 105.700 222.060 ;
        RECT 105.970 221.680 106.330 222.060 ;
        RECT 106.570 221.680 106.930 222.060 ;
        RECT 105.340 221.090 105.700 221.470 ;
        RECT 105.970 221.090 106.330 221.470 ;
        RECT 106.570 221.090 106.930 221.470 ;
        RECT 85.130 220.400 104.330 220.800 ;
        RECT 9.180 220.000 11.480 220.400 ;
        RECT 17.980 220.000 20.280 220.400 ;
        RECT 29.180 220.000 31.480 220.400 ;
        RECT 37.980 220.000 40.280 220.400 ;
        RECT 49.180 220.000 51.480 220.400 ;
        RECT 57.980 220.000 60.280 220.400 ;
        RECT 69.180 220.000 71.480 220.400 ;
        RECT 77.980 220.000 80.280 220.400 ;
        RECT 89.180 220.000 91.480 220.400 ;
        RECT 97.980 220.000 100.280 220.400 ;
        RECT 4.620 197.380 26.020 198.635 ;
        RECT 4.620 183.250 5.940 197.380 ;
        RECT 6.940 195.375 7.400 195.545 ;
        RECT 7.025 194.650 7.315 195.375 ;
        RECT 8.020 193.450 8.190 195.695 ;
        RECT 9.595 195.290 9.770 195.695 ;
        RECT 24.570 195.540 26.020 197.380 ;
        RECT 14.865 195.370 26.020 195.540 ;
        RECT 9.600 193.450 9.770 195.290 ;
        RECT 14.950 194.645 15.240 195.370 ;
        RECT 15.560 194.570 15.890 195.370 ;
        RECT 16.400 194.890 16.730 195.370 ;
        RECT 17.320 194.890 17.560 195.370 ;
        RECT 18.320 194.570 18.650 195.370 ;
        RECT 19.160 194.890 19.490 195.370 ;
        RECT 20.080 194.890 20.320 195.370 ;
        RECT 21.675 194.550 21.905 195.370 ;
        RECT 23.055 194.550 23.285 195.370 ;
        RECT 8.050 190.100 8.340 190.825 ;
        RECT 9.410 190.100 9.720 190.900 ;
        RECT 10.500 190.100 10.885 190.500 ;
        RECT 11.915 190.100 12.300 190.500 ;
        RECT 13.330 190.100 13.715 190.500 ;
        RECT 15.100 190.100 15.485 190.500 ;
        RECT 16.515 190.100 16.900 190.500 ;
        RECT 17.930 190.100 18.315 190.500 ;
        RECT 19.700 190.100 20.085 190.500 ;
        RECT 21.115 190.100 21.500 190.500 ;
        RECT 22.530 190.100 22.915 190.500 ;
        RECT 23.690 190.100 23.980 190.825 ;
        RECT 24.570 190.100 26.020 195.370 ;
        RECT 6.585 189.930 26.020 190.100 ;
        RECT 6.670 189.205 6.960 189.930 ;
        RECT 7.365 189.110 7.595 189.930 ;
        RECT 8.510 189.130 8.820 189.930 ;
        RECT 10.500 189.530 10.885 189.930 ;
        RECT 11.915 189.530 12.300 189.930 ;
        RECT 13.330 189.530 13.715 189.930 ;
        RECT 15.100 189.530 15.485 189.930 ;
        RECT 16.515 189.530 16.900 189.930 ;
        RECT 17.930 189.530 18.315 189.930 ;
        RECT 19.700 189.530 20.085 189.930 ;
        RECT 21.115 189.530 21.500 189.930 ;
        RECT 22.530 189.530 22.915 189.930 ;
        RECT 23.690 189.205 23.980 189.930 ;
        RECT 7.590 184.660 7.880 185.385 ;
        RECT 14.950 184.660 15.240 185.385 ;
        RECT 15.560 184.660 15.890 185.460 ;
        RECT 16.400 184.660 16.730 185.140 ;
        RECT 17.320 184.660 17.560 185.140 ;
        RECT 18.320 184.660 18.650 185.460 ;
        RECT 19.160 184.660 19.490 185.140 ;
        RECT 20.080 184.660 20.320 185.140 ;
        RECT 21.675 184.660 21.905 185.480 ;
        RECT 23.055 184.660 23.285 185.480 ;
        RECT 24.570 184.660 26.020 189.930 ;
        RECT 7.505 184.490 7.965 184.660 ;
        RECT 14.865 184.490 26.020 184.660 ;
        RECT 24.570 183.250 26.020 184.490 ;
        RECT 4.620 182.245 26.020 183.250 ;
        RECT 47.085 182.260 49.385 182.660 ;
        RECT 55.885 182.260 58.185 182.660 ;
        RECT 67.085 182.260 69.385 182.660 ;
        RECT 75.885 182.260 78.185 182.660 ;
        RECT 87.085 182.260 89.385 182.660 ;
        RECT 95.885 182.260 98.185 182.660 ;
        RECT 4.620 182.055 26.015 182.245 ;
        RECT 43.035 181.860 62.235 182.260 ;
        RECT 43.035 178.210 43.435 181.860 ;
        RECT 47.085 181.810 49.385 181.860 ;
        RECT 55.885 181.810 58.185 181.860 ;
        RECT 44.435 180.660 60.835 181.260 ;
        RECT 48.035 180.060 48.385 180.660 ;
        RECT 44.435 179.860 48.385 180.060 ;
        RECT 48.035 179.260 48.385 179.860 ;
        RECT 44.435 179.060 48.385 179.260 ;
        RECT 48.035 178.460 48.385 179.060 ;
        RECT 44.435 178.260 48.385 178.460 ;
        RECT 42.635 175.910 43.485 178.210 ;
        RECT 48.035 177.660 48.385 178.260 ;
        RECT 44.435 177.460 48.385 177.660 ;
        RECT 48.035 176.860 48.385 177.460 ;
        RECT 44.435 176.660 48.385 176.860 ;
        RECT 48.035 176.060 48.385 176.660 ;
        RECT 43.035 169.410 43.435 175.910 ;
        RECT 44.435 175.860 48.385 176.060 ;
        RECT 48.035 175.260 48.385 175.860 ;
        RECT 44.435 175.060 48.385 175.260 ;
        RECT 48.035 174.460 48.385 175.060 ;
        RECT 44.435 174.260 48.385 174.460 ;
        RECT 48.035 173.660 48.385 174.260 ;
        RECT 44.435 173.460 48.385 173.660 ;
        RECT 48.035 173.060 48.385 173.460 ;
        RECT 48.985 173.060 49.185 180.660 ;
        RECT 49.785 173.060 49.985 180.660 ;
        RECT 50.585 173.060 50.785 180.660 ;
        RECT 51.385 173.060 51.585 180.660 ;
        RECT 48.035 171.860 48.385 172.260 ;
        RECT 44.435 171.660 48.385 171.860 ;
        RECT 48.035 171.060 48.385 171.660 ;
        RECT 44.435 170.860 48.385 171.060 ;
        RECT 48.035 170.260 48.385 170.860 ;
        RECT 44.435 170.060 48.385 170.260 ;
        RECT 48.035 169.460 48.385 170.060 ;
        RECT 42.635 167.110 43.485 169.410 ;
        RECT 44.435 169.260 48.385 169.460 ;
        RECT 48.035 168.660 48.385 169.260 ;
        RECT 44.435 168.460 48.385 168.660 ;
        RECT 48.035 167.860 48.385 168.460 ;
        RECT 44.435 167.660 48.385 167.860 ;
        RECT 43.035 163.460 43.435 167.110 ;
        RECT 48.035 167.060 48.385 167.660 ;
        RECT 44.435 166.860 48.385 167.060 ;
        RECT 48.035 166.260 48.385 166.860 ;
        RECT 44.435 166.060 48.385 166.260 ;
        RECT 48.035 165.460 48.385 166.060 ;
        RECT 44.435 165.260 48.385 165.460 ;
        RECT 48.035 164.660 48.385 165.260 ;
        RECT 48.985 164.660 49.185 172.260 ;
        RECT 49.785 164.660 49.985 172.260 ;
        RECT 50.585 164.660 50.785 172.260 ;
        RECT 51.385 164.660 51.585 172.260 ;
        RECT 52.185 164.660 53.085 180.660 ;
        RECT 53.685 173.060 53.885 180.660 ;
        RECT 54.485 173.060 54.685 180.660 ;
        RECT 55.285 173.060 55.485 180.660 ;
        RECT 56.085 173.060 56.285 180.660 ;
        RECT 56.885 180.060 57.235 180.660 ;
        RECT 56.885 179.860 60.835 180.060 ;
        RECT 56.885 179.260 57.235 179.860 ;
        RECT 56.885 179.060 60.835 179.260 ;
        RECT 56.885 178.460 57.235 179.060 ;
        RECT 56.885 178.260 60.835 178.460 ;
        RECT 56.885 177.660 57.235 178.260 ;
        RECT 61.835 178.210 62.235 181.860 ;
        RECT 63.035 181.860 82.235 182.260 ;
        RECT 63.035 178.210 63.435 181.860 ;
        RECT 67.085 181.810 69.385 181.860 ;
        RECT 75.885 181.810 78.185 181.860 ;
        RECT 64.435 180.660 80.835 181.260 ;
        RECT 68.035 180.060 68.385 180.660 ;
        RECT 64.435 179.860 68.385 180.060 ;
        RECT 68.035 179.260 68.385 179.860 ;
        RECT 64.435 179.060 68.385 179.260 ;
        RECT 68.035 178.460 68.385 179.060 ;
        RECT 64.435 178.260 68.385 178.460 ;
        RECT 56.885 177.460 60.835 177.660 ;
        RECT 56.885 176.860 57.235 177.460 ;
        RECT 56.885 176.660 60.835 176.860 ;
        RECT 56.885 176.060 57.235 176.660 ;
        RECT 56.885 175.860 60.835 176.060 ;
        RECT 61.785 175.910 63.485 178.210 ;
        RECT 68.035 177.660 68.385 178.260 ;
        RECT 64.435 177.460 68.385 177.660 ;
        RECT 68.035 176.860 68.385 177.460 ;
        RECT 64.435 176.660 68.385 176.860 ;
        RECT 68.035 176.060 68.385 176.660 ;
        RECT 56.885 175.260 57.235 175.860 ;
        RECT 56.885 175.060 60.835 175.260 ;
        RECT 56.885 174.460 57.235 175.060 ;
        RECT 56.885 174.260 60.835 174.460 ;
        RECT 56.885 173.660 57.235 174.260 ;
        RECT 56.885 173.460 60.835 173.660 ;
        RECT 56.885 173.060 57.235 173.460 ;
        RECT 53.685 164.660 53.885 172.260 ;
        RECT 54.485 164.660 54.685 172.260 ;
        RECT 55.285 164.660 55.485 172.260 ;
        RECT 56.085 164.660 56.285 172.260 ;
        RECT 56.885 171.860 57.235 172.260 ;
        RECT 56.885 171.660 60.835 171.860 ;
        RECT 56.885 171.060 57.235 171.660 ;
        RECT 56.885 170.860 60.835 171.060 ;
        RECT 56.885 170.260 57.235 170.860 ;
        RECT 56.885 170.060 60.835 170.260 ;
        RECT 56.885 169.460 57.235 170.060 ;
        RECT 56.885 169.260 60.835 169.460 ;
        RECT 61.835 169.410 62.235 175.910 ;
        RECT 63.035 169.410 63.435 175.910 ;
        RECT 64.435 175.860 68.385 176.060 ;
        RECT 68.035 175.260 68.385 175.860 ;
        RECT 64.435 175.060 68.385 175.260 ;
        RECT 68.035 174.460 68.385 175.060 ;
        RECT 64.435 174.260 68.385 174.460 ;
        RECT 68.035 173.660 68.385 174.260 ;
        RECT 64.435 173.460 68.385 173.660 ;
        RECT 68.035 173.060 68.385 173.460 ;
        RECT 68.985 173.060 69.185 180.660 ;
        RECT 69.785 173.060 69.985 180.660 ;
        RECT 70.585 173.060 70.785 180.660 ;
        RECT 71.385 173.060 71.585 180.660 ;
        RECT 68.035 171.860 68.385 172.260 ;
        RECT 64.435 171.660 68.385 171.860 ;
        RECT 68.035 171.060 68.385 171.660 ;
        RECT 64.435 170.860 68.385 171.060 ;
        RECT 68.035 170.260 68.385 170.860 ;
        RECT 64.435 170.060 68.385 170.260 ;
        RECT 68.035 169.460 68.385 170.060 ;
        RECT 56.885 168.660 57.235 169.260 ;
        RECT 56.885 168.460 60.835 168.660 ;
        RECT 56.885 167.860 57.235 168.460 ;
        RECT 56.885 167.660 60.835 167.860 ;
        RECT 56.885 167.060 57.235 167.660 ;
        RECT 61.785 167.110 63.485 169.410 ;
        RECT 64.435 169.260 68.385 169.460 ;
        RECT 68.035 168.660 68.385 169.260 ;
        RECT 64.435 168.460 68.385 168.660 ;
        RECT 68.035 167.860 68.385 168.460 ;
        RECT 64.435 167.660 68.385 167.860 ;
        RECT 56.885 166.860 60.835 167.060 ;
        RECT 56.885 166.260 57.235 166.860 ;
        RECT 56.885 166.060 60.835 166.260 ;
        RECT 56.885 165.460 57.235 166.060 ;
        RECT 56.885 165.260 60.835 165.460 ;
        RECT 56.885 164.660 57.235 165.260 ;
        RECT 44.435 164.060 60.835 164.660 ;
        RECT 47.085 163.460 49.385 163.510 ;
        RECT 55.885 163.460 58.185 163.510 ;
        RECT 61.835 163.460 62.235 167.110 ;
        RECT 43.035 163.060 62.235 163.460 ;
        RECT 63.035 163.460 63.435 167.110 ;
        RECT 68.035 167.060 68.385 167.660 ;
        RECT 64.435 166.860 68.385 167.060 ;
        RECT 68.035 166.260 68.385 166.860 ;
        RECT 64.435 166.060 68.385 166.260 ;
        RECT 68.035 165.460 68.385 166.060 ;
        RECT 64.435 165.260 68.385 165.460 ;
        RECT 68.035 164.660 68.385 165.260 ;
        RECT 68.985 164.660 69.185 172.260 ;
        RECT 69.785 164.660 69.985 172.260 ;
        RECT 70.585 164.660 70.785 172.260 ;
        RECT 71.385 164.660 71.585 172.260 ;
        RECT 72.185 164.660 73.085 180.660 ;
        RECT 73.685 173.060 73.885 180.660 ;
        RECT 74.485 173.060 74.685 180.660 ;
        RECT 75.285 173.060 75.485 180.660 ;
        RECT 76.085 173.060 76.285 180.660 ;
        RECT 76.885 180.060 77.235 180.660 ;
        RECT 76.885 179.860 80.835 180.060 ;
        RECT 76.885 179.260 77.235 179.860 ;
        RECT 76.885 179.060 80.835 179.260 ;
        RECT 76.885 178.460 77.235 179.060 ;
        RECT 76.885 178.260 80.835 178.460 ;
        RECT 76.885 177.660 77.235 178.260 ;
        RECT 81.835 178.210 82.235 181.860 ;
        RECT 83.035 181.860 102.235 182.260 ;
        RECT 83.035 178.210 83.435 181.860 ;
        RECT 87.085 181.810 89.385 181.860 ;
        RECT 95.885 181.810 98.185 181.860 ;
        RECT 84.435 180.660 100.835 181.260 ;
        RECT 88.035 180.060 88.385 180.660 ;
        RECT 84.435 179.860 88.385 180.060 ;
        RECT 88.035 179.260 88.385 179.860 ;
        RECT 84.435 179.060 88.385 179.260 ;
        RECT 88.035 178.460 88.385 179.060 ;
        RECT 84.435 178.260 88.385 178.460 ;
        RECT 76.885 177.460 80.835 177.660 ;
        RECT 76.885 176.860 77.235 177.460 ;
        RECT 76.885 176.660 80.835 176.860 ;
        RECT 76.885 176.060 77.235 176.660 ;
        RECT 76.885 175.860 80.835 176.060 ;
        RECT 81.785 175.910 83.485 178.210 ;
        RECT 88.035 177.660 88.385 178.260 ;
        RECT 84.435 177.460 88.385 177.660 ;
        RECT 88.035 176.860 88.385 177.460 ;
        RECT 84.435 176.660 88.385 176.860 ;
        RECT 88.035 176.060 88.385 176.660 ;
        RECT 76.885 175.260 77.235 175.860 ;
        RECT 76.885 175.060 80.835 175.260 ;
        RECT 76.885 174.460 77.235 175.060 ;
        RECT 76.885 174.260 80.835 174.460 ;
        RECT 76.885 173.660 77.235 174.260 ;
        RECT 76.885 173.460 80.835 173.660 ;
        RECT 76.885 173.060 77.235 173.460 ;
        RECT 73.685 164.660 73.885 172.260 ;
        RECT 74.485 164.660 74.685 172.260 ;
        RECT 75.285 164.660 75.485 172.260 ;
        RECT 76.085 164.660 76.285 172.260 ;
        RECT 76.885 171.860 77.235 172.260 ;
        RECT 76.885 171.660 80.835 171.860 ;
        RECT 76.885 171.060 77.235 171.660 ;
        RECT 76.885 170.860 80.835 171.060 ;
        RECT 76.885 170.260 77.235 170.860 ;
        RECT 76.885 170.060 80.835 170.260 ;
        RECT 76.885 169.460 77.235 170.060 ;
        RECT 76.885 169.260 80.835 169.460 ;
        RECT 81.835 169.410 82.235 175.910 ;
        RECT 83.035 169.410 83.435 175.910 ;
        RECT 84.435 175.860 88.385 176.060 ;
        RECT 88.035 175.260 88.385 175.860 ;
        RECT 84.435 175.060 88.385 175.260 ;
        RECT 88.035 174.460 88.385 175.060 ;
        RECT 84.435 174.260 88.385 174.460 ;
        RECT 88.035 173.660 88.385 174.260 ;
        RECT 84.435 173.460 88.385 173.660 ;
        RECT 88.035 173.060 88.385 173.460 ;
        RECT 88.985 173.060 89.185 180.660 ;
        RECT 89.785 173.060 89.985 180.660 ;
        RECT 90.585 173.060 90.785 180.660 ;
        RECT 91.385 173.060 91.585 180.660 ;
        RECT 88.035 171.860 88.385 172.260 ;
        RECT 84.435 171.660 88.385 171.860 ;
        RECT 88.035 171.060 88.385 171.660 ;
        RECT 84.435 170.860 88.385 171.060 ;
        RECT 88.035 170.260 88.385 170.860 ;
        RECT 84.435 170.060 88.385 170.260 ;
        RECT 88.035 169.460 88.385 170.060 ;
        RECT 76.885 168.660 77.235 169.260 ;
        RECT 76.885 168.460 80.835 168.660 ;
        RECT 76.885 167.860 77.235 168.460 ;
        RECT 76.885 167.660 80.835 167.860 ;
        RECT 76.885 167.060 77.235 167.660 ;
        RECT 81.785 167.110 83.485 169.410 ;
        RECT 84.435 169.260 88.385 169.460 ;
        RECT 88.035 168.660 88.385 169.260 ;
        RECT 84.435 168.460 88.385 168.660 ;
        RECT 88.035 167.860 88.385 168.460 ;
        RECT 84.435 167.660 88.385 167.860 ;
        RECT 76.885 166.860 80.835 167.060 ;
        RECT 76.885 166.260 77.235 166.860 ;
        RECT 76.885 166.060 80.835 166.260 ;
        RECT 76.885 165.460 77.235 166.060 ;
        RECT 76.885 165.260 80.835 165.460 ;
        RECT 76.885 164.660 77.235 165.260 ;
        RECT 64.435 164.060 80.835 164.660 ;
        RECT 67.085 163.460 69.385 163.510 ;
        RECT 75.885 163.460 78.185 163.510 ;
        RECT 81.835 163.460 82.235 167.110 ;
        RECT 63.035 163.060 82.235 163.460 ;
        RECT 83.035 163.460 83.435 167.110 ;
        RECT 88.035 167.060 88.385 167.660 ;
        RECT 84.435 166.860 88.385 167.060 ;
        RECT 88.035 166.260 88.385 166.860 ;
        RECT 84.435 166.060 88.385 166.260 ;
        RECT 88.035 165.460 88.385 166.060 ;
        RECT 84.435 165.260 88.385 165.460 ;
        RECT 88.035 164.660 88.385 165.260 ;
        RECT 88.985 164.660 89.185 172.260 ;
        RECT 89.785 164.660 89.985 172.260 ;
        RECT 90.585 164.660 90.785 172.260 ;
        RECT 91.385 164.660 91.585 172.260 ;
        RECT 92.185 164.660 93.085 180.660 ;
        RECT 93.685 173.060 93.885 180.660 ;
        RECT 94.485 173.060 94.685 180.660 ;
        RECT 95.285 173.060 95.485 180.660 ;
        RECT 96.085 173.060 96.285 180.660 ;
        RECT 96.885 180.060 97.235 180.660 ;
        RECT 96.885 179.860 100.835 180.060 ;
        RECT 96.885 179.260 97.235 179.860 ;
        RECT 96.885 179.060 100.835 179.260 ;
        RECT 96.885 178.460 97.235 179.060 ;
        RECT 96.885 178.260 100.835 178.460 ;
        RECT 96.885 177.660 97.235 178.260 ;
        RECT 101.835 178.210 102.235 181.860 ;
        RECT 96.885 177.460 100.835 177.660 ;
        RECT 96.885 176.860 97.235 177.460 ;
        RECT 96.885 176.660 100.835 176.860 ;
        RECT 96.885 176.060 97.235 176.660 ;
        RECT 96.885 175.860 100.835 176.060 ;
        RECT 101.785 175.915 107.140 178.210 ;
        RECT 101.785 175.910 107.005 175.915 ;
        RECT 96.885 175.260 97.235 175.860 ;
        RECT 96.885 175.060 100.835 175.260 ;
        RECT 96.885 174.460 97.235 175.060 ;
        RECT 96.885 174.260 100.835 174.460 ;
        RECT 96.885 173.660 97.235 174.260 ;
        RECT 96.885 173.460 100.835 173.660 ;
        RECT 96.885 173.060 97.235 173.460 ;
        RECT 93.685 164.660 93.885 172.260 ;
        RECT 94.485 164.660 94.685 172.260 ;
        RECT 95.285 164.660 95.485 172.260 ;
        RECT 96.085 164.660 96.285 172.260 ;
        RECT 96.885 171.860 97.235 172.260 ;
        RECT 96.885 171.660 100.835 171.860 ;
        RECT 96.885 171.060 97.235 171.660 ;
        RECT 96.885 170.860 100.835 171.060 ;
        RECT 96.885 170.260 97.235 170.860 ;
        RECT 96.885 170.060 100.835 170.260 ;
        RECT 96.885 169.460 97.235 170.060 ;
        RECT 96.885 169.260 100.835 169.460 ;
        RECT 101.835 169.410 102.235 175.910 ;
        RECT 96.885 168.660 97.235 169.260 ;
        RECT 96.885 168.460 100.835 168.660 ;
        RECT 96.885 167.860 97.235 168.460 ;
        RECT 96.885 167.660 100.835 167.860 ;
        RECT 96.885 167.060 97.235 167.660 ;
        RECT 101.785 167.115 107.140 169.410 ;
        RECT 101.785 167.110 107.005 167.115 ;
        RECT 96.885 166.860 100.835 167.060 ;
        RECT 96.885 166.260 97.235 166.860 ;
        RECT 96.885 166.060 100.835 166.260 ;
        RECT 96.885 165.460 97.235 166.060 ;
        RECT 96.885 165.260 100.835 165.460 ;
        RECT 96.885 164.660 97.235 165.260 ;
        RECT 84.435 164.060 100.835 164.660 ;
        RECT 87.085 163.460 89.385 163.510 ;
        RECT 95.885 163.460 98.185 163.510 ;
        RECT 101.835 163.460 102.235 167.110 ;
        RECT 83.035 163.060 102.235 163.460 ;
        RECT 47.085 162.660 49.385 163.060 ;
        RECT 55.885 162.660 58.185 163.060 ;
        RECT 67.085 162.660 69.385 163.060 ;
        RECT 75.885 162.660 78.185 163.060 ;
        RECT 87.085 162.660 89.385 163.060 ;
        RECT 95.885 162.660 98.185 163.060 ;
        RECT 2.515 161.130 2.875 161.510 ;
        RECT 3.145 161.130 3.505 161.510 ;
        RECT 3.745 161.130 4.105 161.510 ;
        RECT 105.340 161.130 105.700 161.510 ;
        RECT 105.970 161.130 106.330 161.510 ;
        RECT 106.570 161.130 106.930 161.510 ;
        RECT 2.515 160.540 2.875 160.920 ;
        RECT 3.145 160.540 3.505 160.920 ;
        RECT 3.745 160.540 4.105 160.920 ;
        RECT 105.340 160.540 105.700 160.920 ;
        RECT 105.970 160.540 106.330 160.920 ;
        RECT 106.570 160.540 106.930 160.920 ;
        RECT 9.180 159.600 11.480 160.000 ;
        RECT 17.980 159.600 20.280 160.000 ;
        RECT 29.180 159.600 31.480 160.000 ;
        RECT 37.980 159.600 40.280 160.000 ;
        RECT 49.180 159.600 51.480 160.000 ;
        RECT 57.980 159.600 60.280 160.000 ;
        RECT 69.180 159.600 71.480 160.000 ;
        RECT 77.980 159.600 80.280 160.000 ;
        RECT 89.180 159.600 91.480 160.000 ;
        RECT 97.980 159.600 100.280 160.000 ;
        RECT 5.130 159.200 24.330 159.600 ;
        RECT 2.515 157.220 2.875 157.600 ;
        RECT 3.145 157.220 3.505 157.600 ;
        RECT 3.745 157.220 4.105 157.600 ;
        RECT 2.515 156.630 2.875 157.010 ;
        RECT 3.145 156.630 3.505 157.010 ;
        RECT 3.745 156.630 4.105 157.010 ;
        RECT 2.425 155.550 4.235 155.555 ;
        RECT 5.130 155.550 5.530 159.200 ;
        RECT 9.180 159.150 11.480 159.200 ;
        RECT 17.980 159.150 20.280 159.200 ;
        RECT 6.530 158.000 22.930 158.600 ;
        RECT 10.130 157.400 10.480 158.000 ;
        RECT 6.530 157.200 10.480 157.400 ;
        RECT 10.130 156.600 10.480 157.200 ;
        RECT 6.530 156.400 10.480 156.600 ;
        RECT 10.130 155.800 10.480 156.400 ;
        RECT 6.530 155.600 10.480 155.800 ;
        RECT 2.315 153.255 5.580 155.550 ;
        RECT 10.130 155.000 10.480 155.600 ;
        RECT 6.530 154.800 10.480 155.000 ;
        RECT 10.130 154.200 10.480 154.800 ;
        RECT 6.530 154.000 10.480 154.200 ;
        RECT 10.130 153.400 10.480 154.000 ;
        RECT 4.730 153.250 5.580 153.255 ;
        RECT 5.130 146.750 5.530 153.250 ;
        RECT 6.530 153.200 10.480 153.400 ;
        RECT 10.130 152.600 10.480 153.200 ;
        RECT 6.530 152.400 10.480 152.600 ;
        RECT 10.130 151.800 10.480 152.400 ;
        RECT 6.530 151.600 10.480 151.800 ;
        RECT 10.130 151.000 10.480 151.600 ;
        RECT 6.530 150.800 10.480 151.000 ;
        RECT 10.130 150.400 10.480 150.800 ;
        RECT 11.080 150.400 11.280 158.000 ;
        RECT 11.880 150.400 12.080 158.000 ;
        RECT 12.680 150.400 12.880 158.000 ;
        RECT 13.480 150.400 13.680 158.000 ;
        RECT 10.130 149.200 10.480 149.600 ;
        RECT 6.530 149.000 10.480 149.200 ;
        RECT 10.130 148.400 10.480 149.000 ;
        RECT 6.530 148.200 10.480 148.400 ;
        RECT 10.130 147.600 10.480 148.200 ;
        RECT 6.530 147.400 10.480 147.600 ;
        RECT 10.130 146.800 10.480 147.400 ;
        RECT 2.315 144.450 5.580 146.750 ;
        RECT 6.530 146.600 10.480 146.800 ;
        RECT 10.130 146.000 10.480 146.600 ;
        RECT 6.530 145.800 10.480 146.000 ;
        RECT 10.130 145.200 10.480 145.800 ;
        RECT 6.530 145.000 10.480 145.200 ;
        RECT 2.515 142.660 2.875 143.040 ;
        RECT 3.145 142.660 3.505 143.040 ;
        RECT 3.745 142.660 4.105 143.040 ;
        RECT 2.515 142.070 2.875 142.450 ;
        RECT 3.145 142.070 3.505 142.450 ;
        RECT 3.745 142.070 4.105 142.450 ;
        RECT 5.130 140.800 5.530 144.450 ;
        RECT 10.130 144.400 10.480 145.000 ;
        RECT 6.530 144.200 10.480 144.400 ;
        RECT 10.130 143.600 10.480 144.200 ;
        RECT 6.530 143.400 10.480 143.600 ;
        RECT 10.130 142.800 10.480 143.400 ;
        RECT 6.530 142.600 10.480 142.800 ;
        RECT 10.130 142.000 10.480 142.600 ;
        RECT 11.080 142.000 11.280 149.600 ;
        RECT 11.880 142.000 12.080 149.600 ;
        RECT 12.680 142.000 12.880 149.600 ;
        RECT 13.480 142.000 13.680 149.600 ;
        RECT 14.280 142.000 15.180 158.000 ;
        RECT 15.780 150.400 15.980 158.000 ;
        RECT 16.580 150.400 16.780 158.000 ;
        RECT 17.380 150.400 17.580 158.000 ;
        RECT 18.180 150.400 18.380 158.000 ;
        RECT 18.980 157.400 19.330 158.000 ;
        RECT 18.980 157.200 22.930 157.400 ;
        RECT 18.980 156.600 19.330 157.200 ;
        RECT 18.980 156.400 22.930 156.600 ;
        RECT 18.980 155.800 19.330 156.400 ;
        RECT 18.980 155.600 22.930 155.800 ;
        RECT 18.980 155.000 19.330 155.600 ;
        RECT 23.930 155.550 24.330 159.200 ;
        RECT 25.130 159.200 44.330 159.600 ;
        RECT 25.130 155.550 25.530 159.200 ;
        RECT 29.180 159.150 31.480 159.200 ;
        RECT 37.980 159.150 40.280 159.200 ;
        RECT 26.530 158.000 42.930 158.600 ;
        RECT 30.130 157.400 30.480 158.000 ;
        RECT 26.530 157.200 30.480 157.400 ;
        RECT 30.130 156.600 30.480 157.200 ;
        RECT 26.530 156.400 30.480 156.600 ;
        RECT 30.130 155.800 30.480 156.400 ;
        RECT 26.530 155.600 30.480 155.800 ;
        RECT 18.980 154.800 22.930 155.000 ;
        RECT 18.980 154.200 19.330 154.800 ;
        RECT 18.980 154.000 22.930 154.200 ;
        RECT 18.980 153.400 19.330 154.000 ;
        RECT 18.980 153.200 22.930 153.400 ;
        RECT 23.880 153.250 25.580 155.550 ;
        RECT 30.130 155.000 30.480 155.600 ;
        RECT 26.530 154.800 30.480 155.000 ;
        RECT 30.130 154.200 30.480 154.800 ;
        RECT 26.530 154.000 30.480 154.200 ;
        RECT 30.130 153.400 30.480 154.000 ;
        RECT 18.980 152.600 19.330 153.200 ;
        RECT 18.980 152.400 22.930 152.600 ;
        RECT 18.980 151.800 19.330 152.400 ;
        RECT 18.980 151.600 22.930 151.800 ;
        RECT 18.980 151.000 19.330 151.600 ;
        RECT 18.980 150.800 22.930 151.000 ;
        RECT 18.980 150.400 19.330 150.800 ;
        RECT 15.780 142.000 15.980 149.600 ;
        RECT 16.580 142.000 16.780 149.600 ;
        RECT 17.380 142.000 17.580 149.600 ;
        RECT 18.180 142.000 18.380 149.600 ;
        RECT 18.980 149.200 19.330 149.600 ;
        RECT 18.980 149.000 22.930 149.200 ;
        RECT 18.980 148.400 19.330 149.000 ;
        RECT 18.980 148.200 22.930 148.400 ;
        RECT 18.980 147.600 19.330 148.200 ;
        RECT 18.980 147.400 22.930 147.600 ;
        RECT 18.980 146.800 19.330 147.400 ;
        RECT 18.980 146.600 22.930 146.800 ;
        RECT 23.930 146.750 24.330 153.250 ;
        RECT 25.130 146.750 25.530 153.250 ;
        RECT 26.530 153.200 30.480 153.400 ;
        RECT 30.130 152.600 30.480 153.200 ;
        RECT 26.530 152.400 30.480 152.600 ;
        RECT 30.130 151.800 30.480 152.400 ;
        RECT 26.530 151.600 30.480 151.800 ;
        RECT 30.130 151.000 30.480 151.600 ;
        RECT 26.530 150.800 30.480 151.000 ;
        RECT 30.130 150.400 30.480 150.800 ;
        RECT 31.080 150.400 31.280 158.000 ;
        RECT 31.880 150.400 32.080 158.000 ;
        RECT 32.680 150.400 32.880 158.000 ;
        RECT 33.480 150.400 33.680 158.000 ;
        RECT 30.130 149.200 30.480 149.600 ;
        RECT 26.530 149.000 30.480 149.200 ;
        RECT 30.130 148.400 30.480 149.000 ;
        RECT 26.530 148.200 30.480 148.400 ;
        RECT 30.130 147.600 30.480 148.200 ;
        RECT 26.530 147.400 30.480 147.600 ;
        RECT 30.130 146.800 30.480 147.400 ;
        RECT 18.980 146.000 19.330 146.600 ;
        RECT 18.980 145.800 22.930 146.000 ;
        RECT 18.980 145.200 19.330 145.800 ;
        RECT 18.980 145.000 22.930 145.200 ;
        RECT 18.980 144.400 19.330 145.000 ;
        RECT 23.880 144.450 25.580 146.750 ;
        RECT 26.530 146.600 30.480 146.800 ;
        RECT 30.130 146.000 30.480 146.600 ;
        RECT 26.530 145.800 30.480 146.000 ;
        RECT 30.130 145.200 30.480 145.800 ;
        RECT 26.530 145.000 30.480 145.200 ;
        RECT 18.980 144.200 22.930 144.400 ;
        RECT 18.980 143.600 19.330 144.200 ;
        RECT 18.980 143.400 22.930 143.600 ;
        RECT 18.980 142.800 19.330 143.400 ;
        RECT 18.980 142.600 22.930 142.800 ;
        RECT 18.980 142.000 19.330 142.600 ;
        RECT 6.530 141.400 22.930 142.000 ;
        RECT 9.180 140.800 11.480 140.850 ;
        RECT 17.980 140.800 20.280 140.850 ;
        RECT 23.930 140.800 24.330 144.450 ;
        RECT 5.130 140.400 24.330 140.800 ;
        RECT 25.130 140.800 25.530 144.450 ;
        RECT 30.130 144.400 30.480 145.000 ;
        RECT 26.530 144.200 30.480 144.400 ;
        RECT 30.130 143.600 30.480 144.200 ;
        RECT 26.530 143.400 30.480 143.600 ;
        RECT 30.130 142.800 30.480 143.400 ;
        RECT 26.530 142.600 30.480 142.800 ;
        RECT 30.130 142.000 30.480 142.600 ;
        RECT 31.080 142.000 31.280 149.600 ;
        RECT 31.880 142.000 32.080 149.600 ;
        RECT 32.680 142.000 32.880 149.600 ;
        RECT 33.480 142.000 33.680 149.600 ;
        RECT 34.280 142.000 35.180 158.000 ;
        RECT 35.780 150.400 35.980 158.000 ;
        RECT 36.580 150.400 36.780 158.000 ;
        RECT 37.380 150.400 37.580 158.000 ;
        RECT 38.180 150.400 38.380 158.000 ;
        RECT 38.980 157.400 39.330 158.000 ;
        RECT 38.980 157.200 42.930 157.400 ;
        RECT 38.980 156.600 39.330 157.200 ;
        RECT 38.980 156.400 42.930 156.600 ;
        RECT 38.980 155.800 39.330 156.400 ;
        RECT 38.980 155.600 42.930 155.800 ;
        RECT 38.980 155.000 39.330 155.600 ;
        RECT 43.930 155.550 44.330 159.200 ;
        RECT 45.130 159.200 64.330 159.600 ;
        RECT 45.130 155.550 45.530 159.200 ;
        RECT 49.180 159.150 51.480 159.200 ;
        RECT 57.980 159.150 60.280 159.200 ;
        RECT 46.530 158.000 62.930 158.600 ;
        RECT 50.130 157.400 50.480 158.000 ;
        RECT 46.530 157.200 50.480 157.400 ;
        RECT 50.130 156.600 50.480 157.200 ;
        RECT 46.530 156.400 50.480 156.600 ;
        RECT 50.130 155.800 50.480 156.400 ;
        RECT 46.530 155.600 50.480 155.800 ;
        RECT 38.980 154.800 42.930 155.000 ;
        RECT 38.980 154.200 39.330 154.800 ;
        RECT 38.980 154.000 42.930 154.200 ;
        RECT 38.980 153.400 39.330 154.000 ;
        RECT 38.980 153.200 42.930 153.400 ;
        RECT 43.880 153.250 45.580 155.550 ;
        RECT 50.130 155.000 50.480 155.600 ;
        RECT 46.530 154.800 50.480 155.000 ;
        RECT 50.130 154.200 50.480 154.800 ;
        RECT 46.530 154.000 50.480 154.200 ;
        RECT 50.130 153.400 50.480 154.000 ;
        RECT 38.980 152.600 39.330 153.200 ;
        RECT 38.980 152.400 42.930 152.600 ;
        RECT 38.980 151.800 39.330 152.400 ;
        RECT 38.980 151.600 42.930 151.800 ;
        RECT 38.980 151.000 39.330 151.600 ;
        RECT 38.980 150.800 42.930 151.000 ;
        RECT 38.980 150.400 39.330 150.800 ;
        RECT 35.780 142.000 35.980 149.600 ;
        RECT 36.580 142.000 36.780 149.600 ;
        RECT 37.380 142.000 37.580 149.600 ;
        RECT 38.180 142.000 38.380 149.600 ;
        RECT 38.980 149.200 39.330 149.600 ;
        RECT 38.980 149.000 42.930 149.200 ;
        RECT 38.980 148.400 39.330 149.000 ;
        RECT 38.980 148.200 42.930 148.400 ;
        RECT 38.980 147.600 39.330 148.200 ;
        RECT 38.980 147.400 42.930 147.600 ;
        RECT 38.980 146.800 39.330 147.400 ;
        RECT 38.980 146.600 42.930 146.800 ;
        RECT 43.930 146.750 44.330 153.250 ;
        RECT 45.130 146.750 45.530 153.250 ;
        RECT 46.530 153.200 50.480 153.400 ;
        RECT 50.130 152.600 50.480 153.200 ;
        RECT 46.530 152.400 50.480 152.600 ;
        RECT 50.130 151.800 50.480 152.400 ;
        RECT 46.530 151.600 50.480 151.800 ;
        RECT 50.130 151.000 50.480 151.600 ;
        RECT 46.530 150.800 50.480 151.000 ;
        RECT 50.130 150.400 50.480 150.800 ;
        RECT 51.080 150.400 51.280 158.000 ;
        RECT 51.880 150.400 52.080 158.000 ;
        RECT 52.680 150.400 52.880 158.000 ;
        RECT 53.480 150.400 53.680 158.000 ;
        RECT 50.130 149.200 50.480 149.600 ;
        RECT 46.530 149.000 50.480 149.200 ;
        RECT 50.130 148.400 50.480 149.000 ;
        RECT 46.530 148.200 50.480 148.400 ;
        RECT 50.130 147.600 50.480 148.200 ;
        RECT 46.530 147.400 50.480 147.600 ;
        RECT 50.130 146.800 50.480 147.400 ;
        RECT 38.980 146.000 39.330 146.600 ;
        RECT 38.980 145.800 42.930 146.000 ;
        RECT 38.980 145.200 39.330 145.800 ;
        RECT 38.980 145.000 42.930 145.200 ;
        RECT 38.980 144.400 39.330 145.000 ;
        RECT 43.880 144.450 45.580 146.750 ;
        RECT 46.530 146.600 50.480 146.800 ;
        RECT 50.130 146.000 50.480 146.600 ;
        RECT 46.530 145.800 50.480 146.000 ;
        RECT 50.130 145.200 50.480 145.800 ;
        RECT 46.530 145.000 50.480 145.200 ;
        RECT 38.980 144.200 42.930 144.400 ;
        RECT 38.980 143.600 39.330 144.200 ;
        RECT 38.980 143.400 42.930 143.600 ;
        RECT 38.980 142.800 39.330 143.400 ;
        RECT 38.980 142.600 42.930 142.800 ;
        RECT 38.980 142.000 39.330 142.600 ;
        RECT 26.530 141.400 42.930 142.000 ;
        RECT 29.180 140.800 31.480 140.850 ;
        RECT 37.980 140.800 40.280 140.850 ;
        RECT 43.930 140.800 44.330 144.450 ;
        RECT 25.130 140.400 44.330 140.800 ;
        RECT 45.130 140.800 45.530 144.450 ;
        RECT 50.130 144.400 50.480 145.000 ;
        RECT 46.530 144.200 50.480 144.400 ;
        RECT 50.130 143.600 50.480 144.200 ;
        RECT 46.530 143.400 50.480 143.600 ;
        RECT 50.130 142.800 50.480 143.400 ;
        RECT 46.530 142.600 50.480 142.800 ;
        RECT 50.130 142.000 50.480 142.600 ;
        RECT 51.080 142.000 51.280 149.600 ;
        RECT 51.880 142.000 52.080 149.600 ;
        RECT 52.680 142.000 52.880 149.600 ;
        RECT 53.480 142.000 53.680 149.600 ;
        RECT 54.280 142.000 55.180 158.000 ;
        RECT 55.780 150.400 55.980 158.000 ;
        RECT 56.580 150.400 56.780 158.000 ;
        RECT 57.380 150.400 57.580 158.000 ;
        RECT 58.180 150.400 58.380 158.000 ;
        RECT 58.980 157.400 59.330 158.000 ;
        RECT 58.980 157.200 62.930 157.400 ;
        RECT 58.980 156.600 59.330 157.200 ;
        RECT 58.980 156.400 62.930 156.600 ;
        RECT 58.980 155.800 59.330 156.400 ;
        RECT 58.980 155.600 62.930 155.800 ;
        RECT 58.980 155.000 59.330 155.600 ;
        RECT 63.930 155.550 64.330 159.200 ;
        RECT 65.130 159.200 84.330 159.600 ;
        RECT 65.130 155.550 65.530 159.200 ;
        RECT 69.180 159.150 71.480 159.200 ;
        RECT 77.980 159.150 80.280 159.200 ;
        RECT 66.530 158.000 82.930 158.600 ;
        RECT 70.130 157.400 70.480 158.000 ;
        RECT 66.530 157.200 70.480 157.400 ;
        RECT 70.130 156.600 70.480 157.200 ;
        RECT 66.530 156.400 70.480 156.600 ;
        RECT 70.130 155.800 70.480 156.400 ;
        RECT 66.530 155.600 70.480 155.800 ;
        RECT 58.980 154.800 62.930 155.000 ;
        RECT 58.980 154.200 59.330 154.800 ;
        RECT 58.980 154.000 62.930 154.200 ;
        RECT 58.980 153.400 59.330 154.000 ;
        RECT 58.980 153.200 62.930 153.400 ;
        RECT 63.880 153.250 65.580 155.550 ;
        RECT 70.130 155.000 70.480 155.600 ;
        RECT 66.530 154.800 70.480 155.000 ;
        RECT 70.130 154.200 70.480 154.800 ;
        RECT 66.530 154.000 70.480 154.200 ;
        RECT 70.130 153.400 70.480 154.000 ;
        RECT 58.980 152.600 59.330 153.200 ;
        RECT 58.980 152.400 62.930 152.600 ;
        RECT 58.980 151.800 59.330 152.400 ;
        RECT 58.980 151.600 62.930 151.800 ;
        RECT 58.980 151.000 59.330 151.600 ;
        RECT 58.980 150.800 62.930 151.000 ;
        RECT 58.980 150.400 59.330 150.800 ;
        RECT 55.780 142.000 55.980 149.600 ;
        RECT 56.580 142.000 56.780 149.600 ;
        RECT 57.380 142.000 57.580 149.600 ;
        RECT 58.180 142.000 58.380 149.600 ;
        RECT 58.980 149.200 59.330 149.600 ;
        RECT 58.980 149.000 62.930 149.200 ;
        RECT 58.980 148.400 59.330 149.000 ;
        RECT 58.980 148.200 62.930 148.400 ;
        RECT 58.980 147.600 59.330 148.200 ;
        RECT 58.980 147.400 62.930 147.600 ;
        RECT 58.980 146.800 59.330 147.400 ;
        RECT 58.980 146.600 62.930 146.800 ;
        RECT 63.930 146.750 64.330 153.250 ;
        RECT 65.130 146.750 65.530 153.250 ;
        RECT 66.530 153.200 70.480 153.400 ;
        RECT 70.130 152.600 70.480 153.200 ;
        RECT 66.530 152.400 70.480 152.600 ;
        RECT 70.130 151.800 70.480 152.400 ;
        RECT 66.530 151.600 70.480 151.800 ;
        RECT 70.130 151.000 70.480 151.600 ;
        RECT 66.530 150.800 70.480 151.000 ;
        RECT 70.130 150.400 70.480 150.800 ;
        RECT 71.080 150.400 71.280 158.000 ;
        RECT 71.880 150.400 72.080 158.000 ;
        RECT 72.680 150.400 72.880 158.000 ;
        RECT 73.480 150.400 73.680 158.000 ;
        RECT 70.130 149.200 70.480 149.600 ;
        RECT 66.530 149.000 70.480 149.200 ;
        RECT 70.130 148.400 70.480 149.000 ;
        RECT 66.530 148.200 70.480 148.400 ;
        RECT 70.130 147.600 70.480 148.200 ;
        RECT 66.530 147.400 70.480 147.600 ;
        RECT 70.130 146.800 70.480 147.400 ;
        RECT 58.980 146.000 59.330 146.600 ;
        RECT 58.980 145.800 62.930 146.000 ;
        RECT 58.980 145.200 59.330 145.800 ;
        RECT 58.980 145.000 62.930 145.200 ;
        RECT 58.980 144.400 59.330 145.000 ;
        RECT 63.880 144.450 65.580 146.750 ;
        RECT 66.530 146.600 70.480 146.800 ;
        RECT 70.130 146.000 70.480 146.600 ;
        RECT 66.530 145.800 70.480 146.000 ;
        RECT 70.130 145.200 70.480 145.800 ;
        RECT 66.530 145.000 70.480 145.200 ;
        RECT 58.980 144.200 62.930 144.400 ;
        RECT 58.980 143.600 59.330 144.200 ;
        RECT 58.980 143.400 62.930 143.600 ;
        RECT 58.980 142.800 59.330 143.400 ;
        RECT 58.980 142.600 62.930 142.800 ;
        RECT 58.980 142.000 59.330 142.600 ;
        RECT 46.530 141.400 62.930 142.000 ;
        RECT 49.180 140.800 51.480 140.850 ;
        RECT 57.980 140.800 60.280 140.850 ;
        RECT 63.930 140.800 64.330 144.450 ;
        RECT 45.130 140.400 64.330 140.800 ;
        RECT 65.130 140.800 65.530 144.450 ;
        RECT 70.130 144.400 70.480 145.000 ;
        RECT 66.530 144.200 70.480 144.400 ;
        RECT 70.130 143.600 70.480 144.200 ;
        RECT 66.530 143.400 70.480 143.600 ;
        RECT 70.130 142.800 70.480 143.400 ;
        RECT 66.530 142.600 70.480 142.800 ;
        RECT 70.130 142.000 70.480 142.600 ;
        RECT 71.080 142.000 71.280 149.600 ;
        RECT 71.880 142.000 72.080 149.600 ;
        RECT 72.680 142.000 72.880 149.600 ;
        RECT 73.480 142.000 73.680 149.600 ;
        RECT 74.280 142.000 75.180 158.000 ;
        RECT 75.780 150.400 75.980 158.000 ;
        RECT 76.580 150.400 76.780 158.000 ;
        RECT 77.380 150.400 77.580 158.000 ;
        RECT 78.180 150.400 78.380 158.000 ;
        RECT 78.980 157.400 79.330 158.000 ;
        RECT 78.980 157.200 82.930 157.400 ;
        RECT 78.980 156.600 79.330 157.200 ;
        RECT 78.980 156.400 82.930 156.600 ;
        RECT 78.980 155.800 79.330 156.400 ;
        RECT 78.980 155.600 82.930 155.800 ;
        RECT 78.980 155.000 79.330 155.600 ;
        RECT 83.930 155.550 84.330 159.200 ;
        RECT 85.130 159.200 104.330 159.600 ;
        RECT 85.130 155.550 85.530 159.200 ;
        RECT 89.180 159.150 91.480 159.200 ;
        RECT 97.980 159.150 100.280 159.200 ;
        RECT 86.530 158.000 102.930 158.600 ;
        RECT 90.130 157.400 90.480 158.000 ;
        RECT 86.530 157.200 90.480 157.400 ;
        RECT 90.130 156.600 90.480 157.200 ;
        RECT 86.530 156.400 90.480 156.600 ;
        RECT 90.130 155.800 90.480 156.400 ;
        RECT 86.530 155.600 90.480 155.800 ;
        RECT 78.980 154.800 82.930 155.000 ;
        RECT 78.980 154.200 79.330 154.800 ;
        RECT 78.980 154.000 82.930 154.200 ;
        RECT 78.980 153.400 79.330 154.000 ;
        RECT 78.980 153.200 82.930 153.400 ;
        RECT 83.880 153.250 85.580 155.550 ;
        RECT 90.130 155.000 90.480 155.600 ;
        RECT 86.530 154.800 90.480 155.000 ;
        RECT 90.130 154.200 90.480 154.800 ;
        RECT 86.530 154.000 90.480 154.200 ;
        RECT 90.130 153.400 90.480 154.000 ;
        RECT 78.980 152.600 79.330 153.200 ;
        RECT 78.980 152.400 82.930 152.600 ;
        RECT 78.980 151.800 79.330 152.400 ;
        RECT 78.980 151.600 82.930 151.800 ;
        RECT 78.980 151.000 79.330 151.600 ;
        RECT 78.980 150.800 82.930 151.000 ;
        RECT 78.980 150.400 79.330 150.800 ;
        RECT 75.780 142.000 75.980 149.600 ;
        RECT 76.580 142.000 76.780 149.600 ;
        RECT 77.380 142.000 77.580 149.600 ;
        RECT 78.180 142.000 78.380 149.600 ;
        RECT 78.980 149.200 79.330 149.600 ;
        RECT 78.980 149.000 82.930 149.200 ;
        RECT 78.980 148.400 79.330 149.000 ;
        RECT 78.980 148.200 82.930 148.400 ;
        RECT 78.980 147.600 79.330 148.200 ;
        RECT 78.980 147.400 82.930 147.600 ;
        RECT 78.980 146.800 79.330 147.400 ;
        RECT 78.980 146.600 82.930 146.800 ;
        RECT 83.930 146.750 84.330 153.250 ;
        RECT 85.130 146.750 85.530 153.250 ;
        RECT 86.530 153.200 90.480 153.400 ;
        RECT 90.130 152.600 90.480 153.200 ;
        RECT 86.530 152.400 90.480 152.600 ;
        RECT 90.130 151.800 90.480 152.400 ;
        RECT 86.530 151.600 90.480 151.800 ;
        RECT 90.130 151.000 90.480 151.600 ;
        RECT 86.530 150.800 90.480 151.000 ;
        RECT 90.130 150.400 90.480 150.800 ;
        RECT 91.080 150.400 91.280 158.000 ;
        RECT 91.880 150.400 92.080 158.000 ;
        RECT 92.680 150.400 92.880 158.000 ;
        RECT 93.480 150.400 93.680 158.000 ;
        RECT 90.130 149.200 90.480 149.600 ;
        RECT 86.530 149.000 90.480 149.200 ;
        RECT 90.130 148.400 90.480 149.000 ;
        RECT 86.530 148.200 90.480 148.400 ;
        RECT 90.130 147.600 90.480 148.200 ;
        RECT 86.530 147.400 90.480 147.600 ;
        RECT 90.130 146.800 90.480 147.400 ;
        RECT 78.980 146.000 79.330 146.600 ;
        RECT 78.980 145.800 82.930 146.000 ;
        RECT 78.980 145.200 79.330 145.800 ;
        RECT 78.980 145.000 82.930 145.200 ;
        RECT 78.980 144.400 79.330 145.000 ;
        RECT 83.880 144.450 85.580 146.750 ;
        RECT 86.530 146.600 90.480 146.800 ;
        RECT 90.130 146.000 90.480 146.600 ;
        RECT 86.530 145.800 90.480 146.000 ;
        RECT 90.130 145.200 90.480 145.800 ;
        RECT 86.530 145.000 90.480 145.200 ;
        RECT 78.980 144.200 82.930 144.400 ;
        RECT 78.980 143.600 79.330 144.200 ;
        RECT 78.980 143.400 82.930 143.600 ;
        RECT 78.980 142.800 79.330 143.400 ;
        RECT 78.980 142.600 82.930 142.800 ;
        RECT 78.980 142.000 79.330 142.600 ;
        RECT 66.530 141.400 82.930 142.000 ;
        RECT 69.180 140.800 71.480 140.850 ;
        RECT 77.980 140.800 80.280 140.850 ;
        RECT 83.930 140.800 84.330 144.450 ;
        RECT 65.130 140.400 84.330 140.800 ;
        RECT 85.130 140.800 85.530 144.450 ;
        RECT 90.130 144.400 90.480 145.000 ;
        RECT 86.530 144.200 90.480 144.400 ;
        RECT 90.130 143.600 90.480 144.200 ;
        RECT 86.530 143.400 90.480 143.600 ;
        RECT 90.130 142.800 90.480 143.400 ;
        RECT 86.530 142.600 90.480 142.800 ;
        RECT 90.130 142.000 90.480 142.600 ;
        RECT 91.080 142.000 91.280 149.600 ;
        RECT 91.880 142.000 92.080 149.600 ;
        RECT 92.680 142.000 92.880 149.600 ;
        RECT 93.480 142.000 93.680 149.600 ;
        RECT 94.280 142.000 95.180 158.000 ;
        RECT 95.780 150.400 95.980 158.000 ;
        RECT 96.580 150.400 96.780 158.000 ;
        RECT 97.380 150.400 97.580 158.000 ;
        RECT 98.180 150.400 98.380 158.000 ;
        RECT 98.980 157.400 99.330 158.000 ;
        RECT 98.980 157.200 102.930 157.400 ;
        RECT 98.980 156.600 99.330 157.200 ;
        RECT 98.980 156.400 102.930 156.600 ;
        RECT 98.980 155.800 99.330 156.400 ;
        RECT 98.980 155.600 102.930 155.800 ;
        RECT 98.980 155.000 99.330 155.600 ;
        RECT 103.930 155.550 104.330 159.200 ;
        RECT 105.340 157.220 105.700 157.600 ;
        RECT 105.970 157.220 106.330 157.600 ;
        RECT 106.570 157.220 106.930 157.600 ;
        RECT 105.340 156.630 105.700 157.010 ;
        RECT 105.970 156.630 106.330 157.010 ;
        RECT 106.570 156.630 106.930 157.010 ;
        RECT 98.980 154.800 102.930 155.000 ;
        RECT 98.980 154.200 99.330 154.800 ;
        RECT 98.980 154.000 102.930 154.200 ;
        RECT 98.980 153.400 99.330 154.000 ;
        RECT 98.980 153.200 102.930 153.400 ;
        RECT 103.880 153.250 104.730 155.550 ;
        RECT 98.980 152.600 99.330 153.200 ;
        RECT 98.980 152.400 102.930 152.600 ;
        RECT 98.980 151.800 99.330 152.400 ;
        RECT 98.980 151.600 102.930 151.800 ;
        RECT 98.980 151.000 99.330 151.600 ;
        RECT 98.980 150.800 102.930 151.000 ;
        RECT 98.980 150.400 99.330 150.800 ;
        RECT 95.780 142.000 95.980 149.600 ;
        RECT 96.580 142.000 96.780 149.600 ;
        RECT 97.380 142.000 97.580 149.600 ;
        RECT 98.180 142.000 98.380 149.600 ;
        RECT 98.980 149.200 99.330 149.600 ;
        RECT 98.980 149.000 102.930 149.200 ;
        RECT 98.980 148.400 99.330 149.000 ;
        RECT 98.980 148.200 102.930 148.400 ;
        RECT 98.980 147.600 99.330 148.200 ;
        RECT 98.980 147.400 102.930 147.600 ;
        RECT 98.980 146.800 99.330 147.400 ;
        RECT 98.980 146.600 102.930 146.800 ;
        RECT 103.930 146.750 104.330 153.250 ;
        RECT 98.980 146.000 99.330 146.600 ;
        RECT 98.980 145.800 102.930 146.000 ;
        RECT 98.980 145.200 99.330 145.800 ;
        RECT 98.980 145.000 102.930 145.200 ;
        RECT 98.980 144.400 99.330 145.000 ;
        RECT 103.880 144.450 104.730 146.750 ;
        RECT 98.980 144.200 102.930 144.400 ;
        RECT 98.980 143.600 99.330 144.200 ;
        RECT 98.980 143.400 102.930 143.600 ;
        RECT 98.980 142.800 99.330 143.400 ;
        RECT 98.980 142.600 102.930 142.800 ;
        RECT 98.980 142.000 99.330 142.600 ;
        RECT 86.530 141.400 102.930 142.000 ;
        RECT 89.180 140.800 91.480 140.850 ;
        RECT 97.980 140.800 100.280 140.850 ;
        RECT 103.930 140.800 104.330 144.450 ;
        RECT 105.340 142.415 105.700 142.795 ;
        RECT 105.970 142.415 106.330 142.795 ;
        RECT 106.570 142.415 106.930 142.795 ;
        RECT 105.340 141.825 105.700 142.205 ;
        RECT 105.970 141.825 106.330 142.205 ;
        RECT 106.570 141.825 106.930 142.205 ;
        RECT 85.130 140.400 104.330 140.800 ;
        RECT 9.180 139.600 11.480 140.400 ;
        RECT 17.980 139.600 20.280 140.400 ;
        RECT 29.180 139.600 31.480 140.400 ;
        RECT 37.980 139.600 40.280 140.400 ;
        RECT 49.180 139.600 51.480 140.400 ;
        RECT 57.980 139.600 60.280 140.400 ;
        RECT 69.180 139.600 71.480 140.400 ;
        RECT 77.980 139.600 80.280 140.400 ;
        RECT 89.180 139.600 91.480 140.400 ;
        RECT 97.980 139.600 100.280 140.400 ;
        RECT 5.130 139.200 24.330 139.600 ;
        RECT 2.515 137.640 2.875 138.020 ;
        RECT 3.145 137.640 3.505 138.020 ;
        RECT 3.745 137.640 4.105 138.020 ;
        RECT 2.515 137.050 2.875 137.430 ;
        RECT 3.145 137.050 3.505 137.430 ;
        RECT 3.745 137.050 4.105 137.430 ;
        RECT 5.130 135.550 5.530 139.200 ;
        RECT 9.180 139.150 11.480 139.200 ;
        RECT 17.980 139.150 20.280 139.200 ;
        RECT 6.530 138.000 22.930 138.600 ;
        RECT 10.130 137.400 10.480 138.000 ;
        RECT 6.530 137.200 10.480 137.400 ;
        RECT 10.130 136.600 10.480 137.200 ;
        RECT 6.530 136.400 10.480 136.600 ;
        RECT 10.130 135.800 10.480 136.400 ;
        RECT 6.530 135.600 10.480 135.800 ;
        RECT 4.730 135.545 5.580 135.550 ;
        RECT 2.315 133.250 5.580 135.545 ;
        RECT 10.130 135.000 10.480 135.600 ;
        RECT 6.530 134.800 10.480 135.000 ;
        RECT 10.130 134.200 10.480 134.800 ;
        RECT 6.530 134.000 10.480 134.200 ;
        RECT 10.130 133.400 10.480 134.000 ;
        RECT 5.130 126.750 5.530 133.250 ;
        RECT 6.530 133.200 10.480 133.400 ;
        RECT 10.130 132.600 10.480 133.200 ;
        RECT 6.530 132.400 10.480 132.600 ;
        RECT 10.130 131.800 10.480 132.400 ;
        RECT 6.530 131.600 10.480 131.800 ;
        RECT 10.130 131.000 10.480 131.600 ;
        RECT 6.530 130.800 10.480 131.000 ;
        RECT 10.130 130.400 10.480 130.800 ;
        RECT 11.080 130.400 11.280 138.000 ;
        RECT 11.880 130.400 12.080 138.000 ;
        RECT 12.680 130.400 12.880 138.000 ;
        RECT 13.480 130.400 13.680 138.000 ;
        RECT 10.130 129.200 10.480 129.600 ;
        RECT 6.530 129.000 10.480 129.200 ;
        RECT 10.130 128.400 10.480 129.000 ;
        RECT 6.530 128.200 10.480 128.400 ;
        RECT 10.130 127.600 10.480 128.200 ;
        RECT 6.530 127.400 10.480 127.600 ;
        RECT 10.130 126.800 10.480 127.400 ;
        RECT 4.730 126.745 5.580 126.750 ;
        RECT 2.315 124.450 5.580 126.745 ;
        RECT 6.530 126.600 10.480 126.800 ;
        RECT 10.130 126.000 10.480 126.600 ;
        RECT 6.530 125.800 10.480 126.000 ;
        RECT 10.130 125.200 10.480 125.800 ;
        RECT 6.530 125.000 10.480 125.200 ;
        RECT 2.515 122.750 2.875 123.130 ;
        RECT 3.145 122.750 3.505 123.130 ;
        RECT 3.745 122.750 4.105 123.130 ;
        RECT 2.515 122.160 2.875 122.540 ;
        RECT 3.145 122.160 3.505 122.540 ;
        RECT 3.745 122.160 4.105 122.540 ;
        RECT 5.130 120.800 5.530 124.450 ;
        RECT 10.130 124.400 10.480 125.000 ;
        RECT 6.530 124.200 10.480 124.400 ;
        RECT 10.130 123.600 10.480 124.200 ;
        RECT 6.530 123.400 10.480 123.600 ;
        RECT 10.130 122.800 10.480 123.400 ;
        RECT 6.530 122.600 10.480 122.800 ;
        RECT 10.130 122.000 10.480 122.600 ;
        RECT 11.080 122.000 11.280 129.600 ;
        RECT 11.880 122.000 12.080 129.600 ;
        RECT 12.680 122.000 12.880 129.600 ;
        RECT 13.480 122.000 13.680 129.600 ;
        RECT 14.280 122.000 15.180 138.000 ;
        RECT 15.780 130.400 15.980 138.000 ;
        RECT 16.580 130.400 16.780 138.000 ;
        RECT 17.380 130.400 17.580 138.000 ;
        RECT 18.180 130.400 18.380 138.000 ;
        RECT 18.980 137.400 19.330 138.000 ;
        RECT 18.980 137.200 22.930 137.400 ;
        RECT 18.980 136.600 19.330 137.200 ;
        RECT 18.980 136.400 22.930 136.600 ;
        RECT 18.980 135.800 19.330 136.400 ;
        RECT 18.980 135.600 22.930 135.800 ;
        RECT 18.980 135.000 19.330 135.600 ;
        RECT 23.930 135.550 24.330 139.200 ;
        RECT 25.130 139.200 44.330 139.600 ;
        RECT 25.130 135.550 25.530 139.200 ;
        RECT 29.180 139.150 31.480 139.200 ;
        RECT 37.980 139.150 40.280 139.200 ;
        RECT 26.530 138.000 42.930 138.600 ;
        RECT 30.130 137.400 30.480 138.000 ;
        RECT 26.530 137.200 30.480 137.400 ;
        RECT 30.130 136.600 30.480 137.200 ;
        RECT 26.530 136.400 30.480 136.600 ;
        RECT 30.130 135.800 30.480 136.400 ;
        RECT 26.530 135.600 30.480 135.800 ;
        RECT 18.980 134.800 22.930 135.000 ;
        RECT 18.980 134.200 19.330 134.800 ;
        RECT 18.980 134.000 22.930 134.200 ;
        RECT 18.980 133.400 19.330 134.000 ;
        RECT 18.980 133.200 22.930 133.400 ;
        RECT 23.880 133.250 25.580 135.550 ;
        RECT 30.130 135.000 30.480 135.600 ;
        RECT 26.530 134.800 30.480 135.000 ;
        RECT 30.130 134.200 30.480 134.800 ;
        RECT 26.530 134.000 30.480 134.200 ;
        RECT 30.130 133.400 30.480 134.000 ;
        RECT 18.980 132.600 19.330 133.200 ;
        RECT 18.980 132.400 22.930 132.600 ;
        RECT 18.980 131.800 19.330 132.400 ;
        RECT 18.980 131.600 22.930 131.800 ;
        RECT 18.980 131.000 19.330 131.600 ;
        RECT 18.980 130.800 22.930 131.000 ;
        RECT 18.980 130.400 19.330 130.800 ;
        RECT 15.780 122.000 15.980 129.600 ;
        RECT 16.580 122.000 16.780 129.600 ;
        RECT 17.380 122.000 17.580 129.600 ;
        RECT 18.180 122.000 18.380 129.600 ;
        RECT 18.980 129.200 19.330 129.600 ;
        RECT 18.980 129.000 22.930 129.200 ;
        RECT 18.980 128.400 19.330 129.000 ;
        RECT 18.980 128.200 22.930 128.400 ;
        RECT 18.980 127.600 19.330 128.200 ;
        RECT 18.980 127.400 22.930 127.600 ;
        RECT 18.980 126.800 19.330 127.400 ;
        RECT 18.980 126.600 22.930 126.800 ;
        RECT 23.930 126.750 24.330 133.250 ;
        RECT 25.130 126.750 25.530 133.250 ;
        RECT 26.530 133.200 30.480 133.400 ;
        RECT 30.130 132.600 30.480 133.200 ;
        RECT 26.530 132.400 30.480 132.600 ;
        RECT 30.130 131.800 30.480 132.400 ;
        RECT 26.530 131.600 30.480 131.800 ;
        RECT 30.130 131.000 30.480 131.600 ;
        RECT 26.530 130.800 30.480 131.000 ;
        RECT 30.130 130.400 30.480 130.800 ;
        RECT 31.080 130.400 31.280 138.000 ;
        RECT 31.880 130.400 32.080 138.000 ;
        RECT 32.680 130.400 32.880 138.000 ;
        RECT 33.480 130.400 33.680 138.000 ;
        RECT 30.130 129.200 30.480 129.600 ;
        RECT 26.530 129.000 30.480 129.200 ;
        RECT 30.130 128.400 30.480 129.000 ;
        RECT 26.530 128.200 30.480 128.400 ;
        RECT 30.130 127.600 30.480 128.200 ;
        RECT 26.530 127.400 30.480 127.600 ;
        RECT 30.130 126.800 30.480 127.400 ;
        RECT 18.980 126.000 19.330 126.600 ;
        RECT 18.980 125.800 22.930 126.000 ;
        RECT 18.980 125.200 19.330 125.800 ;
        RECT 18.980 125.000 22.930 125.200 ;
        RECT 18.980 124.400 19.330 125.000 ;
        RECT 23.880 124.450 25.580 126.750 ;
        RECT 26.530 126.600 30.480 126.800 ;
        RECT 30.130 126.000 30.480 126.600 ;
        RECT 26.530 125.800 30.480 126.000 ;
        RECT 30.130 125.200 30.480 125.800 ;
        RECT 26.530 125.000 30.480 125.200 ;
        RECT 18.980 124.200 22.930 124.400 ;
        RECT 18.980 123.600 19.330 124.200 ;
        RECT 18.980 123.400 22.930 123.600 ;
        RECT 18.980 122.800 19.330 123.400 ;
        RECT 18.980 122.600 22.930 122.800 ;
        RECT 18.980 122.000 19.330 122.600 ;
        RECT 6.530 121.400 22.930 122.000 ;
        RECT 9.180 120.800 11.480 120.850 ;
        RECT 17.980 120.800 20.280 120.850 ;
        RECT 23.930 120.800 24.330 124.450 ;
        RECT 5.130 120.400 24.330 120.800 ;
        RECT 25.130 120.800 25.530 124.450 ;
        RECT 30.130 124.400 30.480 125.000 ;
        RECT 26.530 124.200 30.480 124.400 ;
        RECT 30.130 123.600 30.480 124.200 ;
        RECT 26.530 123.400 30.480 123.600 ;
        RECT 30.130 122.800 30.480 123.400 ;
        RECT 26.530 122.600 30.480 122.800 ;
        RECT 30.130 122.000 30.480 122.600 ;
        RECT 31.080 122.000 31.280 129.600 ;
        RECT 31.880 122.000 32.080 129.600 ;
        RECT 32.680 122.000 32.880 129.600 ;
        RECT 33.480 122.000 33.680 129.600 ;
        RECT 34.280 122.000 35.180 138.000 ;
        RECT 35.780 130.400 35.980 138.000 ;
        RECT 36.580 130.400 36.780 138.000 ;
        RECT 37.380 130.400 37.580 138.000 ;
        RECT 38.180 130.400 38.380 138.000 ;
        RECT 38.980 137.400 39.330 138.000 ;
        RECT 38.980 137.200 42.930 137.400 ;
        RECT 38.980 136.600 39.330 137.200 ;
        RECT 38.980 136.400 42.930 136.600 ;
        RECT 38.980 135.800 39.330 136.400 ;
        RECT 38.980 135.600 42.930 135.800 ;
        RECT 38.980 135.000 39.330 135.600 ;
        RECT 43.930 135.550 44.330 139.200 ;
        RECT 45.130 139.200 64.330 139.600 ;
        RECT 45.130 135.550 45.530 139.200 ;
        RECT 49.180 139.150 51.480 139.200 ;
        RECT 57.980 139.150 60.280 139.200 ;
        RECT 46.530 138.000 62.930 138.600 ;
        RECT 50.130 137.400 50.480 138.000 ;
        RECT 46.530 137.200 50.480 137.400 ;
        RECT 50.130 136.600 50.480 137.200 ;
        RECT 46.530 136.400 50.480 136.600 ;
        RECT 50.130 135.800 50.480 136.400 ;
        RECT 46.530 135.600 50.480 135.800 ;
        RECT 38.980 134.800 42.930 135.000 ;
        RECT 38.980 134.200 39.330 134.800 ;
        RECT 38.980 134.000 42.930 134.200 ;
        RECT 38.980 133.400 39.330 134.000 ;
        RECT 38.980 133.200 42.930 133.400 ;
        RECT 43.880 133.250 45.580 135.550 ;
        RECT 50.130 135.000 50.480 135.600 ;
        RECT 46.530 134.800 50.480 135.000 ;
        RECT 50.130 134.200 50.480 134.800 ;
        RECT 46.530 134.000 50.480 134.200 ;
        RECT 50.130 133.400 50.480 134.000 ;
        RECT 38.980 132.600 39.330 133.200 ;
        RECT 38.980 132.400 42.930 132.600 ;
        RECT 38.980 131.800 39.330 132.400 ;
        RECT 38.980 131.600 42.930 131.800 ;
        RECT 38.980 131.000 39.330 131.600 ;
        RECT 38.980 130.800 42.930 131.000 ;
        RECT 38.980 130.400 39.330 130.800 ;
        RECT 35.780 122.000 35.980 129.600 ;
        RECT 36.580 122.000 36.780 129.600 ;
        RECT 37.380 122.000 37.580 129.600 ;
        RECT 38.180 122.000 38.380 129.600 ;
        RECT 38.980 129.200 39.330 129.600 ;
        RECT 38.980 129.000 42.930 129.200 ;
        RECT 38.980 128.400 39.330 129.000 ;
        RECT 38.980 128.200 42.930 128.400 ;
        RECT 38.980 127.600 39.330 128.200 ;
        RECT 38.980 127.400 42.930 127.600 ;
        RECT 38.980 126.800 39.330 127.400 ;
        RECT 38.980 126.600 42.930 126.800 ;
        RECT 43.930 126.750 44.330 133.250 ;
        RECT 45.130 126.750 45.530 133.250 ;
        RECT 46.530 133.200 50.480 133.400 ;
        RECT 50.130 132.600 50.480 133.200 ;
        RECT 46.530 132.400 50.480 132.600 ;
        RECT 50.130 131.800 50.480 132.400 ;
        RECT 46.530 131.600 50.480 131.800 ;
        RECT 50.130 131.000 50.480 131.600 ;
        RECT 46.530 130.800 50.480 131.000 ;
        RECT 50.130 130.400 50.480 130.800 ;
        RECT 51.080 130.400 51.280 138.000 ;
        RECT 51.880 130.400 52.080 138.000 ;
        RECT 52.680 130.400 52.880 138.000 ;
        RECT 53.480 130.400 53.680 138.000 ;
        RECT 50.130 129.200 50.480 129.600 ;
        RECT 46.530 129.000 50.480 129.200 ;
        RECT 50.130 128.400 50.480 129.000 ;
        RECT 46.530 128.200 50.480 128.400 ;
        RECT 50.130 127.600 50.480 128.200 ;
        RECT 46.530 127.400 50.480 127.600 ;
        RECT 50.130 126.800 50.480 127.400 ;
        RECT 38.980 126.000 39.330 126.600 ;
        RECT 38.980 125.800 42.930 126.000 ;
        RECT 38.980 125.200 39.330 125.800 ;
        RECT 38.980 125.000 42.930 125.200 ;
        RECT 38.980 124.400 39.330 125.000 ;
        RECT 43.880 124.450 45.580 126.750 ;
        RECT 46.530 126.600 50.480 126.800 ;
        RECT 50.130 126.000 50.480 126.600 ;
        RECT 46.530 125.800 50.480 126.000 ;
        RECT 50.130 125.200 50.480 125.800 ;
        RECT 46.530 125.000 50.480 125.200 ;
        RECT 38.980 124.200 42.930 124.400 ;
        RECT 38.980 123.600 39.330 124.200 ;
        RECT 38.980 123.400 42.930 123.600 ;
        RECT 38.980 122.800 39.330 123.400 ;
        RECT 38.980 122.600 42.930 122.800 ;
        RECT 38.980 122.000 39.330 122.600 ;
        RECT 26.530 121.400 42.930 122.000 ;
        RECT 29.180 120.800 31.480 120.850 ;
        RECT 37.980 120.800 40.280 120.850 ;
        RECT 43.930 120.800 44.330 124.450 ;
        RECT 25.130 120.400 44.330 120.800 ;
        RECT 45.130 120.800 45.530 124.450 ;
        RECT 50.130 124.400 50.480 125.000 ;
        RECT 46.530 124.200 50.480 124.400 ;
        RECT 50.130 123.600 50.480 124.200 ;
        RECT 46.530 123.400 50.480 123.600 ;
        RECT 50.130 122.800 50.480 123.400 ;
        RECT 46.530 122.600 50.480 122.800 ;
        RECT 50.130 122.000 50.480 122.600 ;
        RECT 51.080 122.000 51.280 129.600 ;
        RECT 51.880 122.000 52.080 129.600 ;
        RECT 52.680 122.000 52.880 129.600 ;
        RECT 53.480 122.000 53.680 129.600 ;
        RECT 54.280 122.000 55.180 138.000 ;
        RECT 55.780 130.400 55.980 138.000 ;
        RECT 56.580 130.400 56.780 138.000 ;
        RECT 57.380 130.400 57.580 138.000 ;
        RECT 58.180 130.400 58.380 138.000 ;
        RECT 58.980 137.400 59.330 138.000 ;
        RECT 58.980 137.200 62.930 137.400 ;
        RECT 58.980 136.600 59.330 137.200 ;
        RECT 58.980 136.400 62.930 136.600 ;
        RECT 58.980 135.800 59.330 136.400 ;
        RECT 58.980 135.600 62.930 135.800 ;
        RECT 58.980 135.000 59.330 135.600 ;
        RECT 63.930 135.550 64.330 139.200 ;
        RECT 65.130 139.200 84.330 139.600 ;
        RECT 65.130 135.550 65.530 139.200 ;
        RECT 69.180 139.150 71.480 139.200 ;
        RECT 77.980 139.150 80.280 139.200 ;
        RECT 66.530 138.000 82.930 138.600 ;
        RECT 70.130 137.400 70.480 138.000 ;
        RECT 66.530 137.200 70.480 137.400 ;
        RECT 70.130 136.600 70.480 137.200 ;
        RECT 66.530 136.400 70.480 136.600 ;
        RECT 70.130 135.800 70.480 136.400 ;
        RECT 66.530 135.600 70.480 135.800 ;
        RECT 58.980 134.800 62.930 135.000 ;
        RECT 58.980 134.200 59.330 134.800 ;
        RECT 58.980 134.000 62.930 134.200 ;
        RECT 58.980 133.400 59.330 134.000 ;
        RECT 58.980 133.200 62.930 133.400 ;
        RECT 63.880 133.250 65.580 135.550 ;
        RECT 70.130 135.000 70.480 135.600 ;
        RECT 66.530 134.800 70.480 135.000 ;
        RECT 70.130 134.200 70.480 134.800 ;
        RECT 66.530 134.000 70.480 134.200 ;
        RECT 70.130 133.400 70.480 134.000 ;
        RECT 58.980 132.600 59.330 133.200 ;
        RECT 58.980 132.400 62.930 132.600 ;
        RECT 58.980 131.800 59.330 132.400 ;
        RECT 58.980 131.600 62.930 131.800 ;
        RECT 58.980 131.000 59.330 131.600 ;
        RECT 58.980 130.800 62.930 131.000 ;
        RECT 58.980 130.400 59.330 130.800 ;
        RECT 55.780 122.000 55.980 129.600 ;
        RECT 56.580 122.000 56.780 129.600 ;
        RECT 57.380 122.000 57.580 129.600 ;
        RECT 58.180 122.000 58.380 129.600 ;
        RECT 58.980 129.200 59.330 129.600 ;
        RECT 58.980 129.000 62.930 129.200 ;
        RECT 58.980 128.400 59.330 129.000 ;
        RECT 58.980 128.200 62.930 128.400 ;
        RECT 58.980 127.600 59.330 128.200 ;
        RECT 58.980 127.400 62.930 127.600 ;
        RECT 58.980 126.800 59.330 127.400 ;
        RECT 58.980 126.600 62.930 126.800 ;
        RECT 63.930 126.750 64.330 133.250 ;
        RECT 65.130 126.750 65.530 133.250 ;
        RECT 66.530 133.200 70.480 133.400 ;
        RECT 70.130 132.600 70.480 133.200 ;
        RECT 66.530 132.400 70.480 132.600 ;
        RECT 70.130 131.800 70.480 132.400 ;
        RECT 66.530 131.600 70.480 131.800 ;
        RECT 70.130 131.000 70.480 131.600 ;
        RECT 66.530 130.800 70.480 131.000 ;
        RECT 70.130 130.400 70.480 130.800 ;
        RECT 71.080 130.400 71.280 138.000 ;
        RECT 71.880 130.400 72.080 138.000 ;
        RECT 72.680 130.400 72.880 138.000 ;
        RECT 73.480 130.400 73.680 138.000 ;
        RECT 70.130 129.200 70.480 129.600 ;
        RECT 66.530 129.000 70.480 129.200 ;
        RECT 70.130 128.400 70.480 129.000 ;
        RECT 66.530 128.200 70.480 128.400 ;
        RECT 70.130 127.600 70.480 128.200 ;
        RECT 66.530 127.400 70.480 127.600 ;
        RECT 70.130 126.800 70.480 127.400 ;
        RECT 58.980 126.000 59.330 126.600 ;
        RECT 58.980 125.800 62.930 126.000 ;
        RECT 58.980 125.200 59.330 125.800 ;
        RECT 58.980 125.000 62.930 125.200 ;
        RECT 58.980 124.400 59.330 125.000 ;
        RECT 63.880 124.450 65.580 126.750 ;
        RECT 66.530 126.600 70.480 126.800 ;
        RECT 70.130 126.000 70.480 126.600 ;
        RECT 66.530 125.800 70.480 126.000 ;
        RECT 70.130 125.200 70.480 125.800 ;
        RECT 66.530 125.000 70.480 125.200 ;
        RECT 58.980 124.200 62.930 124.400 ;
        RECT 58.980 123.600 59.330 124.200 ;
        RECT 58.980 123.400 62.930 123.600 ;
        RECT 58.980 122.800 59.330 123.400 ;
        RECT 58.980 122.600 62.930 122.800 ;
        RECT 58.980 122.000 59.330 122.600 ;
        RECT 46.530 121.400 62.930 122.000 ;
        RECT 49.180 120.800 51.480 120.850 ;
        RECT 57.980 120.800 60.280 120.850 ;
        RECT 63.930 120.800 64.330 124.450 ;
        RECT 45.130 120.400 64.330 120.800 ;
        RECT 65.130 120.800 65.530 124.450 ;
        RECT 70.130 124.400 70.480 125.000 ;
        RECT 66.530 124.200 70.480 124.400 ;
        RECT 70.130 123.600 70.480 124.200 ;
        RECT 66.530 123.400 70.480 123.600 ;
        RECT 70.130 122.800 70.480 123.400 ;
        RECT 66.530 122.600 70.480 122.800 ;
        RECT 70.130 122.000 70.480 122.600 ;
        RECT 71.080 122.000 71.280 129.600 ;
        RECT 71.880 122.000 72.080 129.600 ;
        RECT 72.680 122.000 72.880 129.600 ;
        RECT 73.480 122.000 73.680 129.600 ;
        RECT 74.280 122.000 75.180 138.000 ;
        RECT 75.780 130.400 75.980 138.000 ;
        RECT 76.580 130.400 76.780 138.000 ;
        RECT 77.380 130.400 77.580 138.000 ;
        RECT 78.180 130.400 78.380 138.000 ;
        RECT 78.980 137.400 79.330 138.000 ;
        RECT 78.980 137.200 82.930 137.400 ;
        RECT 78.980 136.600 79.330 137.200 ;
        RECT 78.980 136.400 82.930 136.600 ;
        RECT 78.980 135.800 79.330 136.400 ;
        RECT 78.980 135.600 82.930 135.800 ;
        RECT 78.980 135.000 79.330 135.600 ;
        RECT 83.930 135.550 84.330 139.200 ;
        RECT 85.130 139.200 104.330 139.600 ;
        RECT 85.130 135.550 85.530 139.200 ;
        RECT 89.180 139.150 91.480 139.200 ;
        RECT 97.980 139.150 100.280 139.200 ;
        RECT 86.530 138.000 102.930 138.600 ;
        RECT 90.130 137.400 90.480 138.000 ;
        RECT 86.530 137.200 90.480 137.400 ;
        RECT 90.130 136.600 90.480 137.200 ;
        RECT 86.530 136.400 90.480 136.600 ;
        RECT 90.130 135.800 90.480 136.400 ;
        RECT 86.530 135.600 90.480 135.800 ;
        RECT 78.980 134.800 82.930 135.000 ;
        RECT 78.980 134.200 79.330 134.800 ;
        RECT 78.980 134.000 82.930 134.200 ;
        RECT 78.980 133.400 79.330 134.000 ;
        RECT 78.980 133.200 82.930 133.400 ;
        RECT 83.880 133.250 85.580 135.550 ;
        RECT 90.130 135.000 90.480 135.600 ;
        RECT 86.530 134.800 90.480 135.000 ;
        RECT 90.130 134.200 90.480 134.800 ;
        RECT 86.530 134.000 90.480 134.200 ;
        RECT 90.130 133.400 90.480 134.000 ;
        RECT 78.980 132.600 79.330 133.200 ;
        RECT 78.980 132.400 82.930 132.600 ;
        RECT 78.980 131.800 79.330 132.400 ;
        RECT 78.980 131.600 82.930 131.800 ;
        RECT 78.980 131.000 79.330 131.600 ;
        RECT 78.980 130.800 82.930 131.000 ;
        RECT 78.980 130.400 79.330 130.800 ;
        RECT 75.780 122.000 75.980 129.600 ;
        RECT 76.580 122.000 76.780 129.600 ;
        RECT 77.380 122.000 77.580 129.600 ;
        RECT 78.180 122.000 78.380 129.600 ;
        RECT 78.980 129.200 79.330 129.600 ;
        RECT 78.980 129.000 82.930 129.200 ;
        RECT 78.980 128.400 79.330 129.000 ;
        RECT 78.980 128.200 82.930 128.400 ;
        RECT 78.980 127.600 79.330 128.200 ;
        RECT 78.980 127.400 82.930 127.600 ;
        RECT 78.980 126.800 79.330 127.400 ;
        RECT 78.980 126.600 82.930 126.800 ;
        RECT 83.930 126.750 84.330 133.250 ;
        RECT 85.130 126.750 85.530 133.250 ;
        RECT 86.530 133.200 90.480 133.400 ;
        RECT 90.130 132.600 90.480 133.200 ;
        RECT 86.530 132.400 90.480 132.600 ;
        RECT 90.130 131.800 90.480 132.400 ;
        RECT 86.530 131.600 90.480 131.800 ;
        RECT 90.130 131.000 90.480 131.600 ;
        RECT 86.530 130.800 90.480 131.000 ;
        RECT 90.130 130.400 90.480 130.800 ;
        RECT 91.080 130.400 91.280 138.000 ;
        RECT 91.880 130.400 92.080 138.000 ;
        RECT 92.680 130.400 92.880 138.000 ;
        RECT 93.480 130.400 93.680 138.000 ;
        RECT 90.130 129.200 90.480 129.600 ;
        RECT 86.530 129.000 90.480 129.200 ;
        RECT 90.130 128.400 90.480 129.000 ;
        RECT 86.530 128.200 90.480 128.400 ;
        RECT 90.130 127.600 90.480 128.200 ;
        RECT 86.530 127.400 90.480 127.600 ;
        RECT 90.130 126.800 90.480 127.400 ;
        RECT 78.980 126.000 79.330 126.600 ;
        RECT 78.980 125.800 82.930 126.000 ;
        RECT 78.980 125.200 79.330 125.800 ;
        RECT 78.980 125.000 82.930 125.200 ;
        RECT 78.980 124.400 79.330 125.000 ;
        RECT 83.880 124.450 85.580 126.750 ;
        RECT 86.530 126.600 90.480 126.800 ;
        RECT 90.130 126.000 90.480 126.600 ;
        RECT 86.530 125.800 90.480 126.000 ;
        RECT 90.130 125.200 90.480 125.800 ;
        RECT 86.530 125.000 90.480 125.200 ;
        RECT 78.980 124.200 82.930 124.400 ;
        RECT 78.980 123.600 79.330 124.200 ;
        RECT 78.980 123.400 82.930 123.600 ;
        RECT 78.980 122.800 79.330 123.400 ;
        RECT 78.980 122.600 82.930 122.800 ;
        RECT 78.980 122.000 79.330 122.600 ;
        RECT 66.530 121.400 82.930 122.000 ;
        RECT 69.180 120.800 71.480 120.850 ;
        RECT 77.980 120.800 80.280 120.850 ;
        RECT 83.930 120.800 84.330 124.450 ;
        RECT 65.130 120.400 84.330 120.800 ;
        RECT 85.130 120.800 85.530 124.450 ;
        RECT 90.130 124.400 90.480 125.000 ;
        RECT 86.530 124.200 90.480 124.400 ;
        RECT 90.130 123.600 90.480 124.200 ;
        RECT 86.530 123.400 90.480 123.600 ;
        RECT 90.130 122.800 90.480 123.400 ;
        RECT 86.530 122.600 90.480 122.800 ;
        RECT 90.130 122.000 90.480 122.600 ;
        RECT 91.080 122.000 91.280 129.600 ;
        RECT 91.880 122.000 92.080 129.600 ;
        RECT 92.680 122.000 92.880 129.600 ;
        RECT 93.480 122.000 93.680 129.600 ;
        RECT 94.280 122.000 95.180 138.000 ;
        RECT 95.780 130.400 95.980 138.000 ;
        RECT 96.580 130.400 96.780 138.000 ;
        RECT 97.380 130.400 97.580 138.000 ;
        RECT 98.180 130.400 98.380 138.000 ;
        RECT 98.980 137.400 99.330 138.000 ;
        RECT 98.980 137.200 102.930 137.400 ;
        RECT 98.980 136.600 99.330 137.200 ;
        RECT 98.980 136.400 102.930 136.600 ;
        RECT 98.980 135.800 99.330 136.400 ;
        RECT 98.980 135.600 102.930 135.800 ;
        RECT 98.980 135.000 99.330 135.600 ;
        RECT 103.930 135.550 104.330 139.200 ;
        RECT 105.340 136.830 105.700 137.210 ;
        RECT 105.970 136.830 106.330 137.210 ;
        RECT 106.570 136.830 106.930 137.210 ;
        RECT 105.340 136.240 105.700 136.620 ;
        RECT 105.970 136.240 106.330 136.620 ;
        RECT 106.570 136.240 106.930 136.620 ;
        RECT 98.980 134.800 102.930 135.000 ;
        RECT 98.980 134.200 99.330 134.800 ;
        RECT 98.980 134.000 102.930 134.200 ;
        RECT 98.980 133.400 99.330 134.000 ;
        RECT 98.980 133.200 102.930 133.400 ;
        RECT 103.880 133.250 104.730 135.550 ;
        RECT 98.980 132.600 99.330 133.200 ;
        RECT 98.980 132.400 102.930 132.600 ;
        RECT 98.980 131.800 99.330 132.400 ;
        RECT 98.980 131.600 102.930 131.800 ;
        RECT 98.980 131.000 99.330 131.600 ;
        RECT 98.980 130.800 102.930 131.000 ;
        RECT 98.980 130.400 99.330 130.800 ;
        RECT 95.780 122.000 95.980 129.600 ;
        RECT 96.580 122.000 96.780 129.600 ;
        RECT 97.380 122.000 97.580 129.600 ;
        RECT 98.180 122.000 98.380 129.600 ;
        RECT 98.980 129.200 99.330 129.600 ;
        RECT 98.980 129.000 102.930 129.200 ;
        RECT 98.980 128.400 99.330 129.000 ;
        RECT 98.980 128.200 102.930 128.400 ;
        RECT 98.980 127.600 99.330 128.200 ;
        RECT 98.980 127.400 102.930 127.600 ;
        RECT 98.980 126.800 99.330 127.400 ;
        RECT 98.980 126.600 102.930 126.800 ;
        RECT 103.930 126.750 104.330 133.250 ;
        RECT 98.980 126.000 99.330 126.600 ;
        RECT 98.980 125.800 102.930 126.000 ;
        RECT 98.980 125.200 99.330 125.800 ;
        RECT 98.980 125.000 102.930 125.200 ;
        RECT 98.980 124.400 99.330 125.000 ;
        RECT 103.880 124.450 104.730 126.750 ;
        RECT 98.980 124.200 102.930 124.400 ;
        RECT 98.980 123.600 99.330 124.200 ;
        RECT 98.980 123.400 102.930 123.600 ;
        RECT 98.980 122.800 99.330 123.400 ;
        RECT 98.980 122.600 102.930 122.800 ;
        RECT 98.980 122.000 99.330 122.600 ;
        RECT 86.530 121.400 102.930 122.000 ;
        RECT 89.180 120.800 91.480 120.850 ;
        RECT 97.980 120.800 100.280 120.850 ;
        RECT 103.930 120.800 104.330 124.450 ;
        RECT 105.340 122.615 105.700 122.995 ;
        RECT 105.970 122.615 106.330 122.995 ;
        RECT 106.570 122.615 106.930 122.995 ;
        RECT 105.340 122.025 105.700 122.405 ;
        RECT 105.970 122.025 106.330 122.405 ;
        RECT 106.570 122.025 106.930 122.405 ;
        RECT 85.130 120.400 104.330 120.800 ;
        RECT 9.180 119.600 11.480 120.400 ;
        RECT 17.980 119.600 20.280 120.400 ;
        RECT 29.180 119.600 31.480 120.400 ;
        RECT 37.980 119.600 40.280 120.400 ;
        RECT 49.180 119.600 51.480 120.400 ;
        RECT 57.980 119.600 60.280 120.400 ;
        RECT 69.180 119.600 71.480 120.400 ;
        RECT 77.980 119.600 80.280 120.400 ;
        RECT 89.180 119.600 91.480 120.400 ;
        RECT 97.980 119.600 100.280 120.400 ;
        RECT 5.130 119.200 24.330 119.600 ;
        RECT 2.515 117.340 2.875 117.720 ;
        RECT 3.145 117.340 3.505 117.720 ;
        RECT 3.745 117.340 4.105 117.720 ;
        RECT 2.515 116.750 2.875 117.130 ;
        RECT 3.145 116.750 3.505 117.130 ;
        RECT 3.745 116.750 4.105 117.130 ;
        RECT 5.130 115.550 5.530 119.200 ;
        RECT 9.180 119.150 11.480 119.200 ;
        RECT 17.980 119.150 20.280 119.200 ;
        RECT 6.530 118.000 22.930 118.600 ;
        RECT 10.130 117.400 10.480 118.000 ;
        RECT 6.530 117.200 10.480 117.400 ;
        RECT 10.130 116.600 10.480 117.200 ;
        RECT 6.530 116.400 10.480 116.600 ;
        RECT 10.130 115.800 10.480 116.400 ;
        RECT 6.530 115.600 10.480 115.800 ;
        RECT 4.730 115.545 5.580 115.550 ;
        RECT 2.315 113.250 5.580 115.545 ;
        RECT 10.130 115.000 10.480 115.600 ;
        RECT 6.530 114.800 10.480 115.000 ;
        RECT 10.130 114.200 10.480 114.800 ;
        RECT 6.530 114.000 10.480 114.200 ;
        RECT 10.130 113.400 10.480 114.000 ;
        RECT 5.130 106.750 5.530 113.250 ;
        RECT 6.530 113.200 10.480 113.400 ;
        RECT 10.130 112.600 10.480 113.200 ;
        RECT 6.530 112.400 10.480 112.600 ;
        RECT 10.130 111.800 10.480 112.400 ;
        RECT 6.530 111.600 10.480 111.800 ;
        RECT 10.130 111.000 10.480 111.600 ;
        RECT 6.530 110.800 10.480 111.000 ;
        RECT 10.130 110.400 10.480 110.800 ;
        RECT 11.080 110.400 11.280 118.000 ;
        RECT 11.880 110.400 12.080 118.000 ;
        RECT 12.680 110.400 12.880 118.000 ;
        RECT 13.480 110.400 13.680 118.000 ;
        RECT 10.130 109.200 10.480 109.600 ;
        RECT 6.530 109.000 10.480 109.200 ;
        RECT 10.130 108.400 10.480 109.000 ;
        RECT 6.530 108.200 10.480 108.400 ;
        RECT 10.130 107.600 10.480 108.200 ;
        RECT 6.530 107.400 10.480 107.600 ;
        RECT 10.130 106.800 10.480 107.400 ;
        RECT 2.315 104.455 5.580 106.750 ;
        RECT 6.530 106.600 10.480 106.800 ;
        RECT 10.130 106.000 10.480 106.600 ;
        RECT 6.530 105.800 10.480 106.000 ;
        RECT 10.130 105.200 10.480 105.800 ;
        RECT 6.530 105.000 10.480 105.200 ;
        RECT 4.730 104.450 5.580 104.455 ;
        RECT 2.515 102.965 2.875 103.345 ;
        RECT 3.145 102.965 3.505 103.345 ;
        RECT 3.745 102.965 4.105 103.345 ;
        RECT 2.515 102.375 2.875 102.755 ;
        RECT 3.145 102.375 3.505 102.755 ;
        RECT 3.745 102.375 4.105 102.755 ;
        RECT 5.130 100.800 5.530 104.450 ;
        RECT 10.130 104.400 10.480 105.000 ;
        RECT 6.530 104.200 10.480 104.400 ;
        RECT 10.130 103.600 10.480 104.200 ;
        RECT 6.530 103.400 10.480 103.600 ;
        RECT 10.130 102.800 10.480 103.400 ;
        RECT 6.530 102.600 10.480 102.800 ;
        RECT 10.130 102.000 10.480 102.600 ;
        RECT 11.080 102.000 11.280 109.600 ;
        RECT 11.880 102.000 12.080 109.600 ;
        RECT 12.680 102.000 12.880 109.600 ;
        RECT 13.480 102.000 13.680 109.600 ;
        RECT 14.280 102.000 15.180 118.000 ;
        RECT 15.780 110.400 15.980 118.000 ;
        RECT 16.580 110.400 16.780 118.000 ;
        RECT 17.380 110.400 17.580 118.000 ;
        RECT 18.180 110.400 18.380 118.000 ;
        RECT 18.980 117.400 19.330 118.000 ;
        RECT 18.980 117.200 22.930 117.400 ;
        RECT 18.980 116.600 19.330 117.200 ;
        RECT 18.980 116.400 22.930 116.600 ;
        RECT 18.980 115.800 19.330 116.400 ;
        RECT 18.980 115.600 22.930 115.800 ;
        RECT 18.980 115.000 19.330 115.600 ;
        RECT 23.930 115.550 24.330 119.200 ;
        RECT 25.130 119.200 44.330 119.600 ;
        RECT 25.130 115.550 25.530 119.200 ;
        RECT 29.180 119.150 31.480 119.200 ;
        RECT 37.980 119.150 40.280 119.200 ;
        RECT 26.530 118.000 42.930 118.600 ;
        RECT 30.130 117.400 30.480 118.000 ;
        RECT 26.530 117.200 30.480 117.400 ;
        RECT 30.130 116.600 30.480 117.200 ;
        RECT 26.530 116.400 30.480 116.600 ;
        RECT 30.130 115.800 30.480 116.400 ;
        RECT 26.530 115.600 30.480 115.800 ;
        RECT 18.980 114.800 22.930 115.000 ;
        RECT 18.980 114.200 19.330 114.800 ;
        RECT 18.980 114.000 22.930 114.200 ;
        RECT 18.980 113.400 19.330 114.000 ;
        RECT 18.980 113.200 22.930 113.400 ;
        RECT 23.880 113.250 25.580 115.550 ;
        RECT 30.130 115.000 30.480 115.600 ;
        RECT 26.530 114.800 30.480 115.000 ;
        RECT 30.130 114.200 30.480 114.800 ;
        RECT 26.530 114.000 30.480 114.200 ;
        RECT 30.130 113.400 30.480 114.000 ;
        RECT 18.980 112.600 19.330 113.200 ;
        RECT 18.980 112.400 22.930 112.600 ;
        RECT 18.980 111.800 19.330 112.400 ;
        RECT 18.980 111.600 22.930 111.800 ;
        RECT 18.980 111.000 19.330 111.600 ;
        RECT 18.980 110.800 22.930 111.000 ;
        RECT 18.980 110.400 19.330 110.800 ;
        RECT 15.780 102.000 15.980 109.600 ;
        RECT 16.580 102.000 16.780 109.600 ;
        RECT 17.380 102.000 17.580 109.600 ;
        RECT 18.180 102.000 18.380 109.600 ;
        RECT 18.980 109.200 19.330 109.600 ;
        RECT 18.980 109.000 22.930 109.200 ;
        RECT 18.980 108.400 19.330 109.000 ;
        RECT 18.980 108.200 22.930 108.400 ;
        RECT 18.980 107.600 19.330 108.200 ;
        RECT 18.980 107.400 22.930 107.600 ;
        RECT 18.980 106.800 19.330 107.400 ;
        RECT 18.980 106.600 22.930 106.800 ;
        RECT 23.930 106.750 24.330 113.250 ;
        RECT 25.130 106.750 25.530 113.250 ;
        RECT 26.530 113.200 30.480 113.400 ;
        RECT 30.130 112.600 30.480 113.200 ;
        RECT 26.530 112.400 30.480 112.600 ;
        RECT 30.130 111.800 30.480 112.400 ;
        RECT 26.530 111.600 30.480 111.800 ;
        RECT 30.130 111.000 30.480 111.600 ;
        RECT 26.530 110.800 30.480 111.000 ;
        RECT 30.130 110.400 30.480 110.800 ;
        RECT 31.080 110.400 31.280 118.000 ;
        RECT 31.880 110.400 32.080 118.000 ;
        RECT 32.680 110.400 32.880 118.000 ;
        RECT 33.480 110.400 33.680 118.000 ;
        RECT 30.130 109.200 30.480 109.600 ;
        RECT 26.530 109.000 30.480 109.200 ;
        RECT 30.130 108.400 30.480 109.000 ;
        RECT 26.530 108.200 30.480 108.400 ;
        RECT 30.130 107.600 30.480 108.200 ;
        RECT 26.530 107.400 30.480 107.600 ;
        RECT 30.130 106.800 30.480 107.400 ;
        RECT 18.980 106.000 19.330 106.600 ;
        RECT 18.980 105.800 22.930 106.000 ;
        RECT 18.980 105.200 19.330 105.800 ;
        RECT 18.980 105.000 22.930 105.200 ;
        RECT 18.980 104.400 19.330 105.000 ;
        RECT 23.880 104.450 25.580 106.750 ;
        RECT 26.530 106.600 30.480 106.800 ;
        RECT 30.130 106.000 30.480 106.600 ;
        RECT 26.530 105.800 30.480 106.000 ;
        RECT 30.130 105.200 30.480 105.800 ;
        RECT 26.530 105.000 30.480 105.200 ;
        RECT 18.980 104.200 22.930 104.400 ;
        RECT 18.980 103.600 19.330 104.200 ;
        RECT 18.980 103.400 22.930 103.600 ;
        RECT 18.980 102.800 19.330 103.400 ;
        RECT 18.980 102.600 22.930 102.800 ;
        RECT 18.980 102.000 19.330 102.600 ;
        RECT 6.530 101.400 22.930 102.000 ;
        RECT 9.180 100.800 11.480 100.850 ;
        RECT 17.980 100.800 20.280 100.850 ;
        RECT 23.930 100.800 24.330 104.450 ;
        RECT 5.130 100.400 24.330 100.800 ;
        RECT 25.130 100.800 25.530 104.450 ;
        RECT 30.130 104.400 30.480 105.000 ;
        RECT 26.530 104.200 30.480 104.400 ;
        RECT 30.130 103.600 30.480 104.200 ;
        RECT 26.530 103.400 30.480 103.600 ;
        RECT 30.130 102.800 30.480 103.400 ;
        RECT 26.530 102.600 30.480 102.800 ;
        RECT 30.130 102.000 30.480 102.600 ;
        RECT 31.080 102.000 31.280 109.600 ;
        RECT 31.880 102.000 32.080 109.600 ;
        RECT 32.680 102.000 32.880 109.600 ;
        RECT 33.480 102.000 33.680 109.600 ;
        RECT 34.280 102.000 35.180 118.000 ;
        RECT 35.780 110.400 35.980 118.000 ;
        RECT 36.580 110.400 36.780 118.000 ;
        RECT 37.380 110.400 37.580 118.000 ;
        RECT 38.180 110.400 38.380 118.000 ;
        RECT 38.980 117.400 39.330 118.000 ;
        RECT 38.980 117.200 42.930 117.400 ;
        RECT 38.980 116.600 39.330 117.200 ;
        RECT 38.980 116.400 42.930 116.600 ;
        RECT 38.980 115.800 39.330 116.400 ;
        RECT 38.980 115.600 42.930 115.800 ;
        RECT 38.980 115.000 39.330 115.600 ;
        RECT 43.930 115.550 44.330 119.200 ;
        RECT 45.130 119.200 64.330 119.600 ;
        RECT 45.130 115.550 45.530 119.200 ;
        RECT 49.180 119.150 51.480 119.200 ;
        RECT 57.980 119.150 60.280 119.200 ;
        RECT 46.530 118.000 62.930 118.600 ;
        RECT 50.130 117.400 50.480 118.000 ;
        RECT 46.530 117.200 50.480 117.400 ;
        RECT 50.130 116.600 50.480 117.200 ;
        RECT 46.530 116.400 50.480 116.600 ;
        RECT 50.130 115.800 50.480 116.400 ;
        RECT 46.530 115.600 50.480 115.800 ;
        RECT 38.980 114.800 42.930 115.000 ;
        RECT 38.980 114.200 39.330 114.800 ;
        RECT 38.980 114.000 42.930 114.200 ;
        RECT 38.980 113.400 39.330 114.000 ;
        RECT 38.980 113.200 42.930 113.400 ;
        RECT 43.880 113.250 45.580 115.550 ;
        RECT 50.130 115.000 50.480 115.600 ;
        RECT 46.530 114.800 50.480 115.000 ;
        RECT 50.130 114.200 50.480 114.800 ;
        RECT 46.530 114.000 50.480 114.200 ;
        RECT 50.130 113.400 50.480 114.000 ;
        RECT 38.980 112.600 39.330 113.200 ;
        RECT 38.980 112.400 42.930 112.600 ;
        RECT 38.980 111.800 39.330 112.400 ;
        RECT 38.980 111.600 42.930 111.800 ;
        RECT 38.980 111.000 39.330 111.600 ;
        RECT 38.980 110.800 42.930 111.000 ;
        RECT 38.980 110.400 39.330 110.800 ;
        RECT 35.780 102.000 35.980 109.600 ;
        RECT 36.580 102.000 36.780 109.600 ;
        RECT 37.380 102.000 37.580 109.600 ;
        RECT 38.180 102.000 38.380 109.600 ;
        RECT 38.980 109.200 39.330 109.600 ;
        RECT 38.980 109.000 42.930 109.200 ;
        RECT 38.980 108.400 39.330 109.000 ;
        RECT 38.980 108.200 42.930 108.400 ;
        RECT 38.980 107.600 39.330 108.200 ;
        RECT 38.980 107.400 42.930 107.600 ;
        RECT 38.980 106.800 39.330 107.400 ;
        RECT 38.980 106.600 42.930 106.800 ;
        RECT 43.930 106.750 44.330 113.250 ;
        RECT 45.130 106.750 45.530 113.250 ;
        RECT 46.530 113.200 50.480 113.400 ;
        RECT 50.130 112.600 50.480 113.200 ;
        RECT 46.530 112.400 50.480 112.600 ;
        RECT 50.130 111.800 50.480 112.400 ;
        RECT 46.530 111.600 50.480 111.800 ;
        RECT 50.130 111.000 50.480 111.600 ;
        RECT 46.530 110.800 50.480 111.000 ;
        RECT 50.130 110.400 50.480 110.800 ;
        RECT 51.080 110.400 51.280 118.000 ;
        RECT 51.880 110.400 52.080 118.000 ;
        RECT 52.680 110.400 52.880 118.000 ;
        RECT 53.480 110.400 53.680 118.000 ;
        RECT 50.130 109.200 50.480 109.600 ;
        RECT 46.530 109.000 50.480 109.200 ;
        RECT 50.130 108.400 50.480 109.000 ;
        RECT 46.530 108.200 50.480 108.400 ;
        RECT 50.130 107.600 50.480 108.200 ;
        RECT 46.530 107.400 50.480 107.600 ;
        RECT 50.130 106.800 50.480 107.400 ;
        RECT 38.980 106.000 39.330 106.600 ;
        RECT 38.980 105.800 42.930 106.000 ;
        RECT 38.980 105.200 39.330 105.800 ;
        RECT 38.980 105.000 42.930 105.200 ;
        RECT 38.980 104.400 39.330 105.000 ;
        RECT 43.880 104.450 45.580 106.750 ;
        RECT 46.530 106.600 50.480 106.800 ;
        RECT 50.130 106.000 50.480 106.600 ;
        RECT 46.530 105.800 50.480 106.000 ;
        RECT 50.130 105.200 50.480 105.800 ;
        RECT 46.530 105.000 50.480 105.200 ;
        RECT 38.980 104.200 42.930 104.400 ;
        RECT 38.980 103.600 39.330 104.200 ;
        RECT 38.980 103.400 42.930 103.600 ;
        RECT 38.980 102.800 39.330 103.400 ;
        RECT 38.980 102.600 42.930 102.800 ;
        RECT 38.980 102.000 39.330 102.600 ;
        RECT 26.530 101.400 42.930 102.000 ;
        RECT 29.180 100.800 31.480 100.850 ;
        RECT 37.980 100.800 40.280 100.850 ;
        RECT 43.930 100.800 44.330 104.450 ;
        RECT 25.130 100.400 44.330 100.800 ;
        RECT 45.130 100.800 45.530 104.450 ;
        RECT 50.130 104.400 50.480 105.000 ;
        RECT 46.530 104.200 50.480 104.400 ;
        RECT 50.130 103.600 50.480 104.200 ;
        RECT 46.530 103.400 50.480 103.600 ;
        RECT 50.130 102.800 50.480 103.400 ;
        RECT 46.530 102.600 50.480 102.800 ;
        RECT 50.130 102.000 50.480 102.600 ;
        RECT 51.080 102.000 51.280 109.600 ;
        RECT 51.880 102.000 52.080 109.600 ;
        RECT 52.680 102.000 52.880 109.600 ;
        RECT 53.480 102.000 53.680 109.600 ;
        RECT 54.280 102.000 55.180 118.000 ;
        RECT 55.780 110.400 55.980 118.000 ;
        RECT 56.580 110.400 56.780 118.000 ;
        RECT 57.380 110.400 57.580 118.000 ;
        RECT 58.180 110.400 58.380 118.000 ;
        RECT 58.980 117.400 59.330 118.000 ;
        RECT 58.980 117.200 62.930 117.400 ;
        RECT 58.980 116.600 59.330 117.200 ;
        RECT 58.980 116.400 62.930 116.600 ;
        RECT 58.980 115.800 59.330 116.400 ;
        RECT 58.980 115.600 62.930 115.800 ;
        RECT 58.980 115.000 59.330 115.600 ;
        RECT 63.930 115.550 64.330 119.200 ;
        RECT 65.130 119.200 84.330 119.600 ;
        RECT 65.130 115.550 65.530 119.200 ;
        RECT 69.180 119.150 71.480 119.200 ;
        RECT 77.980 119.150 80.280 119.200 ;
        RECT 66.530 118.000 82.930 118.600 ;
        RECT 70.130 117.400 70.480 118.000 ;
        RECT 66.530 117.200 70.480 117.400 ;
        RECT 70.130 116.600 70.480 117.200 ;
        RECT 66.530 116.400 70.480 116.600 ;
        RECT 70.130 115.800 70.480 116.400 ;
        RECT 66.530 115.600 70.480 115.800 ;
        RECT 58.980 114.800 62.930 115.000 ;
        RECT 58.980 114.200 59.330 114.800 ;
        RECT 58.980 114.000 62.930 114.200 ;
        RECT 58.980 113.400 59.330 114.000 ;
        RECT 58.980 113.200 62.930 113.400 ;
        RECT 63.880 113.250 65.580 115.550 ;
        RECT 70.130 115.000 70.480 115.600 ;
        RECT 66.530 114.800 70.480 115.000 ;
        RECT 70.130 114.200 70.480 114.800 ;
        RECT 66.530 114.000 70.480 114.200 ;
        RECT 70.130 113.400 70.480 114.000 ;
        RECT 58.980 112.600 59.330 113.200 ;
        RECT 58.980 112.400 62.930 112.600 ;
        RECT 58.980 111.800 59.330 112.400 ;
        RECT 58.980 111.600 62.930 111.800 ;
        RECT 58.980 111.000 59.330 111.600 ;
        RECT 58.980 110.800 62.930 111.000 ;
        RECT 58.980 110.400 59.330 110.800 ;
        RECT 55.780 102.000 55.980 109.600 ;
        RECT 56.580 102.000 56.780 109.600 ;
        RECT 57.380 102.000 57.580 109.600 ;
        RECT 58.180 102.000 58.380 109.600 ;
        RECT 58.980 109.200 59.330 109.600 ;
        RECT 58.980 109.000 62.930 109.200 ;
        RECT 58.980 108.400 59.330 109.000 ;
        RECT 58.980 108.200 62.930 108.400 ;
        RECT 58.980 107.600 59.330 108.200 ;
        RECT 58.980 107.400 62.930 107.600 ;
        RECT 58.980 106.800 59.330 107.400 ;
        RECT 58.980 106.600 62.930 106.800 ;
        RECT 63.930 106.750 64.330 113.250 ;
        RECT 65.130 106.750 65.530 113.250 ;
        RECT 66.530 113.200 70.480 113.400 ;
        RECT 70.130 112.600 70.480 113.200 ;
        RECT 66.530 112.400 70.480 112.600 ;
        RECT 70.130 111.800 70.480 112.400 ;
        RECT 66.530 111.600 70.480 111.800 ;
        RECT 70.130 111.000 70.480 111.600 ;
        RECT 66.530 110.800 70.480 111.000 ;
        RECT 70.130 110.400 70.480 110.800 ;
        RECT 71.080 110.400 71.280 118.000 ;
        RECT 71.880 110.400 72.080 118.000 ;
        RECT 72.680 110.400 72.880 118.000 ;
        RECT 73.480 110.400 73.680 118.000 ;
        RECT 70.130 109.200 70.480 109.600 ;
        RECT 66.530 109.000 70.480 109.200 ;
        RECT 70.130 108.400 70.480 109.000 ;
        RECT 66.530 108.200 70.480 108.400 ;
        RECT 70.130 107.600 70.480 108.200 ;
        RECT 66.530 107.400 70.480 107.600 ;
        RECT 70.130 106.800 70.480 107.400 ;
        RECT 58.980 106.000 59.330 106.600 ;
        RECT 58.980 105.800 62.930 106.000 ;
        RECT 58.980 105.200 59.330 105.800 ;
        RECT 58.980 105.000 62.930 105.200 ;
        RECT 58.980 104.400 59.330 105.000 ;
        RECT 63.880 104.450 65.580 106.750 ;
        RECT 66.530 106.600 70.480 106.800 ;
        RECT 70.130 106.000 70.480 106.600 ;
        RECT 66.530 105.800 70.480 106.000 ;
        RECT 70.130 105.200 70.480 105.800 ;
        RECT 66.530 105.000 70.480 105.200 ;
        RECT 58.980 104.200 62.930 104.400 ;
        RECT 58.980 103.600 59.330 104.200 ;
        RECT 58.980 103.400 62.930 103.600 ;
        RECT 58.980 102.800 59.330 103.400 ;
        RECT 58.980 102.600 62.930 102.800 ;
        RECT 58.980 102.000 59.330 102.600 ;
        RECT 46.530 101.400 62.930 102.000 ;
        RECT 49.180 100.800 51.480 100.850 ;
        RECT 57.980 100.800 60.280 100.850 ;
        RECT 63.930 100.800 64.330 104.450 ;
        RECT 45.130 100.400 64.330 100.800 ;
        RECT 65.130 100.800 65.530 104.450 ;
        RECT 70.130 104.400 70.480 105.000 ;
        RECT 66.530 104.200 70.480 104.400 ;
        RECT 70.130 103.600 70.480 104.200 ;
        RECT 66.530 103.400 70.480 103.600 ;
        RECT 70.130 102.800 70.480 103.400 ;
        RECT 66.530 102.600 70.480 102.800 ;
        RECT 70.130 102.000 70.480 102.600 ;
        RECT 71.080 102.000 71.280 109.600 ;
        RECT 71.880 102.000 72.080 109.600 ;
        RECT 72.680 102.000 72.880 109.600 ;
        RECT 73.480 102.000 73.680 109.600 ;
        RECT 74.280 102.000 75.180 118.000 ;
        RECT 75.780 110.400 75.980 118.000 ;
        RECT 76.580 110.400 76.780 118.000 ;
        RECT 77.380 110.400 77.580 118.000 ;
        RECT 78.180 110.400 78.380 118.000 ;
        RECT 78.980 117.400 79.330 118.000 ;
        RECT 78.980 117.200 82.930 117.400 ;
        RECT 78.980 116.600 79.330 117.200 ;
        RECT 78.980 116.400 82.930 116.600 ;
        RECT 78.980 115.800 79.330 116.400 ;
        RECT 78.980 115.600 82.930 115.800 ;
        RECT 78.980 115.000 79.330 115.600 ;
        RECT 83.930 115.550 84.330 119.200 ;
        RECT 85.130 119.200 104.330 119.600 ;
        RECT 85.130 115.550 85.530 119.200 ;
        RECT 89.180 119.150 91.480 119.200 ;
        RECT 97.980 119.150 100.280 119.200 ;
        RECT 86.530 118.000 102.930 118.600 ;
        RECT 90.130 117.400 90.480 118.000 ;
        RECT 86.530 117.200 90.480 117.400 ;
        RECT 90.130 116.600 90.480 117.200 ;
        RECT 86.530 116.400 90.480 116.600 ;
        RECT 90.130 115.800 90.480 116.400 ;
        RECT 86.530 115.600 90.480 115.800 ;
        RECT 78.980 114.800 82.930 115.000 ;
        RECT 78.980 114.200 79.330 114.800 ;
        RECT 78.980 114.000 82.930 114.200 ;
        RECT 78.980 113.400 79.330 114.000 ;
        RECT 78.980 113.200 82.930 113.400 ;
        RECT 83.880 113.250 85.580 115.550 ;
        RECT 90.130 115.000 90.480 115.600 ;
        RECT 86.530 114.800 90.480 115.000 ;
        RECT 90.130 114.200 90.480 114.800 ;
        RECT 86.530 114.000 90.480 114.200 ;
        RECT 90.130 113.400 90.480 114.000 ;
        RECT 78.980 112.600 79.330 113.200 ;
        RECT 78.980 112.400 82.930 112.600 ;
        RECT 78.980 111.800 79.330 112.400 ;
        RECT 78.980 111.600 82.930 111.800 ;
        RECT 78.980 111.000 79.330 111.600 ;
        RECT 78.980 110.800 82.930 111.000 ;
        RECT 78.980 110.400 79.330 110.800 ;
        RECT 75.780 102.000 75.980 109.600 ;
        RECT 76.580 102.000 76.780 109.600 ;
        RECT 77.380 102.000 77.580 109.600 ;
        RECT 78.180 102.000 78.380 109.600 ;
        RECT 78.980 109.200 79.330 109.600 ;
        RECT 78.980 109.000 82.930 109.200 ;
        RECT 78.980 108.400 79.330 109.000 ;
        RECT 78.980 108.200 82.930 108.400 ;
        RECT 78.980 107.600 79.330 108.200 ;
        RECT 78.980 107.400 82.930 107.600 ;
        RECT 78.980 106.800 79.330 107.400 ;
        RECT 78.980 106.600 82.930 106.800 ;
        RECT 83.930 106.750 84.330 113.250 ;
        RECT 85.130 106.750 85.530 113.250 ;
        RECT 86.530 113.200 90.480 113.400 ;
        RECT 90.130 112.600 90.480 113.200 ;
        RECT 86.530 112.400 90.480 112.600 ;
        RECT 90.130 111.800 90.480 112.400 ;
        RECT 86.530 111.600 90.480 111.800 ;
        RECT 90.130 111.000 90.480 111.600 ;
        RECT 86.530 110.800 90.480 111.000 ;
        RECT 90.130 110.400 90.480 110.800 ;
        RECT 91.080 110.400 91.280 118.000 ;
        RECT 91.880 110.400 92.080 118.000 ;
        RECT 92.680 110.400 92.880 118.000 ;
        RECT 93.480 110.400 93.680 118.000 ;
        RECT 90.130 109.200 90.480 109.600 ;
        RECT 86.530 109.000 90.480 109.200 ;
        RECT 90.130 108.400 90.480 109.000 ;
        RECT 86.530 108.200 90.480 108.400 ;
        RECT 90.130 107.600 90.480 108.200 ;
        RECT 86.530 107.400 90.480 107.600 ;
        RECT 90.130 106.800 90.480 107.400 ;
        RECT 78.980 106.000 79.330 106.600 ;
        RECT 78.980 105.800 82.930 106.000 ;
        RECT 78.980 105.200 79.330 105.800 ;
        RECT 78.980 105.000 82.930 105.200 ;
        RECT 78.980 104.400 79.330 105.000 ;
        RECT 83.880 104.450 85.580 106.750 ;
        RECT 86.530 106.600 90.480 106.800 ;
        RECT 90.130 106.000 90.480 106.600 ;
        RECT 86.530 105.800 90.480 106.000 ;
        RECT 90.130 105.200 90.480 105.800 ;
        RECT 86.530 105.000 90.480 105.200 ;
        RECT 78.980 104.200 82.930 104.400 ;
        RECT 78.980 103.600 79.330 104.200 ;
        RECT 78.980 103.400 82.930 103.600 ;
        RECT 78.980 102.800 79.330 103.400 ;
        RECT 78.980 102.600 82.930 102.800 ;
        RECT 78.980 102.000 79.330 102.600 ;
        RECT 66.530 101.400 82.930 102.000 ;
        RECT 69.180 100.800 71.480 100.850 ;
        RECT 77.980 100.800 80.280 100.850 ;
        RECT 83.930 100.800 84.330 104.450 ;
        RECT 65.130 100.400 84.330 100.800 ;
        RECT 85.130 100.800 85.530 104.450 ;
        RECT 90.130 104.400 90.480 105.000 ;
        RECT 86.530 104.200 90.480 104.400 ;
        RECT 90.130 103.600 90.480 104.200 ;
        RECT 86.530 103.400 90.480 103.600 ;
        RECT 90.130 102.800 90.480 103.400 ;
        RECT 86.530 102.600 90.480 102.800 ;
        RECT 90.130 102.000 90.480 102.600 ;
        RECT 91.080 102.000 91.280 109.600 ;
        RECT 91.880 102.000 92.080 109.600 ;
        RECT 92.680 102.000 92.880 109.600 ;
        RECT 93.480 102.000 93.680 109.600 ;
        RECT 94.280 102.000 95.180 118.000 ;
        RECT 95.780 110.400 95.980 118.000 ;
        RECT 96.580 110.400 96.780 118.000 ;
        RECT 97.380 110.400 97.580 118.000 ;
        RECT 98.180 110.400 98.380 118.000 ;
        RECT 98.980 117.400 99.330 118.000 ;
        RECT 98.980 117.200 102.930 117.400 ;
        RECT 98.980 116.600 99.330 117.200 ;
        RECT 98.980 116.400 102.930 116.600 ;
        RECT 98.980 115.800 99.330 116.400 ;
        RECT 98.980 115.600 102.930 115.800 ;
        RECT 98.980 115.000 99.330 115.600 ;
        RECT 103.930 115.550 104.330 119.200 ;
        RECT 105.340 116.740 105.700 117.120 ;
        RECT 105.970 116.740 106.330 117.120 ;
        RECT 106.570 116.740 106.930 117.120 ;
        RECT 105.340 116.150 105.700 116.530 ;
        RECT 105.970 116.150 106.330 116.530 ;
        RECT 106.570 116.150 106.930 116.530 ;
        RECT 98.980 114.800 102.930 115.000 ;
        RECT 98.980 114.200 99.330 114.800 ;
        RECT 98.980 114.000 102.930 114.200 ;
        RECT 98.980 113.400 99.330 114.000 ;
        RECT 98.980 113.200 102.930 113.400 ;
        RECT 103.880 113.250 104.730 115.550 ;
        RECT 98.980 112.600 99.330 113.200 ;
        RECT 98.980 112.400 102.930 112.600 ;
        RECT 98.980 111.800 99.330 112.400 ;
        RECT 98.980 111.600 102.930 111.800 ;
        RECT 98.980 111.000 99.330 111.600 ;
        RECT 98.980 110.800 102.930 111.000 ;
        RECT 98.980 110.400 99.330 110.800 ;
        RECT 95.780 102.000 95.980 109.600 ;
        RECT 96.580 102.000 96.780 109.600 ;
        RECT 97.380 102.000 97.580 109.600 ;
        RECT 98.180 102.000 98.380 109.600 ;
        RECT 98.980 109.200 99.330 109.600 ;
        RECT 98.980 109.000 102.930 109.200 ;
        RECT 98.980 108.400 99.330 109.000 ;
        RECT 98.980 108.200 102.930 108.400 ;
        RECT 98.980 107.600 99.330 108.200 ;
        RECT 98.980 107.400 102.930 107.600 ;
        RECT 98.980 106.800 99.330 107.400 ;
        RECT 98.980 106.600 102.930 106.800 ;
        RECT 103.930 106.750 104.330 113.250 ;
        RECT 98.980 106.000 99.330 106.600 ;
        RECT 98.980 105.800 102.930 106.000 ;
        RECT 98.980 105.200 99.330 105.800 ;
        RECT 98.980 105.000 102.930 105.200 ;
        RECT 98.980 104.400 99.330 105.000 ;
        RECT 103.880 104.450 104.730 106.750 ;
        RECT 98.980 104.200 102.930 104.400 ;
        RECT 98.980 103.600 99.330 104.200 ;
        RECT 98.980 103.400 102.930 103.600 ;
        RECT 98.980 102.800 99.330 103.400 ;
        RECT 98.980 102.600 102.930 102.800 ;
        RECT 98.980 102.000 99.330 102.600 ;
        RECT 86.530 101.400 102.930 102.000 ;
        RECT 89.180 100.800 91.480 100.850 ;
        RECT 97.980 100.800 100.280 100.850 ;
        RECT 103.930 100.800 104.330 104.450 ;
        RECT 105.340 102.535 105.700 102.915 ;
        RECT 105.970 102.535 106.330 102.915 ;
        RECT 106.570 102.535 106.930 102.915 ;
        RECT 105.340 101.945 105.700 102.325 ;
        RECT 105.970 101.945 106.330 102.325 ;
        RECT 106.570 101.945 106.930 102.325 ;
        RECT 85.130 100.400 104.330 100.800 ;
        RECT 9.180 99.600 11.480 100.400 ;
        RECT 17.980 99.600 20.280 100.400 ;
        RECT 29.180 99.600 31.480 100.400 ;
        RECT 37.980 99.600 40.280 100.400 ;
        RECT 49.180 99.600 51.480 100.400 ;
        RECT 57.980 99.600 60.280 100.400 ;
        RECT 69.180 99.600 71.480 100.400 ;
        RECT 77.980 99.600 80.280 100.400 ;
        RECT 89.180 99.600 91.480 100.400 ;
        RECT 97.980 99.600 100.280 100.400 ;
        RECT 5.130 99.200 24.330 99.600 ;
        RECT 2.515 97.460 2.875 97.840 ;
        RECT 3.145 97.460 3.505 97.840 ;
        RECT 3.745 97.460 4.105 97.840 ;
        RECT 2.515 96.870 2.875 97.250 ;
        RECT 3.145 96.870 3.505 97.250 ;
        RECT 3.745 96.870 4.105 97.250 ;
        RECT 5.130 95.550 5.530 99.200 ;
        RECT 9.180 99.150 11.480 99.200 ;
        RECT 17.980 99.150 20.280 99.200 ;
        RECT 6.530 98.000 22.930 98.600 ;
        RECT 10.130 97.400 10.480 98.000 ;
        RECT 6.530 97.200 10.480 97.400 ;
        RECT 10.130 96.600 10.480 97.200 ;
        RECT 6.530 96.400 10.480 96.600 ;
        RECT 10.130 95.800 10.480 96.400 ;
        RECT 6.530 95.600 10.480 95.800 ;
        RECT 4.730 95.545 5.580 95.550 ;
        RECT 2.315 93.250 5.580 95.545 ;
        RECT 10.130 95.000 10.480 95.600 ;
        RECT 6.530 94.800 10.480 95.000 ;
        RECT 10.130 94.200 10.480 94.800 ;
        RECT 6.530 94.000 10.480 94.200 ;
        RECT 10.130 93.400 10.480 94.000 ;
        RECT 5.130 86.750 5.530 93.250 ;
        RECT 6.530 93.200 10.480 93.400 ;
        RECT 10.130 92.600 10.480 93.200 ;
        RECT 6.530 92.400 10.480 92.600 ;
        RECT 10.130 91.800 10.480 92.400 ;
        RECT 6.530 91.600 10.480 91.800 ;
        RECT 10.130 91.000 10.480 91.600 ;
        RECT 6.530 90.800 10.480 91.000 ;
        RECT 10.130 90.400 10.480 90.800 ;
        RECT 11.080 90.400 11.280 98.000 ;
        RECT 11.880 90.400 12.080 98.000 ;
        RECT 12.680 90.400 12.880 98.000 ;
        RECT 13.480 90.400 13.680 98.000 ;
        RECT 10.130 89.200 10.480 89.600 ;
        RECT 6.530 89.000 10.480 89.200 ;
        RECT 10.130 88.400 10.480 89.000 ;
        RECT 6.530 88.200 10.480 88.400 ;
        RECT 10.130 87.600 10.480 88.200 ;
        RECT 6.530 87.400 10.480 87.600 ;
        RECT 10.130 86.800 10.480 87.400 ;
        RECT 4.730 86.745 5.580 86.750 ;
        RECT 2.315 84.450 5.580 86.745 ;
        RECT 6.530 86.600 10.480 86.800 ;
        RECT 10.130 86.000 10.480 86.600 ;
        RECT 6.530 85.800 10.480 86.000 ;
        RECT 10.130 85.200 10.480 85.800 ;
        RECT 6.530 85.000 10.480 85.200 ;
        RECT 2.515 83.130 2.875 83.510 ;
        RECT 3.145 83.130 3.505 83.510 ;
        RECT 3.745 83.130 4.105 83.510 ;
        RECT 2.515 82.540 2.875 82.920 ;
        RECT 3.145 82.540 3.505 82.920 ;
        RECT 3.745 82.540 4.105 82.920 ;
        RECT 5.130 80.800 5.530 84.450 ;
        RECT 10.130 84.400 10.480 85.000 ;
        RECT 6.530 84.200 10.480 84.400 ;
        RECT 10.130 83.600 10.480 84.200 ;
        RECT 6.530 83.400 10.480 83.600 ;
        RECT 10.130 82.800 10.480 83.400 ;
        RECT 6.530 82.600 10.480 82.800 ;
        RECT 10.130 82.000 10.480 82.600 ;
        RECT 11.080 82.000 11.280 89.600 ;
        RECT 11.880 82.000 12.080 89.600 ;
        RECT 12.680 82.000 12.880 89.600 ;
        RECT 13.480 82.000 13.680 89.600 ;
        RECT 14.280 82.000 15.180 98.000 ;
        RECT 15.780 90.400 15.980 98.000 ;
        RECT 16.580 90.400 16.780 98.000 ;
        RECT 17.380 90.400 17.580 98.000 ;
        RECT 18.180 90.400 18.380 98.000 ;
        RECT 18.980 97.400 19.330 98.000 ;
        RECT 18.980 97.200 22.930 97.400 ;
        RECT 18.980 96.600 19.330 97.200 ;
        RECT 18.980 96.400 22.930 96.600 ;
        RECT 18.980 95.800 19.330 96.400 ;
        RECT 18.980 95.600 22.930 95.800 ;
        RECT 18.980 95.000 19.330 95.600 ;
        RECT 23.930 95.550 24.330 99.200 ;
        RECT 25.130 99.200 44.330 99.600 ;
        RECT 25.130 95.550 25.530 99.200 ;
        RECT 29.180 99.150 31.480 99.200 ;
        RECT 37.980 99.150 40.280 99.200 ;
        RECT 26.530 98.000 42.930 98.600 ;
        RECT 30.130 97.400 30.480 98.000 ;
        RECT 26.530 97.200 30.480 97.400 ;
        RECT 30.130 96.600 30.480 97.200 ;
        RECT 26.530 96.400 30.480 96.600 ;
        RECT 30.130 95.800 30.480 96.400 ;
        RECT 26.530 95.600 30.480 95.800 ;
        RECT 18.980 94.800 22.930 95.000 ;
        RECT 18.980 94.200 19.330 94.800 ;
        RECT 18.980 94.000 22.930 94.200 ;
        RECT 18.980 93.400 19.330 94.000 ;
        RECT 18.980 93.200 22.930 93.400 ;
        RECT 23.880 93.250 25.580 95.550 ;
        RECT 30.130 95.000 30.480 95.600 ;
        RECT 26.530 94.800 30.480 95.000 ;
        RECT 30.130 94.200 30.480 94.800 ;
        RECT 26.530 94.000 30.480 94.200 ;
        RECT 30.130 93.400 30.480 94.000 ;
        RECT 18.980 92.600 19.330 93.200 ;
        RECT 18.980 92.400 22.930 92.600 ;
        RECT 18.980 91.800 19.330 92.400 ;
        RECT 18.980 91.600 22.930 91.800 ;
        RECT 18.980 91.000 19.330 91.600 ;
        RECT 18.980 90.800 22.930 91.000 ;
        RECT 18.980 90.400 19.330 90.800 ;
        RECT 15.780 82.000 15.980 89.600 ;
        RECT 16.580 82.000 16.780 89.600 ;
        RECT 17.380 82.000 17.580 89.600 ;
        RECT 18.180 82.000 18.380 89.600 ;
        RECT 18.980 89.200 19.330 89.600 ;
        RECT 18.980 89.000 22.930 89.200 ;
        RECT 18.980 88.400 19.330 89.000 ;
        RECT 18.980 88.200 22.930 88.400 ;
        RECT 18.980 87.600 19.330 88.200 ;
        RECT 18.980 87.400 22.930 87.600 ;
        RECT 18.980 86.800 19.330 87.400 ;
        RECT 18.980 86.600 22.930 86.800 ;
        RECT 23.930 86.750 24.330 93.250 ;
        RECT 25.130 86.750 25.530 93.250 ;
        RECT 26.530 93.200 30.480 93.400 ;
        RECT 30.130 92.600 30.480 93.200 ;
        RECT 26.530 92.400 30.480 92.600 ;
        RECT 30.130 91.800 30.480 92.400 ;
        RECT 26.530 91.600 30.480 91.800 ;
        RECT 30.130 91.000 30.480 91.600 ;
        RECT 26.530 90.800 30.480 91.000 ;
        RECT 30.130 90.400 30.480 90.800 ;
        RECT 31.080 90.400 31.280 98.000 ;
        RECT 31.880 90.400 32.080 98.000 ;
        RECT 32.680 90.400 32.880 98.000 ;
        RECT 33.480 90.400 33.680 98.000 ;
        RECT 30.130 89.200 30.480 89.600 ;
        RECT 26.530 89.000 30.480 89.200 ;
        RECT 30.130 88.400 30.480 89.000 ;
        RECT 26.530 88.200 30.480 88.400 ;
        RECT 30.130 87.600 30.480 88.200 ;
        RECT 26.530 87.400 30.480 87.600 ;
        RECT 30.130 86.800 30.480 87.400 ;
        RECT 18.980 86.000 19.330 86.600 ;
        RECT 18.980 85.800 22.930 86.000 ;
        RECT 18.980 85.200 19.330 85.800 ;
        RECT 18.980 85.000 22.930 85.200 ;
        RECT 18.980 84.400 19.330 85.000 ;
        RECT 23.880 84.450 25.580 86.750 ;
        RECT 26.530 86.600 30.480 86.800 ;
        RECT 30.130 86.000 30.480 86.600 ;
        RECT 26.530 85.800 30.480 86.000 ;
        RECT 30.130 85.200 30.480 85.800 ;
        RECT 26.530 85.000 30.480 85.200 ;
        RECT 18.980 84.200 22.930 84.400 ;
        RECT 18.980 83.600 19.330 84.200 ;
        RECT 18.980 83.400 22.930 83.600 ;
        RECT 18.980 82.800 19.330 83.400 ;
        RECT 18.980 82.600 22.930 82.800 ;
        RECT 18.980 82.000 19.330 82.600 ;
        RECT 6.530 81.400 22.930 82.000 ;
        RECT 9.180 80.800 11.480 80.850 ;
        RECT 17.980 80.800 20.280 80.850 ;
        RECT 23.930 80.800 24.330 84.450 ;
        RECT 5.130 80.400 24.330 80.800 ;
        RECT 25.130 80.800 25.530 84.450 ;
        RECT 30.130 84.400 30.480 85.000 ;
        RECT 26.530 84.200 30.480 84.400 ;
        RECT 30.130 83.600 30.480 84.200 ;
        RECT 26.530 83.400 30.480 83.600 ;
        RECT 30.130 82.800 30.480 83.400 ;
        RECT 26.530 82.600 30.480 82.800 ;
        RECT 30.130 82.000 30.480 82.600 ;
        RECT 31.080 82.000 31.280 89.600 ;
        RECT 31.880 82.000 32.080 89.600 ;
        RECT 32.680 82.000 32.880 89.600 ;
        RECT 33.480 82.000 33.680 89.600 ;
        RECT 34.280 82.000 35.180 98.000 ;
        RECT 35.780 90.400 35.980 98.000 ;
        RECT 36.580 90.400 36.780 98.000 ;
        RECT 37.380 90.400 37.580 98.000 ;
        RECT 38.180 90.400 38.380 98.000 ;
        RECT 38.980 97.400 39.330 98.000 ;
        RECT 38.980 97.200 42.930 97.400 ;
        RECT 38.980 96.600 39.330 97.200 ;
        RECT 38.980 96.400 42.930 96.600 ;
        RECT 38.980 95.800 39.330 96.400 ;
        RECT 38.980 95.600 42.930 95.800 ;
        RECT 38.980 95.000 39.330 95.600 ;
        RECT 43.930 95.550 44.330 99.200 ;
        RECT 45.130 99.200 64.330 99.600 ;
        RECT 45.130 95.550 45.530 99.200 ;
        RECT 49.180 99.150 51.480 99.200 ;
        RECT 57.980 99.150 60.280 99.200 ;
        RECT 46.530 98.000 62.930 98.600 ;
        RECT 50.130 97.400 50.480 98.000 ;
        RECT 46.530 97.200 50.480 97.400 ;
        RECT 50.130 96.600 50.480 97.200 ;
        RECT 46.530 96.400 50.480 96.600 ;
        RECT 50.130 95.800 50.480 96.400 ;
        RECT 46.530 95.600 50.480 95.800 ;
        RECT 38.980 94.800 42.930 95.000 ;
        RECT 38.980 94.200 39.330 94.800 ;
        RECT 38.980 94.000 42.930 94.200 ;
        RECT 38.980 93.400 39.330 94.000 ;
        RECT 38.980 93.200 42.930 93.400 ;
        RECT 43.880 93.250 45.580 95.550 ;
        RECT 50.130 95.000 50.480 95.600 ;
        RECT 46.530 94.800 50.480 95.000 ;
        RECT 50.130 94.200 50.480 94.800 ;
        RECT 46.530 94.000 50.480 94.200 ;
        RECT 50.130 93.400 50.480 94.000 ;
        RECT 38.980 92.600 39.330 93.200 ;
        RECT 38.980 92.400 42.930 92.600 ;
        RECT 38.980 91.800 39.330 92.400 ;
        RECT 38.980 91.600 42.930 91.800 ;
        RECT 38.980 91.000 39.330 91.600 ;
        RECT 38.980 90.800 42.930 91.000 ;
        RECT 38.980 90.400 39.330 90.800 ;
        RECT 35.780 82.000 35.980 89.600 ;
        RECT 36.580 82.000 36.780 89.600 ;
        RECT 37.380 82.000 37.580 89.600 ;
        RECT 38.180 82.000 38.380 89.600 ;
        RECT 38.980 89.200 39.330 89.600 ;
        RECT 38.980 89.000 42.930 89.200 ;
        RECT 38.980 88.400 39.330 89.000 ;
        RECT 38.980 88.200 42.930 88.400 ;
        RECT 38.980 87.600 39.330 88.200 ;
        RECT 38.980 87.400 42.930 87.600 ;
        RECT 38.980 86.800 39.330 87.400 ;
        RECT 38.980 86.600 42.930 86.800 ;
        RECT 43.930 86.750 44.330 93.250 ;
        RECT 45.130 86.750 45.530 93.250 ;
        RECT 46.530 93.200 50.480 93.400 ;
        RECT 50.130 92.600 50.480 93.200 ;
        RECT 46.530 92.400 50.480 92.600 ;
        RECT 50.130 91.800 50.480 92.400 ;
        RECT 46.530 91.600 50.480 91.800 ;
        RECT 50.130 91.000 50.480 91.600 ;
        RECT 46.530 90.800 50.480 91.000 ;
        RECT 50.130 90.400 50.480 90.800 ;
        RECT 51.080 90.400 51.280 98.000 ;
        RECT 51.880 90.400 52.080 98.000 ;
        RECT 52.680 90.400 52.880 98.000 ;
        RECT 53.480 90.400 53.680 98.000 ;
        RECT 50.130 89.200 50.480 89.600 ;
        RECT 46.530 89.000 50.480 89.200 ;
        RECT 50.130 88.400 50.480 89.000 ;
        RECT 46.530 88.200 50.480 88.400 ;
        RECT 50.130 87.600 50.480 88.200 ;
        RECT 46.530 87.400 50.480 87.600 ;
        RECT 50.130 86.800 50.480 87.400 ;
        RECT 38.980 86.000 39.330 86.600 ;
        RECT 38.980 85.800 42.930 86.000 ;
        RECT 38.980 85.200 39.330 85.800 ;
        RECT 38.980 85.000 42.930 85.200 ;
        RECT 38.980 84.400 39.330 85.000 ;
        RECT 43.880 84.450 45.580 86.750 ;
        RECT 46.530 86.600 50.480 86.800 ;
        RECT 50.130 86.000 50.480 86.600 ;
        RECT 46.530 85.800 50.480 86.000 ;
        RECT 50.130 85.200 50.480 85.800 ;
        RECT 46.530 85.000 50.480 85.200 ;
        RECT 38.980 84.200 42.930 84.400 ;
        RECT 38.980 83.600 39.330 84.200 ;
        RECT 38.980 83.400 42.930 83.600 ;
        RECT 38.980 82.800 39.330 83.400 ;
        RECT 38.980 82.600 42.930 82.800 ;
        RECT 38.980 82.000 39.330 82.600 ;
        RECT 26.530 81.400 42.930 82.000 ;
        RECT 29.180 80.800 31.480 80.850 ;
        RECT 37.980 80.800 40.280 80.850 ;
        RECT 43.930 80.800 44.330 84.450 ;
        RECT 25.130 80.400 44.330 80.800 ;
        RECT 45.130 80.800 45.530 84.450 ;
        RECT 50.130 84.400 50.480 85.000 ;
        RECT 46.530 84.200 50.480 84.400 ;
        RECT 50.130 83.600 50.480 84.200 ;
        RECT 46.530 83.400 50.480 83.600 ;
        RECT 50.130 82.800 50.480 83.400 ;
        RECT 46.530 82.600 50.480 82.800 ;
        RECT 50.130 82.000 50.480 82.600 ;
        RECT 51.080 82.000 51.280 89.600 ;
        RECT 51.880 82.000 52.080 89.600 ;
        RECT 52.680 82.000 52.880 89.600 ;
        RECT 53.480 82.000 53.680 89.600 ;
        RECT 54.280 82.000 55.180 98.000 ;
        RECT 55.780 90.400 55.980 98.000 ;
        RECT 56.580 90.400 56.780 98.000 ;
        RECT 57.380 90.400 57.580 98.000 ;
        RECT 58.180 90.400 58.380 98.000 ;
        RECT 58.980 97.400 59.330 98.000 ;
        RECT 58.980 97.200 62.930 97.400 ;
        RECT 58.980 96.600 59.330 97.200 ;
        RECT 58.980 96.400 62.930 96.600 ;
        RECT 58.980 95.800 59.330 96.400 ;
        RECT 58.980 95.600 62.930 95.800 ;
        RECT 58.980 95.000 59.330 95.600 ;
        RECT 63.930 95.550 64.330 99.200 ;
        RECT 65.130 99.200 84.330 99.600 ;
        RECT 65.130 95.550 65.530 99.200 ;
        RECT 69.180 99.150 71.480 99.200 ;
        RECT 77.980 99.150 80.280 99.200 ;
        RECT 66.530 98.000 82.930 98.600 ;
        RECT 70.130 97.400 70.480 98.000 ;
        RECT 66.530 97.200 70.480 97.400 ;
        RECT 70.130 96.600 70.480 97.200 ;
        RECT 66.530 96.400 70.480 96.600 ;
        RECT 70.130 95.800 70.480 96.400 ;
        RECT 66.530 95.600 70.480 95.800 ;
        RECT 58.980 94.800 62.930 95.000 ;
        RECT 58.980 94.200 59.330 94.800 ;
        RECT 58.980 94.000 62.930 94.200 ;
        RECT 58.980 93.400 59.330 94.000 ;
        RECT 58.980 93.200 62.930 93.400 ;
        RECT 63.880 93.250 65.580 95.550 ;
        RECT 70.130 95.000 70.480 95.600 ;
        RECT 66.530 94.800 70.480 95.000 ;
        RECT 70.130 94.200 70.480 94.800 ;
        RECT 66.530 94.000 70.480 94.200 ;
        RECT 70.130 93.400 70.480 94.000 ;
        RECT 58.980 92.600 59.330 93.200 ;
        RECT 58.980 92.400 62.930 92.600 ;
        RECT 58.980 91.800 59.330 92.400 ;
        RECT 58.980 91.600 62.930 91.800 ;
        RECT 58.980 91.000 59.330 91.600 ;
        RECT 58.980 90.800 62.930 91.000 ;
        RECT 58.980 90.400 59.330 90.800 ;
        RECT 55.780 82.000 55.980 89.600 ;
        RECT 56.580 82.000 56.780 89.600 ;
        RECT 57.380 82.000 57.580 89.600 ;
        RECT 58.180 82.000 58.380 89.600 ;
        RECT 58.980 89.200 59.330 89.600 ;
        RECT 58.980 89.000 62.930 89.200 ;
        RECT 58.980 88.400 59.330 89.000 ;
        RECT 58.980 88.200 62.930 88.400 ;
        RECT 58.980 87.600 59.330 88.200 ;
        RECT 58.980 87.400 62.930 87.600 ;
        RECT 58.980 86.800 59.330 87.400 ;
        RECT 58.980 86.600 62.930 86.800 ;
        RECT 63.930 86.750 64.330 93.250 ;
        RECT 65.130 86.750 65.530 93.250 ;
        RECT 66.530 93.200 70.480 93.400 ;
        RECT 70.130 92.600 70.480 93.200 ;
        RECT 66.530 92.400 70.480 92.600 ;
        RECT 70.130 91.800 70.480 92.400 ;
        RECT 66.530 91.600 70.480 91.800 ;
        RECT 70.130 91.000 70.480 91.600 ;
        RECT 66.530 90.800 70.480 91.000 ;
        RECT 70.130 90.400 70.480 90.800 ;
        RECT 71.080 90.400 71.280 98.000 ;
        RECT 71.880 90.400 72.080 98.000 ;
        RECT 72.680 90.400 72.880 98.000 ;
        RECT 73.480 90.400 73.680 98.000 ;
        RECT 70.130 89.200 70.480 89.600 ;
        RECT 66.530 89.000 70.480 89.200 ;
        RECT 70.130 88.400 70.480 89.000 ;
        RECT 66.530 88.200 70.480 88.400 ;
        RECT 70.130 87.600 70.480 88.200 ;
        RECT 66.530 87.400 70.480 87.600 ;
        RECT 70.130 86.800 70.480 87.400 ;
        RECT 58.980 86.000 59.330 86.600 ;
        RECT 58.980 85.800 62.930 86.000 ;
        RECT 58.980 85.200 59.330 85.800 ;
        RECT 58.980 85.000 62.930 85.200 ;
        RECT 58.980 84.400 59.330 85.000 ;
        RECT 63.880 84.450 65.580 86.750 ;
        RECT 66.530 86.600 70.480 86.800 ;
        RECT 70.130 86.000 70.480 86.600 ;
        RECT 66.530 85.800 70.480 86.000 ;
        RECT 70.130 85.200 70.480 85.800 ;
        RECT 66.530 85.000 70.480 85.200 ;
        RECT 58.980 84.200 62.930 84.400 ;
        RECT 58.980 83.600 59.330 84.200 ;
        RECT 58.980 83.400 62.930 83.600 ;
        RECT 58.980 82.800 59.330 83.400 ;
        RECT 58.980 82.600 62.930 82.800 ;
        RECT 58.980 82.000 59.330 82.600 ;
        RECT 46.530 81.400 62.930 82.000 ;
        RECT 49.180 80.800 51.480 80.850 ;
        RECT 57.980 80.800 60.280 80.850 ;
        RECT 63.930 80.800 64.330 84.450 ;
        RECT 45.130 80.400 64.330 80.800 ;
        RECT 65.130 80.800 65.530 84.450 ;
        RECT 70.130 84.400 70.480 85.000 ;
        RECT 66.530 84.200 70.480 84.400 ;
        RECT 70.130 83.600 70.480 84.200 ;
        RECT 66.530 83.400 70.480 83.600 ;
        RECT 70.130 82.800 70.480 83.400 ;
        RECT 66.530 82.600 70.480 82.800 ;
        RECT 70.130 82.000 70.480 82.600 ;
        RECT 71.080 82.000 71.280 89.600 ;
        RECT 71.880 82.000 72.080 89.600 ;
        RECT 72.680 82.000 72.880 89.600 ;
        RECT 73.480 82.000 73.680 89.600 ;
        RECT 74.280 82.000 75.180 98.000 ;
        RECT 75.780 90.400 75.980 98.000 ;
        RECT 76.580 90.400 76.780 98.000 ;
        RECT 77.380 90.400 77.580 98.000 ;
        RECT 78.180 90.400 78.380 98.000 ;
        RECT 78.980 97.400 79.330 98.000 ;
        RECT 78.980 97.200 82.930 97.400 ;
        RECT 78.980 96.600 79.330 97.200 ;
        RECT 78.980 96.400 82.930 96.600 ;
        RECT 78.980 95.800 79.330 96.400 ;
        RECT 78.980 95.600 82.930 95.800 ;
        RECT 78.980 95.000 79.330 95.600 ;
        RECT 83.930 95.550 84.330 99.200 ;
        RECT 85.130 99.200 104.330 99.600 ;
        RECT 85.130 95.550 85.530 99.200 ;
        RECT 89.180 99.150 91.480 99.200 ;
        RECT 97.980 99.150 100.280 99.200 ;
        RECT 86.530 98.000 102.930 98.600 ;
        RECT 90.130 97.400 90.480 98.000 ;
        RECT 86.530 97.200 90.480 97.400 ;
        RECT 90.130 96.600 90.480 97.200 ;
        RECT 86.530 96.400 90.480 96.600 ;
        RECT 90.130 95.800 90.480 96.400 ;
        RECT 86.530 95.600 90.480 95.800 ;
        RECT 78.980 94.800 82.930 95.000 ;
        RECT 78.980 94.200 79.330 94.800 ;
        RECT 78.980 94.000 82.930 94.200 ;
        RECT 78.980 93.400 79.330 94.000 ;
        RECT 78.980 93.200 82.930 93.400 ;
        RECT 83.880 93.250 85.580 95.550 ;
        RECT 90.130 95.000 90.480 95.600 ;
        RECT 86.530 94.800 90.480 95.000 ;
        RECT 90.130 94.200 90.480 94.800 ;
        RECT 86.530 94.000 90.480 94.200 ;
        RECT 90.130 93.400 90.480 94.000 ;
        RECT 78.980 92.600 79.330 93.200 ;
        RECT 78.980 92.400 82.930 92.600 ;
        RECT 78.980 91.800 79.330 92.400 ;
        RECT 78.980 91.600 82.930 91.800 ;
        RECT 78.980 91.000 79.330 91.600 ;
        RECT 78.980 90.800 82.930 91.000 ;
        RECT 78.980 90.400 79.330 90.800 ;
        RECT 75.780 82.000 75.980 89.600 ;
        RECT 76.580 82.000 76.780 89.600 ;
        RECT 77.380 82.000 77.580 89.600 ;
        RECT 78.180 82.000 78.380 89.600 ;
        RECT 78.980 89.200 79.330 89.600 ;
        RECT 78.980 89.000 82.930 89.200 ;
        RECT 78.980 88.400 79.330 89.000 ;
        RECT 78.980 88.200 82.930 88.400 ;
        RECT 78.980 87.600 79.330 88.200 ;
        RECT 78.980 87.400 82.930 87.600 ;
        RECT 78.980 86.800 79.330 87.400 ;
        RECT 78.980 86.600 82.930 86.800 ;
        RECT 83.930 86.750 84.330 93.250 ;
        RECT 85.130 86.750 85.530 93.250 ;
        RECT 86.530 93.200 90.480 93.400 ;
        RECT 90.130 92.600 90.480 93.200 ;
        RECT 86.530 92.400 90.480 92.600 ;
        RECT 90.130 91.800 90.480 92.400 ;
        RECT 86.530 91.600 90.480 91.800 ;
        RECT 90.130 91.000 90.480 91.600 ;
        RECT 86.530 90.800 90.480 91.000 ;
        RECT 90.130 90.400 90.480 90.800 ;
        RECT 91.080 90.400 91.280 98.000 ;
        RECT 91.880 90.400 92.080 98.000 ;
        RECT 92.680 90.400 92.880 98.000 ;
        RECT 93.480 90.400 93.680 98.000 ;
        RECT 90.130 89.200 90.480 89.600 ;
        RECT 86.530 89.000 90.480 89.200 ;
        RECT 90.130 88.400 90.480 89.000 ;
        RECT 86.530 88.200 90.480 88.400 ;
        RECT 90.130 87.600 90.480 88.200 ;
        RECT 86.530 87.400 90.480 87.600 ;
        RECT 90.130 86.800 90.480 87.400 ;
        RECT 78.980 86.000 79.330 86.600 ;
        RECT 78.980 85.800 82.930 86.000 ;
        RECT 78.980 85.200 79.330 85.800 ;
        RECT 78.980 85.000 82.930 85.200 ;
        RECT 78.980 84.400 79.330 85.000 ;
        RECT 83.880 84.450 85.580 86.750 ;
        RECT 86.530 86.600 90.480 86.800 ;
        RECT 90.130 86.000 90.480 86.600 ;
        RECT 86.530 85.800 90.480 86.000 ;
        RECT 90.130 85.200 90.480 85.800 ;
        RECT 86.530 85.000 90.480 85.200 ;
        RECT 78.980 84.200 82.930 84.400 ;
        RECT 78.980 83.600 79.330 84.200 ;
        RECT 78.980 83.400 82.930 83.600 ;
        RECT 78.980 82.800 79.330 83.400 ;
        RECT 78.980 82.600 82.930 82.800 ;
        RECT 78.980 82.000 79.330 82.600 ;
        RECT 66.530 81.400 82.930 82.000 ;
        RECT 69.180 80.800 71.480 80.850 ;
        RECT 77.980 80.800 80.280 80.850 ;
        RECT 83.930 80.800 84.330 84.450 ;
        RECT 65.130 80.400 84.330 80.800 ;
        RECT 85.130 80.800 85.530 84.450 ;
        RECT 90.130 84.400 90.480 85.000 ;
        RECT 86.530 84.200 90.480 84.400 ;
        RECT 90.130 83.600 90.480 84.200 ;
        RECT 86.530 83.400 90.480 83.600 ;
        RECT 90.130 82.800 90.480 83.400 ;
        RECT 86.530 82.600 90.480 82.800 ;
        RECT 90.130 82.000 90.480 82.600 ;
        RECT 91.080 82.000 91.280 89.600 ;
        RECT 91.880 82.000 92.080 89.600 ;
        RECT 92.680 82.000 92.880 89.600 ;
        RECT 93.480 82.000 93.680 89.600 ;
        RECT 94.280 82.000 95.180 98.000 ;
        RECT 95.780 90.400 95.980 98.000 ;
        RECT 96.580 90.400 96.780 98.000 ;
        RECT 97.380 90.400 97.580 98.000 ;
        RECT 98.180 90.400 98.380 98.000 ;
        RECT 98.980 97.400 99.330 98.000 ;
        RECT 98.980 97.200 102.930 97.400 ;
        RECT 98.980 96.600 99.330 97.200 ;
        RECT 98.980 96.400 102.930 96.600 ;
        RECT 98.980 95.800 99.330 96.400 ;
        RECT 98.980 95.600 102.930 95.800 ;
        RECT 98.980 95.000 99.330 95.600 ;
        RECT 103.930 95.550 104.330 99.200 ;
        RECT 105.340 96.680 105.700 97.060 ;
        RECT 105.970 96.680 106.330 97.060 ;
        RECT 106.570 96.680 106.930 97.060 ;
        RECT 105.340 96.090 105.700 96.470 ;
        RECT 105.970 96.090 106.330 96.470 ;
        RECT 106.570 96.090 106.930 96.470 ;
        RECT 98.980 94.800 102.930 95.000 ;
        RECT 98.980 94.200 99.330 94.800 ;
        RECT 98.980 94.000 102.930 94.200 ;
        RECT 98.980 93.400 99.330 94.000 ;
        RECT 98.980 93.200 102.930 93.400 ;
        RECT 103.880 93.250 104.730 95.550 ;
        RECT 98.980 92.600 99.330 93.200 ;
        RECT 98.980 92.400 102.930 92.600 ;
        RECT 98.980 91.800 99.330 92.400 ;
        RECT 98.980 91.600 102.930 91.800 ;
        RECT 98.980 91.000 99.330 91.600 ;
        RECT 98.980 90.800 102.930 91.000 ;
        RECT 98.980 90.400 99.330 90.800 ;
        RECT 95.780 82.000 95.980 89.600 ;
        RECT 96.580 82.000 96.780 89.600 ;
        RECT 97.380 82.000 97.580 89.600 ;
        RECT 98.180 82.000 98.380 89.600 ;
        RECT 98.980 89.200 99.330 89.600 ;
        RECT 98.980 89.000 102.930 89.200 ;
        RECT 98.980 88.400 99.330 89.000 ;
        RECT 98.980 88.200 102.930 88.400 ;
        RECT 98.980 87.600 99.330 88.200 ;
        RECT 98.980 87.400 102.930 87.600 ;
        RECT 98.980 86.800 99.330 87.400 ;
        RECT 98.980 86.600 102.930 86.800 ;
        RECT 103.930 86.750 104.330 93.250 ;
        RECT 98.980 86.000 99.330 86.600 ;
        RECT 98.980 85.800 102.930 86.000 ;
        RECT 98.980 85.200 99.330 85.800 ;
        RECT 98.980 85.000 102.930 85.200 ;
        RECT 98.980 84.400 99.330 85.000 ;
        RECT 103.880 84.450 104.730 86.750 ;
        RECT 98.980 84.200 102.930 84.400 ;
        RECT 98.980 83.600 99.330 84.200 ;
        RECT 98.980 83.400 102.930 83.600 ;
        RECT 98.980 82.800 99.330 83.400 ;
        RECT 98.980 82.600 102.930 82.800 ;
        RECT 98.980 82.000 99.330 82.600 ;
        RECT 86.530 81.400 102.930 82.000 ;
        RECT 89.180 80.800 91.480 80.850 ;
        RECT 97.980 80.800 100.280 80.850 ;
        RECT 103.930 80.800 104.330 84.450 ;
        RECT 105.340 82.875 105.700 83.255 ;
        RECT 105.970 82.875 106.330 83.255 ;
        RECT 106.570 82.875 106.930 83.255 ;
        RECT 105.340 82.285 105.700 82.665 ;
        RECT 105.970 82.285 106.330 82.665 ;
        RECT 106.570 82.285 106.930 82.665 ;
        RECT 85.130 80.400 104.330 80.800 ;
        RECT 9.180 79.600 11.480 80.400 ;
        RECT 17.980 79.600 20.280 80.400 ;
        RECT 29.180 79.600 31.480 80.400 ;
        RECT 37.980 79.600 40.280 80.400 ;
        RECT 49.180 79.600 51.480 80.400 ;
        RECT 57.980 79.600 60.280 80.400 ;
        RECT 69.180 79.600 71.480 80.400 ;
        RECT 77.980 79.600 80.280 80.400 ;
        RECT 89.180 79.600 91.480 80.400 ;
        RECT 97.980 79.600 100.280 80.400 ;
        RECT 5.130 79.200 24.330 79.600 ;
        RECT 2.515 77.050 2.875 77.430 ;
        RECT 3.145 77.050 3.505 77.430 ;
        RECT 3.745 77.050 4.105 77.430 ;
        RECT 2.515 76.460 2.875 76.840 ;
        RECT 3.145 76.460 3.505 76.840 ;
        RECT 3.745 76.460 4.105 76.840 ;
        RECT 5.130 75.550 5.530 79.200 ;
        RECT 9.180 79.150 11.480 79.200 ;
        RECT 17.980 79.150 20.280 79.200 ;
        RECT 6.530 78.000 22.930 78.600 ;
        RECT 10.130 77.400 10.480 78.000 ;
        RECT 6.530 77.200 10.480 77.400 ;
        RECT 10.130 76.600 10.480 77.200 ;
        RECT 6.530 76.400 10.480 76.600 ;
        RECT 10.130 75.800 10.480 76.400 ;
        RECT 6.530 75.600 10.480 75.800 ;
        RECT 4.730 75.545 5.580 75.550 ;
        RECT 2.315 73.250 5.580 75.545 ;
        RECT 10.130 75.000 10.480 75.600 ;
        RECT 6.530 74.800 10.480 75.000 ;
        RECT 10.130 74.200 10.480 74.800 ;
        RECT 6.530 74.000 10.480 74.200 ;
        RECT 10.130 73.400 10.480 74.000 ;
        RECT 5.130 66.750 5.530 73.250 ;
        RECT 6.530 73.200 10.480 73.400 ;
        RECT 10.130 72.600 10.480 73.200 ;
        RECT 6.530 72.400 10.480 72.600 ;
        RECT 10.130 71.800 10.480 72.400 ;
        RECT 6.530 71.600 10.480 71.800 ;
        RECT 10.130 71.000 10.480 71.600 ;
        RECT 6.530 70.800 10.480 71.000 ;
        RECT 10.130 70.400 10.480 70.800 ;
        RECT 11.080 70.400 11.280 78.000 ;
        RECT 11.880 70.400 12.080 78.000 ;
        RECT 12.680 70.400 12.880 78.000 ;
        RECT 13.480 70.400 13.680 78.000 ;
        RECT 10.130 69.200 10.480 69.600 ;
        RECT 6.530 69.000 10.480 69.200 ;
        RECT 10.130 68.400 10.480 69.000 ;
        RECT 6.530 68.200 10.480 68.400 ;
        RECT 10.130 67.600 10.480 68.200 ;
        RECT 6.530 67.400 10.480 67.600 ;
        RECT 10.130 66.800 10.480 67.400 ;
        RECT 4.730 66.745 5.580 66.750 ;
        RECT 2.315 64.450 5.580 66.745 ;
        RECT 6.530 66.600 10.480 66.800 ;
        RECT 10.130 66.000 10.480 66.600 ;
        RECT 6.530 65.800 10.480 66.000 ;
        RECT 10.130 65.200 10.480 65.800 ;
        RECT 6.530 65.000 10.480 65.200 ;
        RECT 2.515 62.725 2.875 63.105 ;
        RECT 3.145 62.725 3.505 63.105 ;
        RECT 3.745 62.725 4.105 63.105 ;
        RECT 2.515 62.135 2.875 62.515 ;
        RECT 3.145 62.135 3.505 62.515 ;
        RECT 3.745 62.135 4.105 62.515 ;
        RECT 5.130 60.800 5.530 64.450 ;
        RECT 10.130 64.400 10.480 65.000 ;
        RECT 6.530 64.200 10.480 64.400 ;
        RECT 10.130 63.600 10.480 64.200 ;
        RECT 6.530 63.400 10.480 63.600 ;
        RECT 10.130 62.800 10.480 63.400 ;
        RECT 6.530 62.600 10.480 62.800 ;
        RECT 10.130 62.000 10.480 62.600 ;
        RECT 11.080 62.000 11.280 69.600 ;
        RECT 11.880 62.000 12.080 69.600 ;
        RECT 12.680 62.000 12.880 69.600 ;
        RECT 13.480 62.000 13.680 69.600 ;
        RECT 14.280 62.000 15.180 78.000 ;
        RECT 15.780 70.400 15.980 78.000 ;
        RECT 16.580 70.400 16.780 78.000 ;
        RECT 17.380 70.400 17.580 78.000 ;
        RECT 18.180 70.400 18.380 78.000 ;
        RECT 18.980 77.400 19.330 78.000 ;
        RECT 18.980 77.200 22.930 77.400 ;
        RECT 18.980 76.600 19.330 77.200 ;
        RECT 18.980 76.400 22.930 76.600 ;
        RECT 18.980 75.800 19.330 76.400 ;
        RECT 18.980 75.600 22.930 75.800 ;
        RECT 18.980 75.000 19.330 75.600 ;
        RECT 23.930 75.550 24.330 79.200 ;
        RECT 25.130 79.200 44.330 79.600 ;
        RECT 25.130 75.550 25.530 79.200 ;
        RECT 29.180 79.150 31.480 79.200 ;
        RECT 37.980 79.150 40.280 79.200 ;
        RECT 26.530 78.000 42.930 78.600 ;
        RECT 30.130 77.400 30.480 78.000 ;
        RECT 26.530 77.200 30.480 77.400 ;
        RECT 30.130 76.600 30.480 77.200 ;
        RECT 26.530 76.400 30.480 76.600 ;
        RECT 30.130 75.800 30.480 76.400 ;
        RECT 26.530 75.600 30.480 75.800 ;
        RECT 18.980 74.800 22.930 75.000 ;
        RECT 18.980 74.200 19.330 74.800 ;
        RECT 18.980 74.000 22.930 74.200 ;
        RECT 18.980 73.400 19.330 74.000 ;
        RECT 18.980 73.200 22.930 73.400 ;
        RECT 23.880 73.250 25.580 75.550 ;
        RECT 30.130 75.000 30.480 75.600 ;
        RECT 26.530 74.800 30.480 75.000 ;
        RECT 30.130 74.200 30.480 74.800 ;
        RECT 26.530 74.000 30.480 74.200 ;
        RECT 30.130 73.400 30.480 74.000 ;
        RECT 18.980 72.600 19.330 73.200 ;
        RECT 18.980 72.400 22.930 72.600 ;
        RECT 18.980 71.800 19.330 72.400 ;
        RECT 18.980 71.600 22.930 71.800 ;
        RECT 18.980 71.000 19.330 71.600 ;
        RECT 18.980 70.800 22.930 71.000 ;
        RECT 18.980 70.400 19.330 70.800 ;
        RECT 15.780 62.000 15.980 69.600 ;
        RECT 16.580 62.000 16.780 69.600 ;
        RECT 17.380 62.000 17.580 69.600 ;
        RECT 18.180 62.000 18.380 69.600 ;
        RECT 18.980 69.200 19.330 69.600 ;
        RECT 18.980 69.000 22.930 69.200 ;
        RECT 18.980 68.400 19.330 69.000 ;
        RECT 18.980 68.200 22.930 68.400 ;
        RECT 18.980 67.600 19.330 68.200 ;
        RECT 18.980 67.400 22.930 67.600 ;
        RECT 18.980 66.800 19.330 67.400 ;
        RECT 18.980 66.600 22.930 66.800 ;
        RECT 23.930 66.750 24.330 73.250 ;
        RECT 25.130 66.750 25.530 73.250 ;
        RECT 26.530 73.200 30.480 73.400 ;
        RECT 30.130 72.600 30.480 73.200 ;
        RECT 26.530 72.400 30.480 72.600 ;
        RECT 30.130 71.800 30.480 72.400 ;
        RECT 26.530 71.600 30.480 71.800 ;
        RECT 30.130 71.000 30.480 71.600 ;
        RECT 26.530 70.800 30.480 71.000 ;
        RECT 30.130 70.400 30.480 70.800 ;
        RECT 31.080 70.400 31.280 78.000 ;
        RECT 31.880 70.400 32.080 78.000 ;
        RECT 32.680 70.400 32.880 78.000 ;
        RECT 33.480 70.400 33.680 78.000 ;
        RECT 30.130 69.200 30.480 69.600 ;
        RECT 26.530 69.000 30.480 69.200 ;
        RECT 30.130 68.400 30.480 69.000 ;
        RECT 26.530 68.200 30.480 68.400 ;
        RECT 30.130 67.600 30.480 68.200 ;
        RECT 26.530 67.400 30.480 67.600 ;
        RECT 30.130 66.800 30.480 67.400 ;
        RECT 18.980 66.000 19.330 66.600 ;
        RECT 18.980 65.800 22.930 66.000 ;
        RECT 18.980 65.200 19.330 65.800 ;
        RECT 18.980 65.000 22.930 65.200 ;
        RECT 18.980 64.400 19.330 65.000 ;
        RECT 23.880 64.450 25.580 66.750 ;
        RECT 26.530 66.600 30.480 66.800 ;
        RECT 30.130 66.000 30.480 66.600 ;
        RECT 26.530 65.800 30.480 66.000 ;
        RECT 30.130 65.200 30.480 65.800 ;
        RECT 26.530 65.000 30.480 65.200 ;
        RECT 18.980 64.200 22.930 64.400 ;
        RECT 18.980 63.600 19.330 64.200 ;
        RECT 18.980 63.400 22.930 63.600 ;
        RECT 18.980 62.800 19.330 63.400 ;
        RECT 18.980 62.600 22.930 62.800 ;
        RECT 18.980 62.000 19.330 62.600 ;
        RECT 6.530 61.400 22.930 62.000 ;
        RECT 9.180 60.800 11.480 60.850 ;
        RECT 17.980 60.800 20.280 60.850 ;
        RECT 23.930 60.800 24.330 64.450 ;
        RECT 5.130 60.400 24.330 60.800 ;
        RECT 25.130 60.800 25.530 64.450 ;
        RECT 30.130 64.400 30.480 65.000 ;
        RECT 26.530 64.200 30.480 64.400 ;
        RECT 30.130 63.600 30.480 64.200 ;
        RECT 26.530 63.400 30.480 63.600 ;
        RECT 30.130 62.800 30.480 63.400 ;
        RECT 26.530 62.600 30.480 62.800 ;
        RECT 30.130 62.000 30.480 62.600 ;
        RECT 31.080 62.000 31.280 69.600 ;
        RECT 31.880 62.000 32.080 69.600 ;
        RECT 32.680 62.000 32.880 69.600 ;
        RECT 33.480 62.000 33.680 69.600 ;
        RECT 34.280 62.000 35.180 78.000 ;
        RECT 35.780 70.400 35.980 78.000 ;
        RECT 36.580 70.400 36.780 78.000 ;
        RECT 37.380 70.400 37.580 78.000 ;
        RECT 38.180 70.400 38.380 78.000 ;
        RECT 38.980 77.400 39.330 78.000 ;
        RECT 38.980 77.200 42.930 77.400 ;
        RECT 38.980 76.600 39.330 77.200 ;
        RECT 38.980 76.400 42.930 76.600 ;
        RECT 38.980 75.800 39.330 76.400 ;
        RECT 38.980 75.600 42.930 75.800 ;
        RECT 38.980 75.000 39.330 75.600 ;
        RECT 43.930 75.550 44.330 79.200 ;
        RECT 45.130 79.200 64.330 79.600 ;
        RECT 45.130 75.550 45.530 79.200 ;
        RECT 49.180 79.150 51.480 79.200 ;
        RECT 57.980 79.150 60.280 79.200 ;
        RECT 46.530 78.000 62.930 78.600 ;
        RECT 50.130 77.400 50.480 78.000 ;
        RECT 46.530 77.200 50.480 77.400 ;
        RECT 50.130 76.600 50.480 77.200 ;
        RECT 46.530 76.400 50.480 76.600 ;
        RECT 50.130 75.800 50.480 76.400 ;
        RECT 46.530 75.600 50.480 75.800 ;
        RECT 38.980 74.800 42.930 75.000 ;
        RECT 38.980 74.200 39.330 74.800 ;
        RECT 38.980 74.000 42.930 74.200 ;
        RECT 38.980 73.400 39.330 74.000 ;
        RECT 38.980 73.200 42.930 73.400 ;
        RECT 43.880 73.250 45.580 75.550 ;
        RECT 50.130 75.000 50.480 75.600 ;
        RECT 46.530 74.800 50.480 75.000 ;
        RECT 50.130 74.200 50.480 74.800 ;
        RECT 46.530 74.000 50.480 74.200 ;
        RECT 50.130 73.400 50.480 74.000 ;
        RECT 38.980 72.600 39.330 73.200 ;
        RECT 38.980 72.400 42.930 72.600 ;
        RECT 38.980 71.800 39.330 72.400 ;
        RECT 38.980 71.600 42.930 71.800 ;
        RECT 38.980 71.000 39.330 71.600 ;
        RECT 38.980 70.800 42.930 71.000 ;
        RECT 38.980 70.400 39.330 70.800 ;
        RECT 35.780 62.000 35.980 69.600 ;
        RECT 36.580 62.000 36.780 69.600 ;
        RECT 37.380 62.000 37.580 69.600 ;
        RECT 38.180 62.000 38.380 69.600 ;
        RECT 38.980 69.200 39.330 69.600 ;
        RECT 38.980 69.000 42.930 69.200 ;
        RECT 38.980 68.400 39.330 69.000 ;
        RECT 38.980 68.200 42.930 68.400 ;
        RECT 38.980 67.600 39.330 68.200 ;
        RECT 38.980 67.400 42.930 67.600 ;
        RECT 38.980 66.800 39.330 67.400 ;
        RECT 38.980 66.600 42.930 66.800 ;
        RECT 43.930 66.750 44.330 73.250 ;
        RECT 45.130 66.750 45.530 73.250 ;
        RECT 46.530 73.200 50.480 73.400 ;
        RECT 50.130 72.600 50.480 73.200 ;
        RECT 46.530 72.400 50.480 72.600 ;
        RECT 50.130 71.800 50.480 72.400 ;
        RECT 46.530 71.600 50.480 71.800 ;
        RECT 50.130 71.000 50.480 71.600 ;
        RECT 46.530 70.800 50.480 71.000 ;
        RECT 50.130 70.400 50.480 70.800 ;
        RECT 51.080 70.400 51.280 78.000 ;
        RECT 51.880 70.400 52.080 78.000 ;
        RECT 52.680 70.400 52.880 78.000 ;
        RECT 53.480 70.400 53.680 78.000 ;
        RECT 50.130 69.200 50.480 69.600 ;
        RECT 46.530 69.000 50.480 69.200 ;
        RECT 50.130 68.400 50.480 69.000 ;
        RECT 46.530 68.200 50.480 68.400 ;
        RECT 50.130 67.600 50.480 68.200 ;
        RECT 46.530 67.400 50.480 67.600 ;
        RECT 50.130 66.800 50.480 67.400 ;
        RECT 38.980 66.000 39.330 66.600 ;
        RECT 38.980 65.800 42.930 66.000 ;
        RECT 38.980 65.200 39.330 65.800 ;
        RECT 38.980 65.000 42.930 65.200 ;
        RECT 38.980 64.400 39.330 65.000 ;
        RECT 43.880 64.450 45.580 66.750 ;
        RECT 46.530 66.600 50.480 66.800 ;
        RECT 50.130 66.000 50.480 66.600 ;
        RECT 46.530 65.800 50.480 66.000 ;
        RECT 50.130 65.200 50.480 65.800 ;
        RECT 46.530 65.000 50.480 65.200 ;
        RECT 38.980 64.200 42.930 64.400 ;
        RECT 38.980 63.600 39.330 64.200 ;
        RECT 38.980 63.400 42.930 63.600 ;
        RECT 38.980 62.800 39.330 63.400 ;
        RECT 38.980 62.600 42.930 62.800 ;
        RECT 38.980 62.000 39.330 62.600 ;
        RECT 26.530 61.400 42.930 62.000 ;
        RECT 29.180 60.800 31.480 60.850 ;
        RECT 37.980 60.800 40.280 60.850 ;
        RECT 43.930 60.800 44.330 64.450 ;
        RECT 25.130 60.400 44.330 60.800 ;
        RECT 45.130 60.800 45.530 64.450 ;
        RECT 50.130 64.400 50.480 65.000 ;
        RECT 46.530 64.200 50.480 64.400 ;
        RECT 50.130 63.600 50.480 64.200 ;
        RECT 46.530 63.400 50.480 63.600 ;
        RECT 50.130 62.800 50.480 63.400 ;
        RECT 46.530 62.600 50.480 62.800 ;
        RECT 50.130 62.000 50.480 62.600 ;
        RECT 51.080 62.000 51.280 69.600 ;
        RECT 51.880 62.000 52.080 69.600 ;
        RECT 52.680 62.000 52.880 69.600 ;
        RECT 53.480 62.000 53.680 69.600 ;
        RECT 54.280 62.000 55.180 78.000 ;
        RECT 55.780 70.400 55.980 78.000 ;
        RECT 56.580 70.400 56.780 78.000 ;
        RECT 57.380 70.400 57.580 78.000 ;
        RECT 58.180 70.400 58.380 78.000 ;
        RECT 58.980 77.400 59.330 78.000 ;
        RECT 58.980 77.200 62.930 77.400 ;
        RECT 58.980 76.600 59.330 77.200 ;
        RECT 58.980 76.400 62.930 76.600 ;
        RECT 58.980 75.800 59.330 76.400 ;
        RECT 58.980 75.600 62.930 75.800 ;
        RECT 58.980 75.000 59.330 75.600 ;
        RECT 63.930 75.550 64.330 79.200 ;
        RECT 65.130 79.200 84.330 79.600 ;
        RECT 65.130 75.550 65.530 79.200 ;
        RECT 69.180 79.150 71.480 79.200 ;
        RECT 77.980 79.150 80.280 79.200 ;
        RECT 66.530 78.000 82.930 78.600 ;
        RECT 70.130 77.400 70.480 78.000 ;
        RECT 66.530 77.200 70.480 77.400 ;
        RECT 70.130 76.600 70.480 77.200 ;
        RECT 66.530 76.400 70.480 76.600 ;
        RECT 70.130 75.800 70.480 76.400 ;
        RECT 66.530 75.600 70.480 75.800 ;
        RECT 58.980 74.800 62.930 75.000 ;
        RECT 58.980 74.200 59.330 74.800 ;
        RECT 58.980 74.000 62.930 74.200 ;
        RECT 58.980 73.400 59.330 74.000 ;
        RECT 58.980 73.200 62.930 73.400 ;
        RECT 63.880 73.250 65.580 75.550 ;
        RECT 70.130 75.000 70.480 75.600 ;
        RECT 66.530 74.800 70.480 75.000 ;
        RECT 70.130 74.200 70.480 74.800 ;
        RECT 66.530 74.000 70.480 74.200 ;
        RECT 70.130 73.400 70.480 74.000 ;
        RECT 58.980 72.600 59.330 73.200 ;
        RECT 58.980 72.400 62.930 72.600 ;
        RECT 58.980 71.800 59.330 72.400 ;
        RECT 58.980 71.600 62.930 71.800 ;
        RECT 58.980 71.000 59.330 71.600 ;
        RECT 58.980 70.800 62.930 71.000 ;
        RECT 58.980 70.400 59.330 70.800 ;
        RECT 55.780 62.000 55.980 69.600 ;
        RECT 56.580 62.000 56.780 69.600 ;
        RECT 57.380 62.000 57.580 69.600 ;
        RECT 58.180 62.000 58.380 69.600 ;
        RECT 58.980 69.200 59.330 69.600 ;
        RECT 58.980 69.000 62.930 69.200 ;
        RECT 58.980 68.400 59.330 69.000 ;
        RECT 58.980 68.200 62.930 68.400 ;
        RECT 58.980 67.600 59.330 68.200 ;
        RECT 58.980 67.400 62.930 67.600 ;
        RECT 58.980 66.800 59.330 67.400 ;
        RECT 58.980 66.600 62.930 66.800 ;
        RECT 63.930 66.750 64.330 73.250 ;
        RECT 65.130 66.750 65.530 73.250 ;
        RECT 66.530 73.200 70.480 73.400 ;
        RECT 70.130 72.600 70.480 73.200 ;
        RECT 66.530 72.400 70.480 72.600 ;
        RECT 70.130 71.800 70.480 72.400 ;
        RECT 66.530 71.600 70.480 71.800 ;
        RECT 70.130 71.000 70.480 71.600 ;
        RECT 66.530 70.800 70.480 71.000 ;
        RECT 70.130 70.400 70.480 70.800 ;
        RECT 71.080 70.400 71.280 78.000 ;
        RECT 71.880 70.400 72.080 78.000 ;
        RECT 72.680 70.400 72.880 78.000 ;
        RECT 73.480 70.400 73.680 78.000 ;
        RECT 70.130 69.200 70.480 69.600 ;
        RECT 66.530 69.000 70.480 69.200 ;
        RECT 70.130 68.400 70.480 69.000 ;
        RECT 66.530 68.200 70.480 68.400 ;
        RECT 70.130 67.600 70.480 68.200 ;
        RECT 66.530 67.400 70.480 67.600 ;
        RECT 70.130 66.800 70.480 67.400 ;
        RECT 58.980 66.000 59.330 66.600 ;
        RECT 58.980 65.800 62.930 66.000 ;
        RECT 58.980 65.200 59.330 65.800 ;
        RECT 58.980 65.000 62.930 65.200 ;
        RECT 58.980 64.400 59.330 65.000 ;
        RECT 63.880 64.450 65.580 66.750 ;
        RECT 66.530 66.600 70.480 66.800 ;
        RECT 70.130 66.000 70.480 66.600 ;
        RECT 66.530 65.800 70.480 66.000 ;
        RECT 70.130 65.200 70.480 65.800 ;
        RECT 66.530 65.000 70.480 65.200 ;
        RECT 58.980 64.200 62.930 64.400 ;
        RECT 58.980 63.600 59.330 64.200 ;
        RECT 58.980 63.400 62.930 63.600 ;
        RECT 58.980 62.800 59.330 63.400 ;
        RECT 58.980 62.600 62.930 62.800 ;
        RECT 58.980 62.000 59.330 62.600 ;
        RECT 46.530 61.400 62.930 62.000 ;
        RECT 49.180 60.800 51.480 60.850 ;
        RECT 57.980 60.800 60.280 60.850 ;
        RECT 63.930 60.800 64.330 64.450 ;
        RECT 45.130 60.400 64.330 60.800 ;
        RECT 65.130 60.800 65.530 64.450 ;
        RECT 70.130 64.400 70.480 65.000 ;
        RECT 66.530 64.200 70.480 64.400 ;
        RECT 70.130 63.600 70.480 64.200 ;
        RECT 66.530 63.400 70.480 63.600 ;
        RECT 70.130 62.800 70.480 63.400 ;
        RECT 66.530 62.600 70.480 62.800 ;
        RECT 70.130 62.000 70.480 62.600 ;
        RECT 71.080 62.000 71.280 69.600 ;
        RECT 71.880 62.000 72.080 69.600 ;
        RECT 72.680 62.000 72.880 69.600 ;
        RECT 73.480 62.000 73.680 69.600 ;
        RECT 74.280 62.000 75.180 78.000 ;
        RECT 75.780 70.400 75.980 78.000 ;
        RECT 76.580 70.400 76.780 78.000 ;
        RECT 77.380 70.400 77.580 78.000 ;
        RECT 78.180 70.400 78.380 78.000 ;
        RECT 78.980 77.400 79.330 78.000 ;
        RECT 78.980 77.200 82.930 77.400 ;
        RECT 78.980 76.600 79.330 77.200 ;
        RECT 78.980 76.400 82.930 76.600 ;
        RECT 78.980 75.800 79.330 76.400 ;
        RECT 78.980 75.600 82.930 75.800 ;
        RECT 78.980 75.000 79.330 75.600 ;
        RECT 83.930 75.550 84.330 79.200 ;
        RECT 85.130 79.200 104.330 79.600 ;
        RECT 85.130 75.550 85.530 79.200 ;
        RECT 89.180 79.150 91.480 79.200 ;
        RECT 97.980 79.150 100.280 79.200 ;
        RECT 86.530 78.000 102.930 78.600 ;
        RECT 90.130 77.400 90.480 78.000 ;
        RECT 86.530 77.200 90.480 77.400 ;
        RECT 90.130 76.600 90.480 77.200 ;
        RECT 86.530 76.400 90.480 76.600 ;
        RECT 90.130 75.800 90.480 76.400 ;
        RECT 86.530 75.600 90.480 75.800 ;
        RECT 78.980 74.800 82.930 75.000 ;
        RECT 78.980 74.200 79.330 74.800 ;
        RECT 78.980 74.000 82.930 74.200 ;
        RECT 78.980 73.400 79.330 74.000 ;
        RECT 78.980 73.200 82.930 73.400 ;
        RECT 83.880 73.250 85.580 75.550 ;
        RECT 90.130 75.000 90.480 75.600 ;
        RECT 86.530 74.800 90.480 75.000 ;
        RECT 90.130 74.200 90.480 74.800 ;
        RECT 86.530 74.000 90.480 74.200 ;
        RECT 90.130 73.400 90.480 74.000 ;
        RECT 78.980 72.600 79.330 73.200 ;
        RECT 78.980 72.400 82.930 72.600 ;
        RECT 78.980 71.800 79.330 72.400 ;
        RECT 78.980 71.600 82.930 71.800 ;
        RECT 78.980 71.000 79.330 71.600 ;
        RECT 78.980 70.800 82.930 71.000 ;
        RECT 78.980 70.400 79.330 70.800 ;
        RECT 75.780 62.000 75.980 69.600 ;
        RECT 76.580 62.000 76.780 69.600 ;
        RECT 77.380 62.000 77.580 69.600 ;
        RECT 78.180 62.000 78.380 69.600 ;
        RECT 78.980 69.200 79.330 69.600 ;
        RECT 78.980 69.000 82.930 69.200 ;
        RECT 78.980 68.400 79.330 69.000 ;
        RECT 78.980 68.200 82.930 68.400 ;
        RECT 78.980 67.600 79.330 68.200 ;
        RECT 78.980 67.400 82.930 67.600 ;
        RECT 78.980 66.800 79.330 67.400 ;
        RECT 78.980 66.600 82.930 66.800 ;
        RECT 83.930 66.750 84.330 73.250 ;
        RECT 85.130 66.750 85.530 73.250 ;
        RECT 86.530 73.200 90.480 73.400 ;
        RECT 90.130 72.600 90.480 73.200 ;
        RECT 86.530 72.400 90.480 72.600 ;
        RECT 90.130 71.800 90.480 72.400 ;
        RECT 86.530 71.600 90.480 71.800 ;
        RECT 90.130 71.000 90.480 71.600 ;
        RECT 86.530 70.800 90.480 71.000 ;
        RECT 90.130 70.400 90.480 70.800 ;
        RECT 91.080 70.400 91.280 78.000 ;
        RECT 91.880 70.400 92.080 78.000 ;
        RECT 92.680 70.400 92.880 78.000 ;
        RECT 93.480 70.400 93.680 78.000 ;
        RECT 90.130 69.200 90.480 69.600 ;
        RECT 86.530 69.000 90.480 69.200 ;
        RECT 90.130 68.400 90.480 69.000 ;
        RECT 86.530 68.200 90.480 68.400 ;
        RECT 90.130 67.600 90.480 68.200 ;
        RECT 86.530 67.400 90.480 67.600 ;
        RECT 90.130 66.800 90.480 67.400 ;
        RECT 78.980 66.000 79.330 66.600 ;
        RECT 78.980 65.800 82.930 66.000 ;
        RECT 78.980 65.200 79.330 65.800 ;
        RECT 78.980 65.000 82.930 65.200 ;
        RECT 78.980 64.400 79.330 65.000 ;
        RECT 83.880 64.450 85.580 66.750 ;
        RECT 86.530 66.600 90.480 66.800 ;
        RECT 90.130 66.000 90.480 66.600 ;
        RECT 86.530 65.800 90.480 66.000 ;
        RECT 90.130 65.200 90.480 65.800 ;
        RECT 86.530 65.000 90.480 65.200 ;
        RECT 78.980 64.200 82.930 64.400 ;
        RECT 78.980 63.600 79.330 64.200 ;
        RECT 78.980 63.400 82.930 63.600 ;
        RECT 78.980 62.800 79.330 63.400 ;
        RECT 78.980 62.600 82.930 62.800 ;
        RECT 78.980 62.000 79.330 62.600 ;
        RECT 66.530 61.400 82.930 62.000 ;
        RECT 69.180 60.800 71.480 60.850 ;
        RECT 77.980 60.800 80.280 60.850 ;
        RECT 83.930 60.800 84.330 64.450 ;
        RECT 65.130 60.400 84.330 60.800 ;
        RECT 85.130 60.800 85.530 64.450 ;
        RECT 90.130 64.400 90.480 65.000 ;
        RECT 86.530 64.200 90.480 64.400 ;
        RECT 90.130 63.600 90.480 64.200 ;
        RECT 86.530 63.400 90.480 63.600 ;
        RECT 90.130 62.800 90.480 63.400 ;
        RECT 86.530 62.600 90.480 62.800 ;
        RECT 90.130 62.000 90.480 62.600 ;
        RECT 91.080 62.000 91.280 69.600 ;
        RECT 91.880 62.000 92.080 69.600 ;
        RECT 92.680 62.000 92.880 69.600 ;
        RECT 93.480 62.000 93.680 69.600 ;
        RECT 94.280 62.000 95.180 78.000 ;
        RECT 95.780 70.400 95.980 78.000 ;
        RECT 96.580 70.400 96.780 78.000 ;
        RECT 97.380 70.400 97.580 78.000 ;
        RECT 98.180 70.400 98.380 78.000 ;
        RECT 98.980 77.400 99.330 78.000 ;
        RECT 98.980 77.200 102.930 77.400 ;
        RECT 98.980 76.600 99.330 77.200 ;
        RECT 98.980 76.400 102.930 76.600 ;
        RECT 98.980 75.800 99.330 76.400 ;
        RECT 98.980 75.600 102.930 75.800 ;
        RECT 98.980 75.000 99.330 75.600 ;
        RECT 103.930 75.550 104.330 79.200 ;
        RECT 105.340 76.805 105.700 77.185 ;
        RECT 105.970 76.805 106.330 77.185 ;
        RECT 106.570 76.805 106.930 77.185 ;
        RECT 105.340 76.215 105.700 76.595 ;
        RECT 105.970 76.215 106.330 76.595 ;
        RECT 106.570 76.215 106.930 76.595 ;
        RECT 98.980 74.800 102.930 75.000 ;
        RECT 98.980 74.200 99.330 74.800 ;
        RECT 98.980 74.000 102.930 74.200 ;
        RECT 98.980 73.400 99.330 74.000 ;
        RECT 98.980 73.200 102.930 73.400 ;
        RECT 103.880 73.250 104.730 75.550 ;
        RECT 98.980 72.600 99.330 73.200 ;
        RECT 98.980 72.400 102.930 72.600 ;
        RECT 98.980 71.800 99.330 72.400 ;
        RECT 98.980 71.600 102.930 71.800 ;
        RECT 98.980 71.000 99.330 71.600 ;
        RECT 98.980 70.800 102.930 71.000 ;
        RECT 98.980 70.400 99.330 70.800 ;
        RECT 95.780 62.000 95.980 69.600 ;
        RECT 96.580 62.000 96.780 69.600 ;
        RECT 97.380 62.000 97.580 69.600 ;
        RECT 98.180 62.000 98.380 69.600 ;
        RECT 98.980 69.200 99.330 69.600 ;
        RECT 98.980 69.000 102.930 69.200 ;
        RECT 98.980 68.400 99.330 69.000 ;
        RECT 98.980 68.200 102.930 68.400 ;
        RECT 98.980 67.600 99.330 68.200 ;
        RECT 98.980 67.400 102.930 67.600 ;
        RECT 98.980 66.800 99.330 67.400 ;
        RECT 98.980 66.600 102.930 66.800 ;
        RECT 103.930 66.750 104.330 73.250 ;
        RECT 98.980 66.000 99.330 66.600 ;
        RECT 98.980 65.800 102.930 66.000 ;
        RECT 98.980 65.200 99.330 65.800 ;
        RECT 98.980 65.000 102.930 65.200 ;
        RECT 98.980 64.400 99.330 65.000 ;
        RECT 103.880 64.450 104.730 66.750 ;
        RECT 98.980 64.200 102.930 64.400 ;
        RECT 98.980 63.600 99.330 64.200 ;
        RECT 98.980 63.400 102.930 63.600 ;
        RECT 98.980 62.800 99.330 63.400 ;
        RECT 98.980 62.600 102.930 62.800 ;
        RECT 98.980 62.000 99.330 62.600 ;
        RECT 86.530 61.400 102.930 62.000 ;
        RECT 89.180 60.800 91.480 60.850 ;
        RECT 97.980 60.800 100.280 60.850 ;
        RECT 103.930 60.800 104.330 64.450 ;
        RECT 105.340 62.590 105.700 62.970 ;
        RECT 105.970 62.590 106.330 62.970 ;
        RECT 106.570 62.590 106.930 62.970 ;
        RECT 105.340 62.000 105.700 62.380 ;
        RECT 105.970 62.000 106.330 62.380 ;
        RECT 106.570 62.000 106.930 62.380 ;
        RECT 85.130 60.400 104.330 60.800 ;
        RECT 9.180 59.600 11.480 60.400 ;
        RECT 17.980 59.600 20.280 60.400 ;
        RECT 29.180 59.600 31.480 60.400 ;
        RECT 37.980 59.600 40.280 60.400 ;
        RECT 49.180 59.600 51.480 60.400 ;
        RECT 57.980 59.600 60.280 60.400 ;
        RECT 69.180 59.600 71.480 60.400 ;
        RECT 77.980 59.600 80.280 60.400 ;
        RECT 89.180 59.600 91.480 60.400 ;
        RECT 97.980 59.600 100.280 60.400 ;
        RECT 5.130 59.200 24.330 59.600 ;
        RECT 2.515 57.115 2.875 57.495 ;
        RECT 3.145 57.115 3.505 57.495 ;
        RECT 3.745 57.115 4.105 57.495 ;
        RECT 2.515 56.525 2.875 56.905 ;
        RECT 3.145 56.525 3.505 56.905 ;
        RECT 3.745 56.525 4.105 56.905 ;
        RECT 5.130 55.550 5.530 59.200 ;
        RECT 9.180 59.150 11.480 59.200 ;
        RECT 17.980 59.150 20.280 59.200 ;
        RECT 6.530 58.000 22.930 58.600 ;
        RECT 10.130 57.400 10.480 58.000 ;
        RECT 6.530 57.200 10.480 57.400 ;
        RECT 10.130 56.600 10.480 57.200 ;
        RECT 6.530 56.400 10.480 56.600 ;
        RECT 10.130 55.800 10.480 56.400 ;
        RECT 6.530 55.600 10.480 55.800 ;
        RECT 2.315 53.255 5.580 55.550 ;
        RECT 10.130 55.000 10.480 55.600 ;
        RECT 6.530 54.800 10.480 55.000 ;
        RECT 10.130 54.200 10.480 54.800 ;
        RECT 6.530 54.000 10.480 54.200 ;
        RECT 10.130 53.400 10.480 54.000 ;
        RECT 4.730 53.250 5.580 53.255 ;
        RECT 5.130 46.750 5.530 53.250 ;
        RECT 6.530 53.200 10.480 53.400 ;
        RECT 10.130 52.600 10.480 53.200 ;
        RECT 6.530 52.400 10.480 52.600 ;
        RECT 10.130 51.800 10.480 52.400 ;
        RECT 6.530 51.600 10.480 51.800 ;
        RECT 10.130 51.000 10.480 51.600 ;
        RECT 6.530 50.800 10.480 51.000 ;
        RECT 10.130 50.400 10.480 50.800 ;
        RECT 11.080 50.400 11.280 58.000 ;
        RECT 11.880 50.400 12.080 58.000 ;
        RECT 12.680 50.400 12.880 58.000 ;
        RECT 13.480 50.400 13.680 58.000 ;
        RECT 10.130 49.200 10.480 49.600 ;
        RECT 6.530 49.000 10.480 49.200 ;
        RECT 10.130 48.400 10.480 49.000 ;
        RECT 6.530 48.200 10.480 48.400 ;
        RECT 10.130 47.600 10.480 48.200 ;
        RECT 6.530 47.400 10.480 47.600 ;
        RECT 10.130 46.800 10.480 47.400 ;
        RECT 4.730 46.740 5.580 46.750 ;
        RECT 2.315 44.450 5.580 46.740 ;
        RECT 6.530 46.600 10.480 46.800 ;
        RECT 10.130 46.000 10.480 46.600 ;
        RECT 6.530 45.800 10.480 46.000 ;
        RECT 10.130 45.200 10.480 45.800 ;
        RECT 6.530 45.000 10.480 45.200 ;
        RECT 2.315 44.445 4.730 44.450 ;
        RECT 2.515 42.815 2.875 43.195 ;
        RECT 3.145 42.815 3.505 43.195 ;
        RECT 3.745 42.815 4.105 43.195 ;
        RECT 2.515 42.225 2.875 42.605 ;
        RECT 3.145 42.225 3.505 42.605 ;
        RECT 3.745 42.225 4.105 42.605 ;
        RECT 5.130 40.800 5.530 44.450 ;
        RECT 10.130 44.400 10.480 45.000 ;
        RECT 6.530 44.200 10.480 44.400 ;
        RECT 10.130 43.600 10.480 44.200 ;
        RECT 6.530 43.400 10.480 43.600 ;
        RECT 10.130 42.800 10.480 43.400 ;
        RECT 6.530 42.600 10.480 42.800 ;
        RECT 10.130 42.000 10.480 42.600 ;
        RECT 11.080 42.000 11.280 49.600 ;
        RECT 11.880 42.000 12.080 49.600 ;
        RECT 12.680 42.000 12.880 49.600 ;
        RECT 13.480 42.000 13.680 49.600 ;
        RECT 14.280 42.000 15.180 58.000 ;
        RECT 15.780 50.400 15.980 58.000 ;
        RECT 16.580 50.400 16.780 58.000 ;
        RECT 17.380 50.400 17.580 58.000 ;
        RECT 18.180 50.400 18.380 58.000 ;
        RECT 18.980 57.400 19.330 58.000 ;
        RECT 18.980 57.200 22.930 57.400 ;
        RECT 18.980 56.600 19.330 57.200 ;
        RECT 18.980 56.400 22.930 56.600 ;
        RECT 18.980 55.800 19.330 56.400 ;
        RECT 18.980 55.600 22.930 55.800 ;
        RECT 18.980 55.000 19.330 55.600 ;
        RECT 23.930 55.550 24.330 59.200 ;
        RECT 25.130 59.200 44.330 59.600 ;
        RECT 25.130 55.550 25.530 59.200 ;
        RECT 29.180 59.150 31.480 59.200 ;
        RECT 37.980 59.150 40.280 59.200 ;
        RECT 26.530 58.000 42.930 58.600 ;
        RECT 30.130 57.400 30.480 58.000 ;
        RECT 26.530 57.200 30.480 57.400 ;
        RECT 30.130 56.600 30.480 57.200 ;
        RECT 26.530 56.400 30.480 56.600 ;
        RECT 30.130 55.800 30.480 56.400 ;
        RECT 26.530 55.600 30.480 55.800 ;
        RECT 18.980 54.800 22.930 55.000 ;
        RECT 18.980 54.200 19.330 54.800 ;
        RECT 18.980 54.000 22.930 54.200 ;
        RECT 18.980 53.400 19.330 54.000 ;
        RECT 18.980 53.200 22.930 53.400 ;
        RECT 23.880 53.250 25.580 55.550 ;
        RECT 30.130 55.000 30.480 55.600 ;
        RECT 26.530 54.800 30.480 55.000 ;
        RECT 30.130 54.200 30.480 54.800 ;
        RECT 26.530 54.000 30.480 54.200 ;
        RECT 30.130 53.400 30.480 54.000 ;
        RECT 18.980 52.600 19.330 53.200 ;
        RECT 18.980 52.400 22.930 52.600 ;
        RECT 18.980 51.800 19.330 52.400 ;
        RECT 18.980 51.600 22.930 51.800 ;
        RECT 18.980 51.000 19.330 51.600 ;
        RECT 18.980 50.800 22.930 51.000 ;
        RECT 18.980 50.400 19.330 50.800 ;
        RECT 15.780 42.000 15.980 49.600 ;
        RECT 16.580 42.000 16.780 49.600 ;
        RECT 17.380 42.000 17.580 49.600 ;
        RECT 18.180 42.000 18.380 49.600 ;
        RECT 18.980 49.200 19.330 49.600 ;
        RECT 18.980 49.000 22.930 49.200 ;
        RECT 18.980 48.400 19.330 49.000 ;
        RECT 18.980 48.200 22.930 48.400 ;
        RECT 18.980 47.600 19.330 48.200 ;
        RECT 18.980 47.400 22.930 47.600 ;
        RECT 18.980 46.800 19.330 47.400 ;
        RECT 18.980 46.600 22.930 46.800 ;
        RECT 23.930 46.750 24.330 53.250 ;
        RECT 25.130 46.750 25.530 53.250 ;
        RECT 26.530 53.200 30.480 53.400 ;
        RECT 30.130 52.600 30.480 53.200 ;
        RECT 26.530 52.400 30.480 52.600 ;
        RECT 30.130 51.800 30.480 52.400 ;
        RECT 26.530 51.600 30.480 51.800 ;
        RECT 30.130 51.000 30.480 51.600 ;
        RECT 26.530 50.800 30.480 51.000 ;
        RECT 30.130 50.400 30.480 50.800 ;
        RECT 31.080 50.400 31.280 58.000 ;
        RECT 31.880 50.400 32.080 58.000 ;
        RECT 32.680 50.400 32.880 58.000 ;
        RECT 33.480 50.400 33.680 58.000 ;
        RECT 30.130 49.200 30.480 49.600 ;
        RECT 26.530 49.000 30.480 49.200 ;
        RECT 30.130 48.400 30.480 49.000 ;
        RECT 26.530 48.200 30.480 48.400 ;
        RECT 30.130 47.600 30.480 48.200 ;
        RECT 26.530 47.400 30.480 47.600 ;
        RECT 30.130 46.800 30.480 47.400 ;
        RECT 18.980 46.000 19.330 46.600 ;
        RECT 18.980 45.800 22.930 46.000 ;
        RECT 18.980 45.200 19.330 45.800 ;
        RECT 18.980 45.000 22.930 45.200 ;
        RECT 18.980 44.400 19.330 45.000 ;
        RECT 23.880 44.450 25.580 46.750 ;
        RECT 26.530 46.600 30.480 46.800 ;
        RECT 30.130 46.000 30.480 46.600 ;
        RECT 26.530 45.800 30.480 46.000 ;
        RECT 30.130 45.200 30.480 45.800 ;
        RECT 26.530 45.000 30.480 45.200 ;
        RECT 18.980 44.200 22.930 44.400 ;
        RECT 18.980 43.600 19.330 44.200 ;
        RECT 18.980 43.400 22.930 43.600 ;
        RECT 18.980 42.800 19.330 43.400 ;
        RECT 18.980 42.600 22.930 42.800 ;
        RECT 18.980 42.000 19.330 42.600 ;
        RECT 6.530 41.400 22.930 42.000 ;
        RECT 9.180 40.800 11.480 40.850 ;
        RECT 17.980 40.800 20.280 40.850 ;
        RECT 23.930 40.800 24.330 44.450 ;
        RECT 5.130 40.400 24.330 40.800 ;
        RECT 25.130 40.800 25.530 44.450 ;
        RECT 30.130 44.400 30.480 45.000 ;
        RECT 26.530 44.200 30.480 44.400 ;
        RECT 30.130 43.600 30.480 44.200 ;
        RECT 26.530 43.400 30.480 43.600 ;
        RECT 30.130 42.800 30.480 43.400 ;
        RECT 26.530 42.600 30.480 42.800 ;
        RECT 30.130 42.000 30.480 42.600 ;
        RECT 31.080 42.000 31.280 49.600 ;
        RECT 31.880 42.000 32.080 49.600 ;
        RECT 32.680 42.000 32.880 49.600 ;
        RECT 33.480 42.000 33.680 49.600 ;
        RECT 34.280 42.000 35.180 58.000 ;
        RECT 35.780 50.400 35.980 58.000 ;
        RECT 36.580 50.400 36.780 58.000 ;
        RECT 37.380 50.400 37.580 58.000 ;
        RECT 38.180 50.400 38.380 58.000 ;
        RECT 38.980 57.400 39.330 58.000 ;
        RECT 38.980 57.200 42.930 57.400 ;
        RECT 38.980 56.600 39.330 57.200 ;
        RECT 38.980 56.400 42.930 56.600 ;
        RECT 38.980 55.800 39.330 56.400 ;
        RECT 38.980 55.600 42.930 55.800 ;
        RECT 38.980 55.000 39.330 55.600 ;
        RECT 43.930 55.550 44.330 59.200 ;
        RECT 45.130 59.200 64.330 59.600 ;
        RECT 45.130 55.550 45.530 59.200 ;
        RECT 49.180 59.150 51.480 59.200 ;
        RECT 57.980 59.150 60.280 59.200 ;
        RECT 46.530 58.000 62.930 58.600 ;
        RECT 50.130 57.400 50.480 58.000 ;
        RECT 46.530 57.200 50.480 57.400 ;
        RECT 50.130 56.600 50.480 57.200 ;
        RECT 46.530 56.400 50.480 56.600 ;
        RECT 50.130 55.800 50.480 56.400 ;
        RECT 46.530 55.600 50.480 55.800 ;
        RECT 38.980 54.800 42.930 55.000 ;
        RECT 38.980 54.200 39.330 54.800 ;
        RECT 38.980 54.000 42.930 54.200 ;
        RECT 38.980 53.400 39.330 54.000 ;
        RECT 38.980 53.200 42.930 53.400 ;
        RECT 43.880 53.250 45.580 55.550 ;
        RECT 50.130 55.000 50.480 55.600 ;
        RECT 46.530 54.800 50.480 55.000 ;
        RECT 50.130 54.200 50.480 54.800 ;
        RECT 46.530 54.000 50.480 54.200 ;
        RECT 50.130 53.400 50.480 54.000 ;
        RECT 38.980 52.600 39.330 53.200 ;
        RECT 38.980 52.400 42.930 52.600 ;
        RECT 38.980 51.800 39.330 52.400 ;
        RECT 38.980 51.600 42.930 51.800 ;
        RECT 38.980 51.000 39.330 51.600 ;
        RECT 38.980 50.800 42.930 51.000 ;
        RECT 38.980 50.400 39.330 50.800 ;
        RECT 35.780 42.000 35.980 49.600 ;
        RECT 36.580 42.000 36.780 49.600 ;
        RECT 37.380 42.000 37.580 49.600 ;
        RECT 38.180 42.000 38.380 49.600 ;
        RECT 38.980 49.200 39.330 49.600 ;
        RECT 38.980 49.000 42.930 49.200 ;
        RECT 38.980 48.400 39.330 49.000 ;
        RECT 38.980 48.200 42.930 48.400 ;
        RECT 38.980 47.600 39.330 48.200 ;
        RECT 38.980 47.400 42.930 47.600 ;
        RECT 38.980 46.800 39.330 47.400 ;
        RECT 38.980 46.600 42.930 46.800 ;
        RECT 43.930 46.750 44.330 53.250 ;
        RECT 45.130 46.750 45.530 53.250 ;
        RECT 46.530 53.200 50.480 53.400 ;
        RECT 50.130 52.600 50.480 53.200 ;
        RECT 46.530 52.400 50.480 52.600 ;
        RECT 50.130 51.800 50.480 52.400 ;
        RECT 46.530 51.600 50.480 51.800 ;
        RECT 50.130 51.000 50.480 51.600 ;
        RECT 46.530 50.800 50.480 51.000 ;
        RECT 50.130 50.400 50.480 50.800 ;
        RECT 51.080 50.400 51.280 58.000 ;
        RECT 51.880 50.400 52.080 58.000 ;
        RECT 52.680 50.400 52.880 58.000 ;
        RECT 53.480 50.400 53.680 58.000 ;
        RECT 50.130 49.200 50.480 49.600 ;
        RECT 46.530 49.000 50.480 49.200 ;
        RECT 50.130 48.400 50.480 49.000 ;
        RECT 46.530 48.200 50.480 48.400 ;
        RECT 50.130 47.600 50.480 48.200 ;
        RECT 46.530 47.400 50.480 47.600 ;
        RECT 50.130 46.800 50.480 47.400 ;
        RECT 38.980 46.000 39.330 46.600 ;
        RECT 38.980 45.800 42.930 46.000 ;
        RECT 38.980 45.200 39.330 45.800 ;
        RECT 38.980 45.000 42.930 45.200 ;
        RECT 38.980 44.400 39.330 45.000 ;
        RECT 43.880 44.450 45.580 46.750 ;
        RECT 46.530 46.600 50.480 46.800 ;
        RECT 50.130 46.000 50.480 46.600 ;
        RECT 46.530 45.800 50.480 46.000 ;
        RECT 50.130 45.200 50.480 45.800 ;
        RECT 46.530 45.000 50.480 45.200 ;
        RECT 38.980 44.200 42.930 44.400 ;
        RECT 38.980 43.600 39.330 44.200 ;
        RECT 38.980 43.400 42.930 43.600 ;
        RECT 38.980 42.800 39.330 43.400 ;
        RECT 38.980 42.600 42.930 42.800 ;
        RECT 38.980 42.000 39.330 42.600 ;
        RECT 26.530 41.400 42.930 42.000 ;
        RECT 29.180 40.800 31.480 40.850 ;
        RECT 37.980 40.800 40.280 40.850 ;
        RECT 43.930 40.800 44.330 44.450 ;
        RECT 25.130 40.400 44.330 40.800 ;
        RECT 45.130 40.800 45.530 44.450 ;
        RECT 50.130 44.400 50.480 45.000 ;
        RECT 46.530 44.200 50.480 44.400 ;
        RECT 50.130 43.600 50.480 44.200 ;
        RECT 46.530 43.400 50.480 43.600 ;
        RECT 50.130 42.800 50.480 43.400 ;
        RECT 46.530 42.600 50.480 42.800 ;
        RECT 50.130 42.000 50.480 42.600 ;
        RECT 51.080 42.000 51.280 49.600 ;
        RECT 51.880 42.000 52.080 49.600 ;
        RECT 52.680 42.000 52.880 49.600 ;
        RECT 53.480 42.000 53.680 49.600 ;
        RECT 54.280 42.000 55.180 58.000 ;
        RECT 55.780 50.400 55.980 58.000 ;
        RECT 56.580 50.400 56.780 58.000 ;
        RECT 57.380 50.400 57.580 58.000 ;
        RECT 58.180 50.400 58.380 58.000 ;
        RECT 58.980 57.400 59.330 58.000 ;
        RECT 58.980 57.200 62.930 57.400 ;
        RECT 58.980 56.600 59.330 57.200 ;
        RECT 58.980 56.400 62.930 56.600 ;
        RECT 58.980 55.800 59.330 56.400 ;
        RECT 58.980 55.600 62.930 55.800 ;
        RECT 58.980 55.000 59.330 55.600 ;
        RECT 63.930 55.550 64.330 59.200 ;
        RECT 65.130 59.200 84.330 59.600 ;
        RECT 65.130 55.550 65.530 59.200 ;
        RECT 69.180 59.150 71.480 59.200 ;
        RECT 77.980 59.150 80.280 59.200 ;
        RECT 66.530 58.000 82.930 58.600 ;
        RECT 70.130 57.400 70.480 58.000 ;
        RECT 66.530 57.200 70.480 57.400 ;
        RECT 70.130 56.600 70.480 57.200 ;
        RECT 66.530 56.400 70.480 56.600 ;
        RECT 70.130 55.800 70.480 56.400 ;
        RECT 66.530 55.600 70.480 55.800 ;
        RECT 58.980 54.800 62.930 55.000 ;
        RECT 58.980 54.200 59.330 54.800 ;
        RECT 58.980 54.000 62.930 54.200 ;
        RECT 58.980 53.400 59.330 54.000 ;
        RECT 58.980 53.200 62.930 53.400 ;
        RECT 63.880 53.250 65.580 55.550 ;
        RECT 70.130 55.000 70.480 55.600 ;
        RECT 66.530 54.800 70.480 55.000 ;
        RECT 70.130 54.200 70.480 54.800 ;
        RECT 66.530 54.000 70.480 54.200 ;
        RECT 70.130 53.400 70.480 54.000 ;
        RECT 58.980 52.600 59.330 53.200 ;
        RECT 58.980 52.400 62.930 52.600 ;
        RECT 58.980 51.800 59.330 52.400 ;
        RECT 58.980 51.600 62.930 51.800 ;
        RECT 58.980 51.000 59.330 51.600 ;
        RECT 58.980 50.800 62.930 51.000 ;
        RECT 58.980 50.400 59.330 50.800 ;
        RECT 55.780 42.000 55.980 49.600 ;
        RECT 56.580 42.000 56.780 49.600 ;
        RECT 57.380 42.000 57.580 49.600 ;
        RECT 58.180 42.000 58.380 49.600 ;
        RECT 58.980 49.200 59.330 49.600 ;
        RECT 58.980 49.000 62.930 49.200 ;
        RECT 58.980 48.400 59.330 49.000 ;
        RECT 58.980 48.200 62.930 48.400 ;
        RECT 58.980 47.600 59.330 48.200 ;
        RECT 58.980 47.400 62.930 47.600 ;
        RECT 58.980 46.800 59.330 47.400 ;
        RECT 58.980 46.600 62.930 46.800 ;
        RECT 63.930 46.750 64.330 53.250 ;
        RECT 65.130 46.750 65.530 53.250 ;
        RECT 66.530 53.200 70.480 53.400 ;
        RECT 70.130 52.600 70.480 53.200 ;
        RECT 66.530 52.400 70.480 52.600 ;
        RECT 70.130 51.800 70.480 52.400 ;
        RECT 66.530 51.600 70.480 51.800 ;
        RECT 70.130 51.000 70.480 51.600 ;
        RECT 66.530 50.800 70.480 51.000 ;
        RECT 70.130 50.400 70.480 50.800 ;
        RECT 71.080 50.400 71.280 58.000 ;
        RECT 71.880 50.400 72.080 58.000 ;
        RECT 72.680 50.400 72.880 58.000 ;
        RECT 73.480 50.400 73.680 58.000 ;
        RECT 70.130 49.200 70.480 49.600 ;
        RECT 66.530 49.000 70.480 49.200 ;
        RECT 70.130 48.400 70.480 49.000 ;
        RECT 66.530 48.200 70.480 48.400 ;
        RECT 70.130 47.600 70.480 48.200 ;
        RECT 66.530 47.400 70.480 47.600 ;
        RECT 70.130 46.800 70.480 47.400 ;
        RECT 58.980 46.000 59.330 46.600 ;
        RECT 58.980 45.800 62.930 46.000 ;
        RECT 58.980 45.200 59.330 45.800 ;
        RECT 58.980 45.000 62.930 45.200 ;
        RECT 58.980 44.400 59.330 45.000 ;
        RECT 63.880 44.450 65.580 46.750 ;
        RECT 66.530 46.600 70.480 46.800 ;
        RECT 70.130 46.000 70.480 46.600 ;
        RECT 66.530 45.800 70.480 46.000 ;
        RECT 70.130 45.200 70.480 45.800 ;
        RECT 66.530 45.000 70.480 45.200 ;
        RECT 58.980 44.200 62.930 44.400 ;
        RECT 58.980 43.600 59.330 44.200 ;
        RECT 58.980 43.400 62.930 43.600 ;
        RECT 58.980 42.800 59.330 43.400 ;
        RECT 58.980 42.600 62.930 42.800 ;
        RECT 58.980 42.000 59.330 42.600 ;
        RECT 46.530 41.400 62.930 42.000 ;
        RECT 49.180 40.800 51.480 40.850 ;
        RECT 57.980 40.800 60.280 40.850 ;
        RECT 63.930 40.800 64.330 44.450 ;
        RECT 45.130 40.400 64.330 40.800 ;
        RECT 65.130 40.800 65.530 44.450 ;
        RECT 70.130 44.400 70.480 45.000 ;
        RECT 66.530 44.200 70.480 44.400 ;
        RECT 70.130 43.600 70.480 44.200 ;
        RECT 66.530 43.400 70.480 43.600 ;
        RECT 70.130 42.800 70.480 43.400 ;
        RECT 66.530 42.600 70.480 42.800 ;
        RECT 70.130 42.000 70.480 42.600 ;
        RECT 71.080 42.000 71.280 49.600 ;
        RECT 71.880 42.000 72.080 49.600 ;
        RECT 72.680 42.000 72.880 49.600 ;
        RECT 73.480 42.000 73.680 49.600 ;
        RECT 74.280 42.000 75.180 58.000 ;
        RECT 75.780 50.400 75.980 58.000 ;
        RECT 76.580 50.400 76.780 58.000 ;
        RECT 77.380 50.400 77.580 58.000 ;
        RECT 78.180 50.400 78.380 58.000 ;
        RECT 78.980 57.400 79.330 58.000 ;
        RECT 78.980 57.200 82.930 57.400 ;
        RECT 78.980 56.600 79.330 57.200 ;
        RECT 78.980 56.400 82.930 56.600 ;
        RECT 78.980 55.800 79.330 56.400 ;
        RECT 78.980 55.600 82.930 55.800 ;
        RECT 78.980 55.000 79.330 55.600 ;
        RECT 83.930 55.550 84.330 59.200 ;
        RECT 85.130 59.200 104.330 59.600 ;
        RECT 85.130 55.550 85.530 59.200 ;
        RECT 89.180 59.150 91.480 59.200 ;
        RECT 97.980 59.150 100.280 59.200 ;
        RECT 86.530 58.000 102.930 58.600 ;
        RECT 90.130 57.400 90.480 58.000 ;
        RECT 86.530 57.200 90.480 57.400 ;
        RECT 90.130 56.600 90.480 57.200 ;
        RECT 86.530 56.400 90.480 56.600 ;
        RECT 90.130 55.800 90.480 56.400 ;
        RECT 86.530 55.600 90.480 55.800 ;
        RECT 78.980 54.800 82.930 55.000 ;
        RECT 78.980 54.200 79.330 54.800 ;
        RECT 78.980 54.000 82.930 54.200 ;
        RECT 78.980 53.400 79.330 54.000 ;
        RECT 78.980 53.200 82.930 53.400 ;
        RECT 83.880 53.250 85.580 55.550 ;
        RECT 90.130 55.000 90.480 55.600 ;
        RECT 86.530 54.800 90.480 55.000 ;
        RECT 90.130 54.200 90.480 54.800 ;
        RECT 86.530 54.000 90.480 54.200 ;
        RECT 90.130 53.400 90.480 54.000 ;
        RECT 78.980 52.600 79.330 53.200 ;
        RECT 78.980 52.400 82.930 52.600 ;
        RECT 78.980 51.800 79.330 52.400 ;
        RECT 78.980 51.600 82.930 51.800 ;
        RECT 78.980 51.000 79.330 51.600 ;
        RECT 78.980 50.800 82.930 51.000 ;
        RECT 78.980 50.400 79.330 50.800 ;
        RECT 75.780 42.000 75.980 49.600 ;
        RECT 76.580 42.000 76.780 49.600 ;
        RECT 77.380 42.000 77.580 49.600 ;
        RECT 78.180 42.000 78.380 49.600 ;
        RECT 78.980 49.200 79.330 49.600 ;
        RECT 78.980 49.000 82.930 49.200 ;
        RECT 78.980 48.400 79.330 49.000 ;
        RECT 78.980 48.200 82.930 48.400 ;
        RECT 78.980 47.600 79.330 48.200 ;
        RECT 78.980 47.400 82.930 47.600 ;
        RECT 78.980 46.800 79.330 47.400 ;
        RECT 78.980 46.600 82.930 46.800 ;
        RECT 83.930 46.750 84.330 53.250 ;
        RECT 85.130 46.750 85.530 53.250 ;
        RECT 86.530 53.200 90.480 53.400 ;
        RECT 90.130 52.600 90.480 53.200 ;
        RECT 86.530 52.400 90.480 52.600 ;
        RECT 90.130 51.800 90.480 52.400 ;
        RECT 86.530 51.600 90.480 51.800 ;
        RECT 90.130 51.000 90.480 51.600 ;
        RECT 86.530 50.800 90.480 51.000 ;
        RECT 90.130 50.400 90.480 50.800 ;
        RECT 91.080 50.400 91.280 58.000 ;
        RECT 91.880 50.400 92.080 58.000 ;
        RECT 92.680 50.400 92.880 58.000 ;
        RECT 93.480 50.400 93.680 58.000 ;
        RECT 90.130 49.200 90.480 49.600 ;
        RECT 86.530 49.000 90.480 49.200 ;
        RECT 90.130 48.400 90.480 49.000 ;
        RECT 86.530 48.200 90.480 48.400 ;
        RECT 90.130 47.600 90.480 48.200 ;
        RECT 86.530 47.400 90.480 47.600 ;
        RECT 90.130 46.800 90.480 47.400 ;
        RECT 78.980 46.000 79.330 46.600 ;
        RECT 78.980 45.800 82.930 46.000 ;
        RECT 78.980 45.200 79.330 45.800 ;
        RECT 78.980 45.000 82.930 45.200 ;
        RECT 78.980 44.400 79.330 45.000 ;
        RECT 83.880 44.450 85.580 46.750 ;
        RECT 86.530 46.600 90.480 46.800 ;
        RECT 90.130 46.000 90.480 46.600 ;
        RECT 86.530 45.800 90.480 46.000 ;
        RECT 90.130 45.200 90.480 45.800 ;
        RECT 86.530 45.000 90.480 45.200 ;
        RECT 78.980 44.200 82.930 44.400 ;
        RECT 78.980 43.600 79.330 44.200 ;
        RECT 78.980 43.400 82.930 43.600 ;
        RECT 78.980 42.800 79.330 43.400 ;
        RECT 78.980 42.600 82.930 42.800 ;
        RECT 78.980 42.000 79.330 42.600 ;
        RECT 66.530 41.400 82.930 42.000 ;
        RECT 69.180 40.800 71.480 40.850 ;
        RECT 77.980 40.800 80.280 40.850 ;
        RECT 83.930 40.800 84.330 44.450 ;
        RECT 65.130 40.400 84.330 40.800 ;
        RECT 85.130 40.800 85.530 44.450 ;
        RECT 90.130 44.400 90.480 45.000 ;
        RECT 86.530 44.200 90.480 44.400 ;
        RECT 90.130 43.600 90.480 44.200 ;
        RECT 86.530 43.400 90.480 43.600 ;
        RECT 90.130 42.800 90.480 43.400 ;
        RECT 86.530 42.600 90.480 42.800 ;
        RECT 90.130 42.000 90.480 42.600 ;
        RECT 91.080 42.000 91.280 49.600 ;
        RECT 91.880 42.000 92.080 49.600 ;
        RECT 92.680 42.000 92.880 49.600 ;
        RECT 93.480 42.000 93.680 49.600 ;
        RECT 94.280 42.000 95.180 58.000 ;
        RECT 95.780 50.400 95.980 58.000 ;
        RECT 96.580 50.400 96.780 58.000 ;
        RECT 97.380 50.400 97.580 58.000 ;
        RECT 98.180 50.400 98.380 58.000 ;
        RECT 98.980 57.400 99.330 58.000 ;
        RECT 98.980 57.200 102.930 57.400 ;
        RECT 98.980 56.600 99.330 57.200 ;
        RECT 98.980 56.400 102.930 56.600 ;
        RECT 98.980 55.800 99.330 56.400 ;
        RECT 98.980 55.600 102.930 55.800 ;
        RECT 98.980 55.000 99.330 55.600 ;
        RECT 103.930 55.550 104.330 59.200 ;
        RECT 105.340 56.805 105.700 57.185 ;
        RECT 105.970 56.805 106.330 57.185 ;
        RECT 106.570 56.805 106.930 57.185 ;
        RECT 105.340 56.215 105.700 56.595 ;
        RECT 105.970 56.215 106.330 56.595 ;
        RECT 106.570 56.215 106.930 56.595 ;
        RECT 98.980 54.800 102.930 55.000 ;
        RECT 98.980 54.200 99.330 54.800 ;
        RECT 98.980 54.000 102.930 54.200 ;
        RECT 98.980 53.400 99.330 54.000 ;
        RECT 98.980 53.200 102.930 53.400 ;
        RECT 103.880 53.250 104.730 55.550 ;
        RECT 98.980 52.600 99.330 53.200 ;
        RECT 98.980 52.400 102.930 52.600 ;
        RECT 98.980 51.800 99.330 52.400 ;
        RECT 98.980 51.600 102.930 51.800 ;
        RECT 98.980 51.000 99.330 51.600 ;
        RECT 98.980 50.800 102.930 51.000 ;
        RECT 98.980 50.400 99.330 50.800 ;
        RECT 95.780 42.000 95.980 49.600 ;
        RECT 96.580 42.000 96.780 49.600 ;
        RECT 97.380 42.000 97.580 49.600 ;
        RECT 98.180 42.000 98.380 49.600 ;
        RECT 98.980 49.200 99.330 49.600 ;
        RECT 98.980 49.000 102.930 49.200 ;
        RECT 98.980 48.400 99.330 49.000 ;
        RECT 98.980 48.200 102.930 48.400 ;
        RECT 98.980 47.600 99.330 48.200 ;
        RECT 98.980 47.400 102.930 47.600 ;
        RECT 98.980 46.800 99.330 47.400 ;
        RECT 98.980 46.600 102.930 46.800 ;
        RECT 103.930 46.750 104.330 53.250 ;
        RECT 98.980 46.000 99.330 46.600 ;
        RECT 98.980 45.800 102.930 46.000 ;
        RECT 98.980 45.200 99.330 45.800 ;
        RECT 98.980 45.000 102.930 45.200 ;
        RECT 98.980 44.400 99.330 45.000 ;
        RECT 103.880 44.450 104.730 46.750 ;
        RECT 98.980 44.200 102.930 44.400 ;
        RECT 98.980 43.600 99.330 44.200 ;
        RECT 98.980 43.400 102.930 43.600 ;
        RECT 98.980 42.800 99.330 43.400 ;
        RECT 98.980 42.600 102.930 42.800 ;
        RECT 98.980 42.000 99.330 42.600 ;
        RECT 86.530 41.400 102.930 42.000 ;
        RECT 89.180 40.800 91.480 40.850 ;
        RECT 97.980 40.800 100.280 40.850 ;
        RECT 103.930 40.800 104.330 44.450 ;
        RECT 105.340 42.590 105.700 42.970 ;
        RECT 105.970 42.590 106.330 42.970 ;
        RECT 106.570 42.590 106.930 42.970 ;
        RECT 105.340 42.000 105.700 42.380 ;
        RECT 105.970 42.000 106.330 42.380 ;
        RECT 106.570 42.000 106.930 42.380 ;
        RECT 85.130 40.400 104.330 40.800 ;
        RECT 9.180 39.600 11.480 40.400 ;
        RECT 17.980 39.600 20.280 40.400 ;
        RECT 29.180 39.600 31.480 40.400 ;
        RECT 37.980 39.600 40.280 40.400 ;
        RECT 49.180 39.600 51.480 40.400 ;
        RECT 57.980 39.600 60.280 40.400 ;
        RECT 69.180 39.600 71.480 40.400 ;
        RECT 77.980 39.600 80.280 40.400 ;
        RECT 89.180 39.600 91.480 40.400 ;
        RECT 97.980 39.600 100.280 40.400 ;
        RECT 5.130 39.200 24.330 39.600 ;
        RECT 2.515 37.260 2.875 37.640 ;
        RECT 3.145 37.260 3.505 37.640 ;
        RECT 3.745 37.260 4.105 37.640 ;
        RECT 2.515 36.670 2.875 37.050 ;
        RECT 3.145 36.670 3.505 37.050 ;
        RECT 3.745 36.670 4.105 37.050 ;
        RECT 5.130 35.550 5.530 39.200 ;
        RECT 9.180 39.150 11.480 39.200 ;
        RECT 17.980 39.150 20.280 39.200 ;
        RECT 6.530 38.000 22.930 38.600 ;
        RECT 10.130 37.400 10.480 38.000 ;
        RECT 6.530 37.200 10.480 37.400 ;
        RECT 10.130 36.600 10.480 37.200 ;
        RECT 6.530 36.400 10.480 36.600 ;
        RECT 10.130 35.800 10.480 36.400 ;
        RECT 6.530 35.600 10.480 35.800 ;
        RECT 2.315 33.255 5.580 35.550 ;
        RECT 10.130 35.000 10.480 35.600 ;
        RECT 6.530 34.800 10.480 35.000 ;
        RECT 10.130 34.200 10.480 34.800 ;
        RECT 6.530 34.000 10.480 34.200 ;
        RECT 10.130 33.400 10.480 34.000 ;
        RECT 4.730 33.250 5.580 33.255 ;
        RECT 5.130 26.750 5.530 33.250 ;
        RECT 6.530 33.200 10.480 33.400 ;
        RECT 10.130 32.600 10.480 33.200 ;
        RECT 6.530 32.400 10.480 32.600 ;
        RECT 10.130 31.800 10.480 32.400 ;
        RECT 6.530 31.600 10.480 31.800 ;
        RECT 10.130 31.000 10.480 31.600 ;
        RECT 6.530 30.800 10.480 31.000 ;
        RECT 10.130 30.400 10.480 30.800 ;
        RECT 11.080 30.400 11.280 38.000 ;
        RECT 11.880 30.400 12.080 38.000 ;
        RECT 12.680 30.400 12.880 38.000 ;
        RECT 13.480 30.400 13.680 38.000 ;
        RECT 10.130 29.200 10.480 29.600 ;
        RECT 6.530 29.000 10.480 29.200 ;
        RECT 10.130 28.400 10.480 29.000 ;
        RECT 6.530 28.200 10.480 28.400 ;
        RECT 10.130 27.600 10.480 28.200 ;
        RECT 6.530 27.400 10.480 27.600 ;
        RECT 10.130 26.800 10.480 27.400 ;
        RECT 4.730 26.745 5.580 26.750 ;
        RECT 2.315 24.450 5.580 26.745 ;
        RECT 6.530 26.600 10.480 26.800 ;
        RECT 10.130 26.000 10.480 26.600 ;
        RECT 6.530 25.800 10.480 26.000 ;
        RECT 10.130 25.200 10.480 25.800 ;
        RECT 6.530 25.000 10.480 25.200 ;
        RECT 2.515 23.145 2.875 23.525 ;
        RECT 3.145 23.145 3.505 23.525 ;
        RECT 3.745 23.145 4.105 23.525 ;
        RECT 2.515 22.555 2.875 22.935 ;
        RECT 3.145 22.555 3.505 22.935 ;
        RECT 3.745 22.555 4.105 22.935 ;
        RECT 5.130 20.800 5.530 24.450 ;
        RECT 10.130 24.400 10.480 25.000 ;
        RECT 6.530 24.200 10.480 24.400 ;
        RECT 10.130 23.600 10.480 24.200 ;
        RECT 6.530 23.400 10.480 23.600 ;
        RECT 10.130 22.800 10.480 23.400 ;
        RECT 6.530 22.600 10.480 22.800 ;
        RECT 10.130 22.000 10.480 22.600 ;
        RECT 11.080 22.000 11.280 29.600 ;
        RECT 11.880 22.000 12.080 29.600 ;
        RECT 12.680 22.000 12.880 29.600 ;
        RECT 13.480 22.000 13.680 29.600 ;
        RECT 14.280 22.000 15.180 38.000 ;
        RECT 15.780 30.400 15.980 38.000 ;
        RECT 16.580 30.400 16.780 38.000 ;
        RECT 17.380 30.400 17.580 38.000 ;
        RECT 18.180 30.400 18.380 38.000 ;
        RECT 18.980 37.400 19.330 38.000 ;
        RECT 18.980 37.200 22.930 37.400 ;
        RECT 18.980 36.600 19.330 37.200 ;
        RECT 18.980 36.400 22.930 36.600 ;
        RECT 18.980 35.800 19.330 36.400 ;
        RECT 18.980 35.600 22.930 35.800 ;
        RECT 18.980 35.000 19.330 35.600 ;
        RECT 23.930 35.550 24.330 39.200 ;
        RECT 25.130 39.200 44.330 39.600 ;
        RECT 25.130 35.550 25.530 39.200 ;
        RECT 29.180 39.150 31.480 39.200 ;
        RECT 37.980 39.150 40.280 39.200 ;
        RECT 26.530 38.000 42.930 38.600 ;
        RECT 30.130 37.400 30.480 38.000 ;
        RECT 26.530 37.200 30.480 37.400 ;
        RECT 30.130 36.600 30.480 37.200 ;
        RECT 26.530 36.400 30.480 36.600 ;
        RECT 30.130 35.800 30.480 36.400 ;
        RECT 26.530 35.600 30.480 35.800 ;
        RECT 18.980 34.800 22.930 35.000 ;
        RECT 18.980 34.200 19.330 34.800 ;
        RECT 18.980 34.000 22.930 34.200 ;
        RECT 18.980 33.400 19.330 34.000 ;
        RECT 18.980 33.200 22.930 33.400 ;
        RECT 23.880 33.250 25.580 35.550 ;
        RECT 30.130 35.000 30.480 35.600 ;
        RECT 26.530 34.800 30.480 35.000 ;
        RECT 30.130 34.200 30.480 34.800 ;
        RECT 26.530 34.000 30.480 34.200 ;
        RECT 30.130 33.400 30.480 34.000 ;
        RECT 18.980 32.600 19.330 33.200 ;
        RECT 18.980 32.400 22.930 32.600 ;
        RECT 18.980 31.800 19.330 32.400 ;
        RECT 18.980 31.600 22.930 31.800 ;
        RECT 18.980 31.000 19.330 31.600 ;
        RECT 18.980 30.800 22.930 31.000 ;
        RECT 18.980 30.400 19.330 30.800 ;
        RECT 15.780 22.000 15.980 29.600 ;
        RECT 16.580 22.000 16.780 29.600 ;
        RECT 17.380 22.000 17.580 29.600 ;
        RECT 18.180 22.000 18.380 29.600 ;
        RECT 18.980 29.200 19.330 29.600 ;
        RECT 18.980 29.000 22.930 29.200 ;
        RECT 18.980 28.400 19.330 29.000 ;
        RECT 18.980 28.200 22.930 28.400 ;
        RECT 18.980 27.600 19.330 28.200 ;
        RECT 18.980 27.400 22.930 27.600 ;
        RECT 18.980 26.800 19.330 27.400 ;
        RECT 18.980 26.600 22.930 26.800 ;
        RECT 23.930 26.750 24.330 33.250 ;
        RECT 25.130 26.750 25.530 33.250 ;
        RECT 26.530 33.200 30.480 33.400 ;
        RECT 30.130 32.600 30.480 33.200 ;
        RECT 26.530 32.400 30.480 32.600 ;
        RECT 30.130 31.800 30.480 32.400 ;
        RECT 26.530 31.600 30.480 31.800 ;
        RECT 30.130 31.000 30.480 31.600 ;
        RECT 26.530 30.800 30.480 31.000 ;
        RECT 30.130 30.400 30.480 30.800 ;
        RECT 31.080 30.400 31.280 38.000 ;
        RECT 31.880 30.400 32.080 38.000 ;
        RECT 32.680 30.400 32.880 38.000 ;
        RECT 33.480 30.400 33.680 38.000 ;
        RECT 30.130 29.200 30.480 29.600 ;
        RECT 26.530 29.000 30.480 29.200 ;
        RECT 30.130 28.400 30.480 29.000 ;
        RECT 26.530 28.200 30.480 28.400 ;
        RECT 30.130 27.600 30.480 28.200 ;
        RECT 26.530 27.400 30.480 27.600 ;
        RECT 30.130 26.800 30.480 27.400 ;
        RECT 18.980 26.000 19.330 26.600 ;
        RECT 18.980 25.800 22.930 26.000 ;
        RECT 18.980 25.200 19.330 25.800 ;
        RECT 18.980 25.000 22.930 25.200 ;
        RECT 18.980 24.400 19.330 25.000 ;
        RECT 23.880 24.450 25.580 26.750 ;
        RECT 26.530 26.600 30.480 26.800 ;
        RECT 30.130 26.000 30.480 26.600 ;
        RECT 26.530 25.800 30.480 26.000 ;
        RECT 30.130 25.200 30.480 25.800 ;
        RECT 26.530 25.000 30.480 25.200 ;
        RECT 18.980 24.200 22.930 24.400 ;
        RECT 18.980 23.600 19.330 24.200 ;
        RECT 18.980 23.400 22.930 23.600 ;
        RECT 18.980 22.800 19.330 23.400 ;
        RECT 18.980 22.600 22.930 22.800 ;
        RECT 18.980 22.000 19.330 22.600 ;
        RECT 6.530 21.400 22.930 22.000 ;
        RECT 9.180 20.800 11.480 20.850 ;
        RECT 17.980 20.800 20.280 20.850 ;
        RECT 23.930 20.800 24.330 24.450 ;
        RECT 5.130 20.400 24.330 20.800 ;
        RECT 25.130 20.800 25.530 24.450 ;
        RECT 30.130 24.400 30.480 25.000 ;
        RECT 26.530 24.200 30.480 24.400 ;
        RECT 30.130 23.600 30.480 24.200 ;
        RECT 26.530 23.400 30.480 23.600 ;
        RECT 30.130 22.800 30.480 23.400 ;
        RECT 26.530 22.600 30.480 22.800 ;
        RECT 30.130 22.000 30.480 22.600 ;
        RECT 31.080 22.000 31.280 29.600 ;
        RECT 31.880 22.000 32.080 29.600 ;
        RECT 32.680 22.000 32.880 29.600 ;
        RECT 33.480 22.000 33.680 29.600 ;
        RECT 34.280 22.000 35.180 38.000 ;
        RECT 35.780 30.400 35.980 38.000 ;
        RECT 36.580 30.400 36.780 38.000 ;
        RECT 37.380 30.400 37.580 38.000 ;
        RECT 38.180 30.400 38.380 38.000 ;
        RECT 38.980 37.400 39.330 38.000 ;
        RECT 38.980 37.200 42.930 37.400 ;
        RECT 38.980 36.600 39.330 37.200 ;
        RECT 38.980 36.400 42.930 36.600 ;
        RECT 38.980 35.800 39.330 36.400 ;
        RECT 38.980 35.600 42.930 35.800 ;
        RECT 38.980 35.000 39.330 35.600 ;
        RECT 43.930 35.550 44.330 39.200 ;
        RECT 45.130 39.200 64.330 39.600 ;
        RECT 45.130 35.550 45.530 39.200 ;
        RECT 49.180 39.150 51.480 39.200 ;
        RECT 57.980 39.150 60.280 39.200 ;
        RECT 46.530 38.000 62.930 38.600 ;
        RECT 50.130 37.400 50.480 38.000 ;
        RECT 46.530 37.200 50.480 37.400 ;
        RECT 50.130 36.600 50.480 37.200 ;
        RECT 46.530 36.400 50.480 36.600 ;
        RECT 50.130 35.800 50.480 36.400 ;
        RECT 46.530 35.600 50.480 35.800 ;
        RECT 38.980 34.800 42.930 35.000 ;
        RECT 38.980 34.200 39.330 34.800 ;
        RECT 38.980 34.000 42.930 34.200 ;
        RECT 38.980 33.400 39.330 34.000 ;
        RECT 38.980 33.200 42.930 33.400 ;
        RECT 43.880 33.250 45.580 35.550 ;
        RECT 50.130 35.000 50.480 35.600 ;
        RECT 46.530 34.800 50.480 35.000 ;
        RECT 50.130 34.200 50.480 34.800 ;
        RECT 46.530 34.000 50.480 34.200 ;
        RECT 50.130 33.400 50.480 34.000 ;
        RECT 38.980 32.600 39.330 33.200 ;
        RECT 38.980 32.400 42.930 32.600 ;
        RECT 38.980 31.800 39.330 32.400 ;
        RECT 38.980 31.600 42.930 31.800 ;
        RECT 38.980 31.000 39.330 31.600 ;
        RECT 38.980 30.800 42.930 31.000 ;
        RECT 38.980 30.400 39.330 30.800 ;
        RECT 35.780 22.000 35.980 29.600 ;
        RECT 36.580 22.000 36.780 29.600 ;
        RECT 37.380 22.000 37.580 29.600 ;
        RECT 38.180 22.000 38.380 29.600 ;
        RECT 38.980 29.200 39.330 29.600 ;
        RECT 38.980 29.000 42.930 29.200 ;
        RECT 38.980 28.400 39.330 29.000 ;
        RECT 38.980 28.200 42.930 28.400 ;
        RECT 38.980 27.600 39.330 28.200 ;
        RECT 38.980 27.400 42.930 27.600 ;
        RECT 38.980 26.800 39.330 27.400 ;
        RECT 38.980 26.600 42.930 26.800 ;
        RECT 43.930 26.750 44.330 33.250 ;
        RECT 45.130 26.750 45.530 33.250 ;
        RECT 46.530 33.200 50.480 33.400 ;
        RECT 50.130 32.600 50.480 33.200 ;
        RECT 46.530 32.400 50.480 32.600 ;
        RECT 50.130 31.800 50.480 32.400 ;
        RECT 46.530 31.600 50.480 31.800 ;
        RECT 50.130 31.000 50.480 31.600 ;
        RECT 46.530 30.800 50.480 31.000 ;
        RECT 50.130 30.400 50.480 30.800 ;
        RECT 51.080 30.400 51.280 38.000 ;
        RECT 51.880 30.400 52.080 38.000 ;
        RECT 52.680 30.400 52.880 38.000 ;
        RECT 53.480 30.400 53.680 38.000 ;
        RECT 50.130 29.200 50.480 29.600 ;
        RECT 46.530 29.000 50.480 29.200 ;
        RECT 50.130 28.400 50.480 29.000 ;
        RECT 46.530 28.200 50.480 28.400 ;
        RECT 50.130 27.600 50.480 28.200 ;
        RECT 46.530 27.400 50.480 27.600 ;
        RECT 50.130 26.800 50.480 27.400 ;
        RECT 38.980 26.000 39.330 26.600 ;
        RECT 38.980 25.800 42.930 26.000 ;
        RECT 38.980 25.200 39.330 25.800 ;
        RECT 38.980 25.000 42.930 25.200 ;
        RECT 38.980 24.400 39.330 25.000 ;
        RECT 43.880 24.450 45.580 26.750 ;
        RECT 46.530 26.600 50.480 26.800 ;
        RECT 50.130 26.000 50.480 26.600 ;
        RECT 46.530 25.800 50.480 26.000 ;
        RECT 50.130 25.200 50.480 25.800 ;
        RECT 46.530 25.000 50.480 25.200 ;
        RECT 38.980 24.200 42.930 24.400 ;
        RECT 38.980 23.600 39.330 24.200 ;
        RECT 38.980 23.400 42.930 23.600 ;
        RECT 38.980 22.800 39.330 23.400 ;
        RECT 38.980 22.600 42.930 22.800 ;
        RECT 38.980 22.000 39.330 22.600 ;
        RECT 26.530 21.400 42.930 22.000 ;
        RECT 29.180 20.800 31.480 20.850 ;
        RECT 37.980 20.800 40.280 20.850 ;
        RECT 43.930 20.800 44.330 24.450 ;
        RECT 25.130 20.400 44.330 20.800 ;
        RECT 45.130 20.800 45.530 24.450 ;
        RECT 50.130 24.400 50.480 25.000 ;
        RECT 46.530 24.200 50.480 24.400 ;
        RECT 50.130 23.600 50.480 24.200 ;
        RECT 46.530 23.400 50.480 23.600 ;
        RECT 50.130 22.800 50.480 23.400 ;
        RECT 46.530 22.600 50.480 22.800 ;
        RECT 50.130 22.000 50.480 22.600 ;
        RECT 51.080 22.000 51.280 29.600 ;
        RECT 51.880 22.000 52.080 29.600 ;
        RECT 52.680 22.000 52.880 29.600 ;
        RECT 53.480 22.000 53.680 29.600 ;
        RECT 54.280 22.000 55.180 38.000 ;
        RECT 55.780 30.400 55.980 38.000 ;
        RECT 56.580 30.400 56.780 38.000 ;
        RECT 57.380 30.400 57.580 38.000 ;
        RECT 58.180 30.400 58.380 38.000 ;
        RECT 58.980 37.400 59.330 38.000 ;
        RECT 58.980 37.200 62.930 37.400 ;
        RECT 58.980 36.600 59.330 37.200 ;
        RECT 58.980 36.400 62.930 36.600 ;
        RECT 58.980 35.800 59.330 36.400 ;
        RECT 58.980 35.600 62.930 35.800 ;
        RECT 58.980 35.000 59.330 35.600 ;
        RECT 63.930 35.550 64.330 39.200 ;
        RECT 65.130 39.200 84.330 39.600 ;
        RECT 65.130 35.550 65.530 39.200 ;
        RECT 69.180 39.150 71.480 39.200 ;
        RECT 77.980 39.150 80.280 39.200 ;
        RECT 66.530 38.000 82.930 38.600 ;
        RECT 70.130 37.400 70.480 38.000 ;
        RECT 66.530 37.200 70.480 37.400 ;
        RECT 70.130 36.600 70.480 37.200 ;
        RECT 66.530 36.400 70.480 36.600 ;
        RECT 70.130 35.800 70.480 36.400 ;
        RECT 66.530 35.600 70.480 35.800 ;
        RECT 58.980 34.800 62.930 35.000 ;
        RECT 58.980 34.200 59.330 34.800 ;
        RECT 58.980 34.000 62.930 34.200 ;
        RECT 58.980 33.400 59.330 34.000 ;
        RECT 58.980 33.200 62.930 33.400 ;
        RECT 63.880 33.250 65.580 35.550 ;
        RECT 70.130 35.000 70.480 35.600 ;
        RECT 66.530 34.800 70.480 35.000 ;
        RECT 70.130 34.200 70.480 34.800 ;
        RECT 66.530 34.000 70.480 34.200 ;
        RECT 70.130 33.400 70.480 34.000 ;
        RECT 58.980 32.600 59.330 33.200 ;
        RECT 58.980 32.400 62.930 32.600 ;
        RECT 58.980 31.800 59.330 32.400 ;
        RECT 58.980 31.600 62.930 31.800 ;
        RECT 58.980 31.000 59.330 31.600 ;
        RECT 58.980 30.800 62.930 31.000 ;
        RECT 58.980 30.400 59.330 30.800 ;
        RECT 55.780 22.000 55.980 29.600 ;
        RECT 56.580 22.000 56.780 29.600 ;
        RECT 57.380 22.000 57.580 29.600 ;
        RECT 58.180 22.000 58.380 29.600 ;
        RECT 58.980 29.200 59.330 29.600 ;
        RECT 58.980 29.000 62.930 29.200 ;
        RECT 58.980 28.400 59.330 29.000 ;
        RECT 58.980 28.200 62.930 28.400 ;
        RECT 58.980 27.600 59.330 28.200 ;
        RECT 58.980 27.400 62.930 27.600 ;
        RECT 58.980 26.800 59.330 27.400 ;
        RECT 58.980 26.600 62.930 26.800 ;
        RECT 63.930 26.750 64.330 33.250 ;
        RECT 65.130 26.750 65.530 33.250 ;
        RECT 66.530 33.200 70.480 33.400 ;
        RECT 70.130 32.600 70.480 33.200 ;
        RECT 66.530 32.400 70.480 32.600 ;
        RECT 70.130 31.800 70.480 32.400 ;
        RECT 66.530 31.600 70.480 31.800 ;
        RECT 70.130 31.000 70.480 31.600 ;
        RECT 66.530 30.800 70.480 31.000 ;
        RECT 70.130 30.400 70.480 30.800 ;
        RECT 71.080 30.400 71.280 38.000 ;
        RECT 71.880 30.400 72.080 38.000 ;
        RECT 72.680 30.400 72.880 38.000 ;
        RECT 73.480 30.400 73.680 38.000 ;
        RECT 70.130 29.200 70.480 29.600 ;
        RECT 66.530 29.000 70.480 29.200 ;
        RECT 70.130 28.400 70.480 29.000 ;
        RECT 66.530 28.200 70.480 28.400 ;
        RECT 70.130 27.600 70.480 28.200 ;
        RECT 66.530 27.400 70.480 27.600 ;
        RECT 70.130 26.800 70.480 27.400 ;
        RECT 58.980 26.000 59.330 26.600 ;
        RECT 58.980 25.800 62.930 26.000 ;
        RECT 58.980 25.200 59.330 25.800 ;
        RECT 58.980 25.000 62.930 25.200 ;
        RECT 58.980 24.400 59.330 25.000 ;
        RECT 63.880 24.450 65.580 26.750 ;
        RECT 66.530 26.600 70.480 26.800 ;
        RECT 70.130 26.000 70.480 26.600 ;
        RECT 66.530 25.800 70.480 26.000 ;
        RECT 70.130 25.200 70.480 25.800 ;
        RECT 66.530 25.000 70.480 25.200 ;
        RECT 58.980 24.200 62.930 24.400 ;
        RECT 58.980 23.600 59.330 24.200 ;
        RECT 58.980 23.400 62.930 23.600 ;
        RECT 58.980 22.800 59.330 23.400 ;
        RECT 58.980 22.600 62.930 22.800 ;
        RECT 58.980 22.000 59.330 22.600 ;
        RECT 46.530 21.400 62.930 22.000 ;
        RECT 49.180 20.800 51.480 20.850 ;
        RECT 57.980 20.800 60.280 20.850 ;
        RECT 63.930 20.800 64.330 24.450 ;
        RECT 45.130 20.400 64.330 20.800 ;
        RECT 65.130 20.800 65.530 24.450 ;
        RECT 70.130 24.400 70.480 25.000 ;
        RECT 66.530 24.200 70.480 24.400 ;
        RECT 70.130 23.600 70.480 24.200 ;
        RECT 66.530 23.400 70.480 23.600 ;
        RECT 70.130 22.800 70.480 23.400 ;
        RECT 66.530 22.600 70.480 22.800 ;
        RECT 70.130 22.000 70.480 22.600 ;
        RECT 71.080 22.000 71.280 29.600 ;
        RECT 71.880 22.000 72.080 29.600 ;
        RECT 72.680 22.000 72.880 29.600 ;
        RECT 73.480 22.000 73.680 29.600 ;
        RECT 74.280 22.000 75.180 38.000 ;
        RECT 75.780 30.400 75.980 38.000 ;
        RECT 76.580 30.400 76.780 38.000 ;
        RECT 77.380 30.400 77.580 38.000 ;
        RECT 78.180 30.400 78.380 38.000 ;
        RECT 78.980 37.400 79.330 38.000 ;
        RECT 78.980 37.200 82.930 37.400 ;
        RECT 78.980 36.600 79.330 37.200 ;
        RECT 78.980 36.400 82.930 36.600 ;
        RECT 78.980 35.800 79.330 36.400 ;
        RECT 78.980 35.600 82.930 35.800 ;
        RECT 78.980 35.000 79.330 35.600 ;
        RECT 83.930 35.550 84.330 39.200 ;
        RECT 85.130 39.200 104.330 39.600 ;
        RECT 85.130 35.550 85.530 39.200 ;
        RECT 89.180 39.150 91.480 39.200 ;
        RECT 97.980 39.150 100.280 39.200 ;
        RECT 86.530 38.000 102.930 38.600 ;
        RECT 90.130 37.400 90.480 38.000 ;
        RECT 86.530 37.200 90.480 37.400 ;
        RECT 90.130 36.600 90.480 37.200 ;
        RECT 86.530 36.400 90.480 36.600 ;
        RECT 90.130 35.800 90.480 36.400 ;
        RECT 86.530 35.600 90.480 35.800 ;
        RECT 78.980 34.800 82.930 35.000 ;
        RECT 78.980 34.200 79.330 34.800 ;
        RECT 78.980 34.000 82.930 34.200 ;
        RECT 78.980 33.400 79.330 34.000 ;
        RECT 78.980 33.200 82.930 33.400 ;
        RECT 83.880 33.250 85.580 35.550 ;
        RECT 90.130 35.000 90.480 35.600 ;
        RECT 86.530 34.800 90.480 35.000 ;
        RECT 90.130 34.200 90.480 34.800 ;
        RECT 86.530 34.000 90.480 34.200 ;
        RECT 90.130 33.400 90.480 34.000 ;
        RECT 78.980 32.600 79.330 33.200 ;
        RECT 78.980 32.400 82.930 32.600 ;
        RECT 78.980 31.800 79.330 32.400 ;
        RECT 78.980 31.600 82.930 31.800 ;
        RECT 78.980 31.000 79.330 31.600 ;
        RECT 78.980 30.800 82.930 31.000 ;
        RECT 78.980 30.400 79.330 30.800 ;
        RECT 75.780 22.000 75.980 29.600 ;
        RECT 76.580 22.000 76.780 29.600 ;
        RECT 77.380 22.000 77.580 29.600 ;
        RECT 78.180 22.000 78.380 29.600 ;
        RECT 78.980 29.200 79.330 29.600 ;
        RECT 78.980 29.000 82.930 29.200 ;
        RECT 78.980 28.400 79.330 29.000 ;
        RECT 78.980 28.200 82.930 28.400 ;
        RECT 78.980 27.600 79.330 28.200 ;
        RECT 78.980 27.400 82.930 27.600 ;
        RECT 78.980 26.800 79.330 27.400 ;
        RECT 78.980 26.600 82.930 26.800 ;
        RECT 83.930 26.750 84.330 33.250 ;
        RECT 85.130 26.750 85.530 33.250 ;
        RECT 86.530 33.200 90.480 33.400 ;
        RECT 90.130 32.600 90.480 33.200 ;
        RECT 86.530 32.400 90.480 32.600 ;
        RECT 90.130 31.800 90.480 32.400 ;
        RECT 86.530 31.600 90.480 31.800 ;
        RECT 90.130 31.000 90.480 31.600 ;
        RECT 86.530 30.800 90.480 31.000 ;
        RECT 90.130 30.400 90.480 30.800 ;
        RECT 91.080 30.400 91.280 38.000 ;
        RECT 91.880 30.400 92.080 38.000 ;
        RECT 92.680 30.400 92.880 38.000 ;
        RECT 93.480 30.400 93.680 38.000 ;
        RECT 90.130 29.200 90.480 29.600 ;
        RECT 86.530 29.000 90.480 29.200 ;
        RECT 90.130 28.400 90.480 29.000 ;
        RECT 86.530 28.200 90.480 28.400 ;
        RECT 90.130 27.600 90.480 28.200 ;
        RECT 86.530 27.400 90.480 27.600 ;
        RECT 90.130 26.800 90.480 27.400 ;
        RECT 78.980 26.000 79.330 26.600 ;
        RECT 78.980 25.800 82.930 26.000 ;
        RECT 78.980 25.200 79.330 25.800 ;
        RECT 78.980 25.000 82.930 25.200 ;
        RECT 78.980 24.400 79.330 25.000 ;
        RECT 83.880 24.450 85.580 26.750 ;
        RECT 86.530 26.600 90.480 26.800 ;
        RECT 90.130 26.000 90.480 26.600 ;
        RECT 86.530 25.800 90.480 26.000 ;
        RECT 90.130 25.200 90.480 25.800 ;
        RECT 86.530 25.000 90.480 25.200 ;
        RECT 78.980 24.200 82.930 24.400 ;
        RECT 78.980 23.600 79.330 24.200 ;
        RECT 78.980 23.400 82.930 23.600 ;
        RECT 78.980 22.800 79.330 23.400 ;
        RECT 78.980 22.600 82.930 22.800 ;
        RECT 78.980 22.000 79.330 22.600 ;
        RECT 66.530 21.400 82.930 22.000 ;
        RECT 69.180 20.800 71.480 20.850 ;
        RECT 77.980 20.800 80.280 20.850 ;
        RECT 83.930 20.800 84.330 24.450 ;
        RECT 65.130 20.400 84.330 20.800 ;
        RECT 85.130 20.800 85.530 24.450 ;
        RECT 90.130 24.400 90.480 25.000 ;
        RECT 86.530 24.200 90.480 24.400 ;
        RECT 90.130 23.600 90.480 24.200 ;
        RECT 86.530 23.400 90.480 23.600 ;
        RECT 90.130 22.800 90.480 23.400 ;
        RECT 86.530 22.600 90.480 22.800 ;
        RECT 90.130 22.000 90.480 22.600 ;
        RECT 91.080 22.000 91.280 29.600 ;
        RECT 91.880 22.000 92.080 29.600 ;
        RECT 92.680 22.000 92.880 29.600 ;
        RECT 93.480 22.000 93.680 29.600 ;
        RECT 94.280 22.000 95.180 38.000 ;
        RECT 95.780 30.400 95.980 38.000 ;
        RECT 96.580 30.400 96.780 38.000 ;
        RECT 97.380 30.400 97.580 38.000 ;
        RECT 98.180 30.400 98.380 38.000 ;
        RECT 98.980 37.400 99.330 38.000 ;
        RECT 98.980 37.200 102.930 37.400 ;
        RECT 98.980 36.600 99.330 37.200 ;
        RECT 98.980 36.400 102.930 36.600 ;
        RECT 98.980 35.800 99.330 36.400 ;
        RECT 98.980 35.600 102.930 35.800 ;
        RECT 98.980 35.000 99.330 35.600 ;
        RECT 103.930 35.550 104.330 39.200 ;
        RECT 105.340 36.805 105.700 37.185 ;
        RECT 105.970 36.805 106.330 37.185 ;
        RECT 106.570 36.805 106.930 37.185 ;
        RECT 105.340 36.215 105.700 36.595 ;
        RECT 105.970 36.215 106.330 36.595 ;
        RECT 106.570 36.215 106.930 36.595 ;
        RECT 98.980 34.800 102.930 35.000 ;
        RECT 98.980 34.200 99.330 34.800 ;
        RECT 98.980 34.000 102.930 34.200 ;
        RECT 98.980 33.400 99.330 34.000 ;
        RECT 98.980 33.200 102.930 33.400 ;
        RECT 103.880 33.250 104.730 35.550 ;
        RECT 98.980 32.600 99.330 33.200 ;
        RECT 98.980 32.400 102.930 32.600 ;
        RECT 98.980 31.800 99.330 32.400 ;
        RECT 98.980 31.600 102.930 31.800 ;
        RECT 98.980 31.000 99.330 31.600 ;
        RECT 98.980 30.800 102.930 31.000 ;
        RECT 98.980 30.400 99.330 30.800 ;
        RECT 95.780 22.000 95.980 29.600 ;
        RECT 96.580 22.000 96.780 29.600 ;
        RECT 97.380 22.000 97.580 29.600 ;
        RECT 98.180 22.000 98.380 29.600 ;
        RECT 98.980 29.200 99.330 29.600 ;
        RECT 98.980 29.000 102.930 29.200 ;
        RECT 98.980 28.400 99.330 29.000 ;
        RECT 98.980 28.200 102.930 28.400 ;
        RECT 98.980 27.600 99.330 28.200 ;
        RECT 98.980 27.400 102.930 27.600 ;
        RECT 98.980 26.800 99.330 27.400 ;
        RECT 98.980 26.600 102.930 26.800 ;
        RECT 103.930 26.750 104.330 33.250 ;
        RECT 98.980 26.000 99.330 26.600 ;
        RECT 98.980 25.800 102.930 26.000 ;
        RECT 98.980 25.200 99.330 25.800 ;
        RECT 98.980 25.000 102.930 25.200 ;
        RECT 98.980 24.400 99.330 25.000 ;
        RECT 103.880 24.450 104.730 26.750 ;
        RECT 98.980 24.200 102.930 24.400 ;
        RECT 98.980 23.600 99.330 24.200 ;
        RECT 98.980 23.400 102.930 23.600 ;
        RECT 98.980 22.800 99.330 23.400 ;
        RECT 98.980 22.600 102.930 22.800 ;
        RECT 98.980 22.000 99.330 22.600 ;
        RECT 86.530 21.400 102.930 22.000 ;
        RECT 89.180 20.800 91.480 20.850 ;
        RECT 97.980 20.800 100.280 20.850 ;
        RECT 103.930 20.800 104.330 24.450 ;
        RECT 105.340 22.590 105.700 22.970 ;
        RECT 105.970 22.590 106.330 22.970 ;
        RECT 106.570 22.590 106.930 22.970 ;
        RECT 105.340 22.000 105.700 22.380 ;
        RECT 105.970 22.000 106.330 22.380 ;
        RECT 106.570 22.000 106.930 22.380 ;
        RECT 85.130 20.400 104.330 20.800 ;
        RECT 9.180 19.600 11.480 20.400 ;
        RECT 17.980 19.600 20.280 20.400 ;
        RECT 29.180 19.600 31.480 20.400 ;
        RECT 37.980 19.600 40.280 20.400 ;
        RECT 49.180 19.600 51.480 20.400 ;
        RECT 57.980 19.600 60.280 20.400 ;
        RECT 69.180 19.600 71.480 20.400 ;
        RECT 77.980 19.600 80.280 20.400 ;
        RECT 89.180 19.600 91.480 20.400 ;
        RECT 97.980 19.600 100.280 20.400 ;
        RECT 5.130 19.200 24.330 19.600 ;
        RECT 2.515 17.260 2.875 17.640 ;
        RECT 3.145 17.260 3.505 17.640 ;
        RECT 3.745 17.260 4.105 17.640 ;
        RECT 2.515 16.670 2.875 17.050 ;
        RECT 3.145 16.670 3.505 17.050 ;
        RECT 3.745 16.670 4.105 17.050 ;
        RECT 5.130 15.550 5.530 19.200 ;
        RECT 9.180 19.150 11.480 19.200 ;
        RECT 17.980 19.150 20.280 19.200 ;
        RECT 6.530 18.000 22.930 18.600 ;
        RECT 10.130 17.400 10.480 18.000 ;
        RECT 6.530 17.200 10.480 17.400 ;
        RECT 10.130 16.600 10.480 17.200 ;
        RECT 6.530 16.400 10.480 16.600 ;
        RECT 10.130 15.800 10.480 16.400 ;
        RECT 6.530 15.600 10.480 15.800 ;
        RECT 2.315 13.255 5.580 15.550 ;
        RECT 10.130 15.000 10.480 15.600 ;
        RECT 6.530 14.800 10.480 15.000 ;
        RECT 10.130 14.200 10.480 14.800 ;
        RECT 6.530 14.000 10.480 14.200 ;
        RECT 10.130 13.400 10.480 14.000 ;
        RECT 4.730 13.250 5.580 13.255 ;
        RECT 5.130 6.750 5.530 13.250 ;
        RECT 6.530 13.200 10.480 13.400 ;
        RECT 10.130 12.600 10.480 13.200 ;
        RECT 6.530 12.400 10.480 12.600 ;
        RECT 10.130 11.800 10.480 12.400 ;
        RECT 6.530 11.600 10.480 11.800 ;
        RECT 10.130 11.000 10.480 11.600 ;
        RECT 6.530 10.800 10.480 11.000 ;
        RECT 10.130 10.400 10.480 10.800 ;
        RECT 11.080 10.400 11.280 18.000 ;
        RECT 11.880 10.400 12.080 18.000 ;
        RECT 12.680 10.400 12.880 18.000 ;
        RECT 13.480 10.400 13.680 18.000 ;
        RECT 10.130 9.200 10.480 9.600 ;
        RECT 6.530 9.000 10.480 9.200 ;
        RECT 10.130 8.400 10.480 9.000 ;
        RECT 6.530 8.200 10.480 8.400 ;
        RECT 10.130 7.600 10.480 8.200 ;
        RECT 6.530 7.400 10.480 7.600 ;
        RECT 10.130 6.800 10.480 7.400 ;
        RECT 4.730 6.745 5.580 6.750 ;
        RECT 2.315 4.450 5.580 6.745 ;
        RECT 6.530 6.600 10.480 6.800 ;
        RECT 10.130 6.000 10.480 6.600 ;
        RECT 6.530 5.800 10.480 6.000 ;
        RECT 10.130 5.200 10.480 5.800 ;
        RECT 6.530 5.000 10.480 5.200 ;
        RECT 2.515 3.145 2.875 3.525 ;
        RECT 3.145 3.145 3.505 3.525 ;
        RECT 3.745 3.145 4.105 3.525 ;
        RECT 2.515 2.555 2.875 2.935 ;
        RECT 3.145 2.555 3.505 2.935 ;
        RECT 3.745 2.555 4.105 2.935 ;
        RECT 5.130 0.800 5.530 4.450 ;
        RECT 10.130 4.400 10.480 5.000 ;
        RECT 6.530 4.200 10.480 4.400 ;
        RECT 10.130 3.600 10.480 4.200 ;
        RECT 6.530 3.400 10.480 3.600 ;
        RECT 10.130 2.800 10.480 3.400 ;
        RECT 6.530 2.600 10.480 2.800 ;
        RECT 10.130 2.000 10.480 2.600 ;
        RECT 11.080 2.000 11.280 9.600 ;
        RECT 11.880 2.000 12.080 9.600 ;
        RECT 12.680 2.000 12.880 9.600 ;
        RECT 13.480 2.000 13.680 9.600 ;
        RECT 14.280 2.000 15.180 18.000 ;
        RECT 15.780 10.400 15.980 18.000 ;
        RECT 16.580 10.400 16.780 18.000 ;
        RECT 17.380 10.400 17.580 18.000 ;
        RECT 18.180 10.400 18.380 18.000 ;
        RECT 18.980 17.400 19.330 18.000 ;
        RECT 18.980 17.200 22.930 17.400 ;
        RECT 18.980 16.600 19.330 17.200 ;
        RECT 18.980 16.400 22.930 16.600 ;
        RECT 18.980 15.800 19.330 16.400 ;
        RECT 18.980 15.600 22.930 15.800 ;
        RECT 18.980 15.000 19.330 15.600 ;
        RECT 23.930 15.550 24.330 19.200 ;
        RECT 25.130 19.200 44.330 19.600 ;
        RECT 25.130 15.550 25.530 19.200 ;
        RECT 29.180 19.150 31.480 19.200 ;
        RECT 37.980 19.150 40.280 19.200 ;
        RECT 26.530 18.000 42.930 18.600 ;
        RECT 30.130 17.400 30.480 18.000 ;
        RECT 26.530 17.200 30.480 17.400 ;
        RECT 30.130 16.600 30.480 17.200 ;
        RECT 26.530 16.400 30.480 16.600 ;
        RECT 30.130 15.800 30.480 16.400 ;
        RECT 26.530 15.600 30.480 15.800 ;
        RECT 18.980 14.800 22.930 15.000 ;
        RECT 18.980 14.200 19.330 14.800 ;
        RECT 18.980 14.000 22.930 14.200 ;
        RECT 18.980 13.400 19.330 14.000 ;
        RECT 18.980 13.200 22.930 13.400 ;
        RECT 23.880 13.250 25.580 15.550 ;
        RECT 30.130 15.000 30.480 15.600 ;
        RECT 26.530 14.800 30.480 15.000 ;
        RECT 30.130 14.200 30.480 14.800 ;
        RECT 26.530 14.000 30.480 14.200 ;
        RECT 30.130 13.400 30.480 14.000 ;
        RECT 18.980 12.600 19.330 13.200 ;
        RECT 18.980 12.400 22.930 12.600 ;
        RECT 18.980 11.800 19.330 12.400 ;
        RECT 18.980 11.600 22.930 11.800 ;
        RECT 18.980 11.000 19.330 11.600 ;
        RECT 18.980 10.800 22.930 11.000 ;
        RECT 18.980 10.400 19.330 10.800 ;
        RECT 15.780 2.000 15.980 9.600 ;
        RECT 16.580 2.000 16.780 9.600 ;
        RECT 17.380 2.000 17.580 9.600 ;
        RECT 18.180 2.000 18.380 9.600 ;
        RECT 18.980 9.200 19.330 9.600 ;
        RECT 18.980 9.000 22.930 9.200 ;
        RECT 18.980 8.400 19.330 9.000 ;
        RECT 18.980 8.200 22.930 8.400 ;
        RECT 18.980 7.600 19.330 8.200 ;
        RECT 18.980 7.400 22.930 7.600 ;
        RECT 18.980 6.800 19.330 7.400 ;
        RECT 18.980 6.600 22.930 6.800 ;
        RECT 23.930 6.750 24.330 13.250 ;
        RECT 25.130 6.750 25.530 13.250 ;
        RECT 26.530 13.200 30.480 13.400 ;
        RECT 30.130 12.600 30.480 13.200 ;
        RECT 26.530 12.400 30.480 12.600 ;
        RECT 30.130 11.800 30.480 12.400 ;
        RECT 26.530 11.600 30.480 11.800 ;
        RECT 30.130 11.000 30.480 11.600 ;
        RECT 26.530 10.800 30.480 11.000 ;
        RECT 30.130 10.400 30.480 10.800 ;
        RECT 31.080 10.400 31.280 18.000 ;
        RECT 31.880 10.400 32.080 18.000 ;
        RECT 32.680 10.400 32.880 18.000 ;
        RECT 33.480 10.400 33.680 18.000 ;
        RECT 30.130 9.200 30.480 9.600 ;
        RECT 26.530 9.000 30.480 9.200 ;
        RECT 30.130 8.400 30.480 9.000 ;
        RECT 26.530 8.200 30.480 8.400 ;
        RECT 30.130 7.600 30.480 8.200 ;
        RECT 26.530 7.400 30.480 7.600 ;
        RECT 30.130 6.800 30.480 7.400 ;
        RECT 18.980 6.000 19.330 6.600 ;
        RECT 18.980 5.800 22.930 6.000 ;
        RECT 18.980 5.200 19.330 5.800 ;
        RECT 18.980 5.000 22.930 5.200 ;
        RECT 18.980 4.400 19.330 5.000 ;
        RECT 23.880 4.450 25.580 6.750 ;
        RECT 26.530 6.600 30.480 6.800 ;
        RECT 30.130 6.000 30.480 6.600 ;
        RECT 26.530 5.800 30.480 6.000 ;
        RECT 30.130 5.200 30.480 5.800 ;
        RECT 26.530 5.000 30.480 5.200 ;
        RECT 18.980 4.200 22.930 4.400 ;
        RECT 18.980 3.600 19.330 4.200 ;
        RECT 18.980 3.400 22.930 3.600 ;
        RECT 18.980 2.800 19.330 3.400 ;
        RECT 18.980 2.600 22.930 2.800 ;
        RECT 18.980 2.000 19.330 2.600 ;
        RECT 6.530 1.400 22.930 2.000 ;
        RECT 9.180 0.800 11.480 0.850 ;
        RECT 17.980 0.800 20.280 0.850 ;
        RECT 23.930 0.800 24.330 4.450 ;
        RECT 5.130 0.400 24.330 0.800 ;
        RECT 25.130 0.800 25.530 4.450 ;
        RECT 30.130 4.400 30.480 5.000 ;
        RECT 26.530 4.200 30.480 4.400 ;
        RECT 30.130 3.600 30.480 4.200 ;
        RECT 26.530 3.400 30.480 3.600 ;
        RECT 30.130 2.800 30.480 3.400 ;
        RECT 26.530 2.600 30.480 2.800 ;
        RECT 30.130 2.000 30.480 2.600 ;
        RECT 31.080 2.000 31.280 9.600 ;
        RECT 31.880 2.000 32.080 9.600 ;
        RECT 32.680 2.000 32.880 9.600 ;
        RECT 33.480 2.000 33.680 9.600 ;
        RECT 34.280 2.000 35.180 18.000 ;
        RECT 35.780 10.400 35.980 18.000 ;
        RECT 36.580 10.400 36.780 18.000 ;
        RECT 37.380 10.400 37.580 18.000 ;
        RECT 38.180 10.400 38.380 18.000 ;
        RECT 38.980 17.400 39.330 18.000 ;
        RECT 38.980 17.200 42.930 17.400 ;
        RECT 38.980 16.600 39.330 17.200 ;
        RECT 38.980 16.400 42.930 16.600 ;
        RECT 38.980 15.800 39.330 16.400 ;
        RECT 38.980 15.600 42.930 15.800 ;
        RECT 38.980 15.000 39.330 15.600 ;
        RECT 43.930 15.550 44.330 19.200 ;
        RECT 45.130 19.200 64.330 19.600 ;
        RECT 45.130 15.550 45.530 19.200 ;
        RECT 49.180 19.150 51.480 19.200 ;
        RECT 57.980 19.150 60.280 19.200 ;
        RECT 46.530 18.000 62.930 18.600 ;
        RECT 50.130 17.400 50.480 18.000 ;
        RECT 46.530 17.200 50.480 17.400 ;
        RECT 50.130 16.600 50.480 17.200 ;
        RECT 46.530 16.400 50.480 16.600 ;
        RECT 50.130 15.800 50.480 16.400 ;
        RECT 46.530 15.600 50.480 15.800 ;
        RECT 38.980 14.800 42.930 15.000 ;
        RECT 38.980 14.200 39.330 14.800 ;
        RECT 38.980 14.000 42.930 14.200 ;
        RECT 38.980 13.400 39.330 14.000 ;
        RECT 38.980 13.200 42.930 13.400 ;
        RECT 43.880 13.250 45.580 15.550 ;
        RECT 50.130 15.000 50.480 15.600 ;
        RECT 46.530 14.800 50.480 15.000 ;
        RECT 50.130 14.200 50.480 14.800 ;
        RECT 46.530 14.000 50.480 14.200 ;
        RECT 50.130 13.400 50.480 14.000 ;
        RECT 38.980 12.600 39.330 13.200 ;
        RECT 38.980 12.400 42.930 12.600 ;
        RECT 38.980 11.800 39.330 12.400 ;
        RECT 38.980 11.600 42.930 11.800 ;
        RECT 38.980 11.000 39.330 11.600 ;
        RECT 38.980 10.800 42.930 11.000 ;
        RECT 38.980 10.400 39.330 10.800 ;
        RECT 35.780 2.000 35.980 9.600 ;
        RECT 36.580 2.000 36.780 9.600 ;
        RECT 37.380 2.000 37.580 9.600 ;
        RECT 38.180 2.000 38.380 9.600 ;
        RECT 38.980 9.200 39.330 9.600 ;
        RECT 38.980 9.000 42.930 9.200 ;
        RECT 38.980 8.400 39.330 9.000 ;
        RECT 38.980 8.200 42.930 8.400 ;
        RECT 38.980 7.600 39.330 8.200 ;
        RECT 38.980 7.400 42.930 7.600 ;
        RECT 38.980 6.800 39.330 7.400 ;
        RECT 38.980 6.600 42.930 6.800 ;
        RECT 43.930 6.750 44.330 13.250 ;
        RECT 45.130 6.750 45.530 13.250 ;
        RECT 46.530 13.200 50.480 13.400 ;
        RECT 50.130 12.600 50.480 13.200 ;
        RECT 46.530 12.400 50.480 12.600 ;
        RECT 50.130 11.800 50.480 12.400 ;
        RECT 46.530 11.600 50.480 11.800 ;
        RECT 50.130 11.000 50.480 11.600 ;
        RECT 46.530 10.800 50.480 11.000 ;
        RECT 50.130 10.400 50.480 10.800 ;
        RECT 51.080 10.400 51.280 18.000 ;
        RECT 51.880 10.400 52.080 18.000 ;
        RECT 52.680 10.400 52.880 18.000 ;
        RECT 53.480 10.400 53.680 18.000 ;
        RECT 50.130 9.200 50.480 9.600 ;
        RECT 46.530 9.000 50.480 9.200 ;
        RECT 50.130 8.400 50.480 9.000 ;
        RECT 46.530 8.200 50.480 8.400 ;
        RECT 50.130 7.600 50.480 8.200 ;
        RECT 46.530 7.400 50.480 7.600 ;
        RECT 50.130 6.800 50.480 7.400 ;
        RECT 38.980 6.000 39.330 6.600 ;
        RECT 38.980 5.800 42.930 6.000 ;
        RECT 38.980 5.200 39.330 5.800 ;
        RECT 38.980 5.000 42.930 5.200 ;
        RECT 38.980 4.400 39.330 5.000 ;
        RECT 43.880 4.450 45.580 6.750 ;
        RECT 46.530 6.600 50.480 6.800 ;
        RECT 50.130 6.000 50.480 6.600 ;
        RECT 46.530 5.800 50.480 6.000 ;
        RECT 50.130 5.200 50.480 5.800 ;
        RECT 46.530 5.000 50.480 5.200 ;
        RECT 38.980 4.200 42.930 4.400 ;
        RECT 38.980 3.600 39.330 4.200 ;
        RECT 38.980 3.400 42.930 3.600 ;
        RECT 38.980 2.800 39.330 3.400 ;
        RECT 38.980 2.600 42.930 2.800 ;
        RECT 38.980 2.000 39.330 2.600 ;
        RECT 26.530 1.400 42.930 2.000 ;
        RECT 29.180 0.800 31.480 0.850 ;
        RECT 37.980 0.800 40.280 0.850 ;
        RECT 43.930 0.800 44.330 4.450 ;
        RECT 25.130 0.400 44.330 0.800 ;
        RECT 45.130 0.800 45.530 4.450 ;
        RECT 50.130 4.400 50.480 5.000 ;
        RECT 46.530 4.200 50.480 4.400 ;
        RECT 50.130 3.600 50.480 4.200 ;
        RECT 46.530 3.400 50.480 3.600 ;
        RECT 50.130 2.800 50.480 3.400 ;
        RECT 46.530 2.600 50.480 2.800 ;
        RECT 50.130 2.000 50.480 2.600 ;
        RECT 51.080 2.000 51.280 9.600 ;
        RECT 51.880 2.000 52.080 9.600 ;
        RECT 52.680 2.000 52.880 9.600 ;
        RECT 53.480 2.000 53.680 9.600 ;
        RECT 54.280 2.000 55.180 18.000 ;
        RECT 55.780 10.400 55.980 18.000 ;
        RECT 56.580 10.400 56.780 18.000 ;
        RECT 57.380 10.400 57.580 18.000 ;
        RECT 58.180 10.400 58.380 18.000 ;
        RECT 58.980 17.400 59.330 18.000 ;
        RECT 58.980 17.200 62.930 17.400 ;
        RECT 58.980 16.600 59.330 17.200 ;
        RECT 58.980 16.400 62.930 16.600 ;
        RECT 58.980 15.800 59.330 16.400 ;
        RECT 58.980 15.600 62.930 15.800 ;
        RECT 58.980 15.000 59.330 15.600 ;
        RECT 63.930 15.550 64.330 19.200 ;
        RECT 65.130 19.200 84.330 19.600 ;
        RECT 65.130 15.550 65.530 19.200 ;
        RECT 69.180 19.150 71.480 19.200 ;
        RECT 77.980 19.150 80.280 19.200 ;
        RECT 66.530 18.000 82.930 18.600 ;
        RECT 70.130 17.400 70.480 18.000 ;
        RECT 66.530 17.200 70.480 17.400 ;
        RECT 70.130 16.600 70.480 17.200 ;
        RECT 66.530 16.400 70.480 16.600 ;
        RECT 70.130 15.800 70.480 16.400 ;
        RECT 66.530 15.600 70.480 15.800 ;
        RECT 58.980 14.800 62.930 15.000 ;
        RECT 58.980 14.200 59.330 14.800 ;
        RECT 58.980 14.000 62.930 14.200 ;
        RECT 58.980 13.400 59.330 14.000 ;
        RECT 58.980 13.200 62.930 13.400 ;
        RECT 63.880 13.250 65.580 15.550 ;
        RECT 70.130 15.000 70.480 15.600 ;
        RECT 66.530 14.800 70.480 15.000 ;
        RECT 70.130 14.200 70.480 14.800 ;
        RECT 66.530 14.000 70.480 14.200 ;
        RECT 70.130 13.400 70.480 14.000 ;
        RECT 58.980 12.600 59.330 13.200 ;
        RECT 58.980 12.400 62.930 12.600 ;
        RECT 58.980 11.800 59.330 12.400 ;
        RECT 58.980 11.600 62.930 11.800 ;
        RECT 58.980 11.000 59.330 11.600 ;
        RECT 58.980 10.800 62.930 11.000 ;
        RECT 58.980 10.400 59.330 10.800 ;
        RECT 55.780 2.000 55.980 9.600 ;
        RECT 56.580 2.000 56.780 9.600 ;
        RECT 57.380 2.000 57.580 9.600 ;
        RECT 58.180 2.000 58.380 9.600 ;
        RECT 58.980 9.200 59.330 9.600 ;
        RECT 58.980 9.000 62.930 9.200 ;
        RECT 58.980 8.400 59.330 9.000 ;
        RECT 58.980 8.200 62.930 8.400 ;
        RECT 58.980 7.600 59.330 8.200 ;
        RECT 58.980 7.400 62.930 7.600 ;
        RECT 58.980 6.800 59.330 7.400 ;
        RECT 58.980 6.600 62.930 6.800 ;
        RECT 63.930 6.750 64.330 13.250 ;
        RECT 65.130 6.750 65.530 13.250 ;
        RECT 66.530 13.200 70.480 13.400 ;
        RECT 70.130 12.600 70.480 13.200 ;
        RECT 66.530 12.400 70.480 12.600 ;
        RECT 70.130 11.800 70.480 12.400 ;
        RECT 66.530 11.600 70.480 11.800 ;
        RECT 70.130 11.000 70.480 11.600 ;
        RECT 66.530 10.800 70.480 11.000 ;
        RECT 70.130 10.400 70.480 10.800 ;
        RECT 71.080 10.400 71.280 18.000 ;
        RECT 71.880 10.400 72.080 18.000 ;
        RECT 72.680 10.400 72.880 18.000 ;
        RECT 73.480 10.400 73.680 18.000 ;
        RECT 70.130 9.200 70.480 9.600 ;
        RECT 66.530 9.000 70.480 9.200 ;
        RECT 70.130 8.400 70.480 9.000 ;
        RECT 66.530 8.200 70.480 8.400 ;
        RECT 70.130 7.600 70.480 8.200 ;
        RECT 66.530 7.400 70.480 7.600 ;
        RECT 70.130 6.800 70.480 7.400 ;
        RECT 58.980 6.000 59.330 6.600 ;
        RECT 58.980 5.800 62.930 6.000 ;
        RECT 58.980 5.200 59.330 5.800 ;
        RECT 58.980 5.000 62.930 5.200 ;
        RECT 58.980 4.400 59.330 5.000 ;
        RECT 63.880 4.450 65.580 6.750 ;
        RECT 66.530 6.600 70.480 6.800 ;
        RECT 70.130 6.000 70.480 6.600 ;
        RECT 66.530 5.800 70.480 6.000 ;
        RECT 70.130 5.200 70.480 5.800 ;
        RECT 66.530 5.000 70.480 5.200 ;
        RECT 58.980 4.200 62.930 4.400 ;
        RECT 58.980 3.600 59.330 4.200 ;
        RECT 58.980 3.400 62.930 3.600 ;
        RECT 58.980 2.800 59.330 3.400 ;
        RECT 58.980 2.600 62.930 2.800 ;
        RECT 58.980 2.000 59.330 2.600 ;
        RECT 46.530 1.400 62.930 2.000 ;
        RECT 49.180 0.800 51.480 0.850 ;
        RECT 57.980 0.800 60.280 0.850 ;
        RECT 63.930 0.800 64.330 4.450 ;
        RECT 45.130 0.400 64.330 0.800 ;
        RECT 65.130 0.800 65.530 4.450 ;
        RECT 70.130 4.400 70.480 5.000 ;
        RECT 66.530 4.200 70.480 4.400 ;
        RECT 70.130 3.600 70.480 4.200 ;
        RECT 66.530 3.400 70.480 3.600 ;
        RECT 70.130 2.800 70.480 3.400 ;
        RECT 66.530 2.600 70.480 2.800 ;
        RECT 70.130 2.000 70.480 2.600 ;
        RECT 71.080 2.000 71.280 9.600 ;
        RECT 71.880 2.000 72.080 9.600 ;
        RECT 72.680 2.000 72.880 9.600 ;
        RECT 73.480 2.000 73.680 9.600 ;
        RECT 74.280 2.000 75.180 18.000 ;
        RECT 75.780 10.400 75.980 18.000 ;
        RECT 76.580 10.400 76.780 18.000 ;
        RECT 77.380 10.400 77.580 18.000 ;
        RECT 78.180 10.400 78.380 18.000 ;
        RECT 78.980 17.400 79.330 18.000 ;
        RECT 78.980 17.200 82.930 17.400 ;
        RECT 78.980 16.600 79.330 17.200 ;
        RECT 78.980 16.400 82.930 16.600 ;
        RECT 78.980 15.800 79.330 16.400 ;
        RECT 78.980 15.600 82.930 15.800 ;
        RECT 78.980 15.000 79.330 15.600 ;
        RECT 83.930 15.550 84.330 19.200 ;
        RECT 85.130 19.200 104.330 19.600 ;
        RECT 85.130 15.550 85.530 19.200 ;
        RECT 89.180 19.150 91.480 19.200 ;
        RECT 97.980 19.150 100.280 19.200 ;
        RECT 86.530 18.000 102.930 18.600 ;
        RECT 90.130 17.400 90.480 18.000 ;
        RECT 86.530 17.200 90.480 17.400 ;
        RECT 90.130 16.600 90.480 17.200 ;
        RECT 86.530 16.400 90.480 16.600 ;
        RECT 90.130 15.800 90.480 16.400 ;
        RECT 86.530 15.600 90.480 15.800 ;
        RECT 78.980 14.800 82.930 15.000 ;
        RECT 78.980 14.200 79.330 14.800 ;
        RECT 78.980 14.000 82.930 14.200 ;
        RECT 78.980 13.400 79.330 14.000 ;
        RECT 78.980 13.200 82.930 13.400 ;
        RECT 83.880 13.250 85.580 15.550 ;
        RECT 90.130 15.000 90.480 15.600 ;
        RECT 86.530 14.800 90.480 15.000 ;
        RECT 90.130 14.200 90.480 14.800 ;
        RECT 86.530 14.000 90.480 14.200 ;
        RECT 90.130 13.400 90.480 14.000 ;
        RECT 78.980 12.600 79.330 13.200 ;
        RECT 78.980 12.400 82.930 12.600 ;
        RECT 78.980 11.800 79.330 12.400 ;
        RECT 78.980 11.600 82.930 11.800 ;
        RECT 78.980 11.000 79.330 11.600 ;
        RECT 78.980 10.800 82.930 11.000 ;
        RECT 78.980 10.400 79.330 10.800 ;
        RECT 75.780 2.000 75.980 9.600 ;
        RECT 76.580 2.000 76.780 9.600 ;
        RECT 77.380 2.000 77.580 9.600 ;
        RECT 78.180 2.000 78.380 9.600 ;
        RECT 78.980 9.200 79.330 9.600 ;
        RECT 78.980 9.000 82.930 9.200 ;
        RECT 78.980 8.400 79.330 9.000 ;
        RECT 78.980 8.200 82.930 8.400 ;
        RECT 78.980 7.600 79.330 8.200 ;
        RECT 78.980 7.400 82.930 7.600 ;
        RECT 78.980 6.800 79.330 7.400 ;
        RECT 78.980 6.600 82.930 6.800 ;
        RECT 83.930 6.750 84.330 13.250 ;
        RECT 85.130 6.750 85.530 13.250 ;
        RECT 86.530 13.200 90.480 13.400 ;
        RECT 90.130 12.600 90.480 13.200 ;
        RECT 86.530 12.400 90.480 12.600 ;
        RECT 90.130 11.800 90.480 12.400 ;
        RECT 86.530 11.600 90.480 11.800 ;
        RECT 90.130 11.000 90.480 11.600 ;
        RECT 86.530 10.800 90.480 11.000 ;
        RECT 90.130 10.400 90.480 10.800 ;
        RECT 91.080 10.400 91.280 18.000 ;
        RECT 91.880 10.400 92.080 18.000 ;
        RECT 92.680 10.400 92.880 18.000 ;
        RECT 93.480 10.400 93.680 18.000 ;
        RECT 90.130 9.200 90.480 9.600 ;
        RECT 86.530 9.000 90.480 9.200 ;
        RECT 90.130 8.400 90.480 9.000 ;
        RECT 86.530 8.200 90.480 8.400 ;
        RECT 90.130 7.600 90.480 8.200 ;
        RECT 86.530 7.400 90.480 7.600 ;
        RECT 90.130 6.800 90.480 7.400 ;
        RECT 78.980 6.000 79.330 6.600 ;
        RECT 78.980 5.800 82.930 6.000 ;
        RECT 78.980 5.200 79.330 5.800 ;
        RECT 78.980 5.000 82.930 5.200 ;
        RECT 78.980 4.400 79.330 5.000 ;
        RECT 83.880 4.450 85.580 6.750 ;
        RECT 86.530 6.600 90.480 6.800 ;
        RECT 90.130 6.000 90.480 6.600 ;
        RECT 86.530 5.800 90.480 6.000 ;
        RECT 90.130 5.200 90.480 5.800 ;
        RECT 86.530 5.000 90.480 5.200 ;
        RECT 78.980 4.200 82.930 4.400 ;
        RECT 78.980 3.600 79.330 4.200 ;
        RECT 78.980 3.400 82.930 3.600 ;
        RECT 78.980 2.800 79.330 3.400 ;
        RECT 78.980 2.600 82.930 2.800 ;
        RECT 78.980 2.000 79.330 2.600 ;
        RECT 66.530 1.400 82.930 2.000 ;
        RECT 69.180 0.800 71.480 0.850 ;
        RECT 77.980 0.800 80.280 0.850 ;
        RECT 83.930 0.800 84.330 4.450 ;
        RECT 65.130 0.400 84.330 0.800 ;
        RECT 85.130 0.800 85.530 4.450 ;
        RECT 90.130 4.400 90.480 5.000 ;
        RECT 86.530 4.200 90.480 4.400 ;
        RECT 90.130 3.600 90.480 4.200 ;
        RECT 86.530 3.400 90.480 3.600 ;
        RECT 90.130 2.800 90.480 3.400 ;
        RECT 86.530 2.600 90.480 2.800 ;
        RECT 90.130 2.000 90.480 2.600 ;
        RECT 91.080 2.000 91.280 9.600 ;
        RECT 91.880 2.000 92.080 9.600 ;
        RECT 92.680 2.000 92.880 9.600 ;
        RECT 93.480 2.000 93.680 9.600 ;
        RECT 94.280 2.000 95.180 18.000 ;
        RECT 95.780 10.400 95.980 18.000 ;
        RECT 96.580 10.400 96.780 18.000 ;
        RECT 97.380 10.400 97.580 18.000 ;
        RECT 98.180 10.400 98.380 18.000 ;
        RECT 98.980 17.400 99.330 18.000 ;
        RECT 98.980 17.200 102.930 17.400 ;
        RECT 98.980 16.600 99.330 17.200 ;
        RECT 98.980 16.400 102.930 16.600 ;
        RECT 98.980 15.800 99.330 16.400 ;
        RECT 98.980 15.600 102.930 15.800 ;
        RECT 98.980 15.000 99.330 15.600 ;
        RECT 103.930 15.550 104.330 19.200 ;
        RECT 105.340 16.805 105.700 17.185 ;
        RECT 105.970 16.805 106.330 17.185 ;
        RECT 106.570 16.805 106.930 17.185 ;
        RECT 105.340 16.215 105.700 16.595 ;
        RECT 105.970 16.215 106.330 16.595 ;
        RECT 106.570 16.215 106.930 16.595 ;
        RECT 98.980 14.800 102.930 15.000 ;
        RECT 98.980 14.200 99.330 14.800 ;
        RECT 98.980 14.000 102.930 14.200 ;
        RECT 98.980 13.400 99.330 14.000 ;
        RECT 98.980 13.200 102.930 13.400 ;
        RECT 103.880 13.250 104.730 15.550 ;
        RECT 98.980 12.600 99.330 13.200 ;
        RECT 98.980 12.400 102.930 12.600 ;
        RECT 98.980 11.800 99.330 12.400 ;
        RECT 98.980 11.600 102.930 11.800 ;
        RECT 98.980 11.000 99.330 11.600 ;
        RECT 98.980 10.800 102.930 11.000 ;
        RECT 98.980 10.400 99.330 10.800 ;
        RECT 95.780 2.000 95.980 9.600 ;
        RECT 96.580 2.000 96.780 9.600 ;
        RECT 97.380 2.000 97.580 9.600 ;
        RECT 98.180 2.000 98.380 9.600 ;
        RECT 98.980 9.200 99.330 9.600 ;
        RECT 98.980 9.000 102.930 9.200 ;
        RECT 98.980 8.400 99.330 9.000 ;
        RECT 98.980 8.200 102.930 8.400 ;
        RECT 98.980 7.600 99.330 8.200 ;
        RECT 98.980 7.400 102.930 7.600 ;
        RECT 98.980 6.800 99.330 7.400 ;
        RECT 98.980 6.600 102.930 6.800 ;
        RECT 103.930 6.750 104.330 13.250 ;
        RECT 98.980 6.000 99.330 6.600 ;
        RECT 98.980 5.800 102.930 6.000 ;
        RECT 98.980 5.200 99.330 5.800 ;
        RECT 98.980 5.000 102.930 5.200 ;
        RECT 98.980 4.400 99.330 5.000 ;
        RECT 103.880 4.450 104.730 6.750 ;
        RECT 98.980 4.200 102.930 4.400 ;
        RECT 98.980 3.600 99.330 4.200 ;
        RECT 98.980 3.400 102.930 3.600 ;
        RECT 98.980 2.800 99.330 3.400 ;
        RECT 98.980 2.600 102.930 2.800 ;
        RECT 98.980 2.000 99.330 2.600 ;
        RECT 86.530 1.400 102.930 2.000 ;
        RECT 89.180 0.800 91.480 0.850 ;
        RECT 97.980 0.800 100.280 0.850 ;
        RECT 103.930 0.800 104.330 4.450 ;
        RECT 105.340 2.590 105.700 2.970 ;
        RECT 105.970 2.590 106.330 2.970 ;
        RECT 106.570 2.590 106.930 2.970 ;
        RECT 105.340 2.000 105.700 2.380 ;
        RECT 105.970 2.000 106.330 2.380 ;
        RECT 106.570 2.000 106.930 2.380 ;
        RECT 85.130 0.400 104.330 0.800 ;
        RECT 9.180 0.000 11.480 0.400 ;
        RECT 17.980 0.000 20.280 0.400 ;
        RECT 29.180 0.000 31.480 0.400 ;
        RECT 37.980 0.000 40.280 0.400 ;
        RECT 49.180 0.000 51.480 0.400 ;
        RECT 57.980 0.000 60.280 0.400 ;
        RECT 69.180 0.000 71.480 0.400 ;
        RECT 77.980 0.000 80.280 0.400 ;
        RECT 89.180 0.000 91.480 0.400 ;
        RECT 97.980 0.000 100.280 0.400 ;
      LAYER mcon ;
        RECT 6.830 378.100 7.430 378.600 ;
        RECT 7.630 378.100 8.230 378.600 ;
        RECT 8.430 378.100 9.030 378.600 ;
        RECT 9.230 378.100 9.830 378.600 ;
        RECT 10.030 378.100 10.630 378.600 ;
        RECT 18.830 378.100 19.430 378.600 ;
        RECT 19.630 378.100 20.230 378.600 ;
        RECT 20.430 378.100 21.030 378.600 ;
        RECT 21.230 378.100 21.830 378.600 ;
        RECT 22.030 378.100 22.580 378.600 ;
        RECT 2.520 374.920 2.880 375.300 ;
        RECT 3.130 374.920 3.490 375.300 ;
        RECT 3.760 374.920 4.120 375.300 ;
        RECT 2.520 374.185 2.880 374.565 ;
        RECT 3.130 374.185 3.490 374.565 ;
        RECT 3.760 374.185 4.120 374.565 ;
        RECT 2.520 373.500 2.880 373.880 ;
        RECT 3.130 373.500 3.490 373.880 ;
        RECT 3.760 373.500 4.120 373.880 ;
        RECT 2.520 366.120 2.880 366.500 ;
        RECT 3.130 366.120 3.490 366.500 ;
        RECT 3.760 366.120 4.120 366.500 ;
        RECT 2.520 365.385 2.880 365.765 ;
        RECT 3.130 365.385 3.490 365.765 ;
        RECT 3.760 365.385 4.120 365.765 ;
        RECT 2.520 364.700 2.880 365.080 ;
        RECT 3.130 364.700 3.490 365.080 ;
        RECT 3.760 364.700 4.120 365.080 ;
        RECT 26.830 378.100 27.430 378.600 ;
        RECT 27.630 378.100 28.230 378.600 ;
        RECT 28.430 378.100 29.030 378.600 ;
        RECT 29.230 378.100 29.830 378.600 ;
        RECT 30.030 378.100 30.630 378.600 ;
        RECT 38.830 378.100 39.430 378.600 ;
        RECT 39.630 378.100 40.230 378.600 ;
        RECT 40.430 378.100 41.030 378.600 ;
        RECT 41.230 378.100 41.830 378.600 ;
        RECT 42.030 378.100 42.580 378.600 ;
        RECT 6.830 361.400 7.430 361.900 ;
        RECT 7.630 361.400 8.230 361.900 ;
        RECT 8.430 361.400 9.030 361.900 ;
        RECT 9.230 361.400 9.830 361.900 ;
        RECT 10.030 361.400 10.630 361.900 ;
        RECT 18.830 361.400 19.430 361.900 ;
        RECT 19.630 361.400 20.230 361.900 ;
        RECT 20.430 361.400 21.030 361.900 ;
        RECT 21.230 361.400 21.830 361.900 ;
        RECT 22.030 361.400 22.580 361.900 ;
        RECT 46.830 378.100 47.430 378.600 ;
        RECT 47.630 378.100 48.230 378.600 ;
        RECT 48.430 378.100 49.030 378.600 ;
        RECT 49.230 378.100 49.830 378.600 ;
        RECT 50.030 378.100 50.630 378.600 ;
        RECT 58.830 378.100 59.430 378.600 ;
        RECT 59.630 378.100 60.230 378.600 ;
        RECT 60.430 378.100 61.030 378.600 ;
        RECT 61.230 378.100 61.830 378.600 ;
        RECT 62.030 378.100 62.580 378.600 ;
        RECT 26.830 361.400 27.430 361.900 ;
        RECT 27.630 361.400 28.230 361.900 ;
        RECT 28.430 361.400 29.030 361.900 ;
        RECT 29.230 361.400 29.830 361.900 ;
        RECT 30.030 361.400 30.630 361.900 ;
        RECT 38.830 361.400 39.430 361.900 ;
        RECT 39.630 361.400 40.230 361.900 ;
        RECT 40.430 361.400 41.030 361.900 ;
        RECT 41.230 361.400 41.830 361.900 ;
        RECT 42.030 361.400 42.580 361.900 ;
        RECT 66.830 378.100 67.430 378.600 ;
        RECT 67.630 378.100 68.230 378.600 ;
        RECT 68.430 378.100 69.030 378.600 ;
        RECT 69.230 378.100 69.830 378.600 ;
        RECT 70.030 378.100 70.630 378.600 ;
        RECT 78.830 378.100 79.430 378.600 ;
        RECT 79.630 378.100 80.230 378.600 ;
        RECT 80.430 378.100 81.030 378.600 ;
        RECT 81.230 378.100 81.830 378.600 ;
        RECT 82.030 378.100 82.580 378.600 ;
        RECT 46.830 361.400 47.430 361.900 ;
        RECT 47.630 361.400 48.230 361.900 ;
        RECT 48.430 361.400 49.030 361.900 ;
        RECT 49.230 361.400 49.830 361.900 ;
        RECT 50.030 361.400 50.630 361.900 ;
        RECT 58.830 361.400 59.430 361.900 ;
        RECT 59.630 361.400 60.230 361.900 ;
        RECT 60.430 361.400 61.030 361.900 ;
        RECT 61.230 361.400 61.830 361.900 ;
        RECT 62.030 361.400 62.580 361.900 ;
        RECT 86.830 378.100 87.430 378.600 ;
        RECT 87.630 378.100 88.230 378.600 ;
        RECT 88.430 378.100 89.030 378.600 ;
        RECT 89.230 378.100 89.830 378.600 ;
        RECT 90.030 378.100 90.630 378.600 ;
        RECT 98.830 378.100 99.430 378.600 ;
        RECT 99.630 378.100 100.230 378.600 ;
        RECT 100.430 378.100 101.030 378.600 ;
        RECT 101.230 378.100 101.830 378.600 ;
        RECT 102.030 378.100 102.580 378.600 ;
        RECT 66.830 361.400 67.430 361.900 ;
        RECT 67.630 361.400 68.230 361.900 ;
        RECT 68.430 361.400 69.030 361.900 ;
        RECT 69.230 361.400 69.830 361.900 ;
        RECT 70.030 361.400 70.630 361.900 ;
        RECT 78.830 361.400 79.430 361.900 ;
        RECT 79.630 361.400 80.230 361.900 ;
        RECT 80.430 361.400 81.030 361.900 ;
        RECT 81.230 361.400 81.830 361.900 ;
        RECT 82.030 361.400 82.580 361.900 ;
        RECT 86.830 361.400 87.430 361.900 ;
        RECT 87.630 361.400 88.230 361.900 ;
        RECT 88.430 361.400 89.030 361.900 ;
        RECT 89.230 361.400 89.830 361.900 ;
        RECT 90.030 361.400 90.630 361.900 ;
        RECT 98.830 361.400 99.430 361.900 ;
        RECT 99.630 361.400 100.230 361.900 ;
        RECT 100.430 361.400 101.030 361.900 ;
        RECT 101.230 361.400 101.830 361.900 ;
        RECT 102.030 361.400 102.580 361.900 ;
        RECT 6.830 358.100 7.430 358.600 ;
        RECT 7.630 358.100 8.230 358.600 ;
        RECT 8.430 358.100 9.030 358.600 ;
        RECT 9.230 358.100 9.830 358.600 ;
        RECT 10.030 358.100 10.630 358.600 ;
        RECT 18.830 358.100 19.430 358.600 ;
        RECT 19.630 358.100 20.230 358.600 ;
        RECT 20.430 358.100 21.030 358.600 ;
        RECT 21.230 358.100 21.830 358.600 ;
        RECT 22.030 358.100 22.580 358.600 ;
        RECT 2.520 354.920 2.880 355.300 ;
        RECT 3.130 354.920 3.490 355.300 ;
        RECT 3.760 354.920 4.120 355.300 ;
        RECT 2.520 354.185 2.880 354.565 ;
        RECT 3.130 354.185 3.490 354.565 ;
        RECT 3.760 354.185 4.120 354.565 ;
        RECT 2.520 353.500 2.880 353.880 ;
        RECT 3.130 353.500 3.490 353.880 ;
        RECT 3.760 353.500 4.120 353.880 ;
        RECT 2.520 346.120 2.880 346.500 ;
        RECT 3.130 346.120 3.490 346.500 ;
        RECT 3.760 346.120 4.120 346.500 ;
        RECT 2.520 345.385 2.880 345.765 ;
        RECT 3.130 345.385 3.490 345.765 ;
        RECT 3.760 345.385 4.120 345.765 ;
        RECT 2.520 344.700 2.880 345.080 ;
        RECT 3.130 344.700 3.490 345.080 ;
        RECT 3.760 344.700 4.120 345.080 ;
        RECT 26.830 358.100 27.430 358.600 ;
        RECT 27.630 358.100 28.230 358.600 ;
        RECT 28.430 358.100 29.030 358.600 ;
        RECT 29.230 358.100 29.830 358.600 ;
        RECT 30.030 358.100 30.630 358.600 ;
        RECT 38.830 358.100 39.430 358.600 ;
        RECT 39.630 358.100 40.230 358.600 ;
        RECT 40.430 358.100 41.030 358.600 ;
        RECT 41.230 358.100 41.830 358.600 ;
        RECT 42.030 358.100 42.580 358.600 ;
        RECT 6.830 341.400 7.430 341.900 ;
        RECT 7.630 341.400 8.230 341.900 ;
        RECT 8.430 341.400 9.030 341.900 ;
        RECT 9.230 341.400 9.830 341.900 ;
        RECT 10.030 341.400 10.630 341.900 ;
        RECT 18.830 341.400 19.430 341.900 ;
        RECT 19.630 341.400 20.230 341.900 ;
        RECT 20.430 341.400 21.030 341.900 ;
        RECT 21.230 341.400 21.830 341.900 ;
        RECT 22.030 341.400 22.580 341.900 ;
        RECT 46.830 358.100 47.430 358.600 ;
        RECT 47.630 358.100 48.230 358.600 ;
        RECT 48.430 358.100 49.030 358.600 ;
        RECT 49.230 358.100 49.830 358.600 ;
        RECT 50.030 358.100 50.630 358.600 ;
        RECT 58.830 358.100 59.430 358.600 ;
        RECT 59.630 358.100 60.230 358.600 ;
        RECT 60.430 358.100 61.030 358.600 ;
        RECT 61.230 358.100 61.830 358.600 ;
        RECT 62.030 358.100 62.580 358.600 ;
        RECT 26.830 341.400 27.430 341.900 ;
        RECT 27.630 341.400 28.230 341.900 ;
        RECT 28.430 341.400 29.030 341.900 ;
        RECT 29.230 341.400 29.830 341.900 ;
        RECT 30.030 341.400 30.630 341.900 ;
        RECT 38.830 341.400 39.430 341.900 ;
        RECT 39.630 341.400 40.230 341.900 ;
        RECT 40.430 341.400 41.030 341.900 ;
        RECT 41.230 341.400 41.830 341.900 ;
        RECT 42.030 341.400 42.580 341.900 ;
        RECT 66.830 358.100 67.430 358.600 ;
        RECT 67.630 358.100 68.230 358.600 ;
        RECT 68.430 358.100 69.030 358.600 ;
        RECT 69.230 358.100 69.830 358.600 ;
        RECT 70.030 358.100 70.630 358.600 ;
        RECT 78.830 358.100 79.430 358.600 ;
        RECT 79.630 358.100 80.230 358.600 ;
        RECT 80.430 358.100 81.030 358.600 ;
        RECT 81.230 358.100 81.830 358.600 ;
        RECT 82.030 358.100 82.580 358.600 ;
        RECT 46.830 341.400 47.430 341.900 ;
        RECT 47.630 341.400 48.230 341.900 ;
        RECT 48.430 341.400 49.030 341.900 ;
        RECT 49.230 341.400 49.830 341.900 ;
        RECT 50.030 341.400 50.630 341.900 ;
        RECT 58.830 341.400 59.430 341.900 ;
        RECT 59.630 341.400 60.230 341.900 ;
        RECT 60.430 341.400 61.030 341.900 ;
        RECT 61.230 341.400 61.830 341.900 ;
        RECT 62.030 341.400 62.580 341.900 ;
        RECT 86.830 358.100 87.430 358.600 ;
        RECT 87.630 358.100 88.230 358.600 ;
        RECT 88.430 358.100 89.030 358.600 ;
        RECT 89.230 358.100 89.830 358.600 ;
        RECT 90.030 358.100 90.630 358.600 ;
        RECT 98.830 358.100 99.430 358.600 ;
        RECT 99.630 358.100 100.230 358.600 ;
        RECT 100.430 358.100 101.030 358.600 ;
        RECT 101.230 358.100 101.830 358.600 ;
        RECT 102.030 358.100 102.580 358.600 ;
        RECT 66.830 341.400 67.430 341.900 ;
        RECT 67.630 341.400 68.230 341.900 ;
        RECT 68.430 341.400 69.030 341.900 ;
        RECT 69.230 341.400 69.830 341.900 ;
        RECT 70.030 341.400 70.630 341.900 ;
        RECT 78.830 341.400 79.430 341.900 ;
        RECT 79.630 341.400 80.230 341.900 ;
        RECT 80.430 341.400 81.030 341.900 ;
        RECT 81.230 341.400 81.830 341.900 ;
        RECT 82.030 341.400 82.580 341.900 ;
        RECT 86.830 341.400 87.430 341.900 ;
        RECT 87.630 341.400 88.230 341.900 ;
        RECT 88.430 341.400 89.030 341.900 ;
        RECT 89.230 341.400 89.830 341.900 ;
        RECT 90.030 341.400 90.630 341.900 ;
        RECT 98.830 341.400 99.430 341.900 ;
        RECT 99.630 341.400 100.230 341.900 ;
        RECT 100.430 341.400 101.030 341.900 ;
        RECT 101.230 341.400 101.830 341.900 ;
        RECT 102.030 341.400 102.580 341.900 ;
        RECT 6.830 338.100 7.430 338.600 ;
        RECT 7.630 338.100 8.230 338.600 ;
        RECT 8.430 338.100 9.030 338.600 ;
        RECT 9.230 338.100 9.830 338.600 ;
        RECT 10.030 338.100 10.630 338.600 ;
        RECT 18.830 338.100 19.430 338.600 ;
        RECT 19.630 338.100 20.230 338.600 ;
        RECT 20.430 338.100 21.030 338.600 ;
        RECT 21.230 338.100 21.830 338.600 ;
        RECT 22.030 338.100 22.580 338.600 ;
        RECT 2.520 334.920 2.880 335.300 ;
        RECT 3.130 334.920 3.490 335.300 ;
        RECT 3.760 334.920 4.120 335.300 ;
        RECT 2.520 334.185 2.880 334.565 ;
        RECT 3.130 334.185 3.490 334.565 ;
        RECT 3.760 334.185 4.120 334.565 ;
        RECT 2.520 333.500 2.880 333.880 ;
        RECT 3.130 333.500 3.490 333.880 ;
        RECT 3.760 333.500 4.120 333.880 ;
        RECT 2.520 326.125 2.880 326.505 ;
        RECT 3.130 326.125 3.490 326.505 ;
        RECT 3.760 326.125 4.120 326.505 ;
        RECT 2.520 325.390 2.880 325.770 ;
        RECT 3.130 325.390 3.490 325.770 ;
        RECT 3.760 325.390 4.120 325.770 ;
        RECT 2.520 324.705 2.880 325.085 ;
        RECT 3.130 324.705 3.490 325.085 ;
        RECT 3.760 324.705 4.120 325.085 ;
        RECT 26.830 338.100 27.430 338.600 ;
        RECT 27.630 338.100 28.230 338.600 ;
        RECT 28.430 338.100 29.030 338.600 ;
        RECT 29.230 338.100 29.830 338.600 ;
        RECT 30.030 338.100 30.630 338.600 ;
        RECT 38.830 338.100 39.430 338.600 ;
        RECT 39.630 338.100 40.230 338.600 ;
        RECT 40.430 338.100 41.030 338.600 ;
        RECT 41.230 338.100 41.830 338.600 ;
        RECT 42.030 338.100 42.580 338.600 ;
        RECT 6.830 321.400 7.430 321.900 ;
        RECT 7.630 321.400 8.230 321.900 ;
        RECT 8.430 321.400 9.030 321.900 ;
        RECT 9.230 321.400 9.830 321.900 ;
        RECT 10.030 321.400 10.630 321.900 ;
        RECT 18.830 321.400 19.430 321.900 ;
        RECT 19.630 321.400 20.230 321.900 ;
        RECT 20.430 321.400 21.030 321.900 ;
        RECT 21.230 321.400 21.830 321.900 ;
        RECT 22.030 321.400 22.580 321.900 ;
        RECT 46.830 338.100 47.430 338.600 ;
        RECT 47.630 338.100 48.230 338.600 ;
        RECT 48.430 338.100 49.030 338.600 ;
        RECT 49.230 338.100 49.830 338.600 ;
        RECT 50.030 338.100 50.630 338.600 ;
        RECT 58.830 338.100 59.430 338.600 ;
        RECT 59.630 338.100 60.230 338.600 ;
        RECT 60.430 338.100 61.030 338.600 ;
        RECT 61.230 338.100 61.830 338.600 ;
        RECT 62.030 338.100 62.580 338.600 ;
        RECT 26.830 321.400 27.430 321.900 ;
        RECT 27.630 321.400 28.230 321.900 ;
        RECT 28.430 321.400 29.030 321.900 ;
        RECT 29.230 321.400 29.830 321.900 ;
        RECT 30.030 321.400 30.630 321.900 ;
        RECT 38.830 321.400 39.430 321.900 ;
        RECT 39.630 321.400 40.230 321.900 ;
        RECT 40.430 321.400 41.030 321.900 ;
        RECT 41.230 321.400 41.830 321.900 ;
        RECT 42.030 321.400 42.580 321.900 ;
        RECT 66.830 338.100 67.430 338.600 ;
        RECT 67.630 338.100 68.230 338.600 ;
        RECT 68.430 338.100 69.030 338.600 ;
        RECT 69.230 338.100 69.830 338.600 ;
        RECT 70.030 338.100 70.630 338.600 ;
        RECT 78.830 338.100 79.430 338.600 ;
        RECT 79.630 338.100 80.230 338.600 ;
        RECT 80.430 338.100 81.030 338.600 ;
        RECT 81.230 338.100 81.830 338.600 ;
        RECT 82.030 338.100 82.580 338.600 ;
        RECT 46.830 321.400 47.430 321.900 ;
        RECT 47.630 321.400 48.230 321.900 ;
        RECT 48.430 321.400 49.030 321.900 ;
        RECT 49.230 321.400 49.830 321.900 ;
        RECT 50.030 321.400 50.630 321.900 ;
        RECT 58.830 321.400 59.430 321.900 ;
        RECT 59.630 321.400 60.230 321.900 ;
        RECT 60.430 321.400 61.030 321.900 ;
        RECT 61.230 321.400 61.830 321.900 ;
        RECT 62.030 321.400 62.580 321.900 ;
        RECT 86.830 338.100 87.430 338.600 ;
        RECT 87.630 338.100 88.230 338.600 ;
        RECT 88.430 338.100 89.030 338.600 ;
        RECT 89.230 338.100 89.830 338.600 ;
        RECT 90.030 338.100 90.630 338.600 ;
        RECT 98.830 338.100 99.430 338.600 ;
        RECT 99.630 338.100 100.230 338.600 ;
        RECT 100.430 338.100 101.030 338.600 ;
        RECT 101.230 338.100 101.830 338.600 ;
        RECT 102.030 338.100 102.580 338.600 ;
        RECT 66.830 321.400 67.430 321.900 ;
        RECT 67.630 321.400 68.230 321.900 ;
        RECT 68.430 321.400 69.030 321.900 ;
        RECT 69.230 321.400 69.830 321.900 ;
        RECT 70.030 321.400 70.630 321.900 ;
        RECT 78.830 321.400 79.430 321.900 ;
        RECT 79.630 321.400 80.230 321.900 ;
        RECT 80.430 321.400 81.030 321.900 ;
        RECT 81.230 321.400 81.830 321.900 ;
        RECT 82.030 321.400 82.580 321.900 ;
        RECT 86.830 321.400 87.430 321.900 ;
        RECT 87.630 321.400 88.230 321.900 ;
        RECT 88.430 321.400 89.030 321.900 ;
        RECT 89.230 321.400 89.830 321.900 ;
        RECT 90.030 321.400 90.630 321.900 ;
        RECT 98.830 321.400 99.430 321.900 ;
        RECT 99.630 321.400 100.230 321.900 ;
        RECT 100.430 321.400 101.030 321.900 ;
        RECT 101.230 321.400 101.830 321.900 ;
        RECT 102.030 321.400 102.580 321.900 ;
        RECT 6.830 318.100 7.430 318.600 ;
        RECT 7.630 318.100 8.230 318.600 ;
        RECT 8.430 318.100 9.030 318.600 ;
        RECT 9.230 318.100 9.830 318.600 ;
        RECT 10.030 318.100 10.630 318.600 ;
        RECT 18.830 318.100 19.430 318.600 ;
        RECT 19.630 318.100 20.230 318.600 ;
        RECT 20.430 318.100 21.030 318.600 ;
        RECT 21.230 318.100 21.830 318.600 ;
        RECT 22.030 318.100 22.580 318.600 ;
        RECT 2.520 314.920 2.880 315.300 ;
        RECT 3.130 314.920 3.490 315.300 ;
        RECT 3.760 314.920 4.120 315.300 ;
        RECT 2.520 314.185 2.880 314.565 ;
        RECT 3.130 314.185 3.490 314.565 ;
        RECT 3.760 314.185 4.120 314.565 ;
        RECT 2.520 313.500 2.880 313.880 ;
        RECT 3.130 313.500 3.490 313.880 ;
        RECT 3.760 313.500 4.120 313.880 ;
        RECT 2.520 306.125 2.880 306.505 ;
        RECT 3.130 306.125 3.490 306.505 ;
        RECT 3.760 306.125 4.120 306.505 ;
        RECT 2.520 305.390 2.880 305.770 ;
        RECT 3.130 305.390 3.490 305.770 ;
        RECT 3.760 305.390 4.120 305.770 ;
        RECT 2.520 304.705 2.880 305.085 ;
        RECT 3.130 304.705 3.490 305.085 ;
        RECT 3.760 304.705 4.120 305.085 ;
        RECT 26.830 318.100 27.430 318.600 ;
        RECT 27.630 318.100 28.230 318.600 ;
        RECT 28.430 318.100 29.030 318.600 ;
        RECT 29.230 318.100 29.830 318.600 ;
        RECT 30.030 318.100 30.630 318.600 ;
        RECT 38.830 318.100 39.430 318.600 ;
        RECT 39.630 318.100 40.230 318.600 ;
        RECT 40.430 318.100 41.030 318.600 ;
        RECT 41.230 318.100 41.830 318.600 ;
        RECT 42.030 318.100 42.580 318.600 ;
        RECT 6.830 301.400 7.430 301.900 ;
        RECT 7.630 301.400 8.230 301.900 ;
        RECT 8.430 301.400 9.030 301.900 ;
        RECT 9.230 301.400 9.830 301.900 ;
        RECT 10.030 301.400 10.630 301.900 ;
        RECT 18.830 301.400 19.430 301.900 ;
        RECT 19.630 301.400 20.230 301.900 ;
        RECT 20.430 301.400 21.030 301.900 ;
        RECT 21.230 301.400 21.830 301.900 ;
        RECT 22.030 301.400 22.580 301.900 ;
        RECT 46.830 318.100 47.430 318.600 ;
        RECT 47.630 318.100 48.230 318.600 ;
        RECT 48.430 318.100 49.030 318.600 ;
        RECT 49.230 318.100 49.830 318.600 ;
        RECT 50.030 318.100 50.630 318.600 ;
        RECT 58.830 318.100 59.430 318.600 ;
        RECT 59.630 318.100 60.230 318.600 ;
        RECT 60.430 318.100 61.030 318.600 ;
        RECT 61.230 318.100 61.830 318.600 ;
        RECT 62.030 318.100 62.580 318.600 ;
        RECT 26.830 301.400 27.430 301.900 ;
        RECT 27.630 301.400 28.230 301.900 ;
        RECT 28.430 301.400 29.030 301.900 ;
        RECT 29.230 301.400 29.830 301.900 ;
        RECT 30.030 301.400 30.630 301.900 ;
        RECT 38.830 301.400 39.430 301.900 ;
        RECT 39.630 301.400 40.230 301.900 ;
        RECT 40.430 301.400 41.030 301.900 ;
        RECT 41.230 301.400 41.830 301.900 ;
        RECT 42.030 301.400 42.580 301.900 ;
        RECT 66.830 318.100 67.430 318.600 ;
        RECT 67.630 318.100 68.230 318.600 ;
        RECT 68.430 318.100 69.030 318.600 ;
        RECT 69.230 318.100 69.830 318.600 ;
        RECT 70.030 318.100 70.630 318.600 ;
        RECT 78.830 318.100 79.430 318.600 ;
        RECT 79.630 318.100 80.230 318.600 ;
        RECT 80.430 318.100 81.030 318.600 ;
        RECT 81.230 318.100 81.830 318.600 ;
        RECT 82.030 318.100 82.580 318.600 ;
        RECT 46.830 301.400 47.430 301.900 ;
        RECT 47.630 301.400 48.230 301.900 ;
        RECT 48.430 301.400 49.030 301.900 ;
        RECT 49.230 301.400 49.830 301.900 ;
        RECT 50.030 301.400 50.630 301.900 ;
        RECT 58.830 301.400 59.430 301.900 ;
        RECT 59.630 301.400 60.230 301.900 ;
        RECT 60.430 301.400 61.030 301.900 ;
        RECT 61.230 301.400 61.830 301.900 ;
        RECT 62.030 301.400 62.580 301.900 ;
        RECT 86.830 318.100 87.430 318.600 ;
        RECT 87.630 318.100 88.230 318.600 ;
        RECT 88.430 318.100 89.030 318.600 ;
        RECT 89.230 318.100 89.830 318.600 ;
        RECT 90.030 318.100 90.630 318.600 ;
        RECT 98.830 318.100 99.430 318.600 ;
        RECT 99.630 318.100 100.230 318.600 ;
        RECT 100.430 318.100 101.030 318.600 ;
        RECT 101.230 318.100 101.830 318.600 ;
        RECT 102.030 318.100 102.580 318.600 ;
        RECT 66.830 301.400 67.430 301.900 ;
        RECT 67.630 301.400 68.230 301.900 ;
        RECT 68.430 301.400 69.030 301.900 ;
        RECT 69.230 301.400 69.830 301.900 ;
        RECT 70.030 301.400 70.630 301.900 ;
        RECT 78.830 301.400 79.430 301.900 ;
        RECT 79.630 301.400 80.230 301.900 ;
        RECT 80.430 301.400 81.030 301.900 ;
        RECT 81.230 301.400 81.830 301.900 ;
        RECT 82.030 301.400 82.580 301.900 ;
        RECT 86.830 301.400 87.430 301.900 ;
        RECT 87.630 301.400 88.230 301.900 ;
        RECT 88.430 301.400 89.030 301.900 ;
        RECT 89.230 301.400 89.830 301.900 ;
        RECT 90.030 301.400 90.630 301.900 ;
        RECT 98.830 301.400 99.430 301.900 ;
        RECT 99.630 301.400 100.230 301.900 ;
        RECT 100.430 301.400 101.030 301.900 ;
        RECT 101.230 301.400 101.830 301.900 ;
        RECT 102.030 301.400 102.580 301.900 ;
        RECT 6.830 298.100 7.430 298.600 ;
        RECT 7.630 298.100 8.230 298.600 ;
        RECT 8.430 298.100 9.030 298.600 ;
        RECT 9.230 298.100 9.830 298.600 ;
        RECT 10.030 298.100 10.630 298.600 ;
        RECT 18.830 298.100 19.430 298.600 ;
        RECT 19.630 298.100 20.230 298.600 ;
        RECT 20.430 298.100 21.030 298.600 ;
        RECT 21.230 298.100 21.830 298.600 ;
        RECT 22.030 298.100 22.580 298.600 ;
        RECT 2.520 294.920 2.880 295.300 ;
        RECT 3.130 294.920 3.490 295.300 ;
        RECT 3.760 294.920 4.120 295.300 ;
        RECT 2.520 294.185 2.880 294.565 ;
        RECT 3.130 294.185 3.490 294.565 ;
        RECT 3.760 294.185 4.120 294.565 ;
        RECT 2.520 293.500 2.880 293.880 ;
        RECT 3.130 293.500 3.490 293.880 ;
        RECT 3.760 293.500 4.120 293.880 ;
        RECT 2.520 286.115 2.880 286.495 ;
        RECT 3.130 286.115 3.490 286.495 ;
        RECT 3.760 286.115 4.120 286.495 ;
        RECT 2.520 285.380 2.880 285.760 ;
        RECT 3.130 285.380 3.490 285.760 ;
        RECT 3.760 285.380 4.120 285.760 ;
        RECT 2.520 284.695 2.880 285.075 ;
        RECT 3.130 284.695 3.490 285.075 ;
        RECT 3.760 284.695 4.120 285.075 ;
        RECT 26.830 298.100 27.430 298.600 ;
        RECT 27.630 298.100 28.230 298.600 ;
        RECT 28.430 298.100 29.030 298.600 ;
        RECT 29.230 298.100 29.830 298.600 ;
        RECT 30.030 298.100 30.630 298.600 ;
        RECT 38.830 298.100 39.430 298.600 ;
        RECT 39.630 298.100 40.230 298.600 ;
        RECT 40.430 298.100 41.030 298.600 ;
        RECT 41.230 298.100 41.830 298.600 ;
        RECT 42.030 298.100 42.580 298.600 ;
        RECT 6.830 281.400 7.430 281.900 ;
        RECT 7.630 281.400 8.230 281.900 ;
        RECT 8.430 281.400 9.030 281.900 ;
        RECT 9.230 281.400 9.830 281.900 ;
        RECT 10.030 281.400 10.630 281.900 ;
        RECT 18.830 281.400 19.430 281.900 ;
        RECT 19.630 281.400 20.230 281.900 ;
        RECT 20.430 281.400 21.030 281.900 ;
        RECT 21.230 281.400 21.830 281.900 ;
        RECT 22.030 281.400 22.580 281.900 ;
        RECT 46.830 298.100 47.430 298.600 ;
        RECT 47.630 298.100 48.230 298.600 ;
        RECT 48.430 298.100 49.030 298.600 ;
        RECT 49.230 298.100 49.830 298.600 ;
        RECT 50.030 298.100 50.630 298.600 ;
        RECT 58.830 298.100 59.430 298.600 ;
        RECT 59.630 298.100 60.230 298.600 ;
        RECT 60.430 298.100 61.030 298.600 ;
        RECT 61.230 298.100 61.830 298.600 ;
        RECT 62.030 298.100 62.580 298.600 ;
        RECT 26.830 281.400 27.430 281.900 ;
        RECT 27.630 281.400 28.230 281.900 ;
        RECT 28.430 281.400 29.030 281.900 ;
        RECT 29.230 281.400 29.830 281.900 ;
        RECT 30.030 281.400 30.630 281.900 ;
        RECT 38.830 281.400 39.430 281.900 ;
        RECT 39.630 281.400 40.230 281.900 ;
        RECT 40.430 281.400 41.030 281.900 ;
        RECT 41.230 281.400 41.830 281.900 ;
        RECT 42.030 281.400 42.580 281.900 ;
        RECT 66.830 298.100 67.430 298.600 ;
        RECT 67.630 298.100 68.230 298.600 ;
        RECT 68.430 298.100 69.030 298.600 ;
        RECT 69.230 298.100 69.830 298.600 ;
        RECT 70.030 298.100 70.630 298.600 ;
        RECT 78.830 298.100 79.430 298.600 ;
        RECT 79.630 298.100 80.230 298.600 ;
        RECT 80.430 298.100 81.030 298.600 ;
        RECT 81.230 298.100 81.830 298.600 ;
        RECT 82.030 298.100 82.580 298.600 ;
        RECT 46.830 281.400 47.430 281.900 ;
        RECT 47.630 281.400 48.230 281.900 ;
        RECT 48.430 281.400 49.030 281.900 ;
        RECT 49.230 281.400 49.830 281.900 ;
        RECT 50.030 281.400 50.630 281.900 ;
        RECT 58.830 281.400 59.430 281.900 ;
        RECT 59.630 281.400 60.230 281.900 ;
        RECT 60.430 281.400 61.030 281.900 ;
        RECT 61.230 281.400 61.830 281.900 ;
        RECT 62.030 281.400 62.580 281.900 ;
        RECT 86.830 298.100 87.430 298.600 ;
        RECT 87.630 298.100 88.230 298.600 ;
        RECT 88.430 298.100 89.030 298.600 ;
        RECT 89.230 298.100 89.830 298.600 ;
        RECT 90.030 298.100 90.630 298.600 ;
        RECT 98.830 298.100 99.430 298.600 ;
        RECT 99.630 298.100 100.230 298.600 ;
        RECT 100.430 298.100 101.030 298.600 ;
        RECT 101.230 298.100 101.830 298.600 ;
        RECT 102.030 298.100 102.580 298.600 ;
        RECT 66.830 281.400 67.430 281.900 ;
        RECT 67.630 281.400 68.230 281.900 ;
        RECT 68.430 281.400 69.030 281.900 ;
        RECT 69.230 281.400 69.830 281.900 ;
        RECT 70.030 281.400 70.630 281.900 ;
        RECT 78.830 281.400 79.430 281.900 ;
        RECT 79.630 281.400 80.230 281.900 ;
        RECT 80.430 281.400 81.030 281.900 ;
        RECT 81.230 281.400 81.830 281.900 ;
        RECT 82.030 281.400 82.580 281.900 ;
        RECT 86.830 281.400 87.430 281.900 ;
        RECT 87.630 281.400 88.230 281.900 ;
        RECT 88.430 281.400 89.030 281.900 ;
        RECT 89.230 281.400 89.830 281.900 ;
        RECT 90.030 281.400 90.630 281.900 ;
        RECT 98.830 281.400 99.430 281.900 ;
        RECT 99.630 281.400 100.230 281.900 ;
        RECT 100.430 281.400 101.030 281.900 ;
        RECT 101.230 281.400 101.830 281.900 ;
        RECT 102.030 281.400 102.580 281.900 ;
        RECT 6.830 278.100 7.430 278.600 ;
        RECT 7.630 278.100 8.230 278.600 ;
        RECT 8.430 278.100 9.030 278.600 ;
        RECT 9.230 278.100 9.830 278.600 ;
        RECT 10.030 278.100 10.630 278.600 ;
        RECT 18.830 278.100 19.430 278.600 ;
        RECT 19.630 278.100 20.230 278.600 ;
        RECT 20.430 278.100 21.030 278.600 ;
        RECT 21.230 278.100 21.830 278.600 ;
        RECT 22.030 278.100 22.580 278.600 ;
        RECT 2.520 274.920 2.880 275.300 ;
        RECT 3.130 274.920 3.490 275.300 ;
        RECT 3.760 274.920 4.120 275.300 ;
        RECT 2.520 274.185 2.880 274.565 ;
        RECT 3.130 274.185 3.490 274.565 ;
        RECT 3.760 274.185 4.120 274.565 ;
        RECT 2.520 273.500 2.880 273.880 ;
        RECT 3.130 273.500 3.490 273.880 ;
        RECT 3.760 273.500 4.120 273.880 ;
        RECT 2.520 266.125 2.880 266.505 ;
        RECT 3.130 266.125 3.490 266.505 ;
        RECT 3.760 266.125 4.120 266.505 ;
        RECT 2.520 265.390 2.880 265.770 ;
        RECT 3.130 265.390 3.490 265.770 ;
        RECT 3.760 265.390 4.120 265.770 ;
        RECT 2.520 264.705 2.880 265.085 ;
        RECT 3.130 264.705 3.490 265.085 ;
        RECT 3.760 264.705 4.120 265.085 ;
        RECT 26.830 278.100 27.430 278.600 ;
        RECT 27.630 278.100 28.230 278.600 ;
        RECT 28.430 278.100 29.030 278.600 ;
        RECT 29.230 278.100 29.830 278.600 ;
        RECT 30.030 278.100 30.630 278.600 ;
        RECT 38.830 278.100 39.430 278.600 ;
        RECT 39.630 278.100 40.230 278.600 ;
        RECT 40.430 278.100 41.030 278.600 ;
        RECT 41.230 278.100 41.830 278.600 ;
        RECT 42.030 278.100 42.580 278.600 ;
        RECT 6.830 261.400 7.430 261.900 ;
        RECT 7.630 261.400 8.230 261.900 ;
        RECT 8.430 261.400 9.030 261.900 ;
        RECT 9.230 261.400 9.830 261.900 ;
        RECT 10.030 261.400 10.630 261.900 ;
        RECT 18.830 261.400 19.430 261.900 ;
        RECT 19.630 261.400 20.230 261.900 ;
        RECT 20.430 261.400 21.030 261.900 ;
        RECT 21.230 261.400 21.830 261.900 ;
        RECT 22.030 261.400 22.580 261.900 ;
        RECT 46.830 278.100 47.430 278.600 ;
        RECT 47.630 278.100 48.230 278.600 ;
        RECT 48.430 278.100 49.030 278.600 ;
        RECT 49.230 278.100 49.830 278.600 ;
        RECT 50.030 278.100 50.630 278.600 ;
        RECT 58.830 278.100 59.430 278.600 ;
        RECT 59.630 278.100 60.230 278.600 ;
        RECT 60.430 278.100 61.030 278.600 ;
        RECT 61.230 278.100 61.830 278.600 ;
        RECT 62.030 278.100 62.580 278.600 ;
        RECT 26.830 261.400 27.430 261.900 ;
        RECT 27.630 261.400 28.230 261.900 ;
        RECT 28.430 261.400 29.030 261.900 ;
        RECT 29.230 261.400 29.830 261.900 ;
        RECT 30.030 261.400 30.630 261.900 ;
        RECT 38.830 261.400 39.430 261.900 ;
        RECT 39.630 261.400 40.230 261.900 ;
        RECT 40.430 261.400 41.030 261.900 ;
        RECT 41.230 261.400 41.830 261.900 ;
        RECT 42.030 261.400 42.580 261.900 ;
        RECT 66.830 278.100 67.430 278.600 ;
        RECT 67.630 278.100 68.230 278.600 ;
        RECT 68.430 278.100 69.030 278.600 ;
        RECT 69.230 278.100 69.830 278.600 ;
        RECT 70.030 278.100 70.630 278.600 ;
        RECT 78.830 278.100 79.430 278.600 ;
        RECT 79.630 278.100 80.230 278.600 ;
        RECT 80.430 278.100 81.030 278.600 ;
        RECT 81.230 278.100 81.830 278.600 ;
        RECT 82.030 278.100 82.580 278.600 ;
        RECT 46.830 261.400 47.430 261.900 ;
        RECT 47.630 261.400 48.230 261.900 ;
        RECT 48.430 261.400 49.030 261.900 ;
        RECT 49.230 261.400 49.830 261.900 ;
        RECT 50.030 261.400 50.630 261.900 ;
        RECT 58.830 261.400 59.430 261.900 ;
        RECT 59.630 261.400 60.230 261.900 ;
        RECT 60.430 261.400 61.030 261.900 ;
        RECT 61.230 261.400 61.830 261.900 ;
        RECT 62.030 261.400 62.580 261.900 ;
        RECT 86.830 278.100 87.430 278.600 ;
        RECT 87.630 278.100 88.230 278.600 ;
        RECT 88.430 278.100 89.030 278.600 ;
        RECT 89.230 278.100 89.830 278.600 ;
        RECT 90.030 278.100 90.630 278.600 ;
        RECT 98.830 278.100 99.430 278.600 ;
        RECT 99.630 278.100 100.230 278.600 ;
        RECT 100.430 278.100 101.030 278.600 ;
        RECT 101.230 278.100 101.830 278.600 ;
        RECT 102.030 278.100 102.580 278.600 ;
        RECT 66.830 261.400 67.430 261.900 ;
        RECT 67.630 261.400 68.230 261.900 ;
        RECT 68.430 261.400 69.030 261.900 ;
        RECT 69.230 261.400 69.830 261.900 ;
        RECT 70.030 261.400 70.630 261.900 ;
        RECT 78.830 261.400 79.430 261.900 ;
        RECT 79.630 261.400 80.230 261.900 ;
        RECT 80.430 261.400 81.030 261.900 ;
        RECT 81.230 261.400 81.830 261.900 ;
        RECT 82.030 261.400 82.580 261.900 ;
        RECT 86.830 261.400 87.430 261.900 ;
        RECT 87.630 261.400 88.230 261.900 ;
        RECT 88.430 261.400 89.030 261.900 ;
        RECT 89.230 261.400 89.830 261.900 ;
        RECT 90.030 261.400 90.630 261.900 ;
        RECT 98.830 261.400 99.430 261.900 ;
        RECT 99.630 261.400 100.230 261.900 ;
        RECT 100.430 261.400 101.030 261.900 ;
        RECT 101.230 261.400 101.830 261.900 ;
        RECT 102.030 261.400 102.580 261.900 ;
        RECT 6.830 258.100 7.430 258.600 ;
        RECT 7.630 258.100 8.230 258.600 ;
        RECT 8.430 258.100 9.030 258.600 ;
        RECT 9.230 258.100 9.830 258.600 ;
        RECT 10.030 258.100 10.630 258.600 ;
        RECT 18.830 258.100 19.430 258.600 ;
        RECT 19.630 258.100 20.230 258.600 ;
        RECT 20.430 258.100 21.030 258.600 ;
        RECT 21.230 258.100 21.830 258.600 ;
        RECT 22.030 258.100 22.580 258.600 ;
        RECT 2.520 254.920 2.880 255.300 ;
        RECT 3.130 254.920 3.490 255.300 ;
        RECT 3.760 254.920 4.120 255.300 ;
        RECT 2.520 254.185 2.880 254.565 ;
        RECT 3.130 254.185 3.490 254.565 ;
        RECT 3.760 254.185 4.120 254.565 ;
        RECT 2.520 253.500 2.880 253.880 ;
        RECT 3.130 253.500 3.490 253.880 ;
        RECT 3.760 253.500 4.120 253.880 ;
        RECT 2.520 246.125 2.880 246.505 ;
        RECT 3.130 246.125 3.490 246.505 ;
        RECT 3.760 246.125 4.120 246.505 ;
        RECT 2.520 245.390 2.880 245.770 ;
        RECT 3.130 245.390 3.490 245.770 ;
        RECT 3.760 245.390 4.120 245.770 ;
        RECT 2.520 244.705 2.880 245.085 ;
        RECT 3.130 244.705 3.490 245.085 ;
        RECT 3.760 244.705 4.120 245.085 ;
        RECT 26.830 258.100 27.430 258.600 ;
        RECT 27.630 258.100 28.230 258.600 ;
        RECT 28.430 258.100 29.030 258.600 ;
        RECT 29.230 258.100 29.830 258.600 ;
        RECT 30.030 258.100 30.630 258.600 ;
        RECT 38.830 258.100 39.430 258.600 ;
        RECT 39.630 258.100 40.230 258.600 ;
        RECT 40.430 258.100 41.030 258.600 ;
        RECT 41.230 258.100 41.830 258.600 ;
        RECT 42.030 258.100 42.580 258.600 ;
        RECT 6.830 241.400 7.430 241.900 ;
        RECT 7.630 241.400 8.230 241.900 ;
        RECT 8.430 241.400 9.030 241.900 ;
        RECT 9.230 241.400 9.830 241.900 ;
        RECT 10.030 241.400 10.630 241.900 ;
        RECT 18.830 241.400 19.430 241.900 ;
        RECT 19.630 241.400 20.230 241.900 ;
        RECT 20.430 241.400 21.030 241.900 ;
        RECT 21.230 241.400 21.830 241.900 ;
        RECT 22.030 241.400 22.580 241.900 ;
        RECT 46.830 258.100 47.430 258.600 ;
        RECT 47.630 258.100 48.230 258.600 ;
        RECT 48.430 258.100 49.030 258.600 ;
        RECT 49.230 258.100 49.830 258.600 ;
        RECT 50.030 258.100 50.630 258.600 ;
        RECT 58.830 258.100 59.430 258.600 ;
        RECT 59.630 258.100 60.230 258.600 ;
        RECT 60.430 258.100 61.030 258.600 ;
        RECT 61.230 258.100 61.830 258.600 ;
        RECT 62.030 258.100 62.580 258.600 ;
        RECT 26.830 241.400 27.430 241.900 ;
        RECT 27.630 241.400 28.230 241.900 ;
        RECT 28.430 241.400 29.030 241.900 ;
        RECT 29.230 241.400 29.830 241.900 ;
        RECT 30.030 241.400 30.630 241.900 ;
        RECT 38.830 241.400 39.430 241.900 ;
        RECT 39.630 241.400 40.230 241.900 ;
        RECT 40.430 241.400 41.030 241.900 ;
        RECT 41.230 241.400 41.830 241.900 ;
        RECT 42.030 241.400 42.580 241.900 ;
        RECT 66.830 258.100 67.430 258.600 ;
        RECT 67.630 258.100 68.230 258.600 ;
        RECT 68.430 258.100 69.030 258.600 ;
        RECT 69.230 258.100 69.830 258.600 ;
        RECT 70.030 258.100 70.630 258.600 ;
        RECT 78.830 258.100 79.430 258.600 ;
        RECT 79.630 258.100 80.230 258.600 ;
        RECT 80.430 258.100 81.030 258.600 ;
        RECT 81.230 258.100 81.830 258.600 ;
        RECT 82.030 258.100 82.580 258.600 ;
        RECT 46.830 241.400 47.430 241.900 ;
        RECT 47.630 241.400 48.230 241.900 ;
        RECT 48.430 241.400 49.030 241.900 ;
        RECT 49.230 241.400 49.830 241.900 ;
        RECT 50.030 241.400 50.630 241.900 ;
        RECT 58.830 241.400 59.430 241.900 ;
        RECT 59.630 241.400 60.230 241.900 ;
        RECT 60.430 241.400 61.030 241.900 ;
        RECT 61.230 241.400 61.830 241.900 ;
        RECT 62.030 241.400 62.580 241.900 ;
        RECT 86.830 258.100 87.430 258.600 ;
        RECT 87.630 258.100 88.230 258.600 ;
        RECT 88.430 258.100 89.030 258.600 ;
        RECT 89.230 258.100 89.830 258.600 ;
        RECT 90.030 258.100 90.630 258.600 ;
        RECT 98.830 258.100 99.430 258.600 ;
        RECT 99.630 258.100 100.230 258.600 ;
        RECT 100.430 258.100 101.030 258.600 ;
        RECT 101.230 258.100 101.830 258.600 ;
        RECT 102.030 258.100 102.580 258.600 ;
        RECT 66.830 241.400 67.430 241.900 ;
        RECT 67.630 241.400 68.230 241.900 ;
        RECT 68.430 241.400 69.030 241.900 ;
        RECT 69.230 241.400 69.830 241.900 ;
        RECT 70.030 241.400 70.630 241.900 ;
        RECT 78.830 241.400 79.430 241.900 ;
        RECT 79.630 241.400 80.230 241.900 ;
        RECT 80.430 241.400 81.030 241.900 ;
        RECT 81.230 241.400 81.830 241.900 ;
        RECT 82.030 241.400 82.580 241.900 ;
        RECT 86.830 241.400 87.430 241.900 ;
        RECT 87.630 241.400 88.230 241.900 ;
        RECT 88.430 241.400 89.030 241.900 ;
        RECT 89.230 241.400 89.830 241.900 ;
        RECT 90.030 241.400 90.630 241.900 ;
        RECT 98.830 241.400 99.430 241.900 ;
        RECT 99.630 241.400 100.230 241.900 ;
        RECT 100.430 241.400 101.030 241.900 ;
        RECT 101.230 241.400 101.830 241.900 ;
        RECT 102.030 241.400 102.580 241.900 ;
        RECT 6.830 238.100 7.430 238.600 ;
        RECT 7.630 238.100 8.230 238.600 ;
        RECT 8.430 238.100 9.030 238.600 ;
        RECT 9.230 238.100 9.830 238.600 ;
        RECT 10.030 238.100 10.630 238.600 ;
        RECT 18.830 238.100 19.430 238.600 ;
        RECT 19.630 238.100 20.230 238.600 ;
        RECT 20.430 238.100 21.030 238.600 ;
        RECT 21.230 238.100 21.830 238.600 ;
        RECT 22.030 238.100 22.580 238.600 ;
        RECT 2.520 234.920 2.880 235.300 ;
        RECT 3.130 234.920 3.490 235.300 ;
        RECT 3.760 234.920 4.120 235.300 ;
        RECT 2.520 234.185 2.880 234.565 ;
        RECT 3.130 234.185 3.490 234.565 ;
        RECT 3.760 234.185 4.120 234.565 ;
        RECT 2.520 233.500 2.880 233.880 ;
        RECT 3.130 233.500 3.490 233.880 ;
        RECT 3.760 233.500 4.120 233.880 ;
        RECT 2.520 226.120 2.880 226.500 ;
        RECT 3.130 226.120 3.490 226.500 ;
        RECT 3.760 226.120 4.120 226.500 ;
        RECT 2.520 225.385 2.880 225.765 ;
        RECT 3.130 225.385 3.490 225.765 ;
        RECT 3.760 225.385 4.120 225.765 ;
        RECT 2.520 224.700 2.880 225.080 ;
        RECT 3.130 224.700 3.490 225.080 ;
        RECT 3.760 224.700 4.120 225.080 ;
        RECT 26.830 238.100 27.430 238.600 ;
        RECT 27.630 238.100 28.230 238.600 ;
        RECT 28.430 238.100 29.030 238.600 ;
        RECT 29.230 238.100 29.830 238.600 ;
        RECT 30.030 238.100 30.630 238.600 ;
        RECT 38.830 238.100 39.430 238.600 ;
        RECT 39.630 238.100 40.230 238.600 ;
        RECT 40.430 238.100 41.030 238.600 ;
        RECT 41.230 238.100 41.830 238.600 ;
        RECT 42.030 238.100 42.580 238.600 ;
        RECT 6.830 221.400 7.430 221.900 ;
        RECT 7.630 221.400 8.230 221.900 ;
        RECT 8.430 221.400 9.030 221.900 ;
        RECT 9.230 221.400 9.830 221.900 ;
        RECT 10.030 221.400 10.630 221.900 ;
        RECT 18.830 221.400 19.430 221.900 ;
        RECT 19.630 221.400 20.230 221.900 ;
        RECT 20.430 221.400 21.030 221.900 ;
        RECT 21.230 221.400 21.830 221.900 ;
        RECT 22.030 221.400 22.580 221.900 ;
        RECT 46.830 238.100 47.430 238.600 ;
        RECT 47.630 238.100 48.230 238.600 ;
        RECT 48.430 238.100 49.030 238.600 ;
        RECT 49.230 238.100 49.830 238.600 ;
        RECT 50.030 238.100 50.630 238.600 ;
        RECT 58.830 238.100 59.430 238.600 ;
        RECT 59.630 238.100 60.230 238.600 ;
        RECT 60.430 238.100 61.030 238.600 ;
        RECT 61.230 238.100 61.830 238.600 ;
        RECT 62.030 238.100 62.580 238.600 ;
        RECT 26.830 221.400 27.430 221.900 ;
        RECT 27.630 221.400 28.230 221.900 ;
        RECT 28.430 221.400 29.030 221.900 ;
        RECT 29.230 221.400 29.830 221.900 ;
        RECT 30.030 221.400 30.630 221.900 ;
        RECT 38.830 221.400 39.430 221.900 ;
        RECT 39.630 221.400 40.230 221.900 ;
        RECT 40.430 221.400 41.030 221.900 ;
        RECT 41.230 221.400 41.830 221.900 ;
        RECT 42.030 221.400 42.580 221.900 ;
        RECT 66.830 238.100 67.430 238.600 ;
        RECT 67.630 238.100 68.230 238.600 ;
        RECT 68.430 238.100 69.030 238.600 ;
        RECT 69.230 238.100 69.830 238.600 ;
        RECT 70.030 238.100 70.630 238.600 ;
        RECT 78.830 238.100 79.430 238.600 ;
        RECT 79.630 238.100 80.230 238.600 ;
        RECT 80.430 238.100 81.030 238.600 ;
        RECT 81.230 238.100 81.830 238.600 ;
        RECT 82.030 238.100 82.580 238.600 ;
        RECT 46.830 221.400 47.430 221.900 ;
        RECT 47.630 221.400 48.230 221.900 ;
        RECT 48.430 221.400 49.030 221.900 ;
        RECT 49.230 221.400 49.830 221.900 ;
        RECT 50.030 221.400 50.630 221.900 ;
        RECT 58.830 221.400 59.430 221.900 ;
        RECT 59.630 221.400 60.230 221.900 ;
        RECT 60.430 221.400 61.030 221.900 ;
        RECT 61.230 221.400 61.830 221.900 ;
        RECT 62.030 221.400 62.580 221.900 ;
        RECT 86.830 238.100 87.430 238.600 ;
        RECT 87.630 238.100 88.230 238.600 ;
        RECT 88.430 238.100 89.030 238.600 ;
        RECT 89.230 238.100 89.830 238.600 ;
        RECT 90.030 238.100 90.630 238.600 ;
        RECT 98.830 238.100 99.430 238.600 ;
        RECT 99.630 238.100 100.230 238.600 ;
        RECT 100.430 238.100 101.030 238.600 ;
        RECT 101.230 238.100 101.830 238.600 ;
        RECT 102.030 238.100 102.580 238.600 ;
        RECT 66.830 221.400 67.430 221.900 ;
        RECT 67.630 221.400 68.230 221.900 ;
        RECT 68.430 221.400 69.030 221.900 ;
        RECT 69.230 221.400 69.830 221.900 ;
        RECT 70.030 221.400 70.630 221.900 ;
        RECT 78.830 221.400 79.430 221.900 ;
        RECT 79.630 221.400 80.230 221.900 ;
        RECT 80.430 221.400 81.030 221.900 ;
        RECT 81.230 221.400 81.830 221.900 ;
        RECT 82.030 221.400 82.580 221.900 ;
        RECT 86.830 221.400 87.430 221.900 ;
        RECT 87.630 221.400 88.230 221.900 ;
        RECT 88.430 221.400 89.030 221.900 ;
        RECT 89.230 221.400 89.830 221.900 ;
        RECT 90.030 221.400 90.630 221.900 ;
        RECT 98.830 221.400 99.430 221.900 ;
        RECT 99.630 221.400 100.230 221.900 ;
        RECT 100.430 221.400 101.030 221.900 ;
        RECT 101.230 221.400 101.830 221.900 ;
        RECT 102.030 221.400 102.580 221.900 ;
        RECT 4.705 195.310 5.065 195.685 ;
        RECT 5.490 195.315 5.825 195.690 ;
        RECT 7.085 195.375 7.255 195.545 ;
        RECT 4.720 194.730 5.080 195.105 ;
        RECT 5.490 194.745 5.825 195.120 ;
        RECT 8.020 195.295 8.190 195.625 ;
        RECT 9.600 195.345 9.770 195.620 ;
        RECT 15.010 195.370 15.180 195.540 ;
        RECT 15.470 195.370 15.640 195.540 ;
        RECT 15.930 195.370 16.100 195.540 ;
        RECT 16.390 195.370 16.560 195.540 ;
        RECT 16.850 195.370 17.020 195.540 ;
        RECT 17.310 195.370 17.480 195.540 ;
        RECT 17.770 195.370 17.940 195.540 ;
        RECT 18.230 195.370 18.400 195.540 ;
        RECT 18.690 195.370 18.860 195.540 ;
        RECT 19.150 195.370 19.320 195.540 ;
        RECT 19.610 195.370 19.780 195.540 ;
        RECT 20.070 195.370 20.240 195.540 ;
        RECT 20.530 195.370 20.700 195.540 ;
        RECT 20.990 195.370 21.160 195.540 ;
        RECT 21.450 195.370 21.620 195.540 ;
        RECT 21.910 195.370 22.080 195.540 ;
        RECT 22.370 195.370 22.540 195.540 ;
        RECT 22.830 195.370 23.000 195.540 ;
        RECT 23.290 195.370 23.460 195.540 ;
        RECT 8.020 194.445 8.190 194.720 ;
        RECT 9.600 194.445 9.770 194.720 ;
        RECT 6.730 189.930 6.900 190.100 ;
        RECT 7.190 189.930 7.360 190.100 ;
        RECT 7.650 189.930 7.820 190.100 ;
        RECT 8.110 189.930 8.280 190.100 ;
        RECT 8.570 189.930 8.740 190.100 ;
        RECT 9.030 189.930 9.200 190.100 ;
        RECT 9.490 189.930 9.660 190.100 ;
        RECT 9.950 189.930 10.120 190.100 ;
        RECT 10.410 189.930 10.580 190.100 ;
        RECT 10.870 189.930 11.040 190.100 ;
        RECT 11.330 189.930 11.500 190.100 ;
        RECT 11.790 189.930 11.960 190.100 ;
        RECT 12.250 189.930 12.420 190.100 ;
        RECT 12.710 189.930 12.880 190.100 ;
        RECT 13.170 189.930 13.340 190.100 ;
        RECT 13.630 189.930 13.800 190.100 ;
        RECT 14.090 189.930 14.260 190.100 ;
        RECT 14.550 189.930 14.720 190.100 ;
        RECT 15.010 189.930 15.180 190.100 ;
        RECT 15.470 189.930 15.640 190.100 ;
        RECT 15.930 189.930 16.100 190.100 ;
        RECT 16.390 189.930 16.560 190.100 ;
        RECT 16.850 189.930 17.020 190.100 ;
        RECT 17.310 189.930 17.480 190.100 ;
        RECT 17.770 189.930 17.940 190.100 ;
        RECT 18.230 189.930 18.400 190.100 ;
        RECT 18.690 189.930 18.860 190.100 ;
        RECT 19.150 189.930 19.320 190.100 ;
        RECT 19.610 189.930 19.780 190.100 ;
        RECT 20.070 189.930 20.240 190.100 ;
        RECT 20.530 189.930 20.700 190.100 ;
        RECT 20.990 189.930 21.160 190.100 ;
        RECT 21.450 189.930 21.620 190.100 ;
        RECT 21.910 189.930 22.080 190.100 ;
        RECT 22.370 189.930 22.540 190.100 ;
        RECT 22.830 189.930 23.000 190.100 ;
        RECT 23.290 189.930 23.460 190.100 ;
        RECT 23.750 189.930 23.920 190.100 ;
        RECT 4.735 184.955 5.210 185.395 ;
        RECT 5.400 184.955 5.825 185.395 ;
        RECT 4.735 184.305 5.210 184.745 ;
        RECT 5.405 184.305 5.825 184.745 ;
        RECT 7.650 184.490 7.820 184.660 ;
        RECT 15.010 184.490 15.180 184.660 ;
        RECT 15.470 184.490 15.640 184.660 ;
        RECT 15.930 184.490 16.100 184.660 ;
        RECT 16.390 184.490 16.560 184.660 ;
        RECT 16.850 184.490 17.020 184.660 ;
        RECT 17.310 184.490 17.480 184.660 ;
        RECT 17.770 184.490 17.940 184.660 ;
        RECT 18.230 184.490 18.400 184.660 ;
        RECT 18.690 184.490 18.860 184.660 ;
        RECT 19.150 184.490 19.320 184.660 ;
        RECT 19.610 184.490 19.780 184.660 ;
        RECT 20.070 184.490 20.240 184.660 ;
        RECT 20.530 184.490 20.700 184.660 ;
        RECT 20.990 184.490 21.160 184.660 ;
        RECT 21.450 184.490 21.620 184.660 ;
        RECT 21.910 184.490 22.080 184.660 ;
        RECT 22.370 184.490 22.540 184.660 ;
        RECT 22.830 184.490 23.000 184.660 ;
        RECT 23.290 184.490 23.460 184.660 ;
        RECT 44.735 180.760 45.335 181.260 ;
        RECT 45.535 180.760 46.135 181.260 ;
        RECT 46.335 180.760 46.935 181.260 ;
        RECT 47.135 180.760 47.735 181.260 ;
        RECT 47.935 180.760 48.535 181.260 ;
        RECT 56.735 180.760 57.335 181.260 ;
        RECT 57.535 180.760 58.135 181.260 ;
        RECT 58.335 180.760 58.935 181.260 ;
        RECT 59.135 180.760 59.735 181.260 ;
        RECT 59.935 180.760 60.485 181.260 ;
        RECT 64.735 180.760 65.335 181.260 ;
        RECT 65.535 180.760 66.135 181.260 ;
        RECT 66.335 180.760 66.935 181.260 ;
        RECT 67.135 180.760 67.735 181.260 ;
        RECT 67.935 180.760 68.535 181.260 ;
        RECT 76.735 180.760 77.335 181.260 ;
        RECT 77.535 180.760 78.135 181.260 ;
        RECT 78.335 180.760 78.935 181.260 ;
        RECT 79.135 180.760 79.735 181.260 ;
        RECT 79.935 180.760 80.485 181.260 ;
        RECT 44.735 164.060 45.335 164.560 ;
        RECT 45.535 164.060 46.135 164.560 ;
        RECT 46.335 164.060 46.935 164.560 ;
        RECT 47.135 164.060 47.735 164.560 ;
        RECT 47.935 164.060 48.535 164.560 ;
        RECT 56.735 164.060 57.335 164.560 ;
        RECT 57.535 164.060 58.135 164.560 ;
        RECT 58.335 164.060 58.935 164.560 ;
        RECT 59.135 164.060 59.735 164.560 ;
        RECT 59.935 164.060 60.485 164.560 ;
        RECT 84.735 180.760 85.335 181.260 ;
        RECT 85.535 180.760 86.135 181.260 ;
        RECT 86.335 180.760 86.935 181.260 ;
        RECT 87.135 180.760 87.735 181.260 ;
        RECT 87.935 180.760 88.535 181.260 ;
        RECT 96.735 180.760 97.335 181.260 ;
        RECT 97.535 180.760 98.135 181.260 ;
        RECT 98.335 180.760 98.935 181.260 ;
        RECT 99.135 180.760 99.735 181.260 ;
        RECT 99.935 180.760 100.485 181.260 ;
        RECT 64.735 164.060 65.335 164.560 ;
        RECT 65.535 164.060 66.135 164.560 ;
        RECT 66.335 164.060 66.935 164.560 ;
        RECT 67.135 164.060 67.735 164.560 ;
        RECT 67.935 164.060 68.535 164.560 ;
        RECT 76.735 164.060 77.335 164.560 ;
        RECT 77.535 164.060 78.135 164.560 ;
        RECT 78.335 164.060 78.935 164.560 ;
        RECT 79.135 164.060 79.735 164.560 ;
        RECT 79.935 164.060 80.485 164.560 ;
        RECT 105.345 177.580 105.705 177.960 ;
        RECT 105.955 177.580 106.315 177.960 ;
        RECT 106.585 177.580 106.945 177.960 ;
        RECT 105.345 176.845 105.705 177.225 ;
        RECT 105.955 176.845 106.315 177.225 ;
        RECT 106.585 176.845 106.945 177.225 ;
        RECT 105.345 176.160 105.705 176.540 ;
        RECT 105.955 176.160 106.315 176.540 ;
        RECT 106.585 176.160 106.945 176.540 ;
        RECT 105.345 168.780 105.705 169.160 ;
        RECT 105.955 168.780 106.315 169.160 ;
        RECT 106.585 168.780 106.945 169.160 ;
        RECT 105.345 168.045 105.705 168.425 ;
        RECT 105.955 168.045 106.315 168.425 ;
        RECT 106.585 168.045 106.945 168.425 ;
        RECT 105.345 167.360 105.705 167.740 ;
        RECT 105.955 167.360 106.315 167.740 ;
        RECT 106.585 167.360 106.945 167.740 ;
        RECT 84.735 164.060 85.335 164.560 ;
        RECT 85.535 164.060 86.135 164.560 ;
        RECT 86.335 164.060 86.935 164.560 ;
        RECT 87.135 164.060 87.735 164.560 ;
        RECT 87.935 164.060 88.535 164.560 ;
        RECT 96.735 164.060 97.335 164.560 ;
        RECT 97.535 164.060 98.135 164.560 ;
        RECT 98.335 164.060 98.935 164.560 ;
        RECT 99.135 164.060 99.735 164.560 ;
        RECT 99.935 164.060 100.485 164.560 ;
        RECT 6.830 158.100 7.430 158.600 ;
        RECT 7.630 158.100 8.230 158.600 ;
        RECT 8.430 158.100 9.030 158.600 ;
        RECT 9.230 158.100 9.830 158.600 ;
        RECT 10.030 158.100 10.630 158.600 ;
        RECT 18.830 158.100 19.430 158.600 ;
        RECT 19.630 158.100 20.230 158.600 ;
        RECT 20.430 158.100 21.030 158.600 ;
        RECT 21.230 158.100 21.830 158.600 ;
        RECT 22.030 158.100 22.580 158.600 ;
        RECT 2.520 154.925 2.880 155.305 ;
        RECT 3.130 154.925 3.490 155.305 ;
        RECT 3.760 154.925 4.120 155.305 ;
        RECT 2.520 154.190 2.880 154.570 ;
        RECT 3.130 154.190 3.490 154.570 ;
        RECT 3.760 154.190 4.120 154.570 ;
        RECT 2.520 153.505 2.880 153.885 ;
        RECT 3.130 153.505 3.490 153.885 ;
        RECT 3.760 153.505 4.120 153.885 ;
        RECT 2.520 146.090 2.880 146.470 ;
        RECT 3.130 146.090 3.490 146.470 ;
        RECT 3.760 146.090 4.120 146.470 ;
        RECT 2.520 145.355 2.880 145.735 ;
        RECT 3.130 145.355 3.490 145.735 ;
        RECT 3.760 145.355 4.120 145.735 ;
        RECT 2.520 144.670 2.880 145.050 ;
        RECT 3.130 144.670 3.490 145.050 ;
        RECT 3.760 144.670 4.120 145.050 ;
        RECT 26.830 158.100 27.430 158.600 ;
        RECT 27.630 158.100 28.230 158.600 ;
        RECT 28.430 158.100 29.030 158.600 ;
        RECT 29.230 158.100 29.830 158.600 ;
        RECT 30.030 158.100 30.630 158.600 ;
        RECT 38.830 158.100 39.430 158.600 ;
        RECT 39.630 158.100 40.230 158.600 ;
        RECT 40.430 158.100 41.030 158.600 ;
        RECT 41.230 158.100 41.830 158.600 ;
        RECT 42.030 158.100 42.580 158.600 ;
        RECT 6.830 141.400 7.430 141.900 ;
        RECT 7.630 141.400 8.230 141.900 ;
        RECT 8.430 141.400 9.030 141.900 ;
        RECT 9.230 141.400 9.830 141.900 ;
        RECT 10.030 141.400 10.630 141.900 ;
        RECT 18.830 141.400 19.430 141.900 ;
        RECT 19.630 141.400 20.230 141.900 ;
        RECT 20.430 141.400 21.030 141.900 ;
        RECT 21.230 141.400 21.830 141.900 ;
        RECT 22.030 141.400 22.580 141.900 ;
        RECT 46.830 158.100 47.430 158.600 ;
        RECT 47.630 158.100 48.230 158.600 ;
        RECT 48.430 158.100 49.030 158.600 ;
        RECT 49.230 158.100 49.830 158.600 ;
        RECT 50.030 158.100 50.630 158.600 ;
        RECT 58.830 158.100 59.430 158.600 ;
        RECT 59.630 158.100 60.230 158.600 ;
        RECT 60.430 158.100 61.030 158.600 ;
        RECT 61.230 158.100 61.830 158.600 ;
        RECT 62.030 158.100 62.580 158.600 ;
        RECT 26.830 141.400 27.430 141.900 ;
        RECT 27.630 141.400 28.230 141.900 ;
        RECT 28.430 141.400 29.030 141.900 ;
        RECT 29.230 141.400 29.830 141.900 ;
        RECT 30.030 141.400 30.630 141.900 ;
        RECT 38.830 141.400 39.430 141.900 ;
        RECT 39.630 141.400 40.230 141.900 ;
        RECT 40.430 141.400 41.030 141.900 ;
        RECT 41.230 141.400 41.830 141.900 ;
        RECT 42.030 141.400 42.580 141.900 ;
        RECT 66.830 158.100 67.430 158.600 ;
        RECT 67.630 158.100 68.230 158.600 ;
        RECT 68.430 158.100 69.030 158.600 ;
        RECT 69.230 158.100 69.830 158.600 ;
        RECT 70.030 158.100 70.630 158.600 ;
        RECT 78.830 158.100 79.430 158.600 ;
        RECT 79.630 158.100 80.230 158.600 ;
        RECT 80.430 158.100 81.030 158.600 ;
        RECT 81.230 158.100 81.830 158.600 ;
        RECT 82.030 158.100 82.580 158.600 ;
        RECT 46.830 141.400 47.430 141.900 ;
        RECT 47.630 141.400 48.230 141.900 ;
        RECT 48.430 141.400 49.030 141.900 ;
        RECT 49.230 141.400 49.830 141.900 ;
        RECT 50.030 141.400 50.630 141.900 ;
        RECT 58.830 141.400 59.430 141.900 ;
        RECT 59.630 141.400 60.230 141.900 ;
        RECT 60.430 141.400 61.030 141.900 ;
        RECT 61.230 141.400 61.830 141.900 ;
        RECT 62.030 141.400 62.580 141.900 ;
        RECT 86.830 158.100 87.430 158.600 ;
        RECT 87.630 158.100 88.230 158.600 ;
        RECT 88.430 158.100 89.030 158.600 ;
        RECT 89.230 158.100 89.830 158.600 ;
        RECT 90.030 158.100 90.630 158.600 ;
        RECT 98.830 158.100 99.430 158.600 ;
        RECT 99.630 158.100 100.230 158.600 ;
        RECT 100.430 158.100 101.030 158.600 ;
        RECT 101.230 158.100 101.830 158.600 ;
        RECT 102.030 158.100 102.580 158.600 ;
        RECT 66.830 141.400 67.430 141.900 ;
        RECT 67.630 141.400 68.230 141.900 ;
        RECT 68.430 141.400 69.030 141.900 ;
        RECT 69.230 141.400 69.830 141.900 ;
        RECT 70.030 141.400 70.630 141.900 ;
        RECT 78.830 141.400 79.430 141.900 ;
        RECT 79.630 141.400 80.230 141.900 ;
        RECT 80.430 141.400 81.030 141.900 ;
        RECT 81.230 141.400 81.830 141.900 ;
        RECT 82.030 141.400 82.580 141.900 ;
        RECT 86.830 141.400 87.430 141.900 ;
        RECT 87.630 141.400 88.230 141.900 ;
        RECT 88.430 141.400 89.030 141.900 ;
        RECT 89.230 141.400 89.830 141.900 ;
        RECT 90.030 141.400 90.630 141.900 ;
        RECT 98.830 141.400 99.430 141.900 ;
        RECT 99.630 141.400 100.230 141.900 ;
        RECT 100.430 141.400 101.030 141.900 ;
        RECT 101.230 141.400 101.830 141.900 ;
        RECT 102.030 141.400 102.580 141.900 ;
        RECT 6.830 138.100 7.430 138.600 ;
        RECT 7.630 138.100 8.230 138.600 ;
        RECT 8.430 138.100 9.030 138.600 ;
        RECT 9.230 138.100 9.830 138.600 ;
        RECT 10.030 138.100 10.630 138.600 ;
        RECT 18.830 138.100 19.430 138.600 ;
        RECT 19.630 138.100 20.230 138.600 ;
        RECT 20.430 138.100 21.030 138.600 ;
        RECT 21.230 138.100 21.830 138.600 ;
        RECT 22.030 138.100 22.580 138.600 ;
        RECT 2.520 134.920 2.880 135.300 ;
        RECT 3.130 134.920 3.490 135.300 ;
        RECT 3.760 134.920 4.120 135.300 ;
        RECT 2.520 134.185 2.880 134.565 ;
        RECT 3.130 134.185 3.490 134.565 ;
        RECT 3.760 134.185 4.120 134.565 ;
        RECT 2.520 133.500 2.880 133.880 ;
        RECT 3.130 133.500 3.490 133.880 ;
        RECT 3.760 133.500 4.120 133.880 ;
        RECT 2.520 126.120 2.880 126.500 ;
        RECT 3.130 126.120 3.490 126.500 ;
        RECT 3.760 126.120 4.120 126.500 ;
        RECT 2.520 125.385 2.880 125.765 ;
        RECT 3.130 125.385 3.490 125.765 ;
        RECT 3.760 125.385 4.120 125.765 ;
        RECT 2.520 124.700 2.880 125.080 ;
        RECT 3.130 124.700 3.490 125.080 ;
        RECT 3.760 124.700 4.120 125.080 ;
        RECT 26.830 138.100 27.430 138.600 ;
        RECT 27.630 138.100 28.230 138.600 ;
        RECT 28.430 138.100 29.030 138.600 ;
        RECT 29.230 138.100 29.830 138.600 ;
        RECT 30.030 138.100 30.630 138.600 ;
        RECT 38.830 138.100 39.430 138.600 ;
        RECT 39.630 138.100 40.230 138.600 ;
        RECT 40.430 138.100 41.030 138.600 ;
        RECT 41.230 138.100 41.830 138.600 ;
        RECT 42.030 138.100 42.580 138.600 ;
        RECT 6.830 121.400 7.430 121.900 ;
        RECT 7.630 121.400 8.230 121.900 ;
        RECT 8.430 121.400 9.030 121.900 ;
        RECT 9.230 121.400 9.830 121.900 ;
        RECT 10.030 121.400 10.630 121.900 ;
        RECT 18.830 121.400 19.430 121.900 ;
        RECT 19.630 121.400 20.230 121.900 ;
        RECT 20.430 121.400 21.030 121.900 ;
        RECT 21.230 121.400 21.830 121.900 ;
        RECT 22.030 121.400 22.580 121.900 ;
        RECT 46.830 138.100 47.430 138.600 ;
        RECT 47.630 138.100 48.230 138.600 ;
        RECT 48.430 138.100 49.030 138.600 ;
        RECT 49.230 138.100 49.830 138.600 ;
        RECT 50.030 138.100 50.630 138.600 ;
        RECT 58.830 138.100 59.430 138.600 ;
        RECT 59.630 138.100 60.230 138.600 ;
        RECT 60.430 138.100 61.030 138.600 ;
        RECT 61.230 138.100 61.830 138.600 ;
        RECT 62.030 138.100 62.580 138.600 ;
        RECT 26.830 121.400 27.430 121.900 ;
        RECT 27.630 121.400 28.230 121.900 ;
        RECT 28.430 121.400 29.030 121.900 ;
        RECT 29.230 121.400 29.830 121.900 ;
        RECT 30.030 121.400 30.630 121.900 ;
        RECT 38.830 121.400 39.430 121.900 ;
        RECT 39.630 121.400 40.230 121.900 ;
        RECT 40.430 121.400 41.030 121.900 ;
        RECT 41.230 121.400 41.830 121.900 ;
        RECT 42.030 121.400 42.580 121.900 ;
        RECT 66.830 138.100 67.430 138.600 ;
        RECT 67.630 138.100 68.230 138.600 ;
        RECT 68.430 138.100 69.030 138.600 ;
        RECT 69.230 138.100 69.830 138.600 ;
        RECT 70.030 138.100 70.630 138.600 ;
        RECT 78.830 138.100 79.430 138.600 ;
        RECT 79.630 138.100 80.230 138.600 ;
        RECT 80.430 138.100 81.030 138.600 ;
        RECT 81.230 138.100 81.830 138.600 ;
        RECT 82.030 138.100 82.580 138.600 ;
        RECT 46.830 121.400 47.430 121.900 ;
        RECT 47.630 121.400 48.230 121.900 ;
        RECT 48.430 121.400 49.030 121.900 ;
        RECT 49.230 121.400 49.830 121.900 ;
        RECT 50.030 121.400 50.630 121.900 ;
        RECT 58.830 121.400 59.430 121.900 ;
        RECT 59.630 121.400 60.230 121.900 ;
        RECT 60.430 121.400 61.030 121.900 ;
        RECT 61.230 121.400 61.830 121.900 ;
        RECT 62.030 121.400 62.580 121.900 ;
        RECT 86.830 138.100 87.430 138.600 ;
        RECT 87.630 138.100 88.230 138.600 ;
        RECT 88.430 138.100 89.030 138.600 ;
        RECT 89.230 138.100 89.830 138.600 ;
        RECT 90.030 138.100 90.630 138.600 ;
        RECT 98.830 138.100 99.430 138.600 ;
        RECT 99.630 138.100 100.230 138.600 ;
        RECT 100.430 138.100 101.030 138.600 ;
        RECT 101.230 138.100 101.830 138.600 ;
        RECT 102.030 138.100 102.580 138.600 ;
        RECT 66.830 121.400 67.430 121.900 ;
        RECT 67.630 121.400 68.230 121.900 ;
        RECT 68.430 121.400 69.030 121.900 ;
        RECT 69.230 121.400 69.830 121.900 ;
        RECT 70.030 121.400 70.630 121.900 ;
        RECT 78.830 121.400 79.430 121.900 ;
        RECT 79.630 121.400 80.230 121.900 ;
        RECT 80.430 121.400 81.030 121.900 ;
        RECT 81.230 121.400 81.830 121.900 ;
        RECT 82.030 121.400 82.580 121.900 ;
        RECT 86.830 121.400 87.430 121.900 ;
        RECT 87.630 121.400 88.230 121.900 ;
        RECT 88.430 121.400 89.030 121.900 ;
        RECT 89.230 121.400 89.830 121.900 ;
        RECT 90.030 121.400 90.630 121.900 ;
        RECT 98.830 121.400 99.430 121.900 ;
        RECT 99.630 121.400 100.230 121.900 ;
        RECT 100.430 121.400 101.030 121.900 ;
        RECT 101.230 121.400 101.830 121.900 ;
        RECT 102.030 121.400 102.580 121.900 ;
        RECT 6.830 118.100 7.430 118.600 ;
        RECT 7.630 118.100 8.230 118.600 ;
        RECT 8.430 118.100 9.030 118.600 ;
        RECT 9.230 118.100 9.830 118.600 ;
        RECT 10.030 118.100 10.630 118.600 ;
        RECT 18.830 118.100 19.430 118.600 ;
        RECT 19.630 118.100 20.230 118.600 ;
        RECT 20.430 118.100 21.030 118.600 ;
        RECT 21.230 118.100 21.830 118.600 ;
        RECT 22.030 118.100 22.580 118.600 ;
        RECT 2.520 114.920 2.880 115.300 ;
        RECT 3.130 114.920 3.490 115.300 ;
        RECT 3.760 114.920 4.120 115.300 ;
        RECT 2.520 114.185 2.880 114.565 ;
        RECT 3.130 114.185 3.490 114.565 ;
        RECT 3.760 114.185 4.120 114.565 ;
        RECT 2.520 113.500 2.880 113.880 ;
        RECT 3.130 113.500 3.490 113.880 ;
        RECT 3.760 113.500 4.120 113.880 ;
        RECT 2.520 106.125 2.880 106.505 ;
        RECT 3.130 106.125 3.490 106.505 ;
        RECT 3.760 106.125 4.120 106.505 ;
        RECT 2.520 105.390 2.880 105.770 ;
        RECT 3.130 105.390 3.490 105.770 ;
        RECT 3.760 105.390 4.120 105.770 ;
        RECT 2.520 104.705 2.880 105.085 ;
        RECT 3.130 104.705 3.490 105.085 ;
        RECT 3.760 104.705 4.120 105.085 ;
        RECT 26.830 118.100 27.430 118.600 ;
        RECT 27.630 118.100 28.230 118.600 ;
        RECT 28.430 118.100 29.030 118.600 ;
        RECT 29.230 118.100 29.830 118.600 ;
        RECT 30.030 118.100 30.630 118.600 ;
        RECT 38.830 118.100 39.430 118.600 ;
        RECT 39.630 118.100 40.230 118.600 ;
        RECT 40.430 118.100 41.030 118.600 ;
        RECT 41.230 118.100 41.830 118.600 ;
        RECT 42.030 118.100 42.580 118.600 ;
        RECT 6.830 101.400 7.430 101.900 ;
        RECT 7.630 101.400 8.230 101.900 ;
        RECT 8.430 101.400 9.030 101.900 ;
        RECT 9.230 101.400 9.830 101.900 ;
        RECT 10.030 101.400 10.630 101.900 ;
        RECT 18.830 101.400 19.430 101.900 ;
        RECT 19.630 101.400 20.230 101.900 ;
        RECT 20.430 101.400 21.030 101.900 ;
        RECT 21.230 101.400 21.830 101.900 ;
        RECT 22.030 101.400 22.580 101.900 ;
        RECT 46.830 118.100 47.430 118.600 ;
        RECT 47.630 118.100 48.230 118.600 ;
        RECT 48.430 118.100 49.030 118.600 ;
        RECT 49.230 118.100 49.830 118.600 ;
        RECT 50.030 118.100 50.630 118.600 ;
        RECT 58.830 118.100 59.430 118.600 ;
        RECT 59.630 118.100 60.230 118.600 ;
        RECT 60.430 118.100 61.030 118.600 ;
        RECT 61.230 118.100 61.830 118.600 ;
        RECT 62.030 118.100 62.580 118.600 ;
        RECT 26.830 101.400 27.430 101.900 ;
        RECT 27.630 101.400 28.230 101.900 ;
        RECT 28.430 101.400 29.030 101.900 ;
        RECT 29.230 101.400 29.830 101.900 ;
        RECT 30.030 101.400 30.630 101.900 ;
        RECT 38.830 101.400 39.430 101.900 ;
        RECT 39.630 101.400 40.230 101.900 ;
        RECT 40.430 101.400 41.030 101.900 ;
        RECT 41.230 101.400 41.830 101.900 ;
        RECT 42.030 101.400 42.580 101.900 ;
        RECT 66.830 118.100 67.430 118.600 ;
        RECT 67.630 118.100 68.230 118.600 ;
        RECT 68.430 118.100 69.030 118.600 ;
        RECT 69.230 118.100 69.830 118.600 ;
        RECT 70.030 118.100 70.630 118.600 ;
        RECT 78.830 118.100 79.430 118.600 ;
        RECT 79.630 118.100 80.230 118.600 ;
        RECT 80.430 118.100 81.030 118.600 ;
        RECT 81.230 118.100 81.830 118.600 ;
        RECT 82.030 118.100 82.580 118.600 ;
        RECT 46.830 101.400 47.430 101.900 ;
        RECT 47.630 101.400 48.230 101.900 ;
        RECT 48.430 101.400 49.030 101.900 ;
        RECT 49.230 101.400 49.830 101.900 ;
        RECT 50.030 101.400 50.630 101.900 ;
        RECT 58.830 101.400 59.430 101.900 ;
        RECT 59.630 101.400 60.230 101.900 ;
        RECT 60.430 101.400 61.030 101.900 ;
        RECT 61.230 101.400 61.830 101.900 ;
        RECT 62.030 101.400 62.580 101.900 ;
        RECT 86.830 118.100 87.430 118.600 ;
        RECT 87.630 118.100 88.230 118.600 ;
        RECT 88.430 118.100 89.030 118.600 ;
        RECT 89.230 118.100 89.830 118.600 ;
        RECT 90.030 118.100 90.630 118.600 ;
        RECT 98.830 118.100 99.430 118.600 ;
        RECT 99.630 118.100 100.230 118.600 ;
        RECT 100.430 118.100 101.030 118.600 ;
        RECT 101.230 118.100 101.830 118.600 ;
        RECT 102.030 118.100 102.580 118.600 ;
        RECT 66.830 101.400 67.430 101.900 ;
        RECT 67.630 101.400 68.230 101.900 ;
        RECT 68.430 101.400 69.030 101.900 ;
        RECT 69.230 101.400 69.830 101.900 ;
        RECT 70.030 101.400 70.630 101.900 ;
        RECT 78.830 101.400 79.430 101.900 ;
        RECT 79.630 101.400 80.230 101.900 ;
        RECT 80.430 101.400 81.030 101.900 ;
        RECT 81.230 101.400 81.830 101.900 ;
        RECT 82.030 101.400 82.580 101.900 ;
        RECT 86.830 101.400 87.430 101.900 ;
        RECT 87.630 101.400 88.230 101.900 ;
        RECT 88.430 101.400 89.030 101.900 ;
        RECT 89.230 101.400 89.830 101.900 ;
        RECT 90.030 101.400 90.630 101.900 ;
        RECT 98.830 101.400 99.430 101.900 ;
        RECT 99.630 101.400 100.230 101.900 ;
        RECT 100.430 101.400 101.030 101.900 ;
        RECT 101.230 101.400 101.830 101.900 ;
        RECT 102.030 101.400 102.580 101.900 ;
        RECT 6.830 98.100 7.430 98.600 ;
        RECT 7.630 98.100 8.230 98.600 ;
        RECT 8.430 98.100 9.030 98.600 ;
        RECT 9.230 98.100 9.830 98.600 ;
        RECT 10.030 98.100 10.630 98.600 ;
        RECT 18.830 98.100 19.430 98.600 ;
        RECT 19.630 98.100 20.230 98.600 ;
        RECT 20.430 98.100 21.030 98.600 ;
        RECT 21.230 98.100 21.830 98.600 ;
        RECT 22.030 98.100 22.580 98.600 ;
        RECT 2.520 94.920 2.880 95.300 ;
        RECT 3.130 94.920 3.490 95.300 ;
        RECT 3.760 94.920 4.120 95.300 ;
        RECT 2.520 94.185 2.880 94.565 ;
        RECT 3.130 94.185 3.490 94.565 ;
        RECT 3.760 94.185 4.120 94.565 ;
        RECT 2.520 93.500 2.880 93.880 ;
        RECT 3.130 93.500 3.490 93.880 ;
        RECT 3.760 93.500 4.120 93.880 ;
        RECT 2.520 86.120 2.880 86.500 ;
        RECT 3.130 86.120 3.490 86.500 ;
        RECT 3.760 86.120 4.120 86.500 ;
        RECT 2.520 85.385 2.880 85.765 ;
        RECT 3.130 85.385 3.490 85.765 ;
        RECT 3.760 85.385 4.120 85.765 ;
        RECT 2.520 84.700 2.880 85.080 ;
        RECT 3.130 84.700 3.490 85.080 ;
        RECT 3.760 84.700 4.120 85.080 ;
        RECT 26.830 98.100 27.430 98.600 ;
        RECT 27.630 98.100 28.230 98.600 ;
        RECT 28.430 98.100 29.030 98.600 ;
        RECT 29.230 98.100 29.830 98.600 ;
        RECT 30.030 98.100 30.630 98.600 ;
        RECT 38.830 98.100 39.430 98.600 ;
        RECT 39.630 98.100 40.230 98.600 ;
        RECT 40.430 98.100 41.030 98.600 ;
        RECT 41.230 98.100 41.830 98.600 ;
        RECT 42.030 98.100 42.580 98.600 ;
        RECT 6.830 81.400 7.430 81.900 ;
        RECT 7.630 81.400 8.230 81.900 ;
        RECT 8.430 81.400 9.030 81.900 ;
        RECT 9.230 81.400 9.830 81.900 ;
        RECT 10.030 81.400 10.630 81.900 ;
        RECT 18.830 81.400 19.430 81.900 ;
        RECT 19.630 81.400 20.230 81.900 ;
        RECT 20.430 81.400 21.030 81.900 ;
        RECT 21.230 81.400 21.830 81.900 ;
        RECT 22.030 81.400 22.580 81.900 ;
        RECT 46.830 98.100 47.430 98.600 ;
        RECT 47.630 98.100 48.230 98.600 ;
        RECT 48.430 98.100 49.030 98.600 ;
        RECT 49.230 98.100 49.830 98.600 ;
        RECT 50.030 98.100 50.630 98.600 ;
        RECT 58.830 98.100 59.430 98.600 ;
        RECT 59.630 98.100 60.230 98.600 ;
        RECT 60.430 98.100 61.030 98.600 ;
        RECT 61.230 98.100 61.830 98.600 ;
        RECT 62.030 98.100 62.580 98.600 ;
        RECT 26.830 81.400 27.430 81.900 ;
        RECT 27.630 81.400 28.230 81.900 ;
        RECT 28.430 81.400 29.030 81.900 ;
        RECT 29.230 81.400 29.830 81.900 ;
        RECT 30.030 81.400 30.630 81.900 ;
        RECT 38.830 81.400 39.430 81.900 ;
        RECT 39.630 81.400 40.230 81.900 ;
        RECT 40.430 81.400 41.030 81.900 ;
        RECT 41.230 81.400 41.830 81.900 ;
        RECT 42.030 81.400 42.580 81.900 ;
        RECT 66.830 98.100 67.430 98.600 ;
        RECT 67.630 98.100 68.230 98.600 ;
        RECT 68.430 98.100 69.030 98.600 ;
        RECT 69.230 98.100 69.830 98.600 ;
        RECT 70.030 98.100 70.630 98.600 ;
        RECT 78.830 98.100 79.430 98.600 ;
        RECT 79.630 98.100 80.230 98.600 ;
        RECT 80.430 98.100 81.030 98.600 ;
        RECT 81.230 98.100 81.830 98.600 ;
        RECT 82.030 98.100 82.580 98.600 ;
        RECT 46.830 81.400 47.430 81.900 ;
        RECT 47.630 81.400 48.230 81.900 ;
        RECT 48.430 81.400 49.030 81.900 ;
        RECT 49.230 81.400 49.830 81.900 ;
        RECT 50.030 81.400 50.630 81.900 ;
        RECT 58.830 81.400 59.430 81.900 ;
        RECT 59.630 81.400 60.230 81.900 ;
        RECT 60.430 81.400 61.030 81.900 ;
        RECT 61.230 81.400 61.830 81.900 ;
        RECT 62.030 81.400 62.580 81.900 ;
        RECT 86.830 98.100 87.430 98.600 ;
        RECT 87.630 98.100 88.230 98.600 ;
        RECT 88.430 98.100 89.030 98.600 ;
        RECT 89.230 98.100 89.830 98.600 ;
        RECT 90.030 98.100 90.630 98.600 ;
        RECT 98.830 98.100 99.430 98.600 ;
        RECT 99.630 98.100 100.230 98.600 ;
        RECT 100.430 98.100 101.030 98.600 ;
        RECT 101.230 98.100 101.830 98.600 ;
        RECT 102.030 98.100 102.580 98.600 ;
        RECT 66.830 81.400 67.430 81.900 ;
        RECT 67.630 81.400 68.230 81.900 ;
        RECT 68.430 81.400 69.030 81.900 ;
        RECT 69.230 81.400 69.830 81.900 ;
        RECT 70.030 81.400 70.630 81.900 ;
        RECT 78.830 81.400 79.430 81.900 ;
        RECT 79.630 81.400 80.230 81.900 ;
        RECT 80.430 81.400 81.030 81.900 ;
        RECT 81.230 81.400 81.830 81.900 ;
        RECT 82.030 81.400 82.580 81.900 ;
        RECT 86.830 81.400 87.430 81.900 ;
        RECT 87.630 81.400 88.230 81.900 ;
        RECT 88.430 81.400 89.030 81.900 ;
        RECT 89.230 81.400 89.830 81.900 ;
        RECT 90.030 81.400 90.630 81.900 ;
        RECT 98.830 81.400 99.430 81.900 ;
        RECT 99.630 81.400 100.230 81.900 ;
        RECT 100.430 81.400 101.030 81.900 ;
        RECT 101.230 81.400 101.830 81.900 ;
        RECT 102.030 81.400 102.580 81.900 ;
        RECT 6.830 78.100 7.430 78.600 ;
        RECT 7.630 78.100 8.230 78.600 ;
        RECT 8.430 78.100 9.030 78.600 ;
        RECT 9.230 78.100 9.830 78.600 ;
        RECT 10.030 78.100 10.630 78.600 ;
        RECT 18.830 78.100 19.430 78.600 ;
        RECT 19.630 78.100 20.230 78.600 ;
        RECT 20.430 78.100 21.030 78.600 ;
        RECT 21.230 78.100 21.830 78.600 ;
        RECT 22.030 78.100 22.580 78.600 ;
        RECT 2.520 74.920 2.880 75.300 ;
        RECT 3.130 74.920 3.490 75.300 ;
        RECT 3.760 74.920 4.120 75.300 ;
        RECT 2.520 74.185 2.880 74.565 ;
        RECT 3.130 74.185 3.490 74.565 ;
        RECT 3.760 74.185 4.120 74.565 ;
        RECT 2.520 73.500 2.880 73.880 ;
        RECT 3.130 73.500 3.490 73.880 ;
        RECT 3.760 73.500 4.120 73.880 ;
        RECT 2.520 66.120 2.880 66.500 ;
        RECT 3.130 66.120 3.490 66.500 ;
        RECT 3.760 66.120 4.120 66.500 ;
        RECT 2.520 65.385 2.880 65.765 ;
        RECT 3.130 65.385 3.490 65.765 ;
        RECT 3.760 65.385 4.120 65.765 ;
        RECT 2.520 64.700 2.880 65.080 ;
        RECT 3.130 64.700 3.490 65.080 ;
        RECT 3.760 64.700 4.120 65.080 ;
        RECT 26.830 78.100 27.430 78.600 ;
        RECT 27.630 78.100 28.230 78.600 ;
        RECT 28.430 78.100 29.030 78.600 ;
        RECT 29.230 78.100 29.830 78.600 ;
        RECT 30.030 78.100 30.630 78.600 ;
        RECT 38.830 78.100 39.430 78.600 ;
        RECT 39.630 78.100 40.230 78.600 ;
        RECT 40.430 78.100 41.030 78.600 ;
        RECT 41.230 78.100 41.830 78.600 ;
        RECT 42.030 78.100 42.580 78.600 ;
        RECT 6.830 61.400 7.430 61.900 ;
        RECT 7.630 61.400 8.230 61.900 ;
        RECT 8.430 61.400 9.030 61.900 ;
        RECT 9.230 61.400 9.830 61.900 ;
        RECT 10.030 61.400 10.630 61.900 ;
        RECT 18.830 61.400 19.430 61.900 ;
        RECT 19.630 61.400 20.230 61.900 ;
        RECT 20.430 61.400 21.030 61.900 ;
        RECT 21.230 61.400 21.830 61.900 ;
        RECT 22.030 61.400 22.580 61.900 ;
        RECT 46.830 78.100 47.430 78.600 ;
        RECT 47.630 78.100 48.230 78.600 ;
        RECT 48.430 78.100 49.030 78.600 ;
        RECT 49.230 78.100 49.830 78.600 ;
        RECT 50.030 78.100 50.630 78.600 ;
        RECT 58.830 78.100 59.430 78.600 ;
        RECT 59.630 78.100 60.230 78.600 ;
        RECT 60.430 78.100 61.030 78.600 ;
        RECT 61.230 78.100 61.830 78.600 ;
        RECT 62.030 78.100 62.580 78.600 ;
        RECT 26.830 61.400 27.430 61.900 ;
        RECT 27.630 61.400 28.230 61.900 ;
        RECT 28.430 61.400 29.030 61.900 ;
        RECT 29.230 61.400 29.830 61.900 ;
        RECT 30.030 61.400 30.630 61.900 ;
        RECT 38.830 61.400 39.430 61.900 ;
        RECT 39.630 61.400 40.230 61.900 ;
        RECT 40.430 61.400 41.030 61.900 ;
        RECT 41.230 61.400 41.830 61.900 ;
        RECT 42.030 61.400 42.580 61.900 ;
        RECT 66.830 78.100 67.430 78.600 ;
        RECT 67.630 78.100 68.230 78.600 ;
        RECT 68.430 78.100 69.030 78.600 ;
        RECT 69.230 78.100 69.830 78.600 ;
        RECT 70.030 78.100 70.630 78.600 ;
        RECT 78.830 78.100 79.430 78.600 ;
        RECT 79.630 78.100 80.230 78.600 ;
        RECT 80.430 78.100 81.030 78.600 ;
        RECT 81.230 78.100 81.830 78.600 ;
        RECT 82.030 78.100 82.580 78.600 ;
        RECT 46.830 61.400 47.430 61.900 ;
        RECT 47.630 61.400 48.230 61.900 ;
        RECT 48.430 61.400 49.030 61.900 ;
        RECT 49.230 61.400 49.830 61.900 ;
        RECT 50.030 61.400 50.630 61.900 ;
        RECT 58.830 61.400 59.430 61.900 ;
        RECT 59.630 61.400 60.230 61.900 ;
        RECT 60.430 61.400 61.030 61.900 ;
        RECT 61.230 61.400 61.830 61.900 ;
        RECT 62.030 61.400 62.580 61.900 ;
        RECT 86.830 78.100 87.430 78.600 ;
        RECT 87.630 78.100 88.230 78.600 ;
        RECT 88.430 78.100 89.030 78.600 ;
        RECT 89.230 78.100 89.830 78.600 ;
        RECT 90.030 78.100 90.630 78.600 ;
        RECT 98.830 78.100 99.430 78.600 ;
        RECT 99.630 78.100 100.230 78.600 ;
        RECT 100.430 78.100 101.030 78.600 ;
        RECT 101.230 78.100 101.830 78.600 ;
        RECT 102.030 78.100 102.580 78.600 ;
        RECT 66.830 61.400 67.430 61.900 ;
        RECT 67.630 61.400 68.230 61.900 ;
        RECT 68.430 61.400 69.030 61.900 ;
        RECT 69.230 61.400 69.830 61.900 ;
        RECT 70.030 61.400 70.630 61.900 ;
        RECT 78.830 61.400 79.430 61.900 ;
        RECT 79.630 61.400 80.230 61.900 ;
        RECT 80.430 61.400 81.030 61.900 ;
        RECT 81.230 61.400 81.830 61.900 ;
        RECT 82.030 61.400 82.580 61.900 ;
        RECT 86.830 61.400 87.430 61.900 ;
        RECT 87.630 61.400 88.230 61.900 ;
        RECT 88.430 61.400 89.030 61.900 ;
        RECT 89.230 61.400 89.830 61.900 ;
        RECT 90.030 61.400 90.630 61.900 ;
        RECT 98.830 61.400 99.430 61.900 ;
        RECT 99.630 61.400 100.230 61.900 ;
        RECT 100.430 61.400 101.030 61.900 ;
        RECT 101.230 61.400 101.830 61.900 ;
        RECT 102.030 61.400 102.580 61.900 ;
        RECT 6.830 58.100 7.430 58.600 ;
        RECT 7.630 58.100 8.230 58.600 ;
        RECT 8.430 58.100 9.030 58.600 ;
        RECT 9.230 58.100 9.830 58.600 ;
        RECT 10.030 58.100 10.630 58.600 ;
        RECT 18.830 58.100 19.430 58.600 ;
        RECT 19.630 58.100 20.230 58.600 ;
        RECT 20.430 58.100 21.030 58.600 ;
        RECT 21.230 58.100 21.830 58.600 ;
        RECT 22.030 58.100 22.580 58.600 ;
        RECT 2.520 54.925 2.880 55.305 ;
        RECT 3.130 54.925 3.490 55.305 ;
        RECT 3.760 54.925 4.120 55.305 ;
        RECT 2.520 54.190 2.880 54.570 ;
        RECT 3.130 54.190 3.490 54.570 ;
        RECT 3.760 54.190 4.120 54.570 ;
        RECT 2.520 53.505 2.880 53.885 ;
        RECT 3.130 53.505 3.490 53.885 ;
        RECT 3.760 53.505 4.120 53.885 ;
        RECT 2.520 46.115 2.880 46.495 ;
        RECT 3.130 46.115 3.490 46.495 ;
        RECT 3.760 46.115 4.120 46.495 ;
        RECT 2.520 45.380 2.880 45.760 ;
        RECT 3.130 45.380 3.490 45.760 ;
        RECT 3.760 45.380 4.120 45.760 ;
        RECT 2.520 44.695 2.880 45.075 ;
        RECT 3.130 44.695 3.490 45.075 ;
        RECT 3.760 44.695 4.120 45.075 ;
        RECT 26.830 58.100 27.430 58.600 ;
        RECT 27.630 58.100 28.230 58.600 ;
        RECT 28.430 58.100 29.030 58.600 ;
        RECT 29.230 58.100 29.830 58.600 ;
        RECT 30.030 58.100 30.630 58.600 ;
        RECT 38.830 58.100 39.430 58.600 ;
        RECT 39.630 58.100 40.230 58.600 ;
        RECT 40.430 58.100 41.030 58.600 ;
        RECT 41.230 58.100 41.830 58.600 ;
        RECT 42.030 58.100 42.580 58.600 ;
        RECT 6.830 41.400 7.430 41.900 ;
        RECT 7.630 41.400 8.230 41.900 ;
        RECT 8.430 41.400 9.030 41.900 ;
        RECT 9.230 41.400 9.830 41.900 ;
        RECT 10.030 41.400 10.630 41.900 ;
        RECT 18.830 41.400 19.430 41.900 ;
        RECT 19.630 41.400 20.230 41.900 ;
        RECT 20.430 41.400 21.030 41.900 ;
        RECT 21.230 41.400 21.830 41.900 ;
        RECT 22.030 41.400 22.580 41.900 ;
        RECT 46.830 58.100 47.430 58.600 ;
        RECT 47.630 58.100 48.230 58.600 ;
        RECT 48.430 58.100 49.030 58.600 ;
        RECT 49.230 58.100 49.830 58.600 ;
        RECT 50.030 58.100 50.630 58.600 ;
        RECT 58.830 58.100 59.430 58.600 ;
        RECT 59.630 58.100 60.230 58.600 ;
        RECT 60.430 58.100 61.030 58.600 ;
        RECT 61.230 58.100 61.830 58.600 ;
        RECT 62.030 58.100 62.580 58.600 ;
        RECT 26.830 41.400 27.430 41.900 ;
        RECT 27.630 41.400 28.230 41.900 ;
        RECT 28.430 41.400 29.030 41.900 ;
        RECT 29.230 41.400 29.830 41.900 ;
        RECT 30.030 41.400 30.630 41.900 ;
        RECT 38.830 41.400 39.430 41.900 ;
        RECT 39.630 41.400 40.230 41.900 ;
        RECT 40.430 41.400 41.030 41.900 ;
        RECT 41.230 41.400 41.830 41.900 ;
        RECT 42.030 41.400 42.580 41.900 ;
        RECT 66.830 58.100 67.430 58.600 ;
        RECT 67.630 58.100 68.230 58.600 ;
        RECT 68.430 58.100 69.030 58.600 ;
        RECT 69.230 58.100 69.830 58.600 ;
        RECT 70.030 58.100 70.630 58.600 ;
        RECT 78.830 58.100 79.430 58.600 ;
        RECT 79.630 58.100 80.230 58.600 ;
        RECT 80.430 58.100 81.030 58.600 ;
        RECT 81.230 58.100 81.830 58.600 ;
        RECT 82.030 58.100 82.580 58.600 ;
        RECT 46.830 41.400 47.430 41.900 ;
        RECT 47.630 41.400 48.230 41.900 ;
        RECT 48.430 41.400 49.030 41.900 ;
        RECT 49.230 41.400 49.830 41.900 ;
        RECT 50.030 41.400 50.630 41.900 ;
        RECT 58.830 41.400 59.430 41.900 ;
        RECT 59.630 41.400 60.230 41.900 ;
        RECT 60.430 41.400 61.030 41.900 ;
        RECT 61.230 41.400 61.830 41.900 ;
        RECT 62.030 41.400 62.580 41.900 ;
        RECT 86.830 58.100 87.430 58.600 ;
        RECT 87.630 58.100 88.230 58.600 ;
        RECT 88.430 58.100 89.030 58.600 ;
        RECT 89.230 58.100 89.830 58.600 ;
        RECT 90.030 58.100 90.630 58.600 ;
        RECT 98.830 58.100 99.430 58.600 ;
        RECT 99.630 58.100 100.230 58.600 ;
        RECT 100.430 58.100 101.030 58.600 ;
        RECT 101.230 58.100 101.830 58.600 ;
        RECT 102.030 58.100 102.580 58.600 ;
        RECT 66.830 41.400 67.430 41.900 ;
        RECT 67.630 41.400 68.230 41.900 ;
        RECT 68.430 41.400 69.030 41.900 ;
        RECT 69.230 41.400 69.830 41.900 ;
        RECT 70.030 41.400 70.630 41.900 ;
        RECT 78.830 41.400 79.430 41.900 ;
        RECT 79.630 41.400 80.230 41.900 ;
        RECT 80.430 41.400 81.030 41.900 ;
        RECT 81.230 41.400 81.830 41.900 ;
        RECT 82.030 41.400 82.580 41.900 ;
        RECT 86.830 41.400 87.430 41.900 ;
        RECT 87.630 41.400 88.230 41.900 ;
        RECT 88.430 41.400 89.030 41.900 ;
        RECT 89.230 41.400 89.830 41.900 ;
        RECT 90.030 41.400 90.630 41.900 ;
        RECT 98.830 41.400 99.430 41.900 ;
        RECT 99.630 41.400 100.230 41.900 ;
        RECT 100.430 41.400 101.030 41.900 ;
        RECT 101.230 41.400 101.830 41.900 ;
        RECT 102.030 41.400 102.580 41.900 ;
        RECT 6.830 38.100 7.430 38.600 ;
        RECT 7.630 38.100 8.230 38.600 ;
        RECT 8.430 38.100 9.030 38.600 ;
        RECT 9.230 38.100 9.830 38.600 ;
        RECT 10.030 38.100 10.630 38.600 ;
        RECT 18.830 38.100 19.430 38.600 ;
        RECT 19.630 38.100 20.230 38.600 ;
        RECT 20.430 38.100 21.030 38.600 ;
        RECT 21.230 38.100 21.830 38.600 ;
        RECT 22.030 38.100 22.580 38.600 ;
        RECT 2.520 34.925 2.880 35.305 ;
        RECT 3.130 34.925 3.490 35.305 ;
        RECT 3.760 34.925 4.120 35.305 ;
        RECT 2.520 34.190 2.880 34.570 ;
        RECT 3.130 34.190 3.490 34.570 ;
        RECT 3.760 34.190 4.120 34.570 ;
        RECT 2.520 33.505 2.880 33.885 ;
        RECT 3.130 33.505 3.490 33.885 ;
        RECT 3.760 33.505 4.120 33.885 ;
        RECT 2.520 26.120 2.880 26.500 ;
        RECT 3.130 26.120 3.490 26.500 ;
        RECT 3.760 26.120 4.120 26.500 ;
        RECT 2.520 25.385 2.880 25.765 ;
        RECT 3.130 25.385 3.490 25.765 ;
        RECT 3.760 25.385 4.120 25.765 ;
        RECT 2.520 24.700 2.880 25.080 ;
        RECT 3.130 24.700 3.490 25.080 ;
        RECT 3.760 24.700 4.120 25.080 ;
        RECT 26.830 38.100 27.430 38.600 ;
        RECT 27.630 38.100 28.230 38.600 ;
        RECT 28.430 38.100 29.030 38.600 ;
        RECT 29.230 38.100 29.830 38.600 ;
        RECT 30.030 38.100 30.630 38.600 ;
        RECT 38.830 38.100 39.430 38.600 ;
        RECT 39.630 38.100 40.230 38.600 ;
        RECT 40.430 38.100 41.030 38.600 ;
        RECT 41.230 38.100 41.830 38.600 ;
        RECT 42.030 38.100 42.580 38.600 ;
        RECT 6.830 21.400 7.430 21.900 ;
        RECT 7.630 21.400 8.230 21.900 ;
        RECT 8.430 21.400 9.030 21.900 ;
        RECT 9.230 21.400 9.830 21.900 ;
        RECT 10.030 21.400 10.630 21.900 ;
        RECT 18.830 21.400 19.430 21.900 ;
        RECT 19.630 21.400 20.230 21.900 ;
        RECT 20.430 21.400 21.030 21.900 ;
        RECT 21.230 21.400 21.830 21.900 ;
        RECT 22.030 21.400 22.580 21.900 ;
        RECT 46.830 38.100 47.430 38.600 ;
        RECT 47.630 38.100 48.230 38.600 ;
        RECT 48.430 38.100 49.030 38.600 ;
        RECT 49.230 38.100 49.830 38.600 ;
        RECT 50.030 38.100 50.630 38.600 ;
        RECT 58.830 38.100 59.430 38.600 ;
        RECT 59.630 38.100 60.230 38.600 ;
        RECT 60.430 38.100 61.030 38.600 ;
        RECT 61.230 38.100 61.830 38.600 ;
        RECT 62.030 38.100 62.580 38.600 ;
        RECT 26.830 21.400 27.430 21.900 ;
        RECT 27.630 21.400 28.230 21.900 ;
        RECT 28.430 21.400 29.030 21.900 ;
        RECT 29.230 21.400 29.830 21.900 ;
        RECT 30.030 21.400 30.630 21.900 ;
        RECT 38.830 21.400 39.430 21.900 ;
        RECT 39.630 21.400 40.230 21.900 ;
        RECT 40.430 21.400 41.030 21.900 ;
        RECT 41.230 21.400 41.830 21.900 ;
        RECT 42.030 21.400 42.580 21.900 ;
        RECT 66.830 38.100 67.430 38.600 ;
        RECT 67.630 38.100 68.230 38.600 ;
        RECT 68.430 38.100 69.030 38.600 ;
        RECT 69.230 38.100 69.830 38.600 ;
        RECT 70.030 38.100 70.630 38.600 ;
        RECT 78.830 38.100 79.430 38.600 ;
        RECT 79.630 38.100 80.230 38.600 ;
        RECT 80.430 38.100 81.030 38.600 ;
        RECT 81.230 38.100 81.830 38.600 ;
        RECT 82.030 38.100 82.580 38.600 ;
        RECT 46.830 21.400 47.430 21.900 ;
        RECT 47.630 21.400 48.230 21.900 ;
        RECT 48.430 21.400 49.030 21.900 ;
        RECT 49.230 21.400 49.830 21.900 ;
        RECT 50.030 21.400 50.630 21.900 ;
        RECT 58.830 21.400 59.430 21.900 ;
        RECT 59.630 21.400 60.230 21.900 ;
        RECT 60.430 21.400 61.030 21.900 ;
        RECT 61.230 21.400 61.830 21.900 ;
        RECT 62.030 21.400 62.580 21.900 ;
        RECT 86.830 38.100 87.430 38.600 ;
        RECT 87.630 38.100 88.230 38.600 ;
        RECT 88.430 38.100 89.030 38.600 ;
        RECT 89.230 38.100 89.830 38.600 ;
        RECT 90.030 38.100 90.630 38.600 ;
        RECT 98.830 38.100 99.430 38.600 ;
        RECT 99.630 38.100 100.230 38.600 ;
        RECT 100.430 38.100 101.030 38.600 ;
        RECT 101.230 38.100 101.830 38.600 ;
        RECT 102.030 38.100 102.580 38.600 ;
        RECT 66.830 21.400 67.430 21.900 ;
        RECT 67.630 21.400 68.230 21.900 ;
        RECT 68.430 21.400 69.030 21.900 ;
        RECT 69.230 21.400 69.830 21.900 ;
        RECT 70.030 21.400 70.630 21.900 ;
        RECT 78.830 21.400 79.430 21.900 ;
        RECT 79.630 21.400 80.230 21.900 ;
        RECT 80.430 21.400 81.030 21.900 ;
        RECT 81.230 21.400 81.830 21.900 ;
        RECT 82.030 21.400 82.580 21.900 ;
        RECT 86.830 21.400 87.430 21.900 ;
        RECT 87.630 21.400 88.230 21.900 ;
        RECT 88.430 21.400 89.030 21.900 ;
        RECT 89.230 21.400 89.830 21.900 ;
        RECT 90.030 21.400 90.630 21.900 ;
        RECT 98.830 21.400 99.430 21.900 ;
        RECT 99.630 21.400 100.230 21.900 ;
        RECT 100.430 21.400 101.030 21.900 ;
        RECT 101.230 21.400 101.830 21.900 ;
        RECT 102.030 21.400 102.580 21.900 ;
        RECT 6.830 18.100 7.430 18.600 ;
        RECT 7.630 18.100 8.230 18.600 ;
        RECT 8.430 18.100 9.030 18.600 ;
        RECT 9.230 18.100 9.830 18.600 ;
        RECT 10.030 18.100 10.630 18.600 ;
        RECT 18.830 18.100 19.430 18.600 ;
        RECT 19.630 18.100 20.230 18.600 ;
        RECT 20.430 18.100 21.030 18.600 ;
        RECT 21.230 18.100 21.830 18.600 ;
        RECT 22.030 18.100 22.580 18.600 ;
        RECT 2.520 14.925 2.880 15.305 ;
        RECT 3.130 14.925 3.490 15.305 ;
        RECT 3.760 14.925 4.120 15.305 ;
        RECT 2.520 14.190 2.880 14.570 ;
        RECT 3.130 14.190 3.490 14.570 ;
        RECT 3.760 14.190 4.120 14.570 ;
        RECT 2.520 13.505 2.880 13.885 ;
        RECT 3.130 13.505 3.490 13.885 ;
        RECT 3.760 13.505 4.120 13.885 ;
        RECT 2.520 6.120 2.880 6.500 ;
        RECT 3.130 6.120 3.490 6.500 ;
        RECT 3.760 6.120 4.120 6.500 ;
        RECT 2.520 5.385 2.880 5.765 ;
        RECT 3.130 5.385 3.490 5.765 ;
        RECT 3.760 5.385 4.120 5.765 ;
        RECT 2.520 4.700 2.880 5.080 ;
        RECT 3.130 4.700 3.490 5.080 ;
        RECT 3.760 4.700 4.120 5.080 ;
        RECT 26.830 18.100 27.430 18.600 ;
        RECT 27.630 18.100 28.230 18.600 ;
        RECT 28.430 18.100 29.030 18.600 ;
        RECT 29.230 18.100 29.830 18.600 ;
        RECT 30.030 18.100 30.630 18.600 ;
        RECT 38.830 18.100 39.430 18.600 ;
        RECT 39.630 18.100 40.230 18.600 ;
        RECT 40.430 18.100 41.030 18.600 ;
        RECT 41.230 18.100 41.830 18.600 ;
        RECT 42.030 18.100 42.580 18.600 ;
        RECT 6.830 1.400 7.430 1.900 ;
        RECT 7.630 1.400 8.230 1.900 ;
        RECT 8.430 1.400 9.030 1.900 ;
        RECT 9.230 1.400 9.830 1.900 ;
        RECT 10.030 1.400 10.630 1.900 ;
        RECT 18.830 1.400 19.430 1.900 ;
        RECT 19.630 1.400 20.230 1.900 ;
        RECT 20.430 1.400 21.030 1.900 ;
        RECT 21.230 1.400 21.830 1.900 ;
        RECT 22.030 1.400 22.580 1.900 ;
        RECT 46.830 18.100 47.430 18.600 ;
        RECT 47.630 18.100 48.230 18.600 ;
        RECT 48.430 18.100 49.030 18.600 ;
        RECT 49.230 18.100 49.830 18.600 ;
        RECT 50.030 18.100 50.630 18.600 ;
        RECT 58.830 18.100 59.430 18.600 ;
        RECT 59.630 18.100 60.230 18.600 ;
        RECT 60.430 18.100 61.030 18.600 ;
        RECT 61.230 18.100 61.830 18.600 ;
        RECT 62.030 18.100 62.580 18.600 ;
        RECT 26.830 1.400 27.430 1.900 ;
        RECT 27.630 1.400 28.230 1.900 ;
        RECT 28.430 1.400 29.030 1.900 ;
        RECT 29.230 1.400 29.830 1.900 ;
        RECT 30.030 1.400 30.630 1.900 ;
        RECT 38.830 1.400 39.430 1.900 ;
        RECT 39.630 1.400 40.230 1.900 ;
        RECT 40.430 1.400 41.030 1.900 ;
        RECT 41.230 1.400 41.830 1.900 ;
        RECT 42.030 1.400 42.580 1.900 ;
        RECT 66.830 18.100 67.430 18.600 ;
        RECT 67.630 18.100 68.230 18.600 ;
        RECT 68.430 18.100 69.030 18.600 ;
        RECT 69.230 18.100 69.830 18.600 ;
        RECT 70.030 18.100 70.630 18.600 ;
        RECT 78.830 18.100 79.430 18.600 ;
        RECT 79.630 18.100 80.230 18.600 ;
        RECT 80.430 18.100 81.030 18.600 ;
        RECT 81.230 18.100 81.830 18.600 ;
        RECT 82.030 18.100 82.580 18.600 ;
        RECT 46.830 1.400 47.430 1.900 ;
        RECT 47.630 1.400 48.230 1.900 ;
        RECT 48.430 1.400 49.030 1.900 ;
        RECT 49.230 1.400 49.830 1.900 ;
        RECT 50.030 1.400 50.630 1.900 ;
        RECT 58.830 1.400 59.430 1.900 ;
        RECT 59.630 1.400 60.230 1.900 ;
        RECT 60.430 1.400 61.030 1.900 ;
        RECT 61.230 1.400 61.830 1.900 ;
        RECT 62.030 1.400 62.580 1.900 ;
        RECT 86.830 18.100 87.430 18.600 ;
        RECT 87.630 18.100 88.230 18.600 ;
        RECT 88.430 18.100 89.030 18.600 ;
        RECT 89.230 18.100 89.830 18.600 ;
        RECT 90.030 18.100 90.630 18.600 ;
        RECT 98.830 18.100 99.430 18.600 ;
        RECT 99.630 18.100 100.230 18.600 ;
        RECT 100.430 18.100 101.030 18.600 ;
        RECT 101.230 18.100 101.830 18.600 ;
        RECT 102.030 18.100 102.580 18.600 ;
        RECT 66.830 1.400 67.430 1.900 ;
        RECT 67.630 1.400 68.230 1.900 ;
        RECT 68.430 1.400 69.030 1.900 ;
        RECT 69.230 1.400 69.830 1.900 ;
        RECT 70.030 1.400 70.630 1.900 ;
        RECT 78.830 1.400 79.430 1.900 ;
        RECT 79.630 1.400 80.230 1.900 ;
        RECT 80.430 1.400 81.030 1.900 ;
        RECT 81.230 1.400 81.830 1.900 ;
        RECT 82.030 1.400 82.580 1.900 ;
        RECT 86.830 1.400 87.430 1.900 ;
        RECT 87.630 1.400 88.230 1.900 ;
        RECT 88.430 1.400 89.030 1.900 ;
        RECT 89.230 1.400 89.830 1.900 ;
        RECT 90.030 1.400 90.630 1.900 ;
        RECT 98.830 1.400 99.430 1.900 ;
        RECT 99.630 1.400 100.230 1.900 ;
        RECT 100.430 1.400 101.030 1.900 ;
        RECT 101.230 1.400 101.830 1.900 ;
        RECT 102.030 1.400 102.580 1.900 ;
      LAYER met1 ;
        RECT 4.730 379.850 9.130 380.000 ;
        RECT 20.330 379.850 29.130 380.000 ;
        RECT 40.330 379.850 49.130 380.000 ;
        RECT 60.330 379.850 69.130 380.000 ;
        RECT 80.330 379.850 89.130 380.000 ;
        RECT 4.730 378.950 10.730 379.850 ;
        RECT 20.330 379.800 30.730 379.850 ;
        RECT 40.330 379.800 50.730 379.850 ;
        RECT 60.330 379.800 70.730 379.850 ;
        RECT 80.330 379.800 90.730 379.850 ;
        RECT 100.330 379.800 104.730 380.000 ;
        RECT 4.730 378.800 9.130 378.950 ;
        RECT 4.730 377.385 5.930 378.800 ;
        RECT 9.280 378.650 10.730 378.950 ;
        RECT 2.315 376.110 5.930 377.385 ;
        RECT 4.730 375.600 5.930 376.110 ;
        RECT 6.530 378.450 10.730 378.650 ;
        RECT 18.730 378.950 30.730 379.800 ;
        RECT 18.730 378.900 29.130 378.950 ;
        RECT 18.730 378.650 20.180 378.900 ;
        RECT 20.330 378.800 29.130 378.900 ;
        RECT 18.730 378.450 22.930 378.650 ;
        RECT 6.530 378.300 14.080 378.450 ;
        RECT 15.430 378.300 22.930 378.450 ;
        RECT 6.530 378.000 10.730 378.300 ;
        RECT 2.315 373.250 4.315 375.545 ;
        RECT 6.530 375.150 6.680 378.000 ;
        RECT 7.130 370.450 7.280 378.000 ;
        RECT 7.730 370.450 7.880 378.000 ;
        RECT 8.330 370.450 8.480 378.000 ;
        RECT 8.930 370.450 9.080 378.000 ;
        RECT 9.530 370.450 9.680 378.000 ;
        RECT 10.130 377.850 10.730 378.000 ;
        RECT 18.730 378.000 22.930 378.300 ;
        RECT 18.730 377.850 19.330 378.000 ;
        RECT 10.130 377.700 14.080 377.850 ;
        RECT 15.380 377.700 19.330 377.850 ;
        RECT 10.130 377.250 10.730 377.700 ;
        RECT 18.730 377.250 19.330 377.700 ;
        RECT 10.130 377.100 14.080 377.250 ;
        RECT 15.380 377.100 19.330 377.250 ;
        RECT 10.130 376.650 10.730 377.100 ;
        RECT 18.730 376.650 19.330 377.100 ;
        RECT 10.130 376.500 14.080 376.650 ;
        RECT 15.380 376.500 19.330 376.650 ;
        RECT 10.130 376.050 10.730 376.500 ;
        RECT 18.730 376.050 19.330 376.500 ;
        RECT 10.130 375.900 14.080 376.050 ;
        RECT 15.380 375.900 19.330 376.050 ;
        RECT 10.130 375.450 10.730 375.900 ;
        RECT 18.730 375.450 19.330 375.900 ;
        RECT 10.130 375.300 14.080 375.450 ;
        RECT 15.380 375.300 19.330 375.450 ;
        RECT 10.130 374.850 10.730 375.300 ;
        RECT 18.730 374.850 19.330 375.300 ;
        RECT 10.130 374.700 14.080 374.850 ;
        RECT 15.380 374.700 19.330 374.850 ;
        RECT 10.130 374.250 10.730 374.700 ;
        RECT 18.730 374.250 19.330 374.700 ;
        RECT 10.130 374.100 14.080 374.250 ;
        RECT 15.380 374.100 19.330 374.250 ;
        RECT 10.130 373.650 10.730 374.100 ;
        RECT 18.730 373.650 19.330 374.100 ;
        RECT 10.130 373.500 14.080 373.650 ;
        RECT 15.380 373.500 19.330 373.650 ;
        RECT 10.130 373.050 10.730 373.500 ;
        RECT 18.730 373.050 19.330 373.500 ;
        RECT 10.130 372.900 14.080 373.050 ;
        RECT 15.380 372.900 19.330 373.050 ;
        RECT 10.130 372.450 10.730 372.900 ;
        RECT 18.730 372.450 19.330 372.900 ;
        RECT 10.130 372.300 14.080 372.450 ;
        RECT 15.380 372.300 19.330 372.450 ;
        RECT 10.130 371.850 10.730 372.300 ;
        RECT 18.730 371.850 19.330 372.300 ;
        RECT 10.130 371.700 14.080 371.850 ;
        RECT 15.380 371.700 19.330 371.850 ;
        RECT 10.130 371.250 10.730 371.700 ;
        RECT 18.730 371.250 19.330 371.700 ;
        RECT 10.130 371.100 14.080 371.250 ;
        RECT 15.380 371.100 19.330 371.250 ;
        RECT 10.130 370.650 10.730 371.100 ;
        RECT 18.730 370.650 19.330 371.100 ;
        RECT 10.130 370.450 14.080 370.650 ;
        RECT 15.380 370.450 19.330 370.650 ;
        RECT 19.780 370.450 19.930 378.000 ;
        RECT 20.380 370.450 20.530 378.000 ;
        RECT 20.980 370.450 21.130 378.000 ;
        RECT 21.580 370.450 21.730 378.000 ;
        RECT 22.180 370.450 22.330 378.000 ;
        RECT 22.780 375.150 22.930 378.000 ;
        RECT 23.530 375.600 25.930 378.800 ;
        RECT 29.280 378.650 30.730 378.950 ;
        RECT 26.530 378.450 30.730 378.650 ;
        RECT 38.730 378.950 50.730 379.800 ;
        RECT 38.730 378.900 49.130 378.950 ;
        RECT 38.730 378.650 40.180 378.900 ;
        RECT 40.330 378.800 49.130 378.900 ;
        RECT 38.730 378.450 42.930 378.650 ;
        RECT 26.530 378.300 34.080 378.450 ;
        RECT 35.430 378.300 42.930 378.450 ;
        RECT 26.530 378.000 30.730 378.300 ;
        RECT 26.530 375.150 26.680 378.000 ;
        RECT 27.130 370.450 27.280 378.000 ;
        RECT 27.730 370.450 27.880 378.000 ;
        RECT 28.330 370.450 28.480 378.000 ;
        RECT 28.930 370.450 29.080 378.000 ;
        RECT 29.530 370.450 29.680 378.000 ;
        RECT 30.130 377.850 30.730 378.000 ;
        RECT 38.730 378.000 42.930 378.300 ;
        RECT 38.730 377.850 39.330 378.000 ;
        RECT 30.130 377.700 34.080 377.850 ;
        RECT 35.380 377.700 39.330 377.850 ;
        RECT 30.130 377.250 30.730 377.700 ;
        RECT 38.730 377.250 39.330 377.700 ;
        RECT 30.130 377.100 34.080 377.250 ;
        RECT 35.380 377.100 39.330 377.250 ;
        RECT 30.130 376.650 30.730 377.100 ;
        RECT 38.730 376.650 39.330 377.100 ;
        RECT 30.130 376.500 34.080 376.650 ;
        RECT 35.380 376.500 39.330 376.650 ;
        RECT 30.130 376.050 30.730 376.500 ;
        RECT 38.730 376.050 39.330 376.500 ;
        RECT 30.130 375.900 34.080 376.050 ;
        RECT 35.380 375.900 39.330 376.050 ;
        RECT 30.130 375.450 30.730 375.900 ;
        RECT 38.730 375.450 39.330 375.900 ;
        RECT 30.130 375.300 34.080 375.450 ;
        RECT 35.380 375.300 39.330 375.450 ;
        RECT 30.130 374.850 30.730 375.300 ;
        RECT 38.730 374.850 39.330 375.300 ;
        RECT 30.130 374.700 34.080 374.850 ;
        RECT 35.380 374.700 39.330 374.850 ;
        RECT 30.130 374.250 30.730 374.700 ;
        RECT 38.730 374.250 39.330 374.700 ;
        RECT 30.130 374.100 34.080 374.250 ;
        RECT 35.380 374.100 39.330 374.250 ;
        RECT 30.130 373.650 30.730 374.100 ;
        RECT 38.730 373.650 39.330 374.100 ;
        RECT 30.130 373.500 34.080 373.650 ;
        RECT 35.380 373.500 39.330 373.650 ;
        RECT 30.130 373.050 30.730 373.500 ;
        RECT 38.730 373.050 39.330 373.500 ;
        RECT 30.130 372.900 34.080 373.050 ;
        RECT 35.380 372.900 39.330 373.050 ;
        RECT 30.130 372.450 30.730 372.900 ;
        RECT 38.730 372.450 39.330 372.900 ;
        RECT 30.130 372.300 34.080 372.450 ;
        RECT 35.380 372.300 39.330 372.450 ;
        RECT 30.130 371.850 30.730 372.300 ;
        RECT 38.730 371.850 39.330 372.300 ;
        RECT 30.130 371.700 34.080 371.850 ;
        RECT 35.380 371.700 39.330 371.850 ;
        RECT 30.130 371.250 30.730 371.700 ;
        RECT 38.730 371.250 39.330 371.700 ;
        RECT 30.130 371.100 34.080 371.250 ;
        RECT 35.380 371.100 39.330 371.250 ;
        RECT 30.130 370.650 30.730 371.100 ;
        RECT 38.730 370.650 39.330 371.100 ;
        RECT 30.130 370.450 34.080 370.650 ;
        RECT 35.380 370.450 39.330 370.650 ;
        RECT 39.780 370.450 39.930 378.000 ;
        RECT 40.380 370.450 40.530 378.000 ;
        RECT 40.980 370.450 41.130 378.000 ;
        RECT 41.580 370.450 41.730 378.000 ;
        RECT 42.180 370.450 42.330 378.000 ;
        RECT 42.780 375.150 42.930 378.000 ;
        RECT 43.530 375.600 45.930 378.800 ;
        RECT 49.280 378.650 50.730 378.950 ;
        RECT 46.530 378.450 50.730 378.650 ;
        RECT 58.730 378.950 70.730 379.800 ;
        RECT 58.730 378.900 69.130 378.950 ;
        RECT 58.730 378.650 60.180 378.900 ;
        RECT 60.330 378.800 69.130 378.900 ;
        RECT 58.730 378.450 62.930 378.650 ;
        RECT 46.530 378.300 54.080 378.450 ;
        RECT 55.430 378.300 62.930 378.450 ;
        RECT 46.530 378.000 50.730 378.300 ;
        RECT 46.530 375.150 46.680 378.000 ;
        RECT 47.130 370.450 47.280 378.000 ;
        RECT 47.730 370.450 47.880 378.000 ;
        RECT 48.330 370.450 48.480 378.000 ;
        RECT 48.930 370.450 49.080 378.000 ;
        RECT 49.530 370.450 49.680 378.000 ;
        RECT 50.130 377.850 50.730 378.000 ;
        RECT 58.730 378.000 62.930 378.300 ;
        RECT 58.730 377.850 59.330 378.000 ;
        RECT 50.130 377.700 54.080 377.850 ;
        RECT 55.380 377.700 59.330 377.850 ;
        RECT 50.130 377.250 50.730 377.700 ;
        RECT 58.730 377.250 59.330 377.700 ;
        RECT 50.130 377.100 54.080 377.250 ;
        RECT 55.380 377.100 59.330 377.250 ;
        RECT 50.130 376.650 50.730 377.100 ;
        RECT 58.730 376.650 59.330 377.100 ;
        RECT 50.130 376.500 54.080 376.650 ;
        RECT 55.380 376.500 59.330 376.650 ;
        RECT 50.130 376.050 50.730 376.500 ;
        RECT 58.730 376.050 59.330 376.500 ;
        RECT 50.130 375.900 54.080 376.050 ;
        RECT 55.380 375.900 59.330 376.050 ;
        RECT 50.130 375.450 50.730 375.900 ;
        RECT 58.730 375.450 59.330 375.900 ;
        RECT 50.130 375.300 54.080 375.450 ;
        RECT 55.380 375.300 59.330 375.450 ;
        RECT 50.130 374.850 50.730 375.300 ;
        RECT 58.730 374.850 59.330 375.300 ;
        RECT 50.130 374.700 54.080 374.850 ;
        RECT 55.380 374.700 59.330 374.850 ;
        RECT 50.130 374.250 50.730 374.700 ;
        RECT 58.730 374.250 59.330 374.700 ;
        RECT 50.130 374.100 54.080 374.250 ;
        RECT 55.380 374.100 59.330 374.250 ;
        RECT 50.130 373.650 50.730 374.100 ;
        RECT 58.730 373.650 59.330 374.100 ;
        RECT 50.130 373.500 54.080 373.650 ;
        RECT 55.380 373.500 59.330 373.650 ;
        RECT 50.130 373.050 50.730 373.500 ;
        RECT 58.730 373.050 59.330 373.500 ;
        RECT 50.130 372.900 54.080 373.050 ;
        RECT 55.380 372.900 59.330 373.050 ;
        RECT 50.130 372.450 50.730 372.900 ;
        RECT 58.730 372.450 59.330 372.900 ;
        RECT 50.130 372.300 54.080 372.450 ;
        RECT 55.380 372.300 59.330 372.450 ;
        RECT 50.130 371.850 50.730 372.300 ;
        RECT 58.730 371.850 59.330 372.300 ;
        RECT 50.130 371.700 54.080 371.850 ;
        RECT 55.380 371.700 59.330 371.850 ;
        RECT 50.130 371.250 50.730 371.700 ;
        RECT 58.730 371.250 59.330 371.700 ;
        RECT 50.130 371.100 54.080 371.250 ;
        RECT 55.380 371.100 59.330 371.250 ;
        RECT 50.130 370.650 50.730 371.100 ;
        RECT 58.730 370.650 59.330 371.100 ;
        RECT 50.130 370.450 54.080 370.650 ;
        RECT 55.380 370.450 59.330 370.650 ;
        RECT 59.780 370.450 59.930 378.000 ;
        RECT 60.380 370.450 60.530 378.000 ;
        RECT 60.980 370.450 61.130 378.000 ;
        RECT 61.580 370.450 61.730 378.000 ;
        RECT 62.180 370.450 62.330 378.000 ;
        RECT 62.780 375.150 62.930 378.000 ;
        RECT 63.530 375.600 65.930 378.800 ;
        RECT 69.280 378.650 70.730 378.950 ;
        RECT 66.530 378.450 70.730 378.650 ;
        RECT 78.730 378.950 90.730 379.800 ;
        RECT 78.730 378.900 89.130 378.950 ;
        RECT 78.730 378.650 80.180 378.900 ;
        RECT 80.330 378.800 89.130 378.900 ;
        RECT 78.730 378.450 82.930 378.650 ;
        RECT 66.530 378.300 74.080 378.450 ;
        RECT 75.430 378.300 82.930 378.450 ;
        RECT 66.530 378.000 70.730 378.300 ;
        RECT 66.530 375.150 66.680 378.000 ;
        RECT 67.130 370.450 67.280 378.000 ;
        RECT 67.730 370.450 67.880 378.000 ;
        RECT 68.330 370.450 68.480 378.000 ;
        RECT 68.930 370.450 69.080 378.000 ;
        RECT 69.530 370.450 69.680 378.000 ;
        RECT 70.130 377.850 70.730 378.000 ;
        RECT 78.730 378.000 82.930 378.300 ;
        RECT 78.730 377.850 79.330 378.000 ;
        RECT 70.130 377.700 74.080 377.850 ;
        RECT 75.380 377.700 79.330 377.850 ;
        RECT 70.130 377.250 70.730 377.700 ;
        RECT 78.730 377.250 79.330 377.700 ;
        RECT 70.130 377.100 74.080 377.250 ;
        RECT 75.380 377.100 79.330 377.250 ;
        RECT 70.130 376.650 70.730 377.100 ;
        RECT 78.730 376.650 79.330 377.100 ;
        RECT 70.130 376.500 74.080 376.650 ;
        RECT 75.380 376.500 79.330 376.650 ;
        RECT 70.130 376.050 70.730 376.500 ;
        RECT 78.730 376.050 79.330 376.500 ;
        RECT 70.130 375.900 74.080 376.050 ;
        RECT 75.380 375.900 79.330 376.050 ;
        RECT 70.130 375.450 70.730 375.900 ;
        RECT 78.730 375.450 79.330 375.900 ;
        RECT 70.130 375.300 74.080 375.450 ;
        RECT 75.380 375.300 79.330 375.450 ;
        RECT 70.130 374.850 70.730 375.300 ;
        RECT 78.730 374.850 79.330 375.300 ;
        RECT 70.130 374.700 74.080 374.850 ;
        RECT 75.380 374.700 79.330 374.850 ;
        RECT 70.130 374.250 70.730 374.700 ;
        RECT 78.730 374.250 79.330 374.700 ;
        RECT 70.130 374.100 74.080 374.250 ;
        RECT 75.380 374.100 79.330 374.250 ;
        RECT 70.130 373.650 70.730 374.100 ;
        RECT 78.730 373.650 79.330 374.100 ;
        RECT 70.130 373.500 74.080 373.650 ;
        RECT 75.380 373.500 79.330 373.650 ;
        RECT 70.130 373.050 70.730 373.500 ;
        RECT 78.730 373.050 79.330 373.500 ;
        RECT 70.130 372.900 74.080 373.050 ;
        RECT 75.380 372.900 79.330 373.050 ;
        RECT 70.130 372.450 70.730 372.900 ;
        RECT 78.730 372.450 79.330 372.900 ;
        RECT 70.130 372.300 74.080 372.450 ;
        RECT 75.380 372.300 79.330 372.450 ;
        RECT 70.130 371.850 70.730 372.300 ;
        RECT 78.730 371.850 79.330 372.300 ;
        RECT 70.130 371.700 74.080 371.850 ;
        RECT 75.380 371.700 79.330 371.850 ;
        RECT 70.130 371.250 70.730 371.700 ;
        RECT 78.730 371.250 79.330 371.700 ;
        RECT 70.130 371.100 74.080 371.250 ;
        RECT 75.380 371.100 79.330 371.250 ;
        RECT 70.130 370.650 70.730 371.100 ;
        RECT 78.730 370.650 79.330 371.100 ;
        RECT 70.130 370.450 74.080 370.650 ;
        RECT 75.380 370.450 79.330 370.650 ;
        RECT 79.780 370.450 79.930 378.000 ;
        RECT 80.380 370.450 80.530 378.000 ;
        RECT 80.980 370.450 81.130 378.000 ;
        RECT 81.580 370.450 81.730 378.000 ;
        RECT 82.180 370.450 82.330 378.000 ;
        RECT 82.780 375.150 82.930 378.000 ;
        RECT 83.530 375.600 85.930 378.800 ;
        RECT 89.280 378.650 90.730 378.950 ;
        RECT 86.530 378.450 90.730 378.650 ;
        RECT 98.730 378.900 104.730 379.800 ;
        RECT 98.730 378.650 100.180 378.900 ;
        RECT 100.330 378.800 104.730 378.900 ;
        RECT 98.730 378.450 102.930 378.650 ;
        RECT 86.530 378.300 94.080 378.450 ;
        RECT 95.430 378.300 102.930 378.450 ;
        RECT 86.530 378.000 90.730 378.300 ;
        RECT 86.530 375.150 86.680 378.000 ;
        RECT 87.130 370.450 87.280 378.000 ;
        RECT 87.730 370.450 87.880 378.000 ;
        RECT 88.330 370.450 88.480 378.000 ;
        RECT 88.930 370.450 89.080 378.000 ;
        RECT 89.530 370.450 89.680 378.000 ;
        RECT 90.130 377.850 90.730 378.000 ;
        RECT 98.730 378.000 102.930 378.300 ;
        RECT 98.730 377.850 99.330 378.000 ;
        RECT 90.130 377.700 94.080 377.850 ;
        RECT 95.380 377.700 99.330 377.850 ;
        RECT 90.130 377.250 90.730 377.700 ;
        RECT 98.730 377.250 99.330 377.700 ;
        RECT 90.130 377.100 94.080 377.250 ;
        RECT 95.380 377.100 99.330 377.250 ;
        RECT 90.130 376.650 90.730 377.100 ;
        RECT 98.730 376.650 99.330 377.100 ;
        RECT 90.130 376.500 94.080 376.650 ;
        RECT 95.380 376.500 99.330 376.650 ;
        RECT 90.130 376.050 90.730 376.500 ;
        RECT 98.730 376.050 99.330 376.500 ;
        RECT 90.130 375.900 94.080 376.050 ;
        RECT 95.380 375.900 99.330 376.050 ;
        RECT 90.130 375.450 90.730 375.900 ;
        RECT 98.730 375.450 99.330 375.900 ;
        RECT 90.130 375.300 94.080 375.450 ;
        RECT 95.380 375.300 99.330 375.450 ;
        RECT 90.130 374.850 90.730 375.300 ;
        RECT 98.730 374.850 99.330 375.300 ;
        RECT 90.130 374.700 94.080 374.850 ;
        RECT 95.380 374.700 99.330 374.850 ;
        RECT 90.130 374.250 90.730 374.700 ;
        RECT 98.730 374.250 99.330 374.700 ;
        RECT 90.130 374.100 94.080 374.250 ;
        RECT 95.380 374.100 99.330 374.250 ;
        RECT 90.130 373.650 90.730 374.100 ;
        RECT 98.730 373.650 99.330 374.100 ;
        RECT 90.130 373.500 94.080 373.650 ;
        RECT 95.380 373.500 99.330 373.650 ;
        RECT 90.130 373.050 90.730 373.500 ;
        RECT 98.730 373.050 99.330 373.500 ;
        RECT 90.130 372.900 94.080 373.050 ;
        RECT 95.380 372.900 99.330 373.050 ;
        RECT 90.130 372.450 90.730 372.900 ;
        RECT 98.730 372.450 99.330 372.900 ;
        RECT 90.130 372.300 94.080 372.450 ;
        RECT 95.380 372.300 99.330 372.450 ;
        RECT 90.130 371.850 90.730 372.300 ;
        RECT 98.730 371.850 99.330 372.300 ;
        RECT 90.130 371.700 94.080 371.850 ;
        RECT 95.380 371.700 99.330 371.850 ;
        RECT 90.130 371.250 90.730 371.700 ;
        RECT 98.730 371.250 99.330 371.700 ;
        RECT 90.130 371.100 94.080 371.250 ;
        RECT 95.380 371.100 99.330 371.250 ;
        RECT 90.130 370.650 90.730 371.100 ;
        RECT 98.730 370.650 99.330 371.100 ;
        RECT 90.130 370.450 94.080 370.650 ;
        RECT 95.380 370.450 99.330 370.650 ;
        RECT 99.780 370.450 99.930 378.000 ;
        RECT 100.380 370.450 100.530 378.000 ;
        RECT 100.980 370.450 101.130 378.000 ;
        RECT 101.580 370.450 101.730 378.000 ;
        RECT 102.180 370.450 102.330 378.000 ;
        RECT 102.780 375.150 102.930 378.000 ;
        RECT 103.530 377.585 104.730 378.800 ;
        RECT 103.530 376.310 107.130 377.585 ;
        RECT 103.530 375.600 104.730 376.310 ;
        RECT 2.315 364.450 4.315 366.745 ;
        RECT 4.730 364.020 5.930 364.400 ;
        RECT 2.315 362.745 5.930 364.020 ;
        RECT 4.730 361.200 5.930 362.745 ;
        RECT 6.530 362.000 6.680 364.900 ;
        RECT 7.130 362.000 7.280 369.550 ;
        RECT 7.730 362.000 7.880 369.550 ;
        RECT 8.330 362.000 8.480 369.550 ;
        RECT 8.930 362.000 9.080 369.550 ;
        RECT 9.530 362.000 9.680 369.550 ;
        RECT 10.130 369.350 14.080 369.550 ;
        RECT 15.380 369.350 19.330 369.550 ;
        RECT 10.130 368.900 10.730 369.350 ;
        RECT 18.730 368.900 19.330 369.350 ;
        RECT 10.130 368.750 14.080 368.900 ;
        RECT 15.380 368.750 19.330 368.900 ;
        RECT 10.130 368.300 10.730 368.750 ;
        RECT 18.730 368.300 19.330 368.750 ;
        RECT 10.130 368.150 14.080 368.300 ;
        RECT 15.380 368.150 19.330 368.300 ;
        RECT 10.130 367.700 10.730 368.150 ;
        RECT 18.730 367.700 19.330 368.150 ;
        RECT 10.130 367.550 14.080 367.700 ;
        RECT 15.380 367.550 19.330 367.700 ;
        RECT 10.130 367.100 10.730 367.550 ;
        RECT 18.730 367.100 19.330 367.550 ;
        RECT 10.130 366.950 14.080 367.100 ;
        RECT 15.380 366.950 19.330 367.100 ;
        RECT 10.130 366.500 10.730 366.950 ;
        RECT 18.730 366.500 19.330 366.950 ;
        RECT 10.130 366.350 14.080 366.500 ;
        RECT 15.380 366.350 19.330 366.500 ;
        RECT 10.130 365.900 10.730 366.350 ;
        RECT 18.730 365.900 19.330 366.350 ;
        RECT 10.130 365.750 14.080 365.900 ;
        RECT 15.380 365.750 19.330 365.900 ;
        RECT 10.130 365.300 10.730 365.750 ;
        RECT 18.730 365.300 19.330 365.750 ;
        RECT 10.130 365.150 14.080 365.300 ;
        RECT 15.380 365.150 19.330 365.300 ;
        RECT 10.130 364.700 10.730 365.150 ;
        RECT 18.730 364.700 19.330 365.150 ;
        RECT 10.130 364.550 14.080 364.700 ;
        RECT 15.380 364.550 19.330 364.700 ;
        RECT 10.130 364.100 10.730 364.550 ;
        RECT 18.730 364.100 19.330 364.550 ;
        RECT 10.130 363.950 14.080 364.100 ;
        RECT 15.380 363.950 19.330 364.100 ;
        RECT 10.130 363.500 10.730 363.950 ;
        RECT 18.730 363.500 19.330 363.950 ;
        RECT 10.130 363.350 14.080 363.500 ;
        RECT 15.380 363.350 19.330 363.500 ;
        RECT 10.130 362.900 10.730 363.350 ;
        RECT 18.730 362.900 19.330 363.350 ;
        RECT 10.130 362.750 14.080 362.900 ;
        RECT 15.380 362.750 19.330 362.900 ;
        RECT 10.130 362.300 10.730 362.750 ;
        RECT 18.730 362.300 19.330 362.750 ;
        RECT 10.130 362.150 14.080 362.300 ;
        RECT 15.380 362.150 19.330 362.300 ;
        RECT 10.130 362.000 10.730 362.150 ;
        RECT 6.530 361.700 10.730 362.000 ;
        RECT 18.730 362.000 19.330 362.150 ;
        RECT 19.780 362.000 19.930 369.550 ;
        RECT 20.380 362.000 20.530 369.550 ;
        RECT 20.980 362.000 21.130 369.550 ;
        RECT 21.580 362.000 21.730 369.550 ;
        RECT 22.180 362.000 22.330 369.550 ;
        RECT 22.780 362.000 22.930 364.900 ;
        RECT 18.730 361.700 22.930 362.000 ;
        RECT 6.530 361.550 14.080 361.700 ;
        RECT 15.380 361.550 22.930 361.700 ;
        RECT 6.530 361.350 10.730 361.550 ;
        RECT 4.730 361.050 9.130 361.200 ;
        RECT 9.280 361.050 10.730 361.350 ;
        RECT 4.730 360.150 10.730 361.050 ;
        RECT 18.730 361.350 22.930 361.550 ;
        RECT 18.730 361.050 20.180 361.350 ;
        RECT 23.530 361.200 25.930 364.400 ;
        RECT 26.530 362.000 26.680 364.900 ;
        RECT 27.130 362.000 27.280 369.550 ;
        RECT 27.730 362.000 27.880 369.550 ;
        RECT 28.330 362.000 28.480 369.550 ;
        RECT 28.930 362.000 29.080 369.550 ;
        RECT 29.530 362.000 29.680 369.550 ;
        RECT 30.130 369.350 34.080 369.550 ;
        RECT 35.380 369.350 39.330 369.550 ;
        RECT 30.130 368.900 30.730 369.350 ;
        RECT 38.730 368.900 39.330 369.350 ;
        RECT 30.130 368.750 34.080 368.900 ;
        RECT 35.380 368.750 39.330 368.900 ;
        RECT 30.130 368.300 30.730 368.750 ;
        RECT 38.730 368.300 39.330 368.750 ;
        RECT 30.130 368.150 34.080 368.300 ;
        RECT 35.380 368.150 39.330 368.300 ;
        RECT 30.130 367.700 30.730 368.150 ;
        RECT 38.730 367.700 39.330 368.150 ;
        RECT 30.130 367.550 34.080 367.700 ;
        RECT 35.380 367.550 39.330 367.700 ;
        RECT 30.130 367.100 30.730 367.550 ;
        RECT 38.730 367.100 39.330 367.550 ;
        RECT 30.130 366.950 34.080 367.100 ;
        RECT 35.380 366.950 39.330 367.100 ;
        RECT 30.130 366.500 30.730 366.950 ;
        RECT 38.730 366.500 39.330 366.950 ;
        RECT 30.130 366.350 34.080 366.500 ;
        RECT 35.380 366.350 39.330 366.500 ;
        RECT 30.130 365.900 30.730 366.350 ;
        RECT 38.730 365.900 39.330 366.350 ;
        RECT 30.130 365.750 34.080 365.900 ;
        RECT 35.380 365.750 39.330 365.900 ;
        RECT 30.130 365.300 30.730 365.750 ;
        RECT 38.730 365.300 39.330 365.750 ;
        RECT 30.130 365.150 34.080 365.300 ;
        RECT 35.380 365.150 39.330 365.300 ;
        RECT 30.130 364.700 30.730 365.150 ;
        RECT 38.730 364.700 39.330 365.150 ;
        RECT 30.130 364.550 34.080 364.700 ;
        RECT 35.380 364.550 39.330 364.700 ;
        RECT 30.130 364.100 30.730 364.550 ;
        RECT 38.730 364.100 39.330 364.550 ;
        RECT 30.130 363.950 34.080 364.100 ;
        RECT 35.380 363.950 39.330 364.100 ;
        RECT 30.130 363.500 30.730 363.950 ;
        RECT 38.730 363.500 39.330 363.950 ;
        RECT 30.130 363.350 34.080 363.500 ;
        RECT 35.380 363.350 39.330 363.500 ;
        RECT 30.130 362.900 30.730 363.350 ;
        RECT 38.730 362.900 39.330 363.350 ;
        RECT 30.130 362.750 34.080 362.900 ;
        RECT 35.380 362.750 39.330 362.900 ;
        RECT 30.130 362.300 30.730 362.750 ;
        RECT 38.730 362.300 39.330 362.750 ;
        RECT 30.130 362.150 34.080 362.300 ;
        RECT 35.380 362.150 39.330 362.300 ;
        RECT 30.130 362.000 30.730 362.150 ;
        RECT 26.530 361.700 30.730 362.000 ;
        RECT 38.730 362.000 39.330 362.150 ;
        RECT 39.780 362.000 39.930 369.550 ;
        RECT 40.380 362.000 40.530 369.550 ;
        RECT 40.980 362.000 41.130 369.550 ;
        RECT 41.580 362.000 41.730 369.550 ;
        RECT 42.180 362.000 42.330 369.550 ;
        RECT 42.780 362.000 42.930 364.900 ;
        RECT 38.730 361.700 42.930 362.000 ;
        RECT 26.530 361.550 34.080 361.700 ;
        RECT 35.380 361.550 42.930 361.700 ;
        RECT 26.530 361.350 30.730 361.550 ;
        RECT 20.330 361.050 29.130 361.200 ;
        RECT 29.280 361.050 30.730 361.350 ;
        RECT 18.730 360.150 30.730 361.050 ;
        RECT 38.730 361.350 42.930 361.550 ;
        RECT 38.730 361.050 40.180 361.350 ;
        RECT 43.530 361.200 45.930 364.400 ;
        RECT 46.530 362.000 46.680 364.900 ;
        RECT 47.130 362.000 47.280 369.550 ;
        RECT 47.730 362.000 47.880 369.550 ;
        RECT 48.330 362.000 48.480 369.550 ;
        RECT 48.930 362.000 49.080 369.550 ;
        RECT 49.530 362.000 49.680 369.550 ;
        RECT 50.130 369.350 54.080 369.550 ;
        RECT 55.380 369.350 59.330 369.550 ;
        RECT 50.130 368.900 50.730 369.350 ;
        RECT 58.730 368.900 59.330 369.350 ;
        RECT 50.130 368.750 54.080 368.900 ;
        RECT 55.380 368.750 59.330 368.900 ;
        RECT 50.130 368.300 50.730 368.750 ;
        RECT 58.730 368.300 59.330 368.750 ;
        RECT 50.130 368.150 54.080 368.300 ;
        RECT 55.380 368.150 59.330 368.300 ;
        RECT 50.130 367.700 50.730 368.150 ;
        RECT 58.730 367.700 59.330 368.150 ;
        RECT 50.130 367.550 54.080 367.700 ;
        RECT 55.380 367.550 59.330 367.700 ;
        RECT 50.130 367.100 50.730 367.550 ;
        RECT 58.730 367.100 59.330 367.550 ;
        RECT 50.130 366.950 54.080 367.100 ;
        RECT 55.380 366.950 59.330 367.100 ;
        RECT 50.130 366.500 50.730 366.950 ;
        RECT 58.730 366.500 59.330 366.950 ;
        RECT 50.130 366.350 54.080 366.500 ;
        RECT 55.380 366.350 59.330 366.500 ;
        RECT 50.130 365.900 50.730 366.350 ;
        RECT 58.730 365.900 59.330 366.350 ;
        RECT 50.130 365.750 54.080 365.900 ;
        RECT 55.380 365.750 59.330 365.900 ;
        RECT 50.130 365.300 50.730 365.750 ;
        RECT 58.730 365.300 59.330 365.750 ;
        RECT 50.130 365.150 54.080 365.300 ;
        RECT 55.380 365.150 59.330 365.300 ;
        RECT 50.130 364.700 50.730 365.150 ;
        RECT 58.730 364.700 59.330 365.150 ;
        RECT 50.130 364.550 54.080 364.700 ;
        RECT 55.380 364.550 59.330 364.700 ;
        RECT 50.130 364.100 50.730 364.550 ;
        RECT 58.730 364.100 59.330 364.550 ;
        RECT 50.130 363.950 54.080 364.100 ;
        RECT 55.380 363.950 59.330 364.100 ;
        RECT 50.130 363.500 50.730 363.950 ;
        RECT 58.730 363.500 59.330 363.950 ;
        RECT 50.130 363.350 54.080 363.500 ;
        RECT 55.380 363.350 59.330 363.500 ;
        RECT 50.130 362.900 50.730 363.350 ;
        RECT 58.730 362.900 59.330 363.350 ;
        RECT 50.130 362.750 54.080 362.900 ;
        RECT 55.380 362.750 59.330 362.900 ;
        RECT 50.130 362.300 50.730 362.750 ;
        RECT 58.730 362.300 59.330 362.750 ;
        RECT 50.130 362.150 54.080 362.300 ;
        RECT 55.380 362.150 59.330 362.300 ;
        RECT 50.130 362.000 50.730 362.150 ;
        RECT 46.530 361.700 50.730 362.000 ;
        RECT 58.730 362.000 59.330 362.150 ;
        RECT 59.780 362.000 59.930 369.550 ;
        RECT 60.380 362.000 60.530 369.550 ;
        RECT 60.980 362.000 61.130 369.550 ;
        RECT 61.580 362.000 61.730 369.550 ;
        RECT 62.180 362.000 62.330 369.550 ;
        RECT 62.780 362.000 62.930 364.900 ;
        RECT 58.730 361.700 62.930 362.000 ;
        RECT 46.530 361.550 54.080 361.700 ;
        RECT 55.380 361.550 62.930 361.700 ;
        RECT 46.530 361.350 50.730 361.550 ;
        RECT 40.330 361.050 49.130 361.200 ;
        RECT 49.280 361.050 50.730 361.350 ;
        RECT 38.730 360.150 50.730 361.050 ;
        RECT 58.730 361.350 62.930 361.550 ;
        RECT 58.730 361.050 60.180 361.350 ;
        RECT 63.530 361.200 65.930 364.400 ;
        RECT 66.530 362.000 66.680 364.900 ;
        RECT 67.130 362.000 67.280 369.550 ;
        RECT 67.730 362.000 67.880 369.550 ;
        RECT 68.330 362.000 68.480 369.550 ;
        RECT 68.930 362.000 69.080 369.550 ;
        RECT 69.530 362.000 69.680 369.550 ;
        RECT 70.130 369.350 74.080 369.550 ;
        RECT 75.380 369.350 79.330 369.550 ;
        RECT 70.130 368.900 70.730 369.350 ;
        RECT 78.730 368.900 79.330 369.350 ;
        RECT 70.130 368.750 74.080 368.900 ;
        RECT 75.380 368.750 79.330 368.900 ;
        RECT 70.130 368.300 70.730 368.750 ;
        RECT 78.730 368.300 79.330 368.750 ;
        RECT 70.130 368.150 74.080 368.300 ;
        RECT 75.380 368.150 79.330 368.300 ;
        RECT 70.130 367.700 70.730 368.150 ;
        RECT 78.730 367.700 79.330 368.150 ;
        RECT 70.130 367.550 74.080 367.700 ;
        RECT 75.380 367.550 79.330 367.700 ;
        RECT 70.130 367.100 70.730 367.550 ;
        RECT 78.730 367.100 79.330 367.550 ;
        RECT 70.130 366.950 74.080 367.100 ;
        RECT 75.380 366.950 79.330 367.100 ;
        RECT 70.130 366.500 70.730 366.950 ;
        RECT 78.730 366.500 79.330 366.950 ;
        RECT 70.130 366.350 74.080 366.500 ;
        RECT 75.380 366.350 79.330 366.500 ;
        RECT 70.130 365.900 70.730 366.350 ;
        RECT 78.730 365.900 79.330 366.350 ;
        RECT 70.130 365.750 74.080 365.900 ;
        RECT 75.380 365.750 79.330 365.900 ;
        RECT 70.130 365.300 70.730 365.750 ;
        RECT 78.730 365.300 79.330 365.750 ;
        RECT 70.130 365.150 74.080 365.300 ;
        RECT 75.380 365.150 79.330 365.300 ;
        RECT 70.130 364.700 70.730 365.150 ;
        RECT 78.730 364.700 79.330 365.150 ;
        RECT 70.130 364.550 74.080 364.700 ;
        RECT 75.380 364.550 79.330 364.700 ;
        RECT 70.130 364.100 70.730 364.550 ;
        RECT 78.730 364.100 79.330 364.550 ;
        RECT 70.130 363.950 74.080 364.100 ;
        RECT 75.380 363.950 79.330 364.100 ;
        RECT 70.130 363.500 70.730 363.950 ;
        RECT 78.730 363.500 79.330 363.950 ;
        RECT 70.130 363.350 74.080 363.500 ;
        RECT 75.380 363.350 79.330 363.500 ;
        RECT 70.130 362.900 70.730 363.350 ;
        RECT 78.730 362.900 79.330 363.350 ;
        RECT 70.130 362.750 74.080 362.900 ;
        RECT 75.380 362.750 79.330 362.900 ;
        RECT 70.130 362.300 70.730 362.750 ;
        RECT 78.730 362.300 79.330 362.750 ;
        RECT 70.130 362.150 74.080 362.300 ;
        RECT 75.380 362.150 79.330 362.300 ;
        RECT 70.130 362.000 70.730 362.150 ;
        RECT 66.530 361.700 70.730 362.000 ;
        RECT 78.730 362.000 79.330 362.150 ;
        RECT 79.780 362.000 79.930 369.550 ;
        RECT 80.380 362.000 80.530 369.550 ;
        RECT 80.980 362.000 81.130 369.550 ;
        RECT 81.580 362.000 81.730 369.550 ;
        RECT 82.180 362.000 82.330 369.550 ;
        RECT 82.780 362.000 82.930 364.900 ;
        RECT 78.730 361.700 82.930 362.000 ;
        RECT 66.530 361.550 74.080 361.700 ;
        RECT 75.380 361.550 82.930 361.700 ;
        RECT 66.530 361.350 70.730 361.550 ;
        RECT 60.330 361.050 69.130 361.200 ;
        RECT 69.280 361.050 70.730 361.350 ;
        RECT 58.730 360.150 70.730 361.050 ;
        RECT 78.730 361.350 82.930 361.550 ;
        RECT 78.730 361.050 80.180 361.350 ;
        RECT 83.530 361.200 85.930 364.400 ;
        RECT 86.530 362.000 86.680 364.900 ;
        RECT 87.130 362.000 87.280 369.550 ;
        RECT 87.730 362.000 87.880 369.550 ;
        RECT 88.330 362.000 88.480 369.550 ;
        RECT 88.930 362.000 89.080 369.550 ;
        RECT 89.530 362.000 89.680 369.550 ;
        RECT 90.130 369.350 94.080 369.550 ;
        RECT 95.380 369.350 99.330 369.550 ;
        RECT 90.130 368.900 90.730 369.350 ;
        RECT 98.730 368.900 99.330 369.350 ;
        RECT 90.130 368.750 94.080 368.900 ;
        RECT 95.380 368.750 99.330 368.900 ;
        RECT 90.130 368.300 90.730 368.750 ;
        RECT 98.730 368.300 99.330 368.750 ;
        RECT 90.130 368.150 94.080 368.300 ;
        RECT 95.380 368.150 99.330 368.300 ;
        RECT 90.130 367.700 90.730 368.150 ;
        RECT 98.730 367.700 99.330 368.150 ;
        RECT 90.130 367.550 94.080 367.700 ;
        RECT 95.380 367.550 99.330 367.700 ;
        RECT 90.130 367.100 90.730 367.550 ;
        RECT 98.730 367.100 99.330 367.550 ;
        RECT 90.130 366.950 94.080 367.100 ;
        RECT 95.380 366.950 99.330 367.100 ;
        RECT 90.130 366.500 90.730 366.950 ;
        RECT 98.730 366.500 99.330 366.950 ;
        RECT 90.130 366.350 94.080 366.500 ;
        RECT 95.380 366.350 99.330 366.500 ;
        RECT 90.130 365.900 90.730 366.350 ;
        RECT 98.730 365.900 99.330 366.350 ;
        RECT 90.130 365.750 94.080 365.900 ;
        RECT 95.380 365.750 99.330 365.900 ;
        RECT 90.130 365.300 90.730 365.750 ;
        RECT 98.730 365.300 99.330 365.750 ;
        RECT 90.130 365.150 94.080 365.300 ;
        RECT 95.380 365.150 99.330 365.300 ;
        RECT 90.130 364.700 90.730 365.150 ;
        RECT 98.730 364.700 99.330 365.150 ;
        RECT 90.130 364.550 94.080 364.700 ;
        RECT 95.380 364.550 99.330 364.700 ;
        RECT 90.130 364.100 90.730 364.550 ;
        RECT 98.730 364.100 99.330 364.550 ;
        RECT 90.130 363.950 94.080 364.100 ;
        RECT 95.380 363.950 99.330 364.100 ;
        RECT 90.130 363.500 90.730 363.950 ;
        RECT 98.730 363.500 99.330 363.950 ;
        RECT 90.130 363.350 94.080 363.500 ;
        RECT 95.380 363.350 99.330 363.500 ;
        RECT 90.130 362.900 90.730 363.350 ;
        RECT 98.730 362.900 99.330 363.350 ;
        RECT 90.130 362.750 94.080 362.900 ;
        RECT 95.380 362.750 99.330 362.900 ;
        RECT 90.130 362.300 90.730 362.750 ;
        RECT 98.730 362.300 99.330 362.750 ;
        RECT 90.130 362.150 94.080 362.300 ;
        RECT 95.380 362.150 99.330 362.300 ;
        RECT 90.130 362.000 90.730 362.150 ;
        RECT 86.530 361.700 90.730 362.000 ;
        RECT 98.730 362.000 99.330 362.150 ;
        RECT 99.780 362.000 99.930 369.550 ;
        RECT 100.380 362.000 100.530 369.550 ;
        RECT 100.980 362.000 101.130 369.550 ;
        RECT 101.580 362.000 101.730 369.550 ;
        RECT 102.180 362.000 102.330 369.550 ;
        RECT 102.780 362.000 102.930 364.900 ;
        RECT 98.730 361.700 102.930 362.000 ;
        RECT 86.530 361.550 94.080 361.700 ;
        RECT 95.380 361.550 102.930 361.700 ;
        RECT 86.530 361.350 90.730 361.550 ;
        RECT 80.330 361.050 89.130 361.200 ;
        RECT 89.280 361.050 90.730 361.350 ;
        RECT 78.730 360.150 90.730 361.050 ;
        RECT 98.730 361.350 102.930 361.550 ;
        RECT 103.530 363.600 104.730 364.400 ;
        RECT 103.530 362.325 107.140 363.600 ;
        RECT 98.730 361.050 100.180 361.350 ;
        RECT 103.530 361.200 104.730 362.325 ;
        RECT 100.330 361.050 104.730 361.200 ;
        RECT 98.730 360.150 104.730 361.050 ;
        RECT 4.730 359.850 9.130 360.150 ;
        RECT 20.330 359.850 29.130 360.150 ;
        RECT 40.330 359.850 49.130 360.150 ;
        RECT 60.330 359.850 69.130 360.150 ;
        RECT 80.330 359.850 89.130 360.150 ;
        RECT 4.730 358.950 10.730 359.850 ;
        RECT 20.330 359.800 30.730 359.850 ;
        RECT 40.330 359.800 50.730 359.850 ;
        RECT 60.330 359.800 70.730 359.850 ;
        RECT 80.330 359.800 90.730 359.850 ;
        RECT 100.330 359.800 104.730 360.150 ;
        RECT 4.730 358.800 9.130 358.950 ;
        RECT 4.730 357.385 5.930 358.800 ;
        RECT 9.280 358.650 10.730 358.950 ;
        RECT 2.315 356.110 5.930 357.385 ;
        RECT 4.730 355.600 5.930 356.110 ;
        RECT 6.530 358.450 10.730 358.650 ;
        RECT 18.730 358.950 30.730 359.800 ;
        RECT 18.730 358.900 29.130 358.950 ;
        RECT 18.730 358.650 20.180 358.900 ;
        RECT 20.330 358.800 29.130 358.900 ;
        RECT 18.730 358.450 22.930 358.650 ;
        RECT 6.530 358.300 14.080 358.450 ;
        RECT 15.430 358.300 22.930 358.450 ;
        RECT 6.530 358.000 10.730 358.300 ;
        RECT 2.315 353.250 4.315 355.545 ;
        RECT 6.530 355.150 6.680 358.000 ;
        RECT 7.130 350.450 7.280 358.000 ;
        RECT 7.730 350.450 7.880 358.000 ;
        RECT 8.330 350.450 8.480 358.000 ;
        RECT 8.930 350.450 9.080 358.000 ;
        RECT 9.530 350.450 9.680 358.000 ;
        RECT 10.130 357.850 10.730 358.000 ;
        RECT 18.730 358.000 22.930 358.300 ;
        RECT 18.730 357.850 19.330 358.000 ;
        RECT 10.130 357.700 14.080 357.850 ;
        RECT 15.380 357.700 19.330 357.850 ;
        RECT 10.130 357.250 10.730 357.700 ;
        RECT 18.730 357.250 19.330 357.700 ;
        RECT 10.130 357.100 14.080 357.250 ;
        RECT 15.380 357.100 19.330 357.250 ;
        RECT 10.130 356.650 10.730 357.100 ;
        RECT 18.730 356.650 19.330 357.100 ;
        RECT 10.130 356.500 14.080 356.650 ;
        RECT 15.380 356.500 19.330 356.650 ;
        RECT 10.130 356.050 10.730 356.500 ;
        RECT 18.730 356.050 19.330 356.500 ;
        RECT 10.130 355.900 14.080 356.050 ;
        RECT 15.380 355.900 19.330 356.050 ;
        RECT 10.130 355.450 10.730 355.900 ;
        RECT 18.730 355.450 19.330 355.900 ;
        RECT 10.130 355.300 14.080 355.450 ;
        RECT 15.380 355.300 19.330 355.450 ;
        RECT 10.130 354.850 10.730 355.300 ;
        RECT 18.730 354.850 19.330 355.300 ;
        RECT 10.130 354.700 14.080 354.850 ;
        RECT 15.380 354.700 19.330 354.850 ;
        RECT 10.130 354.250 10.730 354.700 ;
        RECT 18.730 354.250 19.330 354.700 ;
        RECT 10.130 354.100 14.080 354.250 ;
        RECT 15.380 354.100 19.330 354.250 ;
        RECT 10.130 353.650 10.730 354.100 ;
        RECT 18.730 353.650 19.330 354.100 ;
        RECT 10.130 353.500 14.080 353.650 ;
        RECT 15.380 353.500 19.330 353.650 ;
        RECT 10.130 353.050 10.730 353.500 ;
        RECT 18.730 353.050 19.330 353.500 ;
        RECT 10.130 352.900 14.080 353.050 ;
        RECT 15.380 352.900 19.330 353.050 ;
        RECT 10.130 352.450 10.730 352.900 ;
        RECT 18.730 352.450 19.330 352.900 ;
        RECT 10.130 352.300 14.080 352.450 ;
        RECT 15.380 352.300 19.330 352.450 ;
        RECT 10.130 351.850 10.730 352.300 ;
        RECT 18.730 351.850 19.330 352.300 ;
        RECT 10.130 351.700 14.080 351.850 ;
        RECT 15.380 351.700 19.330 351.850 ;
        RECT 10.130 351.250 10.730 351.700 ;
        RECT 18.730 351.250 19.330 351.700 ;
        RECT 10.130 351.100 14.080 351.250 ;
        RECT 15.380 351.100 19.330 351.250 ;
        RECT 10.130 350.650 10.730 351.100 ;
        RECT 18.730 350.650 19.330 351.100 ;
        RECT 10.130 350.450 14.080 350.650 ;
        RECT 15.380 350.450 19.330 350.650 ;
        RECT 19.780 350.450 19.930 358.000 ;
        RECT 20.380 350.450 20.530 358.000 ;
        RECT 20.980 350.450 21.130 358.000 ;
        RECT 21.580 350.450 21.730 358.000 ;
        RECT 22.180 350.450 22.330 358.000 ;
        RECT 22.780 355.150 22.930 358.000 ;
        RECT 23.530 355.600 25.930 358.800 ;
        RECT 29.280 358.650 30.730 358.950 ;
        RECT 26.530 358.450 30.730 358.650 ;
        RECT 38.730 358.950 50.730 359.800 ;
        RECT 38.730 358.900 49.130 358.950 ;
        RECT 38.730 358.650 40.180 358.900 ;
        RECT 40.330 358.800 49.130 358.900 ;
        RECT 38.730 358.450 42.930 358.650 ;
        RECT 26.530 358.300 34.080 358.450 ;
        RECT 35.430 358.300 42.930 358.450 ;
        RECT 26.530 358.000 30.730 358.300 ;
        RECT 26.530 355.150 26.680 358.000 ;
        RECT 27.130 350.450 27.280 358.000 ;
        RECT 27.730 350.450 27.880 358.000 ;
        RECT 28.330 350.450 28.480 358.000 ;
        RECT 28.930 350.450 29.080 358.000 ;
        RECT 29.530 350.450 29.680 358.000 ;
        RECT 30.130 357.850 30.730 358.000 ;
        RECT 38.730 358.000 42.930 358.300 ;
        RECT 38.730 357.850 39.330 358.000 ;
        RECT 30.130 357.700 34.080 357.850 ;
        RECT 35.380 357.700 39.330 357.850 ;
        RECT 30.130 357.250 30.730 357.700 ;
        RECT 38.730 357.250 39.330 357.700 ;
        RECT 30.130 357.100 34.080 357.250 ;
        RECT 35.380 357.100 39.330 357.250 ;
        RECT 30.130 356.650 30.730 357.100 ;
        RECT 38.730 356.650 39.330 357.100 ;
        RECT 30.130 356.500 34.080 356.650 ;
        RECT 35.380 356.500 39.330 356.650 ;
        RECT 30.130 356.050 30.730 356.500 ;
        RECT 38.730 356.050 39.330 356.500 ;
        RECT 30.130 355.900 34.080 356.050 ;
        RECT 35.380 355.900 39.330 356.050 ;
        RECT 30.130 355.450 30.730 355.900 ;
        RECT 38.730 355.450 39.330 355.900 ;
        RECT 30.130 355.300 34.080 355.450 ;
        RECT 35.380 355.300 39.330 355.450 ;
        RECT 30.130 354.850 30.730 355.300 ;
        RECT 38.730 354.850 39.330 355.300 ;
        RECT 30.130 354.700 34.080 354.850 ;
        RECT 35.380 354.700 39.330 354.850 ;
        RECT 30.130 354.250 30.730 354.700 ;
        RECT 38.730 354.250 39.330 354.700 ;
        RECT 30.130 354.100 34.080 354.250 ;
        RECT 35.380 354.100 39.330 354.250 ;
        RECT 30.130 353.650 30.730 354.100 ;
        RECT 38.730 353.650 39.330 354.100 ;
        RECT 30.130 353.500 34.080 353.650 ;
        RECT 35.380 353.500 39.330 353.650 ;
        RECT 30.130 353.050 30.730 353.500 ;
        RECT 38.730 353.050 39.330 353.500 ;
        RECT 30.130 352.900 34.080 353.050 ;
        RECT 35.380 352.900 39.330 353.050 ;
        RECT 30.130 352.450 30.730 352.900 ;
        RECT 38.730 352.450 39.330 352.900 ;
        RECT 30.130 352.300 34.080 352.450 ;
        RECT 35.380 352.300 39.330 352.450 ;
        RECT 30.130 351.850 30.730 352.300 ;
        RECT 38.730 351.850 39.330 352.300 ;
        RECT 30.130 351.700 34.080 351.850 ;
        RECT 35.380 351.700 39.330 351.850 ;
        RECT 30.130 351.250 30.730 351.700 ;
        RECT 38.730 351.250 39.330 351.700 ;
        RECT 30.130 351.100 34.080 351.250 ;
        RECT 35.380 351.100 39.330 351.250 ;
        RECT 30.130 350.650 30.730 351.100 ;
        RECT 38.730 350.650 39.330 351.100 ;
        RECT 30.130 350.450 34.080 350.650 ;
        RECT 35.380 350.450 39.330 350.650 ;
        RECT 39.780 350.450 39.930 358.000 ;
        RECT 40.380 350.450 40.530 358.000 ;
        RECT 40.980 350.450 41.130 358.000 ;
        RECT 41.580 350.450 41.730 358.000 ;
        RECT 42.180 350.450 42.330 358.000 ;
        RECT 42.780 355.150 42.930 358.000 ;
        RECT 43.530 355.600 45.930 358.800 ;
        RECT 49.280 358.650 50.730 358.950 ;
        RECT 46.530 358.450 50.730 358.650 ;
        RECT 58.730 358.950 70.730 359.800 ;
        RECT 58.730 358.900 69.130 358.950 ;
        RECT 58.730 358.650 60.180 358.900 ;
        RECT 60.330 358.800 69.130 358.900 ;
        RECT 58.730 358.450 62.930 358.650 ;
        RECT 46.530 358.300 54.080 358.450 ;
        RECT 55.430 358.300 62.930 358.450 ;
        RECT 46.530 358.000 50.730 358.300 ;
        RECT 46.530 355.150 46.680 358.000 ;
        RECT 47.130 350.450 47.280 358.000 ;
        RECT 47.730 350.450 47.880 358.000 ;
        RECT 48.330 350.450 48.480 358.000 ;
        RECT 48.930 350.450 49.080 358.000 ;
        RECT 49.530 350.450 49.680 358.000 ;
        RECT 50.130 357.850 50.730 358.000 ;
        RECT 58.730 358.000 62.930 358.300 ;
        RECT 58.730 357.850 59.330 358.000 ;
        RECT 50.130 357.700 54.080 357.850 ;
        RECT 55.380 357.700 59.330 357.850 ;
        RECT 50.130 357.250 50.730 357.700 ;
        RECT 58.730 357.250 59.330 357.700 ;
        RECT 50.130 357.100 54.080 357.250 ;
        RECT 55.380 357.100 59.330 357.250 ;
        RECT 50.130 356.650 50.730 357.100 ;
        RECT 58.730 356.650 59.330 357.100 ;
        RECT 50.130 356.500 54.080 356.650 ;
        RECT 55.380 356.500 59.330 356.650 ;
        RECT 50.130 356.050 50.730 356.500 ;
        RECT 58.730 356.050 59.330 356.500 ;
        RECT 50.130 355.900 54.080 356.050 ;
        RECT 55.380 355.900 59.330 356.050 ;
        RECT 50.130 355.450 50.730 355.900 ;
        RECT 58.730 355.450 59.330 355.900 ;
        RECT 50.130 355.300 54.080 355.450 ;
        RECT 55.380 355.300 59.330 355.450 ;
        RECT 50.130 354.850 50.730 355.300 ;
        RECT 58.730 354.850 59.330 355.300 ;
        RECT 50.130 354.700 54.080 354.850 ;
        RECT 55.380 354.700 59.330 354.850 ;
        RECT 50.130 354.250 50.730 354.700 ;
        RECT 58.730 354.250 59.330 354.700 ;
        RECT 50.130 354.100 54.080 354.250 ;
        RECT 55.380 354.100 59.330 354.250 ;
        RECT 50.130 353.650 50.730 354.100 ;
        RECT 58.730 353.650 59.330 354.100 ;
        RECT 50.130 353.500 54.080 353.650 ;
        RECT 55.380 353.500 59.330 353.650 ;
        RECT 50.130 353.050 50.730 353.500 ;
        RECT 58.730 353.050 59.330 353.500 ;
        RECT 50.130 352.900 54.080 353.050 ;
        RECT 55.380 352.900 59.330 353.050 ;
        RECT 50.130 352.450 50.730 352.900 ;
        RECT 58.730 352.450 59.330 352.900 ;
        RECT 50.130 352.300 54.080 352.450 ;
        RECT 55.380 352.300 59.330 352.450 ;
        RECT 50.130 351.850 50.730 352.300 ;
        RECT 58.730 351.850 59.330 352.300 ;
        RECT 50.130 351.700 54.080 351.850 ;
        RECT 55.380 351.700 59.330 351.850 ;
        RECT 50.130 351.250 50.730 351.700 ;
        RECT 58.730 351.250 59.330 351.700 ;
        RECT 50.130 351.100 54.080 351.250 ;
        RECT 55.380 351.100 59.330 351.250 ;
        RECT 50.130 350.650 50.730 351.100 ;
        RECT 58.730 350.650 59.330 351.100 ;
        RECT 50.130 350.450 54.080 350.650 ;
        RECT 55.380 350.450 59.330 350.650 ;
        RECT 59.780 350.450 59.930 358.000 ;
        RECT 60.380 350.450 60.530 358.000 ;
        RECT 60.980 350.450 61.130 358.000 ;
        RECT 61.580 350.450 61.730 358.000 ;
        RECT 62.180 350.450 62.330 358.000 ;
        RECT 62.780 355.150 62.930 358.000 ;
        RECT 63.530 355.600 65.930 358.800 ;
        RECT 69.280 358.650 70.730 358.950 ;
        RECT 66.530 358.450 70.730 358.650 ;
        RECT 78.730 358.950 90.730 359.800 ;
        RECT 78.730 358.900 89.130 358.950 ;
        RECT 78.730 358.650 80.180 358.900 ;
        RECT 80.330 358.800 89.130 358.900 ;
        RECT 78.730 358.450 82.930 358.650 ;
        RECT 66.530 358.300 74.080 358.450 ;
        RECT 75.430 358.300 82.930 358.450 ;
        RECT 66.530 358.000 70.730 358.300 ;
        RECT 66.530 355.150 66.680 358.000 ;
        RECT 67.130 350.450 67.280 358.000 ;
        RECT 67.730 350.450 67.880 358.000 ;
        RECT 68.330 350.450 68.480 358.000 ;
        RECT 68.930 350.450 69.080 358.000 ;
        RECT 69.530 350.450 69.680 358.000 ;
        RECT 70.130 357.850 70.730 358.000 ;
        RECT 78.730 358.000 82.930 358.300 ;
        RECT 78.730 357.850 79.330 358.000 ;
        RECT 70.130 357.700 74.080 357.850 ;
        RECT 75.380 357.700 79.330 357.850 ;
        RECT 70.130 357.250 70.730 357.700 ;
        RECT 78.730 357.250 79.330 357.700 ;
        RECT 70.130 357.100 74.080 357.250 ;
        RECT 75.380 357.100 79.330 357.250 ;
        RECT 70.130 356.650 70.730 357.100 ;
        RECT 78.730 356.650 79.330 357.100 ;
        RECT 70.130 356.500 74.080 356.650 ;
        RECT 75.380 356.500 79.330 356.650 ;
        RECT 70.130 356.050 70.730 356.500 ;
        RECT 78.730 356.050 79.330 356.500 ;
        RECT 70.130 355.900 74.080 356.050 ;
        RECT 75.380 355.900 79.330 356.050 ;
        RECT 70.130 355.450 70.730 355.900 ;
        RECT 78.730 355.450 79.330 355.900 ;
        RECT 70.130 355.300 74.080 355.450 ;
        RECT 75.380 355.300 79.330 355.450 ;
        RECT 70.130 354.850 70.730 355.300 ;
        RECT 78.730 354.850 79.330 355.300 ;
        RECT 70.130 354.700 74.080 354.850 ;
        RECT 75.380 354.700 79.330 354.850 ;
        RECT 70.130 354.250 70.730 354.700 ;
        RECT 78.730 354.250 79.330 354.700 ;
        RECT 70.130 354.100 74.080 354.250 ;
        RECT 75.380 354.100 79.330 354.250 ;
        RECT 70.130 353.650 70.730 354.100 ;
        RECT 78.730 353.650 79.330 354.100 ;
        RECT 70.130 353.500 74.080 353.650 ;
        RECT 75.380 353.500 79.330 353.650 ;
        RECT 70.130 353.050 70.730 353.500 ;
        RECT 78.730 353.050 79.330 353.500 ;
        RECT 70.130 352.900 74.080 353.050 ;
        RECT 75.380 352.900 79.330 353.050 ;
        RECT 70.130 352.450 70.730 352.900 ;
        RECT 78.730 352.450 79.330 352.900 ;
        RECT 70.130 352.300 74.080 352.450 ;
        RECT 75.380 352.300 79.330 352.450 ;
        RECT 70.130 351.850 70.730 352.300 ;
        RECT 78.730 351.850 79.330 352.300 ;
        RECT 70.130 351.700 74.080 351.850 ;
        RECT 75.380 351.700 79.330 351.850 ;
        RECT 70.130 351.250 70.730 351.700 ;
        RECT 78.730 351.250 79.330 351.700 ;
        RECT 70.130 351.100 74.080 351.250 ;
        RECT 75.380 351.100 79.330 351.250 ;
        RECT 70.130 350.650 70.730 351.100 ;
        RECT 78.730 350.650 79.330 351.100 ;
        RECT 70.130 350.450 74.080 350.650 ;
        RECT 75.380 350.450 79.330 350.650 ;
        RECT 79.780 350.450 79.930 358.000 ;
        RECT 80.380 350.450 80.530 358.000 ;
        RECT 80.980 350.450 81.130 358.000 ;
        RECT 81.580 350.450 81.730 358.000 ;
        RECT 82.180 350.450 82.330 358.000 ;
        RECT 82.780 355.150 82.930 358.000 ;
        RECT 83.530 355.600 85.930 358.800 ;
        RECT 89.280 358.650 90.730 358.950 ;
        RECT 86.530 358.450 90.730 358.650 ;
        RECT 98.730 358.900 104.730 359.800 ;
        RECT 98.730 358.650 100.180 358.900 ;
        RECT 100.330 358.800 104.730 358.900 ;
        RECT 98.730 358.450 102.930 358.650 ;
        RECT 86.530 358.300 94.080 358.450 ;
        RECT 95.430 358.300 102.930 358.450 ;
        RECT 86.530 358.000 90.730 358.300 ;
        RECT 86.530 355.150 86.680 358.000 ;
        RECT 87.130 350.450 87.280 358.000 ;
        RECT 87.730 350.450 87.880 358.000 ;
        RECT 88.330 350.450 88.480 358.000 ;
        RECT 88.930 350.450 89.080 358.000 ;
        RECT 89.530 350.450 89.680 358.000 ;
        RECT 90.130 357.850 90.730 358.000 ;
        RECT 98.730 358.000 102.930 358.300 ;
        RECT 98.730 357.850 99.330 358.000 ;
        RECT 90.130 357.700 94.080 357.850 ;
        RECT 95.380 357.700 99.330 357.850 ;
        RECT 90.130 357.250 90.730 357.700 ;
        RECT 98.730 357.250 99.330 357.700 ;
        RECT 90.130 357.100 94.080 357.250 ;
        RECT 95.380 357.100 99.330 357.250 ;
        RECT 90.130 356.650 90.730 357.100 ;
        RECT 98.730 356.650 99.330 357.100 ;
        RECT 90.130 356.500 94.080 356.650 ;
        RECT 95.380 356.500 99.330 356.650 ;
        RECT 90.130 356.050 90.730 356.500 ;
        RECT 98.730 356.050 99.330 356.500 ;
        RECT 90.130 355.900 94.080 356.050 ;
        RECT 95.380 355.900 99.330 356.050 ;
        RECT 90.130 355.450 90.730 355.900 ;
        RECT 98.730 355.450 99.330 355.900 ;
        RECT 90.130 355.300 94.080 355.450 ;
        RECT 95.380 355.300 99.330 355.450 ;
        RECT 90.130 354.850 90.730 355.300 ;
        RECT 98.730 354.850 99.330 355.300 ;
        RECT 90.130 354.700 94.080 354.850 ;
        RECT 95.380 354.700 99.330 354.850 ;
        RECT 90.130 354.250 90.730 354.700 ;
        RECT 98.730 354.250 99.330 354.700 ;
        RECT 90.130 354.100 94.080 354.250 ;
        RECT 95.380 354.100 99.330 354.250 ;
        RECT 90.130 353.650 90.730 354.100 ;
        RECT 98.730 353.650 99.330 354.100 ;
        RECT 90.130 353.500 94.080 353.650 ;
        RECT 95.380 353.500 99.330 353.650 ;
        RECT 90.130 353.050 90.730 353.500 ;
        RECT 98.730 353.050 99.330 353.500 ;
        RECT 90.130 352.900 94.080 353.050 ;
        RECT 95.380 352.900 99.330 353.050 ;
        RECT 90.130 352.450 90.730 352.900 ;
        RECT 98.730 352.450 99.330 352.900 ;
        RECT 90.130 352.300 94.080 352.450 ;
        RECT 95.380 352.300 99.330 352.450 ;
        RECT 90.130 351.850 90.730 352.300 ;
        RECT 98.730 351.850 99.330 352.300 ;
        RECT 90.130 351.700 94.080 351.850 ;
        RECT 95.380 351.700 99.330 351.850 ;
        RECT 90.130 351.250 90.730 351.700 ;
        RECT 98.730 351.250 99.330 351.700 ;
        RECT 90.130 351.100 94.080 351.250 ;
        RECT 95.380 351.100 99.330 351.250 ;
        RECT 90.130 350.650 90.730 351.100 ;
        RECT 98.730 350.650 99.330 351.100 ;
        RECT 90.130 350.450 94.080 350.650 ;
        RECT 95.380 350.450 99.330 350.650 ;
        RECT 99.780 350.450 99.930 358.000 ;
        RECT 100.380 350.450 100.530 358.000 ;
        RECT 100.980 350.450 101.130 358.000 ;
        RECT 101.580 350.450 101.730 358.000 ;
        RECT 102.180 350.450 102.330 358.000 ;
        RECT 102.780 355.150 102.930 358.000 ;
        RECT 103.530 357.585 104.730 358.800 ;
        RECT 103.530 356.310 107.130 357.585 ;
        RECT 103.530 355.600 104.730 356.310 ;
        RECT 2.315 344.450 4.315 346.745 ;
        RECT 4.730 344.020 5.930 344.400 ;
        RECT 2.315 342.745 5.930 344.020 ;
        RECT 4.730 341.200 5.930 342.745 ;
        RECT 6.530 342.000 6.680 344.900 ;
        RECT 7.130 342.000 7.280 349.550 ;
        RECT 7.730 342.000 7.880 349.550 ;
        RECT 8.330 342.000 8.480 349.550 ;
        RECT 8.930 342.000 9.080 349.550 ;
        RECT 9.530 342.000 9.680 349.550 ;
        RECT 10.130 349.350 14.080 349.550 ;
        RECT 15.380 349.350 19.330 349.550 ;
        RECT 10.130 348.900 10.730 349.350 ;
        RECT 18.730 348.900 19.330 349.350 ;
        RECT 10.130 348.750 14.080 348.900 ;
        RECT 15.380 348.750 19.330 348.900 ;
        RECT 10.130 348.300 10.730 348.750 ;
        RECT 18.730 348.300 19.330 348.750 ;
        RECT 10.130 348.150 14.080 348.300 ;
        RECT 15.380 348.150 19.330 348.300 ;
        RECT 10.130 347.700 10.730 348.150 ;
        RECT 18.730 347.700 19.330 348.150 ;
        RECT 10.130 347.550 14.080 347.700 ;
        RECT 15.380 347.550 19.330 347.700 ;
        RECT 10.130 347.100 10.730 347.550 ;
        RECT 18.730 347.100 19.330 347.550 ;
        RECT 10.130 346.950 14.080 347.100 ;
        RECT 15.380 346.950 19.330 347.100 ;
        RECT 10.130 346.500 10.730 346.950 ;
        RECT 18.730 346.500 19.330 346.950 ;
        RECT 10.130 346.350 14.080 346.500 ;
        RECT 15.380 346.350 19.330 346.500 ;
        RECT 10.130 345.900 10.730 346.350 ;
        RECT 18.730 345.900 19.330 346.350 ;
        RECT 10.130 345.750 14.080 345.900 ;
        RECT 15.380 345.750 19.330 345.900 ;
        RECT 10.130 345.300 10.730 345.750 ;
        RECT 18.730 345.300 19.330 345.750 ;
        RECT 10.130 345.150 14.080 345.300 ;
        RECT 15.380 345.150 19.330 345.300 ;
        RECT 10.130 344.700 10.730 345.150 ;
        RECT 18.730 344.700 19.330 345.150 ;
        RECT 10.130 344.550 14.080 344.700 ;
        RECT 15.380 344.550 19.330 344.700 ;
        RECT 10.130 344.100 10.730 344.550 ;
        RECT 18.730 344.100 19.330 344.550 ;
        RECT 10.130 343.950 14.080 344.100 ;
        RECT 15.380 343.950 19.330 344.100 ;
        RECT 10.130 343.500 10.730 343.950 ;
        RECT 18.730 343.500 19.330 343.950 ;
        RECT 10.130 343.350 14.080 343.500 ;
        RECT 15.380 343.350 19.330 343.500 ;
        RECT 10.130 342.900 10.730 343.350 ;
        RECT 18.730 342.900 19.330 343.350 ;
        RECT 10.130 342.750 14.080 342.900 ;
        RECT 15.380 342.750 19.330 342.900 ;
        RECT 10.130 342.300 10.730 342.750 ;
        RECT 18.730 342.300 19.330 342.750 ;
        RECT 10.130 342.150 14.080 342.300 ;
        RECT 15.380 342.150 19.330 342.300 ;
        RECT 10.130 342.000 10.730 342.150 ;
        RECT 6.530 341.700 10.730 342.000 ;
        RECT 18.730 342.000 19.330 342.150 ;
        RECT 19.780 342.000 19.930 349.550 ;
        RECT 20.380 342.000 20.530 349.550 ;
        RECT 20.980 342.000 21.130 349.550 ;
        RECT 21.580 342.000 21.730 349.550 ;
        RECT 22.180 342.000 22.330 349.550 ;
        RECT 22.780 342.000 22.930 344.900 ;
        RECT 18.730 341.700 22.930 342.000 ;
        RECT 6.530 341.550 14.080 341.700 ;
        RECT 15.380 341.550 22.930 341.700 ;
        RECT 6.530 341.350 10.730 341.550 ;
        RECT 4.730 341.050 9.130 341.200 ;
        RECT 9.280 341.050 10.730 341.350 ;
        RECT 4.730 340.150 10.730 341.050 ;
        RECT 18.730 341.350 22.930 341.550 ;
        RECT 18.730 341.050 20.180 341.350 ;
        RECT 23.530 341.200 25.930 344.400 ;
        RECT 26.530 342.000 26.680 344.900 ;
        RECT 27.130 342.000 27.280 349.550 ;
        RECT 27.730 342.000 27.880 349.550 ;
        RECT 28.330 342.000 28.480 349.550 ;
        RECT 28.930 342.000 29.080 349.550 ;
        RECT 29.530 342.000 29.680 349.550 ;
        RECT 30.130 349.350 34.080 349.550 ;
        RECT 35.380 349.350 39.330 349.550 ;
        RECT 30.130 348.900 30.730 349.350 ;
        RECT 38.730 348.900 39.330 349.350 ;
        RECT 30.130 348.750 34.080 348.900 ;
        RECT 35.380 348.750 39.330 348.900 ;
        RECT 30.130 348.300 30.730 348.750 ;
        RECT 38.730 348.300 39.330 348.750 ;
        RECT 30.130 348.150 34.080 348.300 ;
        RECT 35.380 348.150 39.330 348.300 ;
        RECT 30.130 347.700 30.730 348.150 ;
        RECT 38.730 347.700 39.330 348.150 ;
        RECT 30.130 347.550 34.080 347.700 ;
        RECT 35.380 347.550 39.330 347.700 ;
        RECT 30.130 347.100 30.730 347.550 ;
        RECT 38.730 347.100 39.330 347.550 ;
        RECT 30.130 346.950 34.080 347.100 ;
        RECT 35.380 346.950 39.330 347.100 ;
        RECT 30.130 346.500 30.730 346.950 ;
        RECT 38.730 346.500 39.330 346.950 ;
        RECT 30.130 346.350 34.080 346.500 ;
        RECT 35.380 346.350 39.330 346.500 ;
        RECT 30.130 345.900 30.730 346.350 ;
        RECT 38.730 345.900 39.330 346.350 ;
        RECT 30.130 345.750 34.080 345.900 ;
        RECT 35.380 345.750 39.330 345.900 ;
        RECT 30.130 345.300 30.730 345.750 ;
        RECT 38.730 345.300 39.330 345.750 ;
        RECT 30.130 345.150 34.080 345.300 ;
        RECT 35.380 345.150 39.330 345.300 ;
        RECT 30.130 344.700 30.730 345.150 ;
        RECT 38.730 344.700 39.330 345.150 ;
        RECT 30.130 344.550 34.080 344.700 ;
        RECT 35.380 344.550 39.330 344.700 ;
        RECT 30.130 344.100 30.730 344.550 ;
        RECT 38.730 344.100 39.330 344.550 ;
        RECT 30.130 343.950 34.080 344.100 ;
        RECT 35.380 343.950 39.330 344.100 ;
        RECT 30.130 343.500 30.730 343.950 ;
        RECT 38.730 343.500 39.330 343.950 ;
        RECT 30.130 343.350 34.080 343.500 ;
        RECT 35.380 343.350 39.330 343.500 ;
        RECT 30.130 342.900 30.730 343.350 ;
        RECT 38.730 342.900 39.330 343.350 ;
        RECT 30.130 342.750 34.080 342.900 ;
        RECT 35.380 342.750 39.330 342.900 ;
        RECT 30.130 342.300 30.730 342.750 ;
        RECT 38.730 342.300 39.330 342.750 ;
        RECT 30.130 342.150 34.080 342.300 ;
        RECT 35.380 342.150 39.330 342.300 ;
        RECT 30.130 342.000 30.730 342.150 ;
        RECT 26.530 341.700 30.730 342.000 ;
        RECT 38.730 342.000 39.330 342.150 ;
        RECT 39.780 342.000 39.930 349.550 ;
        RECT 40.380 342.000 40.530 349.550 ;
        RECT 40.980 342.000 41.130 349.550 ;
        RECT 41.580 342.000 41.730 349.550 ;
        RECT 42.180 342.000 42.330 349.550 ;
        RECT 42.780 342.000 42.930 344.900 ;
        RECT 38.730 341.700 42.930 342.000 ;
        RECT 26.530 341.550 34.080 341.700 ;
        RECT 35.380 341.550 42.930 341.700 ;
        RECT 26.530 341.350 30.730 341.550 ;
        RECT 20.330 341.050 29.130 341.200 ;
        RECT 29.280 341.050 30.730 341.350 ;
        RECT 18.730 340.150 30.730 341.050 ;
        RECT 38.730 341.350 42.930 341.550 ;
        RECT 38.730 341.050 40.180 341.350 ;
        RECT 43.530 341.200 45.930 344.400 ;
        RECT 46.530 342.000 46.680 344.900 ;
        RECT 47.130 342.000 47.280 349.550 ;
        RECT 47.730 342.000 47.880 349.550 ;
        RECT 48.330 342.000 48.480 349.550 ;
        RECT 48.930 342.000 49.080 349.550 ;
        RECT 49.530 342.000 49.680 349.550 ;
        RECT 50.130 349.350 54.080 349.550 ;
        RECT 55.380 349.350 59.330 349.550 ;
        RECT 50.130 348.900 50.730 349.350 ;
        RECT 58.730 348.900 59.330 349.350 ;
        RECT 50.130 348.750 54.080 348.900 ;
        RECT 55.380 348.750 59.330 348.900 ;
        RECT 50.130 348.300 50.730 348.750 ;
        RECT 58.730 348.300 59.330 348.750 ;
        RECT 50.130 348.150 54.080 348.300 ;
        RECT 55.380 348.150 59.330 348.300 ;
        RECT 50.130 347.700 50.730 348.150 ;
        RECT 58.730 347.700 59.330 348.150 ;
        RECT 50.130 347.550 54.080 347.700 ;
        RECT 55.380 347.550 59.330 347.700 ;
        RECT 50.130 347.100 50.730 347.550 ;
        RECT 58.730 347.100 59.330 347.550 ;
        RECT 50.130 346.950 54.080 347.100 ;
        RECT 55.380 346.950 59.330 347.100 ;
        RECT 50.130 346.500 50.730 346.950 ;
        RECT 58.730 346.500 59.330 346.950 ;
        RECT 50.130 346.350 54.080 346.500 ;
        RECT 55.380 346.350 59.330 346.500 ;
        RECT 50.130 345.900 50.730 346.350 ;
        RECT 58.730 345.900 59.330 346.350 ;
        RECT 50.130 345.750 54.080 345.900 ;
        RECT 55.380 345.750 59.330 345.900 ;
        RECT 50.130 345.300 50.730 345.750 ;
        RECT 58.730 345.300 59.330 345.750 ;
        RECT 50.130 345.150 54.080 345.300 ;
        RECT 55.380 345.150 59.330 345.300 ;
        RECT 50.130 344.700 50.730 345.150 ;
        RECT 58.730 344.700 59.330 345.150 ;
        RECT 50.130 344.550 54.080 344.700 ;
        RECT 55.380 344.550 59.330 344.700 ;
        RECT 50.130 344.100 50.730 344.550 ;
        RECT 58.730 344.100 59.330 344.550 ;
        RECT 50.130 343.950 54.080 344.100 ;
        RECT 55.380 343.950 59.330 344.100 ;
        RECT 50.130 343.500 50.730 343.950 ;
        RECT 58.730 343.500 59.330 343.950 ;
        RECT 50.130 343.350 54.080 343.500 ;
        RECT 55.380 343.350 59.330 343.500 ;
        RECT 50.130 342.900 50.730 343.350 ;
        RECT 58.730 342.900 59.330 343.350 ;
        RECT 50.130 342.750 54.080 342.900 ;
        RECT 55.380 342.750 59.330 342.900 ;
        RECT 50.130 342.300 50.730 342.750 ;
        RECT 58.730 342.300 59.330 342.750 ;
        RECT 50.130 342.150 54.080 342.300 ;
        RECT 55.380 342.150 59.330 342.300 ;
        RECT 50.130 342.000 50.730 342.150 ;
        RECT 46.530 341.700 50.730 342.000 ;
        RECT 58.730 342.000 59.330 342.150 ;
        RECT 59.780 342.000 59.930 349.550 ;
        RECT 60.380 342.000 60.530 349.550 ;
        RECT 60.980 342.000 61.130 349.550 ;
        RECT 61.580 342.000 61.730 349.550 ;
        RECT 62.180 342.000 62.330 349.550 ;
        RECT 62.780 342.000 62.930 344.900 ;
        RECT 58.730 341.700 62.930 342.000 ;
        RECT 46.530 341.550 54.080 341.700 ;
        RECT 55.380 341.550 62.930 341.700 ;
        RECT 46.530 341.350 50.730 341.550 ;
        RECT 40.330 341.050 49.130 341.200 ;
        RECT 49.280 341.050 50.730 341.350 ;
        RECT 38.730 340.150 50.730 341.050 ;
        RECT 58.730 341.350 62.930 341.550 ;
        RECT 58.730 341.050 60.180 341.350 ;
        RECT 63.530 341.200 65.930 344.400 ;
        RECT 66.530 342.000 66.680 344.900 ;
        RECT 67.130 342.000 67.280 349.550 ;
        RECT 67.730 342.000 67.880 349.550 ;
        RECT 68.330 342.000 68.480 349.550 ;
        RECT 68.930 342.000 69.080 349.550 ;
        RECT 69.530 342.000 69.680 349.550 ;
        RECT 70.130 349.350 74.080 349.550 ;
        RECT 75.380 349.350 79.330 349.550 ;
        RECT 70.130 348.900 70.730 349.350 ;
        RECT 78.730 348.900 79.330 349.350 ;
        RECT 70.130 348.750 74.080 348.900 ;
        RECT 75.380 348.750 79.330 348.900 ;
        RECT 70.130 348.300 70.730 348.750 ;
        RECT 78.730 348.300 79.330 348.750 ;
        RECT 70.130 348.150 74.080 348.300 ;
        RECT 75.380 348.150 79.330 348.300 ;
        RECT 70.130 347.700 70.730 348.150 ;
        RECT 78.730 347.700 79.330 348.150 ;
        RECT 70.130 347.550 74.080 347.700 ;
        RECT 75.380 347.550 79.330 347.700 ;
        RECT 70.130 347.100 70.730 347.550 ;
        RECT 78.730 347.100 79.330 347.550 ;
        RECT 70.130 346.950 74.080 347.100 ;
        RECT 75.380 346.950 79.330 347.100 ;
        RECT 70.130 346.500 70.730 346.950 ;
        RECT 78.730 346.500 79.330 346.950 ;
        RECT 70.130 346.350 74.080 346.500 ;
        RECT 75.380 346.350 79.330 346.500 ;
        RECT 70.130 345.900 70.730 346.350 ;
        RECT 78.730 345.900 79.330 346.350 ;
        RECT 70.130 345.750 74.080 345.900 ;
        RECT 75.380 345.750 79.330 345.900 ;
        RECT 70.130 345.300 70.730 345.750 ;
        RECT 78.730 345.300 79.330 345.750 ;
        RECT 70.130 345.150 74.080 345.300 ;
        RECT 75.380 345.150 79.330 345.300 ;
        RECT 70.130 344.700 70.730 345.150 ;
        RECT 78.730 344.700 79.330 345.150 ;
        RECT 70.130 344.550 74.080 344.700 ;
        RECT 75.380 344.550 79.330 344.700 ;
        RECT 70.130 344.100 70.730 344.550 ;
        RECT 78.730 344.100 79.330 344.550 ;
        RECT 70.130 343.950 74.080 344.100 ;
        RECT 75.380 343.950 79.330 344.100 ;
        RECT 70.130 343.500 70.730 343.950 ;
        RECT 78.730 343.500 79.330 343.950 ;
        RECT 70.130 343.350 74.080 343.500 ;
        RECT 75.380 343.350 79.330 343.500 ;
        RECT 70.130 342.900 70.730 343.350 ;
        RECT 78.730 342.900 79.330 343.350 ;
        RECT 70.130 342.750 74.080 342.900 ;
        RECT 75.380 342.750 79.330 342.900 ;
        RECT 70.130 342.300 70.730 342.750 ;
        RECT 78.730 342.300 79.330 342.750 ;
        RECT 70.130 342.150 74.080 342.300 ;
        RECT 75.380 342.150 79.330 342.300 ;
        RECT 70.130 342.000 70.730 342.150 ;
        RECT 66.530 341.700 70.730 342.000 ;
        RECT 78.730 342.000 79.330 342.150 ;
        RECT 79.780 342.000 79.930 349.550 ;
        RECT 80.380 342.000 80.530 349.550 ;
        RECT 80.980 342.000 81.130 349.550 ;
        RECT 81.580 342.000 81.730 349.550 ;
        RECT 82.180 342.000 82.330 349.550 ;
        RECT 82.780 342.000 82.930 344.900 ;
        RECT 78.730 341.700 82.930 342.000 ;
        RECT 66.530 341.550 74.080 341.700 ;
        RECT 75.380 341.550 82.930 341.700 ;
        RECT 66.530 341.350 70.730 341.550 ;
        RECT 60.330 341.050 69.130 341.200 ;
        RECT 69.280 341.050 70.730 341.350 ;
        RECT 58.730 340.150 70.730 341.050 ;
        RECT 78.730 341.350 82.930 341.550 ;
        RECT 78.730 341.050 80.180 341.350 ;
        RECT 83.530 341.200 85.930 344.400 ;
        RECT 86.530 342.000 86.680 344.900 ;
        RECT 87.130 342.000 87.280 349.550 ;
        RECT 87.730 342.000 87.880 349.550 ;
        RECT 88.330 342.000 88.480 349.550 ;
        RECT 88.930 342.000 89.080 349.550 ;
        RECT 89.530 342.000 89.680 349.550 ;
        RECT 90.130 349.350 94.080 349.550 ;
        RECT 95.380 349.350 99.330 349.550 ;
        RECT 90.130 348.900 90.730 349.350 ;
        RECT 98.730 348.900 99.330 349.350 ;
        RECT 90.130 348.750 94.080 348.900 ;
        RECT 95.380 348.750 99.330 348.900 ;
        RECT 90.130 348.300 90.730 348.750 ;
        RECT 98.730 348.300 99.330 348.750 ;
        RECT 90.130 348.150 94.080 348.300 ;
        RECT 95.380 348.150 99.330 348.300 ;
        RECT 90.130 347.700 90.730 348.150 ;
        RECT 98.730 347.700 99.330 348.150 ;
        RECT 90.130 347.550 94.080 347.700 ;
        RECT 95.380 347.550 99.330 347.700 ;
        RECT 90.130 347.100 90.730 347.550 ;
        RECT 98.730 347.100 99.330 347.550 ;
        RECT 90.130 346.950 94.080 347.100 ;
        RECT 95.380 346.950 99.330 347.100 ;
        RECT 90.130 346.500 90.730 346.950 ;
        RECT 98.730 346.500 99.330 346.950 ;
        RECT 90.130 346.350 94.080 346.500 ;
        RECT 95.380 346.350 99.330 346.500 ;
        RECT 90.130 345.900 90.730 346.350 ;
        RECT 98.730 345.900 99.330 346.350 ;
        RECT 90.130 345.750 94.080 345.900 ;
        RECT 95.380 345.750 99.330 345.900 ;
        RECT 90.130 345.300 90.730 345.750 ;
        RECT 98.730 345.300 99.330 345.750 ;
        RECT 90.130 345.150 94.080 345.300 ;
        RECT 95.380 345.150 99.330 345.300 ;
        RECT 90.130 344.700 90.730 345.150 ;
        RECT 98.730 344.700 99.330 345.150 ;
        RECT 90.130 344.550 94.080 344.700 ;
        RECT 95.380 344.550 99.330 344.700 ;
        RECT 90.130 344.100 90.730 344.550 ;
        RECT 98.730 344.100 99.330 344.550 ;
        RECT 90.130 343.950 94.080 344.100 ;
        RECT 95.380 343.950 99.330 344.100 ;
        RECT 90.130 343.500 90.730 343.950 ;
        RECT 98.730 343.500 99.330 343.950 ;
        RECT 90.130 343.350 94.080 343.500 ;
        RECT 95.380 343.350 99.330 343.500 ;
        RECT 90.130 342.900 90.730 343.350 ;
        RECT 98.730 342.900 99.330 343.350 ;
        RECT 90.130 342.750 94.080 342.900 ;
        RECT 95.380 342.750 99.330 342.900 ;
        RECT 90.130 342.300 90.730 342.750 ;
        RECT 98.730 342.300 99.330 342.750 ;
        RECT 90.130 342.150 94.080 342.300 ;
        RECT 95.380 342.150 99.330 342.300 ;
        RECT 90.130 342.000 90.730 342.150 ;
        RECT 86.530 341.700 90.730 342.000 ;
        RECT 98.730 342.000 99.330 342.150 ;
        RECT 99.780 342.000 99.930 349.550 ;
        RECT 100.380 342.000 100.530 349.550 ;
        RECT 100.980 342.000 101.130 349.550 ;
        RECT 101.580 342.000 101.730 349.550 ;
        RECT 102.180 342.000 102.330 349.550 ;
        RECT 102.780 342.000 102.930 344.900 ;
        RECT 98.730 341.700 102.930 342.000 ;
        RECT 86.530 341.550 94.080 341.700 ;
        RECT 95.380 341.550 102.930 341.700 ;
        RECT 86.530 341.350 90.730 341.550 ;
        RECT 80.330 341.050 89.130 341.200 ;
        RECT 89.280 341.050 90.730 341.350 ;
        RECT 78.730 340.150 90.730 341.050 ;
        RECT 98.730 341.350 102.930 341.550 ;
        RECT 103.530 343.600 104.730 344.400 ;
        RECT 103.530 342.325 107.140 343.600 ;
        RECT 98.730 341.050 100.180 341.350 ;
        RECT 103.530 341.200 104.730 342.325 ;
        RECT 100.330 341.050 104.730 341.200 ;
        RECT 98.730 340.150 104.730 341.050 ;
        RECT 4.730 339.850 9.130 340.150 ;
        RECT 20.330 339.850 29.130 340.150 ;
        RECT 40.330 339.850 49.130 340.150 ;
        RECT 60.330 339.850 69.130 340.150 ;
        RECT 80.330 339.850 89.130 340.150 ;
        RECT 4.730 338.950 10.730 339.850 ;
        RECT 20.330 339.800 30.730 339.850 ;
        RECT 40.330 339.800 50.730 339.850 ;
        RECT 60.330 339.800 70.730 339.850 ;
        RECT 80.330 339.800 90.730 339.850 ;
        RECT 100.330 339.800 104.730 340.150 ;
        RECT 4.730 338.800 9.130 338.950 ;
        RECT 4.730 337.375 5.930 338.800 ;
        RECT 9.280 338.650 10.730 338.950 ;
        RECT 2.315 336.100 5.930 337.375 ;
        RECT 4.730 335.600 5.930 336.100 ;
        RECT 6.530 338.450 10.730 338.650 ;
        RECT 18.730 338.950 30.730 339.800 ;
        RECT 18.730 338.900 29.130 338.950 ;
        RECT 18.730 338.650 20.180 338.900 ;
        RECT 20.330 338.800 29.130 338.900 ;
        RECT 18.730 338.450 22.930 338.650 ;
        RECT 6.530 338.300 14.080 338.450 ;
        RECT 15.430 338.300 22.930 338.450 ;
        RECT 6.530 338.000 10.730 338.300 ;
        RECT 2.315 333.250 4.315 335.545 ;
        RECT 6.530 335.150 6.680 338.000 ;
        RECT 7.130 330.450 7.280 338.000 ;
        RECT 7.730 330.450 7.880 338.000 ;
        RECT 8.330 330.450 8.480 338.000 ;
        RECT 8.930 330.450 9.080 338.000 ;
        RECT 9.530 330.450 9.680 338.000 ;
        RECT 10.130 337.850 10.730 338.000 ;
        RECT 18.730 338.000 22.930 338.300 ;
        RECT 18.730 337.850 19.330 338.000 ;
        RECT 10.130 337.700 14.080 337.850 ;
        RECT 15.380 337.700 19.330 337.850 ;
        RECT 10.130 337.250 10.730 337.700 ;
        RECT 18.730 337.250 19.330 337.700 ;
        RECT 10.130 337.100 14.080 337.250 ;
        RECT 15.380 337.100 19.330 337.250 ;
        RECT 10.130 336.650 10.730 337.100 ;
        RECT 18.730 336.650 19.330 337.100 ;
        RECT 10.130 336.500 14.080 336.650 ;
        RECT 15.380 336.500 19.330 336.650 ;
        RECT 10.130 336.050 10.730 336.500 ;
        RECT 18.730 336.050 19.330 336.500 ;
        RECT 10.130 335.900 14.080 336.050 ;
        RECT 15.380 335.900 19.330 336.050 ;
        RECT 10.130 335.450 10.730 335.900 ;
        RECT 18.730 335.450 19.330 335.900 ;
        RECT 10.130 335.300 14.080 335.450 ;
        RECT 15.380 335.300 19.330 335.450 ;
        RECT 10.130 334.850 10.730 335.300 ;
        RECT 18.730 334.850 19.330 335.300 ;
        RECT 10.130 334.700 14.080 334.850 ;
        RECT 15.380 334.700 19.330 334.850 ;
        RECT 10.130 334.250 10.730 334.700 ;
        RECT 18.730 334.250 19.330 334.700 ;
        RECT 10.130 334.100 14.080 334.250 ;
        RECT 15.380 334.100 19.330 334.250 ;
        RECT 10.130 333.650 10.730 334.100 ;
        RECT 18.730 333.650 19.330 334.100 ;
        RECT 10.130 333.500 14.080 333.650 ;
        RECT 15.380 333.500 19.330 333.650 ;
        RECT 10.130 333.050 10.730 333.500 ;
        RECT 18.730 333.050 19.330 333.500 ;
        RECT 10.130 332.900 14.080 333.050 ;
        RECT 15.380 332.900 19.330 333.050 ;
        RECT 10.130 332.450 10.730 332.900 ;
        RECT 18.730 332.450 19.330 332.900 ;
        RECT 10.130 332.300 14.080 332.450 ;
        RECT 15.380 332.300 19.330 332.450 ;
        RECT 10.130 331.850 10.730 332.300 ;
        RECT 18.730 331.850 19.330 332.300 ;
        RECT 10.130 331.700 14.080 331.850 ;
        RECT 15.380 331.700 19.330 331.850 ;
        RECT 10.130 331.250 10.730 331.700 ;
        RECT 18.730 331.250 19.330 331.700 ;
        RECT 10.130 331.100 14.080 331.250 ;
        RECT 15.380 331.100 19.330 331.250 ;
        RECT 10.130 330.650 10.730 331.100 ;
        RECT 18.730 330.650 19.330 331.100 ;
        RECT 10.130 330.450 14.080 330.650 ;
        RECT 15.380 330.450 19.330 330.650 ;
        RECT 19.780 330.450 19.930 338.000 ;
        RECT 20.380 330.450 20.530 338.000 ;
        RECT 20.980 330.450 21.130 338.000 ;
        RECT 21.580 330.450 21.730 338.000 ;
        RECT 22.180 330.450 22.330 338.000 ;
        RECT 22.780 335.150 22.930 338.000 ;
        RECT 23.530 335.600 25.930 338.800 ;
        RECT 29.280 338.650 30.730 338.950 ;
        RECT 26.530 338.450 30.730 338.650 ;
        RECT 38.730 338.950 50.730 339.800 ;
        RECT 38.730 338.900 49.130 338.950 ;
        RECT 38.730 338.650 40.180 338.900 ;
        RECT 40.330 338.800 49.130 338.900 ;
        RECT 38.730 338.450 42.930 338.650 ;
        RECT 26.530 338.300 34.080 338.450 ;
        RECT 35.430 338.300 42.930 338.450 ;
        RECT 26.530 338.000 30.730 338.300 ;
        RECT 26.530 335.150 26.680 338.000 ;
        RECT 27.130 330.450 27.280 338.000 ;
        RECT 27.730 330.450 27.880 338.000 ;
        RECT 28.330 330.450 28.480 338.000 ;
        RECT 28.930 330.450 29.080 338.000 ;
        RECT 29.530 330.450 29.680 338.000 ;
        RECT 30.130 337.850 30.730 338.000 ;
        RECT 38.730 338.000 42.930 338.300 ;
        RECT 38.730 337.850 39.330 338.000 ;
        RECT 30.130 337.700 34.080 337.850 ;
        RECT 35.380 337.700 39.330 337.850 ;
        RECT 30.130 337.250 30.730 337.700 ;
        RECT 38.730 337.250 39.330 337.700 ;
        RECT 30.130 337.100 34.080 337.250 ;
        RECT 35.380 337.100 39.330 337.250 ;
        RECT 30.130 336.650 30.730 337.100 ;
        RECT 38.730 336.650 39.330 337.100 ;
        RECT 30.130 336.500 34.080 336.650 ;
        RECT 35.380 336.500 39.330 336.650 ;
        RECT 30.130 336.050 30.730 336.500 ;
        RECT 38.730 336.050 39.330 336.500 ;
        RECT 30.130 335.900 34.080 336.050 ;
        RECT 35.380 335.900 39.330 336.050 ;
        RECT 30.130 335.450 30.730 335.900 ;
        RECT 38.730 335.450 39.330 335.900 ;
        RECT 30.130 335.300 34.080 335.450 ;
        RECT 35.380 335.300 39.330 335.450 ;
        RECT 30.130 334.850 30.730 335.300 ;
        RECT 38.730 334.850 39.330 335.300 ;
        RECT 30.130 334.700 34.080 334.850 ;
        RECT 35.380 334.700 39.330 334.850 ;
        RECT 30.130 334.250 30.730 334.700 ;
        RECT 38.730 334.250 39.330 334.700 ;
        RECT 30.130 334.100 34.080 334.250 ;
        RECT 35.380 334.100 39.330 334.250 ;
        RECT 30.130 333.650 30.730 334.100 ;
        RECT 38.730 333.650 39.330 334.100 ;
        RECT 30.130 333.500 34.080 333.650 ;
        RECT 35.380 333.500 39.330 333.650 ;
        RECT 30.130 333.050 30.730 333.500 ;
        RECT 38.730 333.050 39.330 333.500 ;
        RECT 30.130 332.900 34.080 333.050 ;
        RECT 35.380 332.900 39.330 333.050 ;
        RECT 30.130 332.450 30.730 332.900 ;
        RECT 38.730 332.450 39.330 332.900 ;
        RECT 30.130 332.300 34.080 332.450 ;
        RECT 35.380 332.300 39.330 332.450 ;
        RECT 30.130 331.850 30.730 332.300 ;
        RECT 38.730 331.850 39.330 332.300 ;
        RECT 30.130 331.700 34.080 331.850 ;
        RECT 35.380 331.700 39.330 331.850 ;
        RECT 30.130 331.250 30.730 331.700 ;
        RECT 38.730 331.250 39.330 331.700 ;
        RECT 30.130 331.100 34.080 331.250 ;
        RECT 35.380 331.100 39.330 331.250 ;
        RECT 30.130 330.650 30.730 331.100 ;
        RECT 38.730 330.650 39.330 331.100 ;
        RECT 30.130 330.450 34.080 330.650 ;
        RECT 35.380 330.450 39.330 330.650 ;
        RECT 39.780 330.450 39.930 338.000 ;
        RECT 40.380 330.450 40.530 338.000 ;
        RECT 40.980 330.450 41.130 338.000 ;
        RECT 41.580 330.450 41.730 338.000 ;
        RECT 42.180 330.450 42.330 338.000 ;
        RECT 42.780 335.150 42.930 338.000 ;
        RECT 43.530 335.600 45.930 338.800 ;
        RECT 49.280 338.650 50.730 338.950 ;
        RECT 46.530 338.450 50.730 338.650 ;
        RECT 58.730 338.950 70.730 339.800 ;
        RECT 58.730 338.900 69.130 338.950 ;
        RECT 58.730 338.650 60.180 338.900 ;
        RECT 60.330 338.800 69.130 338.900 ;
        RECT 58.730 338.450 62.930 338.650 ;
        RECT 46.530 338.300 54.080 338.450 ;
        RECT 55.430 338.300 62.930 338.450 ;
        RECT 46.530 338.000 50.730 338.300 ;
        RECT 46.530 335.150 46.680 338.000 ;
        RECT 47.130 330.450 47.280 338.000 ;
        RECT 47.730 330.450 47.880 338.000 ;
        RECT 48.330 330.450 48.480 338.000 ;
        RECT 48.930 330.450 49.080 338.000 ;
        RECT 49.530 330.450 49.680 338.000 ;
        RECT 50.130 337.850 50.730 338.000 ;
        RECT 58.730 338.000 62.930 338.300 ;
        RECT 58.730 337.850 59.330 338.000 ;
        RECT 50.130 337.700 54.080 337.850 ;
        RECT 55.380 337.700 59.330 337.850 ;
        RECT 50.130 337.250 50.730 337.700 ;
        RECT 58.730 337.250 59.330 337.700 ;
        RECT 50.130 337.100 54.080 337.250 ;
        RECT 55.380 337.100 59.330 337.250 ;
        RECT 50.130 336.650 50.730 337.100 ;
        RECT 58.730 336.650 59.330 337.100 ;
        RECT 50.130 336.500 54.080 336.650 ;
        RECT 55.380 336.500 59.330 336.650 ;
        RECT 50.130 336.050 50.730 336.500 ;
        RECT 58.730 336.050 59.330 336.500 ;
        RECT 50.130 335.900 54.080 336.050 ;
        RECT 55.380 335.900 59.330 336.050 ;
        RECT 50.130 335.450 50.730 335.900 ;
        RECT 58.730 335.450 59.330 335.900 ;
        RECT 50.130 335.300 54.080 335.450 ;
        RECT 55.380 335.300 59.330 335.450 ;
        RECT 50.130 334.850 50.730 335.300 ;
        RECT 58.730 334.850 59.330 335.300 ;
        RECT 50.130 334.700 54.080 334.850 ;
        RECT 55.380 334.700 59.330 334.850 ;
        RECT 50.130 334.250 50.730 334.700 ;
        RECT 58.730 334.250 59.330 334.700 ;
        RECT 50.130 334.100 54.080 334.250 ;
        RECT 55.380 334.100 59.330 334.250 ;
        RECT 50.130 333.650 50.730 334.100 ;
        RECT 58.730 333.650 59.330 334.100 ;
        RECT 50.130 333.500 54.080 333.650 ;
        RECT 55.380 333.500 59.330 333.650 ;
        RECT 50.130 333.050 50.730 333.500 ;
        RECT 58.730 333.050 59.330 333.500 ;
        RECT 50.130 332.900 54.080 333.050 ;
        RECT 55.380 332.900 59.330 333.050 ;
        RECT 50.130 332.450 50.730 332.900 ;
        RECT 58.730 332.450 59.330 332.900 ;
        RECT 50.130 332.300 54.080 332.450 ;
        RECT 55.380 332.300 59.330 332.450 ;
        RECT 50.130 331.850 50.730 332.300 ;
        RECT 58.730 331.850 59.330 332.300 ;
        RECT 50.130 331.700 54.080 331.850 ;
        RECT 55.380 331.700 59.330 331.850 ;
        RECT 50.130 331.250 50.730 331.700 ;
        RECT 58.730 331.250 59.330 331.700 ;
        RECT 50.130 331.100 54.080 331.250 ;
        RECT 55.380 331.100 59.330 331.250 ;
        RECT 50.130 330.650 50.730 331.100 ;
        RECT 58.730 330.650 59.330 331.100 ;
        RECT 50.130 330.450 54.080 330.650 ;
        RECT 55.380 330.450 59.330 330.650 ;
        RECT 59.780 330.450 59.930 338.000 ;
        RECT 60.380 330.450 60.530 338.000 ;
        RECT 60.980 330.450 61.130 338.000 ;
        RECT 61.580 330.450 61.730 338.000 ;
        RECT 62.180 330.450 62.330 338.000 ;
        RECT 62.780 335.150 62.930 338.000 ;
        RECT 63.530 335.600 65.930 338.800 ;
        RECT 69.280 338.650 70.730 338.950 ;
        RECT 66.530 338.450 70.730 338.650 ;
        RECT 78.730 338.950 90.730 339.800 ;
        RECT 78.730 338.900 89.130 338.950 ;
        RECT 78.730 338.650 80.180 338.900 ;
        RECT 80.330 338.800 89.130 338.900 ;
        RECT 78.730 338.450 82.930 338.650 ;
        RECT 66.530 338.300 74.080 338.450 ;
        RECT 75.430 338.300 82.930 338.450 ;
        RECT 66.530 338.000 70.730 338.300 ;
        RECT 66.530 335.150 66.680 338.000 ;
        RECT 67.130 330.450 67.280 338.000 ;
        RECT 67.730 330.450 67.880 338.000 ;
        RECT 68.330 330.450 68.480 338.000 ;
        RECT 68.930 330.450 69.080 338.000 ;
        RECT 69.530 330.450 69.680 338.000 ;
        RECT 70.130 337.850 70.730 338.000 ;
        RECT 78.730 338.000 82.930 338.300 ;
        RECT 78.730 337.850 79.330 338.000 ;
        RECT 70.130 337.700 74.080 337.850 ;
        RECT 75.380 337.700 79.330 337.850 ;
        RECT 70.130 337.250 70.730 337.700 ;
        RECT 78.730 337.250 79.330 337.700 ;
        RECT 70.130 337.100 74.080 337.250 ;
        RECT 75.380 337.100 79.330 337.250 ;
        RECT 70.130 336.650 70.730 337.100 ;
        RECT 78.730 336.650 79.330 337.100 ;
        RECT 70.130 336.500 74.080 336.650 ;
        RECT 75.380 336.500 79.330 336.650 ;
        RECT 70.130 336.050 70.730 336.500 ;
        RECT 78.730 336.050 79.330 336.500 ;
        RECT 70.130 335.900 74.080 336.050 ;
        RECT 75.380 335.900 79.330 336.050 ;
        RECT 70.130 335.450 70.730 335.900 ;
        RECT 78.730 335.450 79.330 335.900 ;
        RECT 70.130 335.300 74.080 335.450 ;
        RECT 75.380 335.300 79.330 335.450 ;
        RECT 70.130 334.850 70.730 335.300 ;
        RECT 78.730 334.850 79.330 335.300 ;
        RECT 70.130 334.700 74.080 334.850 ;
        RECT 75.380 334.700 79.330 334.850 ;
        RECT 70.130 334.250 70.730 334.700 ;
        RECT 78.730 334.250 79.330 334.700 ;
        RECT 70.130 334.100 74.080 334.250 ;
        RECT 75.380 334.100 79.330 334.250 ;
        RECT 70.130 333.650 70.730 334.100 ;
        RECT 78.730 333.650 79.330 334.100 ;
        RECT 70.130 333.500 74.080 333.650 ;
        RECT 75.380 333.500 79.330 333.650 ;
        RECT 70.130 333.050 70.730 333.500 ;
        RECT 78.730 333.050 79.330 333.500 ;
        RECT 70.130 332.900 74.080 333.050 ;
        RECT 75.380 332.900 79.330 333.050 ;
        RECT 70.130 332.450 70.730 332.900 ;
        RECT 78.730 332.450 79.330 332.900 ;
        RECT 70.130 332.300 74.080 332.450 ;
        RECT 75.380 332.300 79.330 332.450 ;
        RECT 70.130 331.850 70.730 332.300 ;
        RECT 78.730 331.850 79.330 332.300 ;
        RECT 70.130 331.700 74.080 331.850 ;
        RECT 75.380 331.700 79.330 331.850 ;
        RECT 70.130 331.250 70.730 331.700 ;
        RECT 78.730 331.250 79.330 331.700 ;
        RECT 70.130 331.100 74.080 331.250 ;
        RECT 75.380 331.100 79.330 331.250 ;
        RECT 70.130 330.650 70.730 331.100 ;
        RECT 78.730 330.650 79.330 331.100 ;
        RECT 70.130 330.450 74.080 330.650 ;
        RECT 75.380 330.450 79.330 330.650 ;
        RECT 79.780 330.450 79.930 338.000 ;
        RECT 80.380 330.450 80.530 338.000 ;
        RECT 80.980 330.450 81.130 338.000 ;
        RECT 81.580 330.450 81.730 338.000 ;
        RECT 82.180 330.450 82.330 338.000 ;
        RECT 82.780 335.150 82.930 338.000 ;
        RECT 83.530 335.600 85.930 338.800 ;
        RECT 89.280 338.650 90.730 338.950 ;
        RECT 86.530 338.450 90.730 338.650 ;
        RECT 98.730 338.900 104.730 339.800 ;
        RECT 98.730 338.650 100.180 338.900 ;
        RECT 100.330 338.800 104.730 338.900 ;
        RECT 98.730 338.450 102.930 338.650 ;
        RECT 86.530 338.300 94.080 338.450 ;
        RECT 95.430 338.300 102.930 338.450 ;
        RECT 86.530 338.000 90.730 338.300 ;
        RECT 86.530 335.150 86.680 338.000 ;
        RECT 87.130 330.450 87.280 338.000 ;
        RECT 87.730 330.450 87.880 338.000 ;
        RECT 88.330 330.450 88.480 338.000 ;
        RECT 88.930 330.450 89.080 338.000 ;
        RECT 89.530 330.450 89.680 338.000 ;
        RECT 90.130 337.850 90.730 338.000 ;
        RECT 98.730 338.000 102.930 338.300 ;
        RECT 98.730 337.850 99.330 338.000 ;
        RECT 90.130 337.700 94.080 337.850 ;
        RECT 95.380 337.700 99.330 337.850 ;
        RECT 90.130 337.250 90.730 337.700 ;
        RECT 98.730 337.250 99.330 337.700 ;
        RECT 90.130 337.100 94.080 337.250 ;
        RECT 95.380 337.100 99.330 337.250 ;
        RECT 90.130 336.650 90.730 337.100 ;
        RECT 98.730 336.650 99.330 337.100 ;
        RECT 90.130 336.500 94.080 336.650 ;
        RECT 95.380 336.500 99.330 336.650 ;
        RECT 90.130 336.050 90.730 336.500 ;
        RECT 98.730 336.050 99.330 336.500 ;
        RECT 90.130 335.900 94.080 336.050 ;
        RECT 95.380 335.900 99.330 336.050 ;
        RECT 90.130 335.450 90.730 335.900 ;
        RECT 98.730 335.450 99.330 335.900 ;
        RECT 90.130 335.300 94.080 335.450 ;
        RECT 95.380 335.300 99.330 335.450 ;
        RECT 90.130 334.850 90.730 335.300 ;
        RECT 98.730 334.850 99.330 335.300 ;
        RECT 90.130 334.700 94.080 334.850 ;
        RECT 95.380 334.700 99.330 334.850 ;
        RECT 90.130 334.250 90.730 334.700 ;
        RECT 98.730 334.250 99.330 334.700 ;
        RECT 90.130 334.100 94.080 334.250 ;
        RECT 95.380 334.100 99.330 334.250 ;
        RECT 90.130 333.650 90.730 334.100 ;
        RECT 98.730 333.650 99.330 334.100 ;
        RECT 90.130 333.500 94.080 333.650 ;
        RECT 95.380 333.500 99.330 333.650 ;
        RECT 90.130 333.050 90.730 333.500 ;
        RECT 98.730 333.050 99.330 333.500 ;
        RECT 90.130 332.900 94.080 333.050 ;
        RECT 95.380 332.900 99.330 333.050 ;
        RECT 90.130 332.450 90.730 332.900 ;
        RECT 98.730 332.450 99.330 332.900 ;
        RECT 90.130 332.300 94.080 332.450 ;
        RECT 95.380 332.300 99.330 332.450 ;
        RECT 90.130 331.850 90.730 332.300 ;
        RECT 98.730 331.850 99.330 332.300 ;
        RECT 90.130 331.700 94.080 331.850 ;
        RECT 95.380 331.700 99.330 331.850 ;
        RECT 90.130 331.250 90.730 331.700 ;
        RECT 98.730 331.250 99.330 331.700 ;
        RECT 90.130 331.100 94.080 331.250 ;
        RECT 95.380 331.100 99.330 331.250 ;
        RECT 90.130 330.650 90.730 331.100 ;
        RECT 98.730 330.650 99.330 331.100 ;
        RECT 90.130 330.450 94.080 330.650 ;
        RECT 95.380 330.450 99.330 330.650 ;
        RECT 99.780 330.450 99.930 338.000 ;
        RECT 100.380 330.450 100.530 338.000 ;
        RECT 100.980 330.450 101.130 338.000 ;
        RECT 101.580 330.450 101.730 338.000 ;
        RECT 102.180 330.450 102.330 338.000 ;
        RECT 102.780 335.150 102.930 338.000 ;
        RECT 103.530 337.585 104.730 338.800 ;
        RECT 103.530 336.310 107.130 337.585 ;
        RECT 103.530 335.600 104.730 336.310 ;
        RECT 2.315 324.455 4.315 326.750 ;
        RECT 4.730 323.675 5.930 324.400 ;
        RECT 2.315 322.400 5.930 323.675 ;
        RECT 4.730 321.200 5.930 322.400 ;
        RECT 6.530 322.000 6.680 324.900 ;
        RECT 7.130 322.000 7.280 329.550 ;
        RECT 7.730 322.000 7.880 329.550 ;
        RECT 8.330 322.000 8.480 329.550 ;
        RECT 8.930 322.000 9.080 329.550 ;
        RECT 9.530 322.000 9.680 329.550 ;
        RECT 10.130 329.350 14.080 329.550 ;
        RECT 15.380 329.350 19.330 329.550 ;
        RECT 10.130 328.900 10.730 329.350 ;
        RECT 18.730 328.900 19.330 329.350 ;
        RECT 10.130 328.750 14.080 328.900 ;
        RECT 15.380 328.750 19.330 328.900 ;
        RECT 10.130 328.300 10.730 328.750 ;
        RECT 18.730 328.300 19.330 328.750 ;
        RECT 10.130 328.150 14.080 328.300 ;
        RECT 15.380 328.150 19.330 328.300 ;
        RECT 10.130 327.700 10.730 328.150 ;
        RECT 18.730 327.700 19.330 328.150 ;
        RECT 10.130 327.550 14.080 327.700 ;
        RECT 15.380 327.550 19.330 327.700 ;
        RECT 10.130 327.100 10.730 327.550 ;
        RECT 18.730 327.100 19.330 327.550 ;
        RECT 10.130 326.950 14.080 327.100 ;
        RECT 15.380 326.950 19.330 327.100 ;
        RECT 10.130 326.500 10.730 326.950 ;
        RECT 18.730 326.500 19.330 326.950 ;
        RECT 10.130 326.350 14.080 326.500 ;
        RECT 15.380 326.350 19.330 326.500 ;
        RECT 10.130 325.900 10.730 326.350 ;
        RECT 18.730 325.900 19.330 326.350 ;
        RECT 10.130 325.750 14.080 325.900 ;
        RECT 15.380 325.750 19.330 325.900 ;
        RECT 10.130 325.300 10.730 325.750 ;
        RECT 18.730 325.300 19.330 325.750 ;
        RECT 10.130 325.150 14.080 325.300 ;
        RECT 15.380 325.150 19.330 325.300 ;
        RECT 10.130 324.700 10.730 325.150 ;
        RECT 18.730 324.700 19.330 325.150 ;
        RECT 10.130 324.550 14.080 324.700 ;
        RECT 15.380 324.550 19.330 324.700 ;
        RECT 10.130 324.100 10.730 324.550 ;
        RECT 18.730 324.100 19.330 324.550 ;
        RECT 10.130 323.950 14.080 324.100 ;
        RECT 15.380 323.950 19.330 324.100 ;
        RECT 10.130 323.500 10.730 323.950 ;
        RECT 18.730 323.500 19.330 323.950 ;
        RECT 10.130 323.350 14.080 323.500 ;
        RECT 15.380 323.350 19.330 323.500 ;
        RECT 10.130 322.900 10.730 323.350 ;
        RECT 18.730 322.900 19.330 323.350 ;
        RECT 10.130 322.750 14.080 322.900 ;
        RECT 15.380 322.750 19.330 322.900 ;
        RECT 10.130 322.300 10.730 322.750 ;
        RECT 18.730 322.300 19.330 322.750 ;
        RECT 10.130 322.150 14.080 322.300 ;
        RECT 15.380 322.150 19.330 322.300 ;
        RECT 10.130 322.000 10.730 322.150 ;
        RECT 6.530 321.700 10.730 322.000 ;
        RECT 18.730 322.000 19.330 322.150 ;
        RECT 19.780 322.000 19.930 329.550 ;
        RECT 20.380 322.000 20.530 329.550 ;
        RECT 20.980 322.000 21.130 329.550 ;
        RECT 21.580 322.000 21.730 329.550 ;
        RECT 22.180 322.000 22.330 329.550 ;
        RECT 22.780 322.000 22.930 324.900 ;
        RECT 18.730 321.700 22.930 322.000 ;
        RECT 6.530 321.550 14.080 321.700 ;
        RECT 15.380 321.550 22.930 321.700 ;
        RECT 6.530 321.350 10.730 321.550 ;
        RECT 4.730 321.050 9.130 321.200 ;
        RECT 9.280 321.050 10.730 321.350 ;
        RECT 4.730 320.150 10.730 321.050 ;
        RECT 18.730 321.350 22.930 321.550 ;
        RECT 18.730 321.050 20.180 321.350 ;
        RECT 23.530 321.200 25.930 324.400 ;
        RECT 26.530 322.000 26.680 324.900 ;
        RECT 27.130 322.000 27.280 329.550 ;
        RECT 27.730 322.000 27.880 329.550 ;
        RECT 28.330 322.000 28.480 329.550 ;
        RECT 28.930 322.000 29.080 329.550 ;
        RECT 29.530 322.000 29.680 329.550 ;
        RECT 30.130 329.350 34.080 329.550 ;
        RECT 35.380 329.350 39.330 329.550 ;
        RECT 30.130 328.900 30.730 329.350 ;
        RECT 38.730 328.900 39.330 329.350 ;
        RECT 30.130 328.750 34.080 328.900 ;
        RECT 35.380 328.750 39.330 328.900 ;
        RECT 30.130 328.300 30.730 328.750 ;
        RECT 38.730 328.300 39.330 328.750 ;
        RECT 30.130 328.150 34.080 328.300 ;
        RECT 35.380 328.150 39.330 328.300 ;
        RECT 30.130 327.700 30.730 328.150 ;
        RECT 38.730 327.700 39.330 328.150 ;
        RECT 30.130 327.550 34.080 327.700 ;
        RECT 35.380 327.550 39.330 327.700 ;
        RECT 30.130 327.100 30.730 327.550 ;
        RECT 38.730 327.100 39.330 327.550 ;
        RECT 30.130 326.950 34.080 327.100 ;
        RECT 35.380 326.950 39.330 327.100 ;
        RECT 30.130 326.500 30.730 326.950 ;
        RECT 38.730 326.500 39.330 326.950 ;
        RECT 30.130 326.350 34.080 326.500 ;
        RECT 35.380 326.350 39.330 326.500 ;
        RECT 30.130 325.900 30.730 326.350 ;
        RECT 38.730 325.900 39.330 326.350 ;
        RECT 30.130 325.750 34.080 325.900 ;
        RECT 35.380 325.750 39.330 325.900 ;
        RECT 30.130 325.300 30.730 325.750 ;
        RECT 38.730 325.300 39.330 325.750 ;
        RECT 30.130 325.150 34.080 325.300 ;
        RECT 35.380 325.150 39.330 325.300 ;
        RECT 30.130 324.700 30.730 325.150 ;
        RECT 38.730 324.700 39.330 325.150 ;
        RECT 30.130 324.550 34.080 324.700 ;
        RECT 35.380 324.550 39.330 324.700 ;
        RECT 30.130 324.100 30.730 324.550 ;
        RECT 38.730 324.100 39.330 324.550 ;
        RECT 30.130 323.950 34.080 324.100 ;
        RECT 35.380 323.950 39.330 324.100 ;
        RECT 30.130 323.500 30.730 323.950 ;
        RECT 38.730 323.500 39.330 323.950 ;
        RECT 30.130 323.350 34.080 323.500 ;
        RECT 35.380 323.350 39.330 323.500 ;
        RECT 30.130 322.900 30.730 323.350 ;
        RECT 38.730 322.900 39.330 323.350 ;
        RECT 30.130 322.750 34.080 322.900 ;
        RECT 35.380 322.750 39.330 322.900 ;
        RECT 30.130 322.300 30.730 322.750 ;
        RECT 38.730 322.300 39.330 322.750 ;
        RECT 30.130 322.150 34.080 322.300 ;
        RECT 35.380 322.150 39.330 322.300 ;
        RECT 30.130 322.000 30.730 322.150 ;
        RECT 26.530 321.700 30.730 322.000 ;
        RECT 38.730 322.000 39.330 322.150 ;
        RECT 39.780 322.000 39.930 329.550 ;
        RECT 40.380 322.000 40.530 329.550 ;
        RECT 40.980 322.000 41.130 329.550 ;
        RECT 41.580 322.000 41.730 329.550 ;
        RECT 42.180 322.000 42.330 329.550 ;
        RECT 42.780 322.000 42.930 324.900 ;
        RECT 38.730 321.700 42.930 322.000 ;
        RECT 26.530 321.550 34.080 321.700 ;
        RECT 35.380 321.550 42.930 321.700 ;
        RECT 26.530 321.350 30.730 321.550 ;
        RECT 20.330 321.050 29.130 321.200 ;
        RECT 29.280 321.050 30.730 321.350 ;
        RECT 18.730 320.150 30.730 321.050 ;
        RECT 38.730 321.350 42.930 321.550 ;
        RECT 38.730 321.050 40.180 321.350 ;
        RECT 43.530 321.200 45.930 324.400 ;
        RECT 46.530 322.000 46.680 324.900 ;
        RECT 47.130 322.000 47.280 329.550 ;
        RECT 47.730 322.000 47.880 329.550 ;
        RECT 48.330 322.000 48.480 329.550 ;
        RECT 48.930 322.000 49.080 329.550 ;
        RECT 49.530 322.000 49.680 329.550 ;
        RECT 50.130 329.350 54.080 329.550 ;
        RECT 55.380 329.350 59.330 329.550 ;
        RECT 50.130 328.900 50.730 329.350 ;
        RECT 58.730 328.900 59.330 329.350 ;
        RECT 50.130 328.750 54.080 328.900 ;
        RECT 55.380 328.750 59.330 328.900 ;
        RECT 50.130 328.300 50.730 328.750 ;
        RECT 58.730 328.300 59.330 328.750 ;
        RECT 50.130 328.150 54.080 328.300 ;
        RECT 55.380 328.150 59.330 328.300 ;
        RECT 50.130 327.700 50.730 328.150 ;
        RECT 58.730 327.700 59.330 328.150 ;
        RECT 50.130 327.550 54.080 327.700 ;
        RECT 55.380 327.550 59.330 327.700 ;
        RECT 50.130 327.100 50.730 327.550 ;
        RECT 58.730 327.100 59.330 327.550 ;
        RECT 50.130 326.950 54.080 327.100 ;
        RECT 55.380 326.950 59.330 327.100 ;
        RECT 50.130 326.500 50.730 326.950 ;
        RECT 58.730 326.500 59.330 326.950 ;
        RECT 50.130 326.350 54.080 326.500 ;
        RECT 55.380 326.350 59.330 326.500 ;
        RECT 50.130 325.900 50.730 326.350 ;
        RECT 58.730 325.900 59.330 326.350 ;
        RECT 50.130 325.750 54.080 325.900 ;
        RECT 55.380 325.750 59.330 325.900 ;
        RECT 50.130 325.300 50.730 325.750 ;
        RECT 58.730 325.300 59.330 325.750 ;
        RECT 50.130 325.150 54.080 325.300 ;
        RECT 55.380 325.150 59.330 325.300 ;
        RECT 50.130 324.700 50.730 325.150 ;
        RECT 58.730 324.700 59.330 325.150 ;
        RECT 50.130 324.550 54.080 324.700 ;
        RECT 55.380 324.550 59.330 324.700 ;
        RECT 50.130 324.100 50.730 324.550 ;
        RECT 58.730 324.100 59.330 324.550 ;
        RECT 50.130 323.950 54.080 324.100 ;
        RECT 55.380 323.950 59.330 324.100 ;
        RECT 50.130 323.500 50.730 323.950 ;
        RECT 58.730 323.500 59.330 323.950 ;
        RECT 50.130 323.350 54.080 323.500 ;
        RECT 55.380 323.350 59.330 323.500 ;
        RECT 50.130 322.900 50.730 323.350 ;
        RECT 58.730 322.900 59.330 323.350 ;
        RECT 50.130 322.750 54.080 322.900 ;
        RECT 55.380 322.750 59.330 322.900 ;
        RECT 50.130 322.300 50.730 322.750 ;
        RECT 58.730 322.300 59.330 322.750 ;
        RECT 50.130 322.150 54.080 322.300 ;
        RECT 55.380 322.150 59.330 322.300 ;
        RECT 50.130 322.000 50.730 322.150 ;
        RECT 46.530 321.700 50.730 322.000 ;
        RECT 58.730 322.000 59.330 322.150 ;
        RECT 59.780 322.000 59.930 329.550 ;
        RECT 60.380 322.000 60.530 329.550 ;
        RECT 60.980 322.000 61.130 329.550 ;
        RECT 61.580 322.000 61.730 329.550 ;
        RECT 62.180 322.000 62.330 329.550 ;
        RECT 62.780 322.000 62.930 324.900 ;
        RECT 58.730 321.700 62.930 322.000 ;
        RECT 46.530 321.550 54.080 321.700 ;
        RECT 55.380 321.550 62.930 321.700 ;
        RECT 46.530 321.350 50.730 321.550 ;
        RECT 40.330 321.050 49.130 321.200 ;
        RECT 49.280 321.050 50.730 321.350 ;
        RECT 38.730 320.150 50.730 321.050 ;
        RECT 58.730 321.350 62.930 321.550 ;
        RECT 58.730 321.050 60.180 321.350 ;
        RECT 63.530 321.200 65.930 324.400 ;
        RECT 66.530 322.000 66.680 324.900 ;
        RECT 67.130 322.000 67.280 329.550 ;
        RECT 67.730 322.000 67.880 329.550 ;
        RECT 68.330 322.000 68.480 329.550 ;
        RECT 68.930 322.000 69.080 329.550 ;
        RECT 69.530 322.000 69.680 329.550 ;
        RECT 70.130 329.350 74.080 329.550 ;
        RECT 75.380 329.350 79.330 329.550 ;
        RECT 70.130 328.900 70.730 329.350 ;
        RECT 78.730 328.900 79.330 329.350 ;
        RECT 70.130 328.750 74.080 328.900 ;
        RECT 75.380 328.750 79.330 328.900 ;
        RECT 70.130 328.300 70.730 328.750 ;
        RECT 78.730 328.300 79.330 328.750 ;
        RECT 70.130 328.150 74.080 328.300 ;
        RECT 75.380 328.150 79.330 328.300 ;
        RECT 70.130 327.700 70.730 328.150 ;
        RECT 78.730 327.700 79.330 328.150 ;
        RECT 70.130 327.550 74.080 327.700 ;
        RECT 75.380 327.550 79.330 327.700 ;
        RECT 70.130 327.100 70.730 327.550 ;
        RECT 78.730 327.100 79.330 327.550 ;
        RECT 70.130 326.950 74.080 327.100 ;
        RECT 75.380 326.950 79.330 327.100 ;
        RECT 70.130 326.500 70.730 326.950 ;
        RECT 78.730 326.500 79.330 326.950 ;
        RECT 70.130 326.350 74.080 326.500 ;
        RECT 75.380 326.350 79.330 326.500 ;
        RECT 70.130 325.900 70.730 326.350 ;
        RECT 78.730 325.900 79.330 326.350 ;
        RECT 70.130 325.750 74.080 325.900 ;
        RECT 75.380 325.750 79.330 325.900 ;
        RECT 70.130 325.300 70.730 325.750 ;
        RECT 78.730 325.300 79.330 325.750 ;
        RECT 70.130 325.150 74.080 325.300 ;
        RECT 75.380 325.150 79.330 325.300 ;
        RECT 70.130 324.700 70.730 325.150 ;
        RECT 78.730 324.700 79.330 325.150 ;
        RECT 70.130 324.550 74.080 324.700 ;
        RECT 75.380 324.550 79.330 324.700 ;
        RECT 70.130 324.100 70.730 324.550 ;
        RECT 78.730 324.100 79.330 324.550 ;
        RECT 70.130 323.950 74.080 324.100 ;
        RECT 75.380 323.950 79.330 324.100 ;
        RECT 70.130 323.500 70.730 323.950 ;
        RECT 78.730 323.500 79.330 323.950 ;
        RECT 70.130 323.350 74.080 323.500 ;
        RECT 75.380 323.350 79.330 323.500 ;
        RECT 70.130 322.900 70.730 323.350 ;
        RECT 78.730 322.900 79.330 323.350 ;
        RECT 70.130 322.750 74.080 322.900 ;
        RECT 75.380 322.750 79.330 322.900 ;
        RECT 70.130 322.300 70.730 322.750 ;
        RECT 78.730 322.300 79.330 322.750 ;
        RECT 70.130 322.150 74.080 322.300 ;
        RECT 75.380 322.150 79.330 322.300 ;
        RECT 70.130 322.000 70.730 322.150 ;
        RECT 66.530 321.700 70.730 322.000 ;
        RECT 78.730 322.000 79.330 322.150 ;
        RECT 79.780 322.000 79.930 329.550 ;
        RECT 80.380 322.000 80.530 329.550 ;
        RECT 80.980 322.000 81.130 329.550 ;
        RECT 81.580 322.000 81.730 329.550 ;
        RECT 82.180 322.000 82.330 329.550 ;
        RECT 82.780 322.000 82.930 324.900 ;
        RECT 78.730 321.700 82.930 322.000 ;
        RECT 66.530 321.550 74.080 321.700 ;
        RECT 75.380 321.550 82.930 321.700 ;
        RECT 66.530 321.350 70.730 321.550 ;
        RECT 60.330 321.050 69.130 321.200 ;
        RECT 69.280 321.050 70.730 321.350 ;
        RECT 58.730 320.150 70.730 321.050 ;
        RECT 78.730 321.350 82.930 321.550 ;
        RECT 78.730 321.050 80.180 321.350 ;
        RECT 83.530 321.200 85.930 324.400 ;
        RECT 86.530 322.000 86.680 324.900 ;
        RECT 87.130 322.000 87.280 329.550 ;
        RECT 87.730 322.000 87.880 329.550 ;
        RECT 88.330 322.000 88.480 329.550 ;
        RECT 88.930 322.000 89.080 329.550 ;
        RECT 89.530 322.000 89.680 329.550 ;
        RECT 90.130 329.350 94.080 329.550 ;
        RECT 95.380 329.350 99.330 329.550 ;
        RECT 90.130 328.900 90.730 329.350 ;
        RECT 98.730 328.900 99.330 329.350 ;
        RECT 90.130 328.750 94.080 328.900 ;
        RECT 95.380 328.750 99.330 328.900 ;
        RECT 90.130 328.300 90.730 328.750 ;
        RECT 98.730 328.300 99.330 328.750 ;
        RECT 90.130 328.150 94.080 328.300 ;
        RECT 95.380 328.150 99.330 328.300 ;
        RECT 90.130 327.700 90.730 328.150 ;
        RECT 98.730 327.700 99.330 328.150 ;
        RECT 90.130 327.550 94.080 327.700 ;
        RECT 95.380 327.550 99.330 327.700 ;
        RECT 90.130 327.100 90.730 327.550 ;
        RECT 98.730 327.100 99.330 327.550 ;
        RECT 90.130 326.950 94.080 327.100 ;
        RECT 95.380 326.950 99.330 327.100 ;
        RECT 90.130 326.500 90.730 326.950 ;
        RECT 98.730 326.500 99.330 326.950 ;
        RECT 90.130 326.350 94.080 326.500 ;
        RECT 95.380 326.350 99.330 326.500 ;
        RECT 90.130 325.900 90.730 326.350 ;
        RECT 98.730 325.900 99.330 326.350 ;
        RECT 90.130 325.750 94.080 325.900 ;
        RECT 95.380 325.750 99.330 325.900 ;
        RECT 90.130 325.300 90.730 325.750 ;
        RECT 98.730 325.300 99.330 325.750 ;
        RECT 90.130 325.150 94.080 325.300 ;
        RECT 95.380 325.150 99.330 325.300 ;
        RECT 90.130 324.700 90.730 325.150 ;
        RECT 98.730 324.700 99.330 325.150 ;
        RECT 90.130 324.550 94.080 324.700 ;
        RECT 95.380 324.550 99.330 324.700 ;
        RECT 90.130 324.100 90.730 324.550 ;
        RECT 98.730 324.100 99.330 324.550 ;
        RECT 90.130 323.950 94.080 324.100 ;
        RECT 95.380 323.950 99.330 324.100 ;
        RECT 90.130 323.500 90.730 323.950 ;
        RECT 98.730 323.500 99.330 323.950 ;
        RECT 90.130 323.350 94.080 323.500 ;
        RECT 95.380 323.350 99.330 323.500 ;
        RECT 90.130 322.900 90.730 323.350 ;
        RECT 98.730 322.900 99.330 323.350 ;
        RECT 90.130 322.750 94.080 322.900 ;
        RECT 95.380 322.750 99.330 322.900 ;
        RECT 90.130 322.300 90.730 322.750 ;
        RECT 98.730 322.300 99.330 322.750 ;
        RECT 90.130 322.150 94.080 322.300 ;
        RECT 95.380 322.150 99.330 322.300 ;
        RECT 90.130 322.000 90.730 322.150 ;
        RECT 86.530 321.700 90.730 322.000 ;
        RECT 98.730 322.000 99.330 322.150 ;
        RECT 99.780 322.000 99.930 329.550 ;
        RECT 100.380 322.000 100.530 329.550 ;
        RECT 100.980 322.000 101.130 329.550 ;
        RECT 101.580 322.000 101.730 329.550 ;
        RECT 102.180 322.000 102.330 329.550 ;
        RECT 102.780 322.000 102.930 324.900 ;
        RECT 98.730 321.700 102.930 322.000 ;
        RECT 86.530 321.550 94.080 321.700 ;
        RECT 95.380 321.550 102.930 321.700 ;
        RECT 86.530 321.350 90.730 321.550 ;
        RECT 80.330 321.050 89.130 321.200 ;
        RECT 89.280 321.050 90.730 321.350 ;
        RECT 78.730 320.150 90.730 321.050 ;
        RECT 98.730 321.350 102.930 321.550 ;
        RECT 103.530 323.600 104.730 324.400 ;
        RECT 103.530 322.325 107.140 323.600 ;
        RECT 98.730 321.050 100.180 321.350 ;
        RECT 103.530 321.200 104.730 322.325 ;
        RECT 100.330 321.050 104.730 321.200 ;
        RECT 98.730 320.150 104.730 321.050 ;
        RECT 4.730 319.850 9.130 320.150 ;
        RECT 20.330 319.850 29.130 320.150 ;
        RECT 40.330 319.850 49.130 320.150 ;
        RECT 60.330 319.850 69.130 320.150 ;
        RECT 80.330 319.850 89.130 320.150 ;
        RECT 4.730 318.950 10.730 319.850 ;
        RECT 20.330 319.800 30.730 319.850 ;
        RECT 40.330 319.800 50.730 319.850 ;
        RECT 60.330 319.800 70.730 319.850 ;
        RECT 80.330 319.800 90.730 319.850 ;
        RECT 100.330 319.800 104.730 320.150 ;
        RECT 4.730 318.800 9.130 318.950 ;
        RECT 4.730 317.785 5.930 318.800 ;
        RECT 9.280 318.650 10.730 318.950 ;
        RECT 2.315 316.510 5.930 317.785 ;
        RECT 4.730 315.600 5.930 316.510 ;
        RECT 6.530 318.450 10.730 318.650 ;
        RECT 18.730 318.950 30.730 319.800 ;
        RECT 18.730 318.900 29.130 318.950 ;
        RECT 18.730 318.650 20.180 318.900 ;
        RECT 20.330 318.800 29.130 318.900 ;
        RECT 18.730 318.450 22.930 318.650 ;
        RECT 6.530 318.300 14.080 318.450 ;
        RECT 15.430 318.300 22.930 318.450 ;
        RECT 6.530 318.000 10.730 318.300 ;
        RECT 2.320 315.340 4.320 315.545 ;
        RECT 2.315 313.250 4.320 315.340 ;
        RECT 6.530 315.150 6.680 318.000 ;
        RECT 7.130 310.450 7.280 318.000 ;
        RECT 7.730 310.450 7.880 318.000 ;
        RECT 8.330 310.450 8.480 318.000 ;
        RECT 8.930 310.450 9.080 318.000 ;
        RECT 9.530 310.450 9.680 318.000 ;
        RECT 10.130 317.850 10.730 318.000 ;
        RECT 18.730 318.000 22.930 318.300 ;
        RECT 18.730 317.850 19.330 318.000 ;
        RECT 10.130 317.700 14.080 317.850 ;
        RECT 15.380 317.700 19.330 317.850 ;
        RECT 10.130 317.250 10.730 317.700 ;
        RECT 18.730 317.250 19.330 317.700 ;
        RECT 10.130 317.100 14.080 317.250 ;
        RECT 15.380 317.100 19.330 317.250 ;
        RECT 10.130 316.650 10.730 317.100 ;
        RECT 18.730 316.650 19.330 317.100 ;
        RECT 10.130 316.500 14.080 316.650 ;
        RECT 15.380 316.500 19.330 316.650 ;
        RECT 10.130 316.050 10.730 316.500 ;
        RECT 18.730 316.050 19.330 316.500 ;
        RECT 10.130 315.900 14.080 316.050 ;
        RECT 15.380 315.900 19.330 316.050 ;
        RECT 10.130 315.450 10.730 315.900 ;
        RECT 18.730 315.450 19.330 315.900 ;
        RECT 10.130 315.300 14.080 315.450 ;
        RECT 15.380 315.300 19.330 315.450 ;
        RECT 10.130 314.850 10.730 315.300 ;
        RECT 18.730 314.850 19.330 315.300 ;
        RECT 10.130 314.700 14.080 314.850 ;
        RECT 15.380 314.700 19.330 314.850 ;
        RECT 10.130 314.250 10.730 314.700 ;
        RECT 18.730 314.250 19.330 314.700 ;
        RECT 10.130 314.100 14.080 314.250 ;
        RECT 15.380 314.100 19.330 314.250 ;
        RECT 10.130 313.650 10.730 314.100 ;
        RECT 18.730 313.650 19.330 314.100 ;
        RECT 10.130 313.500 14.080 313.650 ;
        RECT 15.380 313.500 19.330 313.650 ;
        RECT 10.130 313.050 10.730 313.500 ;
        RECT 18.730 313.050 19.330 313.500 ;
        RECT 10.130 312.900 14.080 313.050 ;
        RECT 15.380 312.900 19.330 313.050 ;
        RECT 10.130 312.450 10.730 312.900 ;
        RECT 18.730 312.450 19.330 312.900 ;
        RECT 10.130 312.300 14.080 312.450 ;
        RECT 15.380 312.300 19.330 312.450 ;
        RECT 10.130 311.850 10.730 312.300 ;
        RECT 18.730 311.850 19.330 312.300 ;
        RECT 10.130 311.700 14.080 311.850 ;
        RECT 15.380 311.700 19.330 311.850 ;
        RECT 10.130 311.250 10.730 311.700 ;
        RECT 18.730 311.250 19.330 311.700 ;
        RECT 10.130 311.100 14.080 311.250 ;
        RECT 15.380 311.100 19.330 311.250 ;
        RECT 10.130 310.650 10.730 311.100 ;
        RECT 18.730 310.650 19.330 311.100 ;
        RECT 10.130 310.450 14.080 310.650 ;
        RECT 15.380 310.450 19.330 310.650 ;
        RECT 19.780 310.450 19.930 318.000 ;
        RECT 20.380 310.450 20.530 318.000 ;
        RECT 20.980 310.450 21.130 318.000 ;
        RECT 21.580 310.450 21.730 318.000 ;
        RECT 22.180 310.450 22.330 318.000 ;
        RECT 22.780 315.150 22.930 318.000 ;
        RECT 23.530 315.600 25.930 318.800 ;
        RECT 29.280 318.650 30.730 318.950 ;
        RECT 26.530 318.450 30.730 318.650 ;
        RECT 38.730 318.950 50.730 319.800 ;
        RECT 38.730 318.900 49.130 318.950 ;
        RECT 38.730 318.650 40.180 318.900 ;
        RECT 40.330 318.800 49.130 318.900 ;
        RECT 38.730 318.450 42.930 318.650 ;
        RECT 26.530 318.300 34.080 318.450 ;
        RECT 35.430 318.300 42.930 318.450 ;
        RECT 26.530 318.000 30.730 318.300 ;
        RECT 26.530 315.150 26.680 318.000 ;
        RECT 27.130 310.450 27.280 318.000 ;
        RECT 27.730 310.450 27.880 318.000 ;
        RECT 28.330 310.450 28.480 318.000 ;
        RECT 28.930 310.450 29.080 318.000 ;
        RECT 29.530 310.450 29.680 318.000 ;
        RECT 30.130 317.850 30.730 318.000 ;
        RECT 38.730 318.000 42.930 318.300 ;
        RECT 38.730 317.850 39.330 318.000 ;
        RECT 30.130 317.700 34.080 317.850 ;
        RECT 35.380 317.700 39.330 317.850 ;
        RECT 30.130 317.250 30.730 317.700 ;
        RECT 38.730 317.250 39.330 317.700 ;
        RECT 30.130 317.100 34.080 317.250 ;
        RECT 35.380 317.100 39.330 317.250 ;
        RECT 30.130 316.650 30.730 317.100 ;
        RECT 38.730 316.650 39.330 317.100 ;
        RECT 30.130 316.500 34.080 316.650 ;
        RECT 35.380 316.500 39.330 316.650 ;
        RECT 30.130 316.050 30.730 316.500 ;
        RECT 38.730 316.050 39.330 316.500 ;
        RECT 30.130 315.900 34.080 316.050 ;
        RECT 35.380 315.900 39.330 316.050 ;
        RECT 30.130 315.450 30.730 315.900 ;
        RECT 38.730 315.450 39.330 315.900 ;
        RECT 30.130 315.300 34.080 315.450 ;
        RECT 35.380 315.300 39.330 315.450 ;
        RECT 30.130 314.850 30.730 315.300 ;
        RECT 38.730 314.850 39.330 315.300 ;
        RECT 30.130 314.700 34.080 314.850 ;
        RECT 35.380 314.700 39.330 314.850 ;
        RECT 30.130 314.250 30.730 314.700 ;
        RECT 38.730 314.250 39.330 314.700 ;
        RECT 30.130 314.100 34.080 314.250 ;
        RECT 35.380 314.100 39.330 314.250 ;
        RECT 30.130 313.650 30.730 314.100 ;
        RECT 38.730 313.650 39.330 314.100 ;
        RECT 30.130 313.500 34.080 313.650 ;
        RECT 35.380 313.500 39.330 313.650 ;
        RECT 30.130 313.050 30.730 313.500 ;
        RECT 38.730 313.050 39.330 313.500 ;
        RECT 30.130 312.900 34.080 313.050 ;
        RECT 35.380 312.900 39.330 313.050 ;
        RECT 30.130 312.450 30.730 312.900 ;
        RECT 38.730 312.450 39.330 312.900 ;
        RECT 30.130 312.300 34.080 312.450 ;
        RECT 35.380 312.300 39.330 312.450 ;
        RECT 30.130 311.850 30.730 312.300 ;
        RECT 38.730 311.850 39.330 312.300 ;
        RECT 30.130 311.700 34.080 311.850 ;
        RECT 35.380 311.700 39.330 311.850 ;
        RECT 30.130 311.250 30.730 311.700 ;
        RECT 38.730 311.250 39.330 311.700 ;
        RECT 30.130 311.100 34.080 311.250 ;
        RECT 35.380 311.100 39.330 311.250 ;
        RECT 30.130 310.650 30.730 311.100 ;
        RECT 38.730 310.650 39.330 311.100 ;
        RECT 30.130 310.450 34.080 310.650 ;
        RECT 35.380 310.450 39.330 310.650 ;
        RECT 39.780 310.450 39.930 318.000 ;
        RECT 40.380 310.450 40.530 318.000 ;
        RECT 40.980 310.450 41.130 318.000 ;
        RECT 41.580 310.450 41.730 318.000 ;
        RECT 42.180 310.450 42.330 318.000 ;
        RECT 42.780 315.150 42.930 318.000 ;
        RECT 43.530 315.600 45.930 318.800 ;
        RECT 49.280 318.650 50.730 318.950 ;
        RECT 46.530 318.450 50.730 318.650 ;
        RECT 58.730 318.950 70.730 319.800 ;
        RECT 58.730 318.900 69.130 318.950 ;
        RECT 58.730 318.650 60.180 318.900 ;
        RECT 60.330 318.800 69.130 318.900 ;
        RECT 58.730 318.450 62.930 318.650 ;
        RECT 46.530 318.300 54.080 318.450 ;
        RECT 55.430 318.300 62.930 318.450 ;
        RECT 46.530 318.000 50.730 318.300 ;
        RECT 46.530 315.150 46.680 318.000 ;
        RECT 47.130 310.450 47.280 318.000 ;
        RECT 47.730 310.450 47.880 318.000 ;
        RECT 48.330 310.450 48.480 318.000 ;
        RECT 48.930 310.450 49.080 318.000 ;
        RECT 49.530 310.450 49.680 318.000 ;
        RECT 50.130 317.850 50.730 318.000 ;
        RECT 58.730 318.000 62.930 318.300 ;
        RECT 58.730 317.850 59.330 318.000 ;
        RECT 50.130 317.700 54.080 317.850 ;
        RECT 55.380 317.700 59.330 317.850 ;
        RECT 50.130 317.250 50.730 317.700 ;
        RECT 58.730 317.250 59.330 317.700 ;
        RECT 50.130 317.100 54.080 317.250 ;
        RECT 55.380 317.100 59.330 317.250 ;
        RECT 50.130 316.650 50.730 317.100 ;
        RECT 58.730 316.650 59.330 317.100 ;
        RECT 50.130 316.500 54.080 316.650 ;
        RECT 55.380 316.500 59.330 316.650 ;
        RECT 50.130 316.050 50.730 316.500 ;
        RECT 58.730 316.050 59.330 316.500 ;
        RECT 50.130 315.900 54.080 316.050 ;
        RECT 55.380 315.900 59.330 316.050 ;
        RECT 50.130 315.450 50.730 315.900 ;
        RECT 58.730 315.450 59.330 315.900 ;
        RECT 50.130 315.300 54.080 315.450 ;
        RECT 55.380 315.300 59.330 315.450 ;
        RECT 50.130 314.850 50.730 315.300 ;
        RECT 58.730 314.850 59.330 315.300 ;
        RECT 50.130 314.700 54.080 314.850 ;
        RECT 55.380 314.700 59.330 314.850 ;
        RECT 50.130 314.250 50.730 314.700 ;
        RECT 58.730 314.250 59.330 314.700 ;
        RECT 50.130 314.100 54.080 314.250 ;
        RECT 55.380 314.100 59.330 314.250 ;
        RECT 50.130 313.650 50.730 314.100 ;
        RECT 58.730 313.650 59.330 314.100 ;
        RECT 50.130 313.500 54.080 313.650 ;
        RECT 55.380 313.500 59.330 313.650 ;
        RECT 50.130 313.050 50.730 313.500 ;
        RECT 58.730 313.050 59.330 313.500 ;
        RECT 50.130 312.900 54.080 313.050 ;
        RECT 55.380 312.900 59.330 313.050 ;
        RECT 50.130 312.450 50.730 312.900 ;
        RECT 58.730 312.450 59.330 312.900 ;
        RECT 50.130 312.300 54.080 312.450 ;
        RECT 55.380 312.300 59.330 312.450 ;
        RECT 50.130 311.850 50.730 312.300 ;
        RECT 58.730 311.850 59.330 312.300 ;
        RECT 50.130 311.700 54.080 311.850 ;
        RECT 55.380 311.700 59.330 311.850 ;
        RECT 50.130 311.250 50.730 311.700 ;
        RECT 58.730 311.250 59.330 311.700 ;
        RECT 50.130 311.100 54.080 311.250 ;
        RECT 55.380 311.100 59.330 311.250 ;
        RECT 50.130 310.650 50.730 311.100 ;
        RECT 58.730 310.650 59.330 311.100 ;
        RECT 50.130 310.450 54.080 310.650 ;
        RECT 55.380 310.450 59.330 310.650 ;
        RECT 59.780 310.450 59.930 318.000 ;
        RECT 60.380 310.450 60.530 318.000 ;
        RECT 60.980 310.450 61.130 318.000 ;
        RECT 61.580 310.450 61.730 318.000 ;
        RECT 62.180 310.450 62.330 318.000 ;
        RECT 62.780 315.150 62.930 318.000 ;
        RECT 63.530 315.600 65.930 318.800 ;
        RECT 69.280 318.650 70.730 318.950 ;
        RECT 66.530 318.450 70.730 318.650 ;
        RECT 78.730 318.950 90.730 319.800 ;
        RECT 78.730 318.900 89.130 318.950 ;
        RECT 78.730 318.650 80.180 318.900 ;
        RECT 80.330 318.800 89.130 318.900 ;
        RECT 78.730 318.450 82.930 318.650 ;
        RECT 66.530 318.300 74.080 318.450 ;
        RECT 75.430 318.300 82.930 318.450 ;
        RECT 66.530 318.000 70.730 318.300 ;
        RECT 66.530 315.150 66.680 318.000 ;
        RECT 67.130 310.450 67.280 318.000 ;
        RECT 67.730 310.450 67.880 318.000 ;
        RECT 68.330 310.450 68.480 318.000 ;
        RECT 68.930 310.450 69.080 318.000 ;
        RECT 69.530 310.450 69.680 318.000 ;
        RECT 70.130 317.850 70.730 318.000 ;
        RECT 78.730 318.000 82.930 318.300 ;
        RECT 78.730 317.850 79.330 318.000 ;
        RECT 70.130 317.700 74.080 317.850 ;
        RECT 75.380 317.700 79.330 317.850 ;
        RECT 70.130 317.250 70.730 317.700 ;
        RECT 78.730 317.250 79.330 317.700 ;
        RECT 70.130 317.100 74.080 317.250 ;
        RECT 75.380 317.100 79.330 317.250 ;
        RECT 70.130 316.650 70.730 317.100 ;
        RECT 78.730 316.650 79.330 317.100 ;
        RECT 70.130 316.500 74.080 316.650 ;
        RECT 75.380 316.500 79.330 316.650 ;
        RECT 70.130 316.050 70.730 316.500 ;
        RECT 78.730 316.050 79.330 316.500 ;
        RECT 70.130 315.900 74.080 316.050 ;
        RECT 75.380 315.900 79.330 316.050 ;
        RECT 70.130 315.450 70.730 315.900 ;
        RECT 78.730 315.450 79.330 315.900 ;
        RECT 70.130 315.300 74.080 315.450 ;
        RECT 75.380 315.300 79.330 315.450 ;
        RECT 70.130 314.850 70.730 315.300 ;
        RECT 78.730 314.850 79.330 315.300 ;
        RECT 70.130 314.700 74.080 314.850 ;
        RECT 75.380 314.700 79.330 314.850 ;
        RECT 70.130 314.250 70.730 314.700 ;
        RECT 78.730 314.250 79.330 314.700 ;
        RECT 70.130 314.100 74.080 314.250 ;
        RECT 75.380 314.100 79.330 314.250 ;
        RECT 70.130 313.650 70.730 314.100 ;
        RECT 78.730 313.650 79.330 314.100 ;
        RECT 70.130 313.500 74.080 313.650 ;
        RECT 75.380 313.500 79.330 313.650 ;
        RECT 70.130 313.050 70.730 313.500 ;
        RECT 78.730 313.050 79.330 313.500 ;
        RECT 70.130 312.900 74.080 313.050 ;
        RECT 75.380 312.900 79.330 313.050 ;
        RECT 70.130 312.450 70.730 312.900 ;
        RECT 78.730 312.450 79.330 312.900 ;
        RECT 70.130 312.300 74.080 312.450 ;
        RECT 75.380 312.300 79.330 312.450 ;
        RECT 70.130 311.850 70.730 312.300 ;
        RECT 78.730 311.850 79.330 312.300 ;
        RECT 70.130 311.700 74.080 311.850 ;
        RECT 75.380 311.700 79.330 311.850 ;
        RECT 70.130 311.250 70.730 311.700 ;
        RECT 78.730 311.250 79.330 311.700 ;
        RECT 70.130 311.100 74.080 311.250 ;
        RECT 75.380 311.100 79.330 311.250 ;
        RECT 70.130 310.650 70.730 311.100 ;
        RECT 78.730 310.650 79.330 311.100 ;
        RECT 70.130 310.450 74.080 310.650 ;
        RECT 75.380 310.450 79.330 310.650 ;
        RECT 79.780 310.450 79.930 318.000 ;
        RECT 80.380 310.450 80.530 318.000 ;
        RECT 80.980 310.450 81.130 318.000 ;
        RECT 81.580 310.450 81.730 318.000 ;
        RECT 82.180 310.450 82.330 318.000 ;
        RECT 82.780 315.150 82.930 318.000 ;
        RECT 83.530 315.600 85.930 318.800 ;
        RECT 89.280 318.650 90.730 318.950 ;
        RECT 86.530 318.450 90.730 318.650 ;
        RECT 98.730 318.900 104.730 319.800 ;
        RECT 98.730 318.650 100.180 318.900 ;
        RECT 100.330 318.800 104.730 318.900 ;
        RECT 98.730 318.450 102.930 318.650 ;
        RECT 86.530 318.300 94.080 318.450 ;
        RECT 95.430 318.300 102.930 318.450 ;
        RECT 86.530 318.000 90.730 318.300 ;
        RECT 86.530 315.150 86.680 318.000 ;
        RECT 87.130 310.450 87.280 318.000 ;
        RECT 87.730 310.450 87.880 318.000 ;
        RECT 88.330 310.450 88.480 318.000 ;
        RECT 88.930 310.450 89.080 318.000 ;
        RECT 89.530 310.450 89.680 318.000 ;
        RECT 90.130 317.850 90.730 318.000 ;
        RECT 98.730 318.000 102.930 318.300 ;
        RECT 98.730 317.850 99.330 318.000 ;
        RECT 90.130 317.700 94.080 317.850 ;
        RECT 95.380 317.700 99.330 317.850 ;
        RECT 90.130 317.250 90.730 317.700 ;
        RECT 98.730 317.250 99.330 317.700 ;
        RECT 90.130 317.100 94.080 317.250 ;
        RECT 95.380 317.100 99.330 317.250 ;
        RECT 90.130 316.650 90.730 317.100 ;
        RECT 98.730 316.650 99.330 317.100 ;
        RECT 90.130 316.500 94.080 316.650 ;
        RECT 95.380 316.500 99.330 316.650 ;
        RECT 90.130 316.050 90.730 316.500 ;
        RECT 98.730 316.050 99.330 316.500 ;
        RECT 90.130 315.900 94.080 316.050 ;
        RECT 95.380 315.900 99.330 316.050 ;
        RECT 90.130 315.450 90.730 315.900 ;
        RECT 98.730 315.450 99.330 315.900 ;
        RECT 90.130 315.300 94.080 315.450 ;
        RECT 95.380 315.300 99.330 315.450 ;
        RECT 90.130 314.850 90.730 315.300 ;
        RECT 98.730 314.850 99.330 315.300 ;
        RECT 90.130 314.700 94.080 314.850 ;
        RECT 95.380 314.700 99.330 314.850 ;
        RECT 90.130 314.250 90.730 314.700 ;
        RECT 98.730 314.250 99.330 314.700 ;
        RECT 90.130 314.100 94.080 314.250 ;
        RECT 95.380 314.100 99.330 314.250 ;
        RECT 90.130 313.650 90.730 314.100 ;
        RECT 98.730 313.650 99.330 314.100 ;
        RECT 90.130 313.500 94.080 313.650 ;
        RECT 95.380 313.500 99.330 313.650 ;
        RECT 90.130 313.050 90.730 313.500 ;
        RECT 98.730 313.050 99.330 313.500 ;
        RECT 90.130 312.900 94.080 313.050 ;
        RECT 95.380 312.900 99.330 313.050 ;
        RECT 90.130 312.450 90.730 312.900 ;
        RECT 98.730 312.450 99.330 312.900 ;
        RECT 90.130 312.300 94.080 312.450 ;
        RECT 95.380 312.300 99.330 312.450 ;
        RECT 90.130 311.850 90.730 312.300 ;
        RECT 98.730 311.850 99.330 312.300 ;
        RECT 90.130 311.700 94.080 311.850 ;
        RECT 95.380 311.700 99.330 311.850 ;
        RECT 90.130 311.250 90.730 311.700 ;
        RECT 98.730 311.250 99.330 311.700 ;
        RECT 90.130 311.100 94.080 311.250 ;
        RECT 95.380 311.100 99.330 311.250 ;
        RECT 90.130 310.650 90.730 311.100 ;
        RECT 98.730 310.650 99.330 311.100 ;
        RECT 90.130 310.450 94.080 310.650 ;
        RECT 95.380 310.450 99.330 310.650 ;
        RECT 99.780 310.450 99.930 318.000 ;
        RECT 100.380 310.450 100.530 318.000 ;
        RECT 100.980 310.450 101.130 318.000 ;
        RECT 101.580 310.450 101.730 318.000 ;
        RECT 102.180 310.450 102.330 318.000 ;
        RECT 102.780 315.150 102.930 318.000 ;
        RECT 103.530 317.585 104.730 318.800 ;
        RECT 103.530 316.310 107.130 317.585 ;
        RECT 103.530 315.600 104.730 316.310 ;
        RECT 2.315 304.455 4.315 306.750 ;
        RECT 4.730 303.545 5.930 304.400 ;
        RECT 2.315 302.270 5.930 303.545 ;
        RECT 4.730 301.200 5.930 302.270 ;
        RECT 6.530 302.000 6.680 304.900 ;
        RECT 7.130 302.000 7.280 309.550 ;
        RECT 7.730 302.000 7.880 309.550 ;
        RECT 8.330 302.000 8.480 309.550 ;
        RECT 8.930 302.000 9.080 309.550 ;
        RECT 9.530 302.000 9.680 309.550 ;
        RECT 10.130 309.350 14.080 309.550 ;
        RECT 15.380 309.350 19.330 309.550 ;
        RECT 10.130 308.900 10.730 309.350 ;
        RECT 18.730 308.900 19.330 309.350 ;
        RECT 10.130 308.750 14.080 308.900 ;
        RECT 15.380 308.750 19.330 308.900 ;
        RECT 10.130 308.300 10.730 308.750 ;
        RECT 18.730 308.300 19.330 308.750 ;
        RECT 10.130 308.150 14.080 308.300 ;
        RECT 15.380 308.150 19.330 308.300 ;
        RECT 10.130 307.700 10.730 308.150 ;
        RECT 18.730 307.700 19.330 308.150 ;
        RECT 10.130 307.550 14.080 307.700 ;
        RECT 15.380 307.550 19.330 307.700 ;
        RECT 10.130 307.100 10.730 307.550 ;
        RECT 18.730 307.100 19.330 307.550 ;
        RECT 10.130 306.950 14.080 307.100 ;
        RECT 15.380 306.950 19.330 307.100 ;
        RECT 10.130 306.500 10.730 306.950 ;
        RECT 18.730 306.500 19.330 306.950 ;
        RECT 10.130 306.350 14.080 306.500 ;
        RECT 15.380 306.350 19.330 306.500 ;
        RECT 10.130 305.900 10.730 306.350 ;
        RECT 18.730 305.900 19.330 306.350 ;
        RECT 10.130 305.750 14.080 305.900 ;
        RECT 15.380 305.750 19.330 305.900 ;
        RECT 10.130 305.300 10.730 305.750 ;
        RECT 18.730 305.300 19.330 305.750 ;
        RECT 10.130 305.150 14.080 305.300 ;
        RECT 15.380 305.150 19.330 305.300 ;
        RECT 10.130 304.700 10.730 305.150 ;
        RECT 18.730 304.700 19.330 305.150 ;
        RECT 10.130 304.550 14.080 304.700 ;
        RECT 15.380 304.550 19.330 304.700 ;
        RECT 10.130 304.100 10.730 304.550 ;
        RECT 18.730 304.100 19.330 304.550 ;
        RECT 10.130 303.950 14.080 304.100 ;
        RECT 15.380 303.950 19.330 304.100 ;
        RECT 10.130 303.500 10.730 303.950 ;
        RECT 18.730 303.500 19.330 303.950 ;
        RECT 10.130 303.350 14.080 303.500 ;
        RECT 15.380 303.350 19.330 303.500 ;
        RECT 10.130 302.900 10.730 303.350 ;
        RECT 18.730 302.900 19.330 303.350 ;
        RECT 10.130 302.750 14.080 302.900 ;
        RECT 15.380 302.750 19.330 302.900 ;
        RECT 10.130 302.300 10.730 302.750 ;
        RECT 18.730 302.300 19.330 302.750 ;
        RECT 10.130 302.150 14.080 302.300 ;
        RECT 15.380 302.150 19.330 302.300 ;
        RECT 10.130 302.000 10.730 302.150 ;
        RECT 6.530 301.700 10.730 302.000 ;
        RECT 18.730 302.000 19.330 302.150 ;
        RECT 19.780 302.000 19.930 309.550 ;
        RECT 20.380 302.000 20.530 309.550 ;
        RECT 20.980 302.000 21.130 309.550 ;
        RECT 21.580 302.000 21.730 309.550 ;
        RECT 22.180 302.000 22.330 309.550 ;
        RECT 22.780 302.000 22.930 304.900 ;
        RECT 18.730 301.700 22.930 302.000 ;
        RECT 6.530 301.550 14.080 301.700 ;
        RECT 15.380 301.550 22.930 301.700 ;
        RECT 6.530 301.350 10.730 301.550 ;
        RECT 4.730 301.050 9.130 301.200 ;
        RECT 9.280 301.050 10.730 301.350 ;
        RECT 4.730 300.150 10.730 301.050 ;
        RECT 18.730 301.350 22.930 301.550 ;
        RECT 18.730 301.050 20.180 301.350 ;
        RECT 23.530 301.200 25.930 304.400 ;
        RECT 26.530 302.000 26.680 304.900 ;
        RECT 27.130 302.000 27.280 309.550 ;
        RECT 27.730 302.000 27.880 309.550 ;
        RECT 28.330 302.000 28.480 309.550 ;
        RECT 28.930 302.000 29.080 309.550 ;
        RECT 29.530 302.000 29.680 309.550 ;
        RECT 30.130 309.350 34.080 309.550 ;
        RECT 35.380 309.350 39.330 309.550 ;
        RECT 30.130 308.900 30.730 309.350 ;
        RECT 38.730 308.900 39.330 309.350 ;
        RECT 30.130 308.750 34.080 308.900 ;
        RECT 35.380 308.750 39.330 308.900 ;
        RECT 30.130 308.300 30.730 308.750 ;
        RECT 38.730 308.300 39.330 308.750 ;
        RECT 30.130 308.150 34.080 308.300 ;
        RECT 35.380 308.150 39.330 308.300 ;
        RECT 30.130 307.700 30.730 308.150 ;
        RECT 38.730 307.700 39.330 308.150 ;
        RECT 30.130 307.550 34.080 307.700 ;
        RECT 35.380 307.550 39.330 307.700 ;
        RECT 30.130 307.100 30.730 307.550 ;
        RECT 38.730 307.100 39.330 307.550 ;
        RECT 30.130 306.950 34.080 307.100 ;
        RECT 35.380 306.950 39.330 307.100 ;
        RECT 30.130 306.500 30.730 306.950 ;
        RECT 38.730 306.500 39.330 306.950 ;
        RECT 30.130 306.350 34.080 306.500 ;
        RECT 35.380 306.350 39.330 306.500 ;
        RECT 30.130 305.900 30.730 306.350 ;
        RECT 38.730 305.900 39.330 306.350 ;
        RECT 30.130 305.750 34.080 305.900 ;
        RECT 35.380 305.750 39.330 305.900 ;
        RECT 30.130 305.300 30.730 305.750 ;
        RECT 38.730 305.300 39.330 305.750 ;
        RECT 30.130 305.150 34.080 305.300 ;
        RECT 35.380 305.150 39.330 305.300 ;
        RECT 30.130 304.700 30.730 305.150 ;
        RECT 38.730 304.700 39.330 305.150 ;
        RECT 30.130 304.550 34.080 304.700 ;
        RECT 35.380 304.550 39.330 304.700 ;
        RECT 30.130 304.100 30.730 304.550 ;
        RECT 38.730 304.100 39.330 304.550 ;
        RECT 30.130 303.950 34.080 304.100 ;
        RECT 35.380 303.950 39.330 304.100 ;
        RECT 30.130 303.500 30.730 303.950 ;
        RECT 38.730 303.500 39.330 303.950 ;
        RECT 30.130 303.350 34.080 303.500 ;
        RECT 35.380 303.350 39.330 303.500 ;
        RECT 30.130 302.900 30.730 303.350 ;
        RECT 38.730 302.900 39.330 303.350 ;
        RECT 30.130 302.750 34.080 302.900 ;
        RECT 35.380 302.750 39.330 302.900 ;
        RECT 30.130 302.300 30.730 302.750 ;
        RECT 38.730 302.300 39.330 302.750 ;
        RECT 30.130 302.150 34.080 302.300 ;
        RECT 35.380 302.150 39.330 302.300 ;
        RECT 30.130 302.000 30.730 302.150 ;
        RECT 26.530 301.700 30.730 302.000 ;
        RECT 38.730 302.000 39.330 302.150 ;
        RECT 39.780 302.000 39.930 309.550 ;
        RECT 40.380 302.000 40.530 309.550 ;
        RECT 40.980 302.000 41.130 309.550 ;
        RECT 41.580 302.000 41.730 309.550 ;
        RECT 42.180 302.000 42.330 309.550 ;
        RECT 42.780 302.000 42.930 304.900 ;
        RECT 38.730 301.700 42.930 302.000 ;
        RECT 26.530 301.550 34.080 301.700 ;
        RECT 35.380 301.550 42.930 301.700 ;
        RECT 26.530 301.350 30.730 301.550 ;
        RECT 20.330 301.050 29.130 301.200 ;
        RECT 29.280 301.050 30.730 301.350 ;
        RECT 18.730 300.150 30.730 301.050 ;
        RECT 38.730 301.350 42.930 301.550 ;
        RECT 38.730 301.050 40.180 301.350 ;
        RECT 43.530 301.200 45.930 304.400 ;
        RECT 46.530 302.000 46.680 304.900 ;
        RECT 47.130 302.000 47.280 309.550 ;
        RECT 47.730 302.000 47.880 309.550 ;
        RECT 48.330 302.000 48.480 309.550 ;
        RECT 48.930 302.000 49.080 309.550 ;
        RECT 49.530 302.000 49.680 309.550 ;
        RECT 50.130 309.350 54.080 309.550 ;
        RECT 55.380 309.350 59.330 309.550 ;
        RECT 50.130 308.900 50.730 309.350 ;
        RECT 58.730 308.900 59.330 309.350 ;
        RECT 50.130 308.750 54.080 308.900 ;
        RECT 55.380 308.750 59.330 308.900 ;
        RECT 50.130 308.300 50.730 308.750 ;
        RECT 58.730 308.300 59.330 308.750 ;
        RECT 50.130 308.150 54.080 308.300 ;
        RECT 55.380 308.150 59.330 308.300 ;
        RECT 50.130 307.700 50.730 308.150 ;
        RECT 58.730 307.700 59.330 308.150 ;
        RECT 50.130 307.550 54.080 307.700 ;
        RECT 55.380 307.550 59.330 307.700 ;
        RECT 50.130 307.100 50.730 307.550 ;
        RECT 58.730 307.100 59.330 307.550 ;
        RECT 50.130 306.950 54.080 307.100 ;
        RECT 55.380 306.950 59.330 307.100 ;
        RECT 50.130 306.500 50.730 306.950 ;
        RECT 58.730 306.500 59.330 306.950 ;
        RECT 50.130 306.350 54.080 306.500 ;
        RECT 55.380 306.350 59.330 306.500 ;
        RECT 50.130 305.900 50.730 306.350 ;
        RECT 58.730 305.900 59.330 306.350 ;
        RECT 50.130 305.750 54.080 305.900 ;
        RECT 55.380 305.750 59.330 305.900 ;
        RECT 50.130 305.300 50.730 305.750 ;
        RECT 58.730 305.300 59.330 305.750 ;
        RECT 50.130 305.150 54.080 305.300 ;
        RECT 55.380 305.150 59.330 305.300 ;
        RECT 50.130 304.700 50.730 305.150 ;
        RECT 58.730 304.700 59.330 305.150 ;
        RECT 50.130 304.550 54.080 304.700 ;
        RECT 55.380 304.550 59.330 304.700 ;
        RECT 50.130 304.100 50.730 304.550 ;
        RECT 58.730 304.100 59.330 304.550 ;
        RECT 50.130 303.950 54.080 304.100 ;
        RECT 55.380 303.950 59.330 304.100 ;
        RECT 50.130 303.500 50.730 303.950 ;
        RECT 58.730 303.500 59.330 303.950 ;
        RECT 50.130 303.350 54.080 303.500 ;
        RECT 55.380 303.350 59.330 303.500 ;
        RECT 50.130 302.900 50.730 303.350 ;
        RECT 58.730 302.900 59.330 303.350 ;
        RECT 50.130 302.750 54.080 302.900 ;
        RECT 55.380 302.750 59.330 302.900 ;
        RECT 50.130 302.300 50.730 302.750 ;
        RECT 58.730 302.300 59.330 302.750 ;
        RECT 50.130 302.150 54.080 302.300 ;
        RECT 55.380 302.150 59.330 302.300 ;
        RECT 50.130 302.000 50.730 302.150 ;
        RECT 46.530 301.700 50.730 302.000 ;
        RECT 58.730 302.000 59.330 302.150 ;
        RECT 59.780 302.000 59.930 309.550 ;
        RECT 60.380 302.000 60.530 309.550 ;
        RECT 60.980 302.000 61.130 309.550 ;
        RECT 61.580 302.000 61.730 309.550 ;
        RECT 62.180 302.000 62.330 309.550 ;
        RECT 62.780 302.000 62.930 304.900 ;
        RECT 58.730 301.700 62.930 302.000 ;
        RECT 46.530 301.550 54.080 301.700 ;
        RECT 55.380 301.550 62.930 301.700 ;
        RECT 46.530 301.350 50.730 301.550 ;
        RECT 40.330 301.050 49.130 301.200 ;
        RECT 49.280 301.050 50.730 301.350 ;
        RECT 38.730 300.150 50.730 301.050 ;
        RECT 58.730 301.350 62.930 301.550 ;
        RECT 58.730 301.050 60.180 301.350 ;
        RECT 63.530 301.200 65.930 304.400 ;
        RECT 66.530 302.000 66.680 304.900 ;
        RECT 67.130 302.000 67.280 309.550 ;
        RECT 67.730 302.000 67.880 309.550 ;
        RECT 68.330 302.000 68.480 309.550 ;
        RECT 68.930 302.000 69.080 309.550 ;
        RECT 69.530 302.000 69.680 309.550 ;
        RECT 70.130 309.350 74.080 309.550 ;
        RECT 75.380 309.350 79.330 309.550 ;
        RECT 70.130 308.900 70.730 309.350 ;
        RECT 78.730 308.900 79.330 309.350 ;
        RECT 70.130 308.750 74.080 308.900 ;
        RECT 75.380 308.750 79.330 308.900 ;
        RECT 70.130 308.300 70.730 308.750 ;
        RECT 78.730 308.300 79.330 308.750 ;
        RECT 70.130 308.150 74.080 308.300 ;
        RECT 75.380 308.150 79.330 308.300 ;
        RECT 70.130 307.700 70.730 308.150 ;
        RECT 78.730 307.700 79.330 308.150 ;
        RECT 70.130 307.550 74.080 307.700 ;
        RECT 75.380 307.550 79.330 307.700 ;
        RECT 70.130 307.100 70.730 307.550 ;
        RECT 78.730 307.100 79.330 307.550 ;
        RECT 70.130 306.950 74.080 307.100 ;
        RECT 75.380 306.950 79.330 307.100 ;
        RECT 70.130 306.500 70.730 306.950 ;
        RECT 78.730 306.500 79.330 306.950 ;
        RECT 70.130 306.350 74.080 306.500 ;
        RECT 75.380 306.350 79.330 306.500 ;
        RECT 70.130 305.900 70.730 306.350 ;
        RECT 78.730 305.900 79.330 306.350 ;
        RECT 70.130 305.750 74.080 305.900 ;
        RECT 75.380 305.750 79.330 305.900 ;
        RECT 70.130 305.300 70.730 305.750 ;
        RECT 78.730 305.300 79.330 305.750 ;
        RECT 70.130 305.150 74.080 305.300 ;
        RECT 75.380 305.150 79.330 305.300 ;
        RECT 70.130 304.700 70.730 305.150 ;
        RECT 78.730 304.700 79.330 305.150 ;
        RECT 70.130 304.550 74.080 304.700 ;
        RECT 75.380 304.550 79.330 304.700 ;
        RECT 70.130 304.100 70.730 304.550 ;
        RECT 78.730 304.100 79.330 304.550 ;
        RECT 70.130 303.950 74.080 304.100 ;
        RECT 75.380 303.950 79.330 304.100 ;
        RECT 70.130 303.500 70.730 303.950 ;
        RECT 78.730 303.500 79.330 303.950 ;
        RECT 70.130 303.350 74.080 303.500 ;
        RECT 75.380 303.350 79.330 303.500 ;
        RECT 70.130 302.900 70.730 303.350 ;
        RECT 78.730 302.900 79.330 303.350 ;
        RECT 70.130 302.750 74.080 302.900 ;
        RECT 75.380 302.750 79.330 302.900 ;
        RECT 70.130 302.300 70.730 302.750 ;
        RECT 78.730 302.300 79.330 302.750 ;
        RECT 70.130 302.150 74.080 302.300 ;
        RECT 75.380 302.150 79.330 302.300 ;
        RECT 70.130 302.000 70.730 302.150 ;
        RECT 66.530 301.700 70.730 302.000 ;
        RECT 78.730 302.000 79.330 302.150 ;
        RECT 79.780 302.000 79.930 309.550 ;
        RECT 80.380 302.000 80.530 309.550 ;
        RECT 80.980 302.000 81.130 309.550 ;
        RECT 81.580 302.000 81.730 309.550 ;
        RECT 82.180 302.000 82.330 309.550 ;
        RECT 82.780 302.000 82.930 304.900 ;
        RECT 78.730 301.700 82.930 302.000 ;
        RECT 66.530 301.550 74.080 301.700 ;
        RECT 75.380 301.550 82.930 301.700 ;
        RECT 66.530 301.350 70.730 301.550 ;
        RECT 60.330 301.050 69.130 301.200 ;
        RECT 69.280 301.050 70.730 301.350 ;
        RECT 58.730 300.150 70.730 301.050 ;
        RECT 78.730 301.350 82.930 301.550 ;
        RECT 78.730 301.050 80.180 301.350 ;
        RECT 83.530 301.200 85.930 304.400 ;
        RECT 86.530 302.000 86.680 304.900 ;
        RECT 87.130 302.000 87.280 309.550 ;
        RECT 87.730 302.000 87.880 309.550 ;
        RECT 88.330 302.000 88.480 309.550 ;
        RECT 88.930 302.000 89.080 309.550 ;
        RECT 89.530 302.000 89.680 309.550 ;
        RECT 90.130 309.350 94.080 309.550 ;
        RECT 95.380 309.350 99.330 309.550 ;
        RECT 90.130 308.900 90.730 309.350 ;
        RECT 98.730 308.900 99.330 309.350 ;
        RECT 90.130 308.750 94.080 308.900 ;
        RECT 95.380 308.750 99.330 308.900 ;
        RECT 90.130 308.300 90.730 308.750 ;
        RECT 98.730 308.300 99.330 308.750 ;
        RECT 90.130 308.150 94.080 308.300 ;
        RECT 95.380 308.150 99.330 308.300 ;
        RECT 90.130 307.700 90.730 308.150 ;
        RECT 98.730 307.700 99.330 308.150 ;
        RECT 90.130 307.550 94.080 307.700 ;
        RECT 95.380 307.550 99.330 307.700 ;
        RECT 90.130 307.100 90.730 307.550 ;
        RECT 98.730 307.100 99.330 307.550 ;
        RECT 90.130 306.950 94.080 307.100 ;
        RECT 95.380 306.950 99.330 307.100 ;
        RECT 90.130 306.500 90.730 306.950 ;
        RECT 98.730 306.500 99.330 306.950 ;
        RECT 90.130 306.350 94.080 306.500 ;
        RECT 95.380 306.350 99.330 306.500 ;
        RECT 90.130 305.900 90.730 306.350 ;
        RECT 98.730 305.900 99.330 306.350 ;
        RECT 90.130 305.750 94.080 305.900 ;
        RECT 95.380 305.750 99.330 305.900 ;
        RECT 90.130 305.300 90.730 305.750 ;
        RECT 98.730 305.300 99.330 305.750 ;
        RECT 90.130 305.150 94.080 305.300 ;
        RECT 95.380 305.150 99.330 305.300 ;
        RECT 90.130 304.700 90.730 305.150 ;
        RECT 98.730 304.700 99.330 305.150 ;
        RECT 90.130 304.550 94.080 304.700 ;
        RECT 95.380 304.550 99.330 304.700 ;
        RECT 90.130 304.100 90.730 304.550 ;
        RECT 98.730 304.100 99.330 304.550 ;
        RECT 90.130 303.950 94.080 304.100 ;
        RECT 95.380 303.950 99.330 304.100 ;
        RECT 90.130 303.500 90.730 303.950 ;
        RECT 98.730 303.500 99.330 303.950 ;
        RECT 90.130 303.350 94.080 303.500 ;
        RECT 95.380 303.350 99.330 303.500 ;
        RECT 90.130 302.900 90.730 303.350 ;
        RECT 98.730 302.900 99.330 303.350 ;
        RECT 90.130 302.750 94.080 302.900 ;
        RECT 95.380 302.750 99.330 302.900 ;
        RECT 90.130 302.300 90.730 302.750 ;
        RECT 98.730 302.300 99.330 302.750 ;
        RECT 90.130 302.150 94.080 302.300 ;
        RECT 95.380 302.150 99.330 302.300 ;
        RECT 90.130 302.000 90.730 302.150 ;
        RECT 86.530 301.700 90.730 302.000 ;
        RECT 98.730 302.000 99.330 302.150 ;
        RECT 99.780 302.000 99.930 309.550 ;
        RECT 100.380 302.000 100.530 309.550 ;
        RECT 100.980 302.000 101.130 309.550 ;
        RECT 101.580 302.000 101.730 309.550 ;
        RECT 102.180 302.000 102.330 309.550 ;
        RECT 102.780 302.000 102.930 304.900 ;
        RECT 98.730 301.700 102.930 302.000 ;
        RECT 86.530 301.550 94.080 301.700 ;
        RECT 95.380 301.550 102.930 301.700 ;
        RECT 86.530 301.350 90.730 301.550 ;
        RECT 80.330 301.050 89.130 301.200 ;
        RECT 89.280 301.050 90.730 301.350 ;
        RECT 78.730 300.150 90.730 301.050 ;
        RECT 98.730 301.350 102.930 301.550 ;
        RECT 103.530 303.600 104.730 304.400 ;
        RECT 103.530 302.325 107.140 303.600 ;
        RECT 98.730 301.050 100.180 301.350 ;
        RECT 103.530 301.200 104.730 302.325 ;
        RECT 100.330 301.050 104.730 301.200 ;
        RECT 98.730 300.150 104.730 301.050 ;
        RECT 4.730 299.850 9.130 300.150 ;
        RECT 20.330 299.850 29.130 300.150 ;
        RECT 40.330 299.850 49.130 300.150 ;
        RECT 60.330 299.850 69.130 300.150 ;
        RECT 80.330 299.850 89.130 300.150 ;
        RECT 4.730 298.950 10.730 299.850 ;
        RECT 20.330 299.800 30.730 299.850 ;
        RECT 40.330 299.800 50.730 299.850 ;
        RECT 60.330 299.800 70.730 299.850 ;
        RECT 80.330 299.800 90.730 299.850 ;
        RECT 100.330 299.800 104.730 300.150 ;
        RECT 4.730 298.800 9.130 298.950 ;
        RECT 4.730 297.530 5.930 298.800 ;
        RECT 9.280 298.650 10.730 298.950 ;
        RECT 2.315 296.255 5.930 297.530 ;
        RECT 4.730 295.600 5.930 296.255 ;
        RECT 6.530 298.450 10.730 298.650 ;
        RECT 18.730 298.950 30.730 299.800 ;
        RECT 18.730 298.900 29.130 298.950 ;
        RECT 18.730 298.650 20.180 298.900 ;
        RECT 20.330 298.800 29.130 298.900 ;
        RECT 18.730 298.450 22.930 298.650 ;
        RECT 6.530 298.300 14.080 298.450 ;
        RECT 15.430 298.300 22.930 298.450 ;
        RECT 6.530 298.000 10.730 298.300 ;
        RECT 2.320 295.340 4.320 295.545 ;
        RECT 2.315 293.250 4.320 295.340 ;
        RECT 6.530 295.150 6.680 298.000 ;
        RECT 7.130 290.450 7.280 298.000 ;
        RECT 7.730 290.450 7.880 298.000 ;
        RECT 8.330 290.450 8.480 298.000 ;
        RECT 8.930 290.450 9.080 298.000 ;
        RECT 9.530 290.450 9.680 298.000 ;
        RECT 10.130 297.850 10.730 298.000 ;
        RECT 18.730 298.000 22.930 298.300 ;
        RECT 18.730 297.850 19.330 298.000 ;
        RECT 10.130 297.700 14.080 297.850 ;
        RECT 15.380 297.700 19.330 297.850 ;
        RECT 10.130 297.250 10.730 297.700 ;
        RECT 18.730 297.250 19.330 297.700 ;
        RECT 10.130 297.100 14.080 297.250 ;
        RECT 15.380 297.100 19.330 297.250 ;
        RECT 10.130 296.650 10.730 297.100 ;
        RECT 18.730 296.650 19.330 297.100 ;
        RECT 10.130 296.500 14.080 296.650 ;
        RECT 15.380 296.500 19.330 296.650 ;
        RECT 10.130 296.050 10.730 296.500 ;
        RECT 18.730 296.050 19.330 296.500 ;
        RECT 10.130 295.900 14.080 296.050 ;
        RECT 15.380 295.900 19.330 296.050 ;
        RECT 10.130 295.450 10.730 295.900 ;
        RECT 18.730 295.450 19.330 295.900 ;
        RECT 10.130 295.300 14.080 295.450 ;
        RECT 15.380 295.300 19.330 295.450 ;
        RECT 10.130 294.850 10.730 295.300 ;
        RECT 18.730 294.850 19.330 295.300 ;
        RECT 10.130 294.700 14.080 294.850 ;
        RECT 15.380 294.700 19.330 294.850 ;
        RECT 10.130 294.250 10.730 294.700 ;
        RECT 18.730 294.250 19.330 294.700 ;
        RECT 10.130 294.100 14.080 294.250 ;
        RECT 15.380 294.100 19.330 294.250 ;
        RECT 10.130 293.650 10.730 294.100 ;
        RECT 18.730 293.650 19.330 294.100 ;
        RECT 10.130 293.500 14.080 293.650 ;
        RECT 15.380 293.500 19.330 293.650 ;
        RECT 10.130 293.050 10.730 293.500 ;
        RECT 18.730 293.050 19.330 293.500 ;
        RECT 10.130 292.900 14.080 293.050 ;
        RECT 15.380 292.900 19.330 293.050 ;
        RECT 10.130 292.450 10.730 292.900 ;
        RECT 18.730 292.450 19.330 292.900 ;
        RECT 10.130 292.300 14.080 292.450 ;
        RECT 15.380 292.300 19.330 292.450 ;
        RECT 10.130 291.850 10.730 292.300 ;
        RECT 18.730 291.850 19.330 292.300 ;
        RECT 10.130 291.700 14.080 291.850 ;
        RECT 15.380 291.700 19.330 291.850 ;
        RECT 10.130 291.250 10.730 291.700 ;
        RECT 18.730 291.250 19.330 291.700 ;
        RECT 10.130 291.100 14.080 291.250 ;
        RECT 15.380 291.100 19.330 291.250 ;
        RECT 10.130 290.650 10.730 291.100 ;
        RECT 18.730 290.650 19.330 291.100 ;
        RECT 10.130 290.450 14.080 290.650 ;
        RECT 15.380 290.450 19.330 290.650 ;
        RECT 19.780 290.450 19.930 298.000 ;
        RECT 20.380 290.450 20.530 298.000 ;
        RECT 20.980 290.450 21.130 298.000 ;
        RECT 21.580 290.450 21.730 298.000 ;
        RECT 22.180 290.450 22.330 298.000 ;
        RECT 22.780 295.150 22.930 298.000 ;
        RECT 23.530 295.600 25.930 298.800 ;
        RECT 29.280 298.650 30.730 298.950 ;
        RECT 26.530 298.450 30.730 298.650 ;
        RECT 38.730 298.950 50.730 299.800 ;
        RECT 38.730 298.900 49.130 298.950 ;
        RECT 38.730 298.650 40.180 298.900 ;
        RECT 40.330 298.800 49.130 298.900 ;
        RECT 38.730 298.450 42.930 298.650 ;
        RECT 26.530 298.300 34.080 298.450 ;
        RECT 35.430 298.300 42.930 298.450 ;
        RECT 26.530 298.000 30.730 298.300 ;
        RECT 26.530 295.150 26.680 298.000 ;
        RECT 27.130 290.450 27.280 298.000 ;
        RECT 27.730 290.450 27.880 298.000 ;
        RECT 28.330 290.450 28.480 298.000 ;
        RECT 28.930 290.450 29.080 298.000 ;
        RECT 29.530 290.450 29.680 298.000 ;
        RECT 30.130 297.850 30.730 298.000 ;
        RECT 38.730 298.000 42.930 298.300 ;
        RECT 38.730 297.850 39.330 298.000 ;
        RECT 30.130 297.700 34.080 297.850 ;
        RECT 35.380 297.700 39.330 297.850 ;
        RECT 30.130 297.250 30.730 297.700 ;
        RECT 38.730 297.250 39.330 297.700 ;
        RECT 30.130 297.100 34.080 297.250 ;
        RECT 35.380 297.100 39.330 297.250 ;
        RECT 30.130 296.650 30.730 297.100 ;
        RECT 38.730 296.650 39.330 297.100 ;
        RECT 30.130 296.500 34.080 296.650 ;
        RECT 35.380 296.500 39.330 296.650 ;
        RECT 30.130 296.050 30.730 296.500 ;
        RECT 38.730 296.050 39.330 296.500 ;
        RECT 30.130 295.900 34.080 296.050 ;
        RECT 35.380 295.900 39.330 296.050 ;
        RECT 30.130 295.450 30.730 295.900 ;
        RECT 38.730 295.450 39.330 295.900 ;
        RECT 30.130 295.300 34.080 295.450 ;
        RECT 35.380 295.300 39.330 295.450 ;
        RECT 30.130 294.850 30.730 295.300 ;
        RECT 38.730 294.850 39.330 295.300 ;
        RECT 30.130 294.700 34.080 294.850 ;
        RECT 35.380 294.700 39.330 294.850 ;
        RECT 30.130 294.250 30.730 294.700 ;
        RECT 38.730 294.250 39.330 294.700 ;
        RECT 30.130 294.100 34.080 294.250 ;
        RECT 35.380 294.100 39.330 294.250 ;
        RECT 30.130 293.650 30.730 294.100 ;
        RECT 38.730 293.650 39.330 294.100 ;
        RECT 30.130 293.500 34.080 293.650 ;
        RECT 35.380 293.500 39.330 293.650 ;
        RECT 30.130 293.050 30.730 293.500 ;
        RECT 38.730 293.050 39.330 293.500 ;
        RECT 30.130 292.900 34.080 293.050 ;
        RECT 35.380 292.900 39.330 293.050 ;
        RECT 30.130 292.450 30.730 292.900 ;
        RECT 38.730 292.450 39.330 292.900 ;
        RECT 30.130 292.300 34.080 292.450 ;
        RECT 35.380 292.300 39.330 292.450 ;
        RECT 30.130 291.850 30.730 292.300 ;
        RECT 38.730 291.850 39.330 292.300 ;
        RECT 30.130 291.700 34.080 291.850 ;
        RECT 35.380 291.700 39.330 291.850 ;
        RECT 30.130 291.250 30.730 291.700 ;
        RECT 38.730 291.250 39.330 291.700 ;
        RECT 30.130 291.100 34.080 291.250 ;
        RECT 35.380 291.100 39.330 291.250 ;
        RECT 30.130 290.650 30.730 291.100 ;
        RECT 38.730 290.650 39.330 291.100 ;
        RECT 30.130 290.450 34.080 290.650 ;
        RECT 35.380 290.450 39.330 290.650 ;
        RECT 39.780 290.450 39.930 298.000 ;
        RECT 40.380 290.450 40.530 298.000 ;
        RECT 40.980 290.450 41.130 298.000 ;
        RECT 41.580 290.450 41.730 298.000 ;
        RECT 42.180 290.450 42.330 298.000 ;
        RECT 42.780 295.150 42.930 298.000 ;
        RECT 43.530 295.600 45.930 298.800 ;
        RECT 49.280 298.650 50.730 298.950 ;
        RECT 46.530 298.450 50.730 298.650 ;
        RECT 58.730 298.950 70.730 299.800 ;
        RECT 58.730 298.900 69.130 298.950 ;
        RECT 58.730 298.650 60.180 298.900 ;
        RECT 60.330 298.800 69.130 298.900 ;
        RECT 58.730 298.450 62.930 298.650 ;
        RECT 46.530 298.300 54.080 298.450 ;
        RECT 55.430 298.300 62.930 298.450 ;
        RECT 46.530 298.000 50.730 298.300 ;
        RECT 46.530 295.150 46.680 298.000 ;
        RECT 47.130 290.450 47.280 298.000 ;
        RECT 47.730 290.450 47.880 298.000 ;
        RECT 48.330 290.450 48.480 298.000 ;
        RECT 48.930 290.450 49.080 298.000 ;
        RECT 49.530 290.450 49.680 298.000 ;
        RECT 50.130 297.850 50.730 298.000 ;
        RECT 58.730 298.000 62.930 298.300 ;
        RECT 58.730 297.850 59.330 298.000 ;
        RECT 50.130 297.700 54.080 297.850 ;
        RECT 55.380 297.700 59.330 297.850 ;
        RECT 50.130 297.250 50.730 297.700 ;
        RECT 58.730 297.250 59.330 297.700 ;
        RECT 50.130 297.100 54.080 297.250 ;
        RECT 55.380 297.100 59.330 297.250 ;
        RECT 50.130 296.650 50.730 297.100 ;
        RECT 58.730 296.650 59.330 297.100 ;
        RECT 50.130 296.500 54.080 296.650 ;
        RECT 55.380 296.500 59.330 296.650 ;
        RECT 50.130 296.050 50.730 296.500 ;
        RECT 58.730 296.050 59.330 296.500 ;
        RECT 50.130 295.900 54.080 296.050 ;
        RECT 55.380 295.900 59.330 296.050 ;
        RECT 50.130 295.450 50.730 295.900 ;
        RECT 58.730 295.450 59.330 295.900 ;
        RECT 50.130 295.300 54.080 295.450 ;
        RECT 55.380 295.300 59.330 295.450 ;
        RECT 50.130 294.850 50.730 295.300 ;
        RECT 58.730 294.850 59.330 295.300 ;
        RECT 50.130 294.700 54.080 294.850 ;
        RECT 55.380 294.700 59.330 294.850 ;
        RECT 50.130 294.250 50.730 294.700 ;
        RECT 58.730 294.250 59.330 294.700 ;
        RECT 50.130 294.100 54.080 294.250 ;
        RECT 55.380 294.100 59.330 294.250 ;
        RECT 50.130 293.650 50.730 294.100 ;
        RECT 58.730 293.650 59.330 294.100 ;
        RECT 50.130 293.500 54.080 293.650 ;
        RECT 55.380 293.500 59.330 293.650 ;
        RECT 50.130 293.050 50.730 293.500 ;
        RECT 58.730 293.050 59.330 293.500 ;
        RECT 50.130 292.900 54.080 293.050 ;
        RECT 55.380 292.900 59.330 293.050 ;
        RECT 50.130 292.450 50.730 292.900 ;
        RECT 58.730 292.450 59.330 292.900 ;
        RECT 50.130 292.300 54.080 292.450 ;
        RECT 55.380 292.300 59.330 292.450 ;
        RECT 50.130 291.850 50.730 292.300 ;
        RECT 58.730 291.850 59.330 292.300 ;
        RECT 50.130 291.700 54.080 291.850 ;
        RECT 55.380 291.700 59.330 291.850 ;
        RECT 50.130 291.250 50.730 291.700 ;
        RECT 58.730 291.250 59.330 291.700 ;
        RECT 50.130 291.100 54.080 291.250 ;
        RECT 55.380 291.100 59.330 291.250 ;
        RECT 50.130 290.650 50.730 291.100 ;
        RECT 58.730 290.650 59.330 291.100 ;
        RECT 50.130 290.450 54.080 290.650 ;
        RECT 55.380 290.450 59.330 290.650 ;
        RECT 59.780 290.450 59.930 298.000 ;
        RECT 60.380 290.450 60.530 298.000 ;
        RECT 60.980 290.450 61.130 298.000 ;
        RECT 61.580 290.450 61.730 298.000 ;
        RECT 62.180 290.450 62.330 298.000 ;
        RECT 62.780 295.150 62.930 298.000 ;
        RECT 63.530 295.600 65.930 298.800 ;
        RECT 69.280 298.650 70.730 298.950 ;
        RECT 66.530 298.450 70.730 298.650 ;
        RECT 78.730 298.950 90.730 299.800 ;
        RECT 78.730 298.900 89.130 298.950 ;
        RECT 78.730 298.650 80.180 298.900 ;
        RECT 80.330 298.800 89.130 298.900 ;
        RECT 78.730 298.450 82.930 298.650 ;
        RECT 66.530 298.300 74.080 298.450 ;
        RECT 75.430 298.300 82.930 298.450 ;
        RECT 66.530 298.000 70.730 298.300 ;
        RECT 66.530 295.150 66.680 298.000 ;
        RECT 67.130 290.450 67.280 298.000 ;
        RECT 67.730 290.450 67.880 298.000 ;
        RECT 68.330 290.450 68.480 298.000 ;
        RECT 68.930 290.450 69.080 298.000 ;
        RECT 69.530 290.450 69.680 298.000 ;
        RECT 70.130 297.850 70.730 298.000 ;
        RECT 78.730 298.000 82.930 298.300 ;
        RECT 78.730 297.850 79.330 298.000 ;
        RECT 70.130 297.700 74.080 297.850 ;
        RECT 75.380 297.700 79.330 297.850 ;
        RECT 70.130 297.250 70.730 297.700 ;
        RECT 78.730 297.250 79.330 297.700 ;
        RECT 70.130 297.100 74.080 297.250 ;
        RECT 75.380 297.100 79.330 297.250 ;
        RECT 70.130 296.650 70.730 297.100 ;
        RECT 78.730 296.650 79.330 297.100 ;
        RECT 70.130 296.500 74.080 296.650 ;
        RECT 75.380 296.500 79.330 296.650 ;
        RECT 70.130 296.050 70.730 296.500 ;
        RECT 78.730 296.050 79.330 296.500 ;
        RECT 70.130 295.900 74.080 296.050 ;
        RECT 75.380 295.900 79.330 296.050 ;
        RECT 70.130 295.450 70.730 295.900 ;
        RECT 78.730 295.450 79.330 295.900 ;
        RECT 70.130 295.300 74.080 295.450 ;
        RECT 75.380 295.300 79.330 295.450 ;
        RECT 70.130 294.850 70.730 295.300 ;
        RECT 78.730 294.850 79.330 295.300 ;
        RECT 70.130 294.700 74.080 294.850 ;
        RECT 75.380 294.700 79.330 294.850 ;
        RECT 70.130 294.250 70.730 294.700 ;
        RECT 78.730 294.250 79.330 294.700 ;
        RECT 70.130 294.100 74.080 294.250 ;
        RECT 75.380 294.100 79.330 294.250 ;
        RECT 70.130 293.650 70.730 294.100 ;
        RECT 78.730 293.650 79.330 294.100 ;
        RECT 70.130 293.500 74.080 293.650 ;
        RECT 75.380 293.500 79.330 293.650 ;
        RECT 70.130 293.050 70.730 293.500 ;
        RECT 78.730 293.050 79.330 293.500 ;
        RECT 70.130 292.900 74.080 293.050 ;
        RECT 75.380 292.900 79.330 293.050 ;
        RECT 70.130 292.450 70.730 292.900 ;
        RECT 78.730 292.450 79.330 292.900 ;
        RECT 70.130 292.300 74.080 292.450 ;
        RECT 75.380 292.300 79.330 292.450 ;
        RECT 70.130 291.850 70.730 292.300 ;
        RECT 78.730 291.850 79.330 292.300 ;
        RECT 70.130 291.700 74.080 291.850 ;
        RECT 75.380 291.700 79.330 291.850 ;
        RECT 70.130 291.250 70.730 291.700 ;
        RECT 78.730 291.250 79.330 291.700 ;
        RECT 70.130 291.100 74.080 291.250 ;
        RECT 75.380 291.100 79.330 291.250 ;
        RECT 70.130 290.650 70.730 291.100 ;
        RECT 78.730 290.650 79.330 291.100 ;
        RECT 70.130 290.450 74.080 290.650 ;
        RECT 75.380 290.450 79.330 290.650 ;
        RECT 79.780 290.450 79.930 298.000 ;
        RECT 80.380 290.450 80.530 298.000 ;
        RECT 80.980 290.450 81.130 298.000 ;
        RECT 81.580 290.450 81.730 298.000 ;
        RECT 82.180 290.450 82.330 298.000 ;
        RECT 82.780 295.150 82.930 298.000 ;
        RECT 83.530 295.600 85.930 298.800 ;
        RECT 89.280 298.650 90.730 298.950 ;
        RECT 86.530 298.450 90.730 298.650 ;
        RECT 98.730 298.900 104.730 299.800 ;
        RECT 98.730 298.650 100.180 298.900 ;
        RECT 100.330 298.800 104.730 298.900 ;
        RECT 98.730 298.450 102.930 298.650 ;
        RECT 86.530 298.300 94.080 298.450 ;
        RECT 95.430 298.300 102.930 298.450 ;
        RECT 86.530 298.000 90.730 298.300 ;
        RECT 86.530 295.150 86.680 298.000 ;
        RECT 87.130 290.450 87.280 298.000 ;
        RECT 87.730 290.450 87.880 298.000 ;
        RECT 88.330 290.450 88.480 298.000 ;
        RECT 88.930 290.450 89.080 298.000 ;
        RECT 89.530 290.450 89.680 298.000 ;
        RECT 90.130 297.850 90.730 298.000 ;
        RECT 98.730 298.000 102.930 298.300 ;
        RECT 98.730 297.850 99.330 298.000 ;
        RECT 90.130 297.700 94.080 297.850 ;
        RECT 95.380 297.700 99.330 297.850 ;
        RECT 90.130 297.250 90.730 297.700 ;
        RECT 98.730 297.250 99.330 297.700 ;
        RECT 90.130 297.100 94.080 297.250 ;
        RECT 95.380 297.100 99.330 297.250 ;
        RECT 90.130 296.650 90.730 297.100 ;
        RECT 98.730 296.650 99.330 297.100 ;
        RECT 90.130 296.500 94.080 296.650 ;
        RECT 95.380 296.500 99.330 296.650 ;
        RECT 90.130 296.050 90.730 296.500 ;
        RECT 98.730 296.050 99.330 296.500 ;
        RECT 90.130 295.900 94.080 296.050 ;
        RECT 95.380 295.900 99.330 296.050 ;
        RECT 90.130 295.450 90.730 295.900 ;
        RECT 98.730 295.450 99.330 295.900 ;
        RECT 90.130 295.300 94.080 295.450 ;
        RECT 95.380 295.300 99.330 295.450 ;
        RECT 90.130 294.850 90.730 295.300 ;
        RECT 98.730 294.850 99.330 295.300 ;
        RECT 90.130 294.700 94.080 294.850 ;
        RECT 95.380 294.700 99.330 294.850 ;
        RECT 90.130 294.250 90.730 294.700 ;
        RECT 98.730 294.250 99.330 294.700 ;
        RECT 90.130 294.100 94.080 294.250 ;
        RECT 95.380 294.100 99.330 294.250 ;
        RECT 90.130 293.650 90.730 294.100 ;
        RECT 98.730 293.650 99.330 294.100 ;
        RECT 90.130 293.500 94.080 293.650 ;
        RECT 95.380 293.500 99.330 293.650 ;
        RECT 90.130 293.050 90.730 293.500 ;
        RECT 98.730 293.050 99.330 293.500 ;
        RECT 90.130 292.900 94.080 293.050 ;
        RECT 95.380 292.900 99.330 293.050 ;
        RECT 90.130 292.450 90.730 292.900 ;
        RECT 98.730 292.450 99.330 292.900 ;
        RECT 90.130 292.300 94.080 292.450 ;
        RECT 95.380 292.300 99.330 292.450 ;
        RECT 90.130 291.850 90.730 292.300 ;
        RECT 98.730 291.850 99.330 292.300 ;
        RECT 90.130 291.700 94.080 291.850 ;
        RECT 95.380 291.700 99.330 291.850 ;
        RECT 90.130 291.250 90.730 291.700 ;
        RECT 98.730 291.250 99.330 291.700 ;
        RECT 90.130 291.100 94.080 291.250 ;
        RECT 95.380 291.100 99.330 291.250 ;
        RECT 90.130 290.650 90.730 291.100 ;
        RECT 98.730 290.650 99.330 291.100 ;
        RECT 90.130 290.450 94.080 290.650 ;
        RECT 95.380 290.450 99.330 290.650 ;
        RECT 99.780 290.450 99.930 298.000 ;
        RECT 100.380 290.450 100.530 298.000 ;
        RECT 100.980 290.450 101.130 298.000 ;
        RECT 101.580 290.450 101.730 298.000 ;
        RECT 102.180 290.450 102.330 298.000 ;
        RECT 102.780 295.150 102.930 298.000 ;
        RECT 103.530 297.855 104.730 298.800 ;
        RECT 103.530 296.580 107.135 297.855 ;
        RECT 103.530 295.600 104.730 296.580 ;
        RECT 2.315 284.445 4.315 286.740 ;
        RECT 4.730 283.645 5.930 284.400 ;
        RECT 2.315 282.370 5.930 283.645 ;
        RECT 4.730 281.200 5.930 282.370 ;
        RECT 6.530 282.000 6.680 284.900 ;
        RECT 7.130 282.000 7.280 289.550 ;
        RECT 7.730 282.000 7.880 289.550 ;
        RECT 8.330 282.000 8.480 289.550 ;
        RECT 8.930 282.000 9.080 289.550 ;
        RECT 9.530 282.000 9.680 289.550 ;
        RECT 10.130 289.350 14.080 289.550 ;
        RECT 15.380 289.350 19.330 289.550 ;
        RECT 10.130 288.900 10.730 289.350 ;
        RECT 18.730 288.900 19.330 289.350 ;
        RECT 10.130 288.750 14.080 288.900 ;
        RECT 15.380 288.750 19.330 288.900 ;
        RECT 10.130 288.300 10.730 288.750 ;
        RECT 18.730 288.300 19.330 288.750 ;
        RECT 10.130 288.150 14.080 288.300 ;
        RECT 15.380 288.150 19.330 288.300 ;
        RECT 10.130 287.700 10.730 288.150 ;
        RECT 18.730 287.700 19.330 288.150 ;
        RECT 10.130 287.550 14.080 287.700 ;
        RECT 15.380 287.550 19.330 287.700 ;
        RECT 10.130 287.100 10.730 287.550 ;
        RECT 18.730 287.100 19.330 287.550 ;
        RECT 10.130 286.950 14.080 287.100 ;
        RECT 15.380 286.950 19.330 287.100 ;
        RECT 10.130 286.500 10.730 286.950 ;
        RECT 18.730 286.500 19.330 286.950 ;
        RECT 10.130 286.350 14.080 286.500 ;
        RECT 15.380 286.350 19.330 286.500 ;
        RECT 10.130 285.900 10.730 286.350 ;
        RECT 18.730 285.900 19.330 286.350 ;
        RECT 10.130 285.750 14.080 285.900 ;
        RECT 15.380 285.750 19.330 285.900 ;
        RECT 10.130 285.300 10.730 285.750 ;
        RECT 18.730 285.300 19.330 285.750 ;
        RECT 10.130 285.150 14.080 285.300 ;
        RECT 15.380 285.150 19.330 285.300 ;
        RECT 10.130 284.700 10.730 285.150 ;
        RECT 18.730 284.700 19.330 285.150 ;
        RECT 10.130 284.550 14.080 284.700 ;
        RECT 15.380 284.550 19.330 284.700 ;
        RECT 10.130 284.100 10.730 284.550 ;
        RECT 18.730 284.100 19.330 284.550 ;
        RECT 10.130 283.950 14.080 284.100 ;
        RECT 15.380 283.950 19.330 284.100 ;
        RECT 10.130 283.500 10.730 283.950 ;
        RECT 18.730 283.500 19.330 283.950 ;
        RECT 10.130 283.350 14.080 283.500 ;
        RECT 15.380 283.350 19.330 283.500 ;
        RECT 10.130 282.900 10.730 283.350 ;
        RECT 18.730 282.900 19.330 283.350 ;
        RECT 10.130 282.750 14.080 282.900 ;
        RECT 15.380 282.750 19.330 282.900 ;
        RECT 10.130 282.300 10.730 282.750 ;
        RECT 18.730 282.300 19.330 282.750 ;
        RECT 10.130 282.150 14.080 282.300 ;
        RECT 15.380 282.150 19.330 282.300 ;
        RECT 10.130 282.000 10.730 282.150 ;
        RECT 6.530 281.700 10.730 282.000 ;
        RECT 18.730 282.000 19.330 282.150 ;
        RECT 19.780 282.000 19.930 289.550 ;
        RECT 20.380 282.000 20.530 289.550 ;
        RECT 20.980 282.000 21.130 289.550 ;
        RECT 21.580 282.000 21.730 289.550 ;
        RECT 22.180 282.000 22.330 289.550 ;
        RECT 22.780 282.000 22.930 284.900 ;
        RECT 18.730 281.700 22.930 282.000 ;
        RECT 6.530 281.550 14.080 281.700 ;
        RECT 15.380 281.550 22.930 281.700 ;
        RECT 6.530 281.350 10.730 281.550 ;
        RECT 4.730 281.050 9.130 281.200 ;
        RECT 9.280 281.050 10.730 281.350 ;
        RECT 4.730 280.150 10.730 281.050 ;
        RECT 18.730 281.350 22.930 281.550 ;
        RECT 18.730 281.050 20.180 281.350 ;
        RECT 23.530 281.200 25.930 284.400 ;
        RECT 26.530 282.000 26.680 284.900 ;
        RECT 27.130 282.000 27.280 289.550 ;
        RECT 27.730 282.000 27.880 289.550 ;
        RECT 28.330 282.000 28.480 289.550 ;
        RECT 28.930 282.000 29.080 289.550 ;
        RECT 29.530 282.000 29.680 289.550 ;
        RECT 30.130 289.350 34.080 289.550 ;
        RECT 35.380 289.350 39.330 289.550 ;
        RECT 30.130 288.900 30.730 289.350 ;
        RECT 38.730 288.900 39.330 289.350 ;
        RECT 30.130 288.750 34.080 288.900 ;
        RECT 35.380 288.750 39.330 288.900 ;
        RECT 30.130 288.300 30.730 288.750 ;
        RECT 38.730 288.300 39.330 288.750 ;
        RECT 30.130 288.150 34.080 288.300 ;
        RECT 35.380 288.150 39.330 288.300 ;
        RECT 30.130 287.700 30.730 288.150 ;
        RECT 38.730 287.700 39.330 288.150 ;
        RECT 30.130 287.550 34.080 287.700 ;
        RECT 35.380 287.550 39.330 287.700 ;
        RECT 30.130 287.100 30.730 287.550 ;
        RECT 38.730 287.100 39.330 287.550 ;
        RECT 30.130 286.950 34.080 287.100 ;
        RECT 35.380 286.950 39.330 287.100 ;
        RECT 30.130 286.500 30.730 286.950 ;
        RECT 38.730 286.500 39.330 286.950 ;
        RECT 30.130 286.350 34.080 286.500 ;
        RECT 35.380 286.350 39.330 286.500 ;
        RECT 30.130 285.900 30.730 286.350 ;
        RECT 38.730 285.900 39.330 286.350 ;
        RECT 30.130 285.750 34.080 285.900 ;
        RECT 35.380 285.750 39.330 285.900 ;
        RECT 30.130 285.300 30.730 285.750 ;
        RECT 38.730 285.300 39.330 285.750 ;
        RECT 30.130 285.150 34.080 285.300 ;
        RECT 35.380 285.150 39.330 285.300 ;
        RECT 30.130 284.700 30.730 285.150 ;
        RECT 38.730 284.700 39.330 285.150 ;
        RECT 30.130 284.550 34.080 284.700 ;
        RECT 35.380 284.550 39.330 284.700 ;
        RECT 30.130 284.100 30.730 284.550 ;
        RECT 38.730 284.100 39.330 284.550 ;
        RECT 30.130 283.950 34.080 284.100 ;
        RECT 35.380 283.950 39.330 284.100 ;
        RECT 30.130 283.500 30.730 283.950 ;
        RECT 38.730 283.500 39.330 283.950 ;
        RECT 30.130 283.350 34.080 283.500 ;
        RECT 35.380 283.350 39.330 283.500 ;
        RECT 30.130 282.900 30.730 283.350 ;
        RECT 38.730 282.900 39.330 283.350 ;
        RECT 30.130 282.750 34.080 282.900 ;
        RECT 35.380 282.750 39.330 282.900 ;
        RECT 30.130 282.300 30.730 282.750 ;
        RECT 38.730 282.300 39.330 282.750 ;
        RECT 30.130 282.150 34.080 282.300 ;
        RECT 35.380 282.150 39.330 282.300 ;
        RECT 30.130 282.000 30.730 282.150 ;
        RECT 26.530 281.700 30.730 282.000 ;
        RECT 38.730 282.000 39.330 282.150 ;
        RECT 39.780 282.000 39.930 289.550 ;
        RECT 40.380 282.000 40.530 289.550 ;
        RECT 40.980 282.000 41.130 289.550 ;
        RECT 41.580 282.000 41.730 289.550 ;
        RECT 42.180 282.000 42.330 289.550 ;
        RECT 42.780 282.000 42.930 284.900 ;
        RECT 38.730 281.700 42.930 282.000 ;
        RECT 26.530 281.550 34.080 281.700 ;
        RECT 35.380 281.550 42.930 281.700 ;
        RECT 26.530 281.350 30.730 281.550 ;
        RECT 20.330 281.050 29.130 281.200 ;
        RECT 29.280 281.050 30.730 281.350 ;
        RECT 18.730 280.150 30.730 281.050 ;
        RECT 38.730 281.350 42.930 281.550 ;
        RECT 38.730 281.050 40.180 281.350 ;
        RECT 43.530 281.200 45.930 284.400 ;
        RECT 46.530 282.000 46.680 284.900 ;
        RECT 47.130 282.000 47.280 289.550 ;
        RECT 47.730 282.000 47.880 289.550 ;
        RECT 48.330 282.000 48.480 289.550 ;
        RECT 48.930 282.000 49.080 289.550 ;
        RECT 49.530 282.000 49.680 289.550 ;
        RECT 50.130 289.350 54.080 289.550 ;
        RECT 55.380 289.350 59.330 289.550 ;
        RECT 50.130 288.900 50.730 289.350 ;
        RECT 58.730 288.900 59.330 289.350 ;
        RECT 50.130 288.750 54.080 288.900 ;
        RECT 55.380 288.750 59.330 288.900 ;
        RECT 50.130 288.300 50.730 288.750 ;
        RECT 58.730 288.300 59.330 288.750 ;
        RECT 50.130 288.150 54.080 288.300 ;
        RECT 55.380 288.150 59.330 288.300 ;
        RECT 50.130 287.700 50.730 288.150 ;
        RECT 58.730 287.700 59.330 288.150 ;
        RECT 50.130 287.550 54.080 287.700 ;
        RECT 55.380 287.550 59.330 287.700 ;
        RECT 50.130 287.100 50.730 287.550 ;
        RECT 58.730 287.100 59.330 287.550 ;
        RECT 50.130 286.950 54.080 287.100 ;
        RECT 55.380 286.950 59.330 287.100 ;
        RECT 50.130 286.500 50.730 286.950 ;
        RECT 58.730 286.500 59.330 286.950 ;
        RECT 50.130 286.350 54.080 286.500 ;
        RECT 55.380 286.350 59.330 286.500 ;
        RECT 50.130 285.900 50.730 286.350 ;
        RECT 58.730 285.900 59.330 286.350 ;
        RECT 50.130 285.750 54.080 285.900 ;
        RECT 55.380 285.750 59.330 285.900 ;
        RECT 50.130 285.300 50.730 285.750 ;
        RECT 58.730 285.300 59.330 285.750 ;
        RECT 50.130 285.150 54.080 285.300 ;
        RECT 55.380 285.150 59.330 285.300 ;
        RECT 50.130 284.700 50.730 285.150 ;
        RECT 58.730 284.700 59.330 285.150 ;
        RECT 50.130 284.550 54.080 284.700 ;
        RECT 55.380 284.550 59.330 284.700 ;
        RECT 50.130 284.100 50.730 284.550 ;
        RECT 58.730 284.100 59.330 284.550 ;
        RECT 50.130 283.950 54.080 284.100 ;
        RECT 55.380 283.950 59.330 284.100 ;
        RECT 50.130 283.500 50.730 283.950 ;
        RECT 58.730 283.500 59.330 283.950 ;
        RECT 50.130 283.350 54.080 283.500 ;
        RECT 55.380 283.350 59.330 283.500 ;
        RECT 50.130 282.900 50.730 283.350 ;
        RECT 58.730 282.900 59.330 283.350 ;
        RECT 50.130 282.750 54.080 282.900 ;
        RECT 55.380 282.750 59.330 282.900 ;
        RECT 50.130 282.300 50.730 282.750 ;
        RECT 58.730 282.300 59.330 282.750 ;
        RECT 50.130 282.150 54.080 282.300 ;
        RECT 55.380 282.150 59.330 282.300 ;
        RECT 50.130 282.000 50.730 282.150 ;
        RECT 46.530 281.700 50.730 282.000 ;
        RECT 58.730 282.000 59.330 282.150 ;
        RECT 59.780 282.000 59.930 289.550 ;
        RECT 60.380 282.000 60.530 289.550 ;
        RECT 60.980 282.000 61.130 289.550 ;
        RECT 61.580 282.000 61.730 289.550 ;
        RECT 62.180 282.000 62.330 289.550 ;
        RECT 62.780 282.000 62.930 284.900 ;
        RECT 58.730 281.700 62.930 282.000 ;
        RECT 46.530 281.550 54.080 281.700 ;
        RECT 55.380 281.550 62.930 281.700 ;
        RECT 46.530 281.350 50.730 281.550 ;
        RECT 40.330 281.050 49.130 281.200 ;
        RECT 49.280 281.050 50.730 281.350 ;
        RECT 38.730 280.150 50.730 281.050 ;
        RECT 58.730 281.350 62.930 281.550 ;
        RECT 58.730 281.050 60.180 281.350 ;
        RECT 63.530 281.200 65.930 284.400 ;
        RECT 66.530 282.000 66.680 284.900 ;
        RECT 67.130 282.000 67.280 289.550 ;
        RECT 67.730 282.000 67.880 289.550 ;
        RECT 68.330 282.000 68.480 289.550 ;
        RECT 68.930 282.000 69.080 289.550 ;
        RECT 69.530 282.000 69.680 289.550 ;
        RECT 70.130 289.350 74.080 289.550 ;
        RECT 75.380 289.350 79.330 289.550 ;
        RECT 70.130 288.900 70.730 289.350 ;
        RECT 78.730 288.900 79.330 289.350 ;
        RECT 70.130 288.750 74.080 288.900 ;
        RECT 75.380 288.750 79.330 288.900 ;
        RECT 70.130 288.300 70.730 288.750 ;
        RECT 78.730 288.300 79.330 288.750 ;
        RECT 70.130 288.150 74.080 288.300 ;
        RECT 75.380 288.150 79.330 288.300 ;
        RECT 70.130 287.700 70.730 288.150 ;
        RECT 78.730 287.700 79.330 288.150 ;
        RECT 70.130 287.550 74.080 287.700 ;
        RECT 75.380 287.550 79.330 287.700 ;
        RECT 70.130 287.100 70.730 287.550 ;
        RECT 78.730 287.100 79.330 287.550 ;
        RECT 70.130 286.950 74.080 287.100 ;
        RECT 75.380 286.950 79.330 287.100 ;
        RECT 70.130 286.500 70.730 286.950 ;
        RECT 78.730 286.500 79.330 286.950 ;
        RECT 70.130 286.350 74.080 286.500 ;
        RECT 75.380 286.350 79.330 286.500 ;
        RECT 70.130 285.900 70.730 286.350 ;
        RECT 78.730 285.900 79.330 286.350 ;
        RECT 70.130 285.750 74.080 285.900 ;
        RECT 75.380 285.750 79.330 285.900 ;
        RECT 70.130 285.300 70.730 285.750 ;
        RECT 78.730 285.300 79.330 285.750 ;
        RECT 70.130 285.150 74.080 285.300 ;
        RECT 75.380 285.150 79.330 285.300 ;
        RECT 70.130 284.700 70.730 285.150 ;
        RECT 78.730 284.700 79.330 285.150 ;
        RECT 70.130 284.550 74.080 284.700 ;
        RECT 75.380 284.550 79.330 284.700 ;
        RECT 70.130 284.100 70.730 284.550 ;
        RECT 78.730 284.100 79.330 284.550 ;
        RECT 70.130 283.950 74.080 284.100 ;
        RECT 75.380 283.950 79.330 284.100 ;
        RECT 70.130 283.500 70.730 283.950 ;
        RECT 78.730 283.500 79.330 283.950 ;
        RECT 70.130 283.350 74.080 283.500 ;
        RECT 75.380 283.350 79.330 283.500 ;
        RECT 70.130 282.900 70.730 283.350 ;
        RECT 78.730 282.900 79.330 283.350 ;
        RECT 70.130 282.750 74.080 282.900 ;
        RECT 75.380 282.750 79.330 282.900 ;
        RECT 70.130 282.300 70.730 282.750 ;
        RECT 78.730 282.300 79.330 282.750 ;
        RECT 70.130 282.150 74.080 282.300 ;
        RECT 75.380 282.150 79.330 282.300 ;
        RECT 70.130 282.000 70.730 282.150 ;
        RECT 66.530 281.700 70.730 282.000 ;
        RECT 78.730 282.000 79.330 282.150 ;
        RECT 79.780 282.000 79.930 289.550 ;
        RECT 80.380 282.000 80.530 289.550 ;
        RECT 80.980 282.000 81.130 289.550 ;
        RECT 81.580 282.000 81.730 289.550 ;
        RECT 82.180 282.000 82.330 289.550 ;
        RECT 82.780 282.000 82.930 284.900 ;
        RECT 78.730 281.700 82.930 282.000 ;
        RECT 66.530 281.550 74.080 281.700 ;
        RECT 75.380 281.550 82.930 281.700 ;
        RECT 66.530 281.350 70.730 281.550 ;
        RECT 60.330 281.050 69.130 281.200 ;
        RECT 69.280 281.050 70.730 281.350 ;
        RECT 58.730 280.150 70.730 281.050 ;
        RECT 78.730 281.350 82.930 281.550 ;
        RECT 78.730 281.050 80.180 281.350 ;
        RECT 83.530 281.200 85.930 284.400 ;
        RECT 86.530 282.000 86.680 284.900 ;
        RECT 87.130 282.000 87.280 289.550 ;
        RECT 87.730 282.000 87.880 289.550 ;
        RECT 88.330 282.000 88.480 289.550 ;
        RECT 88.930 282.000 89.080 289.550 ;
        RECT 89.530 282.000 89.680 289.550 ;
        RECT 90.130 289.350 94.080 289.550 ;
        RECT 95.380 289.350 99.330 289.550 ;
        RECT 90.130 288.900 90.730 289.350 ;
        RECT 98.730 288.900 99.330 289.350 ;
        RECT 90.130 288.750 94.080 288.900 ;
        RECT 95.380 288.750 99.330 288.900 ;
        RECT 90.130 288.300 90.730 288.750 ;
        RECT 98.730 288.300 99.330 288.750 ;
        RECT 90.130 288.150 94.080 288.300 ;
        RECT 95.380 288.150 99.330 288.300 ;
        RECT 90.130 287.700 90.730 288.150 ;
        RECT 98.730 287.700 99.330 288.150 ;
        RECT 90.130 287.550 94.080 287.700 ;
        RECT 95.380 287.550 99.330 287.700 ;
        RECT 90.130 287.100 90.730 287.550 ;
        RECT 98.730 287.100 99.330 287.550 ;
        RECT 90.130 286.950 94.080 287.100 ;
        RECT 95.380 286.950 99.330 287.100 ;
        RECT 90.130 286.500 90.730 286.950 ;
        RECT 98.730 286.500 99.330 286.950 ;
        RECT 90.130 286.350 94.080 286.500 ;
        RECT 95.380 286.350 99.330 286.500 ;
        RECT 90.130 285.900 90.730 286.350 ;
        RECT 98.730 285.900 99.330 286.350 ;
        RECT 90.130 285.750 94.080 285.900 ;
        RECT 95.380 285.750 99.330 285.900 ;
        RECT 90.130 285.300 90.730 285.750 ;
        RECT 98.730 285.300 99.330 285.750 ;
        RECT 90.130 285.150 94.080 285.300 ;
        RECT 95.380 285.150 99.330 285.300 ;
        RECT 90.130 284.700 90.730 285.150 ;
        RECT 98.730 284.700 99.330 285.150 ;
        RECT 90.130 284.550 94.080 284.700 ;
        RECT 95.380 284.550 99.330 284.700 ;
        RECT 90.130 284.100 90.730 284.550 ;
        RECT 98.730 284.100 99.330 284.550 ;
        RECT 90.130 283.950 94.080 284.100 ;
        RECT 95.380 283.950 99.330 284.100 ;
        RECT 90.130 283.500 90.730 283.950 ;
        RECT 98.730 283.500 99.330 283.950 ;
        RECT 90.130 283.350 94.080 283.500 ;
        RECT 95.380 283.350 99.330 283.500 ;
        RECT 90.130 282.900 90.730 283.350 ;
        RECT 98.730 282.900 99.330 283.350 ;
        RECT 90.130 282.750 94.080 282.900 ;
        RECT 95.380 282.750 99.330 282.900 ;
        RECT 90.130 282.300 90.730 282.750 ;
        RECT 98.730 282.300 99.330 282.750 ;
        RECT 90.130 282.150 94.080 282.300 ;
        RECT 95.380 282.150 99.330 282.300 ;
        RECT 90.130 282.000 90.730 282.150 ;
        RECT 86.530 281.700 90.730 282.000 ;
        RECT 98.730 282.000 99.330 282.150 ;
        RECT 99.780 282.000 99.930 289.550 ;
        RECT 100.380 282.000 100.530 289.550 ;
        RECT 100.980 282.000 101.130 289.550 ;
        RECT 101.580 282.000 101.730 289.550 ;
        RECT 102.180 282.000 102.330 289.550 ;
        RECT 102.780 282.000 102.930 284.900 ;
        RECT 98.730 281.700 102.930 282.000 ;
        RECT 86.530 281.550 94.080 281.700 ;
        RECT 95.380 281.550 102.930 281.700 ;
        RECT 86.530 281.350 90.730 281.550 ;
        RECT 80.330 281.050 89.130 281.200 ;
        RECT 89.280 281.050 90.730 281.350 ;
        RECT 78.730 280.150 90.730 281.050 ;
        RECT 98.730 281.350 102.930 281.550 ;
        RECT 103.530 283.275 104.730 284.400 ;
        RECT 103.530 282.000 107.140 283.275 ;
        RECT 98.730 281.050 100.180 281.350 ;
        RECT 103.530 281.200 104.730 282.000 ;
        RECT 100.330 281.050 104.730 281.200 ;
        RECT 98.730 280.150 104.730 281.050 ;
        RECT 4.730 279.850 9.130 280.150 ;
        RECT 20.330 279.850 29.130 280.150 ;
        RECT 40.330 279.850 49.130 280.150 ;
        RECT 60.330 279.850 69.130 280.150 ;
        RECT 80.330 279.850 89.130 280.150 ;
        RECT 4.730 278.950 10.730 279.850 ;
        RECT 20.330 279.800 30.730 279.850 ;
        RECT 40.330 279.800 50.730 279.850 ;
        RECT 60.330 279.800 70.730 279.850 ;
        RECT 80.330 279.800 90.730 279.850 ;
        RECT 100.330 279.800 104.730 280.150 ;
        RECT 4.730 278.800 9.130 278.950 ;
        RECT 4.730 277.610 5.930 278.800 ;
        RECT 9.280 278.650 10.730 278.950 ;
        RECT 2.315 276.335 5.930 277.610 ;
        RECT 4.730 275.600 5.930 276.335 ;
        RECT 6.530 278.450 10.730 278.650 ;
        RECT 18.730 278.950 30.730 279.800 ;
        RECT 18.730 278.900 29.130 278.950 ;
        RECT 18.730 278.650 20.180 278.900 ;
        RECT 20.330 278.800 29.130 278.900 ;
        RECT 18.730 278.450 22.930 278.650 ;
        RECT 6.530 278.300 14.080 278.450 ;
        RECT 15.430 278.300 22.930 278.450 ;
        RECT 6.530 278.000 10.730 278.300 ;
        RECT 2.315 273.250 4.315 275.545 ;
        RECT 6.530 275.150 6.680 278.000 ;
        RECT 7.130 270.450 7.280 278.000 ;
        RECT 7.730 270.450 7.880 278.000 ;
        RECT 8.330 270.450 8.480 278.000 ;
        RECT 8.930 270.450 9.080 278.000 ;
        RECT 9.530 270.450 9.680 278.000 ;
        RECT 10.130 277.850 10.730 278.000 ;
        RECT 18.730 278.000 22.930 278.300 ;
        RECT 18.730 277.850 19.330 278.000 ;
        RECT 10.130 277.700 14.080 277.850 ;
        RECT 15.380 277.700 19.330 277.850 ;
        RECT 10.130 277.250 10.730 277.700 ;
        RECT 18.730 277.250 19.330 277.700 ;
        RECT 10.130 277.100 14.080 277.250 ;
        RECT 15.380 277.100 19.330 277.250 ;
        RECT 10.130 276.650 10.730 277.100 ;
        RECT 18.730 276.650 19.330 277.100 ;
        RECT 10.130 276.500 14.080 276.650 ;
        RECT 15.380 276.500 19.330 276.650 ;
        RECT 10.130 276.050 10.730 276.500 ;
        RECT 18.730 276.050 19.330 276.500 ;
        RECT 10.130 275.900 14.080 276.050 ;
        RECT 15.380 275.900 19.330 276.050 ;
        RECT 10.130 275.450 10.730 275.900 ;
        RECT 18.730 275.450 19.330 275.900 ;
        RECT 10.130 275.300 14.080 275.450 ;
        RECT 15.380 275.300 19.330 275.450 ;
        RECT 10.130 274.850 10.730 275.300 ;
        RECT 18.730 274.850 19.330 275.300 ;
        RECT 10.130 274.700 14.080 274.850 ;
        RECT 15.380 274.700 19.330 274.850 ;
        RECT 10.130 274.250 10.730 274.700 ;
        RECT 18.730 274.250 19.330 274.700 ;
        RECT 10.130 274.100 14.080 274.250 ;
        RECT 15.380 274.100 19.330 274.250 ;
        RECT 10.130 273.650 10.730 274.100 ;
        RECT 18.730 273.650 19.330 274.100 ;
        RECT 10.130 273.500 14.080 273.650 ;
        RECT 15.380 273.500 19.330 273.650 ;
        RECT 10.130 273.050 10.730 273.500 ;
        RECT 18.730 273.050 19.330 273.500 ;
        RECT 10.130 272.900 14.080 273.050 ;
        RECT 15.380 272.900 19.330 273.050 ;
        RECT 10.130 272.450 10.730 272.900 ;
        RECT 18.730 272.450 19.330 272.900 ;
        RECT 10.130 272.300 14.080 272.450 ;
        RECT 15.380 272.300 19.330 272.450 ;
        RECT 10.130 271.850 10.730 272.300 ;
        RECT 18.730 271.850 19.330 272.300 ;
        RECT 10.130 271.700 14.080 271.850 ;
        RECT 15.380 271.700 19.330 271.850 ;
        RECT 10.130 271.250 10.730 271.700 ;
        RECT 18.730 271.250 19.330 271.700 ;
        RECT 10.130 271.100 14.080 271.250 ;
        RECT 15.380 271.100 19.330 271.250 ;
        RECT 10.130 270.650 10.730 271.100 ;
        RECT 18.730 270.650 19.330 271.100 ;
        RECT 10.130 270.450 14.080 270.650 ;
        RECT 15.380 270.450 19.330 270.650 ;
        RECT 19.780 270.450 19.930 278.000 ;
        RECT 20.380 270.450 20.530 278.000 ;
        RECT 20.980 270.450 21.130 278.000 ;
        RECT 21.580 270.450 21.730 278.000 ;
        RECT 22.180 270.450 22.330 278.000 ;
        RECT 22.780 275.150 22.930 278.000 ;
        RECT 23.530 275.600 25.930 278.800 ;
        RECT 29.280 278.650 30.730 278.950 ;
        RECT 26.530 278.450 30.730 278.650 ;
        RECT 38.730 278.950 50.730 279.800 ;
        RECT 38.730 278.900 49.130 278.950 ;
        RECT 38.730 278.650 40.180 278.900 ;
        RECT 40.330 278.800 49.130 278.900 ;
        RECT 38.730 278.450 42.930 278.650 ;
        RECT 26.530 278.300 34.080 278.450 ;
        RECT 35.430 278.300 42.930 278.450 ;
        RECT 26.530 278.000 30.730 278.300 ;
        RECT 26.530 275.150 26.680 278.000 ;
        RECT 27.130 270.450 27.280 278.000 ;
        RECT 27.730 270.450 27.880 278.000 ;
        RECT 28.330 270.450 28.480 278.000 ;
        RECT 28.930 270.450 29.080 278.000 ;
        RECT 29.530 270.450 29.680 278.000 ;
        RECT 30.130 277.850 30.730 278.000 ;
        RECT 38.730 278.000 42.930 278.300 ;
        RECT 38.730 277.850 39.330 278.000 ;
        RECT 30.130 277.700 34.080 277.850 ;
        RECT 35.380 277.700 39.330 277.850 ;
        RECT 30.130 277.250 30.730 277.700 ;
        RECT 38.730 277.250 39.330 277.700 ;
        RECT 30.130 277.100 34.080 277.250 ;
        RECT 35.380 277.100 39.330 277.250 ;
        RECT 30.130 276.650 30.730 277.100 ;
        RECT 38.730 276.650 39.330 277.100 ;
        RECT 30.130 276.500 34.080 276.650 ;
        RECT 35.380 276.500 39.330 276.650 ;
        RECT 30.130 276.050 30.730 276.500 ;
        RECT 38.730 276.050 39.330 276.500 ;
        RECT 30.130 275.900 34.080 276.050 ;
        RECT 35.380 275.900 39.330 276.050 ;
        RECT 30.130 275.450 30.730 275.900 ;
        RECT 38.730 275.450 39.330 275.900 ;
        RECT 30.130 275.300 34.080 275.450 ;
        RECT 35.380 275.300 39.330 275.450 ;
        RECT 30.130 274.850 30.730 275.300 ;
        RECT 38.730 274.850 39.330 275.300 ;
        RECT 30.130 274.700 34.080 274.850 ;
        RECT 35.380 274.700 39.330 274.850 ;
        RECT 30.130 274.250 30.730 274.700 ;
        RECT 38.730 274.250 39.330 274.700 ;
        RECT 30.130 274.100 34.080 274.250 ;
        RECT 35.380 274.100 39.330 274.250 ;
        RECT 30.130 273.650 30.730 274.100 ;
        RECT 38.730 273.650 39.330 274.100 ;
        RECT 30.130 273.500 34.080 273.650 ;
        RECT 35.380 273.500 39.330 273.650 ;
        RECT 30.130 273.050 30.730 273.500 ;
        RECT 38.730 273.050 39.330 273.500 ;
        RECT 30.130 272.900 34.080 273.050 ;
        RECT 35.380 272.900 39.330 273.050 ;
        RECT 30.130 272.450 30.730 272.900 ;
        RECT 38.730 272.450 39.330 272.900 ;
        RECT 30.130 272.300 34.080 272.450 ;
        RECT 35.380 272.300 39.330 272.450 ;
        RECT 30.130 271.850 30.730 272.300 ;
        RECT 38.730 271.850 39.330 272.300 ;
        RECT 30.130 271.700 34.080 271.850 ;
        RECT 35.380 271.700 39.330 271.850 ;
        RECT 30.130 271.250 30.730 271.700 ;
        RECT 38.730 271.250 39.330 271.700 ;
        RECT 30.130 271.100 34.080 271.250 ;
        RECT 35.380 271.100 39.330 271.250 ;
        RECT 30.130 270.650 30.730 271.100 ;
        RECT 38.730 270.650 39.330 271.100 ;
        RECT 30.130 270.450 34.080 270.650 ;
        RECT 35.380 270.450 39.330 270.650 ;
        RECT 39.780 270.450 39.930 278.000 ;
        RECT 40.380 270.450 40.530 278.000 ;
        RECT 40.980 270.450 41.130 278.000 ;
        RECT 41.580 270.450 41.730 278.000 ;
        RECT 42.180 270.450 42.330 278.000 ;
        RECT 42.780 275.150 42.930 278.000 ;
        RECT 43.530 275.600 45.930 278.800 ;
        RECT 49.280 278.650 50.730 278.950 ;
        RECT 46.530 278.450 50.730 278.650 ;
        RECT 58.730 278.950 70.730 279.800 ;
        RECT 58.730 278.900 69.130 278.950 ;
        RECT 58.730 278.650 60.180 278.900 ;
        RECT 60.330 278.800 69.130 278.900 ;
        RECT 58.730 278.450 62.930 278.650 ;
        RECT 46.530 278.300 54.080 278.450 ;
        RECT 55.430 278.300 62.930 278.450 ;
        RECT 46.530 278.000 50.730 278.300 ;
        RECT 46.530 275.150 46.680 278.000 ;
        RECT 47.130 270.450 47.280 278.000 ;
        RECT 47.730 270.450 47.880 278.000 ;
        RECT 48.330 270.450 48.480 278.000 ;
        RECT 48.930 270.450 49.080 278.000 ;
        RECT 49.530 270.450 49.680 278.000 ;
        RECT 50.130 277.850 50.730 278.000 ;
        RECT 58.730 278.000 62.930 278.300 ;
        RECT 58.730 277.850 59.330 278.000 ;
        RECT 50.130 277.700 54.080 277.850 ;
        RECT 55.380 277.700 59.330 277.850 ;
        RECT 50.130 277.250 50.730 277.700 ;
        RECT 58.730 277.250 59.330 277.700 ;
        RECT 50.130 277.100 54.080 277.250 ;
        RECT 55.380 277.100 59.330 277.250 ;
        RECT 50.130 276.650 50.730 277.100 ;
        RECT 58.730 276.650 59.330 277.100 ;
        RECT 50.130 276.500 54.080 276.650 ;
        RECT 55.380 276.500 59.330 276.650 ;
        RECT 50.130 276.050 50.730 276.500 ;
        RECT 58.730 276.050 59.330 276.500 ;
        RECT 50.130 275.900 54.080 276.050 ;
        RECT 55.380 275.900 59.330 276.050 ;
        RECT 50.130 275.450 50.730 275.900 ;
        RECT 58.730 275.450 59.330 275.900 ;
        RECT 50.130 275.300 54.080 275.450 ;
        RECT 55.380 275.300 59.330 275.450 ;
        RECT 50.130 274.850 50.730 275.300 ;
        RECT 58.730 274.850 59.330 275.300 ;
        RECT 50.130 274.700 54.080 274.850 ;
        RECT 55.380 274.700 59.330 274.850 ;
        RECT 50.130 274.250 50.730 274.700 ;
        RECT 58.730 274.250 59.330 274.700 ;
        RECT 50.130 274.100 54.080 274.250 ;
        RECT 55.380 274.100 59.330 274.250 ;
        RECT 50.130 273.650 50.730 274.100 ;
        RECT 58.730 273.650 59.330 274.100 ;
        RECT 50.130 273.500 54.080 273.650 ;
        RECT 55.380 273.500 59.330 273.650 ;
        RECT 50.130 273.050 50.730 273.500 ;
        RECT 58.730 273.050 59.330 273.500 ;
        RECT 50.130 272.900 54.080 273.050 ;
        RECT 55.380 272.900 59.330 273.050 ;
        RECT 50.130 272.450 50.730 272.900 ;
        RECT 58.730 272.450 59.330 272.900 ;
        RECT 50.130 272.300 54.080 272.450 ;
        RECT 55.380 272.300 59.330 272.450 ;
        RECT 50.130 271.850 50.730 272.300 ;
        RECT 58.730 271.850 59.330 272.300 ;
        RECT 50.130 271.700 54.080 271.850 ;
        RECT 55.380 271.700 59.330 271.850 ;
        RECT 50.130 271.250 50.730 271.700 ;
        RECT 58.730 271.250 59.330 271.700 ;
        RECT 50.130 271.100 54.080 271.250 ;
        RECT 55.380 271.100 59.330 271.250 ;
        RECT 50.130 270.650 50.730 271.100 ;
        RECT 58.730 270.650 59.330 271.100 ;
        RECT 50.130 270.450 54.080 270.650 ;
        RECT 55.380 270.450 59.330 270.650 ;
        RECT 59.780 270.450 59.930 278.000 ;
        RECT 60.380 270.450 60.530 278.000 ;
        RECT 60.980 270.450 61.130 278.000 ;
        RECT 61.580 270.450 61.730 278.000 ;
        RECT 62.180 270.450 62.330 278.000 ;
        RECT 62.780 275.150 62.930 278.000 ;
        RECT 63.530 275.600 65.930 278.800 ;
        RECT 69.280 278.650 70.730 278.950 ;
        RECT 66.530 278.450 70.730 278.650 ;
        RECT 78.730 278.950 90.730 279.800 ;
        RECT 78.730 278.900 89.130 278.950 ;
        RECT 78.730 278.650 80.180 278.900 ;
        RECT 80.330 278.800 89.130 278.900 ;
        RECT 78.730 278.450 82.930 278.650 ;
        RECT 66.530 278.300 74.080 278.450 ;
        RECT 75.430 278.300 82.930 278.450 ;
        RECT 66.530 278.000 70.730 278.300 ;
        RECT 66.530 275.150 66.680 278.000 ;
        RECT 67.130 270.450 67.280 278.000 ;
        RECT 67.730 270.450 67.880 278.000 ;
        RECT 68.330 270.450 68.480 278.000 ;
        RECT 68.930 270.450 69.080 278.000 ;
        RECT 69.530 270.450 69.680 278.000 ;
        RECT 70.130 277.850 70.730 278.000 ;
        RECT 78.730 278.000 82.930 278.300 ;
        RECT 78.730 277.850 79.330 278.000 ;
        RECT 70.130 277.700 74.080 277.850 ;
        RECT 75.380 277.700 79.330 277.850 ;
        RECT 70.130 277.250 70.730 277.700 ;
        RECT 78.730 277.250 79.330 277.700 ;
        RECT 70.130 277.100 74.080 277.250 ;
        RECT 75.380 277.100 79.330 277.250 ;
        RECT 70.130 276.650 70.730 277.100 ;
        RECT 78.730 276.650 79.330 277.100 ;
        RECT 70.130 276.500 74.080 276.650 ;
        RECT 75.380 276.500 79.330 276.650 ;
        RECT 70.130 276.050 70.730 276.500 ;
        RECT 78.730 276.050 79.330 276.500 ;
        RECT 70.130 275.900 74.080 276.050 ;
        RECT 75.380 275.900 79.330 276.050 ;
        RECT 70.130 275.450 70.730 275.900 ;
        RECT 78.730 275.450 79.330 275.900 ;
        RECT 70.130 275.300 74.080 275.450 ;
        RECT 75.380 275.300 79.330 275.450 ;
        RECT 70.130 274.850 70.730 275.300 ;
        RECT 78.730 274.850 79.330 275.300 ;
        RECT 70.130 274.700 74.080 274.850 ;
        RECT 75.380 274.700 79.330 274.850 ;
        RECT 70.130 274.250 70.730 274.700 ;
        RECT 78.730 274.250 79.330 274.700 ;
        RECT 70.130 274.100 74.080 274.250 ;
        RECT 75.380 274.100 79.330 274.250 ;
        RECT 70.130 273.650 70.730 274.100 ;
        RECT 78.730 273.650 79.330 274.100 ;
        RECT 70.130 273.500 74.080 273.650 ;
        RECT 75.380 273.500 79.330 273.650 ;
        RECT 70.130 273.050 70.730 273.500 ;
        RECT 78.730 273.050 79.330 273.500 ;
        RECT 70.130 272.900 74.080 273.050 ;
        RECT 75.380 272.900 79.330 273.050 ;
        RECT 70.130 272.450 70.730 272.900 ;
        RECT 78.730 272.450 79.330 272.900 ;
        RECT 70.130 272.300 74.080 272.450 ;
        RECT 75.380 272.300 79.330 272.450 ;
        RECT 70.130 271.850 70.730 272.300 ;
        RECT 78.730 271.850 79.330 272.300 ;
        RECT 70.130 271.700 74.080 271.850 ;
        RECT 75.380 271.700 79.330 271.850 ;
        RECT 70.130 271.250 70.730 271.700 ;
        RECT 78.730 271.250 79.330 271.700 ;
        RECT 70.130 271.100 74.080 271.250 ;
        RECT 75.380 271.100 79.330 271.250 ;
        RECT 70.130 270.650 70.730 271.100 ;
        RECT 78.730 270.650 79.330 271.100 ;
        RECT 70.130 270.450 74.080 270.650 ;
        RECT 75.380 270.450 79.330 270.650 ;
        RECT 79.780 270.450 79.930 278.000 ;
        RECT 80.380 270.450 80.530 278.000 ;
        RECT 80.980 270.450 81.130 278.000 ;
        RECT 81.580 270.450 81.730 278.000 ;
        RECT 82.180 270.450 82.330 278.000 ;
        RECT 82.780 275.150 82.930 278.000 ;
        RECT 83.530 275.600 85.930 278.800 ;
        RECT 89.280 278.650 90.730 278.950 ;
        RECT 86.530 278.450 90.730 278.650 ;
        RECT 98.730 278.900 104.730 279.800 ;
        RECT 98.730 278.650 100.180 278.900 ;
        RECT 100.330 278.800 104.730 278.900 ;
        RECT 98.730 278.450 102.930 278.650 ;
        RECT 86.530 278.300 94.080 278.450 ;
        RECT 95.430 278.300 102.930 278.450 ;
        RECT 86.530 278.000 90.730 278.300 ;
        RECT 86.530 275.150 86.680 278.000 ;
        RECT 87.130 270.450 87.280 278.000 ;
        RECT 87.730 270.450 87.880 278.000 ;
        RECT 88.330 270.450 88.480 278.000 ;
        RECT 88.930 270.450 89.080 278.000 ;
        RECT 89.530 270.450 89.680 278.000 ;
        RECT 90.130 277.850 90.730 278.000 ;
        RECT 98.730 278.000 102.930 278.300 ;
        RECT 98.730 277.850 99.330 278.000 ;
        RECT 90.130 277.700 94.080 277.850 ;
        RECT 95.380 277.700 99.330 277.850 ;
        RECT 90.130 277.250 90.730 277.700 ;
        RECT 98.730 277.250 99.330 277.700 ;
        RECT 90.130 277.100 94.080 277.250 ;
        RECT 95.380 277.100 99.330 277.250 ;
        RECT 90.130 276.650 90.730 277.100 ;
        RECT 98.730 276.650 99.330 277.100 ;
        RECT 90.130 276.500 94.080 276.650 ;
        RECT 95.380 276.500 99.330 276.650 ;
        RECT 90.130 276.050 90.730 276.500 ;
        RECT 98.730 276.050 99.330 276.500 ;
        RECT 90.130 275.900 94.080 276.050 ;
        RECT 95.380 275.900 99.330 276.050 ;
        RECT 90.130 275.450 90.730 275.900 ;
        RECT 98.730 275.450 99.330 275.900 ;
        RECT 90.130 275.300 94.080 275.450 ;
        RECT 95.380 275.300 99.330 275.450 ;
        RECT 90.130 274.850 90.730 275.300 ;
        RECT 98.730 274.850 99.330 275.300 ;
        RECT 90.130 274.700 94.080 274.850 ;
        RECT 95.380 274.700 99.330 274.850 ;
        RECT 90.130 274.250 90.730 274.700 ;
        RECT 98.730 274.250 99.330 274.700 ;
        RECT 90.130 274.100 94.080 274.250 ;
        RECT 95.380 274.100 99.330 274.250 ;
        RECT 90.130 273.650 90.730 274.100 ;
        RECT 98.730 273.650 99.330 274.100 ;
        RECT 90.130 273.500 94.080 273.650 ;
        RECT 95.380 273.500 99.330 273.650 ;
        RECT 90.130 273.050 90.730 273.500 ;
        RECT 98.730 273.050 99.330 273.500 ;
        RECT 90.130 272.900 94.080 273.050 ;
        RECT 95.380 272.900 99.330 273.050 ;
        RECT 90.130 272.450 90.730 272.900 ;
        RECT 98.730 272.450 99.330 272.900 ;
        RECT 90.130 272.300 94.080 272.450 ;
        RECT 95.380 272.300 99.330 272.450 ;
        RECT 90.130 271.850 90.730 272.300 ;
        RECT 98.730 271.850 99.330 272.300 ;
        RECT 90.130 271.700 94.080 271.850 ;
        RECT 95.380 271.700 99.330 271.850 ;
        RECT 90.130 271.250 90.730 271.700 ;
        RECT 98.730 271.250 99.330 271.700 ;
        RECT 90.130 271.100 94.080 271.250 ;
        RECT 95.380 271.100 99.330 271.250 ;
        RECT 90.130 270.650 90.730 271.100 ;
        RECT 98.730 270.650 99.330 271.100 ;
        RECT 90.130 270.450 94.080 270.650 ;
        RECT 95.380 270.450 99.330 270.650 ;
        RECT 99.780 270.450 99.930 278.000 ;
        RECT 100.380 270.450 100.530 278.000 ;
        RECT 100.980 270.450 101.130 278.000 ;
        RECT 101.580 270.450 101.730 278.000 ;
        RECT 102.180 270.450 102.330 278.000 ;
        RECT 102.780 275.150 102.930 278.000 ;
        RECT 103.530 277.360 104.730 278.800 ;
        RECT 103.530 276.085 107.135 277.360 ;
        RECT 103.530 275.600 104.730 276.085 ;
        RECT 2.315 264.455 4.315 266.750 ;
        RECT 4.730 263.780 5.930 264.400 ;
        RECT 2.315 262.505 5.930 263.780 ;
        RECT 4.730 261.200 5.930 262.505 ;
        RECT 6.530 262.000 6.680 264.900 ;
        RECT 7.130 262.000 7.280 269.550 ;
        RECT 7.730 262.000 7.880 269.550 ;
        RECT 8.330 262.000 8.480 269.550 ;
        RECT 8.930 262.000 9.080 269.550 ;
        RECT 9.530 262.000 9.680 269.550 ;
        RECT 10.130 269.350 14.080 269.550 ;
        RECT 15.380 269.350 19.330 269.550 ;
        RECT 10.130 268.900 10.730 269.350 ;
        RECT 18.730 268.900 19.330 269.350 ;
        RECT 10.130 268.750 14.080 268.900 ;
        RECT 15.380 268.750 19.330 268.900 ;
        RECT 10.130 268.300 10.730 268.750 ;
        RECT 18.730 268.300 19.330 268.750 ;
        RECT 10.130 268.150 14.080 268.300 ;
        RECT 15.380 268.150 19.330 268.300 ;
        RECT 10.130 267.700 10.730 268.150 ;
        RECT 18.730 267.700 19.330 268.150 ;
        RECT 10.130 267.550 14.080 267.700 ;
        RECT 15.380 267.550 19.330 267.700 ;
        RECT 10.130 267.100 10.730 267.550 ;
        RECT 18.730 267.100 19.330 267.550 ;
        RECT 10.130 266.950 14.080 267.100 ;
        RECT 15.380 266.950 19.330 267.100 ;
        RECT 10.130 266.500 10.730 266.950 ;
        RECT 18.730 266.500 19.330 266.950 ;
        RECT 10.130 266.350 14.080 266.500 ;
        RECT 15.380 266.350 19.330 266.500 ;
        RECT 10.130 265.900 10.730 266.350 ;
        RECT 18.730 265.900 19.330 266.350 ;
        RECT 10.130 265.750 14.080 265.900 ;
        RECT 15.380 265.750 19.330 265.900 ;
        RECT 10.130 265.300 10.730 265.750 ;
        RECT 18.730 265.300 19.330 265.750 ;
        RECT 10.130 265.150 14.080 265.300 ;
        RECT 15.380 265.150 19.330 265.300 ;
        RECT 10.130 264.700 10.730 265.150 ;
        RECT 18.730 264.700 19.330 265.150 ;
        RECT 10.130 264.550 14.080 264.700 ;
        RECT 15.380 264.550 19.330 264.700 ;
        RECT 10.130 264.100 10.730 264.550 ;
        RECT 18.730 264.100 19.330 264.550 ;
        RECT 10.130 263.950 14.080 264.100 ;
        RECT 15.380 263.950 19.330 264.100 ;
        RECT 10.130 263.500 10.730 263.950 ;
        RECT 18.730 263.500 19.330 263.950 ;
        RECT 10.130 263.350 14.080 263.500 ;
        RECT 15.380 263.350 19.330 263.500 ;
        RECT 10.130 262.900 10.730 263.350 ;
        RECT 18.730 262.900 19.330 263.350 ;
        RECT 10.130 262.750 14.080 262.900 ;
        RECT 15.380 262.750 19.330 262.900 ;
        RECT 10.130 262.300 10.730 262.750 ;
        RECT 18.730 262.300 19.330 262.750 ;
        RECT 10.130 262.150 14.080 262.300 ;
        RECT 15.380 262.150 19.330 262.300 ;
        RECT 10.130 262.000 10.730 262.150 ;
        RECT 6.530 261.700 10.730 262.000 ;
        RECT 18.730 262.000 19.330 262.150 ;
        RECT 19.780 262.000 19.930 269.550 ;
        RECT 20.380 262.000 20.530 269.550 ;
        RECT 20.980 262.000 21.130 269.550 ;
        RECT 21.580 262.000 21.730 269.550 ;
        RECT 22.180 262.000 22.330 269.550 ;
        RECT 22.780 262.000 22.930 264.900 ;
        RECT 18.730 261.700 22.930 262.000 ;
        RECT 6.530 261.550 14.080 261.700 ;
        RECT 15.380 261.550 22.930 261.700 ;
        RECT 6.530 261.350 10.730 261.550 ;
        RECT 4.730 261.050 9.130 261.200 ;
        RECT 9.280 261.050 10.730 261.350 ;
        RECT 4.730 260.150 10.730 261.050 ;
        RECT 18.730 261.350 22.930 261.550 ;
        RECT 18.730 261.050 20.180 261.350 ;
        RECT 23.530 261.200 25.930 264.400 ;
        RECT 26.530 262.000 26.680 264.900 ;
        RECT 27.130 262.000 27.280 269.550 ;
        RECT 27.730 262.000 27.880 269.550 ;
        RECT 28.330 262.000 28.480 269.550 ;
        RECT 28.930 262.000 29.080 269.550 ;
        RECT 29.530 262.000 29.680 269.550 ;
        RECT 30.130 269.350 34.080 269.550 ;
        RECT 35.380 269.350 39.330 269.550 ;
        RECT 30.130 268.900 30.730 269.350 ;
        RECT 38.730 268.900 39.330 269.350 ;
        RECT 30.130 268.750 34.080 268.900 ;
        RECT 35.380 268.750 39.330 268.900 ;
        RECT 30.130 268.300 30.730 268.750 ;
        RECT 38.730 268.300 39.330 268.750 ;
        RECT 30.130 268.150 34.080 268.300 ;
        RECT 35.380 268.150 39.330 268.300 ;
        RECT 30.130 267.700 30.730 268.150 ;
        RECT 38.730 267.700 39.330 268.150 ;
        RECT 30.130 267.550 34.080 267.700 ;
        RECT 35.380 267.550 39.330 267.700 ;
        RECT 30.130 267.100 30.730 267.550 ;
        RECT 38.730 267.100 39.330 267.550 ;
        RECT 30.130 266.950 34.080 267.100 ;
        RECT 35.380 266.950 39.330 267.100 ;
        RECT 30.130 266.500 30.730 266.950 ;
        RECT 38.730 266.500 39.330 266.950 ;
        RECT 30.130 266.350 34.080 266.500 ;
        RECT 35.380 266.350 39.330 266.500 ;
        RECT 30.130 265.900 30.730 266.350 ;
        RECT 38.730 265.900 39.330 266.350 ;
        RECT 30.130 265.750 34.080 265.900 ;
        RECT 35.380 265.750 39.330 265.900 ;
        RECT 30.130 265.300 30.730 265.750 ;
        RECT 38.730 265.300 39.330 265.750 ;
        RECT 30.130 265.150 34.080 265.300 ;
        RECT 35.380 265.150 39.330 265.300 ;
        RECT 30.130 264.700 30.730 265.150 ;
        RECT 38.730 264.700 39.330 265.150 ;
        RECT 30.130 264.550 34.080 264.700 ;
        RECT 35.380 264.550 39.330 264.700 ;
        RECT 30.130 264.100 30.730 264.550 ;
        RECT 38.730 264.100 39.330 264.550 ;
        RECT 30.130 263.950 34.080 264.100 ;
        RECT 35.380 263.950 39.330 264.100 ;
        RECT 30.130 263.500 30.730 263.950 ;
        RECT 38.730 263.500 39.330 263.950 ;
        RECT 30.130 263.350 34.080 263.500 ;
        RECT 35.380 263.350 39.330 263.500 ;
        RECT 30.130 262.900 30.730 263.350 ;
        RECT 38.730 262.900 39.330 263.350 ;
        RECT 30.130 262.750 34.080 262.900 ;
        RECT 35.380 262.750 39.330 262.900 ;
        RECT 30.130 262.300 30.730 262.750 ;
        RECT 38.730 262.300 39.330 262.750 ;
        RECT 30.130 262.150 34.080 262.300 ;
        RECT 35.380 262.150 39.330 262.300 ;
        RECT 30.130 262.000 30.730 262.150 ;
        RECT 26.530 261.700 30.730 262.000 ;
        RECT 38.730 262.000 39.330 262.150 ;
        RECT 39.780 262.000 39.930 269.550 ;
        RECT 40.380 262.000 40.530 269.550 ;
        RECT 40.980 262.000 41.130 269.550 ;
        RECT 41.580 262.000 41.730 269.550 ;
        RECT 42.180 262.000 42.330 269.550 ;
        RECT 42.780 262.000 42.930 264.900 ;
        RECT 38.730 261.700 42.930 262.000 ;
        RECT 26.530 261.550 34.080 261.700 ;
        RECT 35.380 261.550 42.930 261.700 ;
        RECT 26.530 261.350 30.730 261.550 ;
        RECT 20.330 261.050 29.130 261.200 ;
        RECT 29.280 261.050 30.730 261.350 ;
        RECT 18.730 260.150 30.730 261.050 ;
        RECT 38.730 261.350 42.930 261.550 ;
        RECT 38.730 261.050 40.180 261.350 ;
        RECT 43.530 261.200 45.930 264.400 ;
        RECT 46.530 262.000 46.680 264.900 ;
        RECT 47.130 262.000 47.280 269.550 ;
        RECT 47.730 262.000 47.880 269.550 ;
        RECT 48.330 262.000 48.480 269.550 ;
        RECT 48.930 262.000 49.080 269.550 ;
        RECT 49.530 262.000 49.680 269.550 ;
        RECT 50.130 269.350 54.080 269.550 ;
        RECT 55.380 269.350 59.330 269.550 ;
        RECT 50.130 268.900 50.730 269.350 ;
        RECT 58.730 268.900 59.330 269.350 ;
        RECT 50.130 268.750 54.080 268.900 ;
        RECT 55.380 268.750 59.330 268.900 ;
        RECT 50.130 268.300 50.730 268.750 ;
        RECT 58.730 268.300 59.330 268.750 ;
        RECT 50.130 268.150 54.080 268.300 ;
        RECT 55.380 268.150 59.330 268.300 ;
        RECT 50.130 267.700 50.730 268.150 ;
        RECT 58.730 267.700 59.330 268.150 ;
        RECT 50.130 267.550 54.080 267.700 ;
        RECT 55.380 267.550 59.330 267.700 ;
        RECT 50.130 267.100 50.730 267.550 ;
        RECT 58.730 267.100 59.330 267.550 ;
        RECT 50.130 266.950 54.080 267.100 ;
        RECT 55.380 266.950 59.330 267.100 ;
        RECT 50.130 266.500 50.730 266.950 ;
        RECT 58.730 266.500 59.330 266.950 ;
        RECT 50.130 266.350 54.080 266.500 ;
        RECT 55.380 266.350 59.330 266.500 ;
        RECT 50.130 265.900 50.730 266.350 ;
        RECT 58.730 265.900 59.330 266.350 ;
        RECT 50.130 265.750 54.080 265.900 ;
        RECT 55.380 265.750 59.330 265.900 ;
        RECT 50.130 265.300 50.730 265.750 ;
        RECT 58.730 265.300 59.330 265.750 ;
        RECT 50.130 265.150 54.080 265.300 ;
        RECT 55.380 265.150 59.330 265.300 ;
        RECT 50.130 264.700 50.730 265.150 ;
        RECT 58.730 264.700 59.330 265.150 ;
        RECT 50.130 264.550 54.080 264.700 ;
        RECT 55.380 264.550 59.330 264.700 ;
        RECT 50.130 264.100 50.730 264.550 ;
        RECT 58.730 264.100 59.330 264.550 ;
        RECT 50.130 263.950 54.080 264.100 ;
        RECT 55.380 263.950 59.330 264.100 ;
        RECT 50.130 263.500 50.730 263.950 ;
        RECT 58.730 263.500 59.330 263.950 ;
        RECT 50.130 263.350 54.080 263.500 ;
        RECT 55.380 263.350 59.330 263.500 ;
        RECT 50.130 262.900 50.730 263.350 ;
        RECT 58.730 262.900 59.330 263.350 ;
        RECT 50.130 262.750 54.080 262.900 ;
        RECT 55.380 262.750 59.330 262.900 ;
        RECT 50.130 262.300 50.730 262.750 ;
        RECT 58.730 262.300 59.330 262.750 ;
        RECT 50.130 262.150 54.080 262.300 ;
        RECT 55.380 262.150 59.330 262.300 ;
        RECT 50.130 262.000 50.730 262.150 ;
        RECT 46.530 261.700 50.730 262.000 ;
        RECT 58.730 262.000 59.330 262.150 ;
        RECT 59.780 262.000 59.930 269.550 ;
        RECT 60.380 262.000 60.530 269.550 ;
        RECT 60.980 262.000 61.130 269.550 ;
        RECT 61.580 262.000 61.730 269.550 ;
        RECT 62.180 262.000 62.330 269.550 ;
        RECT 62.780 262.000 62.930 264.900 ;
        RECT 58.730 261.700 62.930 262.000 ;
        RECT 46.530 261.550 54.080 261.700 ;
        RECT 55.380 261.550 62.930 261.700 ;
        RECT 46.530 261.350 50.730 261.550 ;
        RECT 40.330 261.050 49.130 261.200 ;
        RECT 49.280 261.050 50.730 261.350 ;
        RECT 38.730 260.150 50.730 261.050 ;
        RECT 58.730 261.350 62.930 261.550 ;
        RECT 58.730 261.050 60.180 261.350 ;
        RECT 63.530 261.200 65.930 264.400 ;
        RECT 66.530 262.000 66.680 264.900 ;
        RECT 67.130 262.000 67.280 269.550 ;
        RECT 67.730 262.000 67.880 269.550 ;
        RECT 68.330 262.000 68.480 269.550 ;
        RECT 68.930 262.000 69.080 269.550 ;
        RECT 69.530 262.000 69.680 269.550 ;
        RECT 70.130 269.350 74.080 269.550 ;
        RECT 75.380 269.350 79.330 269.550 ;
        RECT 70.130 268.900 70.730 269.350 ;
        RECT 78.730 268.900 79.330 269.350 ;
        RECT 70.130 268.750 74.080 268.900 ;
        RECT 75.380 268.750 79.330 268.900 ;
        RECT 70.130 268.300 70.730 268.750 ;
        RECT 78.730 268.300 79.330 268.750 ;
        RECT 70.130 268.150 74.080 268.300 ;
        RECT 75.380 268.150 79.330 268.300 ;
        RECT 70.130 267.700 70.730 268.150 ;
        RECT 78.730 267.700 79.330 268.150 ;
        RECT 70.130 267.550 74.080 267.700 ;
        RECT 75.380 267.550 79.330 267.700 ;
        RECT 70.130 267.100 70.730 267.550 ;
        RECT 78.730 267.100 79.330 267.550 ;
        RECT 70.130 266.950 74.080 267.100 ;
        RECT 75.380 266.950 79.330 267.100 ;
        RECT 70.130 266.500 70.730 266.950 ;
        RECT 78.730 266.500 79.330 266.950 ;
        RECT 70.130 266.350 74.080 266.500 ;
        RECT 75.380 266.350 79.330 266.500 ;
        RECT 70.130 265.900 70.730 266.350 ;
        RECT 78.730 265.900 79.330 266.350 ;
        RECT 70.130 265.750 74.080 265.900 ;
        RECT 75.380 265.750 79.330 265.900 ;
        RECT 70.130 265.300 70.730 265.750 ;
        RECT 78.730 265.300 79.330 265.750 ;
        RECT 70.130 265.150 74.080 265.300 ;
        RECT 75.380 265.150 79.330 265.300 ;
        RECT 70.130 264.700 70.730 265.150 ;
        RECT 78.730 264.700 79.330 265.150 ;
        RECT 70.130 264.550 74.080 264.700 ;
        RECT 75.380 264.550 79.330 264.700 ;
        RECT 70.130 264.100 70.730 264.550 ;
        RECT 78.730 264.100 79.330 264.550 ;
        RECT 70.130 263.950 74.080 264.100 ;
        RECT 75.380 263.950 79.330 264.100 ;
        RECT 70.130 263.500 70.730 263.950 ;
        RECT 78.730 263.500 79.330 263.950 ;
        RECT 70.130 263.350 74.080 263.500 ;
        RECT 75.380 263.350 79.330 263.500 ;
        RECT 70.130 262.900 70.730 263.350 ;
        RECT 78.730 262.900 79.330 263.350 ;
        RECT 70.130 262.750 74.080 262.900 ;
        RECT 75.380 262.750 79.330 262.900 ;
        RECT 70.130 262.300 70.730 262.750 ;
        RECT 78.730 262.300 79.330 262.750 ;
        RECT 70.130 262.150 74.080 262.300 ;
        RECT 75.380 262.150 79.330 262.300 ;
        RECT 70.130 262.000 70.730 262.150 ;
        RECT 66.530 261.700 70.730 262.000 ;
        RECT 78.730 262.000 79.330 262.150 ;
        RECT 79.780 262.000 79.930 269.550 ;
        RECT 80.380 262.000 80.530 269.550 ;
        RECT 80.980 262.000 81.130 269.550 ;
        RECT 81.580 262.000 81.730 269.550 ;
        RECT 82.180 262.000 82.330 269.550 ;
        RECT 82.780 262.000 82.930 264.900 ;
        RECT 78.730 261.700 82.930 262.000 ;
        RECT 66.530 261.550 74.080 261.700 ;
        RECT 75.380 261.550 82.930 261.700 ;
        RECT 66.530 261.350 70.730 261.550 ;
        RECT 60.330 261.050 69.130 261.200 ;
        RECT 69.280 261.050 70.730 261.350 ;
        RECT 58.730 260.150 70.730 261.050 ;
        RECT 78.730 261.350 82.930 261.550 ;
        RECT 78.730 261.050 80.180 261.350 ;
        RECT 83.530 261.200 85.930 264.400 ;
        RECT 86.530 262.000 86.680 264.900 ;
        RECT 87.130 262.000 87.280 269.550 ;
        RECT 87.730 262.000 87.880 269.550 ;
        RECT 88.330 262.000 88.480 269.550 ;
        RECT 88.930 262.000 89.080 269.550 ;
        RECT 89.530 262.000 89.680 269.550 ;
        RECT 90.130 269.350 94.080 269.550 ;
        RECT 95.380 269.350 99.330 269.550 ;
        RECT 90.130 268.900 90.730 269.350 ;
        RECT 98.730 268.900 99.330 269.350 ;
        RECT 90.130 268.750 94.080 268.900 ;
        RECT 95.380 268.750 99.330 268.900 ;
        RECT 90.130 268.300 90.730 268.750 ;
        RECT 98.730 268.300 99.330 268.750 ;
        RECT 90.130 268.150 94.080 268.300 ;
        RECT 95.380 268.150 99.330 268.300 ;
        RECT 90.130 267.700 90.730 268.150 ;
        RECT 98.730 267.700 99.330 268.150 ;
        RECT 90.130 267.550 94.080 267.700 ;
        RECT 95.380 267.550 99.330 267.700 ;
        RECT 90.130 267.100 90.730 267.550 ;
        RECT 98.730 267.100 99.330 267.550 ;
        RECT 90.130 266.950 94.080 267.100 ;
        RECT 95.380 266.950 99.330 267.100 ;
        RECT 90.130 266.500 90.730 266.950 ;
        RECT 98.730 266.500 99.330 266.950 ;
        RECT 90.130 266.350 94.080 266.500 ;
        RECT 95.380 266.350 99.330 266.500 ;
        RECT 90.130 265.900 90.730 266.350 ;
        RECT 98.730 265.900 99.330 266.350 ;
        RECT 90.130 265.750 94.080 265.900 ;
        RECT 95.380 265.750 99.330 265.900 ;
        RECT 90.130 265.300 90.730 265.750 ;
        RECT 98.730 265.300 99.330 265.750 ;
        RECT 90.130 265.150 94.080 265.300 ;
        RECT 95.380 265.150 99.330 265.300 ;
        RECT 90.130 264.700 90.730 265.150 ;
        RECT 98.730 264.700 99.330 265.150 ;
        RECT 90.130 264.550 94.080 264.700 ;
        RECT 95.380 264.550 99.330 264.700 ;
        RECT 90.130 264.100 90.730 264.550 ;
        RECT 98.730 264.100 99.330 264.550 ;
        RECT 90.130 263.950 94.080 264.100 ;
        RECT 95.380 263.950 99.330 264.100 ;
        RECT 90.130 263.500 90.730 263.950 ;
        RECT 98.730 263.500 99.330 263.950 ;
        RECT 90.130 263.350 94.080 263.500 ;
        RECT 95.380 263.350 99.330 263.500 ;
        RECT 90.130 262.900 90.730 263.350 ;
        RECT 98.730 262.900 99.330 263.350 ;
        RECT 90.130 262.750 94.080 262.900 ;
        RECT 95.380 262.750 99.330 262.900 ;
        RECT 90.130 262.300 90.730 262.750 ;
        RECT 98.730 262.300 99.330 262.750 ;
        RECT 90.130 262.150 94.080 262.300 ;
        RECT 95.380 262.150 99.330 262.300 ;
        RECT 90.130 262.000 90.730 262.150 ;
        RECT 86.530 261.700 90.730 262.000 ;
        RECT 98.730 262.000 99.330 262.150 ;
        RECT 99.780 262.000 99.930 269.550 ;
        RECT 100.380 262.000 100.530 269.550 ;
        RECT 100.980 262.000 101.130 269.550 ;
        RECT 101.580 262.000 101.730 269.550 ;
        RECT 102.180 262.000 102.330 269.550 ;
        RECT 102.780 262.000 102.930 264.900 ;
        RECT 98.730 261.700 102.930 262.000 ;
        RECT 86.530 261.550 94.080 261.700 ;
        RECT 95.380 261.550 102.930 261.700 ;
        RECT 86.530 261.350 90.730 261.550 ;
        RECT 80.330 261.050 89.130 261.200 ;
        RECT 89.280 261.050 90.730 261.350 ;
        RECT 78.730 260.150 90.730 261.050 ;
        RECT 98.730 261.350 102.930 261.550 ;
        RECT 103.530 263.000 104.730 264.400 ;
        RECT 103.530 261.725 107.140 263.000 ;
        RECT 98.730 261.050 100.180 261.350 ;
        RECT 103.530 261.200 104.730 261.725 ;
        RECT 100.330 261.050 104.730 261.200 ;
        RECT 98.730 260.150 104.730 261.050 ;
        RECT 4.730 259.850 9.130 260.150 ;
        RECT 20.330 259.850 29.130 260.150 ;
        RECT 40.330 259.850 49.130 260.150 ;
        RECT 60.330 259.850 69.130 260.150 ;
        RECT 80.330 259.850 89.130 260.150 ;
        RECT 4.730 258.950 10.730 259.850 ;
        RECT 20.330 259.800 30.730 259.850 ;
        RECT 40.330 259.800 50.730 259.850 ;
        RECT 60.330 259.800 70.730 259.850 ;
        RECT 80.330 259.800 90.730 259.850 ;
        RECT 100.330 259.800 104.730 260.150 ;
        RECT 4.730 258.800 9.130 258.950 ;
        RECT 4.730 257.845 5.930 258.800 ;
        RECT 9.280 258.650 10.730 258.950 ;
        RECT 2.315 256.570 5.930 257.845 ;
        RECT 4.730 255.600 5.930 256.570 ;
        RECT 6.530 258.450 10.730 258.650 ;
        RECT 18.730 258.950 30.730 259.800 ;
        RECT 18.730 258.900 29.130 258.950 ;
        RECT 18.730 258.650 20.180 258.900 ;
        RECT 20.330 258.800 29.130 258.900 ;
        RECT 18.730 258.450 22.930 258.650 ;
        RECT 6.530 258.300 14.080 258.450 ;
        RECT 15.430 258.300 22.930 258.450 ;
        RECT 6.530 258.000 10.730 258.300 ;
        RECT 2.315 253.250 4.315 255.545 ;
        RECT 6.530 255.150 6.680 258.000 ;
        RECT 7.130 250.450 7.280 258.000 ;
        RECT 7.730 250.450 7.880 258.000 ;
        RECT 8.330 250.450 8.480 258.000 ;
        RECT 8.930 250.450 9.080 258.000 ;
        RECT 9.530 250.450 9.680 258.000 ;
        RECT 10.130 257.850 10.730 258.000 ;
        RECT 18.730 258.000 22.930 258.300 ;
        RECT 18.730 257.850 19.330 258.000 ;
        RECT 10.130 257.700 14.080 257.850 ;
        RECT 15.380 257.700 19.330 257.850 ;
        RECT 10.130 257.250 10.730 257.700 ;
        RECT 18.730 257.250 19.330 257.700 ;
        RECT 10.130 257.100 14.080 257.250 ;
        RECT 15.380 257.100 19.330 257.250 ;
        RECT 10.130 256.650 10.730 257.100 ;
        RECT 18.730 256.650 19.330 257.100 ;
        RECT 10.130 256.500 14.080 256.650 ;
        RECT 15.380 256.500 19.330 256.650 ;
        RECT 10.130 256.050 10.730 256.500 ;
        RECT 18.730 256.050 19.330 256.500 ;
        RECT 10.130 255.900 14.080 256.050 ;
        RECT 15.380 255.900 19.330 256.050 ;
        RECT 10.130 255.450 10.730 255.900 ;
        RECT 18.730 255.450 19.330 255.900 ;
        RECT 10.130 255.300 14.080 255.450 ;
        RECT 15.380 255.300 19.330 255.450 ;
        RECT 10.130 254.850 10.730 255.300 ;
        RECT 18.730 254.850 19.330 255.300 ;
        RECT 10.130 254.700 14.080 254.850 ;
        RECT 15.380 254.700 19.330 254.850 ;
        RECT 10.130 254.250 10.730 254.700 ;
        RECT 18.730 254.250 19.330 254.700 ;
        RECT 10.130 254.100 14.080 254.250 ;
        RECT 15.380 254.100 19.330 254.250 ;
        RECT 10.130 253.650 10.730 254.100 ;
        RECT 18.730 253.650 19.330 254.100 ;
        RECT 10.130 253.500 14.080 253.650 ;
        RECT 15.380 253.500 19.330 253.650 ;
        RECT 10.130 253.050 10.730 253.500 ;
        RECT 18.730 253.050 19.330 253.500 ;
        RECT 10.130 252.900 14.080 253.050 ;
        RECT 15.380 252.900 19.330 253.050 ;
        RECT 10.130 252.450 10.730 252.900 ;
        RECT 18.730 252.450 19.330 252.900 ;
        RECT 10.130 252.300 14.080 252.450 ;
        RECT 15.380 252.300 19.330 252.450 ;
        RECT 10.130 251.850 10.730 252.300 ;
        RECT 18.730 251.850 19.330 252.300 ;
        RECT 10.130 251.700 14.080 251.850 ;
        RECT 15.380 251.700 19.330 251.850 ;
        RECT 10.130 251.250 10.730 251.700 ;
        RECT 18.730 251.250 19.330 251.700 ;
        RECT 10.130 251.100 14.080 251.250 ;
        RECT 15.380 251.100 19.330 251.250 ;
        RECT 10.130 250.650 10.730 251.100 ;
        RECT 18.730 250.650 19.330 251.100 ;
        RECT 10.130 250.450 14.080 250.650 ;
        RECT 15.380 250.450 19.330 250.650 ;
        RECT 19.780 250.450 19.930 258.000 ;
        RECT 20.380 250.450 20.530 258.000 ;
        RECT 20.980 250.450 21.130 258.000 ;
        RECT 21.580 250.450 21.730 258.000 ;
        RECT 22.180 250.450 22.330 258.000 ;
        RECT 22.780 255.150 22.930 258.000 ;
        RECT 23.530 255.600 25.930 258.800 ;
        RECT 29.280 258.650 30.730 258.950 ;
        RECT 26.530 258.450 30.730 258.650 ;
        RECT 38.730 258.950 50.730 259.800 ;
        RECT 38.730 258.900 49.130 258.950 ;
        RECT 38.730 258.650 40.180 258.900 ;
        RECT 40.330 258.800 49.130 258.900 ;
        RECT 38.730 258.450 42.930 258.650 ;
        RECT 26.530 258.300 34.080 258.450 ;
        RECT 35.430 258.300 42.930 258.450 ;
        RECT 26.530 258.000 30.730 258.300 ;
        RECT 26.530 255.150 26.680 258.000 ;
        RECT 27.130 250.450 27.280 258.000 ;
        RECT 27.730 250.450 27.880 258.000 ;
        RECT 28.330 250.450 28.480 258.000 ;
        RECT 28.930 250.450 29.080 258.000 ;
        RECT 29.530 250.450 29.680 258.000 ;
        RECT 30.130 257.850 30.730 258.000 ;
        RECT 38.730 258.000 42.930 258.300 ;
        RECT 38.730 257.850 39.330 258.000 ;
        RECT 30.130 257.700 34.080 257.850 ;
        RECT 35.380 257.700 39.330 257.850 ;
        RECT 30.130 257.250 30.730 257.700 ;
        RECT 38.730 257.250 39.330 257.700 ;
        RECT 30.130 257.100 34.080 257.250 ;
        RECT 35.380 257.100 39.330 257.250 ;
        RECT 30.130 256.650 30.730 257.100 ;
        RECT 38.730 256.650 39.330 257.100 ;
        RECT 30.130 256.500 34.080 256.650 ;
        RECT 35.380 256.500 39.330 256.650 ;
        RECT 30.130 256.050 30.730 256.500 ;
        RECT 38.730 256.050 39.330 256.500 ;
        RECT 30.130 255.900 34.080 256.050 ;
        RECT 35.380 255.900 39.330 256.050 ;
        RECT 30.130 255.450 30.730 255.900 ;
        RECT 38.730 255.450 39.330 255.900 ;
        RECT 30.130 255.300 34.080 255.450 ;
        RECT 35.380 255.300 39.330 255.450 ;
        RECT 30.130 254.850 30.730 255.300 ;
        RECT 38.730 254.850 39.330 255.300 ;
        RECT 30.130 254.700 34.080 254.850 ;
        RECT 35.380 254.700 39.330 254.850 ;
        RECT 30.130 254.250 30.730 254.700 ;
        RECT 38.730 254.250 39.330 254.700 ;
        RECT 30.130 254.100 34.080 254.250 ;
        RECT 35.380 254.100 39.330 254.250 ;
        RECT 30.130 253.650 30.730 254.100 ;
        RECT 38.730 253.650 39.330 254.100 ;
        RECT 30.130 253.500 34.080 253.650 ;
        RECT 35.380 253.500 39.330 253.650 ;
        RECT 30.130 253.050 30.730 253.500 ;
        RECT 38.730 253.050 39.330 253.500 ;
        RECT 30.130 252.900 34.080 253.050 ;
        RECT 35.380 252.900 39.330 253.050 ;
        RECT 30.130 252.450 30.730 252.900 ;
        RECT 38.730 252.450 39.330 252.900 ;
        RECT 30.130 252.300 34.080 252.450 ;
        RECT 35.380 252.300 39.330 252.450 ;
        RECT 30.130 251.850 30.730 252.300 ;
        RECT 38.730 251.850 39.330 252.300 ;
        RECT 30.130 251.700 34.080 251.850 ;
        RECT 35.380 251.700 39.330 251.850 ;
        RECT 30.130 251.250 30.730 251.700 ;
        RECT 38.730 251.250 39.330 251.700 ;
        RECT 30.130 251.100 34.080 251.250 ;
        RECT 35.380 251.100 39.330 251.250 ;
        RECT 30.130 250.650 30.730 251.100 ;
        RECT 38.730 250.650 39.330 251.100 ;
        RECT 30.130 250.450 34.080 250.650 ;
        RECT 35.380 250.450 39.330 250.650 ;
        RECT 39.780 250.450 39.930 258.000 ;
        RECT 40.380 250.450 40.530 258.000 ;
        RECT 40.980 250.450 41.130 258.000 ;
        RECT 41.580 250.450 41.730 258.000 ;
        RECT 42.180 250.450 42.330 258.000 ;
        RECT 42.780 255.150 42.930 258.000 ;
        RECT 43.530 255.600 45.930 258.800 ;
        RECT 49.280 258.650 50.730 258.950 ;
        RECT 46.530 258.450 50.730 258.650 ;
        RECT 58.730 258.950 70.730 259.800 ;
        RECT 58.730 258.900 69.130 258.950 ;
        RECT 58.730 258.650 60.180 258.900 ;
        RECT 60.330 258.800 69.130 258.900 ;
        RECT 58.730 258.450 62.930 258.650 ;
        RECT 46.530 258.300 54.080 258.450 ;
        RECT 55.430 258.300 62.930 258.450 ;
        RECT 46.530 258.000 50.730 258.300 ;
        RECT 46.530 255.150 46.680 258.000 ;
        RECT 47.130 250.450 47.280 258.000 ;
        RECT 47.730 250.450 47.880 258.000 ;
        RECT 48.330 250.450 48.480 258.000 ;
        RECT 48.930 250.450 49.080 258.000 ;
        RECT 49.530 250.450 49.680 258.000 ;
        RECT 50.130 257.850 50.730 258.000 ;
        RECT 58.730 258.000 62.930 258.300 ;
        RECT 58.730 257.850 59.330 258.000 ;
        RECT 50.130 257.700 54.080 257.850 ;
        RECT 55.380 257.700 59.330 257.850 ;
        RECT 50.130 257.250 50.730 257.700 ;
        RECT 58.730 257.250 59.330 257.700 ;
        RECT 50.130 257.100 54.080 257.250 ;
        RECT 55.380 257.100 59.330 257.250 ;
        RECT 50.130 256.650 50.730 257.100 ;
        RECT 58.730 256.650 59.330 257.100 ;
        RECT 50.130 256.500 54.080 256.650 ;
        RECT 55.380 256.500 59.330 256.650 ;
        RECT 50.130 256.050 50.730 256.500 ;
        RECT 58.730 256.050 59.330 256.500 ;
        RECT 50.130 255.900 54.080 256.050 ;
        RECT 55.380 255.900 59.330 256.050 ;
        RECT 50.130 255.450 50.730 255.900 ;
        RECT 58.730 255.450 59.330 255.900 ;
        RECT 50.130 255.300 54.080 255.450 ;
        RECT 55.380 255.300 59.330 255.450 ;
        RECT 50.130 254.850 50.730 255.300 ;
        RECT 58.730 254.850 59.330 255.300 ;
        RECT 50.130 254.700 54.080 254.850 ;
        RECT 55.380 254.700 59.330 254.850 ;
        RECT 50.130 254.250 50.730 254.700 ;
        RECT 58.730 254.250 59.330 254.700 ;
        RECT 50.130 254.100 54.080 254.250 ;
        RECT 55.380 254.100 59.330 254.250 ;
        RECT 50.130 253.650 50.730 254.100 ;
        RECT 58.730 253.650 59.330 254.100 ;
        RECT 50.130 253.500 54.080 253.650 ;
        RECT 55.380 253.500 59.330 253.650 ;
        RECT 50.130 253.050 50.730 253.500 ;
        RECT 58.730 253.050 59.330 253.500 ;
        RECT 50.130 252.900 54.080 253.050 ;
        RECT 55.380 252.900 59.330 253.050 ;
        RECT 50.130 252.450 50.730 252.900 ;
        RECT 58.730 252.450 59.330 252.900 ;
        RECT 50.130 252.300 54.080 252.450 ;
        RECT 55.380 252.300 59.330 252.450 ;
        RECT 50.130 251.850 50.730 252.300 ;
        RECT 58.730 251.850 59.330 252.300 ;
        RECT 50.130 251.700 54.080 251.850 ;
        RECT 55.380 251.700 59.330 251.850 ;
        RECT 50.130 251.250 50.730 251.700 ;
        RECT 58.730 251.250 59.330 251.700 ;
        RECT 50.130 251.100 54.080 251.250 ;
        RECT 55.380 251.100 59.330 251.250 ;
        RECT 50.130 250.650 50.730 251.100 ;
        RECT 58.730 250.650 59.330 251.100 ;
        RECT 50.130 250.450 54.080 250.650 ;
        RECT 55.380 250.450 59.330 250.650 ;
        RECT 59.780 250.450 59.930 258.000 ;
        RECT 60.380 250.450 60.530 258.000 ;
        RECT 60.980 250.450 61.130 258.000 ;
        RECT 61.580 250.450 61.730 258.000 ;
        RECT 62.180 250.450 62.330 258.000 ;
        RECT 62.780 255.150 62.930 258.000 ;
        RECT 63.530 255.600 65.930 258.800 ;
        RECT 69.280 258.650 70.730 258.950 ;
        RECT 66.530 258.450 70.730 258.650 ;
        RECT 78.730 258.950 90.730 259.800 ;
        RECT 78.730 258.900 89.130 258.950 ;
        RECT 78.730 258.650 80.180 258.900 ;
        RECT 80.330 258.800 89.130 258.900 ;
        RECT 78.730 258.450 82.930 258.650 ;
        RECT 66.530 258.300 74.080 258.450 ;
        RECT 75.430 258.300 82.930 258.450 ;
        RECT 66.530 258.000 70.730 258.300 ;
        RECT 66.530 255.150 66.680 258.000 ;
        RECT 67.130 250.450 67.280 258.000 ;
        RECT 67.730 250.450 67.880 258.000 ;
        RECT 68.330 250.450 68.480 258.000 ;
        RECT 68.930 250.450 69.080 258.000 ;
        RECT 69.530 250.450 69.680 258.000 ;
        RECT 70.130 257.850 70.730 258.000 ;
        RECT 78.730 258.000 82.930 258.300 ;
        RECT 78.730 257.850 79.330 258.000 ;
        RECT 70.130 257.700 74.080 257.850 ;
        RECT 75.380 257.700 79.330 257.850 ;
        RECT 70.130 257.250 70.730 257.700 ;
        RECT 78.730 257.250 79.330 257.700 ;
        RECT 70.130 257.100 74.080 257.250 ;
        RECT 75.380 257.100 79.330 257.250 ;
        RECT 70.130 256.650 70.730 257.100 ;
        RECT 78.730 256.650 79.330 257.100 ;
        RECT 70.130 256.500 74.080 256.650 ;
        RECT 75.380 256.500 79.330 256.650 ;
        RECT 70.130 256.050 70.730 256.500 ;
        RECT 78.730 256.050 79.330 256.500 ;
        RECT 70.130 255.900 74.080 256.050 ;
        RECT 75.380 255.900 79.330 256.050 ;
        RECT 70.130 255.450 70.730 255.900 ;
        RECT 78.730 255.450 79.330 255.900 ;
        RECT 70.130 255.300 74.080 255.450 ;
        RECT 75.380 255.300 79.330 255.450 ;
        RECT 70.130 254.850 70.730 255.300 ;
        RECT 78.730 254.850 79.330 255.300 ;
        RECT 70.130 254.700 74.080 254.850 ;
        RECT 75.380 254.700 79.330 254.850 ;
        RECT 70.130 254.250 70.730 254.700 ;
        RECT 78.730 254.250 79.330 254.700 ;
        RECT 70.130 254.100 74.080 254.250 ;
        RECT 75.380 254.100 79.330 254.250 ;
        RECT 70.130 253.650 70.730 254.100 ;
        RECT 78.730 253.650 79.330 254.100 ;
        RECT 70.130 253.500 74.080 253.650 ;
        RECT 75.380 253.500 79.330 253.650 ;
        RECT 70.130 253.050 70.730 253.500 ;
        RECT 78.730 253.050 79.330 253.500 ;
        RECT 70.130 252.900 74.080 253.050 ;
        RECT 75.380 252.900 79.330 253.050 ;
        RECT 70.130 252.450 70.730 252.900 ;
        RECT 78.730 252.450 79.330 252.900 ;
        RECT 70.130 252.300 74.080 252.450 ;
        RECT 75.380 252.300 79.330 252.450 ;
        RECT 70.130 251.850 70.730 252.300 ;
        RECT 78.730 251.850 79.330 252.300 ;
        RECT 70.130 251.700 74.080 251.850 ;
        RECT 75.380 251.700 79.330 251.850 ;
        RECT 70.130 251.250 70.730 251.700 ;
        RECT 78.730 251.250 79.330 251.700 ;
        RECT 70.130 251.100 74.080 251.250 ;
        RECT 75.380 251.100 79.330 251.250 ;
        RECT 70.130 250.650 70.730 251.100 ;
        RECT 78.730 250.650 79.330 251.100 ;
        RECT 70.130 250.450 74.080 250.650 ;
        RECT 75.380 250.450 79.330 250.650 ;
        RECT 79.780 250.450 79.930 258.000 ;
        RECT 80.380 250.450 80.530 258.000 ;
        RECT 80.980 250.450 81.130 258.000 ;
        RECT 81.580 250.450 81.730 258.000 ;
        RECT 82.180 250.450 82.330 258.000 ;
        RECT 82.780 255.150 82.930 258.000 ;
        RECT 83.530 255.600 85.930 258.800 ;
        RECT 89.280 258.650 90.730 258.950 ;
        RECT 86.530 258.450 90.730 258.650 ;
        RECT 98.730 258.900 104.730 259.800 ;
        RECT 98.730 258.650 100.180 258.900 ;
        RECT 100.330 258.800 104.730 258.900 ;
        RECT 98.730 258.450 102.930 258.650 ;
        RECT 86.530 258.300 94.080 258.450 ;
        RECT 95.430 258.300 102.930 258.450 ;
        RECT 86.530 258.000 90.730 258.300 ;
        RECT 86.530 255.150 86.680 258.000 ;
        RECT 87.130 250.450 87.280 258.000 ;
        RECT 87.730 250.450 87.880 258.000 ;
        RECT 88.330 250.450 88.480 258.000 ;
        RECT 88.930 250.450 89.080 258.000 ;
        RECT 89.530 250.450 89.680 258.000 ;
        RECT 90.130 257.850 90.730 258.000 ;
        RECT 98.730 258.000 102.930 258.300 ;
        RECT 98.730 257.850 99.330 258.000 ;
        RECT 90.130 257.700 94.080 257.850 ;
        RECT 95.380 257.700 99.330 257.850 ;
        RECT 90.130 257.250 90.730 257.700 ;
        RECT 98.730 257.250 99.330 257.700 ;
        RECT 90.130 257.100 94.080 257.250 ;
        RECT 95.380 257.100 99.330 257.250 ;
        RECT 90.130 256.650 90.730 257.100 ;
        RECT 98.730 256.650 99.330 257.100 ;
        RECT 90.130 256.500 94.080 256.650 ;
        RECT 95.380 256.500 99.330 256.650 ;
        RECT 90.130 256.050 90.730 256.500 ;
        RECT 98.730 256.050 99.330 256.500 ;
        RECT 90.130 255.900 94.080 256.050 ;
        RECT 95.380 255.900 99.330 256.050 ;
        RECT 90.130 255.450 90.730 255.900 ;
        RECT 98.730 255.450 99.330 255.900 ;
        RECT 90.130 255.300 94.080 255.450 ;
        RECT 95.380 255.300 99.330 255.450 ;
        RECT 90.130 254.850 90.730 255.300 ;
        RECT 98.730 254.850 99.330 255.300 ;
        RECT 90.130 254.700 94.080 254.850 ;
        RECT 95.380 254.700 99.330 254.850 ;
        RECT 90.130 254.250 90.730 254.700 ;
        RECT 98.730 254.250 99.330 254.700 ;
        RECT 90.130 254.100 94.080 254.250 ;
        RECT 95.380 254.100 99.330 254.250 ;
        RECT 90.130 253.650 90.730 254.100 ;
        RECT 98.730 253.650 99.330 254.100 ;
        RECT 90.130 253.500 94.080 253.650 ;
        RECT 95.380 253.500 99.330 253.650 ;
        RECT 90.130 253.050 90.730 253.500 ;
        RECT 98.730 253.050 99.330 253.500 ;
        RECT 90.130 252.900 94.080 253.050 ;
        RECT 95.380 252.900 99.330 253.050 ;
        RECT 90.130 252.450 90.730 252.900 ;
        RECT 98.730 252.450 99.330 252.900 ;
        RECT 90.130 252.300 94.080 252.450 ;
        RECT 95.380 252.300 99.330 252.450 ;
        RECT 90.130 251.850 90.730 252.300 ;
        RECT 98.730 251.850 99.330 252.300 ;
        RECT 90.130 251.700 94.080 251.850 ;
        RECT 95.380 251.700 99.330 251.850 ;
        RECT 90.130 251.250 90.730 251.700 ;
        RECT 98.730 251.250 99.330 251.700 ;
        RECT 90.130 251.100 94.080 251.250 ;
        RECT 95.380 251.100 99.330 251.250 ;
        RECT 90.130 250.650 90.730 251.100 ;
        RECT 98.730 250.650 99.330 251.100 ;
        RECT 90.130 250.450 94.080 250.650 ;
        RECT 95.380 250.450 99.330 250.650 ;
        RECT 99.780 250.450 99.930 258.000 ;
        RECT 100.380 250.450 100.530 258.000 ;
        RECT 100.980 250.450 101.130 258.000 ;
        RECT 101.580 250.450 101.730 258.000 ;
        RECT 102.180 250.450 102.330 258.000 ;
        RECT 102.780 255.150 102.930 258.000 ;
        RECT 103.530 257.325 104.730 258.800 ;
        RECT 103.530 256.050 107.140 257.325 ;
        RECT 103.530 255.600 104.730 256.050 ;
        RECT 2.315 244.455 4.315 246.750 ;
        RECT 4.730 243.735 5.930 244.400 ;
        RECT 2.315 242.460 5.930 243.735 ;
        RECT 4.730 241.200 5.930 242.460 ;
        RECT 6.530 242.000 6.680 244.900 ;
        RECT 7.130 242.000 7.280 249.550 ;
        RECT 7.730 242.000 7.880 249.550 ;
        RECT 8.330 242.000 8.480 249.550 ;
        RECT 8.930 242.000 9.080 249.550 ;
        RECT 9.530 242.000 9.680 249.550 ;
        RECT 10.130 249.350 14.080 249.550 ;
        RECT 15.380 249.350 19.330 249.550 ;
        RECT 10.130 248.900 10.730 249.350 ;
        RECT 18.730 248.900 19.330 249.350 ;
        RECT 10.130 248.750 14.080 248.900 ;
        RECT 15.380 248.750 19.330 248.900 ;
        RECT 10.130 248.300 10.730 248.750 ;
        RECT 18.730 248.300 19.330 248.750 ;
        RECT 10.130 248.150 14.080 248.300 ;
        RECT 15.380 248.150 19.330 248.300 ;
        RECT 10.130 247.700 10.730 248.150 ;
        RECT 18.730 247.700 19.330 248.150 ;
        RECT 10.130 247.550 14.080 247.700 ;
        RECT 15.380 247.550 19.330 247.700 ;
        RECT 10.130 247.100 10.730 247.550 ;
        RECT 18.730 247.100 19.330 247.550 ;
        RECT 10.130 246.950 14.080 247.100 ;
        RECT 15.380 246.950 19.330 247.100 ;
        RECT 10.130 246.500 10.730 246.950 ;
        RECT 18.730 246.500 19.330 246.950 ;
        RECT 10.130 246.350 14.080 246.500 ;
        RECT 15.380 246.350 19.330 246.500 ;
        RECT 10.130 245.900 10.730 246.350 ;
        RECT 18.730 245.900 19.330 246.350 ;
        RECT 10.130 245.750 14.080 245.900 ;
        RECT 15.380 245.750 19.330 245.900 ;
        RECT 10.130 245.300 10.730 245.750 ;
        RECT 18.730 245.300 19.330 245.750 ;
        RECT 10.130 245.150 14.080 245.300 ;
        RECT 15.380 245.150 19.330 245.300 ;
        RECT 10.130 244.700 10.730 245.150 ;
        RECT 18.730 244.700 19.330 245.150 ;
        RECT 10.130 244.550 14.080 244.700 ;
        RECT 15.380 244.550 19.330 244.700 ;
        RECT 10.130 244.100 10.730 244.550 ;
        RECT 18.730 244.100 19.330 244.550 ;
        RECT 10.130 243.950 14.080 244.100 ;
        RECT 15.380 243.950 19.330 244.100 ;
        RECT 10.130 243.500 10.730 243.950 ;
        RECT 18.730 243.500 19.330 243.950 ;
        RECT 10.130 243.350 14.080 243.500 ;
        RECT 15.380 243.350 19.330 243.500 ;
        RECT 10.130 242.900 10.730 243.350 ;
        RECT 18.730 242.900 19.330 243.350 ;
        RECT 10.130 242.750 14.080 242.900 ;
        RECT 15.380 242.750 19.330 242.900 ;
        RECT 10.130 242.300 10.730 242.750 ;
        RECT 18.730 242.300 19.330 242.750 ;
        RECT 10.130 242.150 14.080 242.300 ;
        RECT 15.380 242.150 19.330 242.300 ;
        RECT 10.130 242.000 10.730 242.150 ;
        RECT 6.530 241.700 10.730 242.000 ;
        RECT 18.730 242.000 19.330 242.150 ;
        RECT 19.780 242.000 19.930 249.550 ;
        RECT 20.380 242.000 20.530 249.550 ;
        RECT 20.980 242.000 21.130 249.550 ;
        RECT 21.580 242.000 21.730 249.550 ;
        RECT 22.180 242.000 22.330 249.550 ;
        RECT 22.780 242.000 22.930 244.900 ;
        RECT 18.730 241.700 22.930 242.000 ;
        RECT 6.530 241.550 14.080 241.700 ;
        RECT 15.380 241.550 22.930 241.700 ;
        RECT 6.530 241.350 10.730 241.550 ;
        RECT 4.730 241.050 9.130 241.200 ;
        RECT 9.280 241.050 10.730 241.350 ;
        RECT 4.730 240.150 10.730 241.050 ;
        RECT 18.730 241.350 22.930 241.550 ;
        RECT 18.730 241.050 20.180 241.350 ;
        RECT 23.530 241.200 25.930 244.400 ;
        RECT 26.530 242.000 26.680 244.900 ;
        RECT 27.130 242.000 27.280 249.550 ;
        RECT 27.730 242.000 27.880 249.550 ;
        RECT 28.330 242.000 28.480 249.550 ;
        RECT 28.930 242.000 29.080 249.550 ;
        RECT 29.530 242.000 29.680 249.550 ;
        RECT 30.130 249.350 34.080 249.550 ;
        RECT 35.380 249.350 39.330 249.550 ;
        RECT 30.130 248.900 30.730 249.350 ;
        RECT 38.730 248.900 39.330 249.350 ;
        RECT 30.130 248.750 34.080 248.900 ;
        RECT 35.380 248.750 39.330 248.900 ;
        RECT 30.130 248.300 30.730 248.750 ;
        RECT 38.730 248.300 39.330 248.750 ;
        RECT 30.130 248.150 34.080 248.300 ;
        RECT 35.380 248.150 39.330 248.300 ;
        RECT 30.130 247.700 30.730 248.150 ;
        RECT 38.730 247.700 39.330 248.150 ;
        RECT 30.130 247.550 34.080 247.700 ;
        RECT 35.380 247.550 39.330 247.700 ;
        RECT 30.130 247.100 30.730 247.550 ;
        RECT 38.730 247.100 39.330 247.550 ;
        RECT 30.130 246.950 34.080 247.100 ;
        RECT 35.380 246.950 39.330 247.100 ;
        RECT 30.130 246.500 30.730 246.950 ;
        RECT 38.730 246.500 39.330 246.950 ;
        RECT 30.130 246.350 34.080 246.500 ;
        RECT 35.380 246.350 39.330 246.500 ;
        RECT 30.130 245.900 30.730 246.350 ;
        RECT 38.730 245.900 39.330 246.350 ;
        RECT 30.130 245.750 34.080 245.900 ;
        RECT 35.380 245.750 39.330 245.900 ;
        RECT 30.130 245.300 30.730 245.750 ;
        RECT 38.730 245.300 39.330 245.750 ;
        RECT 30.130 245.150 34.080 245.300 ;
        RECT 35.380 245.150 39.330 245.300 ;
        RECT 30.130 244.700 30.730 245.150 ;
        RECT 38.730 244.700 39.330 245.150 ;
        RECT 30.130 244.550 34.080 244.700 ;
        RECT 35.380 244.550 39.330 244.700 ;
        RECT 30.130 244.100 30.730 244.550 ;
        RECT 38.730 244.100 39.330 244.550 ;
        RECT 30.130 243.950 34.080 244.100 ;
        RECT 35.380 243.950 39.330 244.100 ;
        RECT 30.130 243.500 30.730 243.950 ;
        RECT 38.730 243.500 39.330 243.950 ;
        RECT 30.130 243.350 34.080 243.500 ;
        RECT 35.380 243.350 39.330 243.500 ;
        RECT 30.130 242.900 30.730 243.350 ;
        RECT 38.730 242.900 39.330 243.350 ;
        RECT 30.130 242.750 34.080 242.900 ;
        RECT 35.380 242.750 39.330 242.900 ;
        RECT 30.130 242.300 30.730 242.750 ;
        RECT 38.730 242.300 39.330 242.750 ;
        RECT 30.130 242.150 34.080 242.300 ;
        RECT 35.380 242.150 39.330 242.300 ;
        RECT 30.130 242.000 30.730 242.150 ;
        RECT 26.530 241.700 30.730 242.000 ;
        RECT 38.730 242.000 39.330 242.150 ;
        RECT 39.780 242.000 39.930 249.550 ;
        RECT 40.380 242.000 40.530 249.550 ;
        RECT 40.980 242.000 41.130 249.550 ;
        RECT 41.580 242.000 41.730 249.550 ;
        RECT 42.180 242.000 42.330 249.550 ;
        RECT 42.780 242.000 42.930 244.900 ;
        RECT 38.730 241.700 42.930 242.000 ;
        RECT 26.530 241.550 34.080 241.700 ;
        RECT 35.380 241.550 42.930 241.700 ;
        RECT 26.530 241.350 30.730 241.550 ;
        RECT 20.330 241.050 29.130 241.200 ;
        RECT 29.280 241.050 30.730 241.350 ;
        RECT 18.730 240.150 30.730 241.050 ;
        RECT 38.730 241.350 42.930 241.550 ;
        RECT 38.730 241.050 40.180 241.350 ;
        RECT 43.530 241.200 45.930 244.400 ;
        RECT 46.530 242.000 46.680 244.900 ;
        RECT 47.130 242.000 47.280 249.550 ;
        RECT 47.730 242.000 47.880 249.550 ;
        RECT 48.330 242.000 48.480 249.550 ;
        RECT 48.930 242.000 49.080 249.550 ;
        RECT 49.530 242.000 49.680 249.550 ;
        RECT 50.130 249.350 54.080 249.550 ;
        RECT 55.380 249.350 59.330 249.550 ;
        RECT 50.130 248.900 50.730 249.350 ;
        RECT 58.730 248.900 59.330 249.350 ;
        RECT 50.130 248.750 54.080 248.900 ;
        RECT 55.380 248.750 59.330 248.900 ;
        RECT 50.130 248.300 50.730 248.750 ;
        RECT 58.730 248.300 59.330 248.750 ;
        RECT 50.130 248.150 54.080 248.300 ;
        RECT 55.380 248.150 59.330 248.300 ;
        RECT 50.130 247.700 50.730 248.150 ;
        RECT 58.730 247.700 59.330 248.150 ;
        RECT 50.130 247.550 54.080 247.700 ;
        RECT 55.380 247.550 59.330 247.700 ;
        RECT 50.130 247.100 50.730 247.550 ;
        RECT 58.730 247.100 59.330 247.550 ;
        RECT 50.130 246.950 54.080 247.100 ;
        RECT 55.380 246.950 59.330 247.100 ;
        RECT 50.130 246.500 50.730 246.950 ;
        RECT 58.730 246.500 59.330 246.950 ;
        RECT 50.130 246.350 54.080 246.500 ;
        RECT 55.380 246.350 59.330 246.500 ;
        RECT 50.130 245.900 50.730 246.350 ;
        RECT 58.730 245.900 59.330 246.350 ;
        RECT 50.130 245.750 54.080 245.900 ;
        RECT 55.380 245.750 59.330 245.900 ;
        RECT 50.130 245.300 50.730 245.750 ;
        RECT 58.730 245.300 59.330 245.750 ;
        RECT 50.130 245.150 54.080 245.300 ;
        RECT 55.380 245.150 59.330 245.300 ;
        RECT 50.130 244.700 50.730 245.150 ;
        RECT 58.730 244.700 59.330 245.150 ;
        RECT 50.130 244.550 54.080 244.700 ;
        RECT 55.380 244.550 59.330 244.700 ;
        RECT 50.130 244.100 50.730 244.550 ;
        RECT 58.730 244.100 59.330 244.550 ;
        RECT 50.130 243.950 54.080 244.100 ;
        RECT 55.380 243.950 59.330 244.100 ;
        RECT 50.130 243.500 50.730 243.950 ;
        RECT 58.730 243.500 59.330 243.950 ;
        RECT 50.130 243.350 54.080 243.500 ;
        RECT 55.380 243.350 59.330 243.500 ;
        RECT 50.130 242.900 50.730 243.350 ;
        RECT 58.730 242.900 59.330 243.350 ;
        RECT 50.130 242.750 54.080 242.900 ;
        RECT 55.380 242.750 59.330 242.900 ;
        RECT 50.130 242.300 50.730 242.750 ;
        RECT 58.730 242.300 59.330 242.750 ;
        RECT 50.130 242.150 54.080 242.300 ;
        RECT 55.380 242.150 59.330 242.300 ;
        RECT 50.130 242.000 50.730 242.150 ;
        RECT 46.530 241.700 50.730 242.000 ;
        RECT 58.730 242.000 59.330 242.150 ;
        RECT 59.780 242.000 59.930 249.550 ;
        RECT 60.380 242.000 60.530 249.550 ;
        RECT 60.980 242.000 61.130 249.550 ;
        RECT 61.580 242.000 61.730 249.550 ;
        RECT 62.180 242.000 62.330 249.550 ;
        RECT 62.780 242.000 62.930 244.900 ;
        RECT 58.730 241.700 62.930 242.000 ;
        RECT 46.530 241.550 54.080 241.700 ;
        RECT 55.380 241.550 62.930 241.700 ;
        RECT 46.530 241.350 50.730 241.550 ;
        RECT 40.330 241.050 49.130 241.200 ;
        RECT 49.280 241.050 50.730 241.350 ;
        RECT 38.730 240.150 50.730 241.050 ;
        RECT 58.730 241.350 62.930 241.550 ;
        RECT 58.730 241.050 60.180 241.350 ;
        RECT 63.530 241.200 65.930 244.400 ;
        RECT 66.530 242.000 66.680 244.900 ;
        RECT 67.130 242.000 67.280 249.550 ;
        RECT 67.730 242.000 67.880 249.550 ;
        RECT 68.330 242.000 68.480 249.550 ;
        RECT 68.930 242.000 69.080 249.550 ;
        RECT 69.530 242.000 69.680 249.550 ;
        RECT 70.130 249.350 74.080 249.550 ;
        RECT 75.380 249.350 79.330 249.550 ;
        RECT 70.130 248.900 70.730 249.350 ;
        RECT 78.730 248.900 79.330 249.350 ;
        RECT 70.130 248.750 74.080 248.900 ;
        RECT 75.380 248.750 79.330 248.900 ;
        RECT 70.130 248.300 70.730 248.750 ;
        RECT 78.730 248.300 79.330 248.750 ;
        RECT 70.130 248.150 74.080 248.300 ;
        RECT 75.380 248.150 79.330 248.300 ;
        RECT 70.130 247.700 70.730 248.150 ;
        RECT 78.730 247.700 79.330 248.150 ;
        RECT 70.130 247.550 74.080 247.700 ;
        RECT 75.380 247.550 79.330 247.700 ;
        RECT 70.130 247.100 70.730 247.550 ;
        RECT 78.730 247.100 79.330 247.550 ;
        RECT 70.130 246.950 74.080 247.100 ;
        RECT 75.380 246.950 79.330 247.100 ;
        RECT 70.130 246.500 70.730 246.950 ;
        RECT 78.730 246.500 79.330 246.950 ;
        RECT 70.130 246.350 74.080 246.500 ;
        RECT 75.380 246.350 79.330 246.500 ;
        RECT 70.130 245.900 70.730 246.350 ;
        RECT 78.730 245.900 79.330 246.350 ;
        RECT 70.130 245.750 74.080 245.900 ;
        RECT 75.380 245.750 79.330 245.900 ;
        RECT 70.130 245.300 70.730 245.750 ;
        RECT 78.730 245.300 79.330 245.750 ;
        RECT 70.130 245.150 74.080 245.300 ;
        RECT 75.380 245.150 79.330 245.300 ;
        RECT 70.130 244.700 70.730 245.150 ;
        RECT 78.730 244.700 79.330 245.150 ;
        RECT 70.130 244.550 74.080 244.700 ;
        RECT 75.380 244.550 79.330 244.700 ;
        RECT 70.130 244.100 70.730 244.550 ;
        RECT 78.730 244.100 79.330 244.550 ;
        RECT 70.130 243.950 74.080 244.100 ;
        RECT 75.380 243.950 79.330 244.100 ;
        RECT 70.130 243.500 70.730 243.950 ;
        RECT 78.730 243.500 79.330 243.950 ;
        RECT 70.130 243.350 74.080 243.500 ;
        RECT 75.380 243.350 79.330 243.500 ;
        RECT 70.130 242.900 70.730 243.350 ;
        RECT 78.730 242.900 79.330 243.350 ;
        RECT 70.130 242.750 74.080 242.900 ;
        RECT 75.380 242.750 79.330 242.900 ;
        RECT 70.130 242.300 70.730 242.750 ;
        RECT 78.730 242.300 79.330 242.750 ;
        RECT 70.130 242.150 74.080 242.300 ;
        RECT 75.380 242.150 79.330 242.300 ;
        RECT 70.130 242.000 70.730 242.150 ;
        RECT 66.530 241.700 70.730 242.000 ;
        RECT 78.730 242.000 79.330 242.150 ;
        RECT 79.780 242.000 79.930 249.550 ;
        RECT 80.380 242.000 80.530 249.550 ;
        RECT 80.980 242.000 81.130 249.550 ;
        RECT 81.580 242.000 81.730 249.550 ;
        RECT 82.180 242.000 82.330 249.550 ;
        RECT 82.780 242.000 82.930 244.900 ;
        RECT 78.730 241.700 82.930 242.000 ;
        RECT 66.530 241.550 74.080 241.700 ;
        RECT 75.380 241.550 82.930 241.700 ;
        RECT 66.530 241.350 70.730 241.550 ;
        RECT 60.330 241.050 69.130 241.200 ;
        RECT 69.280 241.050 70.730 241.350 ;
        RECT 58.730 240.150 70.730 241.050 ;
        RECT 78.730 241.350 82.930 241.550 ;
        RECT 78.730 241.050 80.180 241.350 ;
        RECT 83.530 241.200 85.930 244.400 ;
        RECT 86.530 242.000 86.680 244.900 ;
        RECT 87.130 242.000 87.280 249.550 ;
        RECT 87.730 242.000 87.880 249.550 ;
        RECT 88.330 242.000 88.480 249.550 ;
        RECT 88.930 242.000 89.080 249.550 ;
        RECT 89.530 242.000 89.680 249.550 ;
        RECT 90.130 249.350 94.080 249.550 ;
        RECT 95.380 249.350 99.330 249.550 ;
        RECT 90.130 248.900 90.730 249.350 ;
        RECT 98.730 248.900 99.330 249.350 ;
        RECT 90.130 248.750 94.080 248.900 ;
        RECT 95.380 248.750 99.330 248.900 ;
        RECT 90.130 248.300 90.730 248.750 ;
        RECT 98.730 248.300 99.330 248.750 ;
        RECT 90.130 248.150 94.080 248.300 ;
        RECT 95.380 248.150 99.330 248.300 ;
        RECT 90.130 247.700 90.730 248.150 ;
        RECT 98.730 247.700 99.330 248.150 ;
        RECT 90.130 247.550 94.080 247.700 ;
        RECT 95.380 247.550 99.330 247.700 ;
        RECT 90.130 247.100 90.730 247.550 ;
        RECT 98.730 247.100 99.330 247.550 ;
        RECT 90.130 246.950 94.080 247.100 ;
        RECT 95.380 246.950 99.330 247.100 ;
        RECT 90.130 246.500 90.730 246.950 ;
        RECT 98.730 246.500 99.330 246.950 ;
        RECT 90.130 246.350 94.080 246.500 ;
        RECT 95.380 246.350 99.330 246.500 ;
        RECT 90.130 245.900 90.730 246.350 ;
        RECT 98.730 245.900 99.330 246.350 ;
        RECT 90.130 245.750 94.080 245.900 ;
        RECT 95.380 245.750 99.330 245.900 ;
        RECT 90.130 245.300 90.730 245.750 ;
        RECT 98.730 245.300 99.330 245.750 ;
        RECT 90.130 245.150 94.080 245.300 ;
        RECT 95.380 245.150 99.330 245.300 ;
        RECT 90.130 244.700 90.730 245.150 ;
        RECT 98.730 244.700 99.330 245.150 ;
        RECT 90.130 244.550 94.080 244.700 ;
        RECT 95.380 244.550 99.330 244.700 ;
        RECT 90.130 244.100 90.730 244.550 ;
        RECT 98.730 244.100 99.330 244.550 ;
        RECT 90.130 243.950 94.080 244.100 ;
        RECT 95.380 243.950 99.330 244.100 ;
        RECT 90.130 243.500 90.730 243.950 ;
        RECT 98.730 243.500 99.330 243.950 ;
        RECT 90.130 243.350 94.080 243.500 ;
        RECT 95.380 243.350 99.330 243.500 ;
        RECT 90.130 242.900 90.730 243.350 ;
        RECT 98.730 242.900 99.330 243.350 ;
        RECT 90.130 242.750 94.080 242.900 ;
        RECT 95.380 242.750 99.330 242.900 ;
        RECT 90.130 242.300 90.730 242.750 ;
        RECT 98.730 242.300 99.330 242.750 ;
        RECT 90.130 242.150 94.080 242.300 ;
        RECT 95.380 242.150 99.330 242.300 ;
        RECT 90.130 242.000 90.730 242.150 ;
        RECT 86.530 241.700 90.730 242.000 ;
        RECT 98.730 242.000 99.330 242.150 ;
        RECT 99.780 242.000 99.930 249.550 ;
        RECT 100.380 242.000 100.530 249.550 ;
        RECT 100.980 242.000 101.130 249.550 ;
        RECT 101.580 242.000 101.730 249.550 ;
        RECT 102.180 242.000 102.330 249.550 ;
        RECT 102.780 242.000 102.930 244.900 ;
        RECT 98.730 241.700 102.930 242.000 ;
        RECT 86.530 241.550 94.080 241.700 ;
        RECT 95.380 241.550 102.930 241.700 ;
        RECT 86.530 241.350 90.730 241.550 ;
        RECT 80.330 241.050 89.130 241.200 ;
        RECT 89.280 241.050 90.730 241.350 ;
        RECT 78.730 240.150 90.730 241.050 ;
        RECT 98.730 241.350 102.930 241.550 ;
        RECT 103.530 243.530 104.730 244.400 ;
        RECT 103.530 242.255 107.140 243.530 ;
        RECT 98.730 241.050 100.180 241.350 ;
        RECT 103.530 241.200 104.730 242.255 ;
        RECT 100.330 241.050 104.730 241.200 ;
        RECT 98.730 240.150 104.730 241.050 ;
        RECT 4.730 239.850 9.130 240.150 ;
        RECT 20.330 239.850 29.130 240.150 ;
        RECT 40.330 239.850 49.130 240.150 ;
        RECT 60.330 239.850 69.130 240.150 ;
        RECT 80.330 239.850 89.130 240.150 ;
        RECT 4.730 238.950 10.730 239.850 ;
        RECT 20.330 239.800 30.730 239.850 ;
        RECT 40.330 239.800 50.730 239.850 ;
        RECT 60.330 239.800 70.730 239.850 ;
        RECT 80.330 239.800 90.730 239.850 ;
        RECT 100.330 239.800 104.730 240.150 ;
        RECT 4.730 238.800 9.130 238.950 ;
        RECT 4.730 237.970 5.930 238.800 ;
        RECT 9.280 238.650 10.730 238.950 ;
        RECT 2.315 236.695 5.930 237.970 ;
        RECT 4.730 235.600 5.930 236.695 ;
        RECT 6.530 238.450 10.730 238.650 ;
        RECT 18.730 238.950 30.730 239.800 ;
        RECT 18.730 238.900 29.130 238.950 ;
        RECT 18.730 238.650 20.180 238.900 ;
        RECT 20.330 238.800 29.130 238.900 ;
        RECT 18.730 238.450 22.930 238.650 ;
        RECT 6.530 238.300 14.080 238.450 ;
        RECT 15.430 238.300 22.930 238.450 ;
        RECT 6.530 238.000 10.730 238.300 ;
        RECT 2.315 233.250 4.315 235.545 ;
        RECT 6.530 235.150 6.680 238.000 ;
        RECT 7.130 230.450 7.280 238.000 ;
        RECT 7.730 230.450 7.880 238.000 ;
        RECT 8.330 230.450 8.480 238.000 ;
        RECT 8.930 230.450 9.080 238.000 ;
        RECT 9.530 230.450 9.680 238.000 ;
        RECT 10.130 237.850 10.730 238.000 ;
        RECT 18.730 238.000 22.930 238.300 ;
        RECT 18.730 237.850 19.330 238.000 ;
        RECT 10.130 237.700 14.080 237.850 ;
        RECT 15.380 237.700 19.330 237.850 ;
        RECT 10.130 237.250 10.730 237.700 ;
        RECT 18.730 237.250 19.330 237.700 ;
        RECT 10.130 237.100 14.080 237.250 ;
        RECT 15.380 237.100 19.330 237.250 ;
        RECT 10.130 236.650 10.730 237.100 ;
        RECT 18.730 236.650 19.330 237.100 ;
        RECT 10.130 236.500 14.080 236.650 ;
        RECT 15.380 236.500 19.330 236.650 ;
        RECT 10.130 236.050 10.730 236.500 ;
        RECT 18.730 236.050 19.330 236.500 ;
        RECT 10.130 235.900 14.080 236.050 ;
        RECT 15.380 235.900 19.330 236.050 ;
        RECT 10.130 235.450 10.730 235.900 ;
        RECT 18.730 235.450 19.330 235.900 ;
        RECT 10.130 235.300 14.080 235.450 ;
        RECT 15.380 235.300 19.330 235.450 ;
        RECT 10.130 234.850 10.730 235.300 ;
        RECT 18.730 234.850 19.330 235.300 ;
        RECT 10.130 234.700 14.080 234.850 ;
        RECT 15.380 234.700 19.330 234.850 ;
        RECT 10.130 234.250 10.730 234.700 ;
        RECT 18.730 234.250 19.330 234.700 ;
        RECT 10.130 234.100 14.080 234.250 ;
        RECT 15.380 234.100 19.330 234.250 ;
        RECT 10.130 233.650 10.730 234.100 ;
        RECT 18.730 233.650 19.330 234.100 ;
        RECT 10.130 233.500 14.080 233.650 ;
        RECT 15.380 233.500 19.330 233.650 ;
        RECT 10.130 233.050 10.730 233.500 ;
        RECT 18.730 233.050 19.330 233.500 ;
        RECT 10.130 232.900 14.080 233.050 ;
        RECT 15.380 232.900 19.330 233.050 ;
        RECT 10.130 232.450 10.730 232.900 ;
        RECT 18.730 232.450 19.330 232.900 ;
        RECT 10.130 232.300 14.080 232.450 ;
        RECT 15.380 232.300 19.330 232.450 ;
        RECT 10.130 231.850 10.730 232.300 ;
        RECT 18.730 231.850 19.330 232.300 ;
        RECT 10.130 231.700 14.080 231.850 ;
        RECT 15.380 231.700 19.330 231.850 ;
        RECT 10.130 231.250 10.730 231.700 ;
        RECT 18.730 231.250 19.330 231.700 ;
        RECT 10.130 231.100 14.080 231.250 ;
        RECT 15.380 231.100 19.330 231.250 ;
        RECT 10.130 230.650 10.730 231.100 ;
        RECT 18.730 230.650 19.330 231.100 ;
        RECT 10.130 230.450 14.080 230.650 ;
        RECT 15.380 230.450 19.330 230.650 ;
        RECT 19.780 230.450 19.930 238.000 ;
        RECT 20.380 230.450 20.530 238.000 ;
        RECT 20.980 230.450 21.130 238.000 ;
        RECT 21.580 230.450 21.730 238.000 ;
        RECT 22.180 230.450 22.330 238.000 ;
        RECT 22.780 235.150 22.930 238.000 ;
        RECT 23.530 235.600 25.930 238.800 ;
        RECT 29.280 238.650 30.730 238.950 ;
        RECT 26.530 238.450 30.730 238.650 ;
        RECT 38.730 238.950 50.730 239.800 ;
        RECT 38.730 238.900 49.130 238.950 ;
        RECT 38.730 238.650 40.180 238.900 ;
        RECT 40.330 238.800 49.130 238.900 ;
        RECT 38.730 238.450 42.930 238.650 ;
        RECT 26.530 238.300 34.080 238.450 ;
        RECT 35.430 238.300 42.930 238.450 ;
        RECT 26.530 238.000 30.730 238.300 ;
        RECT 26.530 235.150 26.680 238.000 ;
        RECT 27.130 230.450 27.280 238.000 ;
        RECT 27.730 230.450 27.880 238.000 ;
        RECT 28.330 230.450 28.480 238.000 ;
        RECT 28.930 230.450 29.080 238.000 ;
        RECT 29.530 230.450 29.680 238.000 ;
        RECT 30.130 237.850 30.730 238.000 ;
        RECT 38.730 238.000 42.930 238.300 ;
        RECT 38.730 237.850 39.330 238.000 ;
        RECT 30.130 237.700 34.080 237.850 ;
        RECT 35.380 237.700 39.330 237.850 ;
        RECT 30.130 237.250 30.730 237.700 ;
        RECT 38.730 237.250 39.330 237.700 ;
        RECT 30.130 237.100 34.080 237.250 ;
        RECT 35.380 237.100 39.330 237.250 ;
        RECT 30.130 236.650 30.730 237.100 ;
        RECT 38.730 236.650 39.330 237.100 ;
        RECT 30.130 236.500 34.080 236.650 ;
        RECT 35.380 236.500 39.330 236.650 ;
        RECT 30.130 236.050 30.730 236.500 ;
        RECT 38.730 236.050 39.330 236.500 ;
        RECT 30.130 235.900 34.080 236.050 ;
        RECT 35.380 235.900 39.330 236.050 ;
        RECT 30.130 235.450 30.730 235.900 ;
        RECT 38.730 235.450 39.330 235.900 ;
        RECT 30.130 235.300 34.080 235.450 ;
        RECT 35.380 235.300 39.330 235.450 ;
        RECT 30.130 234.850 30.730 235.300 ;
        RECT 38.730 234.850 39.330 235.300 ;
        RECT 30.130 234.700 34.080 234.850 ;
        RECT 35.380 234.700 39.330 234.850 ;
        RECT 30.130 234.250 30.730 234.700 ;
        RECT 38.730 234.250 39.330 234.700 ;
        RECT 30.130 234.100 34.080 234.250 ;
        RECT 35.380 234.100 39.330 234.250 ;
        RECT 30.130 233.650 30.730 234.100 ;
        RECT 38.730 233.650 39.330 234.100 ;
        RECT 30.130 233.500 34.080 233.650 ;
        RECT 35.380 233.500 39.330 233.650 ;
        RECT 30.130 233.050 30.730 233.500 ;
        RECT 38.730 233.050 39.330 233.500 ;
        RECT 30.130 232.900 34.080 233.050 ;
        RECT 35.380 232.900 39.330 233.050 ;
        RECT 30.130 232.450 30.730 232.900 ;
        RECT 38.730 232.450 39.330 232.900 ;
        RECT 30.130 232.300 34.080 232.450 ;
        RECT 35.380 232.300 39.330 232.450 ;
        RECT 30.130 231.850 30.730 232.300 ;
        RECT 38.730 231.850 39.330 232.300 ;
        RECT 30.130 231.700 34.080 231.850 ;
        RECT 35.380 231.700 39.330 231.850 ;
        RECT 30.130 231.250 30.730 231.700 ;
        RECT 38.730 231.250 39.330 231.700 ;
        RECT 30.130 231.100 34.080 231.250 ;
        RECT 35.380 231.100 39.330 231.250 ;
        RECT 30.130 230.650 30.730 231.100 ;
        RECT 38.730 230.650 39.330 231.100 ;
        RECT 30.130 230.450 34.080 230.650 ;
        RECT 35.380 230.450 39.330 230.650 ;
        RECT 39.780 230.450 39.930 238.000 ;
        RECT 40.380 230.450 40.530 238.000 ;
        RECT 40.980 230.450 41.130 238.000 ;
        RECT 41.580 230.450 41.730 238.000 ;
        RECT 42.180 230.450 42.330 238.000 ;
        RECT 42.780 235.150 42.930 238.000 ;
        RECT 43.530 235.600 45.930 238.800 ;
        RECT 49.280 238.650 50.730 238.950 ;
        RECT 46.530 238.450 50.730 238.650 ;
        RECT 58.730 238.950 70.730 239.800 ;
        RECT 58.730 238.900 69.130 238.950 ;
        RECT 58.730 238.650 60.180 238.900 ;
        RECT 60.330 238.800 69.130 238.900 ;
        RECT 58.730 238.450 62.930 238.650 ;
        RECT 46.530 238.300 54.080 238.450 ;
        RECT 55.430 238.300 62.930 238.450 ;
        RECT 46.530 238.000 50.730 238.300 ;
        RECT 46.530 235.150 46.680 238.000 ;
        RECT 47.130 230.450 47.280 238.000 ;
        RECT 47.730 230.450 47.880 238.000 ;
        RECT 48.330 230.450 48.480 238.000 ;
        RECT 48.930 230.450 49.080 238.000 ;
        RECT 49.530 230.450 49.680 238.000 ;
        RECT 50.130 237.850 50.730 238.000 ;
        RECT 58.730 238.000 62.930 238.300 ;
        RECT 58.730 237.850 59.330 238.000 ;
        RECT 50.130 237.700 54.080 237.850 ;
        RECT 55.380 237.700 59.330 237.850 ;
        RECT 50.130 237.250 50.730 237.700 ;
        RECT 58.730 237.250 59.330 237.700 ;
        RECT 50.130 237.100 54.080 237.250 ;
        RECT 55.380 237.100 59.330 237.250 ;
        RECT 50.130 236.650 50.730 237.100 ;
        RECT 58.730 236.650 59.330 237.100 ;
        RECT 50.130 236.500 54.080 236.650 ;
        RECT 55.380 236.500 59.330 236.650 ;
        RECT 50.130 236.050 50.730 236.500 ;
        RECT 58.730 236.050 59.330 236.500 ;
        RECT 50.130 235.900 54.080 236.050 ;
        RECT 55.380 235.900 59.330 236.050 ;
        RECT 50.130 235.450 50.730 235.900 ;
        RECT 58.730 235.450 59.330 235.900 ;
        RECT 50.130 235.300 54.080 235.450 ;
        RECT 55.380 235.300 59.330 235.450 ;
        RECT 50.130 234.850 50.730 235.300 ;
        RECT 58.730 234.850 59.330 235.300 ;
        RECT 50.130 234.700 54.080 234.850 ;
        RECT 55.380 234.700 59.330 234.850 ;
        RECT 50.130 234.250 50.730 234.700 ;
        RECT 58.730 234.250 59.330 234.700 ;
        RECT 50.130 234.100 54.080 234.250 ;
        RECT 55.380 234.100 59.330 234.250 ;
        RECT 50.130 233.650 50.730 234.100 ;
        RECT 58.730 233.650 59.330 234.100 ;
        RECT 50.130 233.500 54.080 233.650 ;
        RECT 55.380 233.500 59.330 233.650 ;
        RECT 50.130 233.050 50.730 233.500 ;
        RECT 58.730 233.050 59.330 233.500 ;
        RECT 50.130 232.900 54.080 233.050 ;
        RECT 55.380 232.900 59.330 233.050 ;
        RECT 50.130 232.450 50.730 232.900 ;
        RECT 58.730 232.450 59.330 232.900 ;
        RECT 50.130 232.300 54.080 232.450 ;
        RECT 55.380 232.300 59.330 232.450 ;
        RECT 50.130 231.850 50.730 232.300 ;
        RECT 58.730 231.850 59.330 232.300 ;
        RECT 50.130 231.700 54.080 231.850 ;
        RECT 55.380 231.700 59.330 231.850 ;
        RECT 50.130 231.250 50.730 231.700 ;
        RECT 58.730 231.250 59.330 231.700 ;
        RECT 50.130 231.100 54.080 231.250 ;
        RECT 55.380 231.100 59.330 231.250 ;
        RECT 50.130 230.650 50.730 231.100 ;
        RECT 58.730 230.650 59.330 231.100 ;
        RECT 50.130 230.450 54.080 230.650 ;
        RECT 55.380 230.450 59.330 230.650 ;
        RECT 59.780 230.450 59.930 238.000 ;
        RECT 60.380 230.450 60.530 238.000 ;
        RECT 60.980 230.450 61.130 238.000 ;
        RECT 61.580 230.450 61.730 238.000 ;
        RECT 62.180 230.450 62.330 238.000 ;
        RECT 62.780 235.150 62.930 238.000 ;
        RECT 63.530 235.600 65.930 238.800 ;
        RECT 69.280 238.650 70.730 238.950 ;
        RECT 66.530 238.450 70.730 238.650 ;
        RECT 78.730 238.950 90.730 239.800 ;
        RECT 78.730 238.900 89.130 238.950 ;
        RECT 78.730 238.650 80.180 238.900 ;
        RECT 80.330 238.800 89.130 238.900 ;
        RECT 78.730 238.450 82.930 238.650 ;
        RECT 66.530 238.300 74.080 238.450 ;
        RECT 75.430 238.300 82.930 238.450 ;
        RECT 66.530 238.000 70.730 238.300 ;
        RECT 66.530 235.150 66.680 238.000 ;
        RECT 67.130 230.450 67.280 238.000 ;
        RECT 67.730 230.450 67.880 238.000 ;
        RECT 68.330 230.450 68.480 238.000 ;
        RECT 68.930 230.450 69.080 238.000 ;
        RECT 69.530 230.450 69.680 238.000 ;
        RECT 70.130 237.850 70.730 238.000 ;
        RECT 78.730 238.000 82.930 238.300 ;
        RECT 78.730 237.850 79.330 238.000 ;
        RECT 70.130 237.700 74.080 237.850 ;
        RECT 75.380 237.700 79.330 237.850 ;
        RECT 70.130 237.250 70.730 237.700 ;
        RECT 78.730 237.250 79.330 237.700 ;
        RECT 70.130 237.100 74.080 237.250 ;
        RECT 75.380 237.100 79.330 237.250 ;
        RECT 70.130 236.650 70.730 237.100 ;
        RECT 78.730 236.650 79.330 237.100 ;
        RECT 70.130 236.500 74.080 236.650 ;
        RECT 75.380 236.500 79.330 236.650 ;
        RECT 70.130 236.050 70.730 236.500 ;
        RECT 78.730 236.050 79.330 236.500 ;
        RECT 70.130 235.900 74.080 236.050 ;
        RECT 75.380 235.900 79.330 236.050 ;
        RECT 70.130 235.450 70.730 235.900 ;
        RECT 78.730 235.450 79.330 235.900 ;
        RECT 70.130 235.300 74.080 235.450 ;
        RECT 75.380 235.300 79.330 235.450 ;
        RECT 70.130 234.850 70.730 235.300 ;
        RECT 78.730 234.850 79.330 235.300 ;
        RECT 70.130 234.700 74.080 234.850 ;
        RECT 75.380 234.700 79.330 234.850 ;
        RECT 70.130 234.250 70.730 234.700 ;
        RECT 78.730 234.250 79.330 234.700 ;
        RECT 70.130 234.100 74.080 234.250 ;
        RECT 75.380 234.100 79.330 234.250 ;
        RECT 70.130 233.650 70.730 234.100 ;
        RECT 78.730 233.650 79.330 234.100 ;
        RECT 70.130 233.500 74.080 233.650 ;
        RECT 75.380 233.500 79.330 233.650 ;
        RECT 70.130 233.050 70.730 233.500 ;
        RECT 78.730 233.050 79.330 233.500 ;
        RECT 70.130 232.900 74.080 233.050 ;
        RECT 75.380 232.900 79.330 233.050 ;
        RECT 70.130 232.450 70.730 232.900 ;
        RECT 78.730 232.450 79.330 232.900 ;
        RECT 70.130 232.300 74.080 232.450 ;
        RECT 75.380 232.300 79.330 232.450 ;
        RECT 70.130 231.850 70.730 232.300 ;
        RECT 78.730 231.850 79.330 232.300 ;
        RECT 70.130 231.700 74.080 231.850 ;
        RECT 75.380 231.700 79.330 231.850 ;
        RECT 70.130 231.250 70.730 231.700 ;
        RECT 78.730 231.250 79.330 231.700 ;
        RECT 70.130 231.100 74.080 231.250 ;
        RECT 75.380 231.100 79.330 231.250 ;
        RECT 70.130 230.650 70.730 231.100 ;
        RECT 78.730 230.650 79.330 231.100 ;
        RECT 70.130 230.450 74.080 230.650 ;
        RECT 75.380 230.450 79.330 230.650 ;
        RECT 79.780 230.450 79.930 238.000 ;
        RECT 80.380 230.450 80.530 238.000 ;
        RECT 80.980 230.450 81.130 238.000 ;
        RECT 81.580 230.450 81.730 238.000 ;
        RECT 82.180 230.450 82.330 238.000 ;
        RECT 82.780 235.150 82.930 238.000 ;
        RECT 83.530 235.600 85.930 238.800 ;
        RECT 89.280 238.650 90.730 238.950 ;
        RECT 86.530 238.450 90.730 238.650 ;
        RECT 98.730 238.900 104.730 239.800 ;
        RECT 98.730 238.650 100.180 238.900 ;
        RECT 100.330 238.800 104.730 238.900 ;
        RECT 98.730 238.450 102.930 238.650 ;
        RECT 86.530 238.300 94.080 238.450 ;
        RECT 95.430 238.300 102.930 238.450 ;
        RECT 86.530 238.000 90.730 238.300 ;
        RECT 86.530 235.150 86.680 238.000 ;
        RECT 87.130 230.450 87.280 238.000 ;
        RECT 87.730 230.450 87.880 238.000 ;
        RECT 88.330 230.450 88.480 238.000 ;
        RECT 88.930 230.450 89.080 238.000 ;
        RECT 89.530 230.450 89.680 238.000 ;
        RECT 90.130 237.850 90.730 238.000 ;
        RECT 98.730 238.000 102.930 238.300 ;
        RECT 98.730 237.850 99.330 238.000 ;
        RECT 90.130 237.700 94.080 237.850 ;
        RECT 95.380 237.700 99.330 237.850 ;
        RECT 90.130 237.250 90.730 237.700 ;
        RECT 98.730 237.250 99.330 237.700 ;
        RECT 90.130 237.100 94.080 237.250 ;
        RECT 95.380 237.100 99.330 237.250 ;
        RECT 90.130 236.650 90.730 237.100 ;
        RECT 98.730 236.650 99.330 237.100 ;
        RECT 90.130 236.500 94.080 236.650 ;
        RECT 95.380 236.500 99.330 236.650 ;
        RECT 90.130 236.050 90.730 236.500 ;
        RECT 98.730 236.050 99.330 236.500 ;
        RECT 90.130 235.900 94.080 236.050 ;
        RECT 95.380 235.900 99.330 236.050 ;
        RECT 90.130 235.450 90.730 235.900 ;
        RECT 98.730 235.450 99.330 235.900 ;
        RECT 90.130 235.300 94.080 235.450 ;
        RECT 95.380 235.300 99.330 235.450 ;
        RECT 90.130 234.850 90.730 235.300 ;
        RECT 98.730 234.850 99.330 235.300 ;
        RECT 90.130 234.700 94.080 234.850 ;
        RECT 95.380 234.700 99.330 234.850 ;
        RECT 90.130 234.250 90.730 234.700 ;
        RECT 98.730 234.250 99.330 234.700 ;
        RECT 90.130 234.100 94.080 234.250 ;
        RECT 95.380 234.100 99.330 234.250 ;
        RECT 90.130 233.650 90.730 234.100 ;
        RECT 98.730 233.650 99.330 234.100 ;
        RECT 90.130 233.500 94.080 233.650 ;
        RECT 95.380 233.500 99.330 233.650 ;
        RECT 90.130 233.050 90.730 233.500 ;
        RECT 98.730 233.050 99.330 233.500 ;
        RECT 90.130 232.900 94.080 233.050 ;
        RECT 95.380 232.900 99.330 233.050 ;
        RECT 90.130 232.450 90.730 232.900 ;
        RECT 98.730 232.450 99.330 232.900 ;
        RECT 90.130 232.300 94.080 232.450 ;
        RECT 95.380 232.300 99.330 232.450 ;
        RECT 90.130 231.850 90.730 232.300 ;
        RECT 98.730 231.850 99.330 232.300 ;
        RECT 90.130 231.700 94.080 231.850 ;
        RECT 95.380 231.700 99.330 231.850 ;
        RECT 90.130 231.250 90.730 231.700 ;
        RECT 98.730 231.250 99.330 231.700 ;
        RECT 90.130 231.100 94.080 231.250 ;
        RECT 95.380 231.100 99.330 231.250 ;
        RECT 90.130 230.650 90.730 231.100 ;
        RECT 98.730 230.650 99.330 231.100 ;
        RECT 90.130 230.450 94.080 230.650 ;
        RECT 95.380 230.450 99.330 230.650 ;
        RECT 99.780 230.450 99.930 238.000 ;
        RECT 100.380 230.450 100.530 238.000 ;
        RECT 100.980 230.450 101.130 238.000 ;
        RECT 101.580 230.450 101.730 238.000 ;
        RECT 102.180 230.450 102.330 238.000 ;
        RECT 102.780 235.150 102.930 238.000 ;
        RECT 103.530 237.765 104.730 238.800 ;
        RECT 103.530 236.490 107.140 237.765 ;
        RECT 103.530 235.600 104.730 236.490 ;
        RECT 2.315 224.455 4.315 226.750 ;
        RECT 2.315 224.450 4.180 224.455 ;
        RECT 4.730 222.670 5.930 224.400 ;
        RECT 2.315 221.395 5.930 222.670 ;
        RECT 4.730 221.200 5.930 221.395 ;
        RECT 6.530 222.000 6.680 224.900 ;
        RECT 7.130 222.000 7.280 229.550 ;
        RECT 7.730 222.000 7.880 229.550 ;
        RECT 8.330 222.000 8.480 229.550 ;
        RECT 8.930 222.000 9.080 229.550 ;
        RECT 9.530 222.000 9.680 229.550 ;
        RECT 10.130 229.350 14.080 229.550 ;
        RECT 15.380 229.350 19.330 229.550 ;
        RECT 10.130 228.900 10.730 229.350 ;
        RECT 18.730 228.900 19.330 229.350 ;
        RECT 10.130 228.750 14.080 228.900 ;
        RECT 15.380 228.750 19.330 228.900 ;
        RECT 10.130 228.300 10.730 228.750 ;
        RECT 18.730 228.300 19.330 228.750 ;
        RECT 10.130 228.150 14.080 228.300 ;
        RECT 15.380 228.150 19.330 228.300 ;
        RECT 10.130 227.700 10.730 228.150 ;
        RECT 18.730 227.700 19.330 228.150 ;
        RECT 10.130 227.550 14.080 227.700 ;
        RECT 15.380 227.550 19.330 227.700 ;
        RECT 10.130 227.100 10.730 227.550 ;
        RECT 18.730 227.100 19.330 227.550 ;
        RECT 10.130 226.950 14.080 227.100 ;
        RECT 15.380 226.950 19.330 227.100 ;
        RECT 10.130 226.500 10.730 226.950 ;
        RECT 18.730 226.500 19.330 226.950 ;
        RECT 10.130 226.350 14.080 226.500 ;
        RECT 15.380 226.350 19.330 226.500 ;
        RECT 10.130 225.900 10.730 226.350 ;
        RECT 18.730 225.900 19.330 226.350 ;
        RECT 10.130 225.750 14.080 225.900 ;
        RECT 15.380 225.750 19.330 225.900 ;
        RECT 10.130 225.300 10.730 225.750 ;
        RECT 18.730 225.300 19.330 225.750 ;
        RECT 10.130 225.150 14.080 225.300 ;
        RECT 15.380 225.150 19.330 225.300 ;
        RECT 10.130 224.700 10.730 225.150 ;
        RECT 18.730 224.700 19.330 225.150 ;
        RECT 10.130 224.550 14.080 224.700 ;
        RECT 15.380 224.550 19.330 224.700 ;
        RECT 10.130 224.100 10.730 224.550 ;
        RECT 18.730 224.100 19.330 224.550 ;
        RECT 10.130 223.950 14.080 224.100 ;
        RECT 15.380 223.950 19.330 224.100 ;
        RECT 10.130 223.500 10.730 223.950 ;
        RECT 18.730 223.500 19.330 223.950 ;
        RECT 10.130 223.350 14.080 223.500 ;
        RECT 15.380 223.350 19.330 223.500 ;
        RECT 10.130 222.900 10.730 223.350 ;
        RECT 18.730 222.900 19.330 223.350 ;
        RECT 10.130 222.750 14.080 222.900 ;
        RECT 15.380 222.750 19.330 222.900 ;
        RECT 10.130 222.300 10.730 222.750 ;
        RECT 18.730 222.300 19.330 222.750 ;
        RECT 10.130 222.150 14.080 222.300 ;
        RECT 15.380 222.150 19.330 222.300 ;
        RECT 10.130 222.000 10.730 222.150 ;
        RECT 6.530 221.700 10.730 222.000 ;
        RECT 18.730 222.000 19.330 222.150 ;
        RECT 19.780 222.000 19.930 229.550 ;
        RECT 20.380 222.000 20.530 229.550 ;
        RECT 20.980 222.000 21.130 229.550 ;
        RECT 21.580 222.000 21.730 229.550 ;
        RECT 22.180 222.000 22.330 229.550 ;
        RECT 22.780 222.000 22.930 224.900 ;
        RECT 18.730 221.700 22.930 222.000 ;
        RECT 6.530 221.550 14.080 221.700 ;
        RECT 15.380 221.550 22.930 221.700 ;
        RECT 6.530 221.350 10.730 221.550 ;
        RECT 4.730 221.050 9.130 221.200 ;
        RECT 9.280 221.050 10.730 221.350 ;
        RECT 4.730 220.150 10.730 221.050 ;
        RECT 18.730 221.350 22.930 221.550 ;
        RECT 18.730 221.050 20.180 221.350 ;
        RECT 23.530 221.200 25.930 224.400 ;
        RECT 26.530 222.000 26.680 224.900 ;
        RECT 27.130 222.000 27.280 229.550 ;
        RECT 27.730 222.000 27.880 229.550 ;
        RECT 28.330 222.000 28.480 229.550 ;
        RECT 28.930 222.000 29.080 229.550 ;
        RECT 29.530 222.000 29.680 229.550 ;
        RECT 30.130 229.350 34.080 229.550 ;
        RECT 35.380 229.350 39.330 229.550 ;
        RECT 30.130 228.900 30.730 229.350 ;
        RECT 38.730 228.900 39.330 229.350 ;
        RECT 30.130 228.750 34.080 228.900 ;
        RECT 35.380 228.750 39.330 228.900 ;
        RECT 30.130 228.300 30.730 228.750 ;
        RECT 38.730 228.300 39.330 228.750 ;
        RECT 30.130 228.150 34.080 228.300 ;
        RECT 35.380 228.150 39.330 228.300 ;
        RECT 30.130 227.700 30.730 228.150 ;
        RECT 38.730 227.700 39.330 228.150 ;
        RECT 30.130 227.550 34.080 227.700 ;
        RECT 35.380 227.550 39.330 227.700 ;
        RECT 30.130 227.100 30.730 227.550 ;
        RECT 38.730 227.100 39.330 227.550 ;
        RECT 30.130 226.950 34.080 227.100 ;
        RECT 35.380 226.950 39.330 227.100 ;
        RECT 30.130 226.500 30.730 226.950 ;
        RECT 38.730 226.500 39.330 226.950 ;
        RECT 30.130 226.350 34.080 226.500 ;
        RECT 35.380 226.350 39.330 226.500 ;
        RECT 30.130 225.900 30.730 226.350 ;
        RECT 38.730 225.900 39.330 226.350 ;
        RECT 30.130 225.750 34.080 225.900 ;
        RECT 35.380 225.750 39.330 225.900 ;
        RECT 30.130 225.300 30.730 225.750 ;
        RECT 38.730 225.300 39.330 225.750 ;
        RECT 30.130 225.150 34.080 225.300 ;
        RECT 35.380 225.150 39.330 225.300 ;
        RECT 30.130 224.700 30.730 225.150 ;
        RECT 38.730 224.700 39.330 225.150 ;
        RECT 30.130 224.550 34.080 224.700 ;
        RECT 35.380 224.550 39.330 224.700 ;
        RECT 30.130 224.100 30.730 224.550 ;
        RECT 38.730 224.100 39.330 224.550 ;
        RECT 30.130 223.950 34.080 224.100 ;
        RECT 35.380 223.950 39.330 224.100 ;
        RECT 30.130 223.500 30.730 223.950 ;
        RECT 38.730 223.500 39.330 223.950 ;
        RECT 30.130 223.350 34.080 223.500 ;
        RECT 35.380 223.350 39.330 223.500 ;
        RECT 30.130 222.900 30.730 223.350 ;
        RECT 38.730 222.900 39.330 223.350 ;
        RECT 30.130 222.750 34.080 222.900 ;
        RECT 35.380 222.750 39.330 222.900 ;
        RECT 30.130 222.300 30.730 222.750 ;
        RECT 38.730 222.300 39.330 222.750 ;
        RECT 30.130 222.150 34.080 222.300 ;
        RECT 35.380 222.150 39.330 222.300 ;
        RECT 30.130 222.000 30.730 222.150 ;
        RECT 26.530 221.700 30.730 222.000 ;
        RECT 38.730 222.000 39.330 222.150 ;
        RECT 39.780 222.000 39.930 229.550 ;
        RECT 40.380 222.000 40.530 229.550 ;
        RECT 40.980 222.000 41.130 229.550 ;
        RECT 41.580 222.000 41.730 229.550 ;
        RECT 42.180 222.000 42.330 229.550 ;
        RECT 42.780 222.000 42.930 224.900 ;
        RECT 38.730 221.700 42.930 222.000 ;
        RECT 26.530 221.550 34.080 221.700 ;
        RECT 35.380 221.550 42.930 221.700 ;
        RECT 26.530 221.350 30.730 221.550 ;
        RECT 20.330 221.050 29.130 221.200 ;
        RECT 29.280 221.050 30.730 221.350 ;
        RECT 18.730 220.150 30.730 221.050 ;
        RECT 38.730 221.350 42.930 221.550 ;
        RECT 38.730 221.050 40.180 221.350 ;
        RECT 43.530 221.200 45.930 224.400 ;
        RECT 46.530 222.000 46.680 224.900 ;
        RECT 47.130 222.000 47.280 229.550 ;
        RECT 47.730 222.000 47.880 229.550 ;
        RECT 48.330 222.000 48.480 229.550 ;
        RECT 48.930 222.000 49.080 229.550 ;
        RECT 49.530 222.000 49.680 229.550 ;
        RECT 50.130 229.350 54.080 229.550 ;
        RECT 55.380 229.350 59.330 229.550 ;
        RECT 50.130 228.900 50.730 229.350 ;
        RECT 58.730 228.900 59.330 229.350 ;
        RECT 50.130 228.750 54.080 228.900 ;
        RECT 55.380 228.750 59.330 228.900 ;
        RECT 50.130 228.300 50.730 228.750 ;
        RECT 58.730 228.300 59.330 228.750 ;
        RECT 50.130 228.150 54.080 228.300 ;
        RECT 55.380 228.150 59.330 228.300 ;
        RECT 50.130 227.700 50.730 228.150 ;
        RECT 58.730 227.700 59.330 228.150 ;
        RECT 50.130 227.550 54.080 227.700 ;
        RECT 55.380 227.550 59.330 227.700 ;
        RECT 50.130 227.100 50.730 227.550 ;
        RECT 58.730 227.100 59.330 227.550 ;
        RECT 50.130 226.950 54.080 227.100 ;
        RECT 55.380 226.950 59.330 227.100 ;
        RECT 50.130 226.500 50.730 226.950 ;
        RECT 58.730 226.500 59.330 226.950 ;
        RECT 50.130 226.350 54.080 226.500 ;
        RECT 55.380 226.350 59.330 226.500 ;
        RECT 50.130 225.900 50.730 226.350 ;
        RECT 58.730 225.900 59.330 226.350 ;
        RECT 50.130 225.750 54.080 225.900 ;
        RECT 55.380 225.750 59.330 225.900 ;
        RECT 50.130 225.300 50.730 225.750 ;
        RECT 58.730 225.300 59.330 225.750 ;
        RECT 50.130 225.150 54.080 225.300 ;
        RECT 55.380 225.150 59.330 225.300 ;
        RECT 50.130 224.700 50.730 225.150 ;
        RECT 58.730 224.700 59.330 225.150 ;
        RECT 50.130 224.550 54.080 224.700 ;
        RECT 55.380 224.550 59.330 224.700 ;
        RECT 50.130 224.100 50.730 224.550 ;
        RECT 58.730 224.100 59.330 224.550 ;
        RECT 50.130 223.950 54.080 224.100 ;
        RECT 55.380 223.950 59.330 224.100 ;
        RECT 50.130 223.500 50.730 223.950 ;
        RECT 58.730 223.500 59.330 223.950 ;
        RECT 50.130 223.350 54.080 223.500 ;
        RECT 55.380 223.350 59.330 223.500 ;
        RECT 50.130 222.900 50.730 223.350 ;
        RECT 58.730 222.900 59.330 223.350 ;
        RECT 50.130 222.750 54.080 222.900 ;
        RECT 55.380 222.750 59.330 222.900 ;
        RECT 50.130 222.300 50.730 222.750 ;
        RECT 58.730 222.300 59.330 222.750 ;
        RECT 50.130 222.150 54.080 222.300 ;
        RECT 55.380 222.150 59.330 222.300 ;
        RECT 50.130 222.000 50.730 222.150 ;
        RECT 46.530 221.700 50.730 222.000 ;
        RECT 58.730 222.000 59.330 222.150 ;
        RECT 59.780 222.000 59.930 229.550 ;
        RECT 60.380 222.000 60.530 229.550 ;
        RECT 60.980 222.000 61.130 229.550 ;
        RECT 61.580 222.000 61.730 229.550 ;
        RECT 62.180 222.000 62.330 229.550 ;
        RECT 62.780 222.000 62.930 224.900 ;
        RECT 58.730 221.700 62.930 222.000 ;
        RECT 46.530 221.550 54.080 221.700 ;
        RECT 55.380 221.550 62.930 221.700 ;
        RECT 46.530 221.350 50.730 221.550 ;
        RECT 40.330 221.050 49.130 221.200 ;
        RECT 49.280 221.050 50.730 221.350 ;
        RECT 38.730 220.150 50.730 221.050 ;
        RECT 58.730 221.350 62.930 221.550 ;
        RECT 58.730 221.050 60.180 221.350 ;
        RECT 63.530 221.200 65.930 224.400 ;
        RECT 66.530 222.000 66.680 224.900 ;
        RECT 67.130 222.000 67.280 229.550 ;
        RECT 67.730 222.000 67.880 229.550 ;
        RECT 68.330 222.000 68.480 229.550 ;
        RECT 68.930 222.000 69.080 229.550 ;
        RECT 69.530 222.000 69.680 229.550 ;
        RECT 70.130 229.350 74.080 229.550 ;
        RECT 75.380 229.350 79.330 229.550 ;
        RECT 70.130 228.900 70.730 229.350 ;
        RECT 78.730 228.900 79.330 229.350 ;
        RECT 70.130 228.750 74.080 228.900 ;
        RECT 75.380 228.750 79.330 228.900 ;
        RECT 70.130 228.300 70.730 228.750 ;
        RECT 78.730 228.300 79.330 228.750 ;
        RECT 70.130 228.150 74.080 228.300 ;
        RECT 75.380 228.150 79.330 228.300 ;
        RECT 70.130 227.700 70.730 228.150 ;
        RECT 78.730 227.700 79.330 228.150 ;
        RECT 70.130 227.550 74.080 227.700 ;
        RECT 75.380 227.550 79.330 227.700 ;
        RECT 70.130 227.100 70.730 227.550 ;
        RECT 78.730 227.100 79.330 227.550 ;
        RECT 70.130 226.950 74.080 227.100 ;
        RECT 75.380 226.950 79.330 227.100 ;
        RECT 70.130 226.500 70.730 226.950 ;
        RECT 78.730 226.500 79.330 226.950 ;
        RECT 70.130 226.350 74.080 226.500 ;
        RECT 75.380 226.350 79.330 226.500 ;
        RECT 70.130 225.900 70.730 226.350 ;
        RECT 78.730 225.900 79.330 226.350 ;
        RECT 70.130 225.750 74.080 225.900 ;
        RECT 75.380 225.750 79.330 225.900 ;
        RECT 70.130 225.300 70.730 225.750 ;
        RECT 78.730 225.300 79.330 225.750 ;
        RECT 70.130 225.150 74.080 225.300 ;
        RECT 75.380 225.150 79.330 225.300 ;
        RECT 70.130 224.700 70.730 225.150 ;
        RECT 78.730 224.700 79.330 225.150 ;
        RECT 70.130 224.550 74.080 224.700 ;
        RECT 75.380 224.550 79.330 224.700 ;
        RECT 70.130 224.100 70.730 224.550 ;
        RECT 78.730 224.100 79.330 224.550 ;
        RECT 70.130 223.950 74.080 224.100 ;
        RECT 75.380 223.950 79.330 224.100 ;
        RECT 70.130 223.500 70.730 223.950 ;
        RECT 78.730 223.500 79.330 223.950 ;
        RECT 70.130 223.350 74.080 223.500 ;
        RECT 75.380 223.350 79.330 223.500 ;
        RECT 70.130 222.900 70.730 223.350 ;
        RECT 78.730 222.900 79.330 223.350 ;
        RECT 70.130 222.750 74.080 222.900 ;
        RECT 75.380 222.750 79.330 222.900 ;
        RECT 70.130 222.300 70.730 222.750 ;
        RECT 78.730 222.300 79.330 222.750 ;
        RECT 70.130 222.150 74.080 222.300 ;
        RECT 75.380 222.150 79.330 222.300 ;
        RECT 70.130 222.000 70.730 222.150 ;
        RECT 66.530 221.700 70.730 222.000 ;
        RECT 78.730 222.000 79.330 222.150 ;
        RECT 79.780 222.000 79.930 229.550 ;
        RECT 80.380 222.000 80.530 229.550 ;
        RECT 80.980 222.000 81.130 229.550 ;
        RECT 81.580 222.000 81.730 229.550 ;
        RECT 82.180 222.000 82.330 229.550 ;
        RECT 82.780 222.000 82.930 224.900 ;
        RECT 78.730 221.700 82.930 222.000 ;
        RECT 66.530 221.550 74.080 221.700 ;
        RECT 75.380 221.550 82.930 221.700 ;
        RECT 66.530 221.350 70.730 221.550 ;
        RECT 60.330 221.050 69.130 221.200 ;
        RECT 69.280 221.050 70.730 221.350 ;
        RECT 58.730 220.150 70.730 221.050 ;
        RECT 78.730 221.350 82.930 221.550 ;
        RECT 78.730 221.050 80.180 221.350 ;
        RECT 83.530 221.200 85.930 224.400 ;
        RECT 86.530 222.000 86.680 224.900 ;
        RECT 87.130 222.000 87.280 229.550 ;
        RECT 87.730 222.000 87.880 229.550 ;
        RECT 88.330 222.000 88.480 229.550 ;
        RECT 88.930 222.000 89.080 229.550 ;
        RECT 89.530 222.000 89.680 229.550 ;
        RECT 90.130 229.350 94.080 229.550 ;
        RECT 95.380 229.350 99.330 229.550 ;
        RECT 90.130 228.900 90.730 229.350 ;
        RECT 98.730 228.900 99.330 229.350 ;
        RECT 90.130 228.750 94.080 228.900 ;
        RECT 95.380 228.750 99.330 228.900 ;
        RECT 90.130 228.300 90.730 228.750 ;
        RECT 98.730 228.300 99.330 228.750 ;
        RECT 90.130 228.150 94.080 228.300 ;
        RECT 95.380 228.150 99.330 228.300 ;
        RECT 90.130 227.700 90.730 228.150 ;
        RECT 98.730 227.700 99.330 228.150 ;
        RECT 90.130 227.550 94.080 227.700 ;
        RECT 95.380 227.550 99.330 227.700 ;
        RECT 90.130 227.100 90.730 227.550 ;
        RECT 98.730 227.100 99.330 227.550 ;
        RECT 90.130 226.950 94.080 227.100 ;
        RECT 95.380 226.950 99.330 227.100 ;
        RECT 90.130 226.500 90.730 226.950 ;
        RECT 98.730 226.500 99.330 226.950 ;
        RECT 90.130 226.350 94.080 226.500 ;
        RECT 95.380 226.350 99.330 226.500 ;
        RECT 90.130 225.900 90.730 226.350 ;
        RECT 98.730 225.900 99.330 226.350 ;
        RECT 90.130 225.750 94.080 225.900 ;
        RECT 95.380 225.750 99.330 225.900 ;
        RECT 90.130 225.300 90.730 225.750 ;
        RECT 98.730 225.300 99.330 225.750 ;
        RECT 90.130 225.150 94.080 225.300 ;
        RECT 95.380 225.150 99.330 225.300 ;
        RECT 90.130 224.700 90.730 225.150 ;
        RECT 98.730 224.700 99.330 225.150 ;
        RECT 90.130 224.550 94.080 224.700 ;
        RECT 95.380 224.550 99.330 224.700 ;
        RECT 90.130 224.100 90.730 224.550 ;
        RECT 98.730 224.100 99.330 224.550 ;
        RECT 90.130 223.950 94.080 224.100 ;
        RECT 95.380 223.950 99.330 224.100 ;
        RECT 90.130 223.500 90.730 223.950 ;
        RECT 98.730 223.500 99.330 223.950 ;
        RECT 90.130 223.350 94.080 223.500 ;
        RECT 95.380 223.350 99.330 223.500 ;
        RECT 90.130 222.900 90.730 223.350 ;
        RECT 98.730 222.900 99.330 223.350 ;
        RECT 90.130 222.750 94.080 222.900 ;
        RECT 95.380 222.750 99.330 222.900 ;
        RECT 90.130 222.300 90.730 222.750 ;
        RECT 98.730 222.300 99.330 222.750 ;
        RECT 90.130 222.150 94.080 222.300 ;
        RECT 95.380 222.150 99.330 222.300 ;
        RECT 90.130 222.000 90.730 222.150 ;
        RECT 86.530 221.700 90.730 222.000 ;
        RECT 98.730 222.000 99.330 222.150 ;
        RECT 99.780 222.000 99.930 229.550 ;
        RECT 100.380 222.000 100.530 229.550 ;
        RECT 100.980 222.000 101.130 229.550 ;
        RECT 101.580 222.000 101.730 229.550 ;
        RECT 102.180 222.000 102.330 229.550 ;
        RECT 102.780 222.000 102.930 224.900 ;
        RECT 98.730 221.700 102.930 222.000 ;
        RECT 86.530 221.550 94.080 221.700 ;
        RECT 95.380 221.550 102.930 221.700 ;
        RECT 86.530 221.350 90.730 221.550 ;
        RECT 80.330 221.050 89.130 221.200 ;
        RECT 89.280 221.050 90.730 221.350 ;
        RECT 78.730 220.150 90.730 221.050 ;
        RECT 98.730 221.350 102.930 221.550 ;
        RECT 103.530 222.185 104.730 224.400 ;
        RECT 98.730 221.050 100.180 221.350 ;
        RECT 103.530 221.200 107.140 222.185 ;
        RECT 100.330 221.050 107.140 221.200 ;
        RECT 98.730 220.910 107.140 221.050 ;
        RECT 98.730 220.150 104.730 220.910 ;
        RECT 4.730 220.000 9.130 220.150 ;
        RECT 20.330 220.000 29.130 220.150 ;
        RECT 40.330 220.000 49.130 220.150 ;
        RECT 60.330 220.000 69.130 220.150 ;
        RECT 80.330 220.000 89.130 220.150 ;
        RECT 100.330 220.000 104.730 220.150 ;
        RECT 4.620 195.695 5.940 195.865 ;
        RECT 6.940 195.695 7.400 195.700 ;
        RECT 2.315 195.215 23.605 195.695 ;
        RECT 4.620 194.615 5.940 195.215 ;
        RECT 7.960 194.410 9.830 194.770 ;
        RECT 2.315 189.775 24.065 190.255 ;
        RECT 4.620 184.815 5.940 185.555 ;
        RECT 2.315 184.335 23.605 184.815 ;
        RECT 4.620 184.175 5.940 184.335 ;
        RECT 42.635 182.510 47.035 182.660 ;
        RECT 58.235 182.510 67.035 182.660 ;
        RECT 78.235 182.510 87.035 182.660 ;
        RECT 42.635 181.610 48.635 182.510 ;
        RECT 58.235 182.460 68.635 182.510 ;
        RECT 78.235 182.460 88.635 182.510 ;
        RECT 98.235 182.460 102.635 182.660 ;
        RECT 42.635 181.460 47.035 181.610 ;
        RECT 42.635 178.260 43.835 181.460 ;
        RECT 47.185 181.310 48.635 181.610 ;
        RECT 44.435 181.110 48.635 181.310 ;
        RECT 56.635 181.610 68.635 182.460 ;
        RECT 56.635 181.560 67.035 181.610 ;
        RECT 56.635 181.310 58.085 181.560 ;
        RECT 58.235 181.460 67.035 181.560 ;
        RECT 56.635 181.110 60.835 181.310 ;
        RECT 44.435 180.960 51.985 181.110 ;
        RECT 53.335 180.960 60.835 181.110 ;
        RECT 44.435 180.660 48.635 180.960 ;
        RECT 44.435 177.810 44.585 180.660 ;
        RECT 45.035 173.110 45.185 180.660 ;
        RECT 45.635 173.110 45.785 180.660 ;
        RECT 46.235 173.110 46.385 180.660 ;
        RECT 46.835 173.110 46.985 180.660 ;
        RECT 47.435 173.110 47.585 180.660 ;
        RECT 48.035 180.510 48.635 180.660 ;
        RECT 56.635 180.660 60.835 180.960 ;
        RECT 56.635 180.510 57.235 180.660 ;
        RECT 48.035 180.360 51.985 180.510 ;
        RECT 53.285 180.360 57.235 180.510 ;
        RECT 48.035 179.910 48.635 180.360 ;
        RECT 56.635 179.910 57.235 180.360 ;
        RECT 48.035 179.760 51.985 179.910 ;
        RECT 53.285 179.760 57.235 179.910 ;
        RECT 48.035 179.310 48.635 179.760 ;
        RECT 56.635 179.310 57.235 179.760 ;
        RECT 48.035 179.160 51.985 179.310 ;
        RECT 53.285 179.160 57.235 179.310 ;
        RECT 48.035 178.710 48.635 179.160 ;
        RECT 56.635 178.710 57.235 179.160 ;
        RECT 48.035 178.560 51.985 178.710 ;
        RECT 53.285 178.560 57.235 178.710 ;
        RECT 48.035 178.110 48.635 178.560 ;
        RECT 56.635 178.110 57.235 178.560 ;
        RECT 48.035 177.960 51.985 178.110 ;
        RECT 53.285 177.960 57.235 178.110 ;
        RECT 48.035 177.510 48.635 177.960 ;
        RECT 56.635 177.510 57.235 177.960 ;
        RECT 48.035 177.360 51.985 177.510 ;
        RECT 53.285 177.360 57.235 177.510 ;
        RECT 48.035 176.910 48.635 177.360 ;
        RECT 56.635 176.910 57.235 177.360 ;
        RECT 48.035 176.760 51.985 176.910 ;
        RECT 53.285 176.760 57.235 176.910 ;
        RECT 48.035 176.310 48.635 176.760 ;
        RECT 56.635 176.310 57.235 176.760 ;
        RECT 48.035 176.160 51.985 176.310 ;
        RECT 53.285 176.160 57.235 176.310 ;
        RECT 48.035 175.710 48.635 176.160 ;
        RECT 56.635 175.710 57.235 176.160 ;
        RECT 48.035 175.560 51.985 175.710 ;
        RECT 53.285 175.560 57.235 175.710 ;
        RECT 48.035 175.110 48.635 175.560 ;
        RECT 56.635 175.110 57.235 175.560 ;
        RECT 48.035 174.960 51.985 175.110 ;
        RECT 53.285 174.960 57.235 175.110 ;
        RECT 48.035 174.510 48.635 174.960 ;
        RECT 56.635 174.510 57.235 174.960 ;
        RECT 48.035 174.360 51.985 174.510 ;
        RECT 53.285 174.360 57.235 174.510 ;
        RECT 48.035 173.910 48.635 174.360 ;
        RECT 56.635 173.910 57.235 174.360 ;
        RECT 48.035 173.760 51.985 173.910 ;
        RECT 53.285 173.760 57.235 173.910 ;
        RECT 48.035 173.310 48.635 173.760 ;
        RECT 56.635 173.310 57.235 173.760 ;
        RECT 48.035 173.110 51.985 173.310 ;
        RECT 53.285 173.110 57.235 173.310 ;
        RECT 57.685 173.110 57.835 180.660 ;
        RECT 58.285 173.110 58.435 180.660 ;
        RECT 58.885 173.110 59.035 180.660 ;
        RECT 59.485 173.110 59.635 180.660 ;
        RECT 60.085 173.110 60.235 180.660 ;
        RECT 60.685 177.810 60.835 180.660 ;
        RECT 61.435 178.260 63.835 181.460 ;
        RECT 67.185 181.310 68.635 181.610 ;
        RECT 64.435 181.110 68.635 181.310 ;
        RECT 76.635 181.610 88.635 182.460 ;
        RECT 76.635 181.560 87.035 181.610 ;
        RECT 76.635 181.310 78.085 181.560 ;
        RECT 78.235 181.460 87.035 181.560 ;
        RECT 76.635 181.110 80.835 181.310 ;
        RECT 64.435 180.960 71.985 181.110 ;
        RECT 73.335 180.960 80.835 181.110 ;
        RECT 64.435 180.660 68.635 180.960 ;
        RECT 64.435 177.810 64.585 180.660 ;
        RECT 65.035 173.110 65.185 180.660 ;
        RECT 65.635 173.110 65.785 180.660 ;
        RECT 66.235 173.110 66.385 180.660 ;
        RECT 66.835 173.110 66.985 180.660 ;
        RECT 67.435 173.110 67.585 180.660 ;
        RECT 68.035 180.510 68.635 180.660 ;
        RECT 76.635 180.660 80.835 180.960 ;
        RECT 76.635 180.510 77.235 180.660 ;
        RECT 68.035 180.360 71.985 180.510 ;
        RECT 73.285 180.360 77.235 180.510 ;
        RECT 68.035 179.910 68.635 180.360 ;
        RECT 76.635 179.910 77.235 180.360 ;
        RECT 68.035 179.760 71.985 179.910 ;
        RECT 73.285 179.760 77.235 179.910 ;
        RECT 68.035 179.310 68.635 179.760 ;
        RECT 76.635 179.310 77.235 179.760 ;
        RECT 68.035 179.160 71.985 179.310 ;
        RECT 73.285 179.160 77.235 179.310 ;
        RECT 68.035 178.710 68.635 179.160 ;
        RECT 76.635 178.710 77.235 179.160 ;
        RECT 68.035 178.560 71.985 178.710 ;
        RECT 73.285 178.560 77.235 178.710 ;
        RECT 68.035 178.110 68.635 178.560 ;
        RECT 76.635 178.110 77.235 178.560 ;
        RECT 68.035 177.960 71.985 178.110 ;
        RECT 73.285 177.960 77.235 178.110 ;
        RECT 68.035 177.510 68.635 177.960 ;
        RECT 76.635 177.510 77.235 177.960 ;
        RECT 68.035 177.360 71.985 177.510 ;
        RECT 73.285 177.360 77.235 177.510 ;
        RECT 68.035 176.910 68.635 177.360 ;
        RECT 76.635 176.910 77.235 177.360 ;
        RECT 68.035 176.760 71.985 176.910 ;
        RECT 73.285 176.760 77.235 176.910 ;
        RECT 68.035 176.310 68.635 176.760 ;
        RECT 76.635 176.310 77.235 176.760 ;
        RECT 68.035 176.160 71.985 176.310 ;
        RECT 73.285 176.160 77.235 176.310 ;
        RECT 68.035 175.710 68.635 176.160 ;
        RECT 76.635 175.710 77.235 176.160 ;
        RECT 68.035 175.560 71.985 175.710 ;
        RECT 73.285 175.560 77.235 175.710 ;
        RECT 68.035 175.110 68.635 175.560 ;
        RECT 76.635 175.110 77.235 175.560 ;
        RECT 68.035 174.960 71.985 175.110 ;
        RECT 73.285 174.960 77.235 175.110 ;
        RECT 68.035 174.510 68.635 174.960 ;
        RECT 76.635 174.510 77.235 174.960 ;
        RECT 68.035 174.360 71.985 174.510 ;
        RECT 73.285 174.360 77.235 174.510 ;
        RECT 68.035 173.910 68.635 174.360 ;
        RECT 76.635 173.910 77.235 174.360 ;
        RECT 68.035 173.760 71.985 173.910 ;
        RECT 73.285 173.760 77.235 173.910 ;
        RECT 68.035 173.310 68.635 173.760 ;
        RECT 76.635 173.310 77.235 173.760 ;
        RECT 68.035 173.110 71.985 173.310 ;
        RECT 73.285 173.110 77.235 173.310 ;
        RECT 77.685 173.110 77.835 180.660 ;
        RECT 78.285 173.110 78.435 180.660 ;
        RECT 78.885 173.110 79.035 180.660 ;
        RECT 79.485 173.110 79.635 180.660 ;
        RECT 80.085 173.110 80.235 180.660 ;
        RECT 80.685 177.810 80.835 180.660 ;
        RECT 81.435 178.260 83.835 181.460 ;
        RECT 87.185 181.310 88.635 181.610 ;
        RECT 84.435 181.110 88.635 181.310 ;
        RECT 96.635 181.560 102.635 182.460 ;
        RECT 96.635 181.310 98.085 181.560 ;
        RECT 98.235 181.460 102.635 181.560 ;
        RECT 96.635 181.110 100.835 181.310 ;
        RECT 84.435 180.960 91.985 181.110 ;
        RECT 93.335 180.960 100.835 181.110 ;
        RECT 84.435 180.660 88.635 180.960 ;
        RECT 84.435 177.810 84.585 180.660 ;
        RECT 85.035 173.110 85.185 180.660 ;
        RECT 85.635 173.110 85.785 180.660 ;
        RECT 86.235 173.110 86.385 180.660 ;
        RECT 86.835 173.110 86.985 180.660 ;
        RECT 87.435 173.110 87.585 180.660 ;
        RECT 88.035 180.510 88.635 180.660 ;
        RECT 96.635 180.660 100.835 180.960 ;
        RECT 96.635 180.510 97.235 180.660 ;
        RECT 88.035 180.360 91.985 180.510 ;
        RECT 93.285 180.360 97.235 180.510 ;
        RECT 88.035 179.910 88.635 180.360 ;
        RECT 96.635 179.910 97.235 180.360 ;
        RECT 88.035 179.760 91.985 179.910 ;
        RECT 93.285 179.760 97.235 179.910 ;
        RECT 88.035 179.310 88.635 179.760 ;
        RECT 96.635 179.310 97.235 179.760 ;
        RECT 88.035 179.160 91.985 179.310 ;
        RECT 93.285 179.160 97.235 179.310 ;
        RECT 88.035 178.710 88.635 179.160 ;
        RECT 96.635 178.710 97.235 179.160 ;
        RECT 88.035 178.560 91.985 178.710 ;
        RECT 93.285 178.560 97.235 178.710 ;
        RECT 88.035 178.110 88.635 178.560 ;
        RECT 96.635 178.110 97.235 178.560 ;
        RECT 88.035 177.960 91.985 178.110 ;
        RECT 93.285 177.960 97.235 178.110 ;
        RECT 88.035 177.510 88.635 177.960 ;
        RECT 96.635 177.510 97.235 177.960 ;
        RECT 88.035 177.360 91.985 177.510 ;
        RECT 93.285 177.360 97.235 177.510 ;
        RECT 88.035 176.910 88.635 177.360 ;
        RECT 96.635 176.910 97.235 177.360 ;
        RECT 88.035 176.760 91.985 176.910 ;
        RECT 93.285 176.760 97.235 176.910 ;
        RECT 88.035 176.310 88.635 176.760 ;
        RECT 96.635 176.310 97.235 176.760 ;
        RECT 88.035 176.160 91.985 176.310 ;
        RECT 93.285 176.160 97.235 176.310 ;
        RECT 88.035 175.710 88.635 176.160 ;
        RECT 96.635 175.710 97.235 176.160 ;
        RECT 88.035 175.560 91.985 175.710 ;
        RECT 93.285 175.560 97.235 175.710 ;
        RECT 88.035 175.110 88.635 175.560 ;
        RECT 96.635 175.110 97.235 175.560 ;
        RECT 88.035 174.960 91.985 175.110 ;
        RECT 93.285 174.960 97.235 175.110 ;
        RECT 88.035 174.510 88.635 174.960 ;
        RECT 96.635 174.510 97.235 174.960 ;
        RECT 88.035 174.360 91.985 174.510 ;
        RECT 93.285 174.360 97.235 174.510 ;
        RECT 88.035 173.910 88.635 174.360 ;
        RECT 96.635 173.910 97.235 174.360 ;
        RECT 88.035 173.760 91.985 173.910 ;
        RECT 93.285 173.760 97.235 173.910 ;
        RECT 88.035 173.310 88.635 173.760 ;
        RECT 96.635 173.310 97.235 173.760 ;
        RECT 88.035 173.110 91.985 173.310 ;
        RECT 93.285 173.110 97.235 173.310 ;
        RECT 97.685 173.110 97.835 180.660 ;
        RECT 98.285 173.110 98.435 180.660 ;
        RECT 98.885 173.110 99.035 180.660 ;
        RECT 99.485 173.110 99.635 180.660 ;
        RECT 100.085 173.110 100.235 180.660 ;
        RECT 100.685 177.810 100.835 180.660 ;
        RECT 101.435 180.990 102.635 181.460 ;
        RECT 101.435 179.715 107.140 180.990 ;
        RECT 101.435 178.260 102.635 179.715 ;
        RECT 105.140 175.915 107.140 178.210 ;
        RECT 105.140 175.910 107.005 175.915 ;
        RECT 42.635 163.860 43.835 167.060 ;
        RECT 44.435 164.660 44.585 167.560 ;
        RECT 45.035 164.660 45.185 172.210 ;
        RECT 45.635 164.660 45.785 172.210 ;
        RECT 46.235 164.660 46.385 172.210 ;
        RECT 46.835 164.660 46.985 172.210 ;
        RECT 47.435 164.660 47.585 172.210 ;
        RECT 48.035 172.010 51.985 172.210 ;
        RECT 53.285 172.010 57.235 172.210 ;
        RECT 48.035 171.560 48.635 172.010 ;
        RECT 56.635 171.560 57.235 172.010 ;
        RECT 48.035 171.410 51.985 171.560 ;
        RECT 53.285 171.410 57.235 171.560 ;
        RECT 48.035 170.960 48.635 171.410 ;
        RECT 56.635 170.960 57.235 171.410 ;
        RECT 48.035 170.810 51.985 170.960 ;
        RECT 53.285 170.810 57.235 170.960 ;
        RECT 48.035 170.360 48.635 170.810 ;
        RECT 56.635 170.360 57.235 170.810 ;
        RECT 48.035 170.210 51.985 170.360 ;
        RECT 53.285 170.210 57.235 170.360 ;
        RECT 48.035 169.760 48.635 170.210 ;
        RECT 56.635 169.760 57.235 170.210 ;
        RECT 48.035 169.610 51.985 169.760 ;
        RECT 53.285 169.610 57.235 169.760 ;
        RECT 48.035 169.160 48.635 169.610 ;
        RECT 56.635 169.160 57.235 169.610 ;
        RECT 48.035 169.010 51.985 169.160 ;
        RECT 53.285 169.010 57.235 169.160 ;
        RECT 48.035 168.560 48.635 169.010 ;
        RECT 56.635 168.560 57.235 169.010 ;
        RECT 48.035 168.410 51.985 168.560 ;
        RECT 53.285 168.410 57.235 168.560 ;
        RECT 48.035 167.960 48.635 168.410 ;
        RECT 56.635 167.960 57.235 168.410 ;
        RECT 48.035 167.810 51.985 167.960 ;
        RECT 53.285 167.810 57.235 167.960 ;
        RECT 48.035 167.360 48.635 167.810 ;
        RECT 56.635 167.360 57.235 167.810 ;
        RECT 48.035 167.210 51.985 167.360 ;
        RECT 53.285 167.210 57.235 167.360 ;
        RECT 48.035 166.760 48.635 167.210 ;
        RECT 56.635 166.760 57.235 167.210 ;
        RECT 48.035 166.610 51.985 166.760 ;
        RECT 53.285 166.610 57.235 166.760 ;
        RECT 48.035 166.160 48.635 166.610 ;
        RECT 56.635 166.160 57.235 166.610 ;
        RECT 48.035 166.010 51.985 166.160 ;
        RECT 53.285 166.010 57.235 166.160 ;
        RECT 48.035 165.560 48.635 166.010 ;
        RECT 56.635 165.560 57.235 166.010 ;
        RECT 48.035 165.410 51.985 165.560 ;
        RECT 53.285 165.410 57.235 165.560 ;
        RECT 48.035 164.960 48.635 165.410 ;
        RECT 56.635 164.960 57.235 165.410 ;
        RECT 48.035 164.810 51.985 164.960 ;
        RECT 53.285 164.810 57.235 164.960 ;
        RECT 48.035 164.660 48.635 164.810 ;
        RECT 44.435 164.360 48.635 164.660 ;
        RECT 56.635 164.660 57.235 164.810 ;
        RECT 57.685 164.660 57.835 172.210 ;
        RECT 58.285 164.660 58.435 172.210 ;
        RECT 58.885 164.660 59.035 172.210 ;
        RECT 59.485 164.660 59.635 172.210 ;
        RECT 60.085 164.660 60.235 172.210 ;
        RECT 60.685 164.660 60.835 167.560 ;
        RECT 56.635 164.360 60.835 164.660 ;
        RECT 44.435 164.210 51.985 164.360 ;
        RECT 53.285 164.210 60.835 164.360 ;
        RECT 44.435 164.010 48.635 164.210 ;
        RECT 42.635 163.710 47.035 163.860 ;
        RECT 47.185 163.710 48.635 164.010 ;
        RECT 42.635 162.810 48.635 163.710 ;
        RECT 56.635 164.010 60.835 164.210 ;
        RECT 56.635 163.710 58.085 164.010 ;
        RECT 61.435 163.860 63.835 167.060 ;
        RECT 64.435 164.660 64.585 167.560 ;
        RECT 65.035 164.660 65.185 172.210 ;
        RECT 65.635 164.660 65.785 172.210 ;
        RECT 66.235 164.660 66.385 172.210 ;
        RECT 66.835 164.660 66.985 172.210 ;
        RECT 67.435 164.660 67.585 172.210 ;
        RECT 68.035 172.010 71.985 172.210 ;
        RECT 73.285 172.010 77.235 172.210 ;
        RECT 68.035 171.560 68.635 172.010 ;
        RECT 76.635 171.560 77.235 172.010 ;
        RECT 68.035 171.410 71.985 171.560 ;
        RECT 73.285 171.410 77.235 171.560 ;
        RECT 68.035 170.960 68.635 171.410 ;
        RECT 76.635 170.960 77.235 171.410 ;
        RECT 68.035 170.810 71.985 170.960 ;
        RECT 73.285 170.810 77.235 170.960 ;
        RECT 68.035 170.360 68.635 170.810 ;
        RECT 76.635 170.360 77.235 170.810 ;
        RECT 68.035 170.210 71.985 170.360 ;
        RECT 73.285 170.210 77.235 170.360 ;
        RECT 68.035 169.760 68.635 170.210 ;
        RECT 76.635 169.760 77.235 170.210 ;
        RECT 68.035 169.610 71.985 169.760 ;
        RECT 73.285 169.610 77.235 169.760 ;
        RECT 68.035 169.160 68.635 169.610 ;
        RECT 76.635 169.160 77.235 169.610 ;
        RECT 68.035 169.010 71.985 169.160 ;
        RECT 73.285 169.010 77.235 169.160 ;
        RECT 68.035 168.560 68.635 169.010 ;
        RECT 76.635 168.560 77.235 169.010 ;
        RECT 68.035 168.410 71.985 168.560 ;
        RECT 73.285 168.410 77.235 168.560 ;
        RECT 68.035 167.960 68.635 168.410 ;
        RECT 76.635 167.960 77.235 168.410 ;
        RECT 68.035 167.810 71.985 167.960 ;
        RECT 73.285 167.810 77.235 167.960 ;
        RECT 68.035 167.360 68.635 167.810 ;
        RECT 76.635 167.360 77.235 167.810 ;
        RECT 68.035 167.210 71.985 167.360 ;
        RECT 73.285 167.210 77.235 167.360 ;
        RECT 68.035 166.760 68.635 167.210 ;
        RECT 76.635 166.760 77.235 167.210 ;
        RECT 68.035 166.610 71.985 166.760 ;
        RECT 73.285 166.610 77.235 166.760 ;
        RECT 68.035 166.160 68.635 166.610 ;
        RECT 76.635 166.160 77.235 166.610 ;
        RECT 68.035 166.010 71.985 166.160 ;
        RECT 73.285 166.010 77.235 166.160 ;
        RECT 68.035 165.560 68.635 166.010 ;
        RECT 76.635 165.560 77.235 166.010 ;
        RECT 68.035 165.410 71.985 165.560 ;
        RECT 73.285 165.410 77.235 165.560 ;
        RECT 68.035 164.960 68.635 165.410 ;
        RECT 76.635 164.960 77.235 165.410 ;
        RECT 68.035 164.810 71.985 164.960 ;
        RECT 73.285 164.810 77.235 164.960 ;
        RECT 68.035 164.660 68.635 164.810 ;
        RECT 64.435 164.360 68.635 164.660 ;
        RECT 76.635 164.660 77.235 164.810 ;
        RECT 77.685 164.660 77.835 172.210 ;
        RECT 78.285 164.660 78.435 172.210 ;
        RECT 78.885 164.660 79.035 172.210 ;
        RECT 79.485 164.660 79.635 172.210 ;
        RECT 80.085 164.660 80.235 172.210 ;
        RECT 80.685 164.660 80.835 167.560 ;
        RECT 76.635 164.360 80.835 164.660 ;
        RECT 64.435 164.210 71.985 164.360 ;
        RECT 73.285 164.210 80.835 164.360 ;
        RECT 64.435 164.010 68.635 164.210 ;
        RECT 58.235 163.710 67.035 163.860 ;
        RECT 67.185 163.710 68.635 164.010 ;
        RECT 56.635 162.810 68.635 163.710 ;
        RECT 76.635 164.010 80.835 164.210 ;
        RECT 76.635 163.710 78.085 164.010 ;
        RECT 81.435 163.860 83.835 167.060 ;
        RECT 84.435 164.660 84.585 167.560 ;
        RECT 85.035 164.660 85.185 172.210 ;
        RECT 85.635 164.660 85.785 172.210 ;
        RECT 86.235 164.660 86.385 172.210 ;
        RECT 86.835 164.660 86.985 172.210 ;
        RECT 87.435 164.660 87.585 172.210 ;
        RECT 88.035 172.010 91.985 172.210 ;
        RECT 93.285 172.010 97.235 172.210 ;
        RECT 88.035 171.560 88.635 172.010 ;
        RECT 96.635 171.560 97.235 172.010 ;
        RECT 88.035 171.410 91.985 171.560 ;
        RECT 93.285 171.410 97.235 171.560 ;
        RECT 88.035 170.960 88.635 171.410 ;
        RECT 96.635 170.960 97.235 171.410 ;
        RECT 88.035 170.810 91.985 170.960 ;
        RECT 93.285 170.810 97.235 170.960 ;
        RECT 88.035 170.360 88.635 170.810 ;
        RECT 96.635 170.360 97.235 170.810 ;
        RECT 88.035 170.210 91.985 170.360 ;
        RECT 93.285 170.210 97.235 170.360 ;
        RECT 88.035 169.760 88.635 170.210 ;
        RECT 96.635 169.760 97.235 170.210 ;
        RECT 88.035 169.610 91.985 169.760 ;
        RECT 93.285 169.610 97.235 169.760 ;
        RECT 88.035 169.160 88.635 169.610 ;
        RECT 96.635 169.160 97.235 169.610 ;
        RECT 88.035 169.010 91.985 169.160 ;
        RECT 93.285 169.010 97.235 169.160 ;
        RECT 88.035 168.560 88.635 169.010 ;
        RECT 96.635 168.560 97.235 169.010 ;
        RECT 88.035 168.410 91.985 168.560 ;
        RECT 93.285 168.410 97.235 168.560 ;
        RECT 88.035 167.960 88.635 168.410 ;
        RECT 96.635 167.960 97.235 168.410 ;
        RECT 88.035 167.810 91.985 167.960 ;
        RECT 93.285 167.810 97.235 167.960 ;
        RECT 88.035 167.360 88.635 167.810 ;
        RECT 96.635 167.360 97.235 167.810 ;
        RECT 88.035 167.210 91.985 167.360 ;
        RECT 93.285 167.210 97.235 167.360 ;
        RECT 88.035 166.760 88.635 167.210 ;
        RECT 96.635 166.760 97.235 167.210 ;
        RECT 88.035 166.610 91.985 166.760 ;
        RECT 93.285 166.610 97.235 166.760 ;
        RECT 88.035 166.160 88.635 166.610 ;
        RECT 96.635 166.160 97.235 166.610 ;
        RECT 88.035 166.010 91.985 166.160 ;
        RECT 93.285 166.010 97.235 166.160 ;
        RECT 88.035 165.560 88.635 166.010 ;
        RECT 96.635 165.560 97.235 166.010 ;
        RECT 88.035 165.410 91.985 165.560 ;
        RECT 93.285 165.410 97.235 165.560 ;
        RECT 88.035 164.960 88.635 165.410 ;
        RECT 96.635 164.960 97.235 165.410 ;
        RECT 88.035 164.810 91.985 164.960 ;
        RECT 93.285 164.810 97.235 164.960 ;
        RECT 88.035 164.660 88.635 164.810 ;
        RECT 84.435 164.360 88.635 164.660 ;
        RECT 96.635 164.660 97.235 164.810 ;
        RECT 97.685 164.660 97.835 172.210 ;
        RECT 98.285 164.660 98.435 172.210 ;
        RECT 98.885 164.660 99.035 172.210 ;
        RECT 99.485 164.660 99.635 172.210 ;
        RECT 100.085 164.660 100.235 172.210 ;
        RECT 100.685 164.660 100.835 167.560 ;
        RECT 105.140 167.115 107.140 169.410 ;
        RECT 105.140 167.110 107.005 167.115 ;
        RECT 96.635 164.360 100.835 164.660 ;
        RECT 84.435 164.210 91.985 164.360 ;
        RECT 93.285 164.210 100.835 164.360 ;
        RECT 84.435 164.010 88.635 164.210 ;
        RECT 78.235 163.710 87.035 163.860 ;
        RECT 87.185 163.710 88.635 164.010 ;
        RECT 76.635 162.810 88.635 163.710 ;
        RECT 96.635 164.010 100.835 164.210 ;
        RECT 101.435 165.715 102.635 167.060 ;
        RECT 101.435 164.440 107.135 165.715 ;
        RECT 96.635 163.710 98.085 164.010 ;
        RECT 101.435 163.860 102.635 164.440 ;
        RECT 98.235 163.710 102.635 163.860 ;
        RECT 96.635 162.810 102.635 163.710 ;
        RECT 42.635 162.660 47.035 162.810 ;
        RECT 58.235 162.660 67.035 162.810 ;
        RECT 78.235 162.660 87.035 162.810 ;
        RECT 98.235 162.660 102.635 162.810 ;
        RECT 2.315 160.365 107.140 161.800 ;
        RECT 2.315 160.360 9.125 160.365 ;
        RECT 11.565 160.360 107.140 160.365 ;
        RECT 4.730 159.850 9.130 160.000 ;
        RECT 20.330 159.850 29.130 160.000 ;
        RECT 40.330 159.850 49.130 160.000 ;
        RECT 60.330 159.850 69.130 160.000 ;
        RECT 80.330 159.850 89.130 160.000 ;
        RECT 4.730 158.950 10.730 159.850 ;
        RECT 20.330 159.800 30.730 159.850 ;
        RECT 40.330 159.800 50.730 159.850 ;
        RECT 60.330 159.800 70.730 159.850 ;
        RECT 80.330 159.800 90.730 159.850 ;
        RECT 100.330 159.800 104.730 160.000 ;
        RECT 4.730 158.800 9.130 158.950 ;
        RECT 4.730 157.725 5.930 158.800 ;
        RECT 9.280 158.650 10.730 158.950 ;
        RECT 2.315 156.450 5.930 157.725 ;
        RECT 4.730 155.600 5.930 156.450 ;
        RECT 6.530 158.450 10.730 158.650 ;
        RECT 18.730 158.950 30.730 159.800 ;
        RECT 18.730 158.900 29.130 158.950 ;
        RECT 18.730 158.650 20.180 158.900 ;
        RECT 20.330 158.800 29.130 158.900 ;
        RECT 18.730 158.450 22.930 158.650 ;
        RECT 6.530 158.300 14.080 158.450 ;
        RECT 15.430 158.300 22.930 158.450 ;
        RECT 6.530 158.000 10.730 158.300 ;
        RECT 2.315 153.255 4.315 155.555 ;
        RECT 6.530 155.150 6.680 158.000 ;
        RECT 7.130 150.450 7.280 158.000 ;
        RECT 7.730 150.450 7.880 158.000 ;
        RECT 8.330 150.450 8.480 158.000 ;
        RECT 8.930 150.450 9.080 158.000 ;
        RECT 9.530 150.450 9.680 158.000 ;
        RECT 10.130 157.850 10.730 158.000 ;
        RECT 18.730 158.000 22.930 158.300 ;
        RECT 18.730 157.850 19.330 158.000 ;
        RECT 10.130 157.700 14.080 157.850 ;
        RECT 15.380 157.700 19.330 157.850 ;
        RECT 10.130 157.250 10.730 157.700 ;
        RECT 18.730 157.250 19.330 157.700 ;
        RECT 10.130 157.100 14.080 157.250 ;
        RECT 15.380 157.100 19.330 157.250 ;
        RECT 10.130 156.650 10.730 157.100 ;
        RECT 18.730 156.650 19.330 157.100 ;
        RECT 10.130 156.500 14.080 156.650 ;
        RECT 15.380 156.500 19.330 156.650 ;
        RECT 10.130 156.050 10.730 156.500 ;
        RECT 18.730 156.050 19.330 156.500 ;
        RECT 10.130 155.900 14.080 156.050 ;
        RECT 15.380 155.900 19.330 156.050 ;
        RECT 10.130 155.450 10.730 155.900 ;
        RECT 18.730 155.450 19.330 155.900 ;
        RECT 10.130 155.300 14.080 155.450 ;
        RECT 15.380 155.300 19.330 155.450 ;
        RECT 10.130 154.850 10.730 155.300 ;
        RECT 18.730 154.850 19.330 155.300 ;
        RECT 10.130 154.700 14.080 154.850 ;
        RECT 15.380 154.700 19.330 154.850 ;
        RECT 10.130 154.250 10.730 154.700 ;
        RECT 18.730 154.250 19.330 154.700 ;
        RECT 10.130 154.100 14.080 154.250 ;
        RECT 15.380 154.100 19.330 154.250 ;
        RECT 10.130 153.650 10.730 154.100 ;
        RECT 18.730 153.650 19.330 154.100 ;
        RECT 10.130 153.500 14.080 153.650 ;
        RECT 15.380 153.500 19.330 153.650 ;
        RECT 10.130 153.050 10.730 153.500 ;
        RECT 18.730 153.050 19.330 153.500 ;
        RECT 10.130 152.900 14.080 153.050 ;
        RECT 15.380 152.900 19.330 153.050 ;
        RECT 10.130 152.450 10.730 152.900 ;
        RECT 18.730 152.450 19.330 152.900 ;
        RECT 10.130 152.300 14.080 152.450 ;
        RECT 15.380 152.300 19.330 152.450 ;
        RECT 10.130 151.850 10.730 152.300 ;
        RECT 18.730 151.850 19.330 152.300 ;
        RECT 10.130 151.700 14.080 151.850 ;
        RECT 15.380 151.700 19.330 151.850 ;
        RECT 10.130 151.250 10.730 151.700 ;
        RECT 18.730 151.250 19.330 151.700 ;
        RECT 10.130 151.100 14.080 151.250 ;
        RECT 15.380 151.100 19.330 151.250 ;
        RECT 10.130 150.650 10.730 151.100 ;
        RECT 18.730 150.650 19.330 151.100 ;
        RECT 10.130 150.450 14.080 150.650 ;
        RECT 15.380 150.450 19.330 150.650 ;
        RECT 19.780 150.450 19.930 158.000 ;
        RECT 20.380 150.450 20.530 158.000 ;
        RECT 20.980 150.450 21.130 158.000 ;
        RECT 21.580 150.450 21.730 158.000 ;
        RECT 22.180 150.450 22.330 158.000 ;
        RECT 22.780 155.150 22.930 158.000 ;
        RECT 23.530 155.600 25.930 158.800 ;
        RECT 29.280 158.650 30.730 158.950 ;
        RECT 26.530 158.450 30.730 158.650 ;
        RECT 38.730 158.950 50.730 159.800 ;
        RECT 38.730 158.900 49.130 158.950 ;
        RECT 38.730 158.650 40.180 158.900 ;
        RECT 40.330 158.800 49.130 158.900 ;
        RECT 38.730 158.450 42.930 158.650 ;
        RECT 26.530 158.300 34.080 158.450 ;
        RECT 35.430 158.300 42.930 158.450 ;
        RECT 26.530 158.000 30.730 158.300 ;
        RECT 26.530 155.150 26.680 158.000 ;
        RECT 27.130 150.450 27.280 158.000 ;
        RECT 27.730 150.450 27.880 158.000 ;
        RECT 28.330 150.450 28.480 158.000 ;
        RECT 28.930 150.450 29.080 158.000 ;
        RECT 29.530 150.450 29.680 158.000 ;
        RECT 30.130 157.850 30.730 158.000 ;
        RECT 38.730 158.000 42.930 158.300 ;
        RECT 38.730 157.850 39.330 158.000 ;
        RECT 30.130 157.700 34.080 157.850 ;
        RECT 35.380 157.700 39.330 157.850 ;
        RECT 30.130 157.250 30.730 157.700 ;
        RECT 38.730 157.250 39.330 157.700 ;
        RECT 30.130 157.100 34.080 157.250 ;
        RECT 35.380 157.100 39.330 157.250 ;
        RECT 30.130 156.650 30.730 157.100 ;
        RECT 38.730 156.650 39.330 157.100 ;
        RECT 30.130 156.500 34.080 156.650 ;
        RECT 35.380 156.500 39.330 156.650 ;
        RECT 30.130 156.050 30.730 156.500 ;
        RECT 38.730 156.050 39.330 156.500 ;
        RECT 30.130 155.900 34.080 156.050 ;
        RECT 35.380 155.900 39.330 156.050 ;
        RECT 30.130 155.450 30.730 155.900 ;
        RECT 38.730 155.450 39.330 155.900 ;
        RECT 30.130 155.300 34.080 155.450 ;
        RECT 35.380 155.300 39.330 155.450 ;
        RECT 30.130 154.850 30.730 155.300 ;
        RECT 38.730 154.850 39.330 155.300 ;
        RECT 30.130 154.700 34.080 154.850 ;
        RECT 35.380 154.700 39.330 154.850 ;
        RECT 30.130 154.250 30.730 154.700 ;
        RECT 38.730 154.250 39.330 154.700 ;
        RECT 30.130 154.100 34.080 154.250 ;
        RECT 35.380 154.100 39.330 154.250 ;
        RECT 30.130 153.650 30.730 154.100 ;
        RECT 38.730 153.650 39.330 154.100 ;
        RECT 30.130 153.500 34.080 153.650 ;
        RECT 35.380 153.500 39.330 153.650 ;
        RECT 30.130 153.050 30.730 153.500 ;
        RECT 38.730 153.050 39.330 153.500 ;
        RECT 30.130 152.900 34.080 153.050 ;
        RECT 35.380 152.900 39.330 153.050 ;
        RECT 30.130 152.450 30.730 152.900 ;
        RECT 38.730 152.450 39.330 152.900 ;
        RECT 30.130 152.300 34.080 152.450 ;
        RECT 35.380 152.300 39.330 152.450 ;
        RECT 30.130 151.850 30.730 152.300 ;
        RECT 38.730 151.850 39.330 152.300 ;
        RECT 30.130 151.700 34.080 151.850 ;
        RECT 35.380 151.700 39.330 151.850 ;
        RECT 30.130 151.250 30.730 151.700 ;
        RECT 38.730 151.250 39.330 151.700 ;
        RECT 30.130 151.100 34.080 151.250 ;
        RECT 35.380 151.100 39.330 151.250 ;
        RECT 30.130 150.650 30.730 151.100 ;
        RECT 38.730 150.650 39.330 151.100 ;
        RECT 30.130 150.450 34.080 150.650 ;
        RECT 35.380 150.450 39.330 150.650 ;
        RECT 39.780 150.450 39.930 158.000 ;
        RECT 40.380 150.450 40.530 158.000 ;
        RECT 40.980 150.450 41.130 158.000 ;
        RECT 41.580 150.450 41.730 158.000 ;
        RECT 42.180 150.450 42.330 158.000 ;
        RECT 42.780 155.150 42.930 158.000 ;
        RECT 43.530 155.600 45.930 158.800 ;
        RECT 49.280 158.650 50.730 158.950 ;
        RECT 46.530 158.450 50.730 158.650 ;
        RECT 58.730 158.950 70.730 159.800 ;
        RECT 58.730 158.900 69.130 158.950 ;
        RECT 58.730 158.650 60.180 158.900 ;
        RECT 60.330 158.800 69.130 158.900 ;
        RECT 58.730 158.450 62.930 158.650 ;
        RECT 46.530 158.300 54.080 158.450 ;
        RECT 55.430 158.300 62.930 158.450 ;
        RECT 46.530 158.000 50.730 158.300 ;
        RECT 46.530 155.150 46.680 158.000 ;
        RECT 47.130 150.450 47.280 158.000 ;
        RECT 47.730 150.450 47.880 158.000 ;
        RECT 48.330 150.450 48.480 158.000 ;
        RECT 48.930 150.450 49.080 158.000 ;
        RECT 49.530 150.450 49.680 158.000 ;
        RECT 50.130 157.850 50.730 158.000 ;
        RECT 58.730 158.000 62.930 158.300 ;
        RECT 58.730 157.850 59.330 158.000 ;
        RECT 50.130 157.700 54.080 157.850 ;
        RECT 55.380 157.700 59.330 157.850 ;
        RECT 50.130 157.250 50.730 157.700 ;
        RECT 58.730 157.250 59.330 157.700 ;
        RECT 50.130 157.100 54.080 157.250 ;
        RECT 55.380 157.100 59.330 157.250 ;
        RECT 50.130 156.650 50.730 157.100 ;
        RECT 58.730 156.650 59.330 157.100 ;
        RECT 50.130 156.500 54.080 156.650 ;
        RECT 55.380 156.500 59.330 156.650 ;
        RECT 50.130 156.050 50.730 156.500 ;
        RECT 58.730 156.050 59.330 156.500 ;
        RECT 50.130 155.900 54.080 156.050 ;
        RECT 55.380 155.900 59.330 156.050 ;
        RECT 50.130 155.450 50.730 155.900 ;
        RECT 58.730 155.450 59.330 155.900 ;
        RECT 50.130 155.300 54.080 155.450 ;
        RECT 55.380 155.300 59.330 155.450 ;
        RECT 50.130 154.850 50.730 155.300 ;
        RECT 58.730 154.850 59.330 155.300 ;
        RECT 50.130 154.700 54.080 154.850 ;
        RECT 55.380 154.700 59.330 154.850 ;
        RECT 50.130 154.250 50.730 154.700 ;
        RECT 58.730 154.250 59.330 154.700 ;
        RECT 50.130 154.100 54.080 154.250 ;
        RECT 55.380 154.100 59.330 154.250 ;
        RECT 50.130 153.650 50.730 154.100 ;
        RECT 58.730 153.650 59.330 154.100 ;
        RECT 50.130 153.500 54.080 153.650 ;
        RECT 55.380 153.500 59.330 153.650 ;
        RECT 50.130 153.050 50.730 153.500 ;
        RECT 58.730 153.050 59.330 153.500 ;
        RECT 50.130 152.900 54.080 153.050 ;
        RECT 55.380 152.900 59.330 153.050 ;
        RECT 50.130 152.450 50.730 152.900 ;
        RECT 58.730 152.450 59.330 152.900 ;
        RECT 50.130 152.300 54.080 152.450 ;
        RECT 55.380 152.300 59.330 152.450 ;
        RECT 50.130 151.850 50.730 152.300 ;
        RECT 58.730 151.850 59.330 152.300 ;
        RECT 50.130 151.700 54.080 151.850 ;
        RECT 55.380 151.700 59.330 151.850 ;
        RECT 50.130 151.250 50.730 151.700 ;
        RECT 58.730 151.250 59.330 151.700 ;
        RECT 50.130 151.100 54.080 151.250 ;
        RECT 55.380 151.100 59.330 151.250 ;
        RECT 50.130 150.650 50.730 151.100 ;
        RECT 58.730 150.650 59.330 151.100 ;
        RECT 50.130 150.450 54.080 150.650 ;
        RECT 55.380 150.450 59.330 150.650 ;
        RECT 59.780 150.450 59.930 158.000 ;
        RECT 60.380 150.450 60.530 158.000 ;
        RECT 60.980 150.450 61.130 158.000 ;
        RECT 61.580 150.450 61.730 158.000 ;
        RECT 62.180 150.450 62.330 158.000 ;
        RECT 62.780 155.150 62.930 158.000 ;
        RECT 63.530 155.600 65.930 158.800 ;
        RECT 69.280 158.650 70.730 158.950 ;
        RECT 66.530 158.450 70.730 158.650 ;
        RECT 78.730 158.950 90.730 159.800 ;
        RECT 78.730 158.900 89.130 158.950 ;
        RECT 78.730 158.650 80.180 158.900 ;
        RECT 80.330 158.800 89.130 158.900 ;
        RECT 78.730 158.450 82.930 158.650 ;
        RECT 66.530 158.300 74.080 158.450 ;
        RECT 75.430 158.300 82.930 158.450 ;
        RECT 66.530 158.000 70.730 158.300 ;
        RECT 66.530 155.150 66.680 158.000 ;
        RECT 67.130 150.450 67.280 158.000 ;
        RECT 67.730 150.450 67.880 158.000 ;
        RECT 68.330 150.450 68.480 158.000 ;
        RECT 68.930 150.450 69.080 158.000 ;
        RECT 69.530 150.450 69.680 158.000 ;
        RECT 70.130 157.850 70.730 158.000 ;
        RECT 78.730 158.000 82.930 158.300 ;
        RECT 78.730 157.850 79.330 158.000 ;
        RECT 70.130 157.700 74.080 157.850 ;
        RECT 75.380 157.700 79.330 157.850 ;
        RECT 70.130 157.250 70.730 157.700 ;
        RECT 78.730 157.250 79.330 157.700 ;
        RECT 70.130 157.100 74.080 157.250 ;
        RECT 75.380 157.100 79.330 157.250 ;
        RECT 70.130 156.650 70.730 157.100 ;
        RECT 78.730 156.650 79.330 157.100 ;
        RECT 70.130 156.500 74.080 156.650 ;
        RECT 75.380 156.500 79.330 156.650 ;
        RECT 70.130 156.050 70.730 156.500 ;
        RECT 78.730 156.050 79.330 156.500 ;
        RECT 70.130 155.900 74.080 156.050 ;
        RECT 75.380 155.900 79.330 156.050 ;
        RECT 70.130 155.450 70.730 155.900 ;
        RECT 78.730 155.450 79.330 155.900 ;
        RECT 70.130 155.300 74.080 155.450 ;
        RECT 75.380 155.300 79.330 155.450 ;
        RECT 70.130 154.850 70.730 155.300 ;
        RECT 78.730 154.850 79.330 155.300 ;
        RECT 70.130 154.700 74.080 154.850 ;
        RECT 75.380 154.700 79.330 154.850 ;
        RECT 70.130 154.250 70.730 154.700 ;
        RECT 78.730 154.250 79.330 154.700 ;
        RECT 70.130 154.100 74.080 154.250 ;
        RECT 75.380 154.100 79.330 154.250 ;
        RECT 70.130 153.650 70.730 154.100 ;
        RECT 78.730 153.650 79.330 154.100 ;
        RECT 70.130 153.500 74.080 153.650 ;
        RECT 75.380 153.500 79.330 153.650 ;
        RECT 70.130 153.050 70.730 153.500 ;
        RECT 78.730 153.050 79.330 153.500 ;
        RECT 70.130 152.900 74.080 153.050 ;
        RECT 75.380 152.900 79.330 153.050 ;
        RECT 70.130 152.450 70.730 152.900 ;
        RECT 78.730 152.450 79.330 152.900 ;
        RECT 70.130 152.300 74.080 152.450 ;
        RECT 75.380 152.300 79.330 152.450 ;
        RECT 70.130 151.850 70.730 152.300 ;
        RECT 78.730 151.850 79.330 152.300 ;
        RECT 70.130 151.700 74.080 151.850 ;
        RECT 75.380 151.700 79.330 151.850 ;
        RECT 70.130 151.250 70.730 151.700 ;
        RECT 78.730 151.250 79.330 151.700 ;
        RECT 70.130 151.100 74.080 151.250 ;
        RECT 75.380 151.100 79.330 151.250 ;
        RECT 70.130 150.650 70.730 151.100 ;
        RECT 78.730 150.650 79.330 151.100 ;
        RECT 70.130 150.450 74.080 150.650 ;
        RECT 75.380 150.450 79.330 150.650 ;
        RECT 79.780 150.450 79.930 158.000 ;
        RECT 80.380 150.450 80.530 158.000 ;
        RECT 80.980 150.450 81.130 158.000 ;
        RECT 81.580 150.450 81.730 158.000 ;
        RECT 82.180 150.450 82.330 158.000 ;
        RECT 82.780 155.150 82.930 158.000 ;
        RECT 83.530 155.600 85.930 158.800 ;
        RECT 89.280 158.650 90.730 158.950 ;
        RECT 86.530 158.450 90.730 158.650 ;
        RECT 98.730 158.900 104.730 159.800 ;
        RECT 98.730 158.650 100.180 158.900 ;
        RECT 100.330 158.800 104.730 158.900 ;
        RECT 98.730 158.450 102.930 158.650 ;
        RECT 86.530 158.300 94.080 158.450 ;
        RECT 95.430 158.300 102.930 158.450 ;
        RECT 86.530 158.000 90.730 158.300 ;
        RECT 86.530 155.150 86.680 158.000 ;
        RECT 87.130 150.450 87.280 158.000 ;
        RECT 87.730 150.450 87.880 158.000 ;
        RECT 88.330 150.450 88.480 158.000 ;
        RECT 88.930 150.450 89.080 158.000 ;
        RECT 89.530 150.450 89.680 158.000 ;
        RECT 90.130 157.850 90.730 158.000 ;
        RECT 98.730 158.000 102.930 158.300 ;
        RECT 98.730 157.850 99.330 158.000 ;
        RECT 90.130 157.700 94.080 157.850 ;
        RECT 95.380 157.700 99.330 157.850 ;
        RECT 90.130 157.250 90.730 157.700 ;
        RECT 98.730 157.250 99.330 157.700 ;
        RECT 90.130 157.100 94.080 157.250 ;
        RECT 95.380 157.100 99.330 157.250 ;
        RECT 90.130 156.650 90.730 157.100 ;
        RECT 98.730 156.650 99.330 157.100 ;
        RECT 90.130 156.500 94.080 156.650 ;
        RECT 95.380 156.500 99.330 156.650 ;
        RECT 90.130 156.050 90.730 156.500 ;
        RECT 98.730 156.050 99.330 156.500 ;
        RECT 90.130 155.900 94.080 156.050 ;
        RECT 95.380 155.900 99.330 156.050 ;
        RECT 90.130 155.450 90.730 155.900 ;
        RECT 98.730 155.450 99.330 155.900 ;
        RECT 90.130 155.300 94.080 155.450 ;
        RECT 95.380 155.300 99.330 155.450 ;
        RECT 90.130 154.850 90.730 155.300 ;
        RECT 98.730 154.850 99.330 155.300 ;
        RECT 90.130 154.700 94.080 154.850 ;
        RECT 95.380 154.700 99.330 154.850 ;
        RECT 90.130 154.250 90.730 154.700 ;
        RECT 98.730 154.250 99.330 154.700 ;
        RECT 90.130 154.100 94.080 154.250 ;
        RECT 95.380 154.100 99.330 154.250 ;
        RECT 90.130 153.650 90.730 154.100 ;
        RECT 98.730 153.650 99.330 154.100 ;
        RECT 90.130 153.500 94.080 153.650 ;
        RECT 95.380 153.500 99.330 153.650 ;
        RECT 90.130 153.050 90.730 153.500 ;
        RECT 98.730 153.050 99.330 153.500 ;
        RECT 90.130 152.900 94.080 153.050 ;
        RECT 95.380 152.900 99.330 153.050 ;
        RECT 90.130 152.450 90.730 152.900 ;
        RECT 98.730 152.450 99.330 152.900 ;
        RECT 90.130 152.300 94.080 152.450 ;
        RECT 95.380 152.300 99.330 152.450 ;
        RECT 90.130 151.850 90.730 152.300 ;
        RECT 98.730 151.850 99.330 152.300 ;
        RECT 90.130 151.700 94.080 151.850 ;
        RECT 95.380 151.700 99.330 151.850 ;
        RECT 90.130 151.250 90.730 151.700 ;
        RECT 98.730 151.250 99.330 151.700 ;
        RECT 90.130 151.100 94.080 151.250 ;
        RECT 95.380 151.100 99.330 151.250 ;
        RECT 90.130 150.650 90.730 151.100 ;
        RECT 98.730 150.650 99.330 151.100 ;
        RECT 90.130 150.450 94.080 150.650 ;
        RECT 95.380 150.450 99.330 150.650 ;
        RECT 99.780 150.450 99.930 158.000 ;
        RECT 100.380 150.450 100.530 158.000 ;
        RECT 100.980 150.450 101.130 158.000 ;
        RECT 101.580 150.450 101.730 158.000 ;
        RECT 102.180 150.450 102.330 158.000 ;
        RECT 102.780 155.150 102.930 158.000 ;
        RECT 103.530 157.725 104.730 158.800 ;
        RECT 103.530 156.450 107.140 157.725 ;
        RECT 103.530 155.600 104.730 156.450 ;
        RECT 2.315 144.450 4.315 146.750 ;
        RECT 4.730 143.165 5.930 144.400 ;
        RECT 2.315 141.890 5.930 143.165 ;
        RECT 4.730 141.200 5.930 141.890 ;
        RECT 6.530 142.000 6.680 144.900 ;
        RECT 7.130 142.000 7.280 149.550 ;
        RECT 7.730 142.000 7.880 149.550 ;
        RECT 8.330 142.000 8.480 149.550 ;
        RECT 8.930 142.000 9.080 149.550 ;
        RECT 9.530 142.000 9.680 149.550 ;
        RECT 10.130 149.350 14.080 149.550 ;
        RECT 15.380 149.350 19.330 149.550 ;
        RECT 10.130 148.900 10.730 149.350 ;
        RECT 18.730 148.900 19.330 149.350 ;
        RECT 10.130 148.750 14.080 148.900 ;
        RECT 15.380 148.750 19.330 148.900 ;
        RECT 10.130 148.300 10.730 148.750 ;
        RECT 18.730 148.300 19.330 148.750 ;
        RECT 10.130 148.150 14.080 148.300 ;
        RECT 15.380 148.150 19.330 148.300 ;
        RECT 10.130 147.700 10.730 148.150 ;
        RECT 18.730 147.700 19.330 148.150 ;
        RECT 10.130 147.550 14.080 147.700 ;
        RECT 15.380 147.550 19.330 147.700 ;
        RECT 10.130 147.100 10.730 147.550 ;
        RECT 18.730 147.100 19.330 147.550 ;
        RECT 10.130 146.950 14.080 147.100 ;
        RECT 15.380 146.950 19.330 147.100 ;
        RECT 10.130 146.500 10.730 146.950 ;
        RECT 18.730 146.500 19.330 146.950 ;
        RECT 10.130 146.350 14.080 146.500 ;
        RECT 15.380 146.350 19.330 146.500 ;
        RECT 10.130 145.900 10.730 146.350 ;
        RECT 18.730 145.900 19.330 146.350 ;
        RECT 10.130 145.750 14.080 145.900 ;
        RECT 15.380 145.750 19.330 145.900 ;
        RECT 10.130 145.300 10.730 145.750 ;
        RECT 18.730 145.300 19.330 145.750 ;
        RECT 10.130 145.150 14.080 145.300 ;
        RECT 15.380 145.150 19.330 145.300 ;
        RECT 10.130 144.700 10.730 145.150 ;
        RECT 18.730 144.700 19.330 145.150 ;
        RECT 10.130 144.550 14.080 144.700 ;
        RECT 15.380 144.550 19.330 144.700 ;
        RECT 10.130 144.100 10.730 144.550 ;
        RECT 18.730 144.100 19.330 144.550 ;
        RECT 10.130 143.950 14.080 144.100 ;
        RECT 15.380 143.950 19.330 144.100 ;
        RECT 10.130 143.500 10.730 143.950 ;
        RECT 18.730 143.500 19.330 143.950 ;
        RECT 10.130 143.350 14.080 143.500 ;
        RECT 15.380 143.350 19.330 143.500 ;
        RECT 10.130 142.900 10.730 143.350 ;
        RECT 18.730 142.900 19.330 143.350 ;
        RECT 10.130 142.750 14.080 142.900 ;
        RECT 15.380 142.750 19.330 142.900 ;
        RECT 10.130 142.300 10.730 142.750 ;
        RECT 18.730 142.300 19.330 142.750 ;
        RECT 10.130 142.150 14.080 142.300 ;
        RECT 15.380 142.150 19.330 142.300 ;
        RECT 10.130 142.000 10.730 142.150 ;
        RECT 6.530 141.700 10.730 142.000 ;
        RECT 18.730 142.000 19.330 142.150 ;
        RECT 19.780 142.000 19.930 149.550 ;
        RECT 20.380 142.000 20.530 149.550 ;
        RECT 20.980 142.000 21.130 149.550 ;
        RECT 21.580 142.000 21.730 149.550 ;
        RECT 22.180 142.000 22.330 149.550 ;
        RECT 22.780 142.000 22.930 144.900 ;
        RECT 18.730 141.700 22.930 142.000 ;
        RECT 6.530 141.550 14.080 141.700 ;
        RECT 15.380 141.550 22.930 141.700 ;
        RECT 6.530 141.350 10.730 141.550 ;
        RECT 4.730 141.050 9.130 141.200 ;
        RECT 9.280 141.050 10.730 141.350 ;
        RECT 4.730 140.150 10.730 141.050 ;
        RECT 18.730 141.350 22.930 141.550 ;
        RECT 18.730 141.050 20.180 141.350 ;
        RECT 23.530 141.200 25.930 144.400 ;
        RECT 26.530 142.000 26.680 144.900 ;
        RECT 27.130 142.000 27.280 149.550 ;
        RECT 27.730 142.000 27.880 149.550 ;
        RECT 28.330 142.000 28.480 149.550 ;
        RECT 28.930 142.000 29.080 149.550 ;
        RECT 29.530 142.000 29.680 149.550 ;
        RECT 30.130 149.350 34.080 149.550 ;
        RECT 35.380 149.350 39.330 149.550 ;
        RECT 30.130 148.900 30.730 149.350 ;
        RECT 38.730 148.900 39.330 149.350 ;
        RECT 30.130 148.750 34.080 148.900 ;
        RECT 35.380 148.750 39.330 148.900 ;
        RECT 30.130 148.300 30.730 148.750 ;
        RECT 38.730 148.300 39.330 148.750 ;
        RECT 30.130 148.150 34.080 148.300 ;
        RECT 35.380 148.150 39.330 148.300 ;
        RECT 30.130 147.700 30.730 148.150 ;
        RECT 38.730 147.700 39.330 148.150 ;
        RECT 30.130 147.550 34.080 147.700 ;
        RECT 35.380 147.550 39.330 147.700 ;
        RECT 30.130 147.100 30.730 147.550 ;
        RECT 38.730 147.100 39.330 147.550 ;
        RECT 30.130 146.950 34.080 147.100 ;
        RECT 35.380 146.950 39.330 147.100 ;
        RECT 30.130 146.500 30.730 146.950 ;
        RECT 38.730 146.500 39.330 146.950 ;
        RECT 30.130 146.350 34.080 146.500 ;
        RECT 35.380 146.350 39.330 146.500 ;
        RECT 30.130 145.900 30.730 146.350 ;
        RECT 38.730 145.900 39.330 146.350 ;
        RECT 30.130 145.750 34.080 145.900 ;
        RECT 35.380 145.750 39.330 145.900 ;
        RECT 30.130 145.300 30.730 145.750 ;
        RECT 38.730 145.300 39.330 145.750 ;
        RECT 30.130 145.150 34.080 145.300 ;
        RECT 35.380 145.150 39.330 145.300 ;
        RECT 30.130 144.700 30.730 145.150 ;
        RECT 38.730 144.700 39.330 145.150 ;
        RECT 30.130 144.550 34.080 144.700 ;
        RECT 35.380 144.550 39.330 144.700 ;
        RECT 30.130 144.100 30.730 144.550 ;
        RECT 38.730 144.100 39.330 144.550 ;
        RECT 30.130 143.950 34.080 144.100 ;
        RECT 35.380 143.950 39.330 144.100 ;
        RECT 30.130 143.500 30.730 143.950 ;
        RECT 38.730 143.500 39.330 143.950 ;
        RECT 30.130 143.350 34.080 143.500 ;
        RECT 35.380 143.350 39.330 143.500 ;
        RECT 30.130 142.900 30.730 143.350 ;
        RECT 38.730 142.900 39.330 143.350 ;
        RECT 30.130 142.750 34.080 142.900 ;
        RECT 35.380 142.750 39.330 142.900 ;
        RECT 30.130 142.300 30.730 142.750 ;
        RECT 38.730 142.300 39.330 142.750 ;
        RECT 30.130 142.150 34.080 142.300 ;
        RECT 35.380 142.150 39.330 142.300 ;
        RECT 30.130 142.000 30.730 142.150 ;
        RECT 26.530 141.700 30.730 142.000 ;
        RECT 38.730 142.000 39.330 142.150 ;
        RECT 39.780 142.000 39.930 149.550 ;
        RECT 40.380 142.000 40.530 149.550 ;
        RECT 40.980 142.000 41.130 149.550 ;
        RECT 41.580 142.000 41.730 149.550 ;
        RECT 42.180 142.000 42.330 149.550 ;
        RECT 42.780 142.000 42.930 144.900 ;
        RECT 38.730 141.700 42.930 142.000 ;
        RECT 26.530 141.550 34.080 141.700 ;
        RECT 35.380 141.550 42.930 141.700 ;
        RECT 26.530 141.350 30.730 141.550 ;
        RECT 20.330 141.050 29.130 141.200 ;
        RECT 29.280 141.050 30.730 141.350 ;
        RECT 18.730 140.150 30.730 141.050 ;
        RECT 38.730 141.350 42.930 141.550 ;
        RECT 38.730 141.050 40.180 141.350 ;
        RECT 43.530 141.200 45.930 144.400 ;
        RECT 46.530 142.000 46.680 144.900 ;
        RECT 47.130 142.000 47.280 149.550 ;
        RECT 47.730 142.000 47.880 149.550 ;
        RECT 48.330 142.000 48.480 149.550 ;
        RECT 48.930 142.000 49.080 149.550 ;
        RECT 49.530 142.000 49.680 149.550 ;
        RECT 50.130 149.350 54.080 149.550 ;
        RECT 55.380 149.350 59.330 149.550 ;
        RECT 50.130 148.900 50.730 149.350 ;
        RECT 58.730 148.900 59.330 149.350 ;
        RECT 50.130 148.750 54.080 148.900 ;
        RECT 55.380 148.750 59.330 148.900 ;
        RECT 50.130 148.300 50.730 148.750 ;
        RECT 58.730 148.300 59.330 148.750 ;
        RECT 50.130 148.150 54.080 148.300 ;
        RECT 55.380 148.150 59.330 148.300 ;
        RECT 50.130 147.700 50.730 148.150 ;
        RECT 58.730 147.700 59.330 148.150 ;
        RECT 50.130 147.550 54.080 147.700 ;
        RECT 55.380 147.550 59.330 147.700 ;
        RECT 50.130 147.100 50.730 147.550 ;
        RECT 58.730 147.100 59.330 147.550 ;
        RECT 50.130 146.950 54.080 147.100 ;
        RECT 55.380 146.950 59.330 147.100 ;
        RECT 50.130 146.500 50.730 146.950 ;
        RECT 58.730 146.500 59.330 146.950 ;
        RECT 50.130 146.350 54.080 146.500 ;
        RECT 55.380 146.350 59.330 146.500 ;
        RECT 50.130 145.900 50.730 146.350 ;
        RECT 58.730 145.900 59.330 146.350 ;
        RECT 50.130 145.750 54.080 145.900 ;
        RECT 55.380 145.750 59.330 145.900 ;
        RECT 50.130 145.300 50.730 145.750 ;
        RECT 58.730 145.300 59.330 145.750 ;
        RECT 50.130 145.150 54.080 145.300 ;
        RECT 55.380 145.150 59.330 145.300 ;
        RECT 50.130 144.700 50.730 145.150 ;
        RECT 58.730 144.700 59.330 145.150 ;
        RECT 50.130 144.550 54.080 144.700 ;
        RECT 55.380 144.550 59.330 144.700 ;
        RECT 50.130 144.100 50.730 144.550 ;
        RECT 58.730 144.100 59.330 144.550 ;
        RECT 50.130 143.950 54.080 144.100 ;
        RECT 55.380 143.950 59.330 144.100 ;
        RECT 50.130 143.500 50.730 143.950 ;
        RECT 58.730 143.500 59.330 143.950 ;
        RECT 50.130 143.350 54.080 143.500 ;
        RECT 55.380 143.350 59.330 143.500 ;
        RECT 50.130 142.900 50.730 143.350 ;
        RECT 58.730 142.900 59.330 143.350 ;
        RECT 50.130 142.750 54.080 142.900 ;
        RECT 55.380 142.750 59.330 142.900 ;
        RECT 50.130 142.300 50.730 142.750 ;
        RECT 58.730 142.300 59.330 142.750 ;
        RECT 50.130 142.150 54.080 142.300 ;
        RECT 55.380 142.150 59.330 142.300 ;
        RECT 50.130 142.000 50.730 142.150 ;
        RECT 46.530 141.700 50.730 142.000 ;
        RECT 58.730 142.000 59.330 142.150 ;
        RECT 59.780 142.000 59.930 149.550 ;
        RECT 60.380 142.000 60.530 149.550 ;
        RECT 60.980 142.000 61.130 149.550 ;
        RECT 61.580 142.000 61.730 149.550 ;
        RECT 62.180 142.000 62.330 149.550 ;
        RECT 62.780 142.000 62.930 144.900 ;
        RECT 58.730 141.700 62.930 142.000 ;
        RECT 46.530 141.550 54.080 141.700 ;
        RECT 55.380 141.550 62.930 141.700 ;
        RECT 46.530 141.350 50.730 141.550 ;
        RECT 40.330 141.050 49.130 141.200 ;
        RECT 49.280 141.050 50.730 141.350 ;
        RECT 38.730 140.150 50.730 141.050 ;
        RECT 58.730 141.350 62.930 141.550 ;
        RECT 58.730 141.050 60.180 141.350 ;
        RECT 63.530 141.200 65.930 144.400 ;
        RECT 66.530 142.000 66.680 144.900 ;
        RECT 67.130 142.000 67.280 149.550 ;
        RECT 67.730 142.000 67.880 149.550 ;
        RECT 68.330 142.000 68.480 149.550 ;
        RECT 68.930 142.000 69.080 149.550 ;
        RECT 69.530 142.000 69.680 149.550 ;
        RECT 70.130 149.350 74.080 149.550 ;
        RECT 75.380 149.350 79.330 149.550 ;
        RECT 70.130 148.900 70.730 149.350 ;
        RECT 78.730 148.900 79.330 149.350 ;
        RECT 70.130 148.750 74.080 148.900 ;
        RECT 75.380 148.750 79.330 148.900 ;
        RECT 70.130 148.300 70.730 148.750 ;
        RECT 78.730 148.300 79.330 148.750 ;
        RECT 70.130 148.150 74.080 148.300 ;
        RECT 75.380 148.150 79.330 148.300 ;
        RECT 70.130 147.700 70.730 148.150 ;
        RECT 78.730 147.700 79.330 148.150 ;
        RECT 70.130 147.550 74.080 147.700 ;
        RECT 75.380 147.550 79.330 147.700 ;
        RECT 70.130 147.100 70.730 147.550 ;
        RECT 78.730 147.100 79.330 147.550 ;
        RECT 70.130 146.950 74.080 147.100 ;
        RECT 75.380 146.950 79.330 147.100 ;
        RECT 70.130 146.500 70.730 146.950 ;
        RECT 78.730 146.500 79.330 146.950 ;
        RECT 70.130 146.350 74.080 146.500 ;
        RECT 75.380 146.350 79.330 146.500 ;
        RECT 70.130 145.900 70.730 146.350 ;
        RECT 78.730 145.900 79.330 146.350 ;
        RECT 70.130 145.750 74.080 145.900 ;
        RECT 75.380 145.750 79.330 145.900 ;
        RECT 70.130 145.300 70.730 145.750 ;
        RECT 78.730 145.300 79.330 145.750 ;
        RECT 70.130 145.150 74.080 145.300 ;
        RECT 75.380 145.150 79.330 145.300 ;
        RECT 70.130 144.700 70.730 145.150 ;
        RECT 78.730 144.700 79.330 145.150 ;
        RECT 70.130 144.550 74.080 144.700 ;
        RECT 75.380 144.550 79.330 144.700 ;
        RECT 70.130 144.100 70.730 144.550 ;
        RECT 78.730 144.100 79.330 144.550 ;
        RECT 70.130 143.950 74.080 144.100 ;
        RECT 75.380 143.950 79.330 144.100 ;
        RECT 70.130 143.500 70.730 143.950 ;
        RECT 78.730 143.500 79.330 143.950 ;
        RECT 70.130 143.350 74.080 143.500 ;
        RECT 75.380 143.350 79.330 143.500 ;
        RECT 70.130 142.900 70.730 143.350 ;
        RECT 78.730 142.900 79.330 143.350 ;
        RECT 70.130 142.750 74.080 142.900 ;
        RECT 75.380 142.750 79.330 142.900 ;
        RECT 70.130 142.300 70.730 142.750 ;
        RECT 78.730 142.300 79.330 142.750 ;
        RECT 70.130 142.150 74.080 142.300 ;
        RECT 75.380 142.150 79.330 142.300 ;
        RECT 70.130 142.000 70.730 142.150 ;
        RECT 66.530 141.700 70.730 142.000 ;
        RECT 78.730 142.000 79.330 142.150 ;
        RECT 79.780 142.000 79.930 149.550 ;
        RECT 80.380 142.000 80.530 149.550 ;
        RECT 80.980 142.000 81.130 149.550 ;
        RECT 81.580 142.000 81.730 149.550 ;
        RECT 82.180 142.000 82.330 149.550 ;
        RECT 82.780 142.000 82.930 144.900 ;
        RECT 78.730 141.700 82.930 142.000 ;
        RECT 66.530 141.550 74.080 141.700 ;
        RECT 75.380 141.550 82.930 141.700 ;
        RECT 66.530 141.350 70.730 141.550 ;
        RECT 60.330 141.050 69.130 141.200 ;
        RECT 69.280 141.050 70.730 141.350 ;
        RECT 58.730 140.150 70.730 141.050 ;
        RECT 78.730 141.350 82.930 141.550 ;
        RECT 78.730 141.050 80.180 141.350 ;
        RECT 83.530 141.200 85.930 144.400 ;
        RECT 86.530 142.000 86.680 144.900 ;
        RECT 87.130 142.000 87.280 149.550 ;
        RECT 87.730 142.000 87.880 149.550 ;
        RECT 88.330 142.000 88.480 149.550 ;
        RECT 88.930 142.000 89.080 149.550 ;
        RECT 89.530 142.000 89.680 149.550 ;
        RECT 90.130 149.350 94.080 149.550 ;
        RECT 95.380 149.350 99.330 149.550 ;
        RECT 90.130 148.900 90.730 149.350 ;
        RECT 98.730 148.900 99.330 149.350 ;
        RECT 90.130 148.750 94.080 148.900 ;
        RECT 95.380 148.750 99.330 148.900 ;
        RECT 90.130 148.300 90.730 148.750 ;
        RECT 98.730 148.300 99.330 148.750 ;
        RECT 90.130 148.150 94.080 148.300 ;
        RECT 95.380 148.150 99.330 148.300 ;
        RECT 90.130 147.700 90.730 148.150 ;
        RECT 98.730 147.700 99.330 148.150 ;
        RECT 90.130 147.550 94.080 147.700 ;
        RECT 95.380 147.550 99.330 147.700 ;
        RECT 90.130 147.100 90.730 147.550 ;
        RECT 98.730 147.100 99.330 147.550 ;
        RECT 90.130 146.950 94.080 147.100 ;
        RECT 95.380 146.950 99.330 147.100 ;
        RECT 90.130 146.500 90.730 146.950 ;
        RECT 98.730 146.500 99.330 146.950 ;
        RECT 90.130 146.350 94.080 146.500 ;
        RECT 95.380 146.350 99.330 146.500 ;
        RECT 90.130 145.900 90.730 146.350 ;
        RECT 98.730 145.900 99.330 146.350 ;
        RECT 90.130 145.750 94.080 145.900 ;
        RECT 95.380 145.750 99.330 145.900 ;
        RECT 90.130 145.300 90.730 145.750 ;
        RECT 98.730 145.300 99.330 145.750 ;
        RECT 90.130 145.150 94.080 145.300 ;
        RECT 95.380 145.150 99.330 145.300 ;
        RECT 90.130 144.700 90.730 145.150 ;
        RECT 98.730 144.700 99.330 145.150 ;
        RECT 90.130 144.550 94.080 144.700 ;
        RECT 95.380 144.550 99.330 144.700 ;
        RECT 90.130 144.100 90.730 144.550 ;
        RECT 98.730 144.100 99.330 144.550 ;
        RECT 90.130 143.950 94.080 144.100 ;
        RECT 95.380 143.950 99.330 144.100 ;
        RECT 90.130 143.500 90.730 143.950 ;
        RECT 98.730 143.500 99.330 143.950 ;
        RECT 90.130 143.350 94.080 143.500 ;
        RECT 95.380 143.350 99.330 143.500 ;
        RECT 90.130 142.900 90.730 143.350 ;
        RECT 98.730 142.900 99.330 143.350 ;
        RECT 90.130 142.750 94.080 142.900 ;
        RECT 95.380 142.750 99.330 142.900 ;
        RECT 90.130 142.300 90.730 142.750 ;
        RECT 98.730 142.300 99.330 142.750 ;
        RECT 90.130 142.150 94.080 142.300 ;
        RECT 95.380 142.150 99.330 142.300 ;
        RECT 90.130 142.000 90.730 142.150 ;
        RECT 86.530 141.700 90.730 142.000 ;
        RECT 98.730 142.000 99.330 142.150 ;
        RECT 99.780 142.000 99.930 149.550 ;
        RECT 100.380 142.000 100.530 149.550 ;
        RECT 100.980 142.000 101.130 149.550 ;
        RECT 101.580 142.000 101.730 149.550 ;
        RECT 102.180 142.000 102.330 149.550 ;
        RECT 102.780 142.000 102.930 144.900 ;
        RECT 98.730 141.700 102.930 142.000 ;
        RECT 86.530 141.550 94.080 141.700 ;
        RECT 95.380 141.550 102.930 141.700 ;
        RECT 86.530 141.350 90.730 141.550 ;
        RECT 80.330 141.050 89.130 141.200 ;
        RECT 89.280 141.050 90.730 141.350 ;
        RECT 78.730 140.150 90.730 141.050 ;
        RECT 98.730 141.350 102.930 141.550 ;
        RECT 103.530 142.920 104.730 144.400 ;
        RECT 103.530 141.645 107.140 142.920 ;
        RECT 98.730 141.050 100.180 141.350 ;
        RECT 103.530 141.200 104.730 141.645 ;
        RECT 100.330 141.050 104.730 141.200 ;
        RECT 98.730 140.150 104.730 141.050 ;
        RECT 4.730 139.850 9.130 140.150 ;
        RECT 20.330 139.850 29.130 140.150 ;
        RECT 40.330 139.850 49.130 140.150 ;
        RECT 60.330 139.850 69.130 140.150 ;
        RECT 80.330 139.850 89.130 140.150 ;
        RECT 4.730 138.950 10.730 139.850 ;
        RECT 20.330 139.800 30.730 139.850 ;
        RECT 40.330 139.800 50.730 139.850 ;
        RECT 60.330 139.800 70.730 139.850 ;
        RECT 80.330 139.800 90.730 139.850 ;
        RECT 100.330 139.800 104.730 140.150 ;
        RECT 4.730 138.800 9.130 138.950 ;
        RECT 4.730 138.145 5.930 138.800 ;
        RECT 9.280 138.650 10.730 138.950 ;
        RECT 2.315 136.870 5.930 138.145 ;
        RECT 4.730 135.600 5.930 136.870 ;
        RECT 6.530 138.450 10.730 138.650 ;
        RECT 18.730 138.950 30.730 139.800 ;
        RECT 18.730 138.900 29.130 138.950 ;
        RECT 18.730 138.650 20.180 138.900 ;
        RECT 20.330 138.800 29.130 138.900 ;
        RECT 18.730 138.450 22.930 138.650 ;
        RECT 6.530 138.300 14.080 138.450 ;
        RECT 15.430 138.300 22.930 138.450 ;
        RECT 6.530 138.000 10.730 138.300 ;
        RECT 2.315 133.250 4.315 135.545 ;
        RECT 6.530 135.150 6.680 138.000 ;
        RECT 7.130 130.450 7.280 138.000 ;
        RECT 7.730 130.450 7.880 138.000 ;
        RECT 8.330 130.450 8.480 138.000 ;
        RECT 8.930 130.450 9.080 138.000 ;
        RECT 9.530 130.450 9.680 138.000 ;
        RECT 10.130 137.850 10.730 138.000 ;
        RECT 18.730 138.000 22.930 138.300 ;
        RECT 18.730 137.850 19.330 138.000 ;
        RECT 10.130 137.700 14.080 137.850 ;
        RECT 15.380 137.700 19.330 137.850 ;
        RECT 10.130 137.250 10.730 137.700 ;
        RECT 18.730 137.250 19.330 137.700 ;
        RECT 10.130 137.100 14.080 137.250 ;
        RECT 15.380 137.100 19.330 137.250 ;
        RECT 10.130 136.650 10.730 137.100 ;
        RECT 18.730 136.650 19.330 137.100 ;
        RECT 10.130 136.500 14.080 136.650 ;
        RECT 15.380 136.500 19.330 136.650 ;
        RECT 10.130 136.050 10.730 136.500 ;
        RECT 18.730 136.050 19.330 136.500 ;
        RECT 10.130 135.900 14.080 136.050 ;
        RECT 15.380 135.900 19.330 136.050 ;
        RECT 10.130 135.450 10.730 135.900 ;
        RECT 18.730 135.450 19.330 135.900 ;
        RECT 10.130 135.300 14.080 135.450 ;
        RECT 15.380 135.300 19.330 135.450 ;
        RECT 10.130 134.850 10.730 135.300 ;
        RECT 18.730 134.850 19.330 135.300 ;
        RECT 10.130 134.700 14.080 134.850 ;
        RECT 15.380 134.700 19.330 134.850 ;
        RECT 10.130 134.250 10.730 134.700 ;
        RECT 18.730 134.250 19.330 134.700 ;
        RECT 10.130 134.100 14.080 134.250 ;
        RECT 15.380 134.100 19.330 134.250 ;
        RECT 10.130 133.650 10.730 134.100 ;
        RECT 18.730 133.650 19.330 134.100 ;
        RECT 10.130 133.500 14.080 133.650 ;
        RECT 15.380 133.500 19.330 133.650 ;
        RECT 10.130 133.050 10.730 133.500 ;
        RECT 18.730 133.050 19.330 133.500 ;
        RECT 10.130 132.900 14.080 133.050 ;
        RECT 15.380 132.900 19.330 133.050 ;
        RECT 10.130 132.450 10.730 132.900 ;
        RECT 18.730 132.450 19.330 132.900 ;
        RECT 10.130 132.300 14.080 132.450 ;
        RECT 15.380 132.300 19.330 132.450 ;
        RECT 10.130 131.850 10.730 132.300 ;
        RECT 18.730 131.850 19.330 132.300 ;
        RECT 10.130 131.700 14.080 131.850 ;
        RECT 15.380 131.700 19.330 131.850 ;
        RECT 10.130 131.250 10.730 131.700 ;
        RECT 18.730 131.250 19.330 131.700 ;
        RECT 10.130 131.100 14.080 131.250 ;
        RECT 15.380 131.100 19.330 131.250 ;
        RECT 10.130 130.650 10.730 131.100 ;
        RECT 18.730 130.650 19.330 131.100 ;
        RECT 10.130 130.450 14.080 130.650 ;
        RECT 15.380 130.450 19.330 130.650 ;
        RECT 19.780 130.450 19.930 138.000 ;
        RECT 20.380 130.450 20.530 138.000 ;
        RECT 20.980 130.450 21.130 138.000 ;
        RECT 21.580 130.450 21.730 138.000 ;
        RECT 22.180 130.450 22.330 138.000 ;
        RECT 22.780 135.150 22.930 138.000 ;
        RECT 23.530 135.600 25.930 138.800 ;
        RECT 29.280 138.650 30.730 138.950 ;
        RECT 26.530 138.450 30.730 138.650 ;
        RECT 38.730 138.950 50.730 139.800 ;
        RECT 38.730 138.900 49.130 138.950 ;
        RECT 38.730 138.650 40.180 138.900 ;
        RECT 40.330 138.800 49.130 138.900 ;
        RECT 38.730 138.450 42.930 138.650 ;
        RECT 26.530 138.300 34.080 138.450 ;
        RECT 35.430 138.300 42.930 138.450 ;
        RECT 26.530 138.000 30.730 138.300 ;
        RECT 26.530 135.150 26.680 138.000 ;
        RECT 27.130 130.450 27.280 138.000 ;
        RECT 27.730 130.450 27.880 138.000 ;
        RECT 28.330 130.450 28.480 138.000 ;
        RECT 28.930 130.450 29.080 138.000 ;
        RECT 29.530 130.450 29.680 138.000 ;
        RECT 30.130 137.850 30.730 138.000 ;
        RECT 38.730 138.000 42.930 138.300 ;
        RECT 38.730 137.850 39.330 138.000 ;
        RECT 30.130 137.700 34.080 137.850 ;
        RECT 35.380 137.700 39.330 137.850 ;
        RECT 30.130 137.250 30.730 137.700 ;
        RECT 38.730 137.250 39.330 137.700 ;
        RECT 30.130 137.100 34.080 137.250 ;
        RECT 35.380 137.100 39.330 137.250 ;
        RECT 30.130 136.650 30.730 137.100 ;
        RECT 38.730 136.650 39.330 137.100 ;
        RECT 30.130 136.500 34.080 136.650 ;
        RECT 35.380 136.500 39.330 136.650 ;
        RECT 30.130 136.050 30.730 136.500 ;
        RECT 38.730 136.050 39.330 136.500 ;
        RECT 30.130 135.900 34.080 136.050 ;
        RECT 35.380 135.900 39.330 136.050 ;
        RECT 30.130 135.450 30.730 135.900 ;
        RECT 38.730 135.450 39.330 135.900 ;
        RECT 30.130 135.300 34.080 135.450 ;
        RECT 35.380 135.300 39.330 135.450 ;
        RECT 30.130 134.850 30.730 135.300 ;
        RECT 38.730 134.850 39.330 135.300 ;
        RECT 30.130 134.700 34.080 134.850 ;
        RECT 35.380 134.700 39.330 134.850 ;
        RECT 30.130 134.250 30.730 134.700 ;
        RECT 38.730 134.250 39.330 134.700 ;
        RECT 30.130 134.100 34.080 134.250 ;
        RECT 35.380 134.100 39.330 134.250 ;
        RECT 30.130 133.650 30.730 134.100 ;
        RECT 38.730 133.650 39.330 134.100 ;
        RECT 30.130 133.500 34.080 133.650 ;
        RECT 35.380 133.500 39.330 133.650 ;
        RECT 30.130 133.050 30.730 133.500 ;
        RECT 38.730 133.050 39.330 133.500 ;
        RECT 30.130 132.900 34.080 133.050 ;
        RECT 35.380 132.900 39.330 133.050 ;
        RECT 30.130 132.450 30.730 132.900 ;
        RECT 38.730 132.450 39.330 132.900 ;
        RECT 30.130 132.300 34.080 132.450 ;
        RECT 35.380 132.300 39.330 132.450 ;
        RECT 30.130 131.850 30.730 132.300 ;
        RECT 38.730 131.850 39.330 132.300 ;
        RECT 30.130 131.700 34.080 131.850 ;
        RECT 35.380 131.700 39.330 131.850 ;
        RECT 30.130 131.250 30.730 131.700 ;
        RECT 38.730 131.250 39.330 131.700 ;
        RECT 30.130 131.100 34.080 131.250 ;
        RECT 35.380 131.100 39.330 131.250 ;
        RECT 30.130 130.650 30.730 131.100 ;
        RECT 38.730 130.650 39.330 131.100 ;
        RECT 30.130 130.450 34.080 130.650 ;
        RECT 35.380 130.450 39.330 130.650 ;
        RECT 39.780 130.450 39.930 138.000 ;
        RECT 40.380 130.450 40.530 138.000 ;
        RECT 40.980 130.450 41.130 138.000 ;
        RECT 41.580 130.450 41.730 138.000 ;
        RECT 42.180 130.450 42.330 138.000 ;
        RECT 42.780 135.150 42.930 138.000 ;
        RECT 43.530 135.600 45.930 138.800 ;
        RECT 49.280 138.650 50.730 138.950 ;
        RECT 46.530 138.450 50.730 138.650 ;
        RECT 58.730 138.950 70.730 139.800 ;
        RECT 58.730 138.900 69.130 138.950 ;
        RECT 58.730 138.650 60.180 138.900 ;
        RECT 60.330 138.800 69.130 138.900 ;
        RECT 58.730 138.450 62.930 138.650 ;
        RECT 46.530 138.300 54.080 138.450 ;
        RECT 55.430 138.300 62.930 138.450 ;
        RECT 46.530 138.000 50.730 138.300 ;
        RECT 46.530 135.150 46.680 138.000 ;
        RECT 47.130 130.450 47.280 138.000 ;
        RECT 47.730 130.450 47.880 138.000 ;
        RECT 48.330 130.450 48.480 138.000 ;
        RECT 48.930 130.450 49.080 138.000 ;
        RECT 49.530 130.450 49.680 138.000 ;
        RECT 50.130 137.850 50.730 138.000 ;
        RECT 58.730 138.000 62.930 138.300 ;
        RECT 58.730 137.850 59.330 138.000 ;
        RECT 50.130 137.700 54.080 137.850 ;
        RECT 55.380 137.700 59.330 137.850 ;
        RECT 50.130 137.250 50.730 137.700 ;
        RECT 58.730 137.250 59.330 137.700 ;
        RECT 50.130 137.100 54.080 137.250 ;
        RECT 55.380 137.100 59.330 137.250 ;
        RECT 50.130 136.650 50.730 137.100 ;
        RECT 58.730 136.650 59.330 137.100 ;
        RECT 50.130 136.500 54.080 136.650 ;
        RECT 55.380 136.500 59.330 136.650 ;
        RECT 50.130 136.050 50.730 136.500 ;
        RECT 58.730 136.050 59.330 136.500 ;
        RECT 50.130 135.900 54.080 136.050 ;
        RECT 55.380 135.900 59.330 136.050 ;
        RECT 50.130 135.450 50.730 135.900 ;
        RECT 58.730 135.450 59.330 135.900 ;
        RECT 50.130 135.300 54.080 135.450 ;
        RECT 55.380 135.300 59.330 135.450 ;
        RECT 50.130 134.850 50.730 135.300 ;
        RECT 58.730 134.850 59.330 135.300 ;
        RECT 50.130 134.700 54.080 134.850 ;
        RECT 55.380 134.700 59.330 134.850 ;
        RECT 50.130 134.250 50.730 134.700 ;
        RECT 58.730 134.250 59.330 134.700 ;
        RECT 50.130 134.100 54.080 134.250 ;
        RECT 55.380 134.100 59.330 134.250 ;
        RECT 50.130 133.650 50.730 134.100 ;
        RECT 58.730 133.650 59.330 134.100 ;
        RECT 50.130 133.500 54.080 133.650 ;
        RECT 55.380 133.500 59.330 133.650 ;
        RECT 50.130 133.050 50.730 133.500 ;
        RECT 58.730 133.050 59.330 133.500 ;
        RECT 50.130 132.900 54.080 133.050 ;
        RECT 55.380 132.900 59.330 133.050 ;
        RECT 50.130 132.450 50.730 132.900 ;
        RECT 58.730 132.450 59.330 132.900 ;
        RECT 50.130 132.300 54.080 132.450 ;
        RECT 55.380 132.300 59.330 132.450 ;
        RECT 50.130 131.850 50.730 132.300 ;
        RECT 58.730 131.850 59.330 132.300 ;
        RECT 50.130 131.700 54.080 131.850 ;
        RECT 55.380 131.700 59.330 131.850 ;
        RECT 50.130 131.250 50.730 131.700 ;
        RECT 58.730 131.250 59.330 131.700 ;
        RECT 50.130 131.100 54.080 131.250 ;
        RECT 55.380 131.100 59.330 131.250 ;
        RECT 50.130 130.650 50.730 131.100 ;
        RECT 58.730 130.650 59.330 131.100 ;
        RECT 50.130 130.450 54.080 130.650 ;
        RECT 55.380 130.450 59.330 130.650 ;
        RECT 59.780 130.450 59.930 138.000 ;
        RECT 60.380 130.450 60.530 138.000 ;
        RECT 60.980 130.450 61.130 138.000 ;
        RECT 61.580 130.450 61.730 138.000 ;
        RECT 62.180 130.450 62.330 138.000 ;
        RECT 62.780 135.150 62.930 138.000 ;
        RECT 63.530 135.600 65.930 138.800 ;
        RECT 69.280 138.650 70.730 138.950 ;
        RECT 66.530 138.450 70.730 138.650 ;
        RECT 78.730 138.950 90.730 139.800 ;
        RECT 78.730 138.900 89.130 138.950 ;
        RECT 78.730 138.650 80.180 138.900 ;
        RECT 80.330 138.800 89.130 138.900 ;
        RECT 78.730 138.450 82.930 138.650 ;
        RECT 66.530 138.300 74.080 138.450 ;
        RECT 75.430 138.300 82.930 138.450 ;
        RECT 66.530 138.000 70.730 138.300 ;
        RECT 66.530 135.150 66.680 138.000 ;
        RECT 67.130 130.450 67.280 138.000 ;
        RECT 67.730 130.450 67.880 138.000 ;
        RECT 68.330 130.450 68.480 138.000 ;
        RECT 68.930 130.450 69.080 138.000 ;
        RECT 69.530 130.450 69.680 138.000 ;
        RECT 70.130 137.850 70.730 138.000 ;
        RECT 78.730 138.000 82.930 138.300 ;
        RECT 78.730 137.850 79.330 138.000 ;
        RECT 70.130 137.700 74.080 137.850 ;
        RECT 75.380 137.700 79.330 137.850 ;
        RECT 70.130 137.250 70.730 137.700 ;
        RECT 78.730 137.250 79.330 137.700 ;
        RECT 70.130 137.100 74.080 137.250 ;
        RECT 75.380 137.100 79.330 137.250 ;
        RECT 70.130 136.650 70.730 137.100 ;
        RECT 78.730 136.650 79.330 137.100 ;
        RECT 70.130 136.500 74.080 136.650 ;
        RECT 75.380 136.500 79.330 136.650 ;
        RECT 70.130 136.050 70.730 136.500 ;
        RECT 78.730 136.050 79.330 136.500 ;
        RECT 70.130 135.900 74.080 136.050 ;
        RECT 75.380 135.900 79.330 136.050 ;
        RECT 70.130 135.450 70.730 135.900 ;
        RECT 78.730 135.450 79.330 135.900 ;
        RECT 70.130 135.300 74.080 135.450 ;
        RECT 75.380 135.300 79.330 135.450 ;
        RECT 70.130 134.850 70.730 135.300 ;
        RECT 78.730 134.850 79.330 135.300 ;
        RECT 70.130 134.700 74.080 134.850 ;
        RECT 75.380 134.700 79.330 134.850 ;
        RECT 70.130 134.250 70.730 134.700 ;
        RECT 78.730 134.250 79.330 134.700 ;
        RECT 70.130 134.100 74.080 134.250 ;
        RECT 75.380 134.100 79.330 134.250 ;
        RECT 70.130 133.650 70.730 134.100 ;
        RECT 78.730 133.650 79.330 134.100 ;
        RECT 70.130 133.500 74.080 133.650 ;
        RECT 75.380 133.500 79.330 133.650 ;
        RECT 70.130 133.050 70.730 133.500 ;
        RECT 78.730 133.050 79.330 133.500 ;
        RECT 70.130 132.900 74.080 133.050 ;
        RECT 75.380 132.900 79.330 133.050 ;
        RECT 70.130 132.450 70.730 132.900 ;
        RECT 78.730 132.450 79.330 132.900 ;
        RECT 70.130 132.300 74.080 132.450 ;
        RECT 75.380 132.300 79.330 132.450 ;
        RECT 70.130 131.850 70.730 132.300 ;
        RECT 78.730 131.850 79.330 132.300 ;
        RECT 70.130 131.700 74.080 131.850 ;
        RECT 75.380 131.700 79.330 131.850 ;
        RECT 70.130 131.250 70.730 131.700 ;
        RECT 78.730 131.250 79.330 131.700 ;
        RECT 70.130 131.100 74.080 131.250 ;
        RECT 75.380 131.100 79.330 131.250 ;
        RECT 70.130 130.650 70.730 131.100 ;
        RECT 78.730 130.650 79.330 131.100 ;
        RECT 70.130 130.450 74.080 130.650 ;
        RECT 75.380 130.450 79.330 130.650 ;
        RECT 79.780 130.450 79.930 138.000 ;
        RECT 80.380 130.450 80.530 138.000 ;
        RECT 80.980 130.450 81.130 138.000 ;
        RECT 81.580 130.450 81.730 138.000 ;
        RECT 82.180 130.450 82.330 138.000 ;
        RECT 82.780 135.150 82.930 138.000 ;
        RECT 83.530 135.600 85.930 138.800 ;
        RECT 89.280 138.650 90.730 138.950 ;
        RECT 86.530 138.450 90.730 138.650 ;
        RECT 98.730 138.900 104.730 139.800 ;
        RECT 98.730 138.650 100.180 138.900 ;
        RECT 100.330 138.800 104.730 138.900 ;
        RECT 98.730 138.450 102.930 138.650 ;
        RECT 86.530 138.300 94.080 138.450 ;
        RECT 95.430 138.300 102.930 138.450 ;
        RECT 86.530 138.000 90.730 138.300 ;
        RECT 86.530 135.150 86.680 138.000 ;
        RECT 87.130 130.450 87.280 138.000 ;
        RECT 87.730 130.450 87.880 138.000 ;
        RECT 88.330 130.450 88.480 138.000 ;
        RECT 88.930 130.450 89.080 138.000 ;
        RECT 89.530 130.450 89.680 138.000 ;
        RECT 90.130 137.850 90.730 138.000 ;
        RECT 98.730 138.000 102.930 138.300 ;
        RECT 98.730 137.850 99.330 138.000 ;
        RECT 90.130 137.700 94.080 137.850 ;
        RECT 95.380 137.700 99.330 137.850 ;
        RECT 90.130 137.250 90.730 137.700 ;
        RECT 98.730 137.250 99.330 137.700 ;
        RECT 90.130 137.100 94.080 137.250 ;
        RECT 95.380 137.100 99.330 137.250 ;
        RECT 90.130 136.650 90.730 137.100 ;
        RECT 98.730 136.650 99.330 137.100 ;
        RECT 90.130 136.500 94.080 136.650 ;
        RECT 95.380 136.500 99.330 136.650 ;
        RECT 90.130 136.050 90.730 136.500 ;
        RECT 98.730 136.050 99.330 136.500 ;
        RECT 90.130 135.900 94.080 136.050 ;
        RECT 95.380 135.900 99.330 136.050 ;
        RECT 90.130 135.450 90.730 135.900 ;
        RECT 98.730 135.450 99.330 135.900 ;
        RECT 90.130 135.300 94.080 135.450 ;
        RECT 95.380 135.300 99.330 135.450 ;
        RECT 90.130 134.850 90.730 135.300 ;
        RECT 98.730 134.850 99.330 135.300 ;
        RECT 90.130 134.700 94.080 134.850 ;
        RECT 95.380 134.700 99.330 134.850 ;
        RECT 90.130 134.250 90.730 134.700 ;
        RECT 98.730 134.250 99.330 134.700 ;
        RECT 90.130 134.100 94.080 134.250 ;
        RECT 95.380 134.100 99.330 134.250 ;
        RECT 90.130 133.650 90.730 134.100 ;
        RECT 98.730 133.650 99.330 134.100 ;
        RECT 90.130 133.500 94.080 133.650 ;
        RECT 95.380 133.500 99.330 133.650 ;
        RECT 90.130 133.050 90.730 133.500 ;
        RECT 98.730 133.050 99.330 133.500 ;
        RECT 90.130 132.900 94.080 133.050 ;
        RECT 95.380 132.900 99.330 133.050 ;
        RECT 90.130 132.450 90.730 132.900 ;
        RECT 98.730 132.450 99.330 132.900 ;
        RECT 90.130 132.300 94.080 132.450 ;
        RECT 95.380 132.300 99.330 132.450 ;
        RECT 90.130 131.850 90.730 132.300 ;
        RECT 98.730 131.850 99.330 132.300 ;
        RECT 90.130 131.700 94.080 131.850 ;
        RECT 95.380 131.700 99.330 131.850 ;
        RECT 90.130 131.250 90.730 131.700 ;
        RECT 98.730 131.250 99.330 131.700 ;
        RECT 90.130 131.100 94.080 131.250 ;
        RECT 95.380 131.100 99.330 131.250 ;
        RECT 90.130 130.650 90.730 131.100 ;
        RECT 98.730 130.650 99.330 131.100 ;
        RECT 90.130 130.450 94.080 130.650 ;
        RECT 95.380 130.450 99.330 130.650 ;
        RECT 99.780 130.450 99.930 138.000 ;
        RECT 100.380 130.450 100.530 138.000 ;
        RECT 100.980 130.450 101.130 138.000 ;
        RECT 101.580 130.450 101.730 138.000 ;
        RECT 102.180 130.450 102.330 138.000 ;
        RECT 102.780 135.150 102.930 138.000 ;
        RECT 103.530 137.335 104.730 138.800 ;
        RECT 103.530 136.060 107.135 137.335 ;
        RECT 103.530 135.600 104.730 136.060 ;
        RECT 2.315 124.450 4.315 126.745 ;
        RECT 4.730 123.255 5.930 124.400 ;
        RECT 2.315 121.980 5.930 123.255 ;
        RECT 4.730 121.200 5.930 121.980 ;
        RECT 6.530 122.000 6.680 124.900 ;
        RECT 7.130 122.000 7.280 129.550 ;
        RECT 7.730 122.000 7.880 129.550 ;
        RECT 8.330 122.000 8.480 129.550 ;
        RECT 8.930 122.000 9.080 129.550 ;
        RECT 9.530 122.000 9.680 129.550 ;
        RECT 10.130 129.350 14.080 129.550 ;
        RECT 15.380 129.350 19.330 129.550 ;
        RECT 10.130 128.900 10.730 129.350 ;
        RECT 18.730 128.900 19.330 129.350 ;
        RECT 10.130 128.750 14.080 128.900 ;
        RECT 15.380 128.750 19.330 128.900 ;
        RECT 10.130 128.300 10.730 128.750 ;
        RECT 18.730 128.300 19.330 128.750 ;
        RECT 10.130 128.150 14.080 128.300 ;
        RECT 15.380 128.150 19.330 128.300 ;
        RECT 10.130 127.700 10.730 128.150 ;
        RECT 18.730 127.700 19.330 128.150 ;
        RECT 10.130 127.550 14.080 127.700 ;
        RECT 15.380 127.550 19.330 127.700 ;
        RECT 10.130 127.100 10.730 127.550 ;
        RECT 18.730 127.100 19.330 127.550 ;
        RECT 10.130 126.950 14.080 127.100 ;
        RECT 15.380 126.950 19.330 127.100 ;
        RECT 10.130 126.500 10.730 126.950 ;
        RECT 18.730 126.500 19.330 126.950 ;
        RECT 10.130 126.350 14.080 126.500 ;
        RECT 15.380 126.350 19.330 126.500 ;
        RECT 10.130 125.900 10.730 126.350 ;
        RECT 18.730 125.900 19.330 126.350 ;
        RECT 10.130 125.750 14.080 125.900 ;
        RECT 15.380 125.750 19.330 125.900 ;
        RECT 10.130 125.300 10.730 125.750 ;
        RECT 18.730 125.300 19.330 125.750 ;
        RECT 10.130 125.150 14.080 125.300 ;
        RECT 15.380 125.150 19.330 125.300 ;
        RECT 10.130 124.700 10.730 125.150 ;
        RECT 18.730 124.700 19.330 125.150 ;
        RECT 10.130 124.550 14.080 124.700 ;
        RECT 15.380 124.550 19.330 124.700 ;
        RECT 10.130 124.100 10.730 124.550 ;
        RECT 18.730 124.100 19.330 124.550 ;
        RECT 10.130 123.950 14.080 124.100 ;
        RECT 15.380 123.950 19.330 124.100 ;
        RECT 10.130 123.500 10.730 123.950 ;
        RECT 18.730 123.500 19.330 123.950 ;
        RECT 10.130 123.350 14.080 123.500 ;
        RECT 15.380 123.350 19.330 123.500 ;
        RECT 10.130 122.900 10.730 123.350 ;
        RECT 18.730 122.900 19.330 123.350 ;
        RECT 10.130 122.750 14.080 122.900 ;
        RECT 15.380 122.750 19.330 122.900 ;
        RECT 10.130 122.300 10.730 122.750 ;
        RECT 18.730 122.300 19.330 122.750 ;
        RECT 10.130 122.150 14.080 122.300 ;
        RECT 15.380 122.150 19.330 122.300 ;
        RECT 10.130 122.000 10.730 122.150 ;
        RECT 6.530 121.700 10.730 122.000 ;
        RECT 18.730 122.000 19.330 122.150 ;
        RECT 19.780 122.000 19.930 129.550 ;
        RECT 20.380 122.000 20.530 129.550 ;
        RECT 20.980 122.000 21.130 129.550 ;
        RECT 21.580 122.000 21.730 129.550 ;
        RECT 22.180 122.000 22.330 129.550 ;
        RECT 22.780 122.000 22.930 124.900 ;
        RECT 18.730 121.700 22.930 122.000 ;
        RECT 6.530 121.550 14.080 121.700 ;
        RECT 15.380 121.550 22.930 121.700 ;
        RECT 6.530 121.350 10.730 121.550 ;
        RECT 4.730 121.050 9.130 121.200 ;
        RECT 9.280 121.050 10.730 121.350 ;
        RECT 4.730 120.150 10.730 121.050 ;
        RECT 18.730 121.350 22.930 121.550 ;
        RECT 18.730 121.050 20.180 121.350 ;
        RECT 23.530 121.200 25.930 124.400 ;
        RECT 26.530 122.000 26.680 124.900 ;
        RECT 27.130 122.000 27.280 129.550 ;
        RECT 27.730 122.000 27.880 129.550 ;
        RECT 28.330 122.000 28.480 129.550 ;
        RECT 28.930 122.000 29.080 129.550 ;
        RECT 29.530 122.000 29.680 129.550 ;
        RECT 30.130 129.350 34.080 129.550 ;
        RECT 35.380 129.350 39.330 129.550 ;
        RECT 30.130 128.900 30.730 129.350 ;
        RECT 38.730 128.900 39.330 129.350 ;
        RECT 30.130 128.750 34.080 128.900 ;
        RECT 35.380 128.750 39.330 128.900 ;
        RECT 30.130 128.300 30.730 128.750 ;
        RECT 38.730 128.300 39.330 128.750 ;
        RECT 30.130 128.150 34.080 128.300 ;
        RECT 35.380 128.150 39.330 128.300 ;
        RECT 30.130 127.700 30.730 128.150 ;
        RECT 38.730 127.700 39.330 128.150 ;
        RECT 30.130 127.550 34.080 127.700 ;
        RECT 35.380 127.550 39.330 127.700 ;
        RECT 30.130 127.100 30.730 127.550 ;
        RECT 38.730 127.100 39.330 127.550 ;
        RECT 30.130 126.950 34.080 127.100 ;
        RECT 35.380 126.950 39.330 127.100 ;
        RECT 30.130 126.500 30.730 126.950 ;
        RECT 38.730 126.500 39.330 126.950 ;
        RECT 30.130 126.350 34.080 126.500 ;
        RECT 35.380 126.350 39.330 126.500 ;
        RECT 30.130 125.900 30.730 126.350 ;
        RECT 38.730 125.900 39.330 126.350 ;
        RECT 30.130 125.750 34.080 125.900 ;
        RECT 35.380 125.750 39.330 125.900 ;
        RECT 30.130 125.300 30.730 125.750 ;
        RECT 38.730 125.300 39.330 125.750 ;
        RECT 30.130 125.150 34.080 125.300 ;
        RECT 35.380 125.150 39.330 125.300 ;
        RECT 30.130 124.700 30.730 125.150 ;
        RECT 38.730 124.700 39.330 125.150 ;
        RECT 30.130 124.550 34.080 124.700 ;
        RECT 35.380 124.550 39.330 124.700 ;
        RECT 30.130 124.100 30.730 124.550 ;
        RECT 38.730 124.100 39.330 124.550 ;
        RECT 30.130 123.950 34.080 124.100 ;
        RECT 35.380 123.950 39.330 124.100 ;
        RECT 30.130 123.500 30.730 123.950 ;
        RECT 38.730 123.500 39.330 123.950 ;
        RECT 30.130 123.350 34.080 123.500 ;
        RECT 35.380 123.350 39.330 123.500 ;
        RECT 30.130 122.900 30.730 123.350 ;
        RECT 38.730 122.900 39.330 123.350 ;
        RECT 30.130 122.750 34.080 122.900 ;
        RECT 35.380 122.750 39.330 122.900 ;
        RECT 30.130 122.300 30.730 122.750 ;
        RECT 38.730 122.300 39.330 122.750 ;
        RECT 30.130 122.150 34.080 122.300 ;
        RECT 35.380 122.150 39.330 122.300 ;
        RECT 30.130 122.000 30.730 122.150 ;
        RECT 26.530 121.700 30.730 122.000 ;
        RECT 38.730 122.000 39.330 122.150 ;
        RECT 39.780 122.000 39.930 129.550 ;
        RECT 40.380 122.000 40.530 129.550 ;
        RECT 40.980 122.000 41.130 129.550 ;
        RECT 41.580 122.000 41.730 129.550 ;
        RECT 42.180 122.000 42.330 129.550 ;
        RECT 42.780 122.000 42.930 124.900 ;
        RECT 38.730 121.700 42.930 122.000 ;
        RECT 26.530 121.550 34.080 121.700 ;
        RECT 35.380 121.550 42.930 121.700 ;
        RECT 26.530 121.350 30.730 121.550 ;
        RECT 20.330 121.050 29.130 121.200 ;
        RECT 29.280 121.050 30.730 121.350 ;
        RECT 18.730 120.150 30.730 121.050 ;
        RECT 38.730 121.350 42.930 121.550 ;
        RECT 38.730 121.050 40.180 121.350 ;
        RECT 43.530 121.200 45.930 124.400 ;
        RECT 46.530 122.000 46.680 124.900 ;
        RECT 47.130 122.000 47.280 129.550 ;
        RECT 47.730 122.000 47.880 129.550 ;
        RECT 48.330 122.000 48.480 129.550 ;
        RECT 48.930 122.000 49.080 129.550 ;
        RECT 49.530 122.000 49.680 129.550 ;
        RECT 50.130 129.350 54.080 129.550 ;
        RECT 55.380 129.350 59.330 129.550 ;
        RECT 50.130 128.900 50.730 129.350 ;
        RECT 58.730 128.900 59.330 129.350 ;
        RECT 50.130 128.750 54.080 128.900 ;
        RECT 55.380 128.750 59.330 128.900 ;
        RECT 50.130 128.300 50.730 128.750 ;
        RECT 58.730 128.300 59.330 128.750 ;
        RECT 50.130 128.150 54.080 128.300 ;
        RECT 55.380 128.150 59.330 128.300 ;
        RECT 50.130 127.700 50.730 128.150 ;
        RECT 58.730 127.700 59.330 128.150 ;
        RECT 50.130 127.550 54.080 127.700 ;
        RECT 55.380 127.550 59.330 127.700 ;
        RECT 50.130 127.100 50.730 127.550 ;
        RECT 58.730 127.100 59.330 127.550 ;
        RECT 50.130 126.950 54.080 127.100 ;
        RECT 55.380 126.950 59.330 127.100 ;
        RECT 50.130 126.500 50.730 126.950 ;
        RECT 58.730 126.500 59.330 126.950 ;
        RECT 50.130 126.350 54.080 126.500 ;
        RECT 55.380 126.350 59.330 126.500 ;
        RECT 50.130 125.900 50.730 126.350 ;
        RECT 58.730 125.900 59.330 126.350 ;
        RECT 50.130 125.750 54.080 125.900 ;
        RECT 55.380 125.750 59.330 125.900 ;
        RECT 50.130 125.300 50.730 125.750 ;
        RECT 58.730 125.300 59.330 125.750 ;
        RECT 50.130 125.150 54.080 125.300 ;
        RECT 55.380 125.150 59.330 125.300 ;
        RECT 50.130 124.700 50.730 125.150 ;
        RECT 58.730 124.700 59.330 125.150 ;
        RECT 50.130 124.550 54.080 124.700 ;
        RECT 55.380 124.550 59.330 124.700 ;
        RECT 50.130 124.100 50.730 124.550 ;
        RECT 58.730 124.100 59.330 124.550 ;
        RECT 50.130 123.950 54.080 124.100 ;
        RECT 55.380 123.950 59.330 124.100 ;
        RECT 50.130 123.500 50.730 123.950 ;
        RECT 58.730 123.500 59.330 123.950 ;
        RECT 50.130 123.350 54.080 123.500 ;
        RECT 55.380 123.350 59.330 123.500 ;
        RECT 50.130 122.900 50.730 123.350 ;
        RECT 58.730 122.900 59.330 123.350 ;
        RECT 50.130 122.750 54.080 122.900 ;
        RECT 55.380 122.750 59.330 122.900 ;
        RECT 50.130 122.300 50.730 122.750 ;
        RECT 58.730 122.300 59.330 122.750 ;
        RECT 50.130 122.150 54.080 122.300 ;
        RECT 55.380 122.150 59.330 122.300 ;
        RECT 50.130 122.000 50.730 122.150 ;
        RECT 46.530 121.700 50.730 122.000 ;
        RECT 58.730 122.000 59.330 122.150 ;
        RECT 59.780 122.000 59.930 129.550 ;
        RECT 60.380 122.000 60.530 129.550 ;
        RECT 60.980 122.000 61.130 129.550 ;
        RECT 61.580 122.000 61.730 129.550 ;
        RECT 62.180 122.000 62.330 129.550 ;
        RECT 62.780 122.000 62.930 124.900 ;
        RECT 58.730 121.700 62.930 122.000 ;
        RECT 46.530 121.550 54.080 121.700 ;
        RECT 55.380 121.550 62.930 121.700 ;
        RECT 46.530 121.350 50.730 121.550 ;
        RECT 40.330 121.050 49.130 121.200 ;
        RECT 49.280 121.050 50.730 121.350 ;
        RECT 38.730 120.150 50.730 121.050 ;
        RECT 58.730 121.350 62.930 121.550 ;
        RECT 58.730 121.050 60.180 121.350 ;
        RECT 63.530 121.200 65.930 124.400 ;
        RECT 66.530 122.000 66.680 124.900 ;
        RECT 67.130 122.000 67.280 129.550 ;
        RECT 67.730 122.000 67.880 129.550 ;
        RECT 68.330 122.000 68.480 129.550 ;
        RECT 68.930 122.000 69.080 129.550 ;
        RECT 69.530 122.000 69.680 129.550 ;
        RECT 70.130 129.350 74.080 129.550 ;
        RECT 75.380 129.350 79.330 129.550 ;
        RECT 70.130 128.900 70.730 129.350 ;
        RECT 78.730 128.900 79.330 129.350 ;
        RECT 70.130 128.750 74.080 128.900 ;
        RECT 75.380 128.750 79.330 128.900 ;
        RECT 70.130 128.300 70.730 128.750 ;
        RECT 78.730 128.300 79.330 128.750 ;
        RECT 70.130 128.150 74.080 128.300 ;
        RECT 75.380 128.150 79.330 128.300 ;
        RECT 70.130 127.700 70.730 128.150 ;
        RECT 78.730 127.700 79.330 128.150 ;
        RECT 70.130 127.550 74.080 127.700 ;
        RECT 75.380 127.550 79.330 127.700 ;
        RECT 70.130 127.100 70.730 127.550 ;
        RECT 78.730 127.100 79.330 127.550 ;
        RECT 70.130 126.950 74.080 127.100 ;
        RECT 75.380 126.950 79.330 127.100 ;
        RECT 70.130 126.500 70.730 126.950 ;
        RECT 78.730 126.500 79.330 126.950 ;
        RECT 70.130 126.350 74.080 126.500 ;
        RECT 75.380 126.350 79.330 126.500 ;
        RECT 70.130 125.900 70.730 126.350 ;
        RECT 78.730 125.900 79.330 126.350 ;
        RECT 70.130 125.750 74.080 125.900 ;
        RECT 75.380 125.750 79.330 125.900 ;
        RECT 70.130 125.300 70.730 125.750 ;
        RECT 78.730 125.300 79.330 125.750 ;
        RECT 70.130 125.150 74.080 125.300 ;
        RECT 75.380 125.150 79.330 125.300 ;
        RECT 70.130 124.700 70.730 125.150 ;
        RECT 78.730 124.700 79.330 125.150 ;
        RECT 70.130 124.550 74.080 124.700 ;
        RECT 75.380 124.550 79.330 124.700 ;
        RECT 70.130 124.100 70.730 124.550 ;
        RECT 78.730 124.100 79.330 124.550 ;
        RECT 70.130 123.950 74.080 124.100 ;
        RECT 75.380 123.950 79.330 124.100 ;
        RECT 70.130 123.500 70.730 123.950 ;
        RECT 78.730 123.500 79.330 123.950 ;
        RECT 70.130 123.350 74.080 123.500 ;
        RECT 75.380 123.350 79.330 123.500 ;
        RECT 70.130 122.900 70.730 123.350 ;
        RECT 78.730 122.900 79.330 123.350 ;
        RECT 70.130 122.750 74.080 122.900 ;
        RECT 75.380 122.750 79.330 122.900 ;
        RECT 70.130 122.300 70.730 122.750 ;
        RECT 78.730 122.300 79.330 122.750 ;
        RECT 70.130 122.150 74.080 122.300 ;
        RECT 75.380 122.150 79.330 122.300 ;
        RECT 70.130 122.000 70.730 122.150 ;
        RECT 66.530 121.700 70.730 122.000 ;
        RECT 78.730 122.000 79.330 122.150 ;
        RECT 79.780 122.000 79.930 129.550 ;
        RECT 80.380 122.000 80.530 129.550 ;
        RECT 80.980 122.000 81.130 129.550 ;
        RECT 81.580 122.000 81.730 129.550 ;
        RECT 82.180 122.000 82.330 129.550 ;
        RECT 82.780 122.000 82.930 124.900 ;
        RECT 78.730 121.700 82.930 122.000 ;
        RECT 66.530 121.550 74.080 121.700 ;
        RECT 75.380 121.550 82.930 121.700 ;
        RECT 66.530 121.350 70.730 121.550 ;
        RECT 60.330 121.050 69.130 121.200 ;
        RECT 69.280 121.050 70.730 121.350 ;
        RECT 58.730 120.150 70.730 121.050 ;
        RECT 78.730 121.350 82.930 121.550 ;
        RECT 78.730 121.050 80.180 121.350 ;
        RECT 83.530 121.200 85.930 124.400 ;
        RECT 86.530 122.000 86.680 124.900 ;
        RECT 87.130 122.000 87.280 129.550 ;
        RECT 87.730 122.000 87.880 129.550 ;
        RECT 88.330 122.000 88.480 129.550 ;
        RECT 88.930 122.000 89.080 129.550 ;
        RECT 89.530 122.000 89.680 129.550 ;
        RECT 90.130 129.350 94.080 129.550 ;
        RECT 95.380 129.350 99.330 129.550 ;
        RECT 90.130 128.900 90.730 129.350 ;
        RECT 98.730 128.900 99.330 129.350 ;
        RECT 90.130 128.750 94.080 128.900 ;
        RECT 95.380 128.750 99.330 128.900 ;
        RECT 90.130 128.300 90.730 128.750 ;
        RECT 98.730 128.300 99.330 128.750 ;
        RECT 90.130 128.150 94.080 128.300 ;
        RECT 95.380 128.150 99.330 128.300 ;
        RECT 90.130 127.700 90.730 128.150 ;
        RECT 98.730 127.700 99.330 128.150 ;
        RECT 90.130 127.550 94.080 127.700 ;
        RECT 95.380 127.550 99.330 127.700 ;
        RECT 90.130 127.100 90.730 127.550 ;
        RECT 98.730 127.100 99.330 127.550 ;
        RECT 90.130 126.950 94.080 127.100 ;
        RECT 95.380 126.950 99.330 127.100 ;
        RECT 90.130 126.500 90.730 126.950 ;
        RECT 98.730 126.500 99.330 126.950 ;
        RECT 90.130 126.350 94.080 126.500 ;
        RECT 95.380 126.350 99.330 126.500 ;
        RECT 90.130 125.900 90.730 126.350 ;
        RECT 98.730 125.900 99.330 126.350 ;
        RECT 90.130 125.750 94.080 125.900 ;
        RECT 95.380 125.750 99.330 125.900 ;
        RECT 90.130 125.300 90.730 125.750 ;
        RECT 98.730 125.300 99.330 125.750 ;
        RECT 90.130 125.150 94.080 125.300 ;
        RECT 95.380 125.150 99.330 125.300 ;
        RECT 90.130 124.700 90.730 125.150 ;
        RECT 98.730 124.700 99.330 125.150 ;
        RECT 90.130 124.550 94.080 124.700 ;
        RECT 95.380 124.550 99.330 124.700 ;
        RECT 90.130 124.100 90.730 124.550 ;
        RECT 98.730 124.100 99.330 124.550 ;
        RECT 90.130 123.950 94.080 124.100 ;
        RECT 95.380 123.950 99.330 124.100 ;
        RECT 90.130 123.500 90.730 123.950 ;
        RECT 98.730 123.500 99.330 123.950 ;
        RECT 90.130 123.350 94.080 123.500 ;
        RECT 95.380 123.350 99.330 123.500 ;
        RECT 90.130 122.900 90.730 123.350 ;
        RECT 98.730 122.900 99.330 123.350 ;
        RECT 90.130 122.750 94.080 122.900 ;
        RECT 95.380 122.750 99.330 122.900 ;
        RECT 90.130 122.300 90.730 122.750 ;
        RECT 98.730 122.300 99.330 122.750 ;
        RECT 90.130 122.150 94.080 122.300 ;
        RECT 95.380 122.150 99.330 122.300 ;
        RECT 90.130 122.000 90.730 122.150 ;
        RECT 86.530 121.700 90.730 122.000 ;
        RECT 98.730 122.000 99.330 122.150 ;
        RECT 99.780 122.000 99.930 129.550 ;
        RECT 100.380 122.000 100.530 129.550 ;
        RECT 100.980 122.000 101.130 129.550 ;
        RECT 101.580 122.000 101.730 129.550 ;
        RECT 102.180 122.000 102.330 129.550 ;
        RECT 102.780 122.000 102.930 124.900 ;
        RECT 98.730 121.700 102.930 122.000 ;
        RECT 86.530 121.550 94.080 121.700 ;
        RECT 95.380 121.550 102.930 121.700 ;
        RECT 86.530 121.350 90.730 121.550 ;
        RECT 80.330 121.050 89.130 121.200 ;
        RECT 89.280 121.050 90.730 121.350 ;
        RECT 78.730 120.150 90.730 121.050 ;
        RECT 98.730 121.350 102.930 121.550 ;
        RECT 103.530 123.120 104.730 124.400 ;
        RECT 103.530 121.845 107.140 123.120 ;
        RECT 98.730 121.050 100.180 121.350 ;
        RECT 103.530 121.200 104.730 121.845 ;
        RECT 100.330 121.050 104.730 121.200 ;
        RECT 98.730 120.150 104.730 121.050 ;
        RECT 4.730 119.850 9.130 120.150 ;
        RECT 20.330 119.850 29.130 120.150 ;
        RECT 40.330 119.850 49.130 120.150 ;
        RECT 60.330 119.850 69.130 120.150 ;
        RECT 80.330 119.850 89.130 120.150 ;
        RECT 4.730 118.950 10.730 119.850 ;
        RECT 20.330 119.800 30.730 119.850 ;
        RECT 40.330 119.800 50.730 119.850 ;
        RECT 60.330 119.800 70.730 119.850 ;
        RECT 80.330 119.800 90.730 119.850 ;
        RECT 100.330 119.800 104.730 120.150 ;
        RECT 4.730 118.800 9.130 118.950 ;
        RECT 4.730 117.845 5.930 118.800 ;
        RECT 9.280 118.650 10.730 118.950 ;
        RECT 2.315 116.570 5.930 117.845 ;
        RECT 4.730 115.600 5.930 116.570 ;
        RECT 6.530 118.450 10.730 118.650 ;
        RECT 18.730 118.950 30.730 119.800 ;
        RECT 18.730 118.900 29.130 118.950 ;
        RECT 18.730 118.650 20.180 118.900 ;
        RECT 20.330 118.800 29.130 118.900 ;
        RECT 18.730 118.450 22.930 118.650 ;
        RECT 6.530 118.300 14.080 118.450 ;
        RECT 15.430 118.300 22.930 118.450 ;
        RECT 6.530 118.000 10.730 118.300 ;
        RECT 2.315 113.250 4.315 115.545 ;
        RECT 6.530 115.150 6.680 118.000 ;
        RECT 7.130 110.450 7.280 118.000 ;
        RECT 7.730 110.450 7.880 118.000 ;
        RECT 8.330 110.450 8.480 118.000 ;
        RECT 8.930 110.450 9.080 118.000 ;
        RECT 9.530 110.450 9.680 118.000 ;
        RECT 10.130 117.850 10.730 118.000 ;
        RECT 18.730 118.000 22.930 118.300 ;
        RECT 18.730 117.850 19.330 118.000 ;
        RECT 10.130 117.700 14.080 117.850 ;
        RECT 15.380 117.700 19.330 117.850 ;
        RECT 10.130 117.250 10.730 117.700 ;
        RECT 18.730 117.250 19.330 117.700 ;
        RECT 10.130 117.100 14.080 117.250 ;
        RECT 15.380 117.100 19.330 117.250 ;
        RECT 10.130 116.650 10.730 117.100 ;
        RECT 18.730 116.650 19.330 117.100 ;
        RECT 10.130 116.500 14.080 116.650 ;
        RECT 15.380 116.500 19.330 116.650 ;
        RECT 10.130 116.050 10.730 116.500 ;
        RECT 18.730 116.050 19.330 116.500 ;
        RECT 10.130 115.900 14.080 116.050 ;
        RECT 15.380 115.900 19.330 116.050 ;
        RECT 10.130 115.450 10.730 115.900 ;
        RECT 18.730 115.450 19.330 115.900 ;
        RECT 10.130 115.300 14.080 115.450 ;
        RECT 15.380 115.300 19.330 115.450 ;
        RECT 10.130 114.850 10.730 115.300 ;
        RECT 18.730 114.850 19.330 115.300 ;
        RECT 10.130 114.700 14.080 114.850 ;
        RECT 15.380 114.700 19.330 114.850 ;
        RECT 10.130 114.250 10.730 114.700 ;
        RECT 18.730 114.250 19.330 114.700 ;
        RECT 10.130 114.100 14.080 114.250 ;
        RECT 15.380 114.100 19.330 114.250 ;
        RECT 10.130 113.650 10.730 114.100 ;
        RECT 18.730 113.650 19.330 114.100 ;
        RECT 10.130 113.500 14.080 113.650 ;
        RECT 15.380 113.500 19.330 113.650 ;
        RECT 10.130 113.050 10.730 113.500 ;
        RECT 18.730 113.050 19.330 113.500 ;
        RECT 10.130 112.900 14.080 113.050 ;
        RECT 15.380 112.900 19.330 113.050 ;
        RECT 10.130 112.450 10.730 112.900 ;
        RECT 18.730 112.450 19.330 112.900 ;
        RECT 10.130 112.300 14.080 112.450 ;
        RECT 15.380 112.300 19.330 112.450 ;
        RECT 10.130 111.850 10.730 112.300 ;
        RECT 18.730 111.850 19.330 112.300 ;
        RECT 10.130 111.700 14.080 111.850 ;
        RECT 15.380 111.700 19.330 111.850 ;
        RECT 10.130 111.250 10.730 111.700 ;
        RECT 18.730 111.250 19.330 111.700 ;
        RECT 10.130 111.100 14.080 111.250 ;
        RECT 15.380 111.100 19.330 111.250 ;
        RECT 10.130 110.650 10.730 111.100 ;
        RECT 18.730 110.650 19.330 111.100 ;
        RECT 10.130 110.450 14.080 110.650 ;
        RECT 15.380 110.450 19.330 110.650 ;
        RECT 19.780 110.450 19.930 118.000 ;
        RECT 20.380 110.450 20.530 118.000 ;
        RECT 20.980 110.450 21.130 118.000 ;
        RECT 21.580 110.450 21.730 118.000 ;
        RECT 22.180 110.450 22.330 118.000 ;
        RECT 22.780 115.150 22.930 118.000 ;
        RECT 23.530 115.600 25.930 118.800 ;
        RECT 29.280 118.650 30.730 118.950 ;
        RECT 26.530 118.450 30.730 118.650 ;
        RECT 38.730 118.950 50.730 119.800 ;
        RECT 38.730 118.900 49.130 118.950 ;
        RECT 38.730 118.650 40.180 118.900 ;
        RECT 40.330 118.800 49.130 118.900 ;
        RECT 38.730 118.450 42.930 118.650 ;
        RECT 26.530 118.300 34.080 118.450 ;
        RECT 35.430 118.300 42.930 118.450 ;
        RECT 26.530 118.000 30.730 118.300 ;
        RECT 26.530 115.150 26.680 118.000 ;
        RECT 27.130 110.450 27.280 118.000 ;
        RECT 27.730 110.450 27.880 118.000 ;
        RECT 28.330 110.450 28.480 118.000 ;
        RECT 28.930 110.450 29.080 118.000 ;
        RECT 29.530 110.450 29.680 118.000 ;
        RECT 30.130 117.850 30.730 118.000 ;
        RECT 38.730 118.000 42.930 118.300 ;
        RECT 38.730 117.850 39.330 118.000 ;
        RECT 30.130 117.700 34.080 117.850 ;
        RECT 35.380 117.700 39.330 117.850 ;
        RECT 30.130 117.250 30.730 117.700 ;
        RECT 38.730 117.250 39.330 117.700 ;
        RECT 30.130 117.100 34.080 117.250 ;
        RECT 35.380 117.100 39.330 117.250 ;
        RECT 30.130 116.650 30.730 117.100 ;
        RECT 38.730 116.650 39.330 117.100 ;
        RECT 30.130 116.500 34.080 116.650 ;
        RECT 35.380 116.500 39.330 116.650 ;
        RECT 30.130 116.050 30.730 116.500 ;
        RECT 38.730 116.050 39.330 116.500 ;
        RECT 30.130 115.900 34.080 116.050 ;
        RECT 35.380 115.900 39.330 116.050 ;
        RECT 30.130 115.450 30.730 115.900 ;
        RECT 38.730 115.450 39.330 115.900 ;
        RECT 30.130 115.300 34.080 115.450 ;
        RECT 35.380 115.300 39.330 115.450 ;
        RECT 30.130 114.850 30.730 115.300 ;
        RECT 38.730 114.850 39.330 115.300 ;
        RECT 30.130 114.700 34.080 114.850 ;
        RECT 35.380 114.700 39.330 114.850 ;
        RECT 30.130 114.250 30.730 114.700 ;
        RECT 38.730 114.250 39.330 114.700 ;
        RECT 30.130 114.100 34.080 114.250 ;
        RECT 35.380 114.100 39.330 114.250 ;
        RECT 30.130 113.650 30.730 114.100 ;
        RECT 38.730 113.650 39.330 114.100 ;
        RECT 30.130 113.500 34.080 113.650 ;
        RECT 35.380 113.500 39.330 113.650 ;
        RECT 30.130 113.050 30.730 113.500 ;
        RECT 38.730 113.050 39.330 113.500 ;
        RECT 30.130 112.900 34.080 113.050 ;
        RECT 35.380 112.900 39.330 113.050 ;
        RECT 30.130 112.450 30.730 112.900 ;
        RECT 38.730 112.450 39.330 112.900 ;
        RECT 30.130 112.300 34.080 112.450 ;
        RECT 35.380 112.300 39.330 112.450 ;
        RECT 30.130 111.850 30.730 112.300 ;
        RECT 38.730 111.850 39.330 112.300 ;
        RECT 30.130 111.700 34.080 111.850 ;
        RECT 35.380 111.700 39.330 111.850 ;
        RECT 30.130 111.250 30.730 111.700 ;
        RECT 38.730 111.250 39.330 111.700 ;
        RECT 30.130 111.100 34.080 111.250 ;
        RECT 35.380 111.100 39.330 111.250 ;
        RECT 30.130 110.650 30.730 111.100 ;
        RECT 38.730 110.650 39.330 111.100 ;
        RECT 30.130 110.450 34.080 110.650 ;
        RECT 35.380 110.450 39.330 110.650 ;
        RECT 39.780 110.450 39.930 118.000 ;
        RECT 40.380 110.450 40.530 118.000 ;
        RECT 40.980 110.450 41.130 118.000 ;
        RECT 41.580 110.450 41.730 118.000 ;
        RECT 42.180 110.450 42.330 118.000 ;
        RECT 42.780 115.150 42.930 118.000 ;
        RECT 43.530 115.600 45.930 118.800 ;
        RECT 49.280 118.650 50.730 118.950 ;
        RECT 46.530 118.450 50.730 118.650 ;
        RECT 58.730 118.950 70.730 119.800 ;
        RECT 58.730 118.900 69.130 118.950 ;
        RECT 58.730 118.650 60.180 118.900 ;
        RECT 60.330 118.800 69.130 118.900 ;
        RECT 58.730 118.450 62.930 118.650 ;
        RECT 46.530 118.300 54.080 118.450 ;
        RECT 55.430 118.300 62.930 118.450 ;
        RECT 46.530 118.000 50.730 118.300 ;
        RECT 46.530 115.150 46.680 118.000 ;
        RECT 47.130 110.450 47.280 118.000 ;
        RECT 47.730 110.450 47.880 118.000 ;
        RECT 48.330 110.450 48.480 118.000 ;
        RECT 48.930 110.450 49.080 118.000 ;
        RECT 49.530 110.450 49.680 118.000 ;
        RECT 50.130 117.850 50.730 118.000 ;
        RECT 58.730 118.000 62.930 118.300 ;
        RECT 58.730 117.850 59.330 118.000 ;
        RECT 50.130 117.700 54.080 117.850 ;
        RECT 55.380 117.700 59.330 117.850 ;
        RECT 50.130 117.250 50.730 117.700 ;
        RECT 58.730 117.250 59.330 117.700 ;
        RECT 50.130 117.100 54.080 117.250 ;
        RECT 55.380 117.100 59.330 117.250 ;
        RECT 50.130 116.650 50.730 117.100 ;
        RECT 58.730 116.650 59.330 117.100 ;
        RECT 50.130 116.500 54.080 116.650 ;
        RECT 55.380 116.500 59.330 116.650 ;
        RECT 50.130 116.050 50.730 116.500 ;
        RECT 58.730 116.050 59.330 116.500 ;
        RECT 50.130 115.900 54.080 116.050 ;
        RECT 55.380 115.900 59.330 116.050 ;
        RECT 50.130 115.450 50.730 115.900 ;
        RECT 58.730 115.450 59.330 115.900 ;
        RECT 50.130 115.300 54.080 115.450 ;
        RECT 55.380 115.300 59.330 115.450 ;
        RECT 50.130 114.850 50.730 115.300 ;
        RECT 58.730 114.850 59.330 115.300 ;
        RECT 50.130 114.700 54.080 114.850 ;
        RECT 55.380 114.700 59.330 114.850 ;
        RECT 50.130 114.250 50.730 114.700 ;
        RECT 58.730 114.250 59.330 114.700 ;
        RECT 50.130 114.100 54.080 114.250 ;
        RECT 55.380 114.100 59.330 114.250 ;
        RECT 50.130 113.650 50.730 114.100 ;
        RECT 58.730 113.650 59.330 114.100 ;
        RECT 50.130 113.500 54.080 113.650 ;
        RECT 55.380 113.500 59.330 113.650 ;
        RECT 50.130 113.050 50.730 113.500 ;
        RECT 58.730 113.050 59.330 113.500 ;
        RECT 50.130 112.900 54.080 113.050 ;
        RECT 55.380 112.900 59.330 113.050 ;
        RECT 50.130 112.450 50.730 112.900 ;
        RECT 58.730 112.450 59.330 112.900 ;
        RECT 50.130 112.300 54.080 112.450 ;
        RECT 55.380 112.300 59.330 112.450 ;
        RECT 50.130 111.850 50.730 112.300 ;
        RECT 58.730 111.850 59.330 112.300 ;
        RECT 50.130 111.700 54.080 111.850 ;
        RECT 55.380 111.700 59.330 111.850 ;
        RECT 50.130 111.250 50.730 111.700 ;
        RECT 58.730 111.250 59.330 111.700 ;
        RECT 50.130 111.100 54.080 111.250 ;
        RECT 55.380 111.100 59.330 111.250 ;
        RECT 50.130 110.650 50.730 111.100 ;
        RECT 58.730 110.650 59.330 111.100 ;
        RECT 50.130 110.450 54.080 110.650 ;
        RECT 55.380 110.450 59.330 110.650 ;
        RECT 59.780 110.450 59.930 118.000 ;
        RECT 60.380 110.450 60.530 118.000 ;
        RECT 60.980 110.450 61.130 118.000 ;
        RECT 61.580 110.450 61.730 118.000 ;
        RECT 62.180 110.450 62.330 118.000 ;
        RECT 62.780 115.150 62.930 118.000 ;
        RECT 63.530 115.600 65.930 118.800 ;
        RECT 69.280 118.650 70.730 118.950 ;
        RECT 66.530 118.450 70.730 118.650 ;
        RECT 78.730 118.950 90.730 119.800 ;
        RECT 78.730 118.900 89.130 118.950 ;
        RECT 78.730 118.650 80.180 118.900 ;
        RECT 80.330 118.800 89.130 118.900 ;
        RECT 78.730 118.450 82.930 118.650 ;
        RECT 66.530 118.300 74.080 118.450 ;
        RECT 75.430 118.300 82.930 118.450 ;
        RECT 66.530 118.000 70.730 118.300 ;
        RECT 66.530 115.150 66.680 118.000 ;
        RECT 67.130 110.450 67.280 118.000 ;
        RECT 67.730 110.450 67.880 118.000 ;
        RECT 68.330 110.450 68.480 118.000 ;
        RECT 68.930 110.450 69.080 118.000 ;
        RECT 69.530 110.450 69.680 118.000 ;
        RECT 70.130 117.850 70.730 118.000 ;
        RECT 78.730 118.000 82.930 118.300 ;
        RECT 78.730 117.850 79.330 118.000 ;
        RECT 70.130 117.700 74.080 117.850 ;
        RECT 75.380 117.700 79.330 117.850 ;
        RECT 70.130 117.250 70.730 117.700 ;
        RECT 78.730 117.250 79.330 117.700 ;
        RECT 70.130 117.100 74.080 117.250 ;
        RECT 75.380 117.100 79.330 117.250 ;
        RECT 70.130 116.650 70.730 117.100 ;
        RECT 78.730 116.650 79.330 117.100 ;
        RECT 70.130 116.500 74.080 116.650 ;
        RECT 75.380 116.500 79.330 116.650 ;
        RECT 70.130 116.050 70.730 116.500 ;
        RECT 78.730 116.050 79.330 116.500 ;
        RECT 70.130 115.900 74.080 116.050 ;
        RECT 75.380 115.900 79.330 116.050 ;
        RECT 70.130 115.450 70.730 115.900 ;
        RECT 78.730 115.450 79.330 115.900 ;
        RECT 70.130 115.300 74.080 115.450 ;
        RECT 75.380 115.300 79.330 115.450 ;
        RECT 70.130 114.850 70.730 115.300 ;
        RECT 78.730 114.850 79.330 115.300 ;
        RECT 70.130 114.700 74.080 114.850 ;
        RECT 75.380 114.700 79.330 114.850 ;
        RECT 70.130 114.250 70.730 114.700 ;
        RECT 78.730 114.250 79.330 114.700 ;
        RECT 70.130 114.100 74.080 114.250 ;
        RECT 75.380 114.100 79.330 114.250 ;
        RECT 70.130 113.650 70.730 114.100 ;
        RECT 78.730 113.650 79.330 114.100 ;
        RECT 70.130 113.500 74.080 113.650 ;
        RECT 75.380 113.500 79.330 113.650 ;
        RECT 70.130 113.050 70.730 113.500 ;
        RECT 78.730 113.050 79.330 113.500 ;
        RECT 70.130 112.900 74.080 113.050 ;
        RECT 75.380 112.900 79.330 113.050 ;
        RECT 70.130 112.450 70.730 112.900 ;
        RECT 78.730 112.450 79.330 112.900 ;
        RECT 70.130 112.300 74.080 112.450 ;
        RECT 75.380 112.300 79.330 112.450 ;
        RECT 70.130 111.850 70.730 112.300 ;
        RECT 78.730 111.850 79.330 112.300 ;
        RECT 70.130 111.700 74.080 111.850 ;
        RECT 75.380 111.700 79.330 111.850 ;
        RECT 70.130 111.250 70.730 111.700 ;
        RECT 78.730 111.250 79.330 111.700 ;
        RECT 70.130 111.100 74.080 111.250 ;
        RECT 75.380 111.100 79.330 111.250 ;
        RECT 70.130 110.650 70.730 111.100 ;
        RECT 78.730 110.650 79.330 111.100 ;
        RECT 70.130 110.450 74.080 110.650 ;
        RECT 75.380 110.450 79.330 110.650 ;
        RECT 79.780 110.450 79.930 118.000 ;
        RECT 80.380 110.450 80.530 118.000 ;
        RECT 80.980 110.450 81.130 118.000 ;
        RECT 81.580 110.450 81.730 118.000 ;
        RECT 82.180 110.450 82.330 118.000 ;
        RECT 82.780 115.150 82.930 118.000 ;
        RECT 83.530 115.600 85.930 118.800 ;
        RECT 89.280 118.650 90.730 118.950 ;
        RECT 86.530 118.450 90.730 118.650 ;
        RECT 98.730 118.900 104.730 119.800 ;
        RECT 98.730 118.650 100.180 118.900 ;
        RECT 100.330 118.800 104.730 118.900 ;
        RECT 98.730 118.450 102.930 118.650 ;
        RECT 86.530 118.300 94.080 118.450 ;
        RECT 95.430 118.300 102.930 118.450 ;
        RECT 86.530 118.000 90.730 118.300 ;
        RECT 86.530 115.150 86.680 118.000 ;
        RECT 87.130 110.450 87.280 118.000 ;
        RECT 87.730 110.450 87.880 118.000 ;
        RECT 88.330 110.450 88.480 118.000 ;
        RECT 88.930 110.450 89.080 118.000 ;
        RECT 89.530 110.450 89.680 118.000 ;
        RECT 90.130 117.850 90.730 118.000 ;
        RECT 98.730 118.000 102.930 118.300 ;
        RECT 98.730 117.850 99.330 118.000 ;
        RECT 90.130 117.700 94.080 117.850 ;
        RECT 95.380 117.700 99.330 117.850 ;
        RECT 90.130 117.250 90.730 117.700 ;
        RECT 98.730 117.250 99.330 117.700 ;
        RECT 90.130 117.100 94.080 117.250 ;
        RECT 95.380 117.100 99.330 117.250 ;
        RECT 90.130 116.650 90.730 117.100 ;
        RECT 98.730 116.650 99.330 117.100 ;
        RECT 90.130 116.500 94.080 116.650 ;
        RECT 95.380 116.500 99.330 116.650 ;
        RECT 90.130 116.050 90.730 116.500 ;
        RECT 98.730 116.050 99.330 116.500 ;
        RECT 90.130 115.900 94.080 116.050 ;
        RECT 95.380 115.900 99.330 116.050 ;
        RECT 90.130 115.450 90.730 115.900 ;
        RECT 98.730 115.450 99.330 115.900 ;
        RECT 90.130 115.300 94.080 115.450 ;
        RECT 95.380 115.300 99.330 115.450 ;
        RECT 90.130 114.850 90.730 115.300 ;
        RECT 98.730 114.850 99.330 115.300 ;
        RECT 90.130 114.700 94.080 114.850 ;
        RECT 95.380 114.700 99.330 114.850 ;
        RECT 90.130 114.250 90.730 114.700 ;
        RECT 98.730 114.250 99.330 114.700 ;
        RECT 90.130 114.100 94.080 114.250 ;
        RECT 95.380 114.100 99.330 114.250 ;
        RECT 90.130 113.650 90.730 114.100 ;
        RECT 98.730 113.650 99.330 114.100 ;
        RECT 90.130 113.500 94.080 113.650 ;
        RECT 95.380 113.500 99.330 113.650 ;
        RECT 90.130 113.050 90.730 113.500 ;
        RECT 98.730 113.050 99.330 113.500 ;
        RECT 90.130 112.900 94.080 113.050 ;
        RECT 95.380 112.900 99.330 113.050 ;
        RECT 90.130 112.450 90.730 112.900 ;
        RECT 98.730 112.450 99.330 112.900 ;
        RECT 90.130 112.300 94.080 112.450 ;
        RECT 95.380 112.300 99.330 112.450 ;
        RECT 90.130 111.850 90.730 112.300 ;
        RECT 98.730 111.850 99.330 112.300 ;
        RECT 90.130 111.700 94.080 111.850 ;
        RECT 95.380 111.700 99.330 111.850 ;
        RECT 90.130 111.250 90.730 111.700 ;
        RECT 98.730 111.250 99.330 111.700 ;
        RECT 90.130 111.100 94.080 111.250 ;
        RECT 95.380 111.100 99.330 111.250 ;
        RECT 90.130 110.650 90.730 111.100 ;
        RECT 98.730 110.650 99.330 111.100 ;
        RECT 90.130 110.450 94.080 110.650 ;
        RECT 95.380 110.450 99.330 110.650 ;
        RECT 99.780 110.450 99.930 118.000 ;
        RECT 100.380 110.450 100.530 118.000 ;
        RECT 100.980 110.450 101.130 118.000 ;
        RECT 101.580 110.450 101.730 118.000 ;
        RECT 102.180 110.450 102.330 118.000 ;
        RECT 102.780 115.150 102.930 118.000 ;
        RECT 103.530 117.245 104.730 118.800 ;
        RECT 103.530 115.970 107.140 117.245 ;
        RECT 103.530 115.600 104.730 115.970 ;
        RECT 2.315 104.455 4.315 106.750 ;
        RECT 4.730 103.470 5.930 104.400 ;
        RECT 2.315 102.195 5.930 103.470 ;
        RECT 4.730 101.200 5.930 102.195 ;
        RECT 6.530 102.000 6.680 104.900 ;
        RECT 7.130 102.000 7.280 109.550 ;
        RECT 7.730 102.000 7.880 109.550 ;
        RECT 8.330 102.000 8.480 109.550 ;
        RECT 8.930 102.000 9.080 109.550 ;
        RECT 9.530 102.000 9.680 109.550 ;
        RECT 10.130 109.350 14.080 109.550 ;
        RECT 15.380 109.350 19.330 109.550 ;
        RECT 10.130 108.900 10.730 109.350 ;
        RECT 18.730 108.900 19.330 109.350 ;
        RECT 10.130 108.750 14.080 108.900 ;
        RECT 15.380 108.750 19.330 108.900 ;
        RECT 10.130 108.300 10.730 108.750 ;
        RECT 18.730 108.300 19.330 108.750 ;
        RECT 10.130 108.150 14.080 108.300 ;
        RECT 15.380 108.150 19.330 108.300 ;
        RECT 10.130 107.700 10.730 108.150 ;
        RECT 18.730 107.700 19.330 108.150 ;
        RECT 10.130 107.550 14.080 107.700 ;
        RECT 15.380 107.550 19.330 107.700 ;
        RECT 10.130 107.100 10.730 107.550 ;
        RECT 18.730 107.100 19.330 107.550 ;
        RECT 10.130 106.950 14.080 107.100 ;
        RECT 15.380 106.950 19.330 107.100 ;
        RECT 10.130 106.500 10.730 106.950 ;
        RECT 18.730 106.500 19.330 106.950 ;
        RECT 10.130 106.350 14.080 106.500 ;
        RECT 15.380 106.350 19.330 106.500 ;
        RECT 10.130 105.900 10.730 106.350 ;
        RECT 18.730 105.900 19.330 106.350 ;
        RECT 10.130 105.750 14.080 105.900 ;
        RECT 15.380 105.750 19.330 105.900 ;
        RECT 10.130 105.300 10.730 105.750 ;
        RECT 18.730 105.300 19.330 105.750 ;
        RECT 10.130 105.150 14.080 105.300 ;
        RECT 15.380 105.150 19.330 105.300 ;
        RECT 10.130 104.700 10.730 105.150 ;
        RECT 18.730 104.700 19.330 105.150 ;
        RECT 10.130 104.550 14.080 104.700 ;
        RECT 15.380 104.550 19.330 104.700 ;
        RECT 10.130 104.100 10.730 104.550 ;
        RECT 18.730 104.100 19.330 104.550 ;
        RECT 10.130 103.950 14.080 104.100 ;
        RECT 15.380 103.950 19.330 104.100 ;
        RECT 10.130 103.500 10.730 103.950 ;
        RECT 18.730 103.500 19.330 103.950 ;
        RECT 10.130 103.350 14.080 103.500 ;
        RECT 15.380 103.350 19.330 103.500 ;
        RECT 10.130 102.900 10.730 103.350 ;
        RECT 18.730 102.900 19.330 103.350 ;
        RECT 10.130 102.750 14.080 102.900 ;
        RECT 15.380 102.750 19.330 102.900 ;
        RECT 10.130 102.300 10.730 102.750 ;
        RECT 18.730 102.300 19.330 102.750 ;
        RECT 10.130 102.150 14.080 102.300 ;
        RECT 15.380 102.150 19.330 102.300 ;
        RECT 10.130 102.000 10.730 102.150 ;
        RECT 6.530 101.700 10.730 102.000 ;
        RECT 18.730 102.000 19.330 102.150 ;
        RECT 19.780 102.000 19.930 109.550 ;
        RECT 20.380 102.000 20.530 109.550 ;
        RECT 20.980 102.000 21.130 109.550 ;
        RECT 21.580 102.000 21.730 109.550 ;
        RECT 22.180 102.000 22.330 109.550 ;
        RECT 22.780 102.000 22.930 104.900 ;
        RECT 18.730 101.700 22.930 102.000 ;
        RECT 6.530 101.550 14.080 101.700 ;
        RECT 15.380 101.550 22.930 101.700 ;
        RECT 6.530 101.350 10.730 101.550 ;
        RECT 4.730 101.050 9.130 101.200 ;
        RECT 9.280 101.050 10.730 101.350 ;
        RECT 4.730 100.150 10.730 101.050 ;
        RECT 18.730 101.350 22.930 101.550 ;
        RECT 18.730 101.050 20.180 101.350 ;
        RECT 23.530 101.200 25.930 104.400 ;
        RECT 26.530 102.000 26.680 104.900 ;
        RECT 27.130 102.000 27.280 109.550 ;
        RECT 27.730 102.000 27.880 109.550 ;
        RECT 28.330 102.000 28.480 109.550 ;
        RECT 28.930 102.000 29.080 109.550 ;
        RECT 29.530 102.000 29.680 109.550 ;
        RECT 30.130 109.350 34.080 109.550 ;
        RECT 35.380 109.350 39.330 109.550 ;
        RECT 30.130 108.900 30.730 109.350 ;
        RECT 38.730 108.900 39.330 109.350 ;
        RECT 30.130 108.750 34.080 108.900 ;
        RECT 35.380 108.750 39.330 108.900 ;
        RECT 30.130 108.300 30.730 108.750 ;
        RECT 38.730 108.300 39.330 108.750 ;
        RECT 30.130 108.150 34.080 108.300 ;
        RECT 35.380 108.150 39.330 108.300 ;
        RECT 30.130 107.700 30.730 108.150 ;
        RECT 38.730 107.700 39.330 108.150 ;
        RECT 30.130 107.550 34.080 107.700 ;
        RECT 35.380 107.550 39.330 107.700 ;
        RECT 30.130 107.100 30.730 107.550 ;
        RECT 38.730 107.100 39.330 107.550 ;
        RECT 30.130 106.950 34.080 107.100 ;
        RECT 35.380 106.950 39.330 107.100 ;
        RECT 30.130 106.500 30.730 106.950 ;
        RECT 38.730 106.500 39.330 106.950 ;
        RECT 30.130 106.350 34.080 106.500 ;
        RECT 35.380 106.350 39.330 106.500 ;
        RECT 30.130 105.900 30.730 106.350 ;
        RECT 38.730 105.900 39.330 106.350 ;
        RECT 30.130 105.750 34.080 105.900 ;
        RECT 35.380 105.750 39.330 105.900 ;
        RECT 30.130 105.300 30.730 105.750 ;
        RECT 38.730 105.300 39.330 105.750 ;
        RECT 30.130 105.150 34.080 105.300 ;
        RECT 35.380 105.150 39.330 105.300 ;
        RECT 30.130 104.700 30.730 105.150 ;
        RECT 38.730 104.700 39.330 105.150 ;
        RECT 30.130 104.550 34.080 104.700 ;
        RECT 35.380 104.550 39.330 104.700 ;
        RECT 30.130 104.100 30.730 104.550 ;
        RECT 38.730 104.100 39.330 104.550 ;
        RECT 30.130 103.950 34.080 104.100 ;
        RECT 35.380 103.950 39.330 104.100 ;
        RECT 30.130 103.500 30.730 103.950 ;
        RECT 38.730 103.500 39.330 103.950 ;
        RECT 30.130 103.350 34.080 103.500 ;
        RECT 35.380 103.350 39.330 103.500 ;
        RECT 30.130 102.900 30.730 103.350 ;
        RECT 38.730 102.900 39.330 103.350 ;
        RECT 30.130 102.750 34.080 102.900 ;
        RECT 35.380 102.750 39.330 102.900 ;
        RECT 30.130 102.300 30.730 102.750 ;
        RECT 38.730 102.300 39.330 102.750 ;
        RECT 30.130 102.150 34.080 102.300 ;
        RECT 35.380 102.150 39.330 102.300 ;
        RECT 30.130 102.000 30.730 102.150 ;
        RECT 26.530 101.700 30.730 102.000 ;
        RECT 38.730 102.000 39.330 102.150 ;
        RECT 39.780 102.000 39.930 109.550 ;
        RECT 40.380 102.000 40.530 109.550 ;
        RECT 40.980 102.000 41.130 109.550 ;
        RECT 41.580 102.000 41.730 109.550 ;
        RECT 42.180 102.000 42.330 109.550 ;
        RECT 42.780 102.000 42.930 104.900 ;
        RECT 38.730 101.700 42.930 102.000 ;
        RECT 26.530 101.550 34.080 101.700 ;
        RECT 35.380 101.550 42.930 101.700 ;
        RECT 26.530 101.350 30.730 101.550 ;
        RECT 20.330 101.050 29.130 101.200 ;
        RECT 29.280 101.050 30.730 101.350 ;
        RECT 18.730 100.150 30.730 101.050 ;
        RECT 38.730 101.350 42.930 101.550 ;
        RECT 38.730 101.050 40.180 101.350 ;
        RECT 43.530 101.200 45.930 104.400 ;
        RECT 46.530 102.000 46.680 104.900 ;
        RECT 47.130 102.000 47.280 109.550 ;
        RECT 47.730 102.000 47.880 109.550 ;
        RECT 48.330 102.000 48.480 109.550 ;
        RECT 48.930 102.000 49.080 109.550 ;
        RECT 49.530 102.000 49.680 109.550 ;
        RECT 50.130 109.350 54.080 109.550 ;
        RECT 55.380 109.350 59.330 109.550 ;
        RECT 50.130 108.900 50.730 109.350 ;
        RECT 58.730 108.900 59.330 109.350 ;
        RECT 50.130 108.750 54.080 108.900 ;
        RECT 55.380 108.750 59.330 108.900 ;
        RECT 50.130 108.300 50.730 108.750 ;
        RECT 58.730 108.300 59.330 108.750 ;
        RECT 50.130 108.150 54.080 108.300 ;
        RECT 55.380 108.150 59.330 108.300 ;
        RECT 50.130 107.700 50.730 108.150 ;
        RECT 58.730 107.700 59.330 108.150 ;
        RECT 50.130 107.550 54.080 107.700 ;
        RECT 55.380 107.550 59.330 107.700 ;
        RECT 50.130 107.100 50.730 107.550 ;
        RECT 58.730 107.100 59.330 107.550 ;
        RECT 50.130 106.950 54.080 107.100 ;
        RECT 55.380 106.950 59.330 107.100 ;
        RECT 50.130 106.500 50.730 106.950 ;
        RECT 58.730 106.500 59.330 106.950 ;
        RECT 50.130 106.350 54.080 106.500 ;
        RECT 55.380 106.350 59.330 106.500 ;
        RECT 50.130 105.900 50.730 106.350 ;
        RECT 58.730 105.900 59.330 106.350 ;
        RECT 50.130 105.750 54.080 105.900 ;
        RECT 55.380 105.750 59.330 105.900 ;
        RECT 50.130 105.300 50.730 105.750 ;
        RECT 58.730 105.300 59.330 105.750 ;
        RECT 50.130 105.150 54.080 105.300 ;
        RECT 55.380 105.150 59.330 105.300 ;
        RECT 50.130 104.700 50.730 105.150 ;
        RECT 58.730 104.700 59.330 105.150 ;
        RECT 50.130 104.550 54.080 104.700 ;
        RECT 55.380 104.550 59.330 104.700 ;
        RECT 50.130 104.100 50.730 104.550 ;
        RECT 58.730 104.100 59.330 104.550 ;
        RECT 50.130 103.950 54.080 104.100 ;
        RECT 55.380 103.950 59.330 104.100 ;
        RECT 50.130 103.500 50.730 103.950 ;
        RECT 58.730 103.500 59.330 103.950 ;
        RECT 50.130 103.350 54.080 103.500 ;
        RECT 55.380 103.350 59.330 103.500 ;
        RECT 50.130 102.900 50.730 103.350 ;
        RECT 58.730 102.900 59.330 103.350 ;
        RECT 50.130 102.750 54.080 102.900 ;
        RECT 55.380 102.750 59.330 102.900 ;
        RECT 50.130 102.300 50.730 102.750 ;
        RECT 58.730 102.300 59.330 102.750 ;
        RECT 50.130 102.150 54.080 102.300 ;
        RECT 55.380 102.150 59.330 102.300 ;
        RECT 50.130 102.000 50.730 102.150 ;
        RECT 46.530 101.700 50.730 102.000 ;
        RECT 58.730 102.000 59.330 102.150 ;
        RECT 59.780 102.000 59.930 109.550 ;
        RECT 60.380 102.000 60.530 109.550 ;
        RECT 60.980 102.000 61.130 109.550 ;
        RECT 61.580 102.000 61.730 109.550 ;
        RECT 62.180 102.000 62.330 109.550 ;
        RECT 62.780 102.000 62.930 104.900 ;
        RECT 58.730 101.700 62.930 102.000 ;
        RECT 46.530 101.550 54.080 101.700 ;
        RECT 55.380 101.550 62.930 101.700 ;
        RECT 46.530 101.350 50.730 101.550 ;
        RECT 40.330 101.050 49.130 101.200 ;
        RECT 49.280 101.050 50.730 101.350 ;
        RECT 38.730 100.150 50.730 101.050 ;
        RECT 58.730 101.350 62.930 101.550 ;
        RECT 58.730 101.050 60.180 101.350 ;
        RECT 63.530 101.200 65.930 104.400 ;
        RECT 66.530 102.000 66.680 104.900 ;
        RECT 67.130 102.000 67.280 109.550 ;
        RECT 67.730 102.000 67.880 109.550 ;
        RECT 68.330 102.000 68.480 109.550 ;
        RECT 68.930 102.000 69.080 109.550 ;
        RECT 69.530 102.000 69.680 109.550 ;
        RECT 70.130 109.350 74.080 109.550 ;
        RECT 75.380 109.350 79.330 109.550 ;
        RECT 70.130 108.900 70.730 109.350 ;
        RECT 78.730 108.900 79.330 109.350 ;
        RECT 70.130 108.750 74.080 108.900 ;
        RECT 75.380 108.750 79.330 108.900 ;
        RECT 70.130 108.300 70.730 108.750 ;
        RECT 78.730 108.300 79.330 108.750 ;
        RECT 70.130 108.150 74.080 108.300 ;
        RECT 75.380 108.150 79.330 108.300 ;
        RECT 70.130 107.700 70.730 108.150 ;
        RECT 78.730 107.700 79.330 108.150 ;
        RECT 70.130 107.550 74.080 107.700 ;
        RECT 75.380 107.550 79.330 107.700 ;
        RECT 70.130 107.100 70.730 107.550 ;
        RECT 78.730 107.100 79.330 107.550 ;
        RECT 70.130 106.950 74.080 107.100 ;
        RECT 75.380 106.950 79.330 107.100 ;
        RECT 70.130 106.500 70.730 106.950 ;
        RECT 78.730 106.500 79.330 106.950 ;
        RECT 70.130 106.350 74.080 106.500 ;
        RECT 75.380 106.350 79.330 106.500 ;
        RECT 70.130 105.900 70.730 106.350 ;
        RECT 78.730 105.900 79.330 106.350 ;
        RECT 70.130 105.750 74.080 105.900 ;
        RECT 75.380 105.750 79.330 105.900 ;
        RECT 70.130 105.300 70.730 105.750 ;
        RECT 78.730 105.300 79.330 105.750 ;
        RECT 70.130 105.150 74.080 105.300 ;
        RECT 75.380 105.150 79.330 105.300 ;
        RECT 70.130 104.700 70.730 105.150 ;
        RECT 78.730 104.700 79.330 105.150 ;
        RECT 70.130 104.550 74.080 104.700 ;
        RECT 75.380 104.550 79.330 104.700 ;
        RECT 70.130 104.100 70.730 104.550 ;
        RECT 78.730 104.100 79.330 104.550 ;
        RECT 70.130 103.950 74.080 104.100 ;
        RECT 75.380 103.950 79.330 104.100 ;
        RECT 70.130 103.500 70.730 103.950 ;
        RECT 78.730 103.500 79.330 103.950 ;
        RECT 70.130 103.350 74.080 103.500 ;
        RECT 75.380 103.350 79.330 103.500 ;
        RECT 70.130 102.900 70.730 103.350 ;
        RECT 78.730 102.900 79.330 103.350 ;
        RECT 70.130 102.750 74.080 102.900 ;
        RECT 75.380 102.750 79.330 102.900 ;
        RECT 70.130 102.300 70.730 102.750 ;
        RECT 78.730 102.300 79.330 102.750 ;
        RECT 70.130 102.150 74.080 102.300 ;
        RECT 75.380 102.150 79.330 102.300 ;
        RECT 70.130 102.000 70.730 102.150 ;
        RECT 66.530 101.700 70.730 102.000 ;
        RECT 78.730 102.000 79.330 102.150 ;
        RECT 79.780 102.000 79.930 109.550 ;
        RECT 80.380 102.000 80.530 109.550 ;
        RECT 80.980 102.000 81.130 109.550 ;
        RECT 81.580 102.000 81.730 109.550 ;
        RECT 82.180 102.000 82.330 109.550 ;
        RECT 82.780 102.000 82.930 104.900 ;
        RECT 78.730 101.700 82.930 102.000 ;
        RECT 66.530 101.550 74.080 101.700 ;
        RECT 75.380 101.550 82.930 101.700 ;
        RECT 66.530 101.350 70.730 101.550 ;
        RECT 60.330 101.050 69.130 101.200 ;
        RECT 69.280 101.050 70.730 101.350 ;
        RECT 58.730 100.150 70.730 101.050 ;
        RECT 78.730 101.350 82.930 101.550 ;
        RECT 78.730 101.050 80.180 101.350 ;
        RECT 83.530 101.200 85.930 104.400 ;
        RECT 86.530 102.000 86.680 104.900 ;
        RECT 87.130 102.000 87.280 109.550 ;
        RECT 87.730 102.000 87.880 109.550 ;
        RECT 88.330 102.000 88.480 109.550 ;
        RECT 88.930 102.000 89.080 109.550 ;
        RECT 89.530 102.000 89.680 109.550 ;
        RECT 90.130 109.350 94.080 109.550 ;
        RECT 95.380 109.350 99.330 109.550 ;
        RECT 90.130 108.900 90.730 109.350 ;
        RECT 98.730 108.900 99.330 109.350 ;
        RECT 90.130 108.750 94.080 108.900 ;
        RECT 95.380 108.750 99.330 108.900 ;
        RECT 90.130 108.300 90.730 108.750 ;
        RECT 98.730 108.300 99.330 108.750 ;
        RECT 90.130 108.150 94.080 108.300 ;
        RECT 95.380 108.150 99.330 108.300 ;
        RECT 90.130 107.700 90.730 108.150 ;
        RECT 98.730 107.700 99.330 108.150 ;
        RECT 90.130 107.550 94.080 107.700 ;
        RECT 95.380 107.550 99.330 107.700 ;
        RECT 90.130 107.100 90.730 107.550 ;
        RECT 98.730 107.100 99.330 107.550 ;
        RECT 90.130 106.950 94.080 107.100 ;
        RECT 95.380 106.950 99.330 107.100 ;
        RECT 90.130 106.500 90.730 106.950 ;
        RECT 98.730 106.500 99.330 106.950 ;
        RECT 90.130 106.350 94.080 106.500 ;
        RECT 95.380 106.350 99.330 106.500 ;
        RECT 90.130 105.900 90.730 106.350 ;
        RECT 98.730 105.900 99.330 106.350 ;
        RECT 90.130 105.750 94.080 105.900 ;
        RECT 95.380 105.750 99.330 105.900 ;
        RECT 90.130 105.300 90.730 105.750 ;
        RECT 98.730 105.300 99.330 105.750 ;
        RECT 90.130 105.150 94.080 105.300 ;
        RECT 95.380 105.150 99.330 105.300 ;
        RECT 90.130 104.700 90.730 105.150 ;
        RECT 98.730 104.700 99.330 105.150 ;
        RECT 90.130 104.550 94.080 104.700 ;
        RECT 95.380 104.550 99.330 104.700 ;
        RECT 90.130 104.100 90.730 104.550 ;
        RECT 98.730 104.100 99.330 104.550 ;
        RECT 90.130 103.950 94.080 104.100 ;
        RECT 95.380 103.950 99.330 104.100 ;
        RECT 90.130 103.500 90.730 103.950 ;
        RECT 98.730 103.500 99.330 103.950 ;
        RECT 90.130 103.350 94.080 103.500 ;
        RECT 95.380 103.350 99.330 103.500 ;
        RECT 90.130 102.900 90.730 103.350 ;
        RECT 98.730 102.900 99.330 103.350 ;
        RECT 90.130 102.750 94.080 102.900 ;
        RECT 95.380 102.750 99.330 102.900 ;
        RECT 90.130 102.300 90.730 102.750 ;
        RECT 98.730 102.300 99.330 102.750 ;
        RECT 90.130 102.150 94.080 102.300 ;
        RECT 95.380 102.150 99.330 102.300 ;
        RECT 90.130 102.000 90.730 102.150 ;
        RECT 86.530 101.700 90.730 102.000 ;
        RECT 98.730 102.000 99.330 102.150 ;
        RECT 99.780 102.000 99.930 109.550 ;
        RECT 100.380 102.000 100.530 109.550 ;
        RECT 100.980 102.000 101.130 109.550 ;
        RECT 101.580 102.000 101.730 109.550 ;
        RECT 102.180 102.000 102.330 109.550 ;
        RECT 102.780 102.000 102.930 104.900 ;
        RECT 98.730 101.700 102.930 102.000 ;
        RECT 86.530 101.550 94.080 101.700 ;
        RECT 95.380 101.550 102.930 101.700 ;
        RECT 86.530 101.350 90.730 101.550 ;
        RECT 80.330 101.050 89.130 101.200 ;
        RECT 89.280 101.050 90.730 101.350 ;
        RECT 78.730 100.150 90.730 101.050 ;
        RECT 98.730 101.350 102.930 101.550 ;
        RECT 103.530 103.040 104.730 104.400 ;
        RECT 103.530 101.765 107.135 103.040 ;
        RECT 98.730 101.050 100.180 101.350 ;
        RECT 103.530 101.200 104.730 101.765 ;
        RECT 100.330 101.050 104.730 101.200 ;
        RECT 98.730 100.150 104.730 101.050 ;
        RECT 4.730 99.850 9.130 100.150 ;
        RECT 20.330 99.850 29.130 100.150 ;
        RECT 40.330 99.850 49.130 100.150 ;
        RECT 60.330 99.850 69.130 100.150 ;
        RECT 80.330 99.850 89.130 100.150 ;
        RECT 4.730 98.950 10.730 99.850 ;
        RECT 20.330 99.800 30.730 99.850 ;
        RECT 40.330 99.800 50.730 99.850 ;
        RECT 60.330 99.800 70.730 99.850 ;
        RECT 80.330 99.800 90.730 99.850 ;
        RECT 100.330 99.800 104.730 100.150 ;
        RECT 4.730 98.800 9.130 98.950 ;
        RECT 4.730 97.965 5.930 98.800 ;
        RECT 9.280 98.650 10.730 98.950 ;
        RECT 2.315 96.690 5.930 97.965 ;
        RECT 4.730 95.600 5.930 96.690 ;
        RECT 6.530 98.450 10.730 98.650 ;
        RECT 18.730 98.950 30.730 99.800 ;
        RECT 18.730 98.900 29.130 98.950 ;
        RECT 18.730 98.650 20.180 98.900 ;
        RECT 20.330 98.800 29.130 98.900 ;
        RECT 18.730 98.450 22.930 98.650 ;
        RECT 6.530 98.300 14.080 98.450 ;
        RECT 15.430 98.300 22.930 98.450 ;
        RECT 6.530 98.000 10.730 98.300 ;
        RECT 2.315 93.250 4.315 95.545 ;
        RECT 6.530 95.150 6.680 98.000 ;
        RECT 7.130 90.450 7.280 98.000 ;
        RECT 7.730 90.450 7.880 98.000 ;
        RECT 8.330 90.450 8.480 98.000 ;
        RECT 8.930 90.450 9.080 98.000 ;
        RECT 9.530 90.450 9.680 98.000 ;
        RECT 10.130 97.850 10.730 98.000 ;
        RECT 18.730 98.000 22.930 98.300 ;
        RECT 18.730 97.850 19.330 98.000 ;
        RECT 10.130 97.700 14.080 97.850 ;
        RECT 15.380 97.700 19.330 97.850 ;
        RECT 10.130 97.250 10.730 97.700 ;
        RECT 18.730 97.250 19.330 97.700 ;
        RECT 10.130 97.100 14.080 97.250 ;
        RECT 15.380 97.100 19.330 97.250 ;
        RECT 10.130 96.650 10.730 97.100 ;
        RECT 18.730 96.650 19.330 97.100 ;
        RECT 10.130 96.500 14.080 96.650 ;
        RECT 15.380 96.500 19.330 96.650 ;
        RECT 10.130 96.050 10.730 96.500 ;
        RECT 18.730 96.050 19.330 96.500 ;
        RECT 10.130 95.900 14.080 96.050 ;
        RECT 15.380 95.900 19.330 96.050 ;
        RECT 10.130 95.450 10.730 95.900 ;
        RECT 18.730 95.450 19.330 95.900 ;
        RECT 10.130 95.300 14.080 95.450 ;
        RECT 15.380 95.300 19.330 95.450 ;
        RECT 10.130 94.850 10.730 95.300 ;
        RECT 18.730 94.850 19.330 95.300 ;
        RECT 10.130 94.700 14.080 94.850 ;
        RECT 15.380 94.700 19.330 94.850 ;
        RECT 10.130 94.250 10.730 94.700 ;
        RECT 18.730 94.250 19.330 94.700 ;
        RECT 10.130 94.100 14.080 94.250 ;
        RECT 15.380 94.100 19.330 94.250 ;
        RECT 10.130 93.650 10.730 94.100 ;
        RECT 18.730 93.650 19.330 94.100 ;
        RECT 10.130 93.500 14.080 93.650 ;
        RECT 15.380 93.500 19.330 93.650 ;
        RECT 10.130 93.050 10.730 93.500 ;
        RECT 18.730 93.050 19.330 93.500 ;
        RECT 10.130 92.900 14.080 93.050 ;
        RECT 15.380 92.900 19.330 93.050 ;
        RECT 10.130 92.450 10.730 92.900 ;
        RECT 18.730 92.450 19.330 92.900 ;
        RECT 10.130 92.300 14.080 92.450 ;
        RECT 15.380 92.300 19.330 92.450 ;
        RECT 10.130 91.850 10.730 92.300 ;
        RECT 18.730 91.850 19.330 92.300 ;
        RECT 10.130 91.700 14.080 91.850 ;
        RECT 15.380 91.700 19.330 91.850 ;
        RECT 10.130 91.250 10.730 91.700 ;
        RECT 18.730 91.250 19.330 91.700 ;
        RECT 10.130 91.100 14.080 91.250 ;
        RECT 15.380 91.100 19.330 91.250 ;
        RECT 10.130 90.650 10.730 91.100 ;
        RECT 18.730 90.650 19.330 91.100 ;
        RECT 10.130 90.450 14.080 90.650 ;
        RECT 15.380 90.450 19.330 90.650 ;
        RECT 19.780 90.450 19.930 98.000 ;
        RECT 20.380 90.450 20.530 98.000 ;
        RECT 20.980 90.450 21.130 98.000 ;
        RECT 21.580 90.450 21.730 98.000 ;
        RECT 22.180 90.450 22.330 98.000 ;
        RECT 22.780 95.150 22.930 98.000 ;
        RECT 23.530 95.600 25.930 98.800 ;
        RECT 29.280 98.650 30.730 98.950 ;
        RECT 26.530 98.450 30.730 98.650 ;
        RECT 38.730 98.950 50.730 99.800 ;
        RECT 38.730 98.900 49.130 98.950 ;
        RECT 38.730 98.650 40.180 98.900 ;
        RECT 40.330 98.800 49.130 98.900 ;
        RECT 38.730 98.450 42.930 98.650 ;
        RECT 26.530 98.300 34.080 98.450 ;
        RECT 35.430 98.300 42.930 98.450 ;
        RECT 26.530 98.000 30.730 98.300 ;
        RECT 26.530 95.150 26.680 98.000 ;
        RECT 27.130 90.450 27.280 98.000 ;
        RECT 27.730 90.450 27.880 98.000 ;
        RECT 28.330 90.450 28.480 98.000 ;
        RECT 28.930 90.450 29.080 98.000 ;
        RECT 29.530 90.450 29.680 98.000 ;
        RECT 30.130 97.850 30.730 98.000 ;
        RECT 38.730 98.000 42.930 98.300 ;
        RECT 38.730 97.850 39.330 98.000 ;
        RECT 30.130 97.700 34.080 97.850 ;
        RECT 35.380 97.700 39.330 97.850 ;
        RECT 30.130 97.250 30.730 97.700 ;
        RECT 38.730 97.250 39.330 97.700 ;
        RECT 30.130 97.100 34.080 97.250 ;
        RECT 35.380 97.100 39.330 97.250 ;
        RECT 30.130 96.650 30.730 97.100 ;
        RECT 38.730 96.650 39.330 97.100 ;
        RECT 30.130 96.500 34.080 96.650 ;
        RECT 35.380 96.500 39.330 96.650 ;
        RECT 30.130 96.050 30.730 96.500 ;
        RECT 38.730 96.050 39.330 96.500 ;
        RECT 30.130 95.900 34.080 96.050 ;
        RECT 35.380 95.900 39.330 96.050 ;
        RECT 30.130 95.450 30.730 95.900 ;
        RECT 38.730 95.450 39.330 95.900 ;
        RECT 30.130 95.300 34.080 95.450 ;
        RECT 35.380 95.300 39.330 95.450 ;
        RECT 30.130 94.850 30.730 95.300 ;
        RECT 38.730 94.850 39.330 95.300 ;
        RECT 30.130 94.700 34.080 94.850 ;
        RECT 35.380 94.700 39.330 94.850 ;
        RECT 30.130 94.250 30.730 94.700 ;
        RECT 38.730 94.250 39.330 94.700 ;
        RECT 30.130 94.100 34.080 94.250 ;
        RECT 35.380 94.100 39.330 94.250 ;
        RECT 30.130 93.650 30.730 94.100 ;
        RECT 38.730 93.650 39.330 94.100 ;
        RECT 30.130 93.500 34.080 93.650 ;
        RECT 35.380 93.500 39.330 93.650 ;
        RECT 30.130 93.050 30.730 93.500 ;
        RECT 38.730 93.050 39.330 93.500 ;
        RECT 30.130 92.900 34.080 93.050 ;
        RECT 35.380 92.900 39.330 93.050 ;
        RECT 30.130 92.450 30.730 92.900 ;
        RECT 38.730 92.450 39.330 92.900 ;
        RECT 30.130 92.300 34.080 92.450 ;
        RECT 35.380 92.300 39.330 92.450 ;
        RECT 30.130 91.850 30.730 92.300 ;
        RECT 38.730 91.850 39.330 92.300 ;
        RECT 30.130 91.700 34.080 91.850 ;
        RECT 35.380 91.700 39.330 91.850 ;
        RECT 30.130 91.250 30.730 91.700 ;
        RECT 38.730 91.250 39.330 91.700 ;
        RECT 30.130 91.100 34.080 91.250 ;
        RECT 35.380 91.100 39.330 91.250 ;
        RECT 30.130 90.650 30.730 91.100 ;
        RECT 38.730 90.650 39.330 91.100 ;
        RECT 30.130 90.450 34.080 90.650 ;
        RECT 35.380 90.450 39.330 90.650 ;
        RECT 39.780 90.450 39.930 98.000 ;
        RECT 40.380 90.450 40.530 98.000 ;
        RECT 40.980 90.450 41.130 98.000 ;
        RECT 41.580 90.450 41.730 98.000 ;
        RECT 42.180 90.450 42.330 98.000 ;
        RECT 42.780 95.150 42.930 98.000 ;
        RECT 43.530 95.600 45.930 98.800 ;
        RECT 49.280 98.650 50.730 98.950 ;
        RECT 46.530 98.450 50.730 98.650 ;
        RECT 58.730 98.950 70.730 99.800 ;
        RECT 58.730 98.900 69.130 98.950 ;
        RECT 58.730 98.650 60.180 98.900 ;
        RECT 60.330 98.800 69.130 98.900 ;
        RECT 58.730 98.450 62.930 98.650 ;
        RECT 46.530 98.300 54.080 98.450 ;
        RECT 55.430 98.300 62.930 98.450 ;
        RECT 46.530 98.000 50.730 98.300 ;
        RECT 46.530 95.150 46.680 98.000 ;
        RECT 47.130 90.450 47.280 98.000 ;
        RECT 47.730 90.450 47.880 98.000 ;
        RECT 48.330 90.450 48.480 98.000 ;
        RECT 48.930 90.450 49.080 98.000 ;
        RECT 49.530 90.450 49.680 98.000 ;
        RECT 50.130 97.850 50.730 98.000 ;
        RECT 58.730 98.000 62.930 98.300 ;
        RECT 58.730 97.850 59.330 98.000 ;
        RECT 50.130 97.700 54.080 97.850 ;
        RECT 55.380 97.700 59.330 97.850 ;
        RECT 50.130 97.250 50.730 97.700 ;
        RECT 58.730 97.250 59.330 97.700 ;
        RECT 50.130 97.100 54.080 97.250 ;
        RECT 55.380 97.100 59.330 97.250 ;
        RECT 50.130 96.650 50.730 97.100 ;
        RECT 58.730 96.650 59.330 97.100 ;
        RECT 50.130 96.500 54.080 96.650 ;
        RECT 55.380 96.500 59.330 96.650 ;
        RECT 50.130 96.050 50.730 96.500 ;
        RECT 58.730 96.050 59.330 96.500 ;
        RECT 50.130 95.900 54.080 96.050 ;
        RECT 55.380 95.900 59.330 96.050 ;
        RECT 50.130 95.450 50.730 95.900 ;
        RECT 58.730 95.450 59.330 95.900 ;
        RECT 50.130 95.300 54.080 95.450 ;
        RECT 55.380 95.300 59.330 95.450 ;
        RECT 50.130 94.850 50.730 95.300 ;
        RECT 58.730 94.850 59.330 95.300 ;
        RECT 50.130 94.700 54.080 94.850 ;
        RECT 55.380 94.700 59.330 94.850 ;
        RECT 50.130 94.250 50.730 94.700 ;
        RECT 58.730 94.250 59.330 94.700 ;
        RECT 50.130 94.100 54.080 94.250 ;
        RECT 55.380 94.100 59.330 94.250 ;
        RECT 50.130 93.650 50.730 94.100 ;
        RECT 58.730 93.650 59.330 94.100 ;
        RECT 50.130 93.500 54.080 93.650 ;
        RECT 55.380 93.500 59.330 93.650 ;
        RECT 50.130 93.050 50.730 93.500 ;
        RECT 58.730 93.050 59.330 93.500 ;
        RECT 50.130 92.900 54.080 93.050 ;
        RECT 55.380 92.900 59.330 93.050 ;
        RECT 50.130 92.450 50.730 92.900 ;
        RECT 58.730 92.450 59.330 92.900 ;
        RECT 50.130 92.300 54.080 92.450 ;
        RECT 55.380 92.300 59.330 92.450 ;
        RECT 50.130 91.850 50.730 92.300 ;
        RECT 58.730 91.850 59.330 92.300 ;
        RECT 50.130 91.700 54.080 91.850 ;
        RECT 55.380 91.700 59.330 91.850 ;
        RECT 50.130 91.250 50.730 91.700 ;
        RECT 58.730 91.250 59.330 91.700 ;
        RECT 50.130 91.100 54.080 91.250 ;
        RECT 55.380 91.100 59.330 91.250 ;
        RECT 50.130 90.650 50.730 91.100 ;
        RECT 58.730 90.650 59.330 91.100 ;
        RECT 50.130 90.450 54.080 90.650 ;
        RECT 55.380 90.450 59.330 90.650 ;
        RECT 59.780 90.450 59.930 98.000 ;
        RECT 60.380 90.450 60.530 98.000 ;
        RECT 60.980 90.450 61.130 98.000 ;
        RECT 61.580 90.450 61.730 98.000 ;
        RECT 62.180 90.450 62.330 98.000 ;
        RECT 62.780 95.150 62.930 98.000 ;
        RECT 63.530 95.600 65.930 98.800 ;
        RECT 69.280 98.650 70.730 98.950 ;
        RECT 66.530 98.450 70.730 98.650 ;
        RECT 78.730 98.950 90.730 99.800 ;
        RECT 78.730 98.900 89.130 98.950 ;
        RECT 78.730 98.650 80.180 98.900 ;
        RECT 80.330 98.800 89.130 98.900 ;
        RECT 78.730 98.450 82.930 98.650 ;
        RECT 66.530 98.300 74.080 98.450 ;
        RECT 75.430 98.300 82.930 98.450 ;
        RECT 66.530 98.000 70.730 98.300 ;
        RECT 66.530 95.150 66.680 98.000 ;
        RECT 67.130 90.450 67.280 98.000 ;
        RECT 67.730 90.450 67.880 98.000 ;
        RECT 68.330 90.450 68.480 98.000 ;
        RECT 68.930 90.450 69.080 98.000 ;
        RECT 69.530 90.450 69.680 98.000 ;
        RECT 70.130 97.850 70.730 98.000 ;
        RECT 78.730 98.000 82.930 98.300 ;
        RECT 78.730 97.850 79.330 98.000 ;
        RECT 70.130 97.700 74.080 97.850 ;
        RECT 75.380 97.700 79.330 97.850 ;
        RECT 70.130 97.250 70.730 97.700 ;
        RECT 78.730 97.250 79.330 97.700 ;
        RECT 70.130 97.100 74.080 97.250 ;
        RECT 75.380 97.100 79.330 97.250 ;
        RECT 70.130 96.650 70.730 97.100 ;
        RECT 78.730 96.650 79.330 97.100 ;
        RECT 70.130 96.500 74.080 96.650 ;
        RECT 75.380 96.500 79.330 96.650 ;
        RECT 70.130 96.050 70.730 96.500 ;
        RECT 78.730 96.050 79.330 96.500 ;
        RECT 70.130 95.900 74.080 96.050 ;
        RECT 75.380 95.900 79.330 96.050 ;
        RECT 70.130 95.450 70.730 95.900 ;
        RECT 78.730 95.450 79.330 95.900 ;
        RECT 70.130 95.300 74.080 95.450 ;
        RECT 75.380 95.300 79.330 95.450 ;
        RECT 70.130 94.850 70.730 95.300 ;
        RECT 78.730 94.850 79.330 95.300 ;
        RECT 70.130 94.700 74.080 94.850 ;
        RECT 75.380 94.700 79.330 94.850 ;
        RECT 70.130 94.250 70.730 94.700 ;
        RECT 78.730 94.250 79.330 94.700 ;
        RECT 70.130 94.100 74.080 94.250 ;
        RECT 75.380 94.100 79.330 94.250 ;
        RECT 70.130 93.650 70.730 94.100 ;
        RECT 78.730 93.650 79.330 94.100 ;
        RECT 70.130 93.500 74.080 93.650 ;
        RECT 75.380 93.500 79.330 93.650 ;
        RECT 70.130 93.050 70.730 93.500 ;
        RECT 78.730 93.050 79.330 93.500 ;
        RECT 70.130 92.900 74.080 93.050 ;
        RECT 75.380 92.900 79.330 93.050 ;
        RECT 70.130 92.450 70.730 92.900 ;
        RECT 78.730 92.450 79.330 92.900 ;
        RECT 70.130 92.300 74.080 92.450 ;
        RECT 75.380 92.300 79.330 92.450 ;
        RECT 70.130 91.850 70.730 92.300 ;
        RECT 78.730 91.850 79.330 92.300 ;
        RECT 70.130 91.700 74.080 91.850 ;
        RECT 75.380 91.700 79.330 91.850 ;
        RECT 70.130 91.250 70.730 91.700 ;
        RECT 78.730 91.250 79.330 91.700 ;
        RECT 70.130 91.100 74.080 91.250 ;
        RECT 75.380 91.100 79.330 91.250 ;
        RECT 70.130 90.650 70.730 91.100 ;
        RECT 78.730 90.650 79.330 91.100 ;
        RECT 70.130 90.450 74.080 90.650 ;
        RECT 75.380 90.450 79.330 90.650 ;
        RECT 79.780 90.450 79.930 98.000 ;
        RECT 80.380 90.450 80.530 98.000 ;
        RECT 80.980 90.450 81.130 98.000 ;
        RECT 81.580 90.450 81.730 98.000 ;
        RECT 82.180 90.450 82.330 98.000 ;
        RECT 82.780 95.150 82.930 98.000 ;
        RECT 83.530 95.600 85.930 98.800 ;
        RECT 89.280 98.650 90.730 98.950 ;
        RECT 86.530 98.450 90.730 98.650 ;
        RECT 98.730 98.900 104.730 99.800 ;
        RECT 98.730 98.650 100.180 98.900 ;
        RECT 100.330 98.800 104.730 98.900 ;
        RECT 98.730 98.450 102.930 98.650 ;
        RECT 86.530 98.300 94.080 98.450 ;
        RECT 95.430 98.300 102.930 98.450 ;
        RECT 86.530 98.000 90.730 98.300 ;
        RECT 86.530 95.150 86.680 98.000 ;
        RECT 87.130 90.450 87.280 98.000 ;
        RECT 87.730 90.450 87.880 98.000 ;
        RECT 88.330 90.450 88.480 98.000 ;
        RECT 88.930 90.450 89.080 98.000 ;
        RECT 89.530 90.450 89.680 98.000 ;
        RECT 90.130 97.850 90.730 98.000 ;
        RECT 98.730 98.000 102.930 98.300 ;
        RECT 98.730 97.850 99.330 98.000 ;
        RECT 90.130 97.700 94.080 97.850 ;
        RECT 95.380 97.700 99.330 97.850 ;
        RECT 90.130 97.250 90.730 97.700 ;
        RECT 98.730 97.250 99.330 97.700 ;
        RECT 90.130 97.100 94.080 97.250 ;
        RECT 95.380 97.100 99.330 97.250 ;
        RECT 90.130 96.650 90.730 97.100 ;
        RECT 98.730 96.650 99.330 97.100 ;
        RECT 90.130 96.500 94.080 96.650 ;
        RECT 95.380 96.500 99.330 96.650 ;
        RECT 90.130 96.050 90.730 96.500 ;
        RECT 98.730 96.050 99.330 96.500 ;
        RECT 90.130 95.900 94.080 96.050 ;
        RECT 95.380 95.900 99.330 96.050 ;
        RECT 90.130 95.450 90.730 95.900 ;
        RECT 98.730 95.450 99.330 95.900 ;
        RECT 90.130 95.300 94.080 95.450 ;
        RECT 95.380 95.300 99.330 95.450 ;
        RECT 90.130 94.850 90.730 95.300 ;
        RECT 98.730 94.850 99.330 95.300 ;
        RECT 90.130 94.700 94.080 94.850 ;
        RECT 95.380 94.700 99.330 94.850 ;
        RECT 90.130 94.250 90.730 94.700 ;
        RECT 98.730 94.250 99.330 94.700 ;
        RECT 90.130 94.100 94.080 94.250 ;
        RECT 95.380 94.100 99.330 94.250 ;
        RECT 90.130 93.650 90.730 94.100 ;
        RECT 98.730 93.650 99.330 94.100 ;
        RECT 90.130 93.500 94.080 93.650 ;
        RECT 95.380 93.500 99.330 93.650 ;
        RECT 90.130 93.050 90.730 93.500 ;
        RECT 98.730 93.050 99.330 93.500 ;
        RECT 90.130 92.900 94.080 93.050 ;
        RECT 95.380 92.900 99.330 93.050 ;
        RECT 90.130 92.450 90.730 92.900 ;
        RECT 98.730 92.450 99.330 92.900 ;
        RECT 90.130 92.300 94.080 92.450 ;
        RECT 95.380 92.300 99.330 92.450 ;
        RECT 90.130 91.850 90.730 92.300 ;
        RECT 98.730 91.850 99.330 92.300 ;
        RECT 90.130 91.700 94.080 91.850 ;
        RECT 95.380 91.700 99.330 91.850 ;
        RECT 90.130 91.250 90.730 91.700 ;
        RECT 98.730 91.250 99.330 91.700 ;
        RECT 90.130 91.100 94.080 91.250 ;
        RECT 95.380 91.100 99.330 91.250 ;
        RECT 90.130 90.650 90.730 91.100 ;
        RECT 98.730 90.650 99.330 91.100 ;
        RECT 90.130 90.450 94.080 90.650 ;
        RECT 95.380 90.450 99.330 90.650 ;
        RECT 99.780 90.450 99.930 98.000 ;
        RECT 100.380 90.450 100.530 98.000 ;
        RECT 100.980 90.450 101.130 98.000 ;
        RECT 101.580 90.450 101.730 98.000 ;
        RECT 102.180 90.450 102.330 98.000 ;
        RECT 102.780 95.150 102.930 98.000 ;
        RECT 103.530 97.185 104.730 98.800 ;
        RECT 103.530 95.910 107.135 97.185 ;
        RECT 103.530 95.600 104.730 95.910 ;
        RECT 2.315 84.450 4.315 86.745 ;
        RECT 4.730 83.635 5.930 84.400 ;
        RECT 2.315 82.360 5.930 83.635 ;
        RECT 4.730 81.200 5.930 82.360 ;
        RECT 6.530 82.000 6.680 84.900 ;
        RECT 7.130 82.000 7.280 89.550 ;
        RECT 7.730 82.000 7.880 89.550 ;
        RECT 8.330 82.000 8.480 89.550 ;
        RECT 8.930 82.000 9.080 89.550 ;
        RECT 9.530 82.000 9.680 89.550 ;
        RECT 10.130 89.350 14.080 89.550 ;
        RECT 15.380 89.350 19.330 89.550 ;
        RECT 10.130 88.900 10.730 89.350 ;
        RECT 18.730 88.900 19.330 89.350 ;
        RECT 10.130 88.750 14.080 88.900 ;
        RECT 15.380 88.750 19.330 88.900 ;
        RECT 10.130 88.300 10.730 88.750 ;
        RECT 18.730 88.300 19.330 88.750 ;
        RECT 10.130 88.150 14.080 88.300 ;
        RECT 15.380 88.150 19.330 88.300 ;
        RECT 10.130 87.700 10.730 88.150 ;
        RECT 18.730 87.700 19.330 88.150 ;
        RECT 10.130 87.550 14.080 87.700 ;
        RECT 15.380 87.550 19.330 87.700 ;
        RECT 10.130 87.100 10.730 87.550 ;
        RECT 18.730 87.100 19.330 87.550 ;
        RECT 10.130 86.950 14.080 87.100 ;
        RECT 15.380 86.950 19.330 87.100 ;
        RECT 10.130 86.500 10.730 86.950 ;
        RECT 18.730 86.500 19.330 86.950 ;
        RECT 10.130 86.350 14.080 86.500 ;
        RECT 15.380 86.350 19.330 86.500 ;
        RECT 10.130 85.900 10.730 86.350 ;
        RECT 18.730 85.900 19.330 86.350 ;
        RECT 10.130 85.750 14.080 85.900 ;
        RECT 15.380 85.750 19.330 85.900 ;
        RECT 10.130 85.300 10.730 85.750 ;
        RECT 18.730 85.300 19.330 85.750 ;
        RECT 10.130 85.150 14.080 85.300 ;
        RECT 15.380 85.150 19.330 85.300 ;
        RECT 10.130 84.700 10.730 85.150 ;
        RECT 18.730 84.700 19.330 85.150 ;
        RECT 10.130 84.550 14.080 84.700 ;
        RECT 15.380 84.550 19.330 84.700 ;
        RECT 10.130 84.100 10.730 84.550 ;
        RECT 18.730 84.100 19.330 84.550 ;
        RECT 10.130 83.950 14.080 84.100 ;
        RECT 15.380 83.950 19.330 84.100 ;
        RECT 10.130 83.500 10.730 83.950 ;
        RECT 18.730 83.500 19.330 83.950 ;
        RECT 10.130 83.350 14.080 83.500 ;
        RECT 15.380 83.350 19.330 83.500 ;
        RECT 10.130 82.900 10.730 83.350 ;
        RECT 18.730 82.900 19.330 83.350 ;
        RECT 10.130 82.750 14.080 82.900 ;
        RECT 15.380 82.750 19.330 82.900 ;
        RECT 10.130 82.300 10.730 82.750 ;
        RECT 18.730 82.300 19.330 82.750 ;
        RECT 10.130 82.150 14.080 82.300 ;
        RECT 15.380 82.150 19.330 82.300 ;
        RECT 10.130 82.000 10.730 82.150 ;
        RECT 6.530 81.700 10.730 82.000 ;
        RECT 18.730 82.000 19.330 82.150 ;
        RECT 19.780 82.000 19.930 89.550 ;
        RECT 20.380 82.000 20.530 89.550 ;
        RECT 20.980 82.000 21.130 89.550 ;
        RECT 21.580 82.000 21.730 89.550 ;
        RECT 22.180 82.000 22.330 89.550 ;
        RECT 22.780 82.000 22.930 84.900 ;
        RECT 18.730 81.700 22.930 82.000 ;
        RECT 6.530 81.550 14.080 81.700 ;
        RECT 15.380 81.550 22.930 81.700 ;
        RECT 6.530 81.350 10.730 81.550 ;
        RECT 4.730 81.050 9.130 81.200 ;
        RECT 9.280 81.050 10.730 81.350 ;
        RECT 4.730 80.150 10.730 81.050 ;
        RECT 18.730 81.350 22.930 81.550 ;
        RECT 18.730 81.050 20.180 81.350 ;
        RECT 23.530 81.200 25.930 84.400 ;
        RECT 26.530 82.000 26.680 84.900 ;
        RECT 27.130 82.000 27.280 89.550 ;
        RECT 27.730 82.000 27.880 89.550 ;
        RECT 28.330 82.000 28.480 89.550 ;
        RECT 28.930 82.000 29.080 89.550 ;
        RECT 29.530 82.000 29.680 89.550 ;
        RECT 30.130 89.350 34.080 89.550 ;
        RECT 35.380 89.350 39.330 89.550 ;
        RECT 30.130 88.900 30.730 89.350 ;
        RECT 38.730 88.900 39.330 89.350 ;
        RECT 30.130 88.750 34.080 88.900 ;
        RECT 35.380 88.750 39.330 88.900 ;
        RECT 30.130 88.300 30.730 88.750 ;
        RECT 38.730 88.300 39.330 88.750 ;
        RECT 30.130 88.150 34.080 88.300 ;
        RECT 35.380 88.150 39.330 88.300 ;
        RECT 30.130 87.700 30.730 88.150 ;
        RECT 38.730 87.700 39.330 88.150 ;
        RECT 30.130 87.550 34.080 87.700 ;
        RECT 35.380 87.550 39.330 87.700 ;
        RECT 30.130 87.100 30.730 87.550 ;
        RECT 38.730 87.100 39.330 87.550 ;
        RECT 30.130 86.950 34.080 87.100 ;
        RECT 35.380 86.950 39.330 87.100 ;
        RECT 30.130 86.500 30.730 86.950 ;
        RECT 38.730 86.500 39.330 86.950 ;
        RECT 30.130 86.350 34.080 86.500 ;
        RECT 35.380 86.350 39.330 86.500 ;
        RECT 30.130 85.900 30.730 86.350 ;
        RECT 38.730 85.900 39.330 86.350 ;
        RECT 30.130 85.750 34.080 85.900 ;
        RECT 35.380 85.750 39.330 85.900 ;
        RECT 30.130 85.300 30.730 85.750 ;
        RECT 38.730 85.300 39.330 85.750 ;
        RECT 30.130 85.150 34.080 85.300 ;
        RECT 35.380 85.150 39.330 85.300 ;
        RECT 30.130 84.700 30.730 85.150 ;
        RECT 38.730 84.700 39.330 85.150 ;
        RECT 30.130 84.550 34.080 84.700 ;
        RECT 35.380 84.550 39.330 84.700 ;
        RECT 30.130 84.100 30.730 84.550 ;
        RECT 38.730 84.100 39.330 84.550 ;
        RECT 30.130 83.950 34.080 84.100 ;
        RECT 35.380 83.950 39.330 84.100 ;
        RECT 30.130 83.500 30.730 83.950 ;
        RECT 38.730 83.500 39.330 83.950 ;
        RECT 30.130 83.350 34.080 83.500 ;
        RECT 35.380 83.350 39.330 83.500 ;
        RECT 30.130 82.900 30.730 83.350 ;
        RECT 38.730 82.900 39.330 83.350 ;
        RECT 30.130 82.750 34.080 82.900 ;
        RECT 35.380 82.750 39.330 82.900 ;
        RECT 30.130 82.300 30.730 82.750 ;
        RECT 38.730 82.300 39.330 82.750 ;
        RECT 30.130 82.150 34.080 82.300 ;
        RECT 35.380 82.150 39.330 82.300 ;
        RECT 30.130 82.000 30.730 82.150 ;
        RECT 26.530 81.700 30.730 82.000 ;
        RECT 38.730 82.000 39.330 82.150 ;
        RECT 39.780 82.000 39.930 89.550 ;
        RECT 40.380 82.000 40.530 89.550 ;
        RECT 40.980 82.000 41.130 89.550 ;
        RECT 41.580 82.000 41.730 89.550 ;
        RECT 42.180 82.000 42.330 89.550 ;
        RECT 42.780 82.000 42.930 84.900 ;
        RECT 38.730 81.700 42.930 82.000 ;
        RECT 26.530 81.550 34.080 81.700 ;
        RECT 35.380 81.550 42.930 81.700 ;
        RECT 26.530 81.350 30.730 81.550 ;
        RECT 20.330 81.050 29.130 81.200 ;
        RECT 29.280 81.050 30.730 81.350 ;
        RECT 18.730 80.150 30.730 81.050 ;
        RECT 38.730 81.350 42.930 81.550 ;
        RECT 38.730 81.050 40.180 81.350 ;
        RECT 43.530 81.200 45.930 84.400 ;
        RECT 46.530 82.000 46.680 84.900 ;
        RECT 47.130 82.000 47.280 89.550 ;
        RECT 47.730 82.000 47.880 89.550 ;
        RECT 48.330 82.000 48.480 89.550 ;
        RECT 48.930 82.000 49.080 89.550 ;
        RECT 49.530 82.000 49.680 89.550 ;
        RECT 50.130 89.350 54.080 89.550 ;
        RECT 55.380 89.350 59.330 89.550 ;
        RECT 50.130 88.900 50.730 89.350 ;
        RECT 58.730 88.900 59.330 89.350 ;
        RECT 50.130 88.750 54.080 88.900 ;
        RECT 55.380 88.750 59.330 88.900 ;
        RECT 50.130 88.300 50.730 88.750 ;
        RECT 58.730 88.300 59.330 88.750 ;
        RECT 50.130 88.150 54.080 88.300 ;
        RECT 55.380 88.150 59.330 88.300 ;
        RECT 50.130 87.700 50.730 88.150 ;
        RECT 58.730 87.700 59.330 88.150 ;
        RECT 50.130 87.550 54.080 87.700 ;
        RECT 55.380 87.550 59.330 87.700 ;
        RECT 50.130 87.100 50.730 87.550 ;
        RECT 58.730 87.100 59.330 87.550 ;
        RECT 50.130 86.950 54.080 87.100 ;
        RECT 55.380 86.950 59.330 87.100 ;
        RECT 50.130 86.500 50.730 86.950 ;
        RECT 58.730 86.500 59.330 86.950 ;
        RECT 50.130 86.350 54.080 86.500 ;
        RECT 55.380 86.350 59.330 86.500 ;
        RECT 50.130 85.900 50.730 86.350 ;
        RECT 58.730 85.900 59.330 86.350 ;
        RECT 50.130 85.750 54.080 85.900 ;
        RECT 55.380 85.750 59.330 85.900 ;
        RECT 50.130 85.300 50.730 85.750 ;
        RECT 58.730 85.300 59.330 85.750 ;
        RECT 50.130 85.150 54.080 85.300 ;
        RECT 55.380 85.150 59.330 85.300 ;
        RECT 50.130 84.700 50.730 85.150 ;
        RECT 58.730 84.700 59.330 85.150 ;
        RECT 50.130 84.550 54.080 84.700 ;
        RECT 55.380 84.550 59.330 84.700 ;
        RECT 50.130 84.100 50.730 84.550 ;
        RECT 58.730 84.100 59.330 84.550 ;
        RECT 50.130 83.950 54.080 84.100 ;
        RECT 55.380 83.950 59.330 84.100 ;
        RECT 50.130 83.500 50.730 83.950 ;
        RECT 58.730 83.500 59.330 83.950 ;
        RECT 50.130 83.350 54.080 83.500 ;
        RECT 55.380 83.350 59.330 83.500 ;
        RECT 50.130 82.900 50.730 83.350 ;
        RECT 58.730 82.900 59.330 83.350 ;
        RECT 50.130 82.750 54.080 82.900 ;
        RECT 55.380 82.750 59.330 82.900 ;
        RECT 50.130 82.300 50.730 82.750 ;
        RECT 58.730 82.300 59.330 82.750 ;
        RECT 50.130 82.150 54.080 82.300 ;
        RECT 55.380 82.150 59.330 82.300 ;
        RECT 50.130 82.000 50.730 82.150 ;
        RECT 46.530 81.700 50.730 82.000 ;
        RECT 58.730 82.000 59.330 82.150 ;
        RECT 59.780 82.000 59.930 89.550 ;
        RECT 60.380 82.000 60.530 89.550 ;
        RECT 60.980 82.000 61.130 89.550 ;
        RECT 61.580 82.000 61.730 89.550 ;
        RECT 62.180 82.000 62.330 89.550 ;
        RECT 62.780 82.000 62.930 84.900 ;
        RECT 58.730 81.700 62.930 82.000 ;
        RECT 46.530 81.550 54.080 81.700 ;
        RECT 55.380 81.550 62.930 81.700 ;
        RECT 46.530 81.350 50.730 81.550 ;
        RECT 40.330 81.050 49.130 81.200 ;
        RECT 49.280 81.050 50.730 81.350 ;
        RECT 38.730 80.150 50.730 81.050 ;
        RECT 58.730 81.350 62.930 81.550 ;
        RECT 58.730 81.050 60.180 81.350 ;
        RECT 63.530 81.200 65.930 84.400 ;
        RECT 66.530 82.000 66.680 84.900 ;
        RECT 67.130 82.000 67.280 89.550 ;
        RECT 67.730 82.000 67.880 89.550 ;
        RECT 68.330 82.000 68.480 89.550 ;
        RECT 68.930 82.000 69.080 89.550 ;
        RECT 69.530 82.000 69.680 89.550 ;
        RECT 70.130 89.350 74.080 89.550 ;
        RECT 75.380 89.350 79.330 89.550 ;
        RECT 70.130 88.900 70.730 89.350 ;
        RECT 78.730 88.900 79.330 89.350 ;
        RECT 70.130 88.750 74.080 88.900 ;
        RECT 75.380 88.750 79.330 88.900 ;
        RECT 70.130 88.300 70.730 88.750 ;
        RECT 78.730 88.300 79.330 88.750 ;
        RECT 70.130 88.150 74.080 88.300 ;
        RECT 75.380 88.150 79.330 88.300 ;
        RECT 70.130 87.700 70.730 88.150 ;
        RECT 78.730 87.700 79.330 88.150 ;
        RECT 70.130 87.550 74.080 87.700 ;
        RECT 75.380 87.550 79.330 87.700 ;
        RECT 70.130 87.100 70.730 87.550 ;
        RECT 78.730 87.100 79.330 87.550 ;
        RECT 70.130 86.950 74.080 87.100 ;
        RECT 75.380 86.950 79.330 87.100 ;
        RECT 70.130 86.500 70.730 86.950 ;
        RECT 78.730 86.500 79.330 86.950 ;
        RECT 70.130 86.350 74.080 86.500 ;
        RECT 75.380 86.350 79.330 86.500 ;
        RECT 70.130 85.900 70.730 86.350 ;
        RECT 78.730 85.900 79.330 86.350 ;
        RECT 70.130 85.750 74.080 85.900 ;
        RECT 75.380 85.750 79.330 85.900 ;
        RECT 70.130 85.300 70.730 85.750 ;
        RECT 78.730 85.300 79.330 85.750 ;
        RECT 70.130 85.150 74.080 85.300 ;
        RECT 75.380 85.150 79.330 85.300 ;
        RECT 70.130 84.700 70.730 85.150 ;
        RECT 78.730 84.700 79.330 85.150 ;
        RECT 70.130 84.550 74.080 84.700 ;
        RECT 75.380 84.550 79.330 84.700 ;
        RECT 70.130 84.100 70.730 84.550 ;
        RECT 78.730 84.100 79.330 84.550 ;
        RECT 70.130 83.950 74.080 84.100 ;
        RECT 75.380 83.950 79.330 84.100 ;
        RECT 70.130 83.500 70.730 83.950 ;
        RECT 78.730 83.500 79.330 83.950 ;
        RECT 70.130 83.350 74.080 83.500 ;
        RECT 75.380 83.350 79.330 83.500 ;
        RECT 70.130 82.900 70.730 83.350 ;
        RECT 78.730 82.900 79.330 83.350 ;
        RECT 70.130 82.750 74.080 82.900 ;
        RECT 75.380 82.750 79.330 82.900 ;
        RECT 70.130 82.300 70.730 82.750 ;
        RECT 78.730 82.300 79.330 82.750 ;
        RECT 70.130 82.150 74.080 82.300 ;
        RECT 75.380 82.150 79.330 82.300 ;
        RECT 70.130 82.000 70.730 82.150 ;
        RECT 66.530 81.700 70.730 82.000 ;
        RECT 78.730 82.000 79.330 82.150 ;
        RECT 79.780 82.000 79.930 89.550 ;
        RECT 80.380 82.000 80.530 89.550 ;
        RECT 80.980 82.000 81.130 89.550 ;
        RECT 81.580 82.000 81.730 89.550 ;
        RECT 82.180 82.000 82.330 89.550 ;
        RECT 82.780 82.000 82.930 84.900 ;
        RECT 78.730 81.700 82.930 82.000 ;
        RECT 66.530 81.550 74.080 81.700 ;
        RECT 75.380 81.550 82.930 81.700 ;
        RECT 66.530 81.350 70.730 81.550 ;
        RECT 60.330 81.050 69.130 81.200 ;
        RECT 69.280 81.050 70.730 81.350 ;
        RECT 58.730 80.150 70.730 81.050 ;
        RECT 78.730 81.350 82.930 81.550 ;
        RECT 78.730 81.050 80.180 81.350 ;
        RECT 83.530 81.200 85.930 84.400 ;
        RECT 86.530 82.000 86.680 84.900 ;
        RECT 87.130 82.000 87.280 89.550 ;
        RECT 87.730 82.000 87.880 89.550 ;
        RECT 88.330 82.000 88.480 89.550 ;
        RECT 88.930 82.000 89.080 89.550 ;
        RECT 89.530 82.000 89.680 89.550 ;
        RECT 90.130 89.350 94.080 89.550 ;
        RECT 95.380 89.350 99.330 89.550 ;
        RECT 90.130 88.900 90.730 89.350 ;
        RECT 98.730 88.900 99.330 89.350 ;
        RECT 90.130 88.750 94.080 88.900 ;
        RECT 95.380 88.750 99.330 88.900 ;
        RECT 90.130 88.300 90.730 88.750 ;
        RECT 98.730 88.300 99.330 88.750 ;
        RECT 90.130 88.150 94.080 88.300 ;
        RECT 95.380 88.150 99.330 88.300 ;
        RECT 90.130 87.700 90.730 88.150 ;
        RECT 98.730 87.700 99.330 88.150 ;
        RECT 90.130 87.550 94.080 87.700 ;
        RECT 95.380 87.550 99.330 87.700 ;
        RECT 90.130 87.100 90.730 87.550 ;
        RECT 98.730 87.100 99.330 87.550 ;
        RECT 90.130 86.950 94.080 87.100 ;
        RECT 95.380 86.950 99.330 87.100 ;
        RECT 90.130 86.500 90.730 86.950 ;
        RECT 98.730 86.500 99.330 86.950 ;
        RECT 90.130 86.350 94.080 86.500 ;
        RECT 95.380 86.350 99.330 86.500 ;
        RECT 90.130 85.900 90.730 86.350 ;
        RECT 98.730 85.900 99.330 86.350 ;
        RECT 90.130 85.750 94.080 85.900 ;
        RECT 95.380 85.750 99.330 85.900 ;
        RECT 90.130 85.300 90.730 85.750 ;
        RECT 98.730 85.300 99.330 85.750 ;
        RECT 90.130 85.150 94.080 85.300 ;
        RECT 95.380 85.150 99.330 85.300 ;
        RECT 90.130 84.700 90.730 85.150 ;
        RECT 98.730 84.700 99.330 85.150 ;
        RECT 90.130 84.550 94.080 84.700 ;
        RECT 95.380 84.550 99.330 84.700 ;
        RECT 90.130 84.100 90.730 84.550 ;
        RECT 98.730 84.100 99.330 84.550 ;
        RECT 90.130 83.950 94.080 84.100 ;
        RECT 95.380 83.950 99.330 84.100 ;
        RECT 90.130 83.500 90.730 83.950 ;
        RECT 98.730 83.500 99.330 83.950 ;
        RECT 90.130 83.350 94.080 83.500 ;
        RECT 95.380 83.350 99.330 83.500 ;
        RECT 90.130 82.900 90.730 83.350 ;
        RECT 98.730 82.900 99.330 83.350 ;
        RECT 90.130 82.750 94.080 82.900 ;
        RECT 95.380 82.750 99.330 82.900 ;
        RECT 90.130 82.300 90.730 82.750 ;
        RECT 98.730 82.300 99.330 82.750 ;
        RECT 90.130 82.150 94.080 82.300 ;
        RECT 95.380 82.150 99.330 82.300 ;
        RECT 90.130 82.000 90.730 82.150 ;
        RECT 86.530 81.700 90.730 82.000 ;
        RECT 98.730 82.000 99.330 82.150 ;
        RECT 99.780 82.000 99.930 89.550 ;
        RECT 100.380 82.000 100.530 89.550 ;
        RECT 100.980 82.000 101.130 89.550 ;
        RECT 101.580 82.000 101.730 89.550 ;
        RECT 102.180 82.000 102.330 89.550 ;
        RECT 102.780 82.000 102.930 84.900 ;
        RECT 98.730 81.700 102.930 82.000 ;
        RECT 86.530 81.550 94.080 81.700 ;
        RECT 95.380 81.550 102.930 81.700 ;
        RECT 86.530 81.350 90.730 81.550 ;
        RECT 80.330 81.050 89.130 81.200 ;
        RECT 89.280 81.050 90.730 81.350 ;
        RECT 78.730 80.150 90.730 81.050 ;
        RECT 98.730 81.350 102.930 81.550 ;
        RECT 103.530 83.380 104.730 84.400 ;
        RECT 103.530 82.105 107.135 83.380 ;
        RECT 98.730 81.050 100.180 81.350 ;
        RECT 103.530 81.200 104.730 82.105 ;
        RECT 100.330 81.050 104.730 81.200 ;
        RECT 98.730 80.150 104.730 81.050 ;
        RECT 4.730 79.850 9.130 80.150 ;
        RECT 20.330 79.850 29.130 80.150 ;
        RECT 40.330 79.850 49.130 80.150 ;
        RECT 60.330 79.850 69.130 80.150 ;
        RECT 80.330 79.850 89.130 80.150 ;
        RECT 4.730 78.950 10.730 79.850 ;
        RECT 20.330 79.800 30.730 79.850 ;
        RECT 40.330 79.800 50.730 79.850 ;
        RECT 60.330 79.800 70.730 79.850 ;
        RECT 80.330 79.800 90.730 79.850 ;
        RECT 100.330 79.800 104.730 80.150 ;
        RECT 4.730 78.800 9.130 78.950 ;
        RECT 4.730 77.555 5.930 78.800 ;
        RECT 9.280 78.650 10.730 78.950 ;
        RECT 2.315 76.280 5.930 77.555 ;
        RECT 4.730 75.600 5.930 76.280 ;
        RECT 6.530 78.450 10.730 78.650 ;
        RECT 18.730 78.950 30.730 79.800 ;
        RECT 18.730 78.900 29.130 78.950 ;
        RECT 18.730 78.650 20.180 78.900 ;
        RECT 20.330 78.800 29.130 78.900 ;
        RECT 18.730 78.450 22.930 78.650 ;
        RECT 6.530 78.300 14.080 78.450 ;
        RECT 15.430 78.300 22.930 78.450 ;
        RECT 6.530 78.000 10.730 78.300 ;
        RECT 2.315 73.250 4.315 75.545 ;
        RECT 6.530 75.150 6.680 78.000 ;
        RECT 7.130 70.450 7.280 78.000 ;
        RECT 7.730 70.450 7.880 78.000 ;
        RECT 8.330 70.450 8.480 78.000 ;
        RECT 8.930 70.450 9.080 78.000 ;
        RECT 9.530 70.450 9.680 78.000 ;
        RECT 10.130 77.850 10.730 78.000 ;
        RECT 18.730 78.000 22.930 78.300 ;
        RECT 18.730 77.850 19.330 78.000 ;
        RECT 10.130 77.700 14.080 77.850 ;
        RECT 15.380 77.700 19.330 77.850 ;
        RECT 10.130 77.250 10.730 77.700 ;
        RECT 18.730 77.250 19.330 77.700 ;
        RECT 10.130 77.100 14.080 77.250 ;
        RECT 15.380 77.100 19.330 77.250 ;
        RECT 10.130 76.650 10.730 77.100 ;
        RECT 18.730 76.650 19.330 77.100 ;
        RECT 10.130 76.500 14.080 76.650 ;
        RECT 15.380 76.500 19.330 76.650 ;
        RECT 10.130 76.050 10.730 76.500 ;
        RECT 18.730 76.050 19.330 76.500 ;
        RECT 10.130 75.900 14.080 76.050 ;
        RECT 15.380 75.900 19.330 76.050 ;
        RECT 10.130 75.450 10.730 75.900 ;
        RECT 18.730 75.450 19.330 75.900 ;
        RECT 10.130 75.300 14.080 75.450 ;
        RECT 15.380 75.300 19.330 75.450 ;
        RECT 10.130 74.850 10.730 75.300 ;
        RECT 18.730 74.850 19.330 75.300 ;
        RECT 10.130 74.700 14.080 74.850 ;
        RECT 15.380 74.700 19.330 74.850 ;
        RECT 10.130 74.250 10.730 74.700 ;
        RECT 18.730 74.250 19.330 74.700 ;
        RECT 10.130 74.100 14.080 74.250 ;
        RECT 15.380 74.100 19.330 74.250 ;
        RECT 10.130 73.650 10.730 74.100 ;
        RECT 18.730 73.650 19.330 74.100 ;
        RECT 10.130 73.500 14.080 73.650 ;
        RECT 15.380 73.500 19.330 73.650 ;
        RECT 10.130 73.050 10.730 73.500 ;
        RECT 18.730 73.050 19.330 73.500 ;
        RECT 10.130 72.900 14.080 73.050 ;
        RECT 15.380 72.900 19.330 73.050 ;
        RECT 10.130 72.450 10.730 72.900 ;
        RECT 18.730 72.450 19.330 72.900 ;
        RECT 10.130 72.300 14.080 72.450 ;
        RECT 15.380 72.300 19.330 72.450 ;
        RECT 10.130 71.850 10.730 72.300 ;
        RECT 18.730 71.850 19.330 72.300 ;
        RECT 10.130 71.700 14.080 71.850 ;
        RECT 15.380 71.700 19.330 71.850 ;
        RECT 10.130 71.250 10.730 71.700 ;
        RECT 18.730 71.250 19.330 71.700 ;
        RECT 10.130 71.100 14.080 71.250 ;
        RECT 15.380 71.100 19.330 71.250 ;
        RECT 10.130 70.650 10.730 71.100 ;
        RECT 18.730 70.650 19.330 71.100 ;
        RECT 10.130 70.450 14.080 70.650 ;
        RECT 15.380 70.450 19.330 70.650 ;
        RECT 19.780 70.450 19.930 78.000 ;
        RECT 20.380 70.450 20.530 78.000 ;
        RECT 20.980 70.450 21.130 78.000 ;
        RECT 21.580 70.450 21.730 78.000 ;
        RECT 22.180 70.450 22.330 78.000 ;
        RECT 22.780 75.150 22.930 78.000 ;
        RECT 23.530 75.600 25.930 78.800 ;
        RECT 29.280 78.650 30.730 78.950 ;
        RECT 26.530 78.450 30.730 78.650 ;
        RECT 38.730 78.950 50.730 79.800 ;
        RECT 38.730 78.900 49.130 78.950 ;
        RECT 38.730 78.650 40.180 78.900 ;
        RECT 40.330 78.800 49.130 78.900 ;
        RECT 38.730 78.450 42.930 78.650 ;
        RECT 26.530 78.300 34.080 78.450 ;
        RECT 35.430 78.300 42.930 78.450 ;
        RECT 26.530 78.000 30.730 78.300 ;
        RECT 26.530 75.150 26.680 78.000 ;
        RECT 27.130 70.450 27.280 78.000 ;
        RECT 27.730 70.450 27.880 78.000 ;
        RECT 28.330 70.450 28.480 78.000 ;
        RECT 28.930 70.450 29.080 78.000 ;
        RECT 29.530 70.450 29.680 78.000 ;
        RECT 30.130 77.850 30.730 78.000 ;
        RECT 38.730 78.000 42.930 78.300 ;
        RECT 38.730 77.850 39.330 78.000 ;
        RECT 30.130 77.700 34.080 77.850 ;
        RECT 35.380 77.700 39.330 77.850 ;
        RECT 30.130 77.250 30.730 77.700 ;
        RECT 38.730 77.250 39.330 77.700 ;
        RECT 30.130 77.100 34.080 77.250 ;
        RECT 35.380 77.100 39.330 77.250 ;
        RECT 30.130 76.650 30.730 77.100 ;
        RECT 38.730 76.650 39.330 77.100 ;
        RECT 30.130 76.500 34.080 76.650 ;
        RECT 35.380 76.500 39.330 76.650 ;
        RECT 30.130 76.050 30.730 76.500 ;
        RECT 38.730 76.050 39.330 76.500 ;
        RECT 30.130 75.900 34.080 76.050 ;
        RECT 35.380 75.900 39.330 76.050 ;
        RECT 30.130 75.450 30.730 75.900 ;
        RECT 38.730 75.450 39.330 75.900 ;
        RECT 30.130 75.300 34.080 75.450 ;
        RECT 35.380 75.300 39.330 75.450 ;
        RECT 30.130 74.850 30.730 75.300 ;
        RECT 38.730 74.850 39.330 75.300 ;
        RECT 30.130 74.700 34.080 74.850 ;
        RECT 35.380 74.700 39.330 74.850 ;
        RECT 30.130 74.250 30.730 74.700 ;
        RECT 38.730 74.250 39.330 74.700 ;
        RECT 30.130 74.100 34.080 74.250 ;
        RECT 35.380 74.100 39.330 74.250 ;
        RECT 30.130 73.650 30.730 74.100 ;
        RECT 38.730 73.650 39.330 74.100 ;
        RECT 30.130 73.500 34.080 73.650 ;
        RECT 35.380 73.500 39.330 73.650 ;
        RECT 30.130 73.050 30.730 73.500 ;
        RECT 38.730 73.050 39.330 73.500 ;
        RECT 30.130 72.900 34.080 73.050 ;
        RECT 35.380 72.900 39.330 73.050 ;
        RECT 30.130 72.450 30.730 72.900 ;
        RECT 38.730 72.450 39.330 72.900 ;
        RECT 30.130 72.300 34.080 72.450 ;
        RECT 35.380 72.300 39.330 72.450 ;
        RECT 30.130 71.850 30.730 72.300 ;
        RECT 38.730 71.850 39.330 72.300 ;
        RECT 30.130 71.700 34.080 71.850 ;
        RECT 35.380 71.700 39.330 71.850 ;
        RECT 30.130 71.250 30.730 71.700 ;
        RECT 38.730 71.250 39.330 71.700 ;
        RECT 30.130 71.100 34.080 71.250 ;
        RECT 35.380 71.100 39.330 71.250 ;
        RECT 30.130 70.650 30.730 71.100 ;
        RECT 38.730 70.650 39.330 71.100 ;
        RECT 30.130 70.450 34.080 70.650 ;
        RECT 35.380 70.450 39.330 70.650 ;
        RECT 39.780 70.450 39.930 78.000 ;
        RECT 40.380 70.450 40.530 78.000 ;
        RECT 40.980 70.450 41.130 78.000 ;
        RECT 41.580 70.450 41.730 78.000 ;
        RECT 42.180 70.450 42.330 78.000 ;
        RECT 42.780 75.150 42.930 78.000 ;
        RECT 43.530 75.600 45.930 78.800 ;
        RECT 49.280 78.650 50.730 78.950 ;
        RECT 46.530 78.450 50.730 78.650 ;
        RECT 58.730 78.950 70.730 79.800 ;
        RECT 58.730 78.900 69.130 78.950 ;
        RECT 58.730 78.650 60.180 78.900 ;
        RECT 60.330 78.800 69.130 78.900 ;
        RECT 58.730 78.450 62.930 78.650 ;
        RECT 46.530 78.300 54.080 78.450 ;
        RECT 55.430 78.300 62.930 78.450 ;
        RECT 46.530 78.000 50.730 78.300 ;
        RECT 46.530 75.150 46.680 78.000 ;
        RECT 47.130 70.450 47.280 78.000 ;
        RECT 47.730 70.450 47.880 78.000 ;
        RECT 48.330 70.450 48.480 78.000 ;
        RECT 48.930 70.450 49.080 78.000 ;
        RECT 49.530 70.450 49.680 78.000 ;
        RECT 50.130 77.850 50.730 78.000 ;
        RECT 58.730 78.000 62.930 78.300 ;
        RECT 58.730 77.850 59.330 78.000 ;
        RECT 50.130 77.700 54.080 77.850 ;
        RECT 55.380 77.700 59.330 77.850 ;
        RECT 50.130 77.250 50.730 77.700 ;
        RECT 58.730 77.250 59.330 77.700 ;
        RECT 50.130 77.100 54.080 77.250 ;
        RECT 55.380 77.100 59.330 77.250 ;
        RECT 50.130 76.650 50.730 77.100 ;
        RECT 58.730 76.650 59.330 77.100 ;
        RECT 50.130 76.500 54.080 76.650 ;
        RECT 55.380 76.500 59.330 76.650 ;
        RECT 50.130 76.050 50.730 76.500 ;
        RECT 58.730 76.050 59.330 76.500 ;
        RECT 50.130 75.900 54.080 76.050 ;
        RECT 55.380 75.900 59.330 76.050 ;
        RECT 50.130 75.450 50.730 75.900 ;
        RECT 58.730 75.450 59.330 75.900 ;
        RECT 50.130 75.300 54.080 75.450 ;
        RECT 55.380 75.300 59.330 75.450 ;
        RECT 50.130 74.850 50.730 75.300 ;
        RECT 58.730 74.850 59.330 75.300 ;
        RECT 50.130 74.700 54.080 74.850 ;
        RECT 55.380 74.700 59.330 74.850 ;
        RECT 50.130 74.250 50.730 74.700 ;
        RECT 58.730 74.250 59.330 74.700 ;
        RECT 50.130 74.100 54.080 74.250 ;
        RECT 55.380 74.100 59.330 74.250 ;
        RECT 50.130 73.650 50.730 74.100 ;
        RECT 58.730 73.650 59.330 74.100 ;
        RECT 50.130 73.500 54.080 73.650 ;
        RECT 55.380 73.500 59.330 73.650 ;
        RECT 50.130 73.050 50.730 73.500 ;
        RECT 58.730 73.050 59.330 73.500 ;
        RECT 50.130 72.900 54.080 73.050 ;
        RECT 55.380 72.900 59.330 73.050 ;
        RECT 50.130 72.450 50.730 72.900 ;
        RECT 58.730 72.450 59.330 72.900 ;
        RECT 50.130 72.300 54.080 72.450 ;
        RECT 55.380 72.300 59.330 72.450 ;
        RECT 50.130 71.850 50.730 72.300 ;
        RECT 58.730 71.850 59.330 72.300 ;
        RECT 50.130 71.700 54.080 71.850 ;
        RECT 55.380 71.700 59.330 71.850 ;
        RECT 50.130 71.250 50.730 71.700 ;
        RECT 58.730 71.250 59.330 71.700 ;
        RECT 50.130 71.100 54.080 71.250 ;
        RECT 55.380 71.100 59.330 71.250 ;
        RECT 50.130 70.650 50.730 71.100 ;
        RECT 58.730 70.650 59.330 71.100 ;
        RECT 50.130 70.450 54.080 70.650 ;
        RECT 55.380 70.450 59.330 70.650 ;
        RECT 59.780 70.450 59.930 78.000 ;
        RECT 60.380 70.450 60.530 78.000 ;
        RECT 60.980 70.450 61.130 78.000 ;
        RECT 61.580 70.450 61.730 78.000 ;
        RECT 62.180 70.450 62.330 78.000 ;
        RECT 62.780 75.150 62.930 78.000 ;
        RECT 63.530 75.600 65.930 78.800 ;
        RECT 69.280 78.650 70.730 78.950 ;
        RECT 66.530 78.450 70.730 78.650 ;
        RECT 78.730 78.950 90.730 79.800 ;
        RECT 78.730 78.900 89.130 78.950 ;
        RECT 78.730 78.650 80.180 78.900 ;
        RECT 80.330 78.800 89.130 78.900 ;
        RECT 78.730 78.450 82.930 78.650 ;
        RECT 66.530 78.300 74.080 78.450 ;
        RECT 75.430 78.300 82.930 78.450 ;
        RECT 66.530 78.000 70.730 78.300 ;
        RECT 66.530 75.150 66.680 78.000 ;
        RECT 67.130 70.450 67.280 78.000 ;
        RECT 67.730 70.450 67.880 78.000 ;
        RECT 68.330 70.450 68.480 78.000 ;
        RECT 68.930 70.450 69.080 78.000 ;
        RECT 69.530 70.450 69.680 78.000 ;
        RECT 70.130 77.850 70.730 78.000 ;
        RECT 78.730 78.000 82.930 78.300 ;
        RECT 78.730 77.850 79.330 78.000 ;
        RECT 70.130 77.700 74.080 77.850 ;
        RECT 75.380 77.700 79.330 77.850 ;
        RECT 70.130 77.250 70.730 77.700 ;
        RECT 78.730 77.250 79.330 77.700 ;
        RECT 70.130 77.100 74.080 77.250 ;
        RECT 75.380 77.100 79.330 77.250 ;
        RECT 70.130 76.650 70.730 77.100 ;
        RECT 78.730 76.650 79.330 77.100 ;
        RECT 70.130 76.500 74.080 76.650 ;
        RECT 75.380 76.500 79.330 76.650 ;
        RECT 70.130 76.050 70.730 76.500 ;
        RECT 78.730 76.050 79.330 76.500 ;
        RECT 70.130 75.900 74.080 76.050 ;
        RECT 75.380 75.900 79.330 76.050 ;
        RECT 70.130 75.450 70.730 75.900 ;
        RECT 78.730 75.450 79.330 75.900 ;
        RECT 70.130 75.300 74.080 75.450 ;
        RECT 75.380 75.300 79.330 75.450 ;
        RECT 70.130 74.850 70.730 75.300 ;
        RECT 78.730 74.850 79.330 75.300 ;
        RECT 70.130 74.700 74.080 74.850 ;
        RECT 75.380 74.700 79.330 74.850 ;
        RECT 70.130 74.250 70.730 74.700 ;
        RECT 78.730 74.250 79.330 74.700 ;
        RECT 70.130 74.100 74.080 74.250 ;
        RECT 75.380 74.100 79.330 74.250 ;
        RECT 70.130 73.650 70.730 74.100 ;
        RECT 78.730 73.650 79.330 74.100 ;
        RECT 70.130 73.500 74.080 73.650 ;
        RECT 75.380 73.500 79.330 73.650 ;
        RECT 70.130 73.050 70.730 73.500 ;
        RECT 78.730 73.050 79.330 73.500 ;
        RECT 70.130 72.900 74.080 73.050 ;
        RECT 75.380 72.900 79.330 73.050 ;
        RECT 70.130 72.450 70.730 72.900 ;
        RECT 78.730 72.450 79.330 72.900 ;
        RECT 70.130 72.300 74.080 72.450 ;
        RECT 75.380 72.300 79.330 72.450 ;
        RECT 70.130 71.850 70.730 72.300 ;
        RECT 78.730 71.850 79.330 72.300 ;
        RECT 70.130 71.700 74.080 71.850 ;
        RECT 75.380 71.700 79.330 71.850 ;
        RECT 70.130 71.250 70.730 71.700 ;
        RECT 78.730 71.250 79.330 71.700 ;
        RECT 70.130 71.100 74.080 71.250 ;
        RECT 75.380 71.100 79.330 71.250 ;
        RECT 70.130 70.650 70.730 71.100 ;
        RECT 78.730 70.650 79.330 71.100 ;
        RECT 70.130 70.450 74.080 70.650 ;
        RECT 75.380 70.450 79.330 70.650 ;
        RECT 79.780 70.450 79.930 78.000 ;
        RECT 80.380 70.450 80.530 78.000 ;
        RECT 80.980 70.450 81.130 78.000 ;
        RECT 81.580 70.450 81.730 78.000 ;
        RECT 82.180 70.450 82.330 78.000 ;
        RECT 82.780 75.150 82.930 78.000 ;
        RECT 83.530 75.600 85.930 78.800 ;
        RECT 89.280 78.650 90.730 78.950 ;
        RECT 86.530 78.450 90.730 78.650 ;
        RECT 98.730 78.900 104.730 79.800 ;
        RECT 98.730 78.650 100.180 78.900 ;
        RECT 100.330 78.800 104.730 78.900 ;
        RECT 98.730 78.450 102.930 78.650 ;
        RECT 86.530 78.300 94.080 78.450 ;
        RECT 95.430 78.300 102.930 78.450 ;
        RECT 86.530 78.000 90.730 78.300 ;
        RECT 86.530 75.150 86.680 78.000 ;
        RECT 87.130 70.450 87.280 78.000 ;
        RECT 87.730 70.450 87.880 78.000 ;
        RECT 88.330 70.450 88.480 78.000 ;
        RECT 88.930 70.450 89.080 78.000 ;
        RECT 89.530 70.450 89.680 78.000 ;
        RECT 90.130 77.850 90.730 78.000 ;
        RECT 98.730 78.000 102.930 78.300 ;
        RECT 98.730 77.850 99.330 78.000 ;
        RECT 90.130 77.700 94.080 77.850 ;
        RECT 95.380 77.700 99.330 77.850 ;
        RECT 90.130 77.250 90.730 77.700 ;
        RECT 98.730 77.250 99.330 77.700 ;
        RECT 90.130 77.100 94.080 77.250 ;
        RECT 95.380 77.100 99.330 77.250 ;
        RECT 90.130 76.650 90.730 77.100 ;
        RECT 98.730 76.650 99.330 77.100 ;
        RECT 90.130 76.500 94.080 76.650 ;
        RECT 95.380 76.500 99.330 76.650 ;
        RECT 90.130 76.050 90.730 76.500 ;
        RECT 98.730 76.050 99.330 76.500 ;
        RECT 90.130 75.900 94.080 76.050 ;
        RECT 95.380 75.900 99.330 76.050 ;
        RECT 90.130 75.450 90.730 75.900 ;
        RECT 98.730 75.450 99.330 75.900 ;
        RECT 90.130 75.300 94.080 75.450 ;
        RECT 95.380 75.300 99.330 75.450 ;
        RECT 90.130 74.850 90.730 75.300 ;
        RECT 98.730 74.850 99.330 75.300 ;
        RECT 90.130 74.700 94.080 74.850 ;
        RECT 95.380 74.700 99.330 74.850 ;
        RECT 90.130 74.250 90.730 74.700 ;
        RECT 98.730 74.250 99.330 74.700 ;
        RECT 90.130 74.100 94.080 74.250 ;
        RECT 95.380 74.100 99.330 74.250 ;
        RECT 90.130 73.650 90.730 74.100 ;
        RECT 98.730 73.650 99.330 74.100 ;
        RECT 90.130 73.500 94.080 73.650 ;
        RECT 95.380 73.500 99.330 73.650 ;
        RECT 90.130 73.050 90.730 73.500 ;
        RECT 98.730 73.050 99.330 73.500 ;
        RECT 90.130 72.900 94.080 73.050 ;
        RECT 95.380 72.900 99.330 73.050 ;
        RECT 90.130 72.450 90.730 72.900 ;
        RECT 98.730 72.450 99.330 72.900 ;
        RECT 90.130 72.300 94.080 72.450 ;
        RECT 95.380 72.300 99.330 72.450 ;
        RECT 90.130 71.850 90.730 72.300 ;
        RECT 98.730 71.850 99.330 72.300 ;
        RECT 90.130 71.700 94.080 71.850 ;
        RECT 95.380 71.700 99.330 71.850 ;
        RECT 90.130 71.250 90.730 71.700 ;
        RECT 98.730 71.250 99.330 71.700 ;
        RECT 90.130 71.100 94.080 71.250 ;
        RECT 95.380 71.100 99.330 71.250 ;
        RECT 90.130 70.650 90.730 71.100 ;
        RECT 98.730 70.650 99.330 71.100 ;
        RECT 90.130 70.450 94.080 70.650 ;
        RECT 95.380 70.450 99.330 70.650 ;
        RECT 99.780 70.450 99.930 78.000 ;
        RECT 100.380 70.450 100.530 78.000 ;
        RECT 100.980 70.450 101.130 78.000 ;
        RECT 101.580 70.450 101.730 78.000 ;
        RECT 102.180 70.450 102.330 78.000 ;
        RECT 102.780 75.150 102.930 78.000 ;
        RECT 103.530 77.310 104.730 78.800 ;
        RECT 103.530 76.035 107.135 77.310 ;
        RECT 103.530 75.600 104.730 76.035 ;
        RECT 2.315 64.450 4.315 66.745 ;
        RECT 4.730 63.230 5.930 64.400 ;
        RECT 2.315 61.955 5.930 63.230 ;
        RECT 4.730 61.200 5.930 61.955 ;
        RECT 6.530 62.000 6.680 64.900 ;
        RECT 7.130 62.000 7.280 69.550 ;
        RECT 7.730 62.000 7.880 69.550 ;
        RECT 8.330 62.000 8.480 69.550 ;
        RECT 8.930 62.000 9.080 69.550 ;
        RECT 9.530 62.000 9.680 69.550 ;
        RECT 10.130 69.350 14.080 69.550 ;
        RECT 15.380 69.350 19.330 69.550 ;
        RECT 10.130 68.900 10.730 69.350 ;
        RECT 18.730 68.900 19.330 69.350 ;
        RECT 10.130 68.750 14.080 68.900 ;
        RECT 15.380 68.750 19.330 68.900 ;
        RECT 10.130 68.300 10.730 68.750 ;
        RECT 18.730 68.300 19.330 68.750 ;
        RECT 10.130 68.150 14.080 68.300 ;
        RECT 15.380 68.150 19.330 68.300 ;
        RECT 10.130 67.700 10.730 68.150 ;
        RECT 18.730 67.700 19.330 68.150 ;
        RECT 10.130 67.550 14.080 67.700 ;
        RECT 15.380 67.550 19.330 67.700 ;
        RECT 10.130 67.100 10.730 67.550 ;
        RECT 18.730 67.100 19.330 67.550 ;
        RECT 10.130 66.950 14.080 67.100 ;
        RECT 15.380 66.950 19.330 67.100 ;
        RECT 10.130 66.500 10.730 66.950 ;
        RECT 18.730 66.500 19.330 66.950 ;
        RECT 10.130 66.350 14.080 66.500 ;
        RECT 15.380 66.350 19.330 66.500 ;
        RECT 10.130 65.900 10.730 66.350 ;
        RECT 18.730 65.900 19.330 66.350 ;
        RECT 10.130 65.750 14.080 65.900 ;
        RECT 15.380 65.750 19.330 65.900 ;
        RECT 10.130 65.300 10.730 65.750 ;
        RECT 18.730 65.300 19.330 65.750 ;
        RECT 10.130 65.150 14.080 65.300 ;
        RECT 15.380 65.150 19.330 65.300 ;
        RECT 10.130 64.700 10.730 65.150 ;
        RECT 18.730 64.700 19.330 65.150 ;
        RECT 10.130 64.550 14.080 64.700 ;
        RECT 15.380 64.550 19.330 64.700 ;
        RECT 10.130 64.100 10.730 64.550 ;
        RECT 18.730 64.100 19.330 64.550 ;
        RECT 10.130 63.950 14.080 64.100 ;
        RECT 15.380 63.950 19.330 64.100 ;
        RECT 10.130 63.500 10.730 63.950 ;
        RECT 18.730 63.500 19.330 63.950 ;
        RECT 10.130 63.350 14.080 63.500 ;
        RECT 15.380 63.350 19.330 63.500 ;
        RECT 10.130 62.900 10.730 63.350 ;
        RECT 18.730 62.900 19.330 63.350 ;
        RECT 10.130 62.750 14.080 62.900 ;
        RECT 15.380 62.750 19.330 62.900 ;
        RECT 10.130 62.300 10.730 62.750 ;
        RECT 18.730 62.300 19.330 62.750 ;
        RECT 10.130 62.150 14.080 62.300 ;
        RECT 15.380 62.150 19.330 62.300 ;
        RECT 10.130 62.000 10.730 62.150 ;
        RECT 6.530 61.700 10.730 62.000 ;
        RECT 18.730 62.000 19.330 62.150 ;
        RECT 19.780 62.000 19.930 69.550 ;
        RECT 20.380 62.000 20.530 69.550 ;
        RECT 20.980 62.000 21.130 69.550 ;
        RECT 21.580 62.000 21.730 69.550 ;
        RECT 22.180 62.000 22.330 69.550 ;
        RECT 22.780 62.000 22.930 64.900 ;
        RECT 18.730 61.700 22.930 62.000 ;
        RECT 6.530 61.550 14.080 61.700 ;
        RECT 15.380 61.550 22.930 61.700 ;
        RECT 6.530 61.350 10.730 61.550 ;
        RECT 4.730 61.050 9.130 61.200 ;
        RECT 9.280 61.050 10.730 61.350 ;
        RECT 4.730 60.150 10.730 61.050 ;
        RECT 18.730 61.350 22.930 61.550 ;
        RECT 18.730 61.050 20.180 61.350 ;
        RECT 23.530 61.200 25.930 64.400 ;
        RECT 26.530 62.000 26.680 64.900 ;
        RECT 27.130 62.000 27.280 69.550 ;
        RECT 27.730 62.000 27.880 69.550 ;
        RECT 28.330 62.000 28.480 69.550 ;
        RECT 28.930 62.000 29.080 69.550 ;
        RECT 29.530 62.000 29.680 69.550 ;
        RECT 30.130 69.350 34.080 69.550 ;
        RECT 35.380 69.350 39.330 69.550 ;
        RECT 30.130 68.900 30.730 69.350 ;
        RECT 38.730 68.900 39.330 69.350 ;
        RECT 30.130 68.750 34.080 68.900 ;
        RECT 35.380 68.750 39.330 68.900 ;
        RECT 30.130 68.300 30.730 68.750 ;
        RECT 38.730 68.300 39.330 68.750 ;
        RECT 30.130 68.150 34.080 68.300 ;
        RECT 35.380 68.150 39.330 68.300 ;
        RECT 30.130 67.700 30.730 68.150 ;
        RECT 38.730 67.700 39.330 68.150 ;
        RECT 30.130 67.550 34.080 67.700 ;
        RECT 35.380 67.550 39.330 67.700 ;
        RECT 30.130 67.100 30.730 67.550 ;
        RECT 38.730 67.100 39.330 67.550 ;
        RECT 30.130 66.950 34.080 67.100 ;
        RECT 35.380 66.950 39.330 67.100 ;
        RECT 30.130 66.500 30.730 66.950 ;
        RECT 38.730 66.500 39.330 66.950 ;
        RECT 30.130 66.350 34.080 66.500 ;
        RECT 35.380 66.350 39.330 66.500 ;
        RECT 30.130 65.900 30.730 66.350 ;
        RECT 38.730 65.900 39.330 66.350 ;
        RECT 30.130 65.750 34.080 65.900 ;
        RECT 35.380 65.750 39.330 65.900 ;
        RECT 30.130 65.300 30.730 65.750 ;
        RECT 38.730 65.300 39.330 65.750 ;
        RECT 30.130 65.150 34.080 65.300 ;
        RECT 35.380 65.150 39.330 65.300 ;
        RECT 30.130 64.700 30.730 65.150 ;
        RECT 38.730 64.700 39.330 65.150 ;
        RECT 30.130 64.550 34.080 64.700 ;
        RECT 35.380 64.550 39.330 64.700 ;
        RECT 30.130 64.100 30.730 64.550 ;
        RECT 38.730 64.100 39.330 64.550 ;
        RECT 30.130 63.950 34.080 64.100 ;
        RECT 35.380 63.950 39.330 64.100 ;
        RECT 30.130 63.500 30.730 63.950 ;
        RECT 38.730 63.500 39.330 63.950 ;
        RECT 30.130 63.350 34.080 63.500 ;
        RECT 35.380 63.350 39.330 63.500 ;
        RECT 30.130 62.900 30.730 63.350 ;
        RECT 38.730 62.900 39.330 63.350 ;
        RECT 30.130 62.750 34.080 62.900 ;
        RECT 35.380 62.750 39.330 62.900 ;
        RECT 30.130 62.300 30.730 62.750 ;
        RECT 38.730 62.300 39.330 62.750 ;
        RECT 30.130 62.150 34.080 62.300 ;
        RECT 35.380 62.150 39.330 62.300 ;
        RECT 30.130 62.000 30.730 62.150 ;
        RECT 26.530 61.700 30.730 62.000 ;
        RECT 38.730 62.000 39.330 62.150 ;
        RECT 39.780 62.000 39.930 69.550 ;
        RECT 40.380 62.000 40.530 69.550 ;
        RECT 40.980 62.000 41.130 69.550 ;
        RECT 41.580 62.000 41.730 69.550 ;
        RECT 42.180 62.000 42.330 69.550 ;
        RECT 42.780 62.000 42.930 64.900 ;
        RECT 38.730 61.700 42.930 62.000 ;
        RECT 26.530 61.550 34.080 61.700 ;
        RECT 35.380 61.550 42.930 61.700 ;
        RECT 26.530 61.350 30.730 61.550 ;
        RECT 20.330 61.050 29.130 61.200 ;
        RECT 29.280 61.050 30.730 61.350 ;
        RECT 18.730 60.150 30.730 61.050 ;
        RECT 38.730 61.350 42.930 61.550 ;
        RECT 38.730 61.050 40.180 61.350 ;
        RECT 43.530 61.200 45.930 64.400 ;
        RECT 46.530 62.000 46.680 64.900 ;
        RECT 47.130 62.000 47.280 69.550 ;
        RECT 47.730 62.000 47.880 69.550 ;
        RECT 48.330 62.000 48.480 69.550 ;
        RECT 48.930 62.000 49.080 69.550 ;
        RECT 49.530 62.000 49.680 69.550 ;
        RECT 50.130 69.350 54.080 69.550 ;
        RECT 55.380 69.350 59.330 69.550 ;
        RECT 50.130 68.900 50.730 69.350 ;
        RECT 58.730 68.900 59.330 69.350 ;
        RECT 50.130 68.750 54.080 68.900 ;
        RECT 55.380 68.750 59.330 68.900 ;
        RECT 50.130 68.300 50.730 68.750 ;
        RECT 58.730 68.300 59.330 68.750 ;
        RECT 50.130 68.150 54.080 68.300 ;
        RECT 55.380 68.150 59.330 68.300 ;
        RECT 50.130 67.700 50.730 68.150 ;
        RECT 58.730 67.700 59.330 68.150 ;
        RECT 50.130 67.550 54.080 67.700 ;
        RECT 55.380 67.550 59.330 67.700 ;
        RECT 50.130 67.100 50.730 67.550 ;
        RECT 58.730 67.100 59.330 67.550 ;
        RECT 50.130 66.950 54.080 67.100 ;
        RECT 55.380 66.950 59.330 67.100 ;
        RECT 50.130 66.500 50.730 66.950 ;
        RECT 58.730 66.500 59.330 66.950 ;
        RECT 50.130 66.350 54.080 66.500 ;
        RECT 55.380 66.350 59.330 66.500 ;
        RECT 50.130 65.900 50.730 66.350 ;
        RECT 58.730 65.900 59.330 66.350 ;
        RECT 50.130 65.750 54.080 65.900 ;
        RECT 55.380 65.750 59.330 65.900 ;
        RECT 50.130 65.300 50.730 65.750 ;
        RECT 58.730 65.300 59.330 65.750 ;
        RECT 50.130 65.150 54.080 65.300 ;
        RECT 55.380 65.150 59.330 65.300 ;
        RECT 50.130 64.700 50.730 65.150 ;
        RECT 58.730 64.700 59.330 65.150 ;
        RECT 50.130 64.550 54.080 64.700 ;
        RECT 55.380 64.550 59.330 64.700 ;
        RECT 50.130 64.100 50.730 64.550 ;
        RECT 58.730 64.100 59.330 64.550 ;
        RECT 50.130 63.950 54.080 64.100 ;
        RECT 55.380 63.950 59.330 64.100 ;
        RECT 50.130 63.500 50.730 63.950 ;
        RECT 58.730 63.500 59.330 63.950 ;
        RECT 50.130 63.350 54.080 63.500 ;
        RECT 55.380 63.350 59.330 63.500 ;
        RECT 50.130 62.900 50.730 63.350 ;
        RECT 58.730 62.900 59.330 63.350 ;
        RECT 50.130 62.750 54.080 62.900 ;
        RECT 55.380 62.750 59.330 62.900 ;
        RECT 50.130 62.300 50.730 62.750 ;
        RECT 58.730 62.300 59.330 62.750 ;
        RECT 50.130 62.150 54.080 62.300 ;
        RECT 55.380 62.150 59.330 62.300 ;
        RECT 50.130 62.000 50.730 62.150 ;
        RECT 46.530 61.700 50.730 62.000 ;
        RECT 58.730 62.000 59.330 62.150 ;
        RECT 59.780 62.000 59.930 69.550 ;
        RECT 60.380 62.000 60.530 69.550 ;
        RECT 60.980 62.000 61.130 69.550 ;
        RECT 61.580 62.000 61.730 69.550 ;
        RECT 62.180 62.000 62.330 69.550 ;
        RECT 62.780 62.000 62.930 64.900 ;
        RECT 58.730 61.700 62.930 62.000 ;
        RECT 46.530 61.550 54.080 61.700 ;
        RECT 55.380 61.550 62.930 61.700 ;
        RECT 46.530 61.350 50.730 61.550 ;
        RECT 40.330 61.050 49.130 61.200 ;
        RECT 49.280 61.050 50.730 61.350 ;
        RECT 38.730 60.150 50.730 61.050 ;
        RECT 58.730 61.350 62.930 61.550 ;
        RECT 58.730 61.050 60.180 61.350 ;
        RECT 63.530 61.200 65.930 64.400 ;
        RECT 66.530 62.000 66.680 64.900 ;
        RECT 67.130 62.000 67.280 69.550 ;
        RECT 67.730 62.000 67.880 69.550 ;
        RECT 68.330 62.000 68.480 69.550 ;
        RECT 68.930 62.000 69.080 69.550 ;
        RECT 69.530 62.000 69.680 69.550 ;
        RECT 70.130 69.350 74.080 69.550 ;
        RECT 75.380 69.350 79.330 69.550 ;
        RECT 70.130 68.900 70.730 69.350 ;
        RECT 78.730 68.900 79.330 69.350 ;
        RECT 70.130 68.750 74.080 68.900 ;
        RECT 75.380 68.750 79.330 68.900 ;
        RECT 70.130 68.300 70.730 68.750 ;
        RECT 78.730 68.300 79.330 68.750 ;
        RECT 70.130 68.150 74.080 68.300 ;
        RECT 75.380 68.150 79.330 68.300 ;
        RECT 70.130 67.700 70.730 68.150 ;
        RECT 78.730 67.700 79.330 68.150 ;
        RECT 70.130 67.550 74.080 67.700 ;
        RECT 75.380 67.550 79.330 67.700 ;
        RECT 70.130 67.100 70.730 67.550 ;
        RECT 78.730 67.100 79.330 67.550 ;
        RECT 70.130 66.950 74.080 67.100 ;
        RECT 75.380 66.950 79.330 67.100 ;
        RECT 70.130 66.500 70.730 66.950 ;
        RECT 78.730 66.500 79.330 66.950 ;
        RECT 70.130 66.350 74.080 66.500 ;
        RECT 75.380 66.350 79.330 66.500 ;
        RECT 70.130 65.900 70.730 66.350 ;
        RECT 78.730 65.900 79.330 66.350 ;
        RECT 70.130 65.750 74.080 65.900 ;
        RECT 75.380 65.750 79.330 65.900 ;
        RECT 70.130 65.300 70.730 65.750 ;
        RECT 78.730 65.300 79.330 65.750 ;
        RECT 70.130 65.150 74.080 65.300 ;
        RECT 75.380 65.150 79.330 65.300 ;
        RECT 70.130 64.700 70.730 65.150 ;
        RECT 78.730 64.700 79.330 65.150 ;
        RECT 70.130 64.550 74.080 64.700 ;
        RECT 75.380 64.550 79.330 64.700 ;
        RECT 70.130 64.100 70.730 64.550 ;
        RECT 78.730 64.100 79.330 64.550 ;
        RECT 70.130 63.950 74.080 64.100 ;
        RECT 75.380 63.950 79.330 64.100 ;
        RECT 70.130 63.500 70.730 63.950 ;
        RECT 78.730 63.500 79.330 63.950 ;
        RECT 70.130 63.350 74.080 63.500 ;
        RECT 75.380 63.350 79.330 63.500 ;
        RECT 70.130 62.900 70.730 63.350 ;
        RECT 78.730 62.900 79.330 63.350 ;
        RECT 70.130 62.750 74.080 62.900 ;
        RECT 75.380 62.750 79.330 62.900 ;
        RECT 70.130 62.300 70.730 62.750 ;
        RECT 78.730 62.300 79.330 62.750 ;
        RECT 70.130 62.150 74.080 62.300 ;
        RECT 75.380 62.150 79.330 62.300 ;
        RECT 70.130 62.000 70.730 62.150 ;
        RECT 66.530 61.700 70.730 62.000 ;
        RECT 78.730 62.000 79.330 62.150 ;
        RECT 79.780 62.000 79.930 69.550 ;
        RECT 80.380 62.000 80.530 69.550 ;
        RECT 80.980 62.000 81.130 69.550 ;
        RECT 81.580 62.000 81.730 69.550 ;
        RECT 82.180 62.000 82.330 69.550 ;
        RECT 82.780 62.000 82.930 64.900 ;
        RECT 78.730 61.700 82.930 62.000 ;
        RECT 66.530 61.550 74.080 61.700 ;
        RECT 75.380 61.550 82.930 61.700 ;
        RECT 66.530 61.350 70.730 61.550 ;
        RECT 60.330 61.050 69.130 61.200 ;
        RECT 69.280 61.050 70.730 61.350 ;
        RECT 58.730 60.150 70.730 61.050 ;
        RECT 78.730 61.350 82.930 61.550 ;
        RECT 78.730 61.050 80.180 61.350 ;
        RECT 83.530 61.200 85.930 64.400 ;
        RECT 86.530 62.000 86.680 64.900 ;
        RECT 87.130 62.000 87.280 69.550 ;
        RECT 87.730 62.000 87.880 69.550 ;
        RECT 88.330 62.000 88.480 69.550 ;
        RECT 88.930 62.000 89.080 69.550 ;
        RECT 89.530 62.000 89.680 69.550 ;
        RECT 90.130 69.350 94.080 69.550 ;
        RECT 95.380 69.350 99.330 69.550 ;
        RECT 90.130 68.900 90.730 69.350 ;
        RECT 98.730 68.900 99.330 69.350 ;
        RECT 90.130 68.750 94.080 68.900 ;
        RECT 95.380 68.750 99.330 68.900 ;
        RECT 90.130 68.300 90.730 68.750 ;
        RECT 98.730 68.300 99.330 68.750 ;
        RECT 90.130 68.150 94.080 68.300 ;
        RECT 95.380 68.150 99.330 68.300 ;
        RECT 90.130 67.700 90.730 68.150 ;
        RECT 98.730 67.700 99.330 68.150 ;
        RECT 90.130 67.550 94.080 67.700 ;
        RECT 95.380 67.550 99.330 67.700 ;
        RECT 90.130 67.100 90.730 67.550 ;
        RECT 98.730 67.100 99.330 67.550 ;
        RECT 90.130 66.950 94.080 67.100 ;
        RECT 95.380 66.950 99.330 67.100 ;
        RECT 90.130 66.500 90.730 66.950 ;
        RECT 98.730 66.500 99.330 66.950 ;
        RECT 90.130 66.350 94.080 66.500 ;
        RECT 95.380 66.350 99.330 66.500 ;
        RECT 90.130 65.900 90.730 66.350 ;
        RECT 98.730 65.900 99.330 66.350 ;
        RECT 90.130 65.750 94.080 65.900 ;
        RECT 95.380 65.750 99.330 65.900 ;
        RECT 90.130 65.300 90.730 65.750 ;
        RECT 98.730 65.300 99.330 65.750 ;
        RECT 90.130 65.150 94.080 65.300 ;
        RECT 95.380 65.150 99.330 65.300 ;
        RECT 90.130 64.700 90.730 65.150 ;
        RECT 98.730 64.700 99.330 65.150 ;
        RECT 90.130 64.550 94.080 64.700 ;
        RECT 95.380 64.550 99.330 64.700 ;
        RECT 90.130 64.100 90.730 64.550 ;
        RECT 98.730 64.100 99.330 64.550 ;
        RECT 90.130 63.950 94.080 64.100 ;
        RECT 95.380 63.950 99.330 64.100 ;
        RECT 90.130 63.500 90.730 63.950 ;
        RECT 98.730 63.500 99.330 63.950 ;
        RECT 90.130 63.350 94.080 63.500 ;
        RECT 95.380 63.350 99.330 63.500 ;
        RECT 90.130 62.900 90.730 63.350 ;
        RECT 98.730 62.900 99.330 63.350 ;
        RECT 90.130 62.750 94.080 62.900 ;
        RECT 95.380 62.750 99.330 62.900 ;
        RECT 90.130 62.300 90.730 62.750 ;
        RECT 98.730 62.300 99.330 62.750 ;
        RECT 90.130 62.150 94.080 62.300 ;
        RECT 95.380 62.150 99.330 62.300 ;
        RECT 90.130 62.000 90.730 62.150 ;
        RECT 86.530 61.700 90.730 62.000 ;
        RECT 98.730 62.000 99.330 62.150 ;
        RECT 99.780 62.000 99.930 69.550 ;
        RECT 100.380 62.000 100.530 69.550 ;
        RECT 100.980 62.000 101.130 69.550 ;
        RECT 101.580 62.000 101.730 69.550 ;
        RECT 102.180 62.000 102.330 69.550 ;
        RECT 102.780 62.000 102.930 64.900 ;
        RECT 98.730 61.700 102.930 62.000 ;
        RECT 86.530 61.550 94.080 61.700 ;
        RECT 95.380 61.550 102.930 61.700 ;
        RECT 86.530 61.350 90.730 61.550 ;
        RECT 80.330 61.050 89.130 61.200 ;
        RECT 89.280 61.050 90.730 61.350 ;
        RECT 78.730 60.150 90.730 61.050 ;
        RECT 98.730 61.350 102.930 61.550 ;
        RECT 103.530 63.095 104.730 64.400 ;
        RECT 103.530 61.820 107.140 63.095 ;
        RECT 98.730 61.050 100.180 61.350 ;
        RECT 103.530 61.200 104.730 61.820 ;
        RECT 100.330 61.050 104.730 61.200 ;
        RECT 98.730 60.150 104.730 61.050 ;
        RECT 4.730 59.850 9.130 60.150 ;
        RECT 20.330 59.850 29.130 60.150 ;
        RECT 40.330 59.850 49.130 60.150 ;
        RECT 60.330 59.850 69.130 60.150 ;
        RECT 80.330 59.850 89.130 60.150 ;
        RECT 4.730 58.950 10.730 59.850 ;
        RECT 20.330 59.800 30.730 59.850 ;
        RECT 40.330 59.800 50.730 59.850 ;
        RECT 60.330 59.800 70.730 59.850 ;
        RECT 80.330 59.800 90.730 59.850 ;
        RECT 100.330 59.800 104.730 60.150 ;
        RECT 4.730 58.800 9.130 58.950 ;
        RECT 4.730 57.620 5.930 58.800 ;
        RECT 9.280 58.650 10.730 58.950 ;
        RECT 2.315 56.345 5.930 57.620 ;
        RECT 4.730 55.600 5.930 56.345 ;
        RECT 6.530 58.450 10.730 58.650 ;
        RECT 18.730 58.950 30.730 59.800 ;
        RECT 18.730 58.900 29.130 58.950 ;
        RECT 18.730 58.650 20.180 58.900 ;
        RECT 20.330 58.800 29.130 58.900 ;
        RECT 18.730 58.450 22.930 58.650 ;
        RECT 6.530 58.300 14.080 58.450 ;
        RECT 15.430 58.300 22.930 58.450 ;
        RECT 6.530 58.000 10.730 58.300 ;
        RECT 2.315 53.255 4.315 55.550 ;
        RECT 6.530 55.150 6.680 58.000 ;
        RECT 7.130 50.450 7.280 58.000 ;
        RECT 7.730 50.450 7.880 58.000 ;
        RECT 8.330 50.450 8.480 58.000 ;
        RECT 8.930 50.450 9.080 58.000 ;
        RECT 9.530 50.450 9.680 58.000 ;
        RECT 10.130 57.850 10.730 58.000 ;
        RECT 18.730 58.000 22.930 58.300 ;
        RECT 18.730 57.850 19.330 58.000 ;
        RECT 10.130 57.700 14.080 57.850 ;
        RECT 15.380 57.700 19.330 57.850 ;
        RECT 10.130 57.250 10.730 57.700 ;
        RECT 18.730 57.250 19.330 57.700 ;
        RECT 10.130 57.100 14.080 57.250 ;
        RECT 15.380 57.100 19.330 57.250 ;
        RECT 10.130 56.650 10.730 57.100 ;
        RECT 18.730 56.650 19.330 57.100 ;
        RECT 10.130 56.500 14.080 56.650 ;
        RECT 15.380 56.500 19.330 56.650 ;
        RECT 10.130 56.050 10.730 56.500 ;
        RECT 18.730 56.050 19.330 56.500 ;
        RECT 10.130 55.900 14.080 56.050 ;
        RECT 15.380 55.900 19.330 56.050 ;
        RECT 10.130 55.450 10.730 55.900 ;
        RECT 18.730 55.450 19.330 55.900 ;
        RECT 10.130 55.300 14.080 55.450 ;
        RECT 15.380 55.300 19.330 55.450 ;
        RECT 10.130 54.850 10.730 55.300 ;
        RECT 18.730 54.850 19.330 55.300 ;
        RECT 10.130 54.700 14.080 54.850 ;
        RECT 15.380 54.700 19.330 54.850 ;
        RECT 10.130 54.250 10.730 54.700 ;
        RECT 18.730 54.250 19.330 54.700 ;
        RECT 10.130 54.100 14.080 54.250 ;
        RECT 15.380 54.100 19.330 54.250 ;
        RECT 10.130 53.650 10.730 54.100 ;
        RECT 18.730 53.650 19.330 54.100 ;
        RECT 10.130 53.500 14.080 53.650 ;
        RECT 15.380 53.500 19.330 53.650 ;
        RECT 10.130 53.050 10.730 53.500 ;
        RECT 18.730 53.050 19.330 53.500 ;
        RECT 10.130 52.900 14.080 53.050 ;
        RECT 15.380 52.900 19.330 53.050 ;
        RECT 10.130 52.450 10.730 52.900 ;
        RECT 18.730 52.450 19.330 52.900 ;
        RECT 10.130 52.300 14.080 52.450 ;
        RECT 15.380 52.300 19.330 52.450 ;
        RECT 10.130 51.850 10.730 52.300 ;
        RECT 18.730 51.850 19.330 52.300 ;
        RECT 10.130 51.700 14.080 51.850 ;
        RECT 15.380 51.700 19.330 51.850 ;
        RECT 10.130 51.250 10.730 51.700 ;
        RECT 18.730 51.250 19.330 51.700 ;
        RECT 10.130 51.100 14.080 51.250 ;
        RECT 15.380 51.100 19.330 51.250 ;
        RECT 10.130 50.650 10.730 51.100 ;
        RECT 18.730 50.650 19.330 51.100 ;
        RECT 10.130 50.450 14.080 50.650 ;
        RECT 15.380 50.450 19.330 50.650 ;
        RECT 19.780 50.450 19.930 58.000 ;
        RECT 20.380 50.450 20.530 58.000 ;
        RECT 20.980 50.450 21.130 58.000 ;
        RECT 21.580 50.450 21.730 58.000 ;
        RECT 22.180 50.450 22.330 58.000 ;
        RECT 22.780 55.150 22.930 58.000 ;
        RECT 23.530 55.600 25.930 58.800 ;
        RECT 29.280 58.650 30.730 58.950 ;
        RECT 26.530 58.450 30.730 58.650 ;
        RECT 38.730 58.950 50.730 59.800 ;
        RECT 38.730 58.900 49.130 58.950 ;
        RECT 38.730 58.650 40.180 58.900 ;
        RECT 40.330 58.800 49.130 58.900 ;
        RECT 38.730 58.450 42.930 58.650 ;
        RECT 26.530 58.300 34.080 58.450 ;
        RECT 35.430 58.300 42.930 58.450 ;
        RECT 26.530 58.000 30.730 58.300 ;
        RECT 26.530 55.150 26.680 58.000 ;
        RECT 27.130 50.450 27.280 58.000 ;
        RECT 27.730 50.450 27.880 58.000 ;
        RECT 28.330 50.450 28.480 58.000 ;
        RECT 28.930 50.450 29.080 58.000 ;
        RECT 29.530 50.450 29.680 58.000 ;
        RECT 30.130 57.850 30.730 58.000 ;
        RECT 38.730 58.000 42.930 58.300 ;
        RECT 38.730 57.850 39.330 58.000 ;
        RECT 30.130 57.700 34.080 57.850 ;
        RECT 35.380 57.700 39.330 57.850 ;
        RECT 30.130 57.250 30.730 57.700 ;
        RECT 38.730 57.250 39.330 57.700 ;
        RECT 30.130 57.100 34.080 57.250 ;
        RECT 35.380 57.100 39.330 57.250 ;
        RECT 30.130 56.650 30.730 57.100 ;
        RECT 38.730 56.650 39.330 57.100 ;
        RECT 30.130 56.500 34.080 56.650 ;
        RECT 35.380 56.500 39.330 56.650 ;
        RECT 30.130 56.050 30.730 56.500 ;
        RECT 38.730 56.050 39.330 56.500 ;
        RECT 30.130 55.900 34.080 56.050 ;
        RECT 35.380 55.900 39.330 56.050 ;
        RECT 30.130 55.450 30.730 55.900 ;
        RECT 38.730 55.450 39.330 55.900 ;
        RECT 30.130 55.300 34.080 55.450 ;
        RECT 35.380 55.300 39.330 55.450 ;
        RECT 30.130 54.850 30.730 55.300 ;
        RECT 38.730 54.850 39.330 55.300 ;
        RECT 30.130 54.700 34.080 54.850 ;
        RECT 35.380 54.700 39.330 54.850 ;
        RECT 30.130 54.250 30.730 54.700 ;
        RECT 38.730 54.250 39.330 54.700 ;
        RECT 30.130 54.100 34.080 54.250 ;
        RECT 35.380 54.100 39.330 54.250 ;
        RECT 30.130 53.650 30.730 54.100 ;
        RECT 38.730 53.650 39.330 54.100 ;
        RECT 30.130 53.500 34.080 53.650 ;
        RECT 35.380 53.500 39.330 53.650 ;
        RECT 30.130 53.050 30.730 53.500 ;
        RECT 38.730 53.050 39.330 53.500 ;
        RECT 30.130 52.900 34.080 53.050 ;
        RECT 35.380 52.900 39.330 53.050 ;
        RECT 30.130 52.450 30.730 52.900 ;
        RECT 38.730 52.450 39.330 52.900 ;
        RECT 30.130 52.300 34.080 52.450 ;
        RECT 35.380 52.300 39.330 52.450 ;
        RECT 30.130 51.850 30.730 52.300 ;
        RECT 38.730 51.850 39.330 52.300 ;
        RECT 30.130 51.700 34.080 51.850 ;
        RECT 35.380 51.700 39.330 51.850 ;
        RECT 30.130 51.250 30.730 51.700 ;
        RECT 38.730 51.250 39.330 51.700 ;
        RECT 30.130 51.100 34.080 51.250 ;
        RECT 35.380 51.100 39.330 51.250 ;
        RECT 30.130 50.650 30.730 51.100 ;
        RECT 38.730 50.650 39.330 51.100 ;
        RECT 30.130 50.450 34.080 50.650 ;
        RECT 35.380 50.450 39.330 50.650 ;
        RECT 39.780 50.450 39.930 58.000 ;
        RECT 40.380 50.450 40.530 58.000 ;
        RECT 40.980 50.450 41.130 58.000 ;
        RECT 41.580 50.450 41.730 58.000 ;
        RECT 42.180 50.450 42.330 58.000 ;
        RECT 42.780 55.150 42.930 58.000 ;
        RECT 43.530 55.600 45.930 58.800 ;
        RECT 49.280 58.650 50.730 58.950 ;
        RECT 46.530 58.450 50.730 58.650 ;
        RECT 58.730 58.950 70.730 59.800 ;
        RECT 58.730 58.900 69.130 58.950 ;
        RECT 58.730 58.650 60.180 58.900 ;
        RECT 60.330 58.800 69.130 58.900 ;
        RECT 58.730 58.450 62.930 58.650 ;
        RECT 46.530 58.300 54.080 58.450 ;
        RECT 55.430 58.300 62.930 58.450 ;
        RECT 46.530 58.000 50.730 58.300 ;
        RECT 46.530 55.150 46.680 58.000 ;
        RECT 47.130 50.450 47.280 58.000 ;
        RECT 47.730 50.450 47.880 58.000 ;
        RECT 48.330 50.450 48.480 58.000 ;
        RECT 48.930 50.450 49.080 58.000 ;
        RECT 49.530 50.450 49.680 58.000 ;
        RECT 50.130 57.850 50.730 58.000 ;
        RECT 58.730 58.000 62.930 58.300 ;
        RECT 58.730 57.850 59.330 58.000 ;
        RECT 50.130 57.700 54.080 57.850 ;
        RECT 55.380 57.700 59.330 57.850 ;
        RECT 50.130 57.250 50.730 57.700 ;
        RECT 58.730 57.250 59.330 57.700 ;
        RECT 50.130 57.100 54.080 57.250 ;
        RECT 55.380 57.100 59.330 57.250 ;
        RECT 50.130 56.650 50.730 57.100 ;
        RECT 58.730 56.650 59.330 57.100 ;
        RECT 50.130 56.500 54.080 56.650 ;
        RECT 55.380 56.500 59.330 56.650 ;
        RECT 50.130 56.050 50.730 56.500 ;
        RECT 58.730 56.050 59.330 56.500 ;
        RECT 50.130 55.900 54.080 56.050 ;
        RECT 55.380 55.900 59.330 56.050 ;
        RECT 50.130 55.450 50.730 55.900 ;
        RECT 58.730 55.450 59.330 55.900 ;
        RECT 50.130 55.300 54.080 55.450 ;
        RECT 55.380 55.300 59.330 55.450 ;
        RECT 50.130 54.850 50.730 55.300 ;
        RECT 58.730 54.850 59.330 55.300 ;
        RECT 50.130 54.700 54.080 54.850 ;
        RECT 55.380 54.700 59.330 54.850 ;
        RECT 50.130 54.250 50.730 54.700 ;
        RECT 58.730 54.250 59.330 54.700 ;
        RECT 50.130 54.100 54.080 54.250 ;
        RECT 55.380 54.100 59.330 54.250 ;
        RECT 50.130 53.650 50.730 54.100 ;
        RECT 58.730 53.650 59.330 54.100 ;
        RECT 50.130 53.500 54.080 53.650 ;
        RECT 55.380 53.500 59.330 53.650 ;
        RECT 50.130 53.050 50.730 53.500 ;
        RECT 58.730 53.050 59.330 53.500 ;
        RECT 50.130 52.900 54.080 53.050 ;
        RECT 55.380 52.900 59.330 53.050 ;
        RECT 50.130 52.450 50.730 52.900 ;
        RECT 58.730 52.450 59.330 52.900 ;
        RECT 50.130 52.300 54.080 52.450 ;
        RECT 55.380 52.300 59.330 52.450 ;
        RECT 50.130 51.850 50.730 52.300 ;
        RECT 58.730 51.850 59.330 52.300 ;
        RECT 50.130 51.700 54.080 51.850 ;
        RECT 55.380 51.700 59.330 51.850 ;
        RECT 50.130 51.250 50.730 51.700 ;
        RECT 58.730 51.250 59.330 51.700 ;
        RECT 50.130 51.100 54.080 51.250 ;
        RECT 55.380 51.100 59.330 51.250 ;
        RECT 50.130 50.650 50.730 51.100 ;
        RECT 58.730 50.650 59.330 51.100 ;
        RECT 50.130 50.450 54.080 50.650 ;
        RECT 55.380 50.450 59.330 50.650 ;
        RECT 59.780 50.450 59.930 58.000 ;
        RECT 60.380 50.450 60.530 58.000 ;
        RECT 60.980 50.450 61.130 58.000 ;
        RECT 61.580 50.450 61.730 58.000 ;
        RECT 62.180 50.450 62.330 58.000 ;
        RECT 62.780 55.150 62.930 58.000 ;
        RECT 63.530 55.600 65.930 58.800 ;
        RECT 69.280 58.650 70.730 58.950 ;
        RECT 66.530 58.450 70.730 58.650 ;
        RECT 78.730 58.950 90.730 59.800 ;
        RECT 78.730 58.900 89.130 58.950 ;
        RECT 78.730 58.650 80.180 58.900 ;
        RECT 80.330 58.800 89.130 58.900 ;
        RECT 78.730 58.450 82.930 58.650 ;
        RECT 66.530 58.300 74.080 58.450 ;
        RECT 75.430 58.300 82.930 58.450 ;
        RECT 66.530 58.000 70.730 58.300 ;
        RECT 66.530 55.150 66.680 58.000 ;
        RECT 67.130 50.450 67.280 58.000 ;
        RECT 67.730 50.450 67.880 58.000 ;
        RECT 68.330 50.450 68.480 58.000 ;
        RECT 68.930 50.450 69.080 58.000 ;
        RECT 69.530 50.450 69.680 58.000 ;
        RECT 70.130 57.850 70.730 58.000 ;
        RECT 78.730 58.000 82.930 58.300 ;
        RECT 78.730 57.850 79.330 58.000 ;
        RECT 70.130 57.700 74.080 57.850 ;
        RECT 75.380 57.700 79.330 57.850 ;
        RECT 70.130 57.250 70.730 57.700 ;
        RECT 78.730 57.250 79.330 57.700 ;
        RECT 70.130 57.100 74.080 57.250 ;
        RECT 75.380 57.100 79.330 57.250 ;
        RECT 70.130 56.650 70.730 57.100 ;
        RECT 78.730 56.650 79.330 57.100 ;
        RECT 70.130 56.500 74.080 56.650 ;
        RECT 75.380 56.500 79.330 56.650 ;
        RECT 70.130 56.050 70.730 56.500 ;
        RECT 78.730 56.050 79.330 56.500 ;
        RECT 70.130 55.900 74.080 56.050 ;
        RECT 75.380 55.900 79.330 56.050 ;
        RECT 70.130 55.450 70.730 55.900 ;
        RECT 78.730 55.450 79.330 55.900 ;
        RECT 70.130 55.300 74.080 55.450 ;
        RECT 75.380 55.300 79.330 55.450 ;
        RECT 70.130 54.850 70.730 55.300 ;
        RECT 78.730 54.850 79.330 55.300 ;
        RECT 70.130 54.700 74.080 54.850 ;
        RECT 75.380 54.700 79.330 54.850 ;
        RECT 70.130 54.250 70.730 54.700 ;
        RECT 78.730 54.250 79.330 54.700 ;
        RECT 70.130 54.100 74.080 54.250 ;
        RECT 75.380 54.100 79.330 54.250 ;
        RECT 70.130 53.650 70.730 54.100 ;
        RECT 78.730 53.650 79.330 54.100 ;
        RECT 70.130 53.500 74.080 53.650 ;
        RECT 75.380 53.500 79.330 53.650 ;
        RECT 70.130 53.050 70.730 53.500 ;
        RECT 78.730 53.050 79.330 53.500 ;
        RECT 70.130 52.900 74.080 53.050 ;
        RECT 75.380 52.900 79.330 53.050 ;
        RECT 70.130 52.450 70.730 52.900 ;
        RECT 78.730 52.450 79.330 52.900 ;
        RECT 70.130 52.300 74.080 52.450 ;
        RECT 75.380 52.300 79.330 52.450 ;
        RECT 70.130 51.850 70.730 52.300 ;
        RECT 78.730 51.850 79.330 52.300 ;
        RECT 70.130 51.700 74.080 51.850 ;
        RECT 75.380 51.700 79.330 51.850 ;
        RECT 70.130 51.250 70.730 51.700 ;
        RECT 78.730 51.250 79.330 51.700 ;
        RECT 70.130 51.100 74.080 51.250 ;
        RECT 75.380 51.100 79.330 51.250 ;
        RECT 70.130 50.650 70.730 51.100 ;
        RECT 78.730 50.650 79.330 51.100 ;
        RECT 70.130 50.450 74.080 50.650 ;
        RECT 75.380 50.450 79.330 50.650 ;
        RECT 79.780 50.450 79.930 58.000 ;
        RECT 80.380 50.450 80.530 58.000 ;
        RECT 80.980 50.450 81.130 58.000 ;
        RECT 81.580 50.450 81.730 58.000 ;
        RECT 82.180 50.450 82.330 58.000 ;
        RECT 82.780 55.150 82.930 58.000 ;
        RECT 83.530 55.600 85.930 58.800 ;
        RECT 89.280 58.650 90.730 58.950 ;
        RECT 86.530 58.450 90.730 58.650 ;
        RECT 98.730 58.900 104.730 59.800 ;
        RECT 98.730 58.650 100.180 58.900 ;
        RECT 100.330 58.800 104.730 58.900 ;
        RECT 98.730 58.450 102.930 58.650 ;
        RECT 86.530 58.300 94.080 58.450 ;
        RECT 95.430 58.300 102.930 58.450 ;
        RECT 86.530 58.000 90.730 58.300 ;
        RECT 86.530 55.150 86.680 58.000 ;
        RECT 87.130 50.450 87.280 58.000 ;
        RECT 87.730 50.450 87.880 58.000 ;
        RECT 88.330 50.450 88.480 58.000 ;
        RECT 88.930 50.450 89.080 58.000 ;
        RECT 89.530 50.450 89.680 58.000 ;
        RECT 90.130 57.850 90.730 58.000 ;
        RECT 98.730 58.000 102.930 58.300 ;
        RECT 98.730 57.850 99.330 58.000 ;
        RECT 90.130 57.700 94.080 57.850 ;
        RECT 95.380 57.700 99.330 57.850 ;
        RECT 90.130 57.250 90.730 57.700 ;
        RECT 98.730 57.250 99.330 57.700 ;
        RECT 90.130 57.100 94.080 57.250 ;
        RECT 95.380 57.100 99.330 57.250 ;
        RECT 90.130 56.650 90.730 57.100 ;
        RECT 98.730 56.650 99.330 57.100 ;
        RECT 90.130 56.500 94.080 56.650 ;
        RECT 95.380 56.500 99.330 56.650 ;
        RECT 90.130 56.050 90.730 56.500 ;
        RECT 98.730 56.050 99.330 56.500 ;
        RECT 90.130 55.900 94.080 56.050 ;
        RECT 95.380 55.900 99.330 56.050 ;
        RECT 90.130 55.450 90.730 55.900 ;
        RECT 98.730 55.450 99.330 55.900 ;
        RECT 90.130 55.300 94.080 55.450 ;
        RECT 95.380 55.300 99.330 55.450 ;
        RECT 90.130 54.850 90.730 55.300 ;
        RECT 98.730 54.850 99.330 55.300 ;
        RECT 90.130 54.700 94.080 54.850 ;
        RECT 95.380 54.700 99.330 54.850 ;
        RECT 90.130 54.250 90.730 54.700 ;
        RECT 98.730 54.250 99.330 54.700 ;
        RECT 90.130 54.100 94.080 54.250 ;
        RECT 95.380 54.100 99.330 54.250 ;
        RECT 90.130 53.650 90.730 54.100 ;
        RECT 98.730 53.650 99.330 54.100 ;
        RECT 90.130 53.500 94.080 53.650 ;
        RECT 95.380 53.500 99.330 53.650 ;
        RECT 90.130 53.050 90.730 53.500 ;
        RECT 98.730 53.050 99.330 53.500 ;
        RECT 90.130 52.900 94.080 53.050 ;
        RECT 95.380 52.900 99.330 53.050 ;
        RECT 90.130 52.450 90.730 52.900 ;
        RECT 98.730 52.450 99.330 52.900 ;
        RECT 90.130 52.300 94.080 52.450 ;
        RECT 95.380 52.300 99.330 52.450 ;
        RECT 90.130 51.850 90.730 52.300 ;
        RECT 98.730 51.850 99.330 52.300 ;
        RECT 90.130 51.700 94.080 51.850 ;
        RECT 95.380 51.700 99.330 51.850 ;
        RECT 90.130 51.250 90.730 51.700 ;
        RECT 98.730 51.250 99.330 51.700 ;
        RECT 90.130 51.100 94.080 51.250 ;
        RECT 95.380 51.100 99.330 51.250 ;
        RECT 90.130 50.650 90.730 51.100 ;
        RECT 98.730 50.650 99.330 51.100 ;
        RECT 90.130 50.450 94.080 50.650 ;
        RECT 95.380 50.450 99.330 50.650 ;
        RECT 99.780 50.450 99.930 58.000 ;
        RECT 100.380 50.450 100.530 58.000 ;
        RECT 100.980 50.450 101.130 58.000 ;
        RECT 101.580 50.450 101.730 58.000 ;
        RECT 102.180 50.450 102.330 58.000 ;
        RECT 102.780 55.150 102.930 58.000 ;
        RECT 103.530 57.310 104.730 58.800 ;
        RECT 103.530 56.035 107.135 57.310 ;
        RECT 103.530 55.600 104.730 56.035 ;
        RECT 2.315 44.445 4.315 46.740 ;
        RECT 4.730 43.320 5.930 44.400 ;
        RECT 2.315 42.045 5.930 43.320 ;
        RECT 4.730 41.200 5.930 42.045 ;
        RECT 6.530 42.000 6.680 44.900 ;
        RECT 7.130 42.000 7.280 49.550 ;
        RECT 7.730 42.000 7.880 49.550 ;
        RECT 8.330 42.000 8.480 49.550 ;
        RECT 8.930 42.000 9.080 49.550 ;
        RECT 9.530 42.000 9.680 49.550 ;
        RECT 10.130 49.350 14.080 49.550 ;
        RECT 15.380 49.350 19.330 49.550 ;
        RECT 10.130 48.900 10.730 49.350 ;
        RECT 18.730 48.900 19.330 49.350 ;
        RECT 10.130 48.750 14.080 48.900 ;
        RECT 15.380 48.750 19.330 48.900 ;
        RECT 10.130 48.300 10.730 48.750 ;
        RECT 18.730 48.300 19.330 48.750 ;
        RECT 10.130 48.150 14.080 48.300 ;
        RECT 15.380 48.150 19.330 48.300 ;
        RECT 10.130 47.700 10.730 48.150 ;
        RECT 18.730 47.700 19.330 48.150 ;
        RECT 10.130 47.550 14.080 47.700 ;
        RECT 15.380 47.550 19.330 47.700 ;
        RECT 10.130 47.100 10.730 47.550 ;
        RECT 18.730 47.100 19.330 47.550 ;
        RECT 10.130 46.950 14.080 47.100 ;
        RECT 15.380 46.950 19.330 47.100 ;
        RECT 10.130 46.500 10.730 46.950 ;
        RECT 18.730 46.500 19.330 46.950 ;
        RECT 10.130 46.350 14.080 46.500 ;
        RECT 15.380 46.350 19.330 46.500 ;
        RECT 10.130 45.900 10.730 46.350 ;
        RECT 18.730 45.900 19.330 46.350 ;
        RECT 10.130 45.750 14.080 45.900 ;
        RECT 15.380 45.750 19.330 45.900 ;
        RECT 10.130 45.300 10.730 45.750 ;
        RECT 18.730 45.300 19.330 45.750 ;
        RECT 10.130 45.150 14.080 45.300 ;
        RECT 15.380 45.150 19.330 45.300 ;
        RECT 10.130 44.700 10.730 45.150 ;
        RECT 18.730 44.700 19.330 45.150 ;
        RECT 10.130 44.550 14.080 44.700 ;
        RECT 15.380 44.550 19.330 44.700 ;
        RECT 10.130 44.100 10.730 44.550 ;
        RECT 18.730 44.100 19.330 44.550 ;
        RECT 10.130 43.950 14.080 44.100 ;
        RECT 15.380 43.950 19.330 44.100 ;
        RECT 10.130 43.500 10.730 43.950 ;
        RECT 18.730 43.500 19.330 43.950 ;
        RECT 10.130 43.350 14.080 43.500 ;
        RECT 15.380 43.350 19.330 43.500 ;
        RECT 10.130 42.900 10.730 43.350 ;
        RECT 18.730 42.900 19.330 43.350 ;
        RECT 10.130 42.750 14.080 42.900 ;
        RECT 15.380 42.750 19.330 42.900 ;
        RECT 10.130 42.300 10.730 42.750 ;
        RECT 18.730 42.300 19.330 42.750 ;
        RECT 10.130 42.150 14.080 42.300 ;
        RECT 15.380 42.150 19.330 42.300 ;
        RECT 10.130 42.000 10.730 42.150 ;
        RECT 6.530 41.700 10.730 42.000 ;
        RECT 18.730 42.000 19.330 42.150 ;
        RECT 19.780 42.000 19.930 49.550 ;
        RECT 20.380 42.000 20.530 49.550 ;
        RECT 20.980 42.000 21.130 49.550 ;
        RECT 21.580 42.000 21.730 49.550 ;
        RECT 22.180 42.000 22.330 49.550 ;
        RECT 22.780 42.000 22.930 44.900 ;
        RECT 18.730 41.700 22.930 42.000 ;
        RECT 6.530 41.550 14.080 41.700 ;
        RECT 15.380 41.550 22.930 41.700 ;
        RECT 6.530 41.350 10.730 41.550 ;
        RECT 4.730 41.050 9.130 41.200 ;
        RECT 9.280 41.050 10.730 41.350 ;
        RECT 4.730 40.150 10.730 41.050 ;
        RECT 18.730 41.350 22.930 41.550 ;
        RECT 18.730 41.050 20.180 41.350 ;
        RECT 23.530 41.200 25.930 44.400 ;
        RECT 26.530 42.000 26.680 44.900 ;
        RECT 27.130 42.000 27.280 49.550 ;
        RECT 27.730 42.000 27.880 49.550 ;
        RECT 28.330 42.000 28.480 49.550 ;
        RECT 28.930 42.000 29.080 49.550 ;
        RECT 29.530 42.000 29.680 49.550 ;
        RECT 30.130 49.350 34.080 49.550 ;
        RECT 35.380 49.350 39.330 49.550 ;
        RECT 30.130 48.900 30.730 49.350 ;
        RECT 38.730 48.900 39.330 49.350 ;
        RECT 30.130 48.750 34.080 48.900 ;
        RECT 35.380 48.750 39.330 48.900 ;
        RECT 30.130 48.300 30.730 48.750 ;
        RECT 38.730 48.300 39.330 48.750 ;
        RECT 30.130 48.150 34.080 48.300 ;
        RECT 35.380 48.150 39.330 48.300 ;
        RECT 30.130 47.700 30.730 48.150 ;
        RECT 38.730 47.700 39.330 48.150 ;
        RECT 30.130 47.550 34.080 47.700 ;
        RECT 35.380 47.550 39.330 47.700 ;
        RECT 30.130 47.100 30.730 47.550 ;
        RECT 38.730 47.100 39.330 47.550 ;
        RECT 30.130 46.950 34.080 47.100 ;
        RECT 35.380 46.950 39.330 47.100 ;
        RECT 30.130 46.500 30.730 46.950 ;
        RECT 38.730 46.500 39.330 46.950 ;
        RECT 30.130 46.350 34.080 46.500 ;
        RECT 35.380 46.350 39.330 46.500 ;
        RECT 30.130 45.900 30.730 46.350 ;
        RECT 38.730 45.900 39.330 46.350 ;
        RECT 30.130 45.750 34.080 45.900 ;
        RECT 35.380 45.750 39.330 45.900 ;
        RECT 30.130 45.300 30.730 45.750 ;
        RECT 38.730 45.300 39.330 45.750 ;
        RECT 30.130 45.150 34.080 45.300 ;
        RECT 35.380 45.150 39.330 45.300 ;
        RECT 30.130 44.700 30.730 45.150 ;
        RECT 38.730 44.700 39.330 45.150 ;
        RECT 30.130 44.550 34.080 44.700 ;
        RECT 35.380 44.550 39.330 44.700 ;
        RECT 30.130 44.100 30.730 44.550 ;
        RECT 38.730 44.100 39.330 44.550 ;
        RECT 30.130 43.950 34.080 44.100 ;
        RECT 35.380 43.950 39.330 44.100 ;
        RECT 30.130 43.500 30.730 43.950 ;
        RECT 38.730 43.500 39.330 43.950 ;
        RECT 30.130 43.350 34.080 43.500 ;
        RECT 35.380 43.350 39.330 43.500 ;
        RECT 30.130 42.900 30.730 43.350 ;
        RECT 38.730 42.900 39.330 43.350 ;
        RECT 30.130 42.750 34.080 42.900 ;
        RECT 35.380 42.750 39.330 42.900 ;
        RECT 30.130 42.300 30.730 42.750 ;
        RECT 38.730 42.300 39.330 42.750 ;
        RECT 30.130 42.150 34.080 42.300 ;
        RECT 35.380 42.150 39.330 42.300 ;
        RECT 30.130 42.000 30.730 42.150 ;
        RECT 26.530 41.700 30.730 42.000 ;
        RECT 38.730 42.000 39.330 42.150 ;
        RECT 39.780 42.000 39.930 49.550 ;
        RECT 40.380 42.000 40.530 49.550 ;
        RECT 40.980 42.000 41.130 49.550 ;
        RECT 41.580 42.000 41.730 49.550 ;
        RECT 42.180 42.000 42.330 49.550 ;
        RECT 42.780 42.000 42.930 44.900 ;
        RECT 38.730 41.700 42.930 42.000 ;
        RECT 26.530 41.550 34.080 41.700 ;
        RECT 35.380 41.550 42.930 41.700 ;
        RECT 26.530 41.350 30.730 41.550 ;
        RECT 20.330 41.050 29.130 41.200 ;
        RECT 29.280 41.050 30.730 41.350 ;
        RECT 18.730 40.150 30.730 41.050 ;
        RECT 38.730 41.350 42.930 41.550 ;
        RECT 38.730 41.050 40.180 41.350 ;
        RECT 43.530 41.200 45.930 44.400 ;
        RECT 46.530 42.000 46.680 44.900 ;
        RECT 47.130 42.000 47.280 49.550 ;
        RECT 47.730 42.000 47.880 49.550 ;
        RECT 48.330 42.000 48.480 49.550 ;
        RECT 48.930 42.000 49.080 49.550 ;
        RECT 49.530 42.000 49.680 49.550 ;
        RECT 50.130 49.350 54.080 49.550 ;
        RECT 55.380 49.350 59.330 49.550 ;
        RECT 50.130 48.900 50.730 49.350 ;
        RECT 58.730 48.900 59.330 49.350 ;
        RECT 50.130 48.750 54.080 48.900 ;
        RECT 55.380 48.750 59.330 48.900 ;
        RECT 50.130 48.300 50.730 48.750 ;
        RECT 58.730 48.300 59.330 48.750 ;
        RECT 50.130 48.150 54.080 48.300 ;
        RECT 55.380 48.150 59.330 48.300 ;
        RECT 50.130 47.700 50.730 48.150 ;
        RECT 58.730 47.700 59.330 48.150 ;
        RECT 50.130 47.550 54.080 47.700 ;
        RECT 55.380 47.550 59.330 47.700 ;
        RECT 50.130 47.100 50.730 47.550 ;
        RECT 58.730 47.100 59.330 47.550 ;
        RECT 50.130 46.950 54.080 47.100 ;
        RECT 55.380 46.950 59.330 47.100 ;
        RECT 50.130 46.500 50.730 46.950 ;
        RECT 58.730 46.500 59.330 46.950 ;
        RECT 50.130 46.350 54.080 46.500 ;
        RECT 55.380 46.350 59.330 46.500 ;
        RECT 50.130 45.900 50.730 46.350 ;
        RECT 58.730 45.900 59.330 46.350 ;
        RECT 50.130 45.750 54.080 45.900 ;
        RECT 55.380 45.750 59.330 45.900 ;
        RECT 50.130 45.300 50.730 45.750 ;
        RECT 58.730 45.300 59.330 45.750 ;
        RECT 50.130 45.150 54.080 45.300 ;
        RECT 55.380 45.150 59.330 45.300 ;
        RECT 50.130 44.700 50.730 45.150 ;
        RECT 58.730 44.700 59.330 45.150 ;
        RECT 50.130 44.550 54.080 44.700 ;
        RECT 55.380 44.550 59.330 44.700 ;
        RECT 50.130 44.100 50.730 44.550 ;
        RECT 58.730 44.100 59.330 44.550 ;
        RECT 50.130 43.950 54.080 44.100 ;
        RECT 55.380 43.950 59.330 44.100 ;
        RECT 50.130 43.500 50.730 43.950 ;
        RECT 58.730 43.500 59.330 43.950 ;
        RECT 50.130 43.350 54.080 43.500 ;
        RECT 55.380 43.350 59.330 43.500 ;
        RECT 50.130 42.900 50.730 43.350 ;
        RECT 58.730 42.900 59.330 43.350 ;
        RECT 50.130 42.750 54.080 42.900 ;
        RECT 55.380 42.750 59.330 42.900 ;
        RECT 50.130 42.300 50.730 42.750 ;
        RECT 58.730 42.300 59.330 42.750 ;
        RECT 50.130 42.150 54.080 42.300 ;
        RECT 55.380 42.150 59.330 42.300 ;
        RECT 50.130 42.000 50.730 42.150 ;
        RECT 46.530 41.700 50.730 42.000 ;
        RECT 58.730 42.000 59.330 42.150 ;
        RECT 59.780 42.000 59.930 49.550 ;
        RECT 60.380 42.000 60.530 49.550 ;
        RECT 60.980 42.000 61.130 49.550 ;
        RECT 61.580 42.000 61.730 49.550 ;
        RECT 62.180 42.000 62.330 49.550 ;
        RECT 62.780 42.000 62.930 44.900 ;
        RECT 58.730 41.700 62.930 42.000 ;
        RECT 46.530 41.550 54.080 41.700 ;
        RECT 55.380 41.550 62.930 41.700 ;
        RECT 46.530 41.350 50.730 41.550 ;
        RECT 40.330 41.050 49.130 41.200 ;
        RECT 49.280 41.050 50.730 41.350 ;
        RECT 38.730 40.150 50.730 41.050 ;
        RECT 58.730 41.350 62.930 41.550 ;
        RECT 58.730 41.050 60.180 41.350 ;
        RECT 63.530 41.200 65.930 44.400 ;
        RECT 66.530 42.000 66.680 44.900 ;
        RECT 67.130 42.000 67.280 49.550 ;
        RECT 67.730 42.000 67.880 49.550 ;
        RECT 68.330 42.000 68.480 49.550 ;
        RECT 68.930 42.000 69.080 49.550 ;
        RECT 69.530 42.000 69.680 49.550 ;
        RECT 70.130 49.350 74.080 49.550 ;
        RECT 75.380 49.350 79.330 49.550 ;
        RECT 70.130 48.900 70.730 49.350 ;
        RECT 78.730 48.900 79.330 49.350 ;
        RECT 70.130 48.750 74.080 48.900 ;
        RECT 75.380 48.750 79.330 48.900 ;
        RECT 70.130 48.300 70.730 48.750 ;
        RECT 78.730 48.300 79.330 48.750 ;
        RECT 70.130 48.150 74.080 48.300 ;
        RECT 75.380 48.150 79.330 48.300 ;
        RECT 70.130 47.700 70.730 48.150 ;
        RECT 78.730 47.700 79.330 48.150 ;
        RECT 70.130 47.550 74.080 47.700 ;
        RECT 75.380 47.550 79.330 47.700 ;
        RECT 70.130 47.100 70.730 47.550 ;
        RECT 78.730 47.100 79.330 47.550 ;
        RECT 70.130 46.950 74.080 47.100 ;
        RECT 75.380 46.950 79.330 47.100 ;
        RECT 70.130 46.500 70.730 46.950 ;
        RECT 78.730 46.500 79.330 46.950 ;
        RECT 70.130 46.350 74.080 46.500 ;
        RECT 75.380 46.350 79.330 46.500 ;
        RECT 70.130 45.900 70.730 46.350 ;
        RECT 78.730 45.900 79.330 46.350 ;
        RECT 70.130 45.750 74.080 45.900 ;
        RECT 75.380 45.750 79.330 45.900 ;
        RECT 70.130 45.300 70.730 45.750 ;
        RECT 78.730 45.300 79.330 45.750 ;
        RECT 70.130 45.150 74.080 45.300 ;
        RECT 75.380 45.150 79.330 45.300 ;
        RECT 70.130 44.700 70.730 45.150 ;
        RECT 78.730 44.700 79.330 45.150 ;
        RECT 70.130 44.550 74.080 44.700 ;
        RECT 75.380 44.550 79.330 44.700 ;
        RECT 70.130 44.100 70.730 44.550 ;
        RECT 78.730 44.100 79.330 44.550 ;
        RECT 70.130 43.950 74.080 44.100 ;
        RECT 75.380 43.950 79.330 44.100 ;
        RECT 70.130 43.500 70.730 43.950 ;
        RECT 78.730 43.500 79.330 43.950 ;
        RECT 70.130 43.350 74.080 43.500 ;
        RECT 75.380 43.350 79.330 43.500 ;
        RECT 70.130 42.900 70.730 43.350 ;
        RECT 78.730 42.900 79.330 43.350 ;
        RECT 70.130 42.750 74.080 42.900 ;
        RECT 75.380 42.750 79.330 42.900 ;
        RECT 70.130 42.300 70.730 42.750 ;
        RECT 78.730 42.300 79.330 42.750 ;
        RECT 70.130 42.150 74.080 42.300 ;
        RECT 75.380 42.150 79.330 42.300 ;
        RECT 70.130 42.000 70.730 42.150 ;
        RECT 66.530 41.700 70.730 42.000 ;
        RECT 78.730 42.000 79.330 42.150 ;
        RECT 79.780 42.000 79.930 49.550 ;
        RECT 80.380 42.000 80.530 49.550 ;
        RECT 80.980 42.000 81.130 49.550 ;
        RECT 81.580 42.000 81.730 49.550 ;
        RECT 82.180 42.000 82.330 49.550 ;
        RECT 82.780 42.000 82.930 44.900 ;
        RECT 78.730 41.700 82.930 42.000 ;
        RECT 66.530 41.550 74.080 41.700 ;
        RECT 75.380 41.550 82.930 41.700 ;
        RECT 66.530 41.350 70.730 41.550 ;
        RECT 60.330 41.050 69.130 41.200 ;
        RECT 69.280 41.050 70.730 41.350 ;
        RECT 58.730 40.150 70.730 41.050 ;
        RECT 78.730 41.350 82.930 41.550 ;
        RECT 78.730 41.050 80.180 41.350 ;
        RECT 83.530 41.200 85.930 44.400 ;
        RECT 86.530 42.000 86.680 44.900 ;
        RECT 87.130 42.000 87.280 49.550 ;
        RECT 87.730 42.000 87.880 49.550 ;
        RECT 88.330 42.000 88.480 49.550 ;
        RECT 88.930 42.000 89.080 49.550 ;
        RECT 89.530 42.000 89.680 49.550 ;
        RECT 90.130 49.350 94.080 49.550 ;
        RECT 95.380 49.350 99.330 49.550 ;
        RECT 90.130 48.900 90.730 49.350 ;
        RECT 98.730 48.900 99.330 49.350 ;
        RECT 90.130 48.750 94.080 48.900 ;
        RECT 95.380 48.750 99.330 48.900 ;
        RECT 90.130 48.300 90.730 48.750 ;
        RECT 98.730 48.300 99.330 48.750 ;
        RECT 90.130 48.150 94.080 48.300 ;
        RECT 95.380 48.150 99.330 48.300 ;
        RECT 90.130 47.700 90.730 48.150 ;
        RECT 98.730 47.700 99.330 48.150 ;
        RECT 90.130 47.550 94.080 47.700 ;
        RECT 95.380 47.550 99.330 47.700 ;
        RECT 90.130 47.100 90.730 47.550 ;
        RECT 98.730 47.100 99.330 47.550 ;
        RECT 90.130 46.950 94.080 47.100 ;
        RECT 95.380 46.950 99.330 47.100 ;
        RECT 90.130 46.500 90.730 46.950 ;
        RECT 98.730 46.500 99.330 46.950 ;
        RECT 90.130 46.350 94.080 46.500 ;
        RECT 95.380 46.350 99.330 46.500 ;
        RECT 90.130 45.900 90.730 46.350 ;
        RECT 98.730 45.900 99.330 46.350 ;
        RECT 90.130 45.750 94.080 45.900 ;
        RECT 95.380 45.750 99.330 45.900 ;
        RECT 90.130 45.300 90.730 45.750 ;
        RECT 98.730 45.300 99.330 45.750 ;
        RECT 90.130 45.150 94.080 45.300 ;
        RECT 95.380 45.150 99.330 45.300 ;
        RECT 90.130 44.700 90.730 45.150 ;
        RECT 98.730 44.700 99.330 45.150 ;
        RECT 90.130 44.550 94.080 44.700 ;
        RECT 95.380 44.550 99.330 44.700 ;
        RECT 90.130 44.100 90.730 44.550 ;
        RECT 98.730 44.100 99.330 44.550 ;
        RECT 90.130 43.950 94.080 44.100 ;
        RECT 95.380 43.950 99.330 44.100 ;
        RECT 90.130 43.500 90.730 43.950 ;
        RECT 98.730 43.500 99.330 43.950 ;
        RECT 90.130 43.350 94.080 43.500 ;
        RECT 95.380 43.350 99.330 43.500 ;
        RECT 90.130 42.900 90.730 43.350 ;
        RECT 98.730 42.900 99.330 43.350 ;
        RECT 90.130 42.750 94.080 42.900 ;
        RECT 95.380 42.750 99.330 42.900 ;
        RECT 90.130 42.300 90.730 42.750 ;
        RECT 98.730 42.300 99.330 42.750 ;
        RECT 90.130 42.150 94.080 42.300 ;
        RECT 95.380 42.150 99.330 42.300 ;
        RECT 90.130 42.000 90.730 42.150 ;
        RECT 86.530 41.700 90.730 42.000 ;
        RECT 98.730 42.000 99.330 42.150 ;
        RECT 99.780 42.000 99.930 49.550 ;
        RECT 100.380 42.000 100.530 49.550 ;
        RECT 100.980 42.000 101.130 49.550 ;
        RECT 101.580 42.000 101.730 49.550 ;
        RECT 102.180 42.000 102.330 49.550 ;
        RECT 102.780 42.000 102.930 44.900 ;
        RECT 98.730 41.700 102.930 42.000 ;
        RECT 86.530 41.550 94.080 41.700 ;
        RECT 95.380 41.550 102.930 41.700 ;
        RECT 86.530 41.350 90.730 41.550 ;
        RECT 80.330 41.050 89.130 41.200 ;
        RECT 89.280 41.050 90.730 41.350 ;
        RECT 78.730 40.150 90.730 41.050 ;
        RECT 98.730 41.350 102.930 41.550 ;
        RECT 103.530 43.095 104.730 44.400 ;
        RECT 103.530 41.820 107.140 43.095 ;
        RECT 98.730 41.050 100.180 41.350 ;
        RECT 103.530 41.200 104.730 41.820 ;
        RECT 100.330 41.050 104.730 41.200 ;
        RECT 98.730 40.150 104.730 41.050 ;
        RECT 4.730 39.850 9.130 40.150 ;
        RECT 20.330 39.850 29.130 40.150 ;
        RECT 40.330 39.850 49.130 40.150 ;
        RECT 60.330 39.850 69.130 40.150 ;
        RECT 80.330 39.850 89.130 40.150 ;
        RECT 4.730 38.950 10.730 39.850 ;
        RECT 20.330 39.800 30.730 39.850 ;
        RECT 40.330 39.800 50.730 39.850 ;
        RECT 60.330 39.800 70.730 39.850 ;
        RECT 80.330 39.800 90.730 39.850 ;
        RECT 100.330 39.800 104.730 40.150 ;
        RECT 4.730 38.800 9.130 38.950 ;
        RECT 4.730 37.765 5.930 38.800 ;
        RECT 9.280 38.650 10.730 38.950 ;
        RECT 2.315 36.490 5.930 37.765 ;
        RECT 4.730 35.600 5.930 36.490 ;
        RECT 6.530 38.450 10.730 38.650 ;
        RECT 18.730 38.950 30.730 39.800 ;
        RECT 18.730 38.900 29.130 38.950 ;
        RECT 18.730 38.650 20.180 38.900 ;
        RECT 20.330 38.800 29.130 38.900 ;
        RECT 18.730 38.450 22.930 38.650 ;
        RECT 6.530 38.300 14.080 38.450 ;
        RECT 15.430 38.300 22.930 38.450 ;
        RECT 6.530 38.000 10.730 38.300 ;
        RECT 2.315 33.255 4.315 35.550 ;
        RECT 6.530 35.150 6.680 38.000 ;
        RECT 7.130 30.450 7.280 38.000 ;
        RECT 7.730 30.450 7.880 38.000 ;
        RECT 8.330 30.450 8.480 38.000 ;
        RECT 8.930 30.450 9.080 38.000 ;
        RECT 9.530 30.450 9.680 38.000 ;
        RECT 10.130 37.850 10.730 38.000 ;
        RECT 18.730 38.000 22.930 38.300 ;
        RECT 18.730 37.850 19.330 38.000 ;
        RECT 10.130 37.700 14.080 37.850 ;
        RECT 15.380 37.700 19.330 37.850 ;
        RECT 10.130 37.250 10.730 37.700 ;
        RECT 18.730 37.250 19.330 37.700 ;
        RECT 10.130 37.100 14.080 37.250 ;
        RECT 15.380 37.100 19.330 37.250 ;
        RECT 10.130 36.650 10.730 37.100 ;
        RECT 18.730 36.650 19.330 37.100 ;
        RECT 10.130 36.500 14.080 36.650 ;
        RECT 15.380 36.500 19.330 36.650 ;
        RECT 10.130 36.050 10.730 36.500 ;
        RECT 18.730 36.050 19.330 36.500 ;
        RECT 10.130 35.900 14.080 36.050 ;
        RECT 15.380 35.900 19.330 36.050 ;
        RECT 10.130 35.450 10.730 35.900 ;
        RECT 18.730 35.450 19.330 35.900 ;
        RECT 10.130 35.300 14.080 35.450 ;
        RECT 15.380 35.300 19.330 35.450 ;
        RECT 10.130 34.850 10.730 35.300 ;
        RECT 18.730 34.850 19.330 35.300 ;
        RECT 10.130 34.700 14.080 34.850 ;
        RECT 15.380 34.700 19.330 34.850 ;
        RECT 10.130 34.250 10.730 34.700 ;
        RECT 18.730 34.250 19.330 34.700 ;
        RECT 10.130 34.100 14.080 34.250 ;
        RECT 15.380 34.100 19.330 34.250 ;
        RECT 10.130 33.650 10.730 34.100 ;
        RECT 18.730 33.650 19.330 34.100 ;
        RECT 10.130 33.500 14.080 33.650 ;
        RECT 15.380 33.500 19.330 33.650 ;
        RECT 10.130 33.050 10.730 33.500 ;
        RECT 18.730 33.050 19.330 33.500 ;
        RECT 10.130 32.900 14.080 33.050 ;
        RECT 15.380 32.900 19.330 33.050 ;
        RECT 10.130 32.450 10.730 32.900 ;
        RECT 18.730 32.450 19.330 32.900 ;
        RECT 10.130 32.300 14.080 32.450 ;
        RECT 15.380 32.300 19.330 32.450 ;
        RECT 10.130 31.850 10.730 32.300 ;
        RECT 18.730 31.850 19.330 32.300 ;
        RECT 10.130 31.700 14.080 31.850 ;
        RECT 15.380 31.700 19.330 31.850 ;
        RECT 10.130 31.250 10.730 31.700 ;
        RECT 18.730 31.250 19.330 31.700 ;
        RECT 10.130 31.100 14.080 31.250 ;
        RECT 15.380 31.100 19.330 31.250 ;
        RECT 10.130 30.650 10.730 31.100 ;
        RECT 18.730 30.650 19.330 31.100 ;
        RECT 10.130 30.450 14.080 30.650 ;
        RECT 15.380 30.450 19.330 30.650 ;
        RECT 19.780 30.450 19.930 38.000 ;
        RECT 20.380 30.450 20.530 38.000 ;
        RECT 20.980 30.450 21.130 38.000 ;
        RECT 21.580 30.450 21.730 38.000 ;
        RECT 22.180 30.450 22.330 38.000 ;
        RECT 22.780 35.150 22.930 38.000 ;
        RECT 23.530 35.600 25.930 38.800 ;
        RECT 29.280 38.650 30.730 38.950 ;
        RECT 26.530 38.450 30.730 38.650 ;
        RECT 38.730 38.950 50.730 39.800 ;
        RECT 38.730 38.900 49.130 38.950 ;
        RECT 38.730 38.650 40.180 38.900 ;
        RECT 40.330 38.800 49.130 38.900 ;
        RECT 38.730 38.450 42.930 38.650 ;
        RECT 26.530 38.300 34.080 38.450 ;
        RECT 35.430 38.300 42.930 38.450 ;
        RECT 26.530 38.000 30.730 38.300 ;
        RECT 26.530 35.150 26.680 38.000 ;
        RECT 27.130 30.450 27.280 38.000 ;
        RECT 27.730 30.450 27.880 38.000 ;
        RECT 28.330 30.450 28.480 38.000 ;
        RECT 28.930 30.450 29.080 38.000 ;
        RECT 29.530 30.450 29.680 38.000 ;
        RECT 30.130 37.850 30.730 38.000 ;
        RECT 38.730 38.000 42.930 38.300 ;
        RECT 38.730 37.850 39.330 38.000 ;
        RECT 30.130 37.700 34.080 37.850 ;
        RECT 35.380 37.700 39.330 37.850 ;
        RECT 30.130 37.250 30.730 37.700 ;
        RECT 38.730 37.250 39.330 37.700 ;
        RECT 30.130 37.100 34.080 37.250 ;
        RECT 35.380 37.100 39.330 37.250 ;
        RECT 30.130 36.650 30.730 37.100 ;
        RECT 38.730 36.650 39.330 37.100 ;
        RECT 30.130 36.500 34.080 36.650 ;
        RECT 35.380 36.500 39.330 36.650 ;
        RECT 30.130 36.050 30.730 36.500 ;
        RECT 38.730 36.050 39.330 36.500 ;
        RECT 30.130 35.900 34.080 36.050 ;
        RECT 35.380 35.900 39.330 36.050 ;
        RECT 30.130 35.450 30.730 35.900 ;
        RECT 38.730 35.450 39.330 35.900 ;
        RECT 30.130 35.300 34.080 35.450 ;
        RECT 35.380 35.300 39.330 35.450 ;
        RECT 30.130 34.850 30.730 35.300 ;
        RECT 38.730 34.850 39.330 35.300 ;
        RECT 30.130 34.700 34.080 34.850 ;
        RECT 35.380 34.700 39.330 34.850 ;
        RECT 30.130 34.250 30.730 34.700 ;
        RECT 38.730 34.250 39.330 34.700 ;
        RECT 30.130 34.100 34.080 34.250 ;
        RECT 35.380 34.100 39.330 34.250 ;
        RECT 30.130 33.650 30.730 34.100 ;
        RECT 38.730 33.650 39.330 34.100 ;
        RECT 30.130 33.500 34.080 33.650 ;
        RECT 35.380 33.500 39.330 33.650 ;
        RECT 30.130 33.050 30.730 33.500 ;
        RECT 38.730 33.050 39.330 33.500 ;
        RECT 30.130 32.900 34.080 33.050 ;
        RECT 35.380 32.900 39.330 33.050 ;
        RECT 30.130 32.450 30.730 32.900 ;
        RECT 38.730 32.450 39.330 32.900 ;
        RECT 30.130 32.300 34.080 32.450 ;
        RECT 35.380 32.300 39.330 32.450 ;
        RECT 30.130 31.850 30.730 32.300 ;
        RECT 38.730 31.850 39.330 32.300 ;
        RECT 30.130 31.700 34.080 31.850 ;
        RECT 35.380 31.700 39.330 31.850 ;
        RECT 30.130 31.250 30.730 31.700 ;
        RECT 38.730 31.250 39.330 31.700 ;
        RECT 30.130 31.100 34.080 31.250 ;
        RECT 35.380 31.100 39.330 31.250 ;
        RECT 30.130 30.650 30.730 31.100 ;
        RECT 38.730 30.650 39.330 31.100 ;
        RECT 30.130 30.450 34.080 30.650 ;
        RECT 35.380 30.450 39.330 30.650 ;
        RECT 39.780 30.450 39.930 38.000 ;
        RECT 40.380 30.450 40.530 38.000 ;
        RECT 40.980 30.450 41.130 38.000 ;
        RECT 41.580 30.450 41.730 38.000 ;
        RECT 42.180 30.450 42.330 38.000 ;
        RECT 42.780 35.150 42.930 38.000 ;
        RECT 43.530 35.600 45.930 38.800 ;
        RECT 49.280 38.650 50.730 38.950 ;
        RECT 46.530 38.450 50.730 38.650 ;
        RECT 58.730 38.950 70.730 39.800 ;
        RECT 58.730 38.900 69.130 38.950 ;
        RECT 58.730 38.650 60.180 38.900 ;
        RECT 60.330 38.800 69.130 38.900 ;
        RECT 58.730 38.450 62.930 38.650 ;
        RECT 46.530 38.300 54.080 38.450 ;
        RECT 55.430 38.300 62.930 38.450 ;
        RECT 46.530 38.000 50.730 38.300 ;
        RECT 46.530 35.150 46.680 38.000 ;
        RECT 47.130 30.450 47.280 38.000 ;
        RECT 47.730 30.450 47.880 38.000 ;
        RECT 48.330 30.450 48.480 38.000 ;
        RECT 48.930 30.450 49.080 38.000 ;
        RECT 49.530 30.450 49.680 38.000 ;
        RECT 50.130 37.850 50.730 38.000 ;
        RECT 58.730 38.000 62.930 38.300 ;
        RECT 58.730 37.850 59.330 38.000 ;
        RECT 50.130 37.700 54.080 37.850 ;
        RECT 55.380 37.700 59.330 37.850 ;
        RECT 50.130 37.250 50.730 37.700 ;
        RECT 58.730 37.250 59.330 37.700 ;
        RECT 50.130 37.100 54.080 37.250 ;
        RECT 55.380 37.100 59.330 37.250 ;
        RECT 50.130 36.650 50.730 37.100 ;
        RECT 58.730 36.650 59.330 37.100 ;
        RECT 50.130 36.500 54.080 36.650 ;
        RECT 55.380 36.500 59.330 36.650 ;
        RECT 50.130 36.050 50.730 36.500 ;
        RECT 58.730 36.050 59.330 36.500 ;
        RECT 50.130 35.900 54.080 36.050 ;
        RECT 55.380 35.900 59.330 36.050 ;
        RECT 50.130 35.450 50.730 35.900 ;
        RECT 58.730 35.450 59.330 35.900 ;
        RECT 50.130 35.300 54.080 35.450 ;
        RECT 55.380 35.300 59.330 35.450 ;
        RECT 50.130 34.850 50.730 35.300 ;
        RECT 58.730 34.850 59.330 35.300 ;
        RECT 50.130 34.700 54.080 34.850 ;
        RECT 55.380 34.700 59.330 34.850 ;
        RECT 50.130 34.250 50.730 34.700 ;
        RECT 58.730 34.250 59.330 34.700 ;
        RECT 50.130 34.100 54.080 34.250 ;
        RECT 55.380 34.100 59.330 34.250 ;
        RECT 50.130 33.650 50.730 34.100 ;
        RECT 58.730 33.650 59.330 34.100 ;
        RECT 50.130 33.500 54.080 33.650 ;
        RECT 55.380 33.500 59.330 33.650 ;
        RECT 50.130 33.050 50.730 33.500 ;
        RECT 58.730 33.050 59.330 33.500 ;
        RECT 50.130 32.900 54.080 33.050 ;
        RECT 55.380 32.900 59.330 33.050 ;
        RECT 50.130 32.450 50.730 32.900 ;
        RECT 58.730 32.450 59.330 32.900 ;
        RECT 50.130 32.300 54.080 32.450 ;
        RECT 55.380 32.300 59.330 32.450 ;
        RECT 50.130 31.850 50.730 32.300 ;
        RECT 58.730 31.850 59.330 32.300 ;
        RECT 50.130 31.700 54.080 31.850 ;
        RECT 55.380 31.700 59.330 31.850 ;
        RECT 50.130 31.250 50.730 31.700 ;
        RECT 58.730 31.250 59.330 31.700 ;
        RECT 50.130 31.100 54.080 31.250 ;
        RECT 55.380 31.100 59.330 31.250 ;
        RECT 50.130 30.650 50.730 31.100 ;
        RECT 58.730 30.650 59.330 31.100 ;
        RECT 50.130 30.450 54.080 30.650 ;
        RECT 55.380 30.450 59.330 30.650 ;
        RECT 59.780 30.450 59.930 38.000 ;
        RECT 60.380 30.450 60.530 38.000 ;
        RECT 60.980 30.450 61.130 38.000 ;
        RECT 61.580 30.450 61.730 38.000 ;
        RECT 62.180 30.450 62.330 38.000 ;
        RECT 62.780 35.150 62.930 38.000 ;
        RECT 63.530 35.600 65.930 38.800 ;
        RECT 69.280 38.650 70.730 38.950 ;
        RECT 66.530 38.450 70.730 38.650 ;
        RECT 78.730 38.950 90.730 39.800 ;
        RECT 78.730 38.900 89.130 38.950 ;
        RECT 78.730 38.650 80.180 38.900 ;
        RECT 80.330 38.800 89.130 38.900 ;
        RECT 78.730 38.450 82.930 38.650 ;
        RECT 66.530 38.300 74.080 38.450 ;
        RECT 75.430 38.300 82.930 38.450 ;
        RECT 66.530 38.000 70.730 38.300 ;
        RECT 66.530 35.150 66.680 38.000 ;
        RECT 67.130 30.450 67.280 38.000 ;
        RECT 67.730 30.450 67.880 38.000 ;
        RECT 68.330 30.450 68.480 38.000 ;
        RECT 68.930 30.450 69.080 38.000 ;
        RECT 69.530 30.450 69.680 38.000 ;
        RECT 70.130 37.850 70.730 38.000 ;
        RECT 78.730 38.000 82.930 38.300 ;
        RECT 78.730 37.850 79.330 38.000 ;
        RECT 70.130 37.700 74.080 37.850 ;
        RECT 75.380 37.700 79.330 37.850 ;
        RECT 70.130 37.250 70.730 37.700 ;
        RECT 78.730 37.250 79.330 37.700 ;
        RECT 70.130 37.100 74.080 37.250 ;
        RECT 75.380 37.100 79.330 37.250 ;
        RECT 70.130 36.650 70.730 37.100 ;
        RECT 78.730 36.650 79.330 37.100 ;
        RECT 70.130 36.500 74.080 36.650 ;
        RECT 75.380 36.500 79.330 36.650 ;
        RECT 70.130 36.050 70.730 36.500 ;
        RECT 78.730 36.050 79.330 36.500 ;
        RECT 70.130 35.900 74.080 36.050 ;
        RECT 75.380 35.900 79.330 36.050 ;
        RECT 70.130 35.450 70.730 35.900 ;
        RECT 78.730 35.450 79.330 35.900 ;
        RECT 70.130 35.300 74.080 35.450 ;
        RECT 75.380 35.300 79.330 35.450 ;
        RECT 70.130 34.850 70.730 35.300 ;
        RECT 78.730 34.850 79.330 35.300 ;
        RECT 70.130 34.700 74.080 34.850 ;
        RECT 75.380 34.700 79.330 34.850 ;
        RECT 70.130 34.250 70.730 34.700 ;
        RECT 78.730 34.250 79.330 34.700 ;
        RECT 70.130 34.100 74.080 34.250 ;
        RECT 75.380 34.100 79.330 34.250 ;
        RECT 70.130 33.650 70.730 34.100 ;
        RECT 78.730 33.650 79.330 34.100 ;
        RECT 70.130 33.500 74.080 33.650 ;
        RECT 75.380 33.500 79.330 33.650 ;
        RECT 70.130 33.050 70.730 33.500 ;
        RECT 78.730 33.050 79.330 33.500 ;
        RECT 70.130 32.900 74.080 33.050 ;
        RECT 75.380 32.900 79.330 33.050 ;
        RECT 70.130 32.450 70.730 32.900 ;
        RECT 78.730 32.450 79.330 32.900 ;
        RECT 70.130 32.300 74.080 32.450 ;
        RECT 75.380 32.300 79.330 32.450 ;
        RECT 70.130 31.850 70.730 32.300 ;
        RECT 78.730 31.850 79.330 32.300 ;
        RECT 70.130 31.700 74.080 31.850 ;
        RECT 75.380 31.700 79.330 31.850 ;
        RECT 70.130 31.250 70.730 31.700 ;
        RECT 78.730 31.250 79.330 31.700 ;
        RECT 70.130 31.100 74.080 31.250 ;
        RECT 75.380 31.100 79.330 31.250 ;
        RECT 70.130 30.650 70.730 31.100 ;
        RECT 78.730 30.650 79.330 31.100 ;
        RECT 70.130 30.450 74.080 30.650 ;
        RECT 75.380 30.450 79.330 30.650 ;
        RECT 79.780 30.450 79.930 38.000 ;
        RECT 80.380 30.450 80.530 38.000 ;
        RECT 80.980 30.450 81.130 38.000 ;
        RECT 81.580 30.450 81.730 38.000 ;
        RECT 82.180 30.450 82.330 38.000 ;
        RECT 82.780 35.150 82.930 38.000 ;
        RECT 83.530 35.600 85.930 38.800 ;
        RECT 89.280 38.650 90.730 38.950 ;
        RECT 86.530 38.450 90.730 38.650 ;
        RECT 98.730 38.900 104.730 39.800 ;
        RECT 98.730 38.650 100.180 38.900 ;
        RECT 100.330 38.800 104.730 38.900 ;
        RECT 98.730 38.450 102.930 38.650 ;
        RECT 86.530 38.300 94.080 38.450 ;
        RECT 95.430 38.300 102.930 38.450 ;
        RECT 86.530 38.000 90.730 38.300 ;
        RECT 86.530 35.150 86.680 38.000 ;
        RECT 87.130 30.450 87.280 38.000 ;
        RECT 87.730 30.450 87.880 38.000 ;
        RECT 88.330 30.450 88.480 38.000 ;
        RECT 88.930 30.450 89.080 38.000 ;
        RECT 89.530 30.450 89.680 38.000 ;
        RECT 90.130 37.850 90.730 38.000 ;
        RECT 98.730 38.000 102.930 38.300 ;
        RECT 98.730 37.850 99.330 38.000 ;
        RECT 90.130 37.700 94.080 37.850 ;
        RECT 95.380 37.700 99.330 37.850 ;
        RECT 90.130 37.250 90.730 37.700 ;
        RECT 98.730 37.250 99.330 37.700 ;
        RECT 90.130 37.100 94.080 37.250 ;
        RECT 95.380 37.100 99.330 37.250 ;
        RECT 90.130 36.650 90.730 37.100 ;
        RECT 98.730 36.650 99.330 37.100 ;
        RECT 90.130 36.500 94.080 36.650 ;
        RECT 95.380 36.500 99.330 36.650 ;
        RECT 90.130 36.050 90.730 36.500 ;
        RECT 98.730 36.050 99.330 36.500 ;
        RECT 90.130 35.900 94.080 36.050 ;
        RECT 95.380 35.900 99.330 36.050 ;
        RECT 90.130 35.450 90.730 35.900 ;
        RECT 98.730 35.450 99.330 35.900 ;
        RECT 90.130 35.300 94.080 35.450 ;
        RECT 95.380 35.300 99.330 35.450 ;
        RECT 90.130 34.850 90.730 35.300 ;
        RECT 98.730 34.850 99.330 35.300 ;
        RECT 90.130 34.700 94.080 34.850 ;
        RECT 95.380 34.700 99.330 34.850 ;
        RECT 90.130 34.250 90.730 34.700 ;
        RECT 98.730 34.250 99.330 34.700 ;
        RECT 90.130 34.100 94.080 34.250 ;
        RECT 95.380 34.100 99.330 34.250 ;
        RECT 90.130 33.650 90.730 34.100 ;
        RECT 98.730 33.650 99.330 34.100 ;
        RECT 90.130 33.500 94.080 33.650 ;
        RECT 95.380 33.500 99.330 33.650 ;
        RECT 90.130 33.050 90.730 33.500 ;
        RECT 98.730 33.050 99.330 33.500 ;
        RECT 90.130 32.900 94.080 33.050 ;
        RECT 95.380 32.900 99.330 33.050 ;
        RECT 90.130 32.450 90.730 32.900 ;
        RECT 98.730 32.450 99.330 32.900 ;
        RECT 90.130 32.300 94.080 32.450 ;
        RECT 95.380 32.300 99.330 32.450 ;
        RECT 90.130 31.850 90.730 32.300 ;
        RECT 98.730 31.850 99.330 32.300 ;
        RECT 90.130 31.700 94.080 31.850 ;
        RECT 95.380 31.700 99.330 31.850 ;
        RECT 90.130 31.250 90.730 31.700 ;
        RECT 98.730 31.250 99.330 31.700 ;
        RECT 90.130 31.100 94.080 31.250 ;
        RECT 95.380 31.100 99.330 31.250 ;
        RECT 90.130 30.650 90.730 31.100 ;
        RECT 98.730 30.650 99.330 31.100 ;
        RECT 90.130 30.450 94.080 30.650 ;
        RECT 95.380 30.450 99.330 30.650 ;
        RECT 99.780 30.450 99.930 38.000 ;
        RECT 100.380 30.450 100.530 38.000 ;
        RECT 100.980 30.450 101.130 38.000 ;
        RECT 101.580 30.450 101.730 38.000 ;
        RECT 102.180 30.450 102.330 38.000 ;
        RECT 102.780 35.150 102.930 38.000 ;
        RECT 103.530 37.310 104.730 38.800 ;
        RECT 103.530 36.035 107.135 37.310 ;
        RECT 103.530 35.600 104.730 36.035 ;
        RECT 2.315 24.450 4.315 26.745 ;
        RECT 4.730 23.650 5.930 24.400 ;
        RECT 2.315 22.375 5.930 23.650 ;
        RECT 4.730 21.200 5.930 22.375 ;
        RECT 6.530 22.000 6.680 24.900 ;
        RECT 7.130 22.000 7.280 29.550 ;
        RECT 7.730 22.000 7.880 29.550 ;
        RECT 8.330 22.000 8.480 29.550 ;
        RECT 8.930 22.000 9.080 29.550 ;
        RECT 9.530 22.000 9.680 29.550 ;
        RECT 10.130 29.350 14.080 29.550 ;
        RECT 15.380 29.350 19.330 29.550 ;
        RECT 10.130 28.900 10.730 29.350 ;
        RECT 18.730 28.900 19.330 29.350 ;
        RECT 10.130 28.750 14.080 28.900 ;
        RECT 15.380 28.750 19.330 28.900 ;
        RECT 10.130 28.300 10.730 28.750 ;
        RECT 18.730 28.300 19.330 28.750 ;
        RECT 10.130 28.150 14.080 28.300 ;
        RECT 15.380 28.150 19.330 28.300 ;
        RECT 10.130 27.700 10.730 28.150 ;
        RECT 18.730 27.700 19.330 28.150 ;
        RECT 10.130 27.550 14.080 27.700 ;
        RECT 15.380 27.550 19.330 27.700 ;
        RECT 10.130 27.100 10.730 27.550 ;
        RECT 18.730 27.100 19.330 27.550 ;
        RECT 10.130 26.950 14.080 27.100 ;
        RECT 15.380 26.950 19.330 27.100 ;
        RECT 10.130 26.500 10.730 26.950 ;
        RECT 18.730 26.500 19.330 26.950 ;
        RECT 10.130 26.350 14.080 26.500 ;
        RECT 15.380 26.350 19.330 26.500 ;
        RECT 10.130 25.900 10.730 26.350 ;
        RECT 18.730 25.900 19.330 26.350 ;
        RECT 10.130 25.750 14.080 25.900 ;
        RECT 15.380 25.750 19.330 25.900 ;
        RECT 10.130 25.300 10.730 25.750 ;
        RECT 18.730 25.300 19.330 25.750 ;
        RECT 10.130 25.150 14.080 25.300 ;
        RECT 15.380 25.150 19.330 25.300 ;
        RECT 10.130 24.700 10.730 25.150 ;
        RECT 18.730 24.700 19.330 25.150 ;
        RECT 10.130 24.550 14.080 24.700 ;
        RECT 15.380 24.550 19.330 24.700 ;
        RECT 10.130 24.100 10.730 24.550 ;
        RECT 18.730 24.100 19.330 24.550 ;
        RECT 10.130 23.950 14.080 24.100 ;
        RECT 15.380 23.950 19.330 24.100 ;
        RECT 10.130 23.500 10.730 23.950 ;
        RECT 18.730 23.500 19.330 23.950 ;
        RECT 10.130 23.350 14.080 23.500 ;
        RECT 15.380 23.350 19.330 23.500 ;
        RECT 10.130 22.900 10.730 23.350 ;
        RECT 18.730 22.900 19.330 23.350 ;
        RECT 10.130 22.750 14.080 22.900 ;
        RECT 15.380 22.750 19.330 22.900 ;
        RECT 10.130 22.300 10.730 22.750 ;
        RECT 18.730 22.300 19.330 22.750 ;
        RECT 10.130 22.150 14.080 22.300 ;
        RECT 15.380 22.150 19.330 22.300 ;
        RECT 10.130 22.000 10.730 22.150 ;
        RECT 6.530 21.700 10.730 22.000 ;
        RECT 18.730 22.000 19.330 22.150 ;
        RECT 19.780 22.000 19.930 29.550 ;
        RECT 20.380 22.000 20.530 29.550 ;
        RECT 20.980 22.000 21.130 29.550 ;
        RECT 21.580 22.000 21.730 29.550 ;
        RECT 22.180 22.000 22.330 29.550 ;
        RECT 22.780 22.000 22.930 24.900 ;
        RECT 18.730 21.700 22.930 22.000 ;
        RECT 6.530 21.550 14.080 21.700 ;
        RECT 15.380 21.550 22.930 21.700 ;
        RECT 6.530 21.350 10.730 21.550 ;
        RECT 4.730 21.050 9.130 21.200 ;
        RECT 9.280 21.050 10.730 21.350 ;
        RECT 4.730 20.150 10.730 21.050 ;
        RECT 18.730 21.350 22.930 21.550 ;
        RECT 18.730 21.050 20.180 21.350 ;
        RECT 23.530 21.200 25.930 24.400 ;
        RECT 26.530 22.000 26.680 24.900 ;
        RECT 27.130 22.000 27.280 29.550 ;
        RECT 27.730 22.000 27.880 29.550 ;
        RECT 28.330 22.000 28.480 29.550 ;
        RECT 28.930 22.000 29.080 29.550 ;
        RECT 29.530 22.000 29.680 29.550 ;
        RECT 30.130 29.350 34.080 29.550 ;
        RECT 35.380 29.350 39.330 29.550 ;
        RECT 30.130 28.900 30.730 29.350 ;
        RECT 38.730 28.900 39.330 29.350 ;
        RECT 30.130 28.750 34.080 28.900 ;
        RECT 35.380 28.750 39.330 28.900 ;
        RECT 30.130 28.300 30.730 28.750 ;
        RECT 38.730 28.300 39.330 28.750 ;
        RECT 30.130 28.150 34.080 28.300 ;
        RECT 35.380 28.150 39.330 28.300 ;
        RECT 30.130 27.700 30.730 28.150 ;
        RECT 38.730 27.700 39.330 28.150 ;
        RECT 30.130 27.550 34.080 27.700 ;
        RECT 35.380 27.550 39.330 27.700 ;
        RECT 30.130 27.100 30.730 27.550 ;
        RECT 38.730 27.100 39.330 27.550 ;
        RECT 30.130 26.950 34.080 27.100 ;
        RECT 35.380 26.950 39.330 27.100 ;
        RECT 30.130 26.500 30.730 26.950 ;
        RECT 38.730 26.500 39.330 26.950 ;
        RECT 30.130 26.350 34.080 26.500 ;
        RECT 35.380 26.350 39.330 26.500 ;
        RECT 30.130 25.900 30.730 26.350 ;
        RECT 38.730 25.900 39.330 26.350 ;
        RECT 30.130 25.750 34.080 25.900 ;
        RECT 35.380 25.750 39.330 25.900 ;
        RECT 30.130 25.300 30.730 25.750 ;
        RECT 38.730 25.300 39.330 25.750 ;
        RECT 30.130 25.150 34.080 25.300 ;
        RECT 35.380 25.150 39.330 25.300 ;
        RECT 30.130 24.700 30.730 25.150 ;
        RECT 38.730 24.700 39.330 25.150 ;
        RECT 30.130 24.550 34.080 24.700 ;
        RECT 35.380 24.550 39.330 24.700 ;
        RECT 30.130 24.100 30.730 24.550 ;
        RECT 38.730 24.100 39.330 24.550 ;
        RECT 30.130 23.950 34.080 24.100 ;
        RECT 35.380 23.950 39.330 24.100 ;
        RECT 30.130 23.500 30.730 23.950 ;
        RECT 38.730 23.500 39.330 23.950 ;
        RECT 30.130 23.350 34.080 23.500 ;
        RECT 35.380 23.350 39.330 23.500 ;
        RECT 30.130 22.900 30.730 23.350 ;
        RECT 38.730 22.900 39.330 23.350 ;
        RECT 30.130 22.750 34.080 22.900 ;
        RECT 35.380 22.750 39.330 22.900 ;
        RECT 30.130 22.300 30.730 22.750 ;
        RECT 38.730 22.300 39.330 22.750 ;
        RECT 30.130 22.150 34.080 22.300 ;
        RECT 35.380 22.150 39.330 22.300 ;
        RECT 30.130 22.000 30.730 22.150 ;
        RECT 26.530 21.700 30.730 22.000 ;
        RECT 38.730 22.000 39.330 22.150 ;
        RECT 39.780 22.000 39.930 29.550 ;
        RECT 40.380 22.000 40.530 29.550 ;
        RECT 40.980 22.000 41.130 29.550 ;
        RECT 41.580 22.000 41.730 29.550 ;
        RECT 42.180 22.000 42.330 29.550 ;
        RECT 42.780 22.000 42.930 24.900 ;
        RECT 38.730 21.700 42.930 22.000 ;
        RECT 26.530 21.550 34.080 21.700 ;
        RECT 35.380 21.550 42.930 21.700 ;
        RECT 26.530 21.350 30.730 21.550 ;
        RECT 20.330 21.050 29.130 21.200 ;
        RECT 29.280 21.050 30.730 21.350 ;
        RECT 18.730 20.150 30.730 21.050 ;
        RECT 38.730 21.350 42.930 21.550 ;
        RECT 38.730 21.050 40.180 21.350 ;
        RECT 43.530 21.200 45.930 24.400 ;
        RECT 46.530 22.000 46.680 24.900 ;
        RECT 47.130 22.000 47.280 29.550 ;
        RECT 47.730 22.000 47.880 29.550 ;
        RECT 48.330 22.000 48.480 29.550 ;
        RECT 48.930 22.000 49.080 29.550 ;
        RECT 49.530 22.000 49.680 29.550 ;
        RECT 50.130 29.350 54.080 29.550 ;
        RECT 55.380 29.350 59.330 29.550 ;
        RECT 50.130 28.900 50.730 29.350 ;
        RECT 58.730 28.900 59.330 29.350 ;
        RECT 50.130 28.750 54.080 28.900 ;
        RECT 55.380 28.750 59.330 28.900 ;
        RECT 50.130 28.300 50.730 28.750 ;
        RECT 58.730 28.300 59.330 28.750 ;
        RECT 50.130 28.150 54.080 28.300 ;
        RECT 55.380 28.150 59.330 28.300 ;
        RECT 50.130 27.700 50.730 28.150 ;
        RECT 58.730 27.700 59.330 28.150 ;
        RECT 50.130 27.550 54.080 27.700 ;
        RECT 55.380 27.550 59.330 27.700 ;
        RECT 50.130 27.100 50.730 27.550 ;
        RECT 58.730 27.100 59.330 27.550 ;
        RECT 50.130 26.950 54.080 27.100 ;
        RECT 55.380 26.950 59.330 27.100 ;
        RECT 50.130 26.500 50.730 26.950 ;
        RECT 58.730 26.500 59.330 26.950 ;
        RECT 50.130 26.350 54.080 26.500 ;
        RECT 55.380 26.350 59.330 26.500 ;
        RECT 50.130 25.900 50.730 26.350 ;
        RECT 58.730 25.900 59.330 26.350 ;
        RECT 50.130 25.750 54.080 25.900 ;
        RECT 55.380 25.750 59.330 25.900 ;
        RECT 50.130 25.300 50.730 25.750 ;
        RECT 58.730 25.300 59.330 25.750 ;
        RECT 50.130 25.150 54.080 25.300 ;
        RECT 55.380 25.150 59.330 25.300 ;
        RECT 50.130 24.700 50.730 25.150 ;
        RECT 58.730 24.700 59.330 25.150 ;
        RECT 50.130 24.550 54.080 24.700 ;
        RECT 55.380 24.550 59.330 24.700 ;
        RECT 50.130 24.100 50.730 24.550 ;
        RECT 58.730 24.100 59.330 24.550 ;
        RECT 50.130 23.950 54.080 24.100 ;
        RECT 55.380 23.950 59.330 24.100 ;
        RECT 50.130 23.500 50.730 23.950 ;
        RECT 58.730 23.500 59.330 23.950 ;
        RECT 50.130 23.350 54.080 23.500 ;
        RECT 55.380 23.350 59.330 23.500 ;
        RECT 50.130 22.900 50.730 23.350 ;
        RECT 58.730 22.900 59.330 23.350 ;
        RECT 50.130 22.750 54.080 22.900 ;
        RECT 55.380 22.750 59.330 22.900 ;
        RECT 50.130 22.300 50.730 22.750 ;
        RECT 58.730 22.300 59.330 22.750 ;
        RECT 50.130 22.150 54.080 22.300 ;
        RECT 55.380 22.150 59.330 22.300 ;
        RECT 50.130 22.000 50.730 22.150 ;
        RECT 46.530 21.700 50.730 22.000 ;
        RECT 58.730 22.000 59.330 22.150 ;
        RECT 59.780 22.000 59.930 29.550 ;
        RECT 60.380 22.000 60.530 29.550 ;
        RECT 60.980 22.000 61.130 29.550 ;
        RECT 61.580 22.000 61.730 29.550 ;
        RECT 62.180 22.000 62.330 29.550 ;
        RECT 62.780 22.000 62.930 24.900 ;
        RECT 58.730 21.700 62.930 22.000 ;
        RECT 46.530 21.550 54.080 21.700 ;
        RECT 55.380 21.550 62.930 21.700 ;
        RECT 46.530 21.350 50.730 21.550 ;
        RECT 40.330 21.050 49.130 21.200 ;
        RECT 49.280 21.050 50.730 21.350 ;
        RECT 38.730 20.150 50.730 21.050 ;
        RECT 58.730 21.350 62.930 21.550 ;
        RECT 58.730 21.050 60.180 21.350 ;
        RECT 63.530 21.200 65.930 24.400 ;
        RECT 66.530 22.000 66.680 24.900 ;
        RECT 67.130 22.000 67.280 29.550 ;
        RECT 67.730 22.000 67.880 29.550 ;
        RECT 68.330 22.000 68.480 29.550 ;
        RECT 68.930 22.000 69.080 29.550 ;
        RECT 69.530 22.000 69.680 29.550 ;
        RECT 70.130 29.350 74.080 29.550 ;
        RECT 75.380 29.350 79.330 29.550 ;
        RECT 70.130 28.900 70.730 29.350 ;
        RECT 78.730 28.900 79.330 29.350 ;
        RECT 70.130 28.750 74.080 28.900 ;
        RECT 75.380 28.750 79.330 28.900 ;
        RECT 70.130 28.300 70.730 28.750 ;
        RECT 78.730 28.300 79.330 28.750 ;
        RECT 70.130 28.150 74.080 28.300 ;
        RECT 75.380 28.150 79.330 28.300 ;
        RECT 70.130 27.700 70.730 28.150 ;
        RECT 78.730 27.700 79.330 28.150 ;
        RECT 70.130 27.550 74.080 27.700 ;
        RECT 75.380 27.550 79.330 27.700 ;
        RECT 70.130 27.100 70.730 27.550 ;
        RECT 78.730 27.100 79.330 27.550 ;
        RECT 70.130 26.950 74.080 27.100 ;
        RECT 75.380 26.950 79.330 27.100 ;
        RECT 70.130 26.500 70.730 26.950 ;
        RECT 78.730 26.500 79.330 26.950 ;
        RECT 70.130 26.350 74.080 26.500 ;
        RECT 75.380 26.350 79.330 26.500 ;
        RECT 70.130 25.900 70.730 26.350 ;
        RECT 78.730 25.900 79.330 26.350 ;
        RECT 70.130 25.750 74.080 25.900 ;
        RECT 75.380 25.750 79.330 25.900 ;
        RECT 70.130 25.300 70.730 25.750 ;
        RECT 78.730 25.300 79.330 25.750 ;
        RECT 70.130 25.150 74.080 25.300 ;
        RECT 75.380 25.150 79.330 25.300 ;
        RECT 70.130 24.700 70.730 25.150 ;
        RECT 78.730 24.700 79.330 25.150 ;
        RECT 70.130 24.550 74.080 24.700 ;
        RECT 75.380 24.550 79.330 24.700 ;
        RECT 70.130 24.100 70.730 24.550 ;
        RECT 78.730 24.100 79.330 24.550 ;
        RECT 70.130 23.950 74.080 24.100 ;
        RECT 75.380 23.950 79.330 24.100 ;
        RECT 70.130 23.500 70.730 23.950 ;
        RECT 78.730 23.500 79.330 23.950 ;
        RECT 70.130 23.350 74.080 23.500 ;
        RECT 75.380 23.350 79.330 23.500 ;
        RECT 70.130 22.900 70.730 23.350 ;
        RECT 78.730 22.900 79.330 23.350 ;
        RECT 70.130 22.750 74.080 22.900 ;
        RECT 75.380 22.750 79.330 22.900 ;
        RECT 70.130 22.300 70.730 22.750 ;
        RECT 78.730 22.300 79.330 22.750 ;
        RECT 70.130 22.150 74.080 22.300 ;
        RECT 75.380 22.150 79.330 22.300 ;
        RECT 70.130 22.000 70.730 22.150 ;
        RECT 66.530 21.700 70.730 22.000 ;
        RECT 78.730 22.000 79.330 22.150 ;
        RECT 79.780 22.000 79.930 29.550 ;
        RECT 80.380 22.000 80.530 29.550 ;
        RECT 80.980 22.000 81.130 29.550 ;
        RECT 81.580 22.000 81.730 29.550 ;
        RECT 82.180 22.000 82.330 29.550 ;
        RECT 82.780 22.000 82.930 24.900 ;
        RECT 78.730 21.700 82.930 22.000 ;
        RECT 66.530 21.550 74.080 21.700 ;
        RECT 75.380 21.550 82.930 21.700 ;
        RECT 66.530 21.350 70.730 21.550 ;
        RECT 60.330 21.050 69.130 21.200 ;
        RECT 69.280 21.050 70.730 21.350 ;
        RECT 58.730 20.150 70.730 21.050 ;
        RECT 78.730 21.350 82.930 21.550 ;
        RECT 78.730 21.050 80.180 21.350 ;
        RECT 83.530 21.200 85.930 24.400 ;
        RECT 86.530 22.000 86.680 24.900 ;
        RECT 87.130 22.000 87.280 29.550 ;
        RECT 87.730 22.000 87.880 29.550 ;
        RECT 88.330 22.000 88.480 29.550 ;
        RECT 88.930 22.000 89.080 29.550 ;
        RECT 89.530 22.000 89.680 29.550 ;
        RECT 90.130 29.350 94.080 29.550 ;
        RECT 95.380 29.350 99.330 29.550 ;
        RECT 90.130 28.900 90.730 29.350 ;
        RECT 98.730 28.900 99.330 29.350 ;
        RECT 90.130 28.750 94.080 28.900 ;
        RECT 95.380 28.750 99.330 28.900 ;
        RECT 90.130 28.300 90.730 28.750 ;
        RECT 98.730 28.300 99.330 28.750 ;
        RECT 90.130 28.150 94.080 28.300 ;
        RECT 95.380 28.150 99.330 28.300 ;
        RECT 90.130 27.700 90.730 28.150 ;
        RECT 98.730 27.700 99.330 28.150 ;
        RECT 90.130 27.550 94.080 27.700 ;
        RECT 95.380 27.550 99.330 27.700 ;
        RECT 90.130 27.100 90.730 27.550 ;
        RECT 98.730 27.100 99.330 27.550 ;
        RECT 90.130 26.950 94.080 27.100 ;
        RECT 95.380 26.950 99.330 27.100 ;
        RECT 90.130 26.500 90.730 26.950 ;
        RECT 98.730 26.500 99.330 26.950 ;
        RECT 90.130 26.350 94.080 26.500 ;
        RECT 95.380 26.350 99.330 26.500 ;
        RECT 90.130 25.900 90.730 26.350 ;
        RECT 98.730 25.900 99.330 26.350 ;
        RECT 90.130 25.750 94.080 25.900 ;
        RECT 95.380 25.750 99.330 25.900 ;
        RECT 90.130 25.300 90.730 25.750 ;
        RECT 98.730 25.300 99.330 25.750 ;
        RECT 90.130 25.150 94.080 25.300 ;
        RECT 95.380 25.150 99.330 25.300 ;
        RECT 90.130 24.700 90.730 25.150 ;
        RECT 98.730 24.700 99.330 25.150 ;
        RECT 90.130 24.550 94.080 24.700 ;
        RECT 95.380 24.550 99.330 24.700 ;
        RECT 90.130 24.100 90.730 24.550 ;
        RECT 98.730 24.100 99.330 24.550 ;
        RECT 90.130 23.950 94.080 24.100 ;
        RECT 95.380 23.950 99.330 24.100 ;
        RECT 90.130 23.500 90.730 23.950 ;
        RECT 98.730 23.500 99.330 23.950 ;
        RECT 90.130 23.350 94.080 23.500 ;
        RECT 95.380 23.350 99.330 23.500 ;
        RECT 90.130 22.900 90.730 23.350 ;
        RECT 98.730 22.900 99.330 23.350 ;
        RECT 90.130 22.750 94.080 22.900 ;
        RECT 95.380 22.750 99.330 22.900 ;
        RECT 90.130 22.300 90.730 22.750 ;
        RECT 98.730 22.300 99.330 22.750 ;
        RECT 90.130 22.150 94.080 22.300 ;
        RECT 95.380 22.150 99.330 22.300 ;
        RECT 90.130 22.000 90.730 22.150 ;
        RECT 86.530 21.700 90.730 22.000 ;
        RECT 98.730 22.000 99.330 22.150 ;
        RECT 99.780 22.000 99.930 29.550 ;
        RECT 100.380 22.000 100.530 29.550 ;
        RECT 100.980 22.000 101.130 29.550 ;
        RECT 101.580 22.000 101.730 29.550 ;
        RECT 102.180 22.000 102.330 29.550 ;
        RECT 102.780 22.000 102.930 24.900 ;
        RECT 98.730 21.700 102.930 22.000 ;
        RECT 86.530 21.550 94.080 21.700 ;
        RECT 95.380 21.550 102.930 21.700 ;
        RECT 86.530 21.350 90.730 21.550 ;
        RECT 80.330 21.050 89.130 21.200 ;
        RECT 89.280 21.050 90.730 21.350 ;
        RECT 78.730 20.150 90.730 21.050 ;
        RECT 98.730 21.350 102.930 21.550 ;
        RECT 103.530 23.095 104.730 24.400 ;
        RECT 103.530 21.820 107.140 23.095 ;
        RECT 98.730 21.050 100.180 21.350 ;
        RECT 103.530 21.200 104.730 21.820 ;
        RECT 100.330 21.050 104.730 21.200 ;
        RECT 98.730 20.150 104.730 21.050 ;
        RECT 4.730 19.850 9.130 20.150 ;
        RECT 20.330 19.850 29.130 20.150 ;
        RECT 40.330 19.850 49.130 20.150 ;
        RECT 60.330 19.850 69.130 20.150 ;
        RECT 80.330 19.850 89.130 20.150 ;
        RECT 4.730 18.950 10.730 19.850 ;
        RECT 20.330 19.800 30.730 19.850 ;
        RECT 40.330 19.800 50.730 19.850 ;
        RECT 60.330 19.800 70.730 19.850 ;
        RECT 80.330 19.800 90.730 19.850 ;
        RECT 100.330 19.800 104.730 20.150 ;
        RECT 4.730 18.800 9.130 18.950 ;
        RECT 4.730 17.765 5.930 18.800 ;
        RECT 9.280 18.650 10.730 18.950 ;
        RECT 2.315 16.490 5.930 17.765 ;
        RECT 4.730 15.600 5.930 16.490 ;
        RECT 6.530 18.450 10.730 18.650 ;
        RECT 18.730 18.950 30.730 19.800 ;
        RECT 18.730 18.900 29.130 18.950 ;
        RECT 18.730 18.650 20.180 18.900 ;
        RECT 20.330 18.800 29.130 18.900 ;
        RECT 18.730 18.450 22.930 18.650 ;
        RECT 6.530 18.300 14.080 18.450 ;
        RECT 15.430 18.300 22.930 18.450 ;
        RECT 6.530 18.000 10.730 18.300 ;
        RECT 2.315 13.255 4.315 15.550 ;
        RECT 6.530 15.150 6.680 18.000 ;
        RECT 7.130 10.450 7.280 18.000 ;
        RECT 7.730 10.450 7.880 18.000 ;
        RECT 8.330 10.450 8.480 18.000 ;
        RECT 8.930 10.450 9.080 18.000 ;
        RECT 9.530 10.450 9.680 18.000 ;
        RECT 10.130 17.850 10.730 18.000 ;
        RECT 18.730 18.000 22.930 18.300 ;
        RECT 18.730 17.850 19.330 18.000 ;
        RECT 10.130 17.700 14.080 17.850 ;
        RECT 15.380 17.700 19.330 17.850 ;
        RECT 10.130 17.250 10.730 17.700 ;
        RECT 18.730 17.250 19.330 17.700 ;
        RECT 10.130 17.100 14.080 17.250 ;
        RECT 15.380 17.100 19.330 17.250 ;
        RECT 10.130 16.650 10.730 17.100 ;
        RECT 18.730 16.650 19.330 17.100 ;
        RECT 10.130 16.500 14.080 16.650 ;
        RECT 15.380 16.500 19.330 16.650 ;
        RECT 10.130 16.050 10.730 16.500 ;
        RECT 18.730 16.050 19.330 16.500 ;
        RECT 10.130 15.900 14.080 16.050 ;
        RECT 15.380 15.900 19.330 16.050 ;
        RECT 10.130 15.450 10.730 15.900 ;
        RECT 18.730 15.450 19.330 15.900 ;
        RECT 10.130 15.300 14.080 15.450 ;
        RECT 15.380 15.300 19.330 15.450 ;
        RECT 10.130 14.850 10.730 15.300 ;
        RECT 18.730 14.850 19.330 15.300 ;
        RECT 10.130 14.700 14.080 14.850 ;
        RECT 15.380 14.700 19.330 14.850 ;
        RECT 10.130 14.250 10.730 14.700 ;
        RECT 18.730 14.250 19.330 14.700 ;
        RECT 10.130 14.100 14.080 14.250 ;
        RECT 15.380 14.100 19.330 14.250 ;
        RECT 10.130 13.650 10.730 14.100 ;
        RECT 18.730 13.650 19.330 14.100 ;
        RECT 10.130 13.500 14.080 13.650 ;
        RECT 15.380 13.500 19.330 13.650 ;
        RECT 10.130 13.050 10.730 13.500 ;
        RECT 18.730 13.050 19.330 13.500 ;
        RECT 10.130 12.900 14.080 13.050 ;
        RECT 15.380 12.900 19.330 13.050 ;
        RECT 10.130 12.450 10.730 12.900 ;
        RECT 18.730 12.450 19.330 12.900 ;
        RECT 10.130 12.300 14.080 12.450 ;
        RECT 15.380 12.300 19.330 12.450 ;
        RECT 10.130 11.850 10.730 12.300 ;
        RECT 18.730 11.850 19.330 12.300 ;
        RECT 10.130 11.700 14.080 11.850 ;
        RECT 15.380 11.700 19.330 11.850 ;
        RECT 10.130 11.250 10.730 11.700 ;
        RECT 18.730 11.250 19.330 11.700 ;
        RECT 10.130 11.100 14.080 11.250 ;
        RECT 15.380 11.100 19.330 11.250 ;
        RECT 10.130 10.650 10.730 11.100 ;
        RECT 18.730 10.650 19.330 11.100 ;
        RECT 10.130 10.450 14.080 10.650 ;
        RECT 15.380 10.450 19.330 10.650 ;
        RECT 19.780 10.450 19.930 18.000 ;
        RECT 20.380 10.450 20.530 18.000 ;
        RECT 20.980 10.450 21.130 18.000 ;
        RECT 21.580 10.450 21.730 18.000 ;
        RECT 22.180 10.450 22.330 18.000 ;
        RECT 22.780 15.150 22.930 18.000 ;
        RECT 23.530 15.600 25.930 18.800 ;
        RECT 29.280 18.650 30.730 18.950 ;
        RECT 26.530 18.450 30.730 18.650 ;
        RECT 38.730 18.950 50.730 19.800 ;
        RECT 38.730 18.900 49.130 18.950 ;
        RECT 38.730 18.650 40.180 18.900 ;
        RECT 40.330 18.800 49.130 18.900 ;
        RECT 38.730 18.450 42.930 18.650 ;
        RECT 26.530 18.300 34.080 18.450 ;
        RECT 35.430 18.300 42.930 18.450 ;
        RECT 26.530 18.000 30.730 18.300 ;
        RECT 26.530 15.150 26.680 18.000 ;
        RECT 27.130 10.450 27.280 18.000 ;
        RECT 27.730 10.450 27.880 18.000 ;
        RECT 28.330 10.450 28.480 18.000 ;
        RECT 28.930 10.450 29.080 18.000 ;
        RECT 29.530 10.450 29.680 18.000 ;
        RECT 30.130 17.850 30.730 18.000 ;
        RECT 38.730 18.000 42.930 18.300 ;
        RECT 38.730 17.850 39.330 18.000 ;
        RECT 30.130 17.700 34.080 17.850 ;
        RECT 35.380 17.700 39.330 17.850 ;
        RECT 30.130 17.250 30.730 17.700 ;
        RECT 38.730 17.250 39.330 17.700 ;
        RECT 30.130 17.100 34.080 17.250 ;
        RECT 35.380 17.100 39.330 17.250 ;
        RECT 30.130 16.650 30.730 17.100 ;
        RECT 38.730 16.650 39.330 17.100 ;
        RECT 30.130 16.500 34.080 16.650 ;
        RECT 35.380 16.500 39.330 16.650 ;
        RECT 30.130 16.050 30.730 16.500 ;
        RECT 38.730 16.050 39.330 16.500 ;
        RECT 30.130 15.900 34.080 16.050 ;
        RECT 35.380 15.900 39.330 16.050 ;
        RECT 30.130 15.450 30.730 15.900 ;
        RECT 38.730 15.450 39.330 15.900 ;
        RECT 30.130 15.300 34.080 15.450 ;
        RECT 35.380 15.300 39.330 15.450 ;
        RECT 30.130 14.850 30.730 15.300 ;
        RECT 38.730 14.850 39.330 15.300 ;
        RECT 30.130 14.700 34.080 14.850 ;
        RECT 35.380 14.700 39.330 14.850 ;
        RECT 30.130 14.250 30.730 14.700 ;
        RECT 38.730 14.250 39.330 14.700 ;
        RECT 30.130 14.100 34.080 14.250 ;
        RECT 35.380 14.100 39.330 14.250 ;
        RECT 30.130 13.650 30.730 14.100 ;
        RECT 38.730 13.650 39.330 14.100 ;
        RECT 30.130 13.500 34.080 13.650 ;
        RECT 35.380 13.500 39.330 13.650 ;
        RECT 30.130 13.050 30.730 13.500 ;
        RECT 38.730 13.050 39.330 13.500 ;
        RECT 30.130 12.900 34.080 13.050 ;
        RECT 35.380 12.900 39.330 13.050 ;
        RECT 30.130 12.450 30.730 12.900 ;
        RECT 38.730 12.450 39.330 12.900 ;
        RECT 30.130 12.300 34.080 12.450 ;
        RECT 35.380 12.300 39.330 12.450 ;
        RECT 30.130 11.850 30.730 12.300 ;
        RECT 38.730 11.850 39.330 12.300 ;
        RECT 30.130 11.700 34.080 11.850 ;
        RECT 35.380 11.700 39.330 11.850 ;
        RECT 30.130 11.250 30.730 11.700 ;
        RECT 38.730 11.250 39.330 11.700 ;
        RECT 30.130 11.100 34.080 11.250 ;
        RECT 35.380 11.100 39.330 11.250 ;
        RECT 30.130 10.650 30.730 11.100 ;
        RECT 38.730 10.650 39.330 11.100 ;
        RECT 30.130 10.450 34.080 10.650 ;
        RECT 35.380 10.450 39.330 10.650 ;
        RECT 39.780 10.450 39.930 18.000 ;
        RECT 40.380 10.450 40.530 18.000 ;
        RECT 40.980 10.450 41.130 18.000 ;
        RECT 41.580 10.450 41.730 18.000 ;
        RECT 42.180 10.450 42.330 18.000 ;
        RECT 42.780 15.150 42.930 18.000 ;
        RECT 43.530 15.600 45.930 18.800 ;
        RECT 49.280 18.650 50.730 18.950 ;
        RECT 46.530 18.450 50.730 18.650 ;
        RECT 58.730 18.950 70.730 19.800 ;
        RECT 58.730 18.900 69.130 18.950 ;
        RECT 58.730 18.650 60.180 18.900 ;
        RECT 60.330 18.800 69.130 18.900 ;
        RECT 58.730 18.450 62.930 18.650 ;
        RECT 46.530 18.300 54.080 18.450 ;
        RECT 55.430 18.300 62.930 18.450 ;
        RECT 46.530 18.000 50.730 18.300 ;
        RECT 46.530 15.150 46.680 18.000 ;
        RECT 47.130 10.450 47.280 18.000 ;
        RECT 47.730 10.450 47.880 18.000 ;
        RECT 48.330 10.450 48.480 18.000 ;
        RECT 48.930 10.450 49.080 18.000 ;
        RECT 49.530 10.450 49.680 18.000 ;
        RECT 50.130 17.850 50.730 18.000 ;
        RECT 58.730 18.000 62.930 18.300 ;
        RECT 58.730 17.850 59.330 18.000 ;
        RECT 50.130 17.700 54.080 17.850 ;
        RECT 55.380 17.700 59.330 17.850 ;
        RECT 50.130 17.250 50.730 17.700 ;
        RECT 58.730 17.250 59.330 17.700 ;
        RECT 50.130 17.100 54.080 17.250 ;
        RECT 55.380 17.100 59.330 17.250 ;
        RECT 50.130 16.650 50.730 17.100 ;
        RECT 58.730 16.650 59.330 17.100 ;
        RECT 50.130 16.500 54.080 16.650 ;
        RECT 55.380 16.500 59.330 16.650 ;
        RECT 50.130 16.050 50.730 16.500 ;
        RECT 58.730 16.050 59.330 16.500 ;
        RECT 50.130 15.900 54.080 16.050 ;
        RECT 55.380 15.900 59.330 16.050 ;
        RECT 50.130 15.450 50.730 15.900 ;
        RECT 58.730 15.450 59.330 15.900 ;
        RECT 50.130 15.300 54.080 15.450 ;
        RECT 55.380 15.300 59.330 15.450 ;
        RECT 50.130 14.850 50.730 15.300 ;
        RECT 58.730 14.850 59.330 15.300 ;
        RECT 50.130 14.700 54.080 14.850 ;
        RECT 55.380 14.700 59.330 14.850 ;
        RECT 50.130 14.250 50.730 14.700 ;
        RECT 58.730 14.250 59.330 14.700 ;
        RECT 50.130 14.100 54.080 14.250 ;
        RECT 55.380 14.100 59.330 14.250 ;
        RECT 50.130 13.650 50.730 14.100 ;
        RECT 58.730 13.650 59.330 14.100 ;
        RECT 50.130 13.500 54.080 13.650 ;
        RECT 55.380 13.500 59.330 13.650 ;
        RECT 50.130 13.050 50.730 13.500 ;
        RECT 58.730 13.050 59.330 13.500 ;
        RECT 50.130 12.900 54.080 13.050 ;
        RECT 55.380 12.900 59.330 13.050 ;
        RECT 50.130 12.450 50.730 12.900 ;
        RECT 58.730 12.450 59.330 12.900 ;
        RECT 50.130 12.300 54.080 12.450 ;
        RECT 55.380 12.300 59.330 12.450 ;
        RECT 50.130 11.850 50.730 12.300 ;
        RECT 58.730 11.850 59.330 12.300 ;
        RECT 50.130 11.700 54.080 11.850 ;
        RECT 55.380 11.700 59.330 11.850 ;
        RECT 50.130 11.250 50.730 11.700 ;
        RECT 58.730 11.250 59.330 11.700 ;
        RECT 50.130 11.100 54.080 11.250 ;
        RECT 55.380 11.100 59.330 11.250 ;
        RECT 50.130 10.650 50.730 11.100 ;
        RECT 58.730 10.650 59.330 11.100 ;
        RECT 50.130 10.450 54.080 10.650 ;
        RECT 55.380 10.450 59.330 10.650 ;
        RECT 59.780 10.450 59.930 18.000 ;
        RECT 60.380 10.450 60.530 18.000 ;
        RECT 60.980 10.450 61.130 18.000 ;
        RECT 61.580 10.450 61.730 18.000 ;
        RECT 62.180 10.450 62.330 18.000 ;
        RECT 62.780 15.150 62.930 18.000 ;
        RECT 63.530 15.600 65.930 18.800 ;
        RECT 69.280 18.650 70.730 18.950 ;
        RECT 66.530 18.450 70.730 18.650 ;
        RECT 78.730 18.950 90.730 19.800 ;
        RECT 78.730 18.900 89.130 18.950 ;
        RECT 78.730 18.650 80.180 18.900 ;
        RECT 80.330 18.800 89.130 18.900 ;
        RECT 78.730 18.450 82.930 18.650 ;
        RECT 66.530 18.300 74.080 18.450 ;
        RECT 75.430 18.300 82.930 18.450 ;
        RECT 66.530 18.000 70.730 18.300 ;
        RECT 66.530 15.150 66.680 18.000 ;
        RECT 67.130 10.450 67.280 18.000 ;
        RECT 67.730 10.450 67.880 18.000 ;
        RECT 68.330 10.450 68.480 18.000 ;
        RECT 68.930 10.450 69.080 18.000 ;
        RECT 69.530 10.450 69.680 18.000 ;
        RECT 70.130 17.850 70.730 18.000 ;
        RECT 78.730 18.000 82.930 18.300 ;
        RECT 78.730 17.850 79.330 18.000 ;
        RECT 70.130 17.700 74.080 17.850 ;
        RECT 75.380 17.700 79.330 17.850 ;
        RECT 70.130 17.250 70.730 17.700 ;
        RECT 78.730 17.250 79.330 17.700 ;
        RECT 70.130 17.100 74.080 17.250 ;
        RECT 75.380 17.100 79.330 17.250 ;
        RECT 70.130 16.650 70.730 17.100 ;
        RECT 78.730 16.650 79.330 17.100 ;
        RECT 70.130 16.500 74.080 16.650 ;
        RECT 75.380 16.500 79.330 16.650 ;
        RECT 70.130 16.050 70.730 16.500 ;
        RECT 78.730 16.050 79.330 16.500 ;
        RECT 70.130 15.900 74.080 16.050 ;
        RECT 75.380 15.900 79.330 16.050 ;
        RECT 70.130 15.450 70.730 15.900 ;
        RECT 78.730 15.450 79.330 15.900 ;
        RECT 70.130 15.300 74.080 15.450 ;
        RECT 75.380 15.300 79.330 15.450 ;
        RECT 70.130 14.850 70.730 15.300 ;
        RECT 78.730 14.850 79.330 15.300 ;
        RECT 70.130 14.700 74.080 14.850 ;
        RECT 75.380 14.700 79.330 14.850 ;
        RECT 70.130 14.250 70.730 14.700 ;
        RECT 78.730 14.250 79.330 14.700 ;
        RECT 70.130 14.100 74.080 14.250 ;
        RECT 75.380 14.100 79.330 14.250 ;
        RECT 70.130 13.650 70.730 14.100 ;
        RECT 78.730 13.650 79.330 14.100 ;
        RECT 70.130 13.500 74.080 13.650 ;
        RECT 75.380 13.500 79.330 13.650 ;
        RECT 70.130 13.050 70.730 13.500 ;
        RECT 78.730 13.050 79.330 13.500 ;
        RECT 70.130 12.900 74.080 13.050 ;
        RECT 75.380 12.900 79.330 13.050 ;
        RECT 70.130 12.450 70.730 12.900 ;
        RECT 78.730 12.450 79.330 12.900 ;
        RECT 70.130 12.300 74.080 12.450 ;
        RECT 75.380 12.300 79.330 12.450 ;
        RECT 70.130 11.850 70.730 12.300 ;
        RECT 78.730 11.850 79.330 12.300 ;
        RECT 70.130 11.700 74.080 11.850 ;
        RECT 75.380 11.700 79.330 11.850 ;
        RECT 70.130 11.250 70.730 11.700 ;
        RECT 78.730 11.250 79.330 11.700 ;
        RECT 70.130 11.100 74.080 11.250 ;
        RECT 75.380 11.100 79.330 11.250 ;
        RECT 70.130 10.650 70.730 11.100 ;
        RECT 78.730 10.650 79.330 11.100 ;
        RECT 70.130 10.450 74.080 10.650 ;
        RECT 75.380 10.450 79.330 10.650 ;
        RECT 79.780 10.450 79.930 18.000 ;
        RECT 80.380 10.450 80.530 18.000 ;
        RECT 80.980 10.450 81.130 18.000 ;
        RECT 81.580 10.450 81.730 18.000 ;
        RECT 82.180 10.450 82.330 18.000 ;
        RECT 82.780 15.150 82.930 18.000 ;
        RECT 83.530 15.600 85.930 18.800 ;
        RECT 89.280 18.650 90.730 18.950 ;
        RECT 86.530 18.450 90.730 18.650 ;
        RECT 98.730 18.900 104.730 19.800 ;
        RECT 98.730 18.650 100.180 18.900 ;
        RECT 100.330 18.800 104.730 18.900 ;
        RECT 98.730 18.450 102.930 18.650 ;
        RECT 86.530 18.300 94.080 18.450 ;
        RECT 95.430 18.300 102.930 18.450 ;
        RECT 86.530 18.000 90.730 18.300 ;
        RECT 86.530 15.150 86.680 18.000 ;
        RECT 87.130 10.450 87.280 18.000 ;
        RECT 87.730 10.450 87.880 18.000 ;
        RECT 88.330 10.450 88.480 18.000 ;
        RECT 88.930 10.450 89.080 18.000 ;
        RECT 89.530 10.450 89.680 18.000 ;
        RECT 90.130 17.850 90.730 18.000 ;
        RECT 98.730 18.000 102.930 18.300 ;
        RECT 98.730 17.850 99.330 18.000 ;
        RECT 90.130 17.700 94.080 17.850 ;
        RECT 95.380 17.700 99.330 17.850 ;
        RECT 90.130 17.250 90.730 17.700 ;
        RECT 98.730 17.250 99.330 17.700 ;
        RECT 90.130 17.100 94.080 17.250 ;
        RECT 95.380 17.100 99.330 17.250 ;
        RECT 90.130 16.650 90.730 17.100 ;
        RECT 98.730 16.650 99.330 17.100 ;
        RECT 90.130 16.500 94.080 16.650 ;
        RECT 95.380 16.500 99.330 16.650 ;
        RECT 90.130 16.050 90.730 16.500 ;
        RECT 98.730 16.050 99.330 16.500 ;
        RECT 90.130 15.900 94.080 16.050 ;
        RECT 95.380 15.900 99.330 16.050 ;
        RECT 90.130 15.450 90.730 15.900 ;
        RECT 98.730 15.450 99.330 15.900 ;
        RECT 90.130 15.300 94.080 15.450 ;
        RECT 95.380 15.300 99.330 15.450 ;
        RECT 90.130 14.850 90.730 15.300 ;
        RECT 98.730 14.850 99.330 15.300 ;
        RECT 90.130 14.700 94.080 14.850 ;
        RECT 95.380 14.700 99.330 14.850 ;
        RECT 90.130 14.250 90.730 14.700 ;
        RECT 98.730 14.250 99.330 14.700 ;
        RECT 90.130 14.100 94.080 14.250 ;
        RECT 95.380 14.100 99.330 14.250 ;
        RECT 90.130 13.650 90.730 14.100 ;
        RECT 98.730 13.650 99.330 14.100 ;
        RECT 90.130 13.500 94.080 13.650 ;
        RECT 95.380 13.500 99.330 13.650 ;
        RECT 90.130 13.050 90.730 13.500 ;
        RECT 98.730 13.050 99.330 13.500 ;
        RECT 90.130 12.900 94.080 13.050 ;
        RECT 95.380 12.900 99.330 13.050 ;
        RECT 90.130 12.450 90.730 12.900 ;
        RECT 98.730 12.450 99.330 12.900 ;
        RECT 90.130 12.300 94.080 12.450 ;
        RECT 95.380 12.300 99.330 12.450 ;
        RECT 90.130 11.850 90.730 12.300 ;
        RECT 98.730 11.850 99.330 12.300 ;
        RECT 90.130 11.700 94.080 11.850 ;
        RECT 95.380 11.700 99.330 11.850 ;
        RECT 90.130 11.250 90.730 11.700 ;
        RECT 98.730 11.250 99.330 11.700 ;
        RECT 90.130 11.100 94.080 11.250 ;
        RECT 95.380 11.100 99.330 11.250 ;
        RECT 90.130 10.650 90.730 11.100 ;
        RECT 98.730 10.650 99.330 11.100 ;
        RECT 90.130 10.450 94.080 10.650 ;
        RECT 95.380 10.450 99.330 10.650 ;
        RECT 99.780 10.450 99.930 18.000 ;
        RECT 100.380 10.450 100.530 18.000 ;
        RECT 100.980 10.450 101.130 18.000 ;
        RECT 101.580 10.450 101.730 18.000 ;
        RECT 102.180 10.450 102.330 18.000 ;
        RECT 102.780 15.150 102.930 18.000 ;
        RECT 103.530 17.310 104.730 18.800 ;
        RECT 103.530 16.035 107.135 17.310 ;
        RECT 103.530 15.600 104.730 16.035 ;
        RECT 2.315 4.450 4.315 6.745 ;
        RECT 4.730 3.650 5.930 4.400 ;
        RECT 2.315 2.375 5.930 3.650 ;
        RECT 4.730 1.200 5.930 2.375 ;
        RECT 6.530 2.000 6.680 4.900 ;
        RECT 7.130 2.000 7.280 9.550 ;
        RECT 7.730 2.000 7.880 9.550 ;
        RECT 8.330 2.000 8.480 9.550 ;
        RECT 8.930 2.000 9.080 9.550 ;
        RECT 9.530 2.000 9.680 9.550 ;
        RECT 10.130 9.350 14.080 9.550 ;
        RECT 15.380 9.350 19.330 9.550 ;
        RECT 10.130 8.900 10.730 9.350 ;
        RECT 18.730 8.900 19.330 9.350 ;
        RECT 10.130 8.750 14.080 8.900 ;
        RECT 15.380 8.750 19.330 8.900 ;
        RECT 10.130 8.300 10.730 8.750 ;
        RECT 18.730 8.300 19.330 8.750 ;
        RECT 10.130 8.150 14.080 8.300 ;
        RECT 15.380 8.150 19.330 8.300 ;
        RECT 10.130 7.700 10.730 8.150 ;
        RECT 18.730 7.700 19.330 8.150 ;
        RECT 10.130 7.550 14.080 7.700 ;
        RECT 15.380 7.550 19.330 7.700 ;
        RECT 10.130 7.100 10.730 7.550 ;
        RECT 18.730 7.100 19.330 7.550 ;
        RECT 10.130 6.950 14.080 7.100 ;
        RECT 15.380 6.950 19.330 7.100 ;
        RECT 10.130 6.500 10.730 6.950 ;
        RECT 18.730 6.500 19.330 6.950 ;
        RECT 10.130 6.350 14.080 6.500 ;
        RECT 15.380 6.350 19.330 6.500 ;
        RECT 10.130 5.900 10.730 6.350 ;
        RECT 18.730 5.900 19.330 6.350 ;
        RECT 10.130 5.750 14.080 5.900 ;
        RECT 15.380 5.750 19.330 5.900 ;
        RECT 10.130 5.300 10.730 5.750 ;
        RECT 18.730 5.300 19.330 5.750 ;
        RECT 10.130 5.150 14.080 5.300 ;
        RECT 15.380 5.150 19.330 5.300 ;
        RECT 10.130 4.700 10.730 5.150 ;
        RECT 18.730 4.700 19.330 5.150 ;
        RECT 10.130 4.550 14.080 4.700 ;
        RECT 15.380 4.550 19.330 4.700 ;
        RECT 10.130 4.100 10.730 4.550 ;
        RECT 18.730 4.100 19.330 4.550 ;
        RECT 10.130 3.950 14.080 4.100 ;
        RECT 15.380 3.950 19.330 4.100 ;
        RECT 10.130 3.500 10.730 3.950 ;
        RECT 18.730 3.500 19.330 3.950 ;
        RECT 10.130 3.350 14.080 3.500 ;
        RECT 15.380 3.350 19.330 3.500 ;
        RECT 10.130 2.900 10.730 3.350 ;
        RECT 18.730 2.900 19.330 3.350 ;
        RECT 10.130 2.750 14.080 2.900 ;
        RECT 15.380 2.750 19.330 2.900 ;
        RECT 10.130 2.300 10.730 2.750 ;
        RECT 18.730 2.300 19.330 2.750 ;
        RECT 10.130 2.150 14.080 2.300 ;
        RECT 15.380 2.150 19.330 2.300 ;
        RECT 10.130 2.000 10.730 2.150 ;
        RECT 6.530 1.700 10.730 2.000 ;
        RECT 18.730 2.000 19.330 2.150 ;
        RECT 19.780 2.000 19.930 9.550 ;
        RECT 20.380 2.000 20.530 9.550 ;
        RECT 20.980 2.000 21.130 9.550 ;
        RECT 21.580 2.000 21.730 9.550 ;
        RECT 22.180 2.000 22.330 9.550 ;
        RECT 22.780 2.000 22.930 4.900 ;
        RECT 18.730 1.700 22.930 2.000 ;
        RECT 6.530 1.550 14.080 1.700 ;
        RECT 15.380 1.550 22.930 1.700 ;
        RECT 6.530 1.350 10.730 1.550 ;
        RECT 4.730 1.050 9.130 1.200 ;
        RECT 9.280 1.050 10.730 1.350 ;
        RECT 4.730 0.150 10.730 1.050 ;
        RECT 18.730 1.350 22.930 1.550 ;
        RECT 18.730 1.050 20.180 1.350 ;
        RECT 23.530 1.200 25.930 4.400 ;
        RECT 26.530 2.000 26.680 4.900 ;
        RECT 27.130 2.000 27.280 9.550 ;
        RECT 27.730 2.000 27.880 9.550 ;
        RECT 28.330 2.000 28.480 9.550 ;
        RECT 28.930 2.000 29.080 9.550 ;
        RECT 29.530 2.000 29.680 9.550 ;
        RECT 30.130 9.350 34.080 9.550 ;
        RECT 35.380 9.350 39.330 9.550 ;
        RECT 30.130 8.900 30.730 9.350 ;
        RECT 38.730 8.900 39.330 9.350 ;
        RECT 30.130 8.750 34.080 8.900 ;
        RECT 35.380 8.750 39.330 8.900 ;
        RECT 30.130 8.300 30.730 8.750 ;
        RECT 38.730 8.300 39.330 8.750 ;
        RECT 30.130 8.150 34.080 8.300 ;
        RECT 35.380 8.150 39.330 8.300 ;
        RECT 30.130 7.700 30.730 8.150 ;
        RECT 38.730 7.700 39.330 8.150 ;
        RECT 30.130 7.550 34.080 7.700 ;
        RECT 35.380 7.550 39.330 7.700 ;
        RECT 30.130 7.100 30.730 7.550 ;
        RECT 38.730 7.100 39.330 7.550 ;
        RECT 30.130 6.950 34.080 7.100 ;
        RECT 35.380 6.950 39.330 7.100 ;
        RECT 30.130 6.500 30.730 6.950 ;
        RECT 38.730 6.500 39.330 6.950 ;
        RECT 30.130 6.350 34.080 6.500 ;
        RECT 35.380 6.350 39.330 6.500 ;
        RECT 30.130 5.900 30.730 6.350 ;
        RECT 38.730 5.900 39.330 6.350 ;
        RECT 30.130 5.750 34.080 5.900 ;
        RECT 35.380 5.750 39.330 5.900 ;
        RECT 30.130 5.300 30.730 5.750 ;
        RECT 38.730 5.300 39.330 5.750 ;
        RECT 30.130 5.150 34.080 5.300 ;
        RECT 35.380 5.150 39.330 5.300 ;
        RECT 30.130 4.700 30.730 5.150 ;
        RECT 38.730 4.700 39.330 5.150 ;
        RECT 30.130 4.550 34.080 4.700 ;
        RECT 35.380 4.550 39.330 4.700 ;
        RECT 30.130 4.100 30.730 4.550 ;
        RECT 38.730 4.100 39.330 4.550 ;
        RECT 30.130 3.950 34.080 4.100 ;
        RECT 35.380 3.950 39.330 4.100 ;
        RECT 30.130 3.500 30.730 3.950 ;
        RECT 38.730 3.500 39.330 3.950 ;
        RECT 30.130 3.350 34.080 3.500 ;
        RECT 35.380 3.350 39.330 3.500 ;
        RECT 30.130 2.900 30.730 3.350 ;
        RECT 38.730 2.900 39.330 3.350 ;
        RECT 30.130 2.750 34.080 2.900 ;
        RECT 35.380 2.750 39.330 2.900 ;
        RECT 30.130 2.300 30.730 2.750 ;
        RECT 38.730 2.300 39.330 2.750 ;
        RECT 30.130 2.150 34.080 2.300 ;
        RECT 35.380 2.150 39.330 2.300 ;
        RECT 30.130 2.000 30.730 2.150 ;
        RECT 26.530 1.700 30.730 2.000 ;
        RECT 38.730 2.000 39.330 2.150 ;
        RECT 39.780 2.000 39.930 9.550 ;
        RECT 40.380 2.000 40.530 9.550 ;
        RECT 40.980 2.000 41.130 9.550 ;
        RECT 41.580 2.000 41.730 9.550 ;
        RECT 42.180 2.000 42.330 9.550 ;
        RECT 42.780 2.000 42.930 4.900 ;
        RECT 38.730 1.700 42.930 2.000 ;
        RECT 26.530 1.550 34.080 1.700 ;
        RECT 35.380 1.550 42.930 1.700 ;
        RECT 26.530 1.350 30.730 1.550 ;
        RECT 20.330 1.050 29.130 1.200 ;
        RECT 29.280 1.050 30.730 1.350 ;
        RECT 18.730 0.150 30.730 1.050 ;
        RECT 38.730 1.350 42.930 1.550 ;
        RECT 38.730 1.050 40.180 1.350 ;
        RECT 43.530 1.200 45.930 4.400 ;
        RECT 46.530 2.000 46.680 4.900 ;
        RECT 47.130 2.000 47.280 9.550 ;
        RECT 47.730 2.000 47.880 9.550 ;
        RECT 48.330 2.000 48.480 9.550 ;
        RECT 48.930 2.000 49.080 9.550 ;
        RECT 49.530 2.000 49.680 9.550 ;
        RECT 50.130 9.350 54.080 9.550 ;
        RECT 55.380 9.350 59.330 9.550 ;
        RECT 50.130 8.900 50.730 9.350 ;
        RECT 58.730 8.900 59.330 9.350 ;
        RECT 50.130 8.750 54.080 8.900 ;
        RECT 55.380 8.750 59.330 8.900 ;
        RECT 50.130 8.300 50.730 8.750 ;
        RECT 58.730 8.300 59.330 8.750 ;
        RECT 50.130 8.150 54.080 8.300 ;
        RECT 55.380 8.150 59.330 8.300 ;
        RECT 50.130 7.700 50.730 8.150 ;
        RECT 58.730 7.700 59.330 8.150 ;
        RECT 50.130 7.550 54.080 7.700 ;
        RECT 55.380 7.550 59.330 7.700 ;
        RECT 50.130 7.100 50.730 7.550 ;
        RECT 58.730 7.100 59.330 7.550 ;
        RECT 50.130 6.950 54.080 7.100 ;
        RECT 55.380 6.950 59.330 7.100 ;
        RECT 50.130 6.500 50.730 6.950 ;
        RECT 58.730 6.500 59.330 6.950 ;
        RECT 50.130 6.350 54.080 6.500 ;
        RECT 55.380 6.350 59.330 6.500 ;
        RECT 50.130 5.900 50.730 6.350 ;
        RECT 58.730 5.900 59.330 6.350 ;
        RECT 50.130 5.750 54.080 5.900 ;
        RECT 55.380 5.750 59.330 5.900 ;
        RECT 50.130 5.300 50.730 5.750 ;
        RECT 58.730 5.300 59.330 5.750 ;
        RECT 50.130 5.150 54.080 5.300 ;
        RECT 55.380 5.150 59.330 5.300 ;
        RECT 50.130 4.700 50.730 5.150 ;
        RECT 58.730 4.700 59.330 5.150 ;
        RECT 50.130 4.550 54.080 4.700 ;
        RECT 55.380 4.550 59.330 4.700 ;
        RECT 50.130 4.100 50.730 4.550 ;
        RECT 58.730 4.100 59.330 4.550 ;
        RECT 50.130 3.950 54.080 4.100 ;
        RECT 55.380 3.950 59.330 4.100 ;
        RECT 50.130 3.500 50.730 3.950 ;
        RECT 58.730 3.500 59.330 3.950 ;
        RECT 50.130 3.350 54.080 3.500 ;
        RECT 55.380 3.350 59.330 3.500 ;
        RECT 50.130 2.900 50.730 3.350 ;
        RECT 58.730 2.900 59.330 3.350 ;
        RECT 50.130 2.750 54.080 2.900 ;
        RECT 55.380 2.750 59.330 2.900 ;
        RECT 50.130 2.300 50.730 2.750 ;
        RECT 58.730 2.300 59.330 2.750 ;
        RECT 50.130 2.150 54.080 2.300 ;
        RECT 55.380 2.150 59.330 2.300 ;
        RECT 50.130 2.000 50.730 2.150 ;
        RECT 46.530 1.700 50.730 2.000 ;
        RECT 58.730 2.000 59.330 2.150 ;
        RECT 59.780 2.000 59.930 9.550 ;
        RECT 60.380 2.000 60.530 9.550 ;
        RECT 60.980 2.000 61.130 9.550 ;
        RECT 61.580 2.000 61.730 9.550 ;
        RECT 62.180 2.000 62.330 9.550 ;
        RECT 62.780 2.000 62.930 4.900 ;
        RECT 58.730 1.700 62.930 2.000 ;
        RECT 46.530 1.550 54.080 1.700 ;
        RECT 55.380 1.550 62.930 1.700 ;
        RECT 46.530 1.350 50.730 1.550 ;
        RECT 40.330 1.050 49.130 1.200 ;
        RECT 49.280 1.050 50.730 1.350 ;
        RECT 38.730 0.150 50.730 1.050 ;
        RECT 58.730 1.350 62.930 1.550 ;
        RECT 58.730 1.050 60.180 1.350 ;
        RECT 63.530 1.200 65.930 4.400 ;
        RECT 66.530 2.000 66.680 4.900 ;
        RECT 67.130 2.000 67.280 9.550 ;
        RECT 67.730 2.000 67.880 9.550 ;
        RECT 68.330 2.000 68.480 9.550 ;
        RECT 68.930 2.000 69.080 9.550 ;
        RECT 69.530 2.000 69.680 9.550 ;
        RECT 70.130 9.350 74.080 9.550 ;
        RECT 75.380 9.350 79.330 9.550 ;
        RECT 70.130 8.900 70.730 9.350 ;
        RECT 78.730 8.900 79.330 9.350 ;
        RECT 70.130 8.750 74.080 8.900 ;
        RECT 75.380 8.750 79.330 8.900 ;
        RECT 70.130 8.300 70.730 8.750 ;
        RECT 78.730 8.300 79.330 8.750 ;
        RECT 70.130 8.150 74.080 8.300 ;
        RECT 75.380 8.150 79.330 8.300 ;
        RECT 70.130 7.700 70.730 8.150 ;
        RECT 78.730 7.700 79.330 8.150 ;
        RECT 70.130 7.550 74.080 7.700 ;
        RECT 75.380 7.550 79.330 7.700 ;
        RECT 70.130 7.100 70.730 7.550 ;
        RECT 78.730 7.100 79.330 7.550 ;
        RECT 70.130 6.950 74.080 7.100 ;
        RECT 75.380 6.950 79.330 7.100 ;
        RECT 70.130 6.500 70.730 6.950 ;
        RECT 78.730 6.500 79.330 6.950 ;
        RECT 70.130 6.350 74.080 6.500 ;
        RECT 75.380 6.350 79.330 6.500 ;
        RECT 70.130 5.900 70.730 6.350 ;
        RECT 78.730 5.900 79.330 6.350 ;
        RECT 70.130 5.750 74.080 5.900 ;
        RECT 75.380 5.750 79.330 5.900 ;
        RECT 70.130 5.300 70.730 5.750 ;
        RECT 78.730 5.300 79.330 5.750 ;
        RECT 70.130 5.150 74.080 5.300 ;
        RECT 75.380 5.150 79.330 5.300 ;
        RECT 70.130 4.700 70.730 5.150 ;
        RECT 78.730 4.700 79.330 5.150 ;
        RECT 70.130 4.550 74.080 4.700 ;
        RECT 75.380 4.550 79.330 4.700 ;
        RECT 70.130 4.100 70.730 4.550 ;
        RECT 78.730 4.100 79.330 4.550 ;
        RECT 70.130 3.950 74.080 4.100 ;
        RECT 75.380 3.950 79.330 4.100 ;
        RECT 70.130 3.500 70.730 3.950 ;
        RECT 78.730 3.500 79.330 3.950 ;
        RECT 70.130 3.350 74.080 3.500 ;
        RECT 75.380 3.350 79.330 3.500 ;
        RECT 70.130 2.900 70.730 3.350 ;
        RECT 78.730 2.900 79.330 3.350 ;
        RECT 70.130 2.750 74.080 2.900 ;
        RECT 75.380 2.750 79.330 2.900 ;
        RECT 70.130 2.300 70.730 2.750 ;
        RECT 78.730 2.300 79.330 2.750 ;
        RECT 70.130 2.150 74.080 2.300 ;
        RECT 75.380 2.150 79.330 2.300 ;
        RECT 70.130 2.000 70.730 2.150 ;
        RECT 66.530 1.700 70.730 2.000 ;
        RECT 78.730 2.000 79.330 2.150 ;
        RECT 79.780 2.000 79.930 9.550 ;
        RECT 80.380 2.000 80.530 9.550 ;
        RECT 80.980 2.000 81.130 9.550 ;
        RECT 81.580 2.000 81.730 9.550 ;
        RECT 82.180 2.000 82.330 9.550 ;
        RECT 82.780 2.000 82.930 4.900 ;
        RECT 78.730 1.700 82.930 2.000 ;
        RECT 66.530 1.550 74.080 1.700 ;
        RECT 75.380 1.550 82.930 1.700 ;
        RECT 66.530 1.350 70.730 1.550 ;
        RECT 60.330 1.050 69.130 1.200 ;
        RECT 69.280 1.050 70.730 1.350 ;
        RECT 58.730 0.150 70.730 1.050 ;
        RECT 78.730 1.350 82.930 1.550 ;
        RECT 78.730 1.050 80.180 1.350 ;
        RECT 83.530 1.200 85.930 4.400 ;
        RECT 86.530 2.000 86.680 4.900 ;
        RECT 87.130 2.000 87.280 9.550 ;
        RECT 87.730 2.000 87.880 9.550 ;
        RECT 88.330 2.000 88.480 9.550 ;
        RECT 88.930 2.000 89.080 9.550 ;
        RECT 89.530 2.000 89.680 9.550 ;
        RECT 90.130 9.350 94.080 9.550 ;
        RECT 95.380 9.350 99.330 9.550 ;
        RECT 90.130 8.900 90.730 9.350 ;
        RECT 98.730 8.900 99.330 9.350 ;
        RECT 90.130 8.750 94.080 8.900 ;
        RECT 95.380 8.750 99.330 8.900 ;
        RECT 90.130 8.300 90.730 8.750 ;
        RECT 98.730 8.300 99.330 8.750 ;
        RECT 90.130 8.150 94.080 8.300 ;
        RECT 95.380 8.150 99.330 8.300 ;
        RECT 90.130 7.700 90.730 8.150 ;
        RECT 98.730 7.700 99.330 8.150 ;
        RECT 90.130 7.550 94.080 7.700 ;
        RECT 95.380 7.550 99.330 7.700 ;
        RECT 90.130 7.100 90.730 7.550 ;
        RECT 98.730 7.100 99.330 7.550 ;
        RECT 90.130 6.950 94.080 7.100 ;
        RECT 95.380 6.950 99.330 7.100 ;
        RECT 90.130 6.500 90.730 6.950 ;
        RECT 98.730 6.500 99.330 6.950 ;
        RECT 90.130 6.350 94.080 6.500 ;
        RECT 95.380 6.350 99.330 6.500 ;
        RECT 90.130 5.900 90.730 6.350 ;
        RECT 98.730 5.900 99.330 6.350 ;
        RECT 90.130 5.750 94.080 5.900 ;
        RECT 95.380 5.750 99.330 5.900 ;
        RECT 90.130 5.300 90.730 5.750 ;
        RECT 98.730 5.300 99.330 5.750 ;
        RECT 90.130 5.150 94.080 5.300 ;
        RECT 95.380 5.150 99.330 5.300 ;
        RECT 90.130 4.700 90.730 5.150 ;
        RECT 98.730 4.700 99.330 5.150 ;
        RECT 90.130 4.550 94.080 4.700 ;
        RECT 95.380 4.550 99.330 4.700 ;
        RECT 90.130 4.100 90.730 4.550 ;
        RECT 98.730 4.100 99.330 4.550 ;
        RECT 90.130 3.950 94.080 4.100 ;
        RECT 95.380 3.950 99.330 4.100 ;
        RECT 90.130 3.500 90.730 3.950 ;
        RECT 98.730 3.500 99.330 3.950 ;
        RECT 90.130 3.350 94.080 3.500 ;
        RECT 95.380 3.350 99.330 3.500 ;
        RECT 90.130 2.900 90.730 3.350 ;
        RECT 98.730 2.900 99.330 3.350 ;
        RECT 90.130 2.750 94.080 2.900 ;
        RECT 95.380 2.750 99.330 2.900 ;
        RECT 90.130 2.300 90.730 2.750 ;
        RECT 98.730 2.300 99.330 2.750 ;
        RECT 90.130 2.150 94.080 2.300 ;
        RECT 95.380 2.150 99.330 2.300 ;
        RECT 90.130 2.000 90.730 2.150 ;
        RECT 86.530 1.700 90.730 2.000 ;
        RECT 98.730 2.000 99.330 2.150 ;
        RECT 99.780 2.000 99.930 9.550 ;
        RECT 100.380 2.000 100.530 9.550 ;
        RECT 100.980 2.000 101.130 9.550 ;
        RECT 101.580 2.000 101.730 9.550 ;
        RECT 102.180 2.000 102.330 9.550 ;
        RECT 102.780 2.000 102.930 4.900 ;
        RECT 98.730 1.700 102.930 2.000 ;
        RECT 86.530 1.550 94.080 1.700 ;
        RECT 95.380 1.550 102.930 1.700 ;
        RECT 86.530 1.350 90.730 1.550 ;
        RECT 80.330 1.050 89.130 1.200 ;
        RECT 89.280 1.050 90.730 1.350 ;
        RECT 78.730 0.150 90.730 1.050 ;
        RECT 98.730 1.350 102.930 1.550 ;
        RECT 103.530 3.095 104.730 4.400 ;
        RECT 103.530 1.820 107.140 3.095 ;
        RECT 98.730 1.050 100.180 1.350 ;
        RECT 103.530 1.200 104.730 1.820 ;
        RECT 100.330 1.050 104.730 1.200 ;
        RECT 98.730 0.150 104.730 1.050 ;
        RECT 4.730 0.000 9.130 0.150 ;
        RECT 20.330 0.000 29.130 0.150 ;
        RECT 40.330 0.000 49.130 0.150 ;
        RECT 60.330 0.000 69.130 0.150 ;
        RECT 80.330 0.000 89.130 0.150 ;
        RECT 100.330 0.000 104.730 0.150 ;
      LAYER via ;
        RECT 4.830 378.900 5.830 379.900 ;
        RECT 6.430 378.900 7.430 379.900 ;
        RECT 8.030 378.900 9.030 379.900 ;
        RECT 4.830 377.300 5.830 378.300 ;
        RECT 2.515 376.880 2.875 377.260 ;
        RECT 3.145 376.880 3.505 377.260 ;
        RECT 3.745 376.880 4.105 377.260 ;
        RECT 2.515 376.290 2.875 376.670 ;
        RECT 3.145 376.290 3.505 376.670 ;
        RECT 3.745 376.290 4.105 376.670 ;
        RECT 4.830 375.700 5.830 376.700 ;
        RECT 20.430 378.900 21.430 379.900 ;
        RECT 22.030 378.900 23.030 379.900 ;
        RECT 23.630 378.900 24.630 379.900 ;
        RECT 24.830 378.900 25.830 379.900 ;
        RECT 26.430 378.900 27.430 379.900 ;
        RECT 28.030 378.900 29.030 379.900 ;
        RECT 2.520 374.920 2.880 375.300 ;
        RECT 3.130 374.920 3.490 375.300 ;
        RECT 3.760 374.920 4.120 375.300 ;
        RECT 2.520 374.185 2.880 374.565 ;
        RECT 3.130 374.185 3.490 374.565 ;
        RECT 3.760 374.185 4.120 374.565 ;
        RECT 2.520 373.500 2.880 373.880 ;
        RECT 3.130 373.500 3.490 373.880 ;
        RECT 3.760 373.500 4.120 373.880 ;
        RECT 23.630 377.300 24.630 378.300 ;
        RECT 24.830 377.300 25.830 378.300 ;
        RECT 23.630 375.700 24.630 376.700 ;
        RECT 24.830 375.700 25.830 376.700 ;
        RECT 40.430 378.900 41.430 379.900 ;
        RECT 42.030 378.900 43.030 379.900 ;
        RECT 43.630 378.900 44.630 379.900 ;
        RECT 44.830 378.900 45.830 379.900 ;
        RECT 46.430 378.900 47.430 379.900 ;
        RECT 48.030 378.900 49.030 379.900 ;
        RECT 43.630 377.300 44.630 378.300 ;
        RECT 44.830 377.300 45.830 378.300 ;
        RECT 43.630 375.700 44.630 376.700 ;
        RECT 44.830 375.700 45.830 376.700 ;
        RECT 60.430 378.900 61.430 379.900 ;
        RECT 62.030 378.900 63.030 379.900 ;
        RECT 63.630 378.900 64.630 379.900 ;
        RECT 64.830 378.900 65.830 379.900 ;
        RECT 66.430 378.900 67.430 379.900 ;
        RECT 68.030 378.900 69.030 379.900 ;
        RECT 63.630 377.300 64.630 378.300 ;
        RECT 64.830 377.300 65.830 378.300 ;
        RECT 63.630 375.700 64.630 376.700 ;
        RECT 64.830 375.700 65.830 376.700 ;
        RECT 80.430 378.900 81.430 379.900 ;
        RECT 82.030 378.900 83.030 379.900 ;
        RECT 83.630 378.900 84.630 379.900 ;
        RECT 84.830 378.900 85.830 379.900 ;
        RECT 86.430 378.900 87.430 379.900 ;
        RECT 88.030 378.900 89.030 379.900 ;
        RECT 83.630 377.300 84.630 378.300 ;
        RECT 84.830 377.300 85.830 378.300 ;
        RECT 83.630 375.700 84.630 376.700 ;
        RECT 84.830 375.700 85.830 376.700 ;
        RECT 100.430 378.900 101.430 379.900 ;
        RECT 102.030 378.900 103.030 379.900 ;
        RECT 103.630 378.900 104.630 379.900 ;
        RECT 103.630 377.300 104.630 378.300 ;
        RECT 105.340 377.080 105.700 377.460 ;
        RECT 105.970 377.080 106.330 377.460 ;
        RECT 106.570 377.080 106.930 377.460 ;
        RECT 103.630 375.700 104.630 376.700 ;
        RECT 105.340 376.490 105.700 376.870 ;
        RECT 105.970 376.490 106.330 376.870 ;
        RECT 106.570 376.490 106.930 376.870 ;
        RECT 2.520 366.120 2.880 366.500 ;
        RECT 3.130 366.120 3.490 366.500 ;
        RECT 3.760 366.120 4.120 366.500 ;
        RECT 2.520 365.385 2.880 365.765 ;
        RECT 3.130 365.385 3.490 365.765 ;
        RECT 3.760 365.385 4.120 365.765 ;
        RECT 2.520 364.700 2.880 365.080 ;
        RECT 3.130 364.700 3.490 365.080 ;
        RECT 3.760 364.700 4.120 365.080 ;
        RECT 2.515 363.515 2.875 363.895 ;
        RECT 3.145 363.515 3.505 363.895 ;
        RECT 3.745 363.515 4.105 363.895 ;
        RECT 2.515 362.925 2.875 363.305 ;
        RECT 3.145 362.925 3.505 363.305 ;
        RECT 3.745 362.925 4.105 363.305 ;
        RECT 4.830 363.300 5.830 364.300 ;
        RECT 4.830 361.700 5.830 362.700 ;
        RECT 4.830 360.100 5.830 361.100 ;
        RECT 6.430 360.100 7.430 361.100 ;
        RECT 8.030 360.100 9.030 361.100 ;
        RECT 23.630 363.300 24.630 364.300 ;
        RECT 24.830 363.300 25.830 364.300 ;
        RECT 23.630 361.700 24.630 362.700 ;
        RECT 24.830 361.700 25.830 362.700 ;
        RECT 4.830 358.900 5.830 359.900 ;
        RECT 6.430 358.900 7.430 359.900 ;
        RECT 8.030 358.900 9.030 359.900 ;
        RECT 20.430 360.100 21.430 361.100 ;
        RECT 22.030 360.100 23.030 361.100 ;
        RECT 23.630 360.100 24.630 361.100 ;
        RECT 24.830 360.100 25.830 361.100 ;
        RECT 26.430 360.100 27.430 361.100 ;
        RECT 28.030 360.100 29.030 361.100 ;
        RECT 43.630 363.300 44.630 364.300 ;
        RECT 44.830 363.300 45.830 364.300 ;
        RECT 43.630 361.700 44.630 362.700 ;
        RECT 44.830 361.700 45.830 362.700 ;
        RECT 4.830 357.300 5.830 358.300 ;
        RECT 2.515 356.880 2.875 357.260 ;
        RECT 3.145 356.880 3.505 357.260 ;
        RECT 3.745 356.880 4.105 357.260 ;
        RECT 2.515 356.290 2.875 356.670 ;
        RECT 3.145 356.290 3.505 356.670 ;
        RECT 3.745 356.290 4.105 356.670 ;
        RECT 4.830 355.700 5.830 356.700 ;
        RECT 20.430 358.900 21.430 359.900 ;
        RECT 22.030 358.900 23.030 359.900 ;
        RECT 23.630 358.900 24.630 359.900 ;
        RECT 24.830 358.900 25.830 359.900 ;
        RECT 26.430 358.900 27.430 359.900 ;
        RECT 28.030 358.900 29.030 359.900 ;
        RECT 40.430 360.100 41.430 361.100 ;
        RECT 42.030 360.100 43.030 361.100 ;
        RECT 43.630 360.100 44.630 361.100 ;
        RECT 44.830 360.100 45.830 361.100 ;
        RECT 46.430 360.100 47.430 361.100 ;
        RECT 48.030 360.100 49.030 361.100 ;
        RECT 63.630 363.300 64.630 364.300 ;
        RECT 64.830 363.300 65.830 364.300 ;
        RECT 63.630 361.700 64.630 362.700 ;
        RECT 64.830 361.700 65.830 362.700 ;
        RECT 2.520 354.920 2.880 355.300 ;
        RECT 3.130 354.920 3.490 355.300 ;
        RECT 3.760 354.920 4.120 355.300 ;
        RECT 2.520 354.185 2.880 354.565 ;
        RECT 3.130 354.185 3.490 354.565 ;
        RECT 3.760 354.185 4.120 354.565 ;
        RECT 2.520 353.500 2.880 353.880 ;
        RECT 3.130 353.500 3.490 353.880 ;
        RECT 3.760 353.500 4.120 353.880 ;
        RECT 23.630 357.300 24.630 358.300 ;
        RECT 24.830 357.300 25.830 358.300 ;
        RECT 23.630 355.700 24.630 356.700 ;
        RECT 24.830 355.700 25.830 356.700 ;
        RECT 40.430 358.900 41.430 359.900 ;
        RECT 42.030 358.900 43.030 359.900 ;
        RECT 43.630 358.900 44.630 359.900 ;
        RECT 44.830 358.900 45.830 359.900 ;
        RECT 46.430 358.900 47.430 359.900 ;
        RECT 48.030 358.900 49.030 359.900 ;
        RECT 60.430 360.100 61.430 361.100 ;
        RECT 62.030 360.100 63.030 361.100 ;
        RECT 63.630 360.100 64.630 361.100 ;
        RECT 64.830 360.100 65.830 361.100 ;
        RECT 66.430 360.100 67.430 361.100 ;
        RECT 68.030 360.100 69.030 361.100 ;
        RECT 83.630 363.300 84.630 364.300 ;
        RECT 84.830 363.300 85.830 364.300 ;
        RECT 83.630 361.700 84.630 362.700 ;
        RECT 84.830 361.700 85.830 362.700 ;
        RECT 43.630 357.300 44.630 358.300 ;
        RECT 44.830 357.300 45.830 358.300 ;
        RECT 43.630 355.700 44.630 356.700 ;
        RECT 44.830 355.700 45.830 356.700 ;
        RECT 60.430 358.900 61.430 359.900 ;
        RECT 62.030 358.900 63.030 359.900 ;
        RECT 63.630 358.900 64.630 359.900 ;
        RECT 64.830 358.900 65.830 359.900 ;
        RECT 66.430 358.900 67.430 359.900 ;
        RECT 68.030 358.900 69.030 359.900 ;
        RECT 80.430 360.100 81.430 361.100 ;
        RECT 82.030 360.100 83.030 361.100 ;
        RECT 83.630 360.100 84.630 361.100 ;
        RECT 84.830 360.100 85.830 361.100 ;
        RECT 86.430 360.100 87.430 361.100 ;
        RECT 88.030 360.100 89.030 361.100 ;
        RECT 103.630 363.300 104.630 364.300 ;
        RECT 105.340 363.095 105.700 363.475 ;
        RECT 105.970 363.095 106.330 363.475 ;
        RECT 106.570 363.095 106.930 363.475 ;
        RECT 103.630 361.700 104.630 362.700 ;
        RECT 105.340 362.505 105.700 362.885 ;
        RECT 105.970 362.505 106.330 362.885 ;
        RECT 106.570 362.505 106.930 362.885 ;
        RECT 63.630 357.300 64.630 358.300 ;
        RECT 64.830 357.300 65.830 358.300 ;
        RECT 63.630 355.700 64.630 356.700 ;
        RECT 64.830 355.700 65.830 356.700 ;
        RECT 80.430 358.900 81.430 359.900 ;
        RECT 82.030 358.900 83.030 359.900 ;
        RECT 83.630 358.900 84.630 359.900 ;
        RECT 84.830 358.900 85.830 359.900 ;
        RECT 86.430 358.900 87.430 359.900 ;
        RECT 88.030 358.900 89.030 359.900 ;
        RECT 100.430 360.100 101.430 361.100 ;
        RECT 102.030 360.100 103.030 361.100 ;
        RECT 103.630 360.100 104.630 361.100 ;
        RECT 83.630 357.300 84.630 358.300 ;
        RECT 84.830 357.300 85.830 358.300 ;
        RECT 83.630 355.700 84.630 356.700 ;
        RECT 84.830 355.700 85.830 356.700 ;
        RECT 100.430 358.900 101.430 359.900 ;
        RECT 102.030 358.900 103.030 359.900 ;
        RECT 103.630 358.900 104.630 359.900 ;
        RECT 103.630 357.300 104.630 358.300 ;
        RECT 105.340 357.080 105.700 357.460 ;
        RECT 105.970 357.080 106.330 357.460 ;
        RECT 106.570 357.080 106.930 357.460 ;
        RECT 103.630 355.700 104.630 356.700 ;
        RECT 105.340 356.490 105.700 356.870 ;
        RECT 105.970 356.490 106.330 356.870 ;
        RECT 106.570 356.490 106.930 356.870 ;
        RECT 2.520 346.120 2.880 346.500 ;
        RECT 3.130 346.120 3.490 346.500 ;
        RECT 3.760 346.120 4.120 346.500 ;
        RECT 2.520 345.385 2.880 345.765 ;
        RECT 3.130 345.385 3.490 345.765 ;
        RECT 3.760 345.385 4.120 345.765 ;
        RECT 2.520 344.700 2.880 345.080 ;
        RECT 3.130 344.700 3.490 345.080 ;
        RECT 3.760 344.700 4.120 345.080 ;
        RECT 2.515 343.515 2.875 343.895 ;
        RECT 3.145 343.515 3.505 343.895 ;
        RECT 3.745 343.515 4.105 343.895 ;
        RECT 2.515 342.925 2.875 343.305 ;
        RECT 3.145 342.925 3.505 343.305 ;
        RECT 3.745 342.925 4.105 343.305 ;
        RECT 4.830 343.300 5.830 344.300 ;
        RECT 4.830 341.700 5.830 342.700 ;
        RECT 4.830 340.100 5.830 341.100 ;
        RECT 6.430 340.100 7.430 341.100 ;
        RECT 8.030 340.100 9.030 341.100 ;
        RECT 23.630 343.300 24.630 344.300 ;
        RECT 24.830 343.300 25.830 344.300 ;
        RECT 23.630 341.700 24.630 342.700 ;
        RECT 24.830 341.700 25.830 342.700 ;
        RECT 4.830 338.900 5.830 339.900 ;
        RECT 6.430 338.900 7.430 339.900 ;
        RECT 8.030 338.900 9.030 339.900 ;
        RECT 20.430 340.100 21.430 341.100 ;
        RECT 22.030 340.100 23.030 341.100 ;
        RECT 23.630 340.100 24.630 341.100 ;
        RECT 24.830 340.100 25.830 341.100 ;
        RECT 26.430 340.100 27.430 341.100 ;
        RECT 28.030 340.100 29.030 341.100 ;
        RECT 43.630 343.300 44.630 344.300 ;
        RECT 44.830 343.300 45.830 344.300 ;
        RECT 43.630 341.700 44.630 342.700 ;
        RECT 44.830 341.700 45.830 342.700 ;
        RECT 4.830 337.300 5.830 338.300 ;
        RECT 2.515 336.870 2.875 337.250 ;
        RECT 3.145 336.870 3.505 337.250 ;
        RECT 3.745 336.870 4.105 337.250 ;
        RECT 2.515 336.280 2.875 336.660 ;
        RECT 3.145 336.280 3.505 336.660 ;
        RECT 3.745 336.280 4.105 336.660 ;
        RECT 4.830 335.700 5.830 336.700 ;
        RECT 20.430 338.900 21.430 339.900 ;
        RECT 22.030 338.900 23.030 339.900 ;
        RECT 23.630 338.900 24.630 339.900 ;
        RECT 24.830 338.900 25.830 339.900 ;
        RECT 26.430 338.900 27.430 339.900 ;
        RECT 28.030 338.900 29.030 339.900 ;
        RECT 40.430 340.100 41.430 341.100 ;
        RECT 42.030 340.100 43.030 341.100 ;
        RECT 43.630 340.100 44.630 341.100 ;
        RECT 44.830 340.100 45.830 341.100 ;
        RECT 46.430 340.100 47.430 341.100 ;
        RECT 48.030 340.100 49.030 341.100 ;
        RECT 63.630 343.300 64.630 344.300 ;
        RECT 64.830 343.300 65.830 344.300 ;
        RECT 63.630 341.700 64.630 342.700 ;
        RECT 64.830 341.700 65.830 342.700 ;
        RECT 2.520 334.920 2.880 335.300 ;
        RECT 3.130 334.920 3.490 335.300 ;
        RECT 3.760 334.920 4.120 335.300 ;
        RECT 2.520 334.185 2.880 334.565 ;
        RECT 3.130 334.185 3.490 334.565 ;
        RECT 3.760 334.185 4.120 334.565 ;
        RECT 2.520 333.500 2.880 333.880 ;
        RECT 3.130 333.500 3.490 333.880 ;
        RECT 3.760 333.500 4.120 333.880 ;
        RECT 23.630 337.300 24.630 338.300 ;
        RECT 24.830 337.300 25.830 338.300 ;
        RECT 23.630 335.700 24.630 336.700 ;
        RECT 24.830 335.700 25.830 336.700 ;
        RECT 40.430 338.900 41.430 339.900 ;
        RECT 42.030 338.900 43.030 339.900 ;
        RECT 43.630 338.900 44.630 339.900 ;
        RECT 44.830 338.900 45.830 339.900 ;
        RECT 46.430 338.900 47.430 339.900 ;
        RECT 48.030 338.900 49.030 339.900 ;
        RECT 60.430 340.100 61.430 341.100 ;
        RECT 62.030 340.100 63.030 341.100 ;
        RECT 63.630 340.100 64.630 341.100 ;
        RECT 64.830 340.100 65.830 341.100 ;
        RECT 66.430 340.100 67.430 341.100 ;
        RECT 68.030 340.100 69.030 341.100 ;
        RECT 83.630 343.300 84.630 344.300 ;
        RECT 84.830 343.300 85.830 344.300 ;
        RECT 83.630 341.700 84.630 342.700 ;
        RECT 84.830 341.700 85.830 342.700 ;
        RECT 43.630 337.300 44.630 338.300 ;
        RECT 44.830 337.300 45.830 338.300 ;
        RECT 43.630 335.700 44.630 336.700 ;
        RECT 44.830 335.700 45.830 336.700 ;
        RECT 60.430 338.900 61.430 339.900 ;
        RECT 62.030 338.900 63.030 339.900 ;
        RECT 63.630 338.900 64.630 339.900 ;
        RECT 64.830 338.900 65.830 339.900 ;
        RECT 66.430 338.900 67.430 339.900 ;
        RECT 68.030 338.900 69.030 339.900 ;
        RECT 80.430 340.100 81.430 341.100 ;
        RECT 82.030 340.100 83.030 341.100 ;
        RECT 83.630 340.100 84.630 341.100 ;
        RECT 84.830 340.100 85.830 341.100 ;
        RECT 86.430 340.100 87.430 341.100 ;
        RECT 88.030 340.100 89.030 341.100 ;
        RECT 103.630 343.300 104.630 344.300 ;
        RECT 105.340 343.095 105.700 343.475 ;
        RECT 105.970 343.095 106.330 343.475 ;
        RECT 106.570 343.095 106.930 343.475 ;
        RECT 103.630 341.700 104.630 342.700 ;
        RECT 105.340 342.505 105.700 342.885 ;
        RECT 105.970 342.505 106.330 342.885 ;
        RECT 106.570 342.505 106.930 342.885 ;
        RECT 63.630 337.300 64.630 338.300 ;
        RECT 64.830 337.300 65.830 338.300 ;
        RECT 63.630 335.700 64.630 336.700 ;
        RECT 64.830 335.700 65.830 336.700 ;
        RECT 80.430 338.900 81.430 339.900 ;
        RECT 82.030 338.900 83.030 339.900 ;
        RECT 83.630 338.900 84.630 339.900 ;
        RECT 84.830 338.900 85.830 339.900 ;
        RECT 86.430 338.900 87.430 339.900 ;
        RECT 88.030 338.900 89.030 339.900 ;
        RECT 100.430 340.100 101.430 341.100 ;
        RECT 102.030 340.100 103.030 341.100 ;
        RECT 103.630 340.100 104.630 341.100 ;
        RECT 83.630 337.300 84.630 338.300 ;
        RECT 84.830 337.300 85.830 338.300 ;
        RECT 83.630 335.700 84.630 336.700 ;
        RECT 84.830 335.700 85.830 336.700 ;
        RECT 100.430 338.900 101.430 339.900 ;
        RECT 102.030 338.900 103.030 339.900 ;
        RECT 103.630 338.900 104.630 339.900 ;
        RECT 103.630 337.300 104.630 338.300 ;
        RECT 105.340 337.080 105.700 337.460 ;
        RECT 105.970 337.080 106.330 337.460 ;
        RECT 106.570 337.080 106.930 337.460 ;
        RECT 103.630 335.700 104.630 336.700 ;
        RECT 105.340 336.490 105.700 336.870 ;
        RECT 105.970 336.490 106.330 336.870 ;
        RECT 106.570 336.490 106.930 336.870 ;
        RECT 2.520 326.125 2.880 326.505 ;
        RECT 3.130 326.125 3.490 326.505 ;
        RECT 3.760 326.125 4.120 326.505 ;
        RECT 2.520 325.390 2.880 325.770 ;
        RECT 3.130 325.390 3.490 325.770 ;
        RECT 3.760 325.390 4.120 325.770 ;
        RECT 2.520 324.705 2.880 325.085 ;
        RECT 3.130 324.705 3.490 325.085 ;
        RECT 3.760 324.705 4.120 325.085 ;
        RECT 2.515 323.170 2.875 323.550 ;
        RECT 3.145 323.170 3.505 323.550 ;
        RECT 3.745 323.170 4.105 323.550 ;
        RECT 4.830 323.300 5.830 324.300 ;
        RECT 2.515 322.580 2.875 322.960 ;
        RECT 3.145 322.580 3.505 322.960 ;
        RECT 3.745 322.580 4.105 322.960 ;
        RECT 4.830 321.700 5.830 322.700 ;
        RECT 4.830 320.100 5.830 321.100 ;
        RECT 6.430 320.100 7.430 321.100 ;
        RECT 8.030 320.100 9.030 321.100 ;
        RECT 23.630 323.300 24.630 324.300 ;
        RECT 24.830 323.300 25.830 324.300 ;
        RECT 23.630 321.700 24.630 322.700 ;
        RECT 24.830 321.700 25.830 322.700 ;
        RECT 4.830 318.900 5.830 319.900 ;
        RECT 6.430 318.900 7.430 319.900 ;
        RECT 8.030 318.900 9.030 319.900 ;
        RECT 20.430 320.100 21.430 321.100 ;
        RECT 22.030 320.100 23.030 321.100 ;
        RECT 23.630 320.100 24.630 321.100 ;
        RECT 24.830 320.100 25.830 321.100 ;
        RECT 26.430 320.100 27.430 321.100 ;
        RECT 28.030 320.100 29.030 321.100 ;
        RECT 43.630 323.300 44.630 324.300 ;
        RECT 44.830 323.300 45.830 324.300 ;
        RECT 43.630 321.700 44.630 322.700 ;
        RECT 44.830 321.700 45.830 322.700 ;
        RECT 2.515 317.280 2.875 317.660 ;
        RECT 3.145 317.280 3.505 317.660 ;
        RECT 3.745 317.280 4.105 317.660 ;
        RECT 4.830 317.300 5.830 318.300 ;
        RECT 2.515 316.690 2.875 317.070 ;
        RECT 3.145 316.690 3.505 317.070 ;
        RECT 3.745 316.690 4.105 317.070 ;
        RECT 4.830 315.700 5.830 316.700 ;
        RECT 20.430 318.900 21.430 319.900 ;
        RECT 22.030 318.900 23.030 319.900 ;
        RECT 23.630 318.900 24.630 319.900 ;
        RECT 24.830 318.900 25.830 319.900 ;
        RECT 26.430 318.900 27.430 319.900 ;
        RECT 28.030 318.900 29.030 319.900 ;
        RECT 40.430 320.100 41.430 321.100 ;
        RECT 42.030 320.100 43.030 321.100 ;
        RECT 43.630 320.100 44.630 321.100 ;
        RECT 44.830 320.100 45.830 321.100 ;
        RECT 46.430 320.100 47.430 321.100 ;
        RECT 48.030 320.100 49.030 321.100 ;
        RECT 63.630 323.300 64.630 324.300 ;
        RECT 64.830 323.300 65.830 324.300 ;
        RECT 63.630 321.700 64.630 322.700 ;
        RECT 64.830 321.700 65.830 322.700 ;
        RECT 2.520 314.920 2.880 315.300 ;
        RECT 3.130 314.920 3.490 315.300 ;
        RECT 3.760 314.920 4.120 315.300 ;
        RECT 2.520 314.185 2.880 314.565 ;
        RECT 3.130 314.185 3.490 314.565 ;
        RECT 3.760 314.185 4.120 314.565 ;
        RECT 2.520 313.500 2.880 313.880 ;
        RECT 3.130 313.500 3.490 313.880 ;
        RECT 3.760 313.500 4.120 313.880 ;
        RECT 23.630 317.300 24.630 318.300 ;
        RECT 24.830 317.300 25.830 318.300 ;
        RECT 23.630 315.700 24.630 316.700 ;
        RECT 24.830 315.700 25.830 316.700 ;
        RECT 40.430 318.900 41.430 319.900 ;
        RECT 42.030 318.900 43.030 319.900 ;
        RECT 43.630 318.900 44.630 319.900 ;
        RECT 44.830 318.900 45.830 319.900 ;
        RECT 46.430 318.900 47.430 319.900 ;
        RECT 48.030 318.900 49.030 319.900 ;
        RECT 60.430 320.100 61.430 321.100 ;
        RECT 62.030 320.100 63.030 321.100 ;
        RECT 63.630 320.100 64.630 321.100 ;
        RECT 64.830 320.100 65.830 321.100 ;
        RECT 66.430 320.100 67.430 321.100 ;
        RECT 68.030 320.100 69.030 321.100 ;
        RECT 83.630 323.300 84.630 324.300 ;
        RECT 84.830 323.300 85.830 324.300 ;
        RECT 83.630 321.700 84.630 322.700 ;
        RECT 84.830 321.700 85.830 322.700 ;
        RECT 43.630 317.300 44.630 318.300 ;
        RECT 44.830 317.300 45.830 318.300 ;
        RECT 43.630 315.700 44.630 316.700 ;
        RECT 44.830 315.700 45.830 316.700 ;
        RECT 60.430 318.900 61.430 319.900 ;
        RECT 62.030 318.900 63.030 319.900 ;
        RECT 63.630 318.900 64.630 319.900 ;
        RECT 64.830 318.900 65.830 319.900 ;
        RECT 66.430 318.900 67.430 319.900 ;
        RECT 68.030 318.900 69.030 319.900 ;
        RECT 80.430 320.100 81.430 321.100 ;
        RECT 82.030 320.100 83.030 321.100 ;
        RECT 83.630 320.100 84.630 321.100 ;
        RECT 84.830 320.100 85.830 321.100 ;
        RECT 86.430 320.100 87.430 321.100 ;
        RECT 88.030 320.100 89.030 321.100 ;
        RECT 103.630 323.300 104.630 324.300 ;
        RECT 105.340 323.095 105.700 323.475 ;
        RECT 105.970 323.095 106.330 323.475 ;
        RECT 106.570 323.095 106.930 323.475 ;
        RECT 103.630 321.700 104.630 322.700 ;
        RECT 105.340 322.505 105.700 322.885 ;
        RECT 105.970 322.505 106.330 322.885 ;
        RECT 106.570 322.505 106.930 322.885 ;
        RECT 63.630 317.300 64.630 318.300 ;
        RECT 64.830 317.300 65.830 318.300 ;
        RECT 63.630 315.700 64.630 316.700 ;
        RECT 64.830 315.700 65.830 316.700 ;
        RECT 80.430 318.900 81.430 319.900 ;
        RECT 82.030 318.900 83.030 319.900 ;
        RECT 83.630 318.900 84.630 319.900 ;
        RECT 84.830 318.900 85.830 319.900 ;
        RECT 86.430 318.900 87.430 319.900 ;
        RECT 88.030 318.900 89.030 319.900 ;
        RECT 100.430 320.100 101.430 321.100 ;
        RECT 102.030 320.100 103.030 321.100 ;
        RECT 103.630 320.100 104.630 321.100 ;
        RECT 83.630 317.300 84.630 318.300 ;
        RECT 84.830 317.300 85.830 318.300 ;
        RECT 83.630 315.700 84.630 316.700 ;
        RECT 84.830 315.700 85.830 316.700 ;
        RECT 100.430 318.900 101.430 319.900 ;
        RECT 102.030 318.900 103.030 319.900 ;
        RECT 103.630 318.900 104.630 319.900 ;
        RECT 103.630 317.300 104.630 318.300 ;
        RECT 105.340 317.080 105.700 317.460 ;
        RECT 105.970 317.080 106.330 317.460 ;
        RECT 106.570 317.080 106.930 317.460 ;
        RECT 103.630 315.700 104.630 316.700 ;
        RECT 105.340 316.490 105.700 316.870 ;
        RECT 105.970 316.490 106.330 316.870 ;
        RECT 106.570 316.490 106.930 316.870 ;
        RECT 2.520 306.125 2.880 306.505 ;
        RECT 3.130 306.125 3.490 306.505 ;
        RECT 3.760 306.125 4.120 306.505 ;
        RECT 2.520 305.390 2.880 305.770 ;
        RECT 3.130 305.390 3.490 305.770 ;
        RECT 3.760 305.390 4.120 305.770 ;
        RECT 2.520 304.705 2.880 305.085 ;
        RECT 3.130 304.705 3.490 305.085 ;
        RECT 3.760 304.705 4.120 305.085 ;
        RECT 2.515 303.040 2.875 303.420 ;
        RECT 3.145 303.040 3.505 303.420 ;
        RECT 3.745 303.040 4.105 303.420 ;
        RECT 4.830 303.300 5.830 304.300 ;
        RECT 2.515 302.450 2.875 302.830 ;
        RECT 3.145 302.450 3.505 302.830 ;
        RECT 3.745 302.450 4.105 302.830 ;
        RECT 4.830 301.700 5.830 302.700 ;
        RECT 4.830 300.100 5.830 301.100 ;
        RECT 6.430 300.100 7.430 301.100 ;
        RECT 8.030 300.100 9.030 301.100 ;
        RECT 23.630 303.300 24.630 304.300 ;
        RECT 24.830 303.300 25.830 304.300 ;
        RECT 23.630 301.700 24.630 302.700 ;
        RECT 24.830 301.700 25.830 302.700 ;
        RECT 4.830 298.900 5.830 299.900 ;
        RECT 6.430 298.900 7.430 299.900 ;
        RECT 8.030 298.900 9.030 299.900 ;
        RECT 20.430 300.100 21.430 301.100 ;
        RECT 22.030 300.100 23.030 301.100 ;
        RECT 23.630 300.100 24.630 301.100 ;
        RECT 24.830 300.100 25.830 301.100 ;
        RECT 26.430 300.100 27.430 301.100 ;
        RECT 28.030 300.100 29.030 301.100 ;
        RECT 43.630 303.300 44.630 304.300 ;
        RECT 44.830 303.300 45.830 304.300 ;
        RECT 43.630 301.700 44.630 302.700 ;
        RECT 44.830 301.700 45.830 302.700 ;
        RECT 2.515 297.025 2.875 297.405 ;
        RECT 3.145 297.025 3.505 297.405 ;
        RECT 3.745 297.025 4.105 297.405 ;
        RECT 4.830 297.300 5.830 298.300 ;
        RECT 2.515 296.435 2.875 296.815 ;
        RECT 3.145 296.435 3.505 296.815 ;
        RECT 3.745 296.435 4.105 296.815 ;
        RECT 4.830 295.700 5.830 296.700 ;
        RECT 20.430 298.900 21.430 299.900 ;
        RECT 22.030 298.900 23.030 299.900 ;
        RECT 23.630 298.900 24.630 299.900 ;
        RECT 24.830 298.900 25.830 299.900 ;
        RECT 26.430 298.900 27.430 299.900 ;
        RECT 28.030 298.900 29.030 299.900 ;
        RECT 40.430 300.100 41.430 301.100 ;
        RECT 42.030 300.100 43.030 301.100 ;
        RECT 43.630 300.100 44.630 301.100 ;
        RECT 44.830 300.100 45.830 301.100 ;
        RECT 46.430 300.100 47.430 301.100 ;
        RECT 48.030 300.100 49.030 301.100 ;
        RECT 63.630 303.300 64.630 304.300 ;
        RECT 64.830 303.300 65.830 304.300 ;
        RECT 63.630 301.700 64.630 302.700 ;
        RECT 64.830 301.700 65.830 302.700 ;
        RECT 2.520 294.920 2.880 295.300 ;
        RECT 3.130 294.920 3.490 295.300 ;
        RECT 3.760 294.920 4.120 295.300 ;
        RECT 2.520 294.185 2.880 294.565 ;
        RECT 3.130 294.185 3.490 294.565 ;
        RECT 3.760 294.185 4.120 294.565 ;
        RECT 2.520 293.500 2.880 293.880 ;
        RECT 3.130 293.500 3.490 293.880 ;
        RECT 3.760 293.500 4.120 293.880 ;
        RECT 23.630 297.300 24.630 298.300 ;
        RECT 24.830 297.300 25.830 298.300 ;
        RECT 23.630 295.700 24.630 296.700 ;
        RECT 24.830 295.700 25.830 296.700 ;
        RECT 40.430 298.900 41.430 299.900 ;
        RECT 42.030 298.900 43.030 299.900 ;
        RECT 43.630 298.900 44.630 299.900 ;
        RECT 44.830 298.900 45.830 299.900 ;
        RECT 46.430 298.900 47.430 299.900 ;
        RECT 48.030 298.900 49.030 299.900 ;
        RECT 60.430 300.100 61.430 301.100 ;
        RECT 62.030 300.100 63.030 301.100 ;
        RECT 63.630 300.100 64.630 301.100 ;
        RECT 64.830 300.100 65.830 301.100 ;
        RECT 66.430 300.100 67.430 301.100 ;
        RECT 68.030 300.100 69.030 301.100 ;
        RECT 83.630 303.300 84.630 304.300 ;
        RECT 84.830 303.300 85.830 304.300 ;
        RECT 83.630 301.700 84.630 302.700 ;
        RECT 84.830 301.700 85.830 302.700 ;
        RECT 43.630 297.300 44.630 298.300 ;
        RECT 44.830 297.300 45.830 298.300 ;
        RECT 43.630 295.700 44.630 296.700 ;
        RECT 44.830 295.700 45.830 296.700 ;
        RECT 60.430 298.900 61.430 299.900 ;
        RECT 62.030 298.900 63.030 299.900 ;
        RECT 63.630 298.900 64.630 299.900 ;
        RECT 64.830 298.900 65.830 299.900 ;
        RECT 66.430 298.900 67.430 299.900 ;
        RECT 68.030 298.900 69.030 299.900 ;
        RECT 80.430 300.100 81.430 301.100 ;
        RECT 82.030 300.100 83.030 301.100 ;
        RECT 83.630 300.100 84.630 301.100 ;
        RECT 84.830 300.100 85.830 301.100 ;
        RECT 86.430 300.100 87.430 301.100 ;
        RECT 88.030 300.100 89.030 301.100 ;
        RECT 103.630 303.300 104.630 304.300 ;
        RECT 105.340 303.095 105.700 303.475 ;
        RECT 105.970 303.095 106.330 303.475 ;
        RECT 106.570 303.095 106.930 303.475 ;
        RECT 103.630 301.700 104.630 302.700 ;
        RECT 105.340 302.505 105.700 302.885 ;
        RECT 105.970 302.505 106.330 302.885 ;
        RECT 106.570 302.505 106.930 302.885 ;
        RECT 63.630 297.300 64.630 298.300 ;
        RECT 64.830 297.300 65.830 298.300 ;
        RECT 63.630 295.700 64.630 296.700 ;
        RECT 64.830 295.700 65.830 296.700 ;
        RECT 80.430 298.900 81.430 299.900 ;
        RECT 82.030 298.900 83.030 299.900 ;
        RECT 83.630 298.900 84.630 299.900 ;
        RECT 84.830 298.900 85.830 299.900 ;
        RECT 86.430 298.900 87.430 299.900 ;
        RECT 88.030 298.900 89.030 299.900 ;
        RECT 100.430 300.100 101.430 301.100 ;
        RECT 102.030 300.100 103.030 301.100 ;
        RECT 103.630 300.100 104.630 301.100 ;
        RECT 83.630 297.300 84.630 298.300 ;
        RECT 84.830 297.300 85.830 298.300 ;
        RECT 83.630 295.700 84.630 296.700 ;
        RECT 84.830 295.700 85.830 296.700 ;
        RECT 100.430 298.900 101.430 299.900 ;
        RECT 102.030 298.900 103.030 299.900 ;
        RECT 103.630 298.900 104.630 299.900 ;
        RECT 103.630 297.300 104.630 298.300 ;
        RECT 105.340 297.350 105.700 297.730 ;
        RECT 105.970 297.350 106.330 297.730 ;
        RECT 106.570 297.350 106.930 297.730 ;
        RECT 105.340 296.760 105.700 297.140 ;
        RECT 105.970 296.760 106.330 297.140 ;
        RECT 106.570 296.760 106.930 297.140 ;
        RECT 103.630 295.700 104.630 296.700 ;
        RECT 2.520 286.115 2.880 286.495 ;
        RECT 3.130 286.115 3.490 286.495 ;
        RECT 3.760 286.115 4.120 286.495 ;
        RECT 2.520 285.380 2.880 285.760 ;
        RECT 3.130 285.380 3.490 285.760 ;
        RECT 3.760 285.380 4.120 285.760 ;
        RECT 2.520 284.695 2.880 285.075 ;
        RECT 3.130 284.695 3.490 285.075 ;
        RECT 3.760 284.695 4.120 285.075 ;
        RECT 2.515 283.140 2.875 283.520 ;
        RECT 3.145 283.140 3.505 283.520 ;
        RECT 3.745 283.140 4.105 283.520 ;
        RECT 4.830 283.300 5.830 284.300 ;
        RECT 2.515 282.550 2.875 282.930 ;
        RECT 3.145 282.550 3.505 282.930 ;
        RECT 3.745 282.550 4.105 282.930 ;
        RECT 4.830 281.700 5.830 282.700 ;
        RECT 4.830 280.100 5.830 281.100 ;
        RECT 6.430 280.100 7.430 281.100 ;
        RECT 8.030 280.100 9.030 281.100 ;
        RECT 23.630 283.300 24.630 284.300 ;
        RECT 24.830 283.300 25.830 284.300 ;
        RECT 23.630 281.700 24.630 282.700 ;
        RECT 24.830 281.700 25.830 282.700 ;
        RECT 4.830 278.900 5.830 279.900 ;
        RECT 6.430 278.900 7.430 279.900 ;
        RECT 8.030 278.900 9.030 279.900 ;
        RECT 20.430 280.100 21.430 281.100 ;
        RECT 22.030 280.100 23.030 281.100 ;
        RECT 23.630 280.100 24.630 281.100 ;
        RECT 24.830 280.100 25.830 281.100 ;
        RECT 26.430 280.100 27.430 281.100 ;
        RECT 28.030 280.100 29.030 281.100 ;
        RECT 43.630 283.300 44.630 284.300 ;
        RECT 44.830 283.300 45.830 284.300 ;
        RECT 43.630 281.700 44.630 282.700 ;
        RECT 44.830 281.700 45.830 282.700 ;
        RECT 2.515 277.105 2.875 277.485 ;
        RECT 3.145 277.105 3.505 277.485 ;
        RECT 3.745 277.105 4.105 277.485 ;
        RECT 4.830 277.300 5.830 278.300 ;
        RECT 2.515 276.515 2.875 276.895 ;
        RECT 3.145 276.515 3.505 276.895 ;
        RECT 3.745 276.515 4.105 276.895 ;
        RECT 4.830 275.700 5.830 276.700 ;
        RECT 20.430 278.900 21.430 279.900 ;
        RECT 22.030 278.900 23.030 279.900 ;
        RECT 23.630 278.900 24.630 279.900 ;
        RECT 24.830 278.900 25.830 279.900 ;
        RECT 26.430 278.900 27.430 279.900 ;
        RECT 28.030 278.900 29.030 279.900 ;
        RECT 40.430 280.100 41.430 281.100 ;
        RECT 42.030 280.100 43.030 281.100 ;
        RECT 43.630 280.100 44.630 281.100 ;
        RECT 44.830 280.100 45.830 281.100 ;
        RECT 46.430 280.100 47.430 281.100 ;
        RECT 48.030 280.100 49.030 281.100 ;
        RECT 63.630 283.300 64.630 284.300 ;
        RECT 64.830 283.300 65.830 284.300 ;
        RECT 63.630 281.700 64.630 282.700 ;
        RECT 64.830 281.700 65.830 282.700 ;
        RECT 2.520 274.920 2.880 275.300 ;
        RECT 3.130 274.920 3.490 275.300 ;
        RECT 3.760 274.920 4.120 275.300 ;
        RECT 2.520 274.185 2.880 274.565 ;
        RECT 3.130 274.185 3.490 274.565 ;
        RECT 3.760 274.185 4.120 274.565 ;
        RECT 2.520 273.500 2.880 273.880 ;
        RECT 3.130 273.500 3.490 273.880 ;
        RECT 3.760 273.500 4.120 273.880 ;
        RECT 23.630 277.300 24.630 278.300 ;
        RECT 24.830 277.300 25.830 278.300 ;
        RECT 23.630 275.700 24.630 276.700 ;
        RECT 24.830 275.700 25.830 276.700 ;
        RECT 40.430 278.900 41.430 279.900 ;
        RECT 42.030 278.900 43.030 279.900 ;
        RECT 43.630 278.900 44.630 279.900 ;
        RECT 44.830 278.900 45.830 279.900 ;
        RECT 46.430 278.900 47.430 279.900 ;
        RECT 48.030 278.900 49.030 279.900 ;
        RECT 60.430 280.100 61.430 281.100 ;
        RECT 62.030 280.100 63.030 281.100 ;
        RECT 63.630 280.100 64.630 281.100 ;
        RECT 64.830 280.100 65.830 281.100 ;
        RECT 66.430 280.100 67.430 281.100 ;
        RECT 68.030 280.100 69.030 281.100 ;
        RECT 83.630 283.300 84.630 284.300 ;
        RECT 84.830 283.300 85.830 284.300 ;
        RECT 83.630 281.700 84.630 282.700 ;
        RECT 84.830 281.700 85.830 282.700 ;
        RECT 43.630 277.300 44.630 278.300 ;
        RECT 44.830 277.300 45.830 278.300 ;
        RECT 43.630 275.700 44.630 276.700 ;
        RECT 44.830 275.700 45.830 276.700 ;
        RECT 60.430 278.900 61.430 279.900 ;
        RECT 62.030 278.900 63.030 279.900 ;
        RECT 63.630 278.900 64.630 279.900 ;
        RECT 64.830 278.900 65.830 279.900 ;
        RECT 66.430 278.900 67.430 279.900 ;
        RECT 68.030 278.900 69.030 279.900 ;
        RECT 80.430 280.100 81.430 281.100 ;
        RECT 82.030 280.100 83.030 281.100 ;
        RECT 83.630 280.100 84.630 281.100 ;
        RECT 84.830 280.100 85.830 281.100 ;
        RECT 86.430 280.100 87.430 281.100 ;
        RECT 88.030 280.100 89.030 281.100 ;
        RECT 103.630 283.300 104.630 284.300 ;
        RECT 105.340 282.770 105.700 283.150 ;
        RECT 105.970 282.770 106.330 283.150 ;
        RECT 106.570 282.770 106.930 283.150 ;
        RECT 103.630 281.700 104.630 282.700 ;
        RECT 105.340 282.180 105.700 282.560 ;
        RECT 105.970 282.180 106.330 282.560 ;
        RECT 106.570 282.180 106.930 282.560 ;
        RECT 63.630 277.300 64.630 278.300 ;
        RECT 64.830 277.300 65.830 278.300 ;
        RECT 63.630 275.700 64.630 276.700 ;
        RECT 64.830 275.700 65.830 276.700 ;
        RECT 80.430 278.900 81.430 279.900 ;
        RECT 82.030 278.900 83.030 279.900 ;
        RECT 83.630 278.900 84.630 279.900 ;
        RECT 84.830 278.900 85.830 279.900 ;
        RECT 86.430 278.900 87.430 279.900 ;
        RECT 88.030 278.900 89.030 279.900 ;
        RECT 100.430 280.100 101.430 281.100 ;
        RECT 102.030 280.100 103.030 281.100 ;
        RECT 103.630 280.100 104.630 281.100 ;
        RECT 83.630 277.300 84.630 278.300 ;
        RECT 84.830 277.300 85.830 278.300 ;
        RECT 83.630 275.700 84.630 276.700 ;
        RECT 84.830 275.700 85.830 276.700 ;
        RECT 100.430 278.900 101.430 279.900 ;
        RECT 102.030 278.900 103.030 279.900 ;
        RECT 103.630 278.900 104.630 279.900 ;
        RECT 103.630 277.300 104.630 278.300 ;
        RECT 105.340 276.855 105.700 277.235 ;
        RECT 105.970 276.855 106.330 277.235 ;
        RECT 106.570 276.855 106.930 277.235 ;
        RECT 103.630 275.700 104.630 276.700 ;
        RECT 105.340 276.265 105.700 276.645 ;
        RECT 105.970 276.265 106.330 276.645 ;
        RECT 106.570 276.265 106.930 276.645 ;
        RECT 2.520 266.125 2.880 266.505 ;
        RECT 3.130 266.125 3.490 266.505 ;
        RECT 3.760 266.125 4.120 266.505 ;
        RECT 2.520 265.390 2.880 265.770 ;
        RECT 3.130 265.390 3.490 265.770 ;
        RECT 3.760 265.390 4.120 265.770 ;
        RECT 2.520 264.705 2.880 265.085 ;
        RECT 3.130 264.705 3.490 265.085 ;
        RECT 3.760 264.705 4.120 265.085 ;
        RECT 2.515 263.275 2.875 263.655 ;
        RECT 3.145 263.275 3.505 263.655 ;
        RECT 3.745 263.275 4.105 263.655 ;
        RECT 4.830 263.300 5.830 264.300 ;
        RECT 2.515 262.685 2.875 263.065 ;
        RECT 3.145 262.685 3.505 263.065 ;
        RECT 3.745 262.685 4.105 263.065 ;
        RECT 4.830 261.700 5.830 262.700 ;
        RECT 4.830 260.100 5.830 261.100 ;
        RECT 6.430 260.100 7.430 261.100 ;
        RECT 8.030 260.100 9.030 261.100 ;
        RECT 23.630 263.300 24.630 264.300 ;
        RECT 24.830 263.300 25.830 264.300 ;
        RECT 23.630 261.700 24.630 262.700 ;
        RECT 24.830 261.700 25.830 262.700 ;
        RECT 4.830 258.900 5.830 259.900 ;
        RECT 6.430 258.900 7.430 259.900 ;
        RECT 8.030 258.900 9.030 259.900 ;
        RECT 20.430 260.100 21.430 261.100 ;
        RECT 22.030 260.100 23.030 261.100 ;
        RECT 23.630 260.100 24.630 261.100 ;
        RECT 24.830 260.100 25.830 261.100 ;
        RECT 26.430 260.100 27.430 261.100 ;
        RECT 28.030 260.100 29.030 261.100 ;
        RECT 43.630 263.300 44.630 264.300 ;
        RECT 44.830 263.300 45.830 264.300 ;
        RECT 43.630 261.700 44.630 262.700 ;
        RECT 44.830 261.700 45.830 262.700 ;
        RECT 2.515 257.340 2.875 257.720 ;
        RECT 3.145 257.340 3.505 257.720 ;
        RECT 3.745 257.340 4.105 257.720 ;
        RECT 4.830 257.300 5.830 258.300 ;
        RECT 2.515 256.750 2.875 257.130 ;
        RECT 3.145 256.750 3.505 257.130 ;
        RECT 3.745 256.750 4.105 257.130 ;
        RECT 4.830 255.700 5.830 256.700 ;
        RECT 20.430 258.900 21.430 259.900 ;
        RECT 22.030 258.900 23.030 259.900 ;
        RECT 23.630 258.900 24.630 259.900 ;
        RECT 24.830 258.900 25.830 259.900 ;
        RECT 26.430 258.900 27.430 259.900 ;
        RECT 28.030 258.900 29.030 259.900 ;
        RECT 40.430 260.100 41.430 261.100 ;
        RECT 42.030 260.100 43.030 261.100 ;
        RECT 43.630 260.100 44.630 261.100 ;
        RECT 44.830 260.100 45.830 261.100 ;
        RECT 46.430 260.100 47.430 261.100 ;
        RECT 48.030 260.100 49.030 261.100 ;
        RECT 63.630 263.300 64.630 264.300 ;
        RECT 64.830 263.300 65.830 264.300 ;
        RECT 63.630 261.700 64.630 262.700 ;
        RECT 64.830 261.700 65.830 262.700 ;
        RECT 2.520 254.920 2.880 255.300 ;
        RECT 3.130 254.920 3.490 255.300 ;
        RECT 3.760 254.920 4.120 255.300 ;
        RECT 2.520 254.185 2.880 254.565 ;
        RECT 3.130 254.185 3.490 254.565 ;
        RECT 3.760 254.185 4.120 254.565 ;
        RECT 2.520 253.500 2.880 253.880 ;
        RECT 3.130 253.500 3.490 253.880 ;
        RECT 3.760 253.500 4.120 253.880 ;
        RECT 23.630 257.300 24.630 258.300 ;
        RECT 24.830 257.300 25.830 258.300 ;
        RECT 23.630 255.700 24.630 256.700 ;
        RECT 24.830 255.700 25.830 256.700 ;
        RECT 40.430 258.900 41.430 259.900 ;
        RECT 42.030 258.900 43.030 259.900 ;
        RECT 43.630 258.900 44.630 259.900 ;
        RECT 44.830 258.900 45.830 259.900 ;
        RECT 46.430 258.900 47.430 259.900 ;
        RECT 48.030 258.900 49.030 259.900 ;
        RECT 60.430 260.100 61.430 261.100 ;
        RECT 62.030 260.100 63.030 261.100 ;
        RECT 63.630 260.100 64.630 261.100 ;
        RECT 64.830 260.100 65.830 261.100 ;
        RECT 66.430 260.100 67.430 261.100 ;
        RECT 68.030 260.100 69.030 261.100 ;
        RECT 83.630 263.300 84.630 264.300 ;
        RECT 84.830 263.300 85.830 264.300 ;
        RECT 83.630 261.700 84.630 262.700 ;
        RECT 84.830 261.700 85.830 262.700 ;
        RECT 43.630 257.300 44.630 258.300 ;
        RECT 44.830 257.300 45.830 258.300 ;
        RECT 43.630 255.700 44.630 256.700 ;
        RECT 44.830 255.700 45.830 256.700 ;
        RECT 60.430 258.900 61.430 259.900 ;
        RECT 62.030 258.900 63.030 259.900 ;
        RECT 63.630 258.900 64.630 259.900 ;
        RECT 64.830 258.900 65.830 259.900 ;
        RECT 66.430 258.900 67.430 259.900 ;
        RECT 68.030 258.900 69.030 259.900 ;
        RECT 80.430 260.100 81.430 261.100 ;
        RECT 82.030 260.100 83.030 261.100 ;
        RECT 83.630 260.100 84.630 261.100 ;
        RECT 84.830 260.100 85.830 261.100 ;
        RECT 86.430 260.100 87.430 261.100 ;
        RECT 88.030 260.100 89.030 261.100 ;
        RECT 103.630 263.300 104.630 264.300 ;
        RECT 103.630 261.700 104.630 262.700 ;
        RECT 105.340 262.495 105.700 262.875 ;
        RECT 105.970 262.495 106.330 262.875 ;
        RECT 106.570 262.495 106.930 262.875 ;
        RECT 105.340 261.905 105.700 262.285 ;
        RECT 105.970 261.905 106.330 262.285 ;
        RECT 106.570 261.905 106.930 262.285 ;
        RECT 63.630 257.300 64.630 258.300 ;
        RECT 64.830 257.300 65.830 258.300 ;
        RECT 63.630 255.700 64.630 256.700 ;
        RECT 64.830 255.700 65.830 256.700 ;
        RECT 80.430 258.900 81.430 259.900 ;
        RECT 82.030 258.900 83.030 259.900 ;
        RECT 83.630 258.900 84.630 259.900 ;
        RECT 84.830 258.900 85.830 259.900 ;
        RECT 86.430 258.900 87.430 259.900 ;
        RECT 88.030 258.900 89.030 259.900 ;
        RECT 100.430 260.100 101.430 261.100 ;
        RECT 102.030 260.100 103.030 261.100 ;
        RECT 103.630 260.100 104.630 261.100 ;
        RECT 83.630 257.300 84.630 258.300 ;
        RECT 84.830 257.300 85.830 258.300 ;
        RECT 83.630 255.700 84.630 256.700 ;
        RECT 84.830 255.700 85.830 256.700 ;
        RECT 100.430 258.900 101.430 259.900 ;
        RECT 102.030 258.900 103.030 259.900 ;
        RECT 103.630 258.900 104.630 259.900 ;
        RECT 103.630 257.300 104.630 258.300 ;
        RECT 105.340 256.820 105.700 257.200 ;
        RECT 105.970 256.820 106.330 257.200 ;
        RECT 106.570 256.820 106.930 257.200 ;
        RECT 103.630 255.700 104.630 256.700 ;
        RECT 105.340 256.230 105.700 256.610 ;
        RECT 105.970 256.230 106.330 256.610 ;
        RECT 106.570 256.230 106.930 256.610 ;
        RECT 2.520 246.125 2.880 246.505 ;
        RECT 3.130 246.125 3.490 246.505 ;
        RECT 3.760 246.125 4.120 246.505 ;
        RECT 2.520 245.390 2.880 245.770 ;
        RECT 3.130 245.390 3.490 245.770 ;
        RECT 3.760 245.390 4.120 245.770 ;
        RECT 2.520 244.705 2.880 245.085 ;
        RECT 3.130 244.705 3.490 245.085 ;
        RECT 3.760 244.705 4.120 245.085 ;
        RECT 2.515 243.230 2.875 243.610 ;
        RECT 3.145 243.230 3.505 243.610 ;
        RECT 3.745 243.230 4.105 243.610 ;
        RECT 4.830 243.300 5.830 244.300 ;
        RECT 2.515 242.640 2.875 243.020 ;
        RECT 3.145 242.640 3.505 243.020 ;
        RECT 3.745 242.640 4.105 243.020 ;
        RECT 4.830 241.700 5.830 242.700 ;
        RECT 4.830 240.100 5.830 241.100 ;
        RECT 6.430 240.100 7.430 241.100 ;
        RECT 8.030 240.100 9.030 241.100 ;
        RECT 23.630 243.300 24.630 244.300 ;
        RECT 24.830 243.300 25.830 244.300 ;
        RECT 23.630 241.700 24.630 242.700 ;
        RECT 24.830 241.700 25.830 242.700 ;
        RECT 4.830 238.900 5.830 239.900 ;
        RECT 6.430 238.900 7.430 239.900 ;
        RECT 8.030 238.900 9.030 239.900 ;
        RECT 20.430 240.100 21.430 241.100 ;
        RECT 22.030 240.100 23.030 241.100 ;
        RECT 23.630 240.100 24.630 241.100 ;
        RECT 24.830 240.100 25.830 241.100 ;
        RECT 26.430 240.100 27.430 241.100 ;
        RECT 28.030 240.100 29.030 241.100 ;
        RECT 43.630 243.300 44.630 244.300 ;
        RECT 44.830 243.300 45.830 244.300 ;
        RECT 43.630 241.700 44.630 242.700 ;
        RECT 44.830 241.700 45.830 242.700 ;
        RECT 2.515 237.465 2.875 237.845 ;
        RECT 3.145 237.465 3.505 237.845 ;
        RECT 3.745 237.465 4.105 237.845 ;
        RECT 4.830 237.300 5.830 238.300 ;
        RECT 2.515 236.875 2.875 237.255 ;
        RECT 3.145 236.875 3.505 237.255 ;
        RECT 3.745 236.875 4.105 237.255 ;
        RECT 4.830 235.700 5.830 236.700 ;
        RECT 20.430 238.900 21.430 239.900 ;
        RECT 22.030 238.900 23.030 239.900 ;
        RECT 23.630 238.900 24.630 239.900 ;
        RECT 24.830 238.900 25.830 239.900 ;
        RECT 26.430 238.900 27.430 239.900 ;
        RECT 28.030 238.900 29.030 239.900 ;
        RECT 40.430 240.100 41.430 241.100 ;
        RECT 42.030 240.100 43.030 241.100 ;
        RECT 43.630 240.100 44.630 241.100 ;
        RECT 44.830 240.100 45.830 241.100 ;
        RECT 46.430 240.100 47.430 241.100 ;
        RECT 48.030 240.100 49.030 241.100 ;
        RECT 63.630 243.300 64.630 244.300 ;
        RECT 64.830 243.300 65.830 244.300 ;
        RECT 63.630 241.700 64.630 242.700 ;
        RECT 64.830 241.700 65.830 242.700 ;
        RECT 2.520 234.920 2.880 235.300 ;
        RECT 3.130 234.920 3.490 235.300 ;
        RECT 3.760 234.920 4.120 235.300 ;
        RECT 2.520 234.185 2.880 234.565 ;
        RECT 3.130 234.185 3.490 234.565 ;
        RECT 3.760 234.185 4.120 234.565 ;
        RECT 2.520 233.500 2.880 233.880 ;
        RECT 3.130 233.500 3.490 233.880 ;
        RECT 3.760 233.500 4.120 233.880 ;
        RECT 23.630 237.300 24.630 238.300 ;
        RECT 24.830 237.300 25.830 238.300 ;
        RECT 23.630 235.700 24.630 236.700 ;
        RECT 24.830 235.700 25.830 236.700 ;
        RECT 40.430 238.900 41.430 239.900 ;
        RECT 42.030 238.900 43.030 239.900 ;
        RECT 43.630 238.900 44.630 239.900 ;
        RECT 44.830 238.900 45.830 239.900 ;
        RECT 46.430 238.900 47.430 239.900 ;
        RECT 48.030 238.900 49.030 239.900 ;
        RECT 60.430 240.100 61.430 241.100 ;
        RECT 62.030 240.100 63.030 241.100 ;
        RECT 63.630 240.100 64.630 241.100 ;
        RECT 64.830 240.100 65.830 241.100 ;
        RECT 66.430 240.100 67.430 241.100 ;
        RECT 68.030 240.100 69.030 241.100 ;
        RECT 83.630 243.300 84.630 244.300 ;
        RECT 84.830 243.300 85.830 244.300 ;
        RECT 83.630 241.700 84.630 242.700 ;
        RECT 84.830 241.700 85.830 242.700 ;
        RECT 43.630 237.300 44.630 238.300 ;
        RECT 44.830 237.300 45.830 238.300 ;
        RECT 43.630 235.700 44.630 236.700 ;
        RECT 44.830 235.700 45.830 236.700 ;
        RECT 60.430 238.900 61.430 239.900 ;
        RECT 62.030 238.900 63.030 239.900 ;
        RECT 63.630 238.900 64.630 239.900 ;
        RECT 64.830 238.900 65.830 239.900 ;
        RECT 66.430 238.900 67.430 239.900 ;
        RECT 68.030 238.900 69.030 239.900 ;
        RECT 80.430 240.100 81.430 241.100 ;
        RECT 82.030 240.100 83.030 241.100 ;
        RECT 83.630 240.100 84.630 241.100 ;
        RECT 84.830 240.100 85.830 241.100 ;
        RECT 86.430 240.100 87.430 241.100 ;
        RECT 88.030 240.100 89.030 241.100 ;
        RECT 103.630 243.300 104.630 244.300 ;
        RECT 105.340 243.025 105.700 243.405 ;
        RECT 105.970 243.025 106.330 243.405 ;
        RECT 106.570 243.025 106.930 243.405 ;
        RECT 103.630 241.700 104.630 242.700 ;
        RECT 105.340 242.435 105.700 242.815 ;
        RECT 105.970 242.435 106.330 242.815 ;
        RECT 106.570 242.435 106.930 242.815 ;
        RECT 63.630 237.300 64.630 238.300 ;
        RECT 64.830 237.300 65.830 238.300 ;
        RECT 63.630 235.700 64.630 236.700 ;
        RECT 64.830 235.700 65.830 236.700 ;
        RECT 80.430 238.900 81.430 239.900 ;
        RECT 82.030 238.900 83.030 239.900 ;
        RECT 83.630 238.900 84.630 239.900 ;
        RECT 84.830 238.900 85.830 239.900 ;
        RECT 86.430 238.900 87.430 239.900 ;
        RECT 88.030 238.900 89.030 239.900 ;
        RECT 100.430 240.100 101.430 241.100 ;
        RECT 102.030 240.100 103.030 241.100 ;
        RECT 103.630 240.100 104.630 241.100 ;
        RECT 83.630 237.300 84.630 238.300 ;
        RECT 84.830 237.300 85.830 238.300 ;
        RECT 83.630 235.700 84.630 236.700 ;
        RECT 84.830 235.700 85.830 236.700 ;
        RECT 100.430 238.900 101.430 239.900 ;
        RECT 102.030 238.900 103.030 239.900 ;
        RECT 103.630 238.900 104.630 239.900 ;
        RECT 103.630 237.300 104.630 238.300 ;
        RECT 105.340 237.260 105.700 237.640 ;
        RECT 105.970 237.260 106.330 237.640 ;
        RECT 106.570 237.260 106.930 237.640 ;
        RECT 103.630 235.700 104.630 236.700 ;
        RECT 105.340 236.670 105.700 237.050 ;
        RECT 105.970 236.670 106.330 237.050 ;
        RECT 106.570 236.670 106.930 237.050 ;
        RECT 2.520 226.120 2.880 226.500 ;
        RECT 3.130 226.120 3.490 226.500 ;
        RECT 3.760 226.120 4.120 226.500 ;
        RECT 2.520 225.385 2.880 225.765 ;
        RECT 3.130 225.385 3.490 225.765 ;
        RECT 3.760 225.385 4.120 225.765 ;
        RECT 2.520 224.700 2.880 225.080 ;
        RECT 3.130 224.700 3.490 225.080 ;
        RECT 3.760 224.700 4.120 225.080 ;
        RECT 4.830 223.300 5.830 224.300 ;
        RECT 2.515 222.165 2.875 222.545 ;
        RECT 3.145 222.165 3.505 222.545 ;
        RECT 3.745 222.165 4.105 222.545 ;
        RECT 2.515 221.575 2.875 221.955 ;
        RECT 3.145 221.575 3.505 221.955 ;
        RECT 3.745 221.575 4.105 221.955 ;
        RECT 4.830 221.700 5.830 222.700 ;
        RECT 4.830 220.100 5.830 221.100 ;
        RECT 6.430 220.100 7.430 221.100 ;
        RECT 8.030 220.100 9.030 221.100 ;
        RECT 23.630 223.300 24.630 224.300 ;
        RECT 24.830 223.300 25.830 224.300 ;
        RECT 23.630 221.700 24.630 222.700 ;
        RECT 24.830 221.700 25.830 222.700 ;
        RECT 20.430 220.100 21.430 221.100 ;
        RECT 22.030 220.100 23.030 221.100 ;
        RECT 23.630 220.100 24.630 221.100 ;
        RECT 24.830 220.100 25.830 221.100 ;
        RECT 26.430 220.100 27.430 221.100 ;
        RECT 28.030 220.100 29.030 221.100 ;
        RECT 43.630 223.300 44.630 224.300 ;
        RECT 44.830 223.300 45.830 224.300 ;
        RECT 43.630 221.700 44.630 222.700 ;
        RECT 44.830 221.700 45.830 222.700 ;
        RECT 40.430 220.100 41.430 221.100 ;
        RECT 42.030 220.100 43.030 221.100 ;
        RECT 43.630 220.100 44.630 221.100 ;
        RECT 44.830 220.100 45.830 221.100 ;
        RECT 46.430 220.100 47.430 221.100 ;
        RECT 48.030 220.100 49.030 221.100 ;
        RECT 63.630 223.300 64.630 224.300 ;
        RECT 64.830 223.300 65.830 224.300 ;
        RECT 63.630 221.700 64.630 222.700 ;
        RECT 64.830 221.700 65.830 222.700 ;
        RECT 60.430 220.100 61.430 221.100 ;
        RECT 62.030 220.100 63.030 221.100 ;
        RECT 63.630 220.100 64.630 221.100 ;
        RECT 64.830 220.100 65.830 221.100 ;
        RECT 66.430 220.100 67.430 221.100 ;
        RECT 68.030 220.100 69.030 221.100 ;
        RECT 83.630 223.300 84.630 224.300 ;
        RECT 84.830 223.300 85.830 224.300 ;
        RECT 83.630 221.700 84.630 222.700 ;
        RECT 84.830 221.700 85.830 222.700 ;
        RECT 80.430 220.100 81.430 221.100 ;
        RECT 82.030 220.100 83.030 221.100 ;
        RECT 83.630 220.100 84.630 221.100 ;
        RECT 84.830 220.100 85.830 221.100 ;
        RECT 86.430 220.100 87.430 221.100 ;
        RECT 88.030 220.100 89.030 221.100 ;
        RECT 103.630 223.300 104.630 224.300 ;
        RECT 103.630 221.700 104.630 222.700 ;
        RECT 105.340 221.680 105.700 222.060 ;
        RECT 105.970 221.680 106.330 222.060 ;
        RECT 106.570 221.680 106.930 222.060 ;
        RECT 100.430 220.100 101.430 221.100 ;
        RECT 102.030 220.100 103.030 221.100 ;
        RECT 103.630 220.100 104.630 221.100 ;
        RECT 105.340 221.090 105.700 221.470 ;
        RECT 105.970 221.090 106.330 221.470 ;
        RECT 106.570 221.090 106.930 221.470 ;
        RECT 2.395 195.260 2.805 195.650 ;
        RECT 2.965 195.260 3.375 195.650 ;
        RECT 3.535 195.260 3.945 195.650 ;
        RECT 2.395 189.820 2.805 190.210 ;
        RECT 2.965 189.820 3.375 190.210 ;
        RECT 3.535 189.820 3.945 190.210 ;
        RECT 2.395 184.380 2.805 184.770 ;
        RECT 2.965 184.380 3.375 184.770 ;
        RECT 3.535 184.380 3.945 184.770 ;
        RECT 42.735 181.560 43.735 182.560 ;
        RECT 44.335 181.560 45.335 182.560 ;
        RECT 45.935 181.560 46.935 182.560 ;
        RECT 42.735 179.960 43.735 180.960 ;
        RECT 42.735 178.360 43.735 179.360 ;
        RECT 58.335 181.560 59.335 182.560 ;
        RECT 59.935 181.560 60.935 182.560 ;
        RECT 61.535 181.560 62.535 182.560 ;
        RECT 62.735 181.560 63.735 182.560 ;
        RECT 64.335 181.560 65.335 182.560 ;
        RECT 65.935 181.560 66.935 182.560 ;
        RECT 61.535 179.960 62.535 180.960 ;
        RECT 62.735 179.960 63.735 180.960 ;
        RECT 61.535 178.360 62.535 179.360 ;
        RECT 62.735 178.360 63.735 179.360 ;
        RECT 78.335 181.560 79.335 182.560 ;
        RECT 79.935 181.560 80.935 182.560 ;
        RECT 81.535 181.560 82.535 182.560 ;
        RECT 82.735 181.560 83.735 182.560 ;
        RECT 84.335 181.560 85.335 182.560 ;
        RECT 85.935 181.560 86.935 182.560 ;
        RECT 81.535 179.960 82.535 180.960 ;
        RECT 82.735 179.960 83.735 180.960 ;
        RECT 81.535 178.360 82.535 179.360 ;
        RECT 82.735 178.360 83.735 179.360 ;
        RECT 98.335 181.560 99.335 182.560 ;
        RECT 99.935 181.560 100.935 182.560 ;
        RECT 101.535 181.560 102.535 182.560 ;
        RECT 101.535 179.960 102.535 180.960 ;
        RECT 105.305 180.460 105.705 180.860 ;
        RECT 105.930 180.460 106.330 180.860 ;
        RECT 106.555 180.460 106.955 180.860 ;
        RECT 105.300 179.860 105.700 180.260 ;
        RECT 105.925 179.860 106.325 180.260 ;
        RECT 106.550 179.860 106.950 180.260 ;
        RECT 101.535 178.360 102.535 179.360 ;
        RECT 105.345 177.580 105.705 177.960 ;
        RECT 105.955 177.580 106.315 177.960 ;
        RECT 106.585 177.580 106.945 177.960 ;
        RECT 105.345 176.845 105.705 177.225 ;
        RECT 105.955 176.845 106.315 177.225 ;
        RECT 106.585 176.845 106.945 177.225 ;
        RECT 105.345 176.160 105.705 176.540 ;
        RECT 105.955 176.160 106.315 176.540 ;
        RECT 106.585 176.160 106.945 176.540 ;
        RECT 42.735 165.960 43.735 166.960 ;
        RECT 42.735 164.360 43.735 165.360 ;
        RECT 42.735 162.760 43.735 163.760 ;
        RECT 44.335 162.760 45.335 163.760 ;
        RECT 45.935 162.760 46.935 163.760 ;
        RECT 61.535 165.960 62.535 166.960 ;
        RECT 62.735 165.960 63.735 166.960 ;
        RECT 61.535 164.360 62.535 165.360 ;
        RECT 62.735 164.360 63.735 165.360 ;
        RECT 58.335 162.760 59.335 163.760 ;
        RECT 59.935 162.760 60.935 163.760 ;
        RECT 61.535 162.760 62.535 163.760 ;
        RECT 62.735 162.760 63.735 163.760 ;
        RECT 64.335 162.760 65.335 163.760 ;
        RECT 65.935 162.760 66.935 163.760 ;
        RECT 81.535 165.960 82.535 166.960 ;
        RECT 82.735 165.960 83.735 166.960 ;
        RECT 81.535 164.360 82.535 165.360 ;
        RECT 82.735 164.360 83.735 165.360 ;
        RECT 105.345 168.780 105.705 169.160 ;
        RECT 105.955 168.780 106.315 169.160 ;
        RECT 106.585 168.780 106.945 169.160 ;
        RECT 105.345 168.045 105.705 168.425 ;
        RECT 105.955 168.045 106.315 168.425 ;
        RECT 106.585 168.045 106.945 168.425 ;
        RECT 105.345 167.360 105.705 167.740 ;
        RECT 105.955 167.360 106.315 167.740 ;
        RECT 106.585 167.360 106.945 167.740 ;
        RECT 78.335 162.760 79.335 163.760 ;
        RECT 79.935 162.760 80.935 163.760 ;
        RECT 81.535 162.760 82.535 163.760 ;
        RECT 82.735 162.760 83.735 163.760 ;
        RECT 84.335 162.760 85.335 163.760 ;
        RECT 85.935 162.760 86.935 163.760 ;
        RECT 101.535 165.960 102.535 166.960 ;
        RECT 101.535 164.360 102.535 165.360 ;
        RECT 105.300 165.185 105.700 165.585 ;
        RECT 105.925 165.185 106.325 165.585 ;
        RECT 106.550 165.185 106.950 165.585 ;
        RECT 105.295 164.585 105.695 164.985 ;
        RECT 105.920 164.585 106.320 164.985 ;
        RECT 106.545 164.585 106.945 164.985 ;
        RECT 98.335 162.760 99.335 163.760 ;
        RECT 99.935 162.760 100.935 163.760 ;
        RECT 101.535 162.760 102.535 163.760 ;
        RECT 2.515 161.130 2.875 161.510 ;
        RECT 3.145 161.130 3.505 161.510 ;
        RECT 3.745 161.130 4.105 161.510 ;
        RECT 105.340 161.130 105.700 161.510 ;
        RECT 105.970 161.130 106.330 161.510 ;
        RECT 106.570 161.130 106.930 161.510 ;
        RECT 2.515 160.540 2.875 160.920 ;
        RECT 3.145 160.540 3.505 160.920 ;
        RECT 3.745 160.540 4.105 160.920 ;
        RECT 105.340 160.540 105.700 160.920 ;
        RECT 105.970 160.540 106.330 160.920 ;
        RECT 106.570 160.540 106.930 160.920 ;
        RECT 4.830 158.900 5.830 159.900 ;
        RECT 6.430 158.900 7.430 159.900 ;
        RECT 8.030 158.900 9.030 159.900 ;
        RECT 2.515 157.220 2.875 157.600 ;
        RECT 3.145 157.220 3.505 157.600 ;
        RECT 3.745 157.220 4.105 157.600 ;
        RECT 4.830 157.300 5.830 158.300 ;
        RECT 2.515 156.630 2.875 157.010 ;
        RECT 3.145 156.630 3.505 157.010 ;
        RECT 3.745 156.630 4.105 157.010 ;
        RECT 4.830 155.700 5.830 156.700 ;
        RECT 20.430 158.900 21.430 159.900 ;
        RECT 22.030 158.900 23.030 159.900 ;
        RECT 23.630 158.900 24.630 159.900 ;
        RECT 24.830 158.900 25.830 159.900 ;
        RECT 26.430 158.900 27.430 159.900 ;
        RECT 28.030 158.900 29.030 159.900 ;
        RECT 2.520 154.925 2.880 155.305 ;
        RECT 3.130 154.925 3.490 155.305 ;
        RECT 3.760 154.925 4.120 155.305 ;
        RECT 2.520 154.190 2.880 154.570 ;
        RECT 3.130 154.190 3.490 154.570 ;
        RECT 3.760 154.190 4.120 154.570 ;
        RECT 2.520 153.505 2.880 153.885 ;
        RECT 3.130 153.505 3.490 153.885 ;
        RECT 3.760 153.505 4.120 153.885 ;
        RECT 23.630 157.300 24.630 158.300 ;
        RECT 24.830 157.300 25.830 158.300 ;
        RECT 23.630 155.700 24.630 156.700 ;
        RECT 24.830 155.700 25.830 156.700 ;
        RECT 40.430 158.900 41.430 159.900 ;
        RECT 42.030 158.900 43.030 159.900 ;
        RECT 43.630 158.900 44.630 159.900 ;
        RECT 44.830 158.900 45.830 159.900 ;
        RECT 46.430 158.900 47.430 159.900 ;
        RECT 48.030 158.900 49.030 159.900 ;
        RECT 43.630 157.300 44.630 158.300 ;
        RECT 44.830 157.300 45.830 158.300 ;
        RECT 43.630 155.700 44.630 156.700 ;
        RECT 44.830 155.700 45.830 156.700 ;
        RECT 60.430 158.900 61.430 159.900 ;
        RECT 62.030 158.900 63.030 159.900 ;
        RECT 63.630 158.900 64.630 159.900 ;
        RECT 64.830 158.900 65.830 159.900 ;
        RECT 66.430 158.900 67.430 159.900 ;
        RECT 68.030 158.900 69.030 159.900 ;
        RECT 63.630 157.300 64.630 158.300 ;
        RECT 64.830 157.300 65.830 158.300 ;
        RECT 63.630 155.700 64.630 156.700 ;
        RECT 64.830 155.700 65.830 156.700 ;
        RECT 80.430 158.900 81.430 159.900 ;
        RECT 82.030 158.900 83.030 159.900 ;
        RECT 83.630 158.900 84.630 159.900 ;
        RECT 84.830 158.900 85.830 159.900 ;
        RECT 86.430 158.900 87.430 159.900 ;
        RECT 88.030 158.900 89.030 159.900 ;
        RECT 83.630 157.300 84.630 158.300 ;
        RECT 84.830 157.300 85.830 158.300 ;
        RECT 83.630 155.700 84.630 156.700 ;
        RECT 84.830 155.700 85.830 156.700 ;
        RECT 100.430 158.900 101.430 159.900 ;
        RECT 102.030 158.900 103.030 159.900 ;
        RECT 103.630 158.900 104.630 159.900 ;
        RECT 103.630 157.300 104.630 158.300 ;
        RECT 105.340 157.220 105.700 157.600 ;
        RECT 105.970 157.220 106.330 157.600 ;
        RECT 106.570 157.220 106.930 157.600 ;
        RECT 103.630 155.700 104.630 156.700 ;
        RECT 105.340 156.630 105.700 157.010 ;
        RECT 105.970 156.630 106.330 157.010 ;
        RECT 106.570 156.630 106.930 157.010 ;
        RECT 2.520 146.090 2.880 146.470 ;
        RECT 3.130 146.090 3.490 146.470 ;
        RECT 3.760 146.090 4.120 146.470 ;
        RECT 2.520 145.355 2.880 145.735 ;
        RECT 3.130 145.355 3.490 145.735 ;
        RECT 3.760 145.355 4.120 145.735 ;
        RECT 2.520 144.670 2.880 145.050 ;
        RECT 3.130 144.670 3.490 145.050 ;
        RECT 3.760 144.670 4.120 145.050 ;
        RECT 4.830 143.300 5.830 144.300 ;
        RECT 2.515 142.660 2.875 143.040 ;
        RECT 3.145 142.660 3.505 143.040 ;
        RECT 3.745 142.660 4.105 143.040 ;
        RECT 2.515 142.070 2.875 142.450 ;
        RECT 3.145 142.070 3.505 142.450 ;
        RECT 3.745 142.070 4.105 142.450 ;
        RECT 4.830 141.700 5.830 142.700 ;
        RECT 4.830 140.100 5.830 141.100 ;
        RECT 6.430 140.100 7.430 141.100 ;
        RECT 8.030 140.100 9.030 141.100 ;
        RECT 23.630 143.300 24.630 144.300 ;
        RECT 24.830 143.300 25.830 144.300 ;
        RECT 23.630 141.700 24.630 142.700 ;
        RECT 24.830 141.700 25.830 142.700 ;
        RECT 4.830 138.900 5.830 139.900 ;
        RECT 6.430 138.900 7.430 139.900 ;
        RECT 8.030 138.900 9.030 139.900 ;
        RECT 20.430 140.100 21.430 141.100 ;
        RECT 22.030 140.100 23.030 141.100 ;
        RECT 23.630 140.100 24.630 141.100 ;
        RECT 24.830 140.100 25.830 141.100 ;
        RECT 26.430 140.100 27.430 141.100 ;
        RECT 28.030 140.100 29.030 141.100 ;
        RECT 43.630 143.300 44.630 144.300 ;
        RECT 44.830 143.300 45.830 144.300 ;
        RECT 43.630 141.700 44.630 142.700 ;
        RECT 44.830 141.700 45.830 142.700 ;
        RECT 2.515 137.640 2.875 138.020 ;
        RECT 3.145 137.640 3.505 138.020 ;
        RECT 3.745 137.640 4.105 138.020 ;
        RECT 2.515 137.050 2.875 137.430 ;
        RECT 3.145 137.050 3.505 137.430 ;
        RECT 3.745 137.050 4.105 137.430 ;
        RECT 4.830 137.300 5.830 138.300 ;
        RECT 4.830 135.700 5.830 136.700 ;
        RECT 20.430 138.900 21.430 139.900 ;
        RECT 22.030 138.900 23.030 139.900 ;
        RECT 23.630 138.900 24.630 139.900 ;
        RECT 24.830 138.900 25.830 139.900 ;
        RECT 26.430 138.900 27.430 139.900 ;
        RECT 28.030 138.900 29.030 139.900 ;
        RECT 40.430 140.100 41.430 141.100 ;
        RECT 42.030 140.100 43.030 141.100 ;
        RECT 43.630 140.100 44.630 141.100 ;
        RECT 44.830 140.100 45.830 141.100 ;
        RECT 46.430 140.100 47.430 141.100 ;
        RECT 48.030 140.100 49.030 141.100 ;
        RECT 63.630 143.300 64.630 144.300 ;
        RECT 64.830 143.300 65.830 144.300 ;
        RECT 63.630 141.700 64.630 142.700 ;
        RECT 64.830 141.700 65.830 142.700 ;
        RECT 2.520 134.920 2.880 135.300 ;
        RECT 3.130 134.920 3.490 135.300 ;
        RECT 3.760 134.920 4.120 135.300 ;
        RECT 2.520 134.185 2.880 134.565 ;
        RECT 3.130 134.185 3.490 134.565 ;
        RECT 3.760 134.185 4.120 134.565 ;
        RECT 2.520 133.500 2.880 133.880 ;
        RECT 3.130 133.500 3.490 133.880 ;
        RECT 3.760 133.500 4.120 133.880 ;
        RECT 23.630 137.300 24.630 138.300 ;
        RECT 24.830 137.300 25.830 138.300 ;
        RECT 23.630 135.700 24.630 136.700 ;
        RECT 24.830 135.700 25.830 136.700 ;
        RECT 40.430 138.900 41.430 139.900 ;
        RECT 42.030 138.900 43.030 139.900 ;
        RECT 43.630 138.900 44.630 139.900 ;
        RECT 44.830 138.900 45.830 139.900 ;
        RECT 46.430 138.900 47.430 139.900 ;
        RECT 48.030 138.900 49.030 139.900 ;
        RECT 60.430 140.100 61.430 141.100 ;
        RECT 62.030 140.100 63.030 141.100 ;
        RECT 63.630 140.100 64.630 141.100 ;
        RECT 64.830 140.100 65.830 141.100 ;
        RECT 66.430 140.100 67.430 141.100 ;
        RECT 68.030 140.100 69.030 141.100 ;
        RECT 83.630 143.300 84.630 144.300 ;
        RECT 84.830 143.300 85.830 144.300 ;
        RECT 83.630 141.700 84.630 142.700 ;
        RECT 84.830 141.700 85.830 142.700 ;
        RECT 43.630 137.300 44.630 138.300 ;
        RECT 44.830 137.300 45.830 138.300 ;
        RECT 43.630 135.700 44.630 136.700 ;
        RECT 44.830 135.700 45.830 136.700 ;
        RECT 60.430 138.900 61.430 139.900 ;
        RECT 62.030 138.900 63.030 139.900 ;
        RECT 63.630 138.900 64.630 139.900 ;
        RECT 64.830 138.900 65.830 139.900 ;
        RECT 66.430 138.900 67.430 139.900 ;
        RECT 68.030 138.900 69.030 139.900 ;
        RECT 80.430 140.100 81.430 141.100 ;
        RECT 82.030 140.100 83.030 141.100 ;
        RECT 83.630 140.100 84.630 141.100 ;
        RECT 84.830 140.100 85.830 141.100 ;
        RECT 86.430 140.100 87.430 141.100 ;
        RECT 88.030 140.100 89.030 141.100 ;
        RECT 103.630 143.300 104.630 144.300 ;
        RECT 103.630 141.700 104.630 142.700 ;
        RECT 105.340 142.415 105.700 142.795 ;
        RECT 105.970 142.415 106.330 142.795 ;
        RECT 106.570 142.415 106.930 142.795 ;
        RECT 105.340 141.825 105.700 142.205 ;
        RECT 105.970 141.825 106.330 142.205 ;
        RECT 106.570 141.825 106.930 142.205 ;
        RECT 63.630 137.300 64.630 138.300 ;
        RECT 64.830 137.300 65.830 138.300 ;
        RECT 63.630 135.700 64.630 136.700 ;
        RECT 64.830 135.700 65.830 136.700 ;
        RECT 80.430 138.900 81.430 139.900 ;
        RECT 82.030 138.900 83.030 139.900 ;
        RECT 83.630 138.900 84.630 139.900 ;
        RECT 84.830 138.900 85.830 139.900 ;
        RECT 86.430 138.900 87.430 139.900 ;
        RECT 88.030 138.900 89.030 139.900 ;
        RECT 100.430 140.100 101.430 141.100 ;
        RECT 102.030 140.100 103.030 141.100 ;
        RECT 103.630 140.100 104.630 141.100 ;
        RECT 83.630 137.300 84.630 138.300 ;
        RECT 84.830 137.300 85.830 138.300 ;
        RECT 83.630 135.700 84.630 136.700 ;
        RECT 84.830 135.700 85.830 136.700 ;
        RECT 100.430 138.900 101.430 139.900 ;
        RECT 102.030 138.900 103.030 139.900 ;
        RECT 103.630 138.900 104.630 139.900 ;
        RECT 103.630 137.300 104.630 138.300 ;
        RECT 105.340 136.830 105.700 137.210 ;
        RECT 105.970 136.830 106.330 137.210 ;
        RECT 106.570 136.830 106.930 137.210 ;
        RECT 103.630 135.700 104.630 136.700 ;
        RECT 105.340 136.240 105.700 136.620 ;
        RECT 105.970 136.240 106.330 136.620 ;
        RECT 106.570 136.240 106.930 136.620 ;
        RECT 2.520 126.120 2.880 126.500 ;
        RECT 3.130 126.120 3.490 126.500 ;
        RECT 3.760 126.120 4.120 126.500 ;
        RECT 2.520 125.385 2.880 125.765 ;
        RECT 3.130 125.385 3.490 125.765 ;
        RECT 3.760 125.385 4.120 125.765 ;
        RECT 2.520 124.700 2.880 125.080 ;
        RECT 3.130 124.700 3.490 125.080 ;
        RECT 3.760 124.700 4.120 125.080 ;
        RECT 4.830 123.300 5.830 124.300 ;
        RECT 2.515 122.750 2.875 123.130 ;
        RECT 3.145 122.750 3.505 123.130 ;
        RECT 3.745 122.750 4.105 123.130 ;
        RECT 2.515 122.160 2.875 122.540 ;
        RECT 3.145 122.160 3.505 122.540 ;
        RECT 3.745 122.160 4.105 122.540 ;
        RECT 4.830 121.700 5.830 122.700 ;
        RECT 4.830 120.100 5.830 121.100 ;
        RECT 6.430 120.100 7.430 121.100 ;
        RECT 8.030 120.100 9.030 121.100 ;
        RECT 23.630 123.300 24.630 124.300 ;
        RECT 24.830 123.300 25.830 124.300 ;
        RECT 23.630 121.700 24.630 122.700 ;
        RECT 24.830 121.700 25.830 122.700 ;
        RECT 4.830 118.900 5.830 119.900 ;
        RECT 6.430 118.900 7.430 119.900 ;
        RECT 8.030 118.900 9.030 119.900 ;
        RECT 20.430 120.100 21.430 121.100 ;
        RECT 22.030 120.100 23.030 121.100 ;
        RECT 23.630 120.100 24.630 121.100 ;
        RECT 24.830 120.100 25.830 121.100 ;
        RECT 26.430 120.100 27.430 121.100 ;
        RECT 28.030 120.100 29.030 121.100 ;
        RECT 43.630 123.300 44.630 124.300 ;
        RECT 44.830 123.300 45.830 124.300 ;
        RECT 43.630 121.700 44.630 122.700 ;
        RECT 44.830 121.700 45.830 122.700 ;
        RECT 2.515 117.340 2.875 117.720 ;
        RECT 3.145 117.340 3.505 117.720 ;
        RECT 3.745 117.340 4.105 117.720 ;
        RECT 4.830 117.300 5.830 118.300 ;
        RECT 2.515 116.750 2.875 117.130 ;
        RECT 3.145 116.750 3.505 117.130 ;
        RECT 3.745 116.750 4.105 117.130 ;
        RECT 4.830 115.700 5.830 116.700 ;
        RECT 20.430 118.900 21.430 119.900 ;
        RECT 22.030 118.900 23.030 119.900 ;
        RECT 23.630 118.900 24.630 119.900 ;
        RECT 24.830 118.900 25.830 119.900 ;
        RECT 26.430 118.900 27.430 119.900 ;
        RECT 28.030 118.900 29.030 119.900 ;
        RECT 40.430 120.100 41.430 121.100 ;
        RECT 42.030 120.100 43.030 121.100 ;
        RECT 43.630 120.100 44.630 121.100 ;
        RECT 44.830 120.100 45.830 121.100 ;
        RECT 46.430 120.100 47.430 121.100 ;
        RECT 48.030 120.100 49.030 121.100 ;
        RECT 63.630 123.300 64.630 124.300 ;
        RECT 64.830 123.300 65.830 124.300 ;
        RECT 63.630 121.700 64.630 122.700 ;
        RECT 64.830 121.700 65.830 122.700 ;
        RECT 2.520 114.920 2.880 115.300 ;
        RECT 3.130 114.920 3.490 115.300 ;
        RECT 3.760 114.920 4.120 115.300 ;
        RECT 2.520 114.185 2.880 114.565 ;
        RECT 3.130 114.185 3.490 114.565 ;
        RECT 3.760 114.185 4.120 114.565 ;
        RECT 2.520 113.500 2.880 113.880 ;
        RECT 3.130 113.500 3.490 113.880 ;
        RECT 3.760 113.500 4.120 113.880 ;
        RECT 23.630 117.300 24.630 118.300 ;
        RECT 24.830 117.300 25.830 118.300 ;
        RECT 23.630 115.700 24.630 116.700 ;
        RECT 24.830 115.700 25.830 116.700 ;
        RECT 40.430 118.900 41.430 119.900 ;
        RECT 42.030 118.900 43.030 119.900 ;
        RECT 43.630 118.900 44.630 119.900 ;
        RECT 44.830 118.900 45.830 119.900 ;
        RECT 46.430 118.900 47.430 119.900 ;
        RECT 48.030 118.900 49.030 119.900 ;
        RECT 60.430 120.100 61.430 121.100 ;
        RECT 62.030 120.100 63.030 121.100 ;
        RECT 63.630 120.100 64.630 121.100 ;
        RECT 64.830 120.100 65.830 121.100 ;
        RECT 66.430 120.100 67.430 121.100 ;
        RECT 68.030 120.100 69.030 121.100 ;
        RECT 83.630 123.300 84.630 124.300 ;
        RECT 84.830 123.300 85.830 124.300 ;
        RECT 83.630 121.700 84.630 122.700 ;
        RECT 84.830 121.700 85.830 122.700 ;
        RECT 43.630 117.300 44.630 118.300 ;
        RECT 44.830 117.300 45.830 118.300 ;
        RECT 43.630 115.700 44.630 116.700 ;
        RECT 44.830 115.700 45.830 116.700 ;
        RECT 60.430 118.900 61.430 119.900 ;
        RECT 62.030 118.900 63.030 119.900 ;
        RECT 63.630 118.900 64.630 119.900 ;
        RECT 64.830 118.900 65.830 119.900 ;
        RECT 66.430 118.900 67.430 119.900 ;
        RECT 68.030 118.900 69.030 119.900 ;
        RECT 80.430 120.100 81.430 121.100 ;
        RECT 82.030 120.100 83.030 121.100 ;
        RECT 83.630 120.100 84.630 121.100 ;
        RECT 84.830 120.100 85.830 121.100 ;
        RECT 86.430 120.100 87.430 121.100 ;
        RECT 88.030 120.100 89.030 121.100 ;
        RECT 103.630 123.300 104.630 124.300 ;
        RECT 103.630 121.700 104.630 122.700 ;
        RECT 105.340 122.615 105.700 122.995 ;
        RECT 105.970 122.615 106.330 122.995 ;
        RECT 106.570 122.615 106.930 122.995 ;
        RECT 105.340 122.025 105.700 122.405 ;
        RECT 105.970 122.025 106.330 122.405 ;
        RECT 106.570 122.025 106.930 122.405 ;
        RECT 63.630 117.300 64.630 118.300 ;
        RECT 64.830 117.300 65.830 118.300 ;
        RECT 63.630 115.700 64.630 116.700 ;
        RECT 64.830 115.700 65.830 116.700 ;
        RECT 80.430 118.900 81.430 119.900 ;
        RECT 82.030 118.900 83.030 119.900 ;
        RECT 83.630 118.900 84.630 119.900 ;
        RECT 84.830 118.900 85.830 119.900 ;
        RECT 86.430 118.900 87.430 119.900 ;
        RECT 88.030 118.900 89.030 119.900 ;
        RECT 100.430 120.100 101.430 121.100 ;
        RECT 102.030 120.100 103.030 121.100 ;
        RECT 103.630 120.100 104.630 121.100 ;
        RECT 83.630 117.300 84.630 118.300 ;
        RECT 84.830 117.300 85.830 118.300 ;
        RECT 83.630 115.700 84.630 116.700 ;
        RECT 84.830 115.700 85.830 116.700 ;
        RECT 100.430 118.900 101.430 119.900 ;
        RECT 102.030 118.900 103.030 119.900 ;
        RECT 103.630 118.900 104.630 119.900 ;
        RECT 103.630 117.300 104.630 118.300 ;
        RECT 105.340 116.740 105.700 117.120 ;
        RECT 105.970 116.740 106.330 117.120 ;
        RECT 106.570 116.740 106.930 117.120 ;
        RECT 103.630 115.700 104.630 116.700 ;
        RECT 105.340 116.150 105.700 116.530 ;
        RECT 105.970 116.150 106.330 116.530 ;
        RECT 106.570 116.150 106.930 116.530 ;
        RECT 2.520 106.125 2.880 106.505 ;
        RECT 3.130 106.125 3.490 106.505 ;
        RECT 3.760 106.125 4.120 106.505 ;
        RECT 2.520 105.390 2.880 105.770 ;
        RECT 3.130 105.390 3.490 105.770 ;
        RECT 3.760 105.390 4.120 105.770 ;
        RECT 2.520 104.705 2.880 105.085 ;
        RECT 3.130 104.705 3.490 105.085 ;
        RECT 3.760 104.705 4.120 105.085 ;
        RECT 2.515 102.965 2.875 103.345 ;
        RECT 3.145 102.965 3.505 103.345 ;
        RECT 3.745 102.965 4.105 103.345 ;
        RECT 4.830 103.300 5.830 104.300 ;
        RECT 2.515 102.375 2.875 102.755 ;
        RECT 3.145 102.375 3.505 102.755 ;
        RECT 3.745 102.375 4.105 102.755 ;
        RECT 4.830 101.700 5.830 102.700 ;
        RECT 4.830 100.100 5.830 101.100 ;
        RECT 6.430 100.100 7.430 101.100 ;
        RECT 8.030 100.100 9.030 101.100 ;
        RECT 23.630 103.300 24.630 104.300 ;
        RECT 24.830 103.300 25.830 104.300 ;
        RECT 23.630 101.700 24.630 102.700 ;
        RECT 24.830 101.700 25.830 102.700 ;
        RECT 4.830 98.900 5.830 99.900 ;
        RECT 6.430 98.900 7.430 99.900 ;
        RECT 8.030 98.900 9.030 99.900 ;
        RECT 20.430 100.100 21.430 101.100 ;
        RECT 22.030 100.100 23.030 101.100 ;
        RECT 23.630 100.100 24.630 101.100 ;
        RECT 24.830 100.100 25.830 101.100 ;
        RECT 26.430 100.100 27.430 101.100 ;
        RECT 28.030 100.100 29.030 101.100 ;
        RECT 43.630 103.300 44.630 104.300 ;
        RECT 44.830 103.300 45.830 104.300 ;
        RECT 43.630 101.700 44.630 102.700 ;
        RECT 44.830 101.700 45.830 102.700 ;
        RECT 2.515 97.460 2.875 97.840 ;
        RECT 3.145 97.460 3.505 97.840 ;
        RECT 3.745 97.460 4.105 97.840 ;
        RECT 4.830 97.300 5.830 98.300 ;
        RECT 2.515 96.870 2.875 97.250 ;
        RECT 3.145 96.870 3.505 97.250 ;
        RECT 3.745 96.870 4.105 97.250 ;
        RECT 4.830 95.700 5.830 96.700 ;
        RECT 20.430 98.900 21.430 99.900 ;
        RECT 22.030 98.900 23.030 99.900 ;
        RECT 23.630 98.900 24.630 99.900 ;
        RECT 24.830 98.900 25.830 99.900 ;
        RECT 26.430 98.900 27.430 99.900 ;
        RECT 28.030 98.900 29.030 99.900 ;
        RECT 40.430 100.100 41.430 101.100 ;
        RECT 42.030 100.100 43.030 101.100 ;
        RECT 43.630 100.100 44.630 101.100 ;
        RECT 44.830 100.100 45.830 101.100 ;
        RECT 46.430 100.100 47.430 101.100 ;
        RECT 48.030 100.100 49.030 101.100 ;
        RECT 63.630 103.300 64.630 104.300 ;
        RECT 64.830 103.300 65.830 104.300 ;
        RECT 63.630 101.700 64.630 102.700 ;
        RECT 64.830 101.700 65.830 102.700 ;
        RECT 2.520 94.920 2.880 95.300 ;
        RECT 3.130 94.920 3.490 95.300 ;
        RECT 3.760 94.920 4.120 95.300 ;
        RECT 2.520 94.185 2.880 94.565 ;
        RECT 3.130 94.185 3.490 94.565 ;
        RECT 3.760 94.185 4.120 94.565 ;
        RECT 2.520 93.500 2.880 93.880 ;
        RECT 3.130 93.500 3.490 93.880 ;
        RECT 3.760 93.500 4.120 93.880 ;
        RECT 23.630 97.300 24.630 98.300 ;
        RECT 24.830 97.300 25.830 98.300 ;
        RECT 23.630 95.700 24.630 96.700 ;
        RECT 24.830 95.700 25.830 96.700 ;
        RECT 40.430 98.900 41.430 99.900 ;
        RECT 42.030 98.900 43.030 99.900 ;
        RECT 43.630 98.900 44.630 99.900 ;
        RECT 44.830 98.900 45.830 99.900 ;
        RECT 46.430 98.900 47.430 99.900 ;
        RECT 48.030 98.900 49.030 99.900 ;
        RECT 60.430 100.100 61.430 101.100 ;
        RECT 62.030 100.100 63.030 101.100 ;
        RECT 63.630 100.100 64.630 101.100 ;
        RECT 64.830 100.100 65.830 101.100 ;
        RECT 66.430 100.100 67.430 101.100 ;
        RECT 68.030 100.100 69.030 101.100 ;
        RECT 83.630 103.300 84.630 104.300 ;
        RECT 84.830 103.300 85.830 104.300 ;
        RECT 83.630 101.700 84.630 102.700 ;
        RECT 84.830 101.700 85.830 102.700 ;
        RECT 43.630 97.300 44.630 98.300 ;
        RECT 44.830 97.300 45.830 98.300 ;
        RECT 43.630 95.700 44.630 96.700 ;
        RECT 44.830 95.700 45.830 96.700 ;
        RECT 60.430 98.900 61.430 99.900 ;
        RECT 62.030 98.900 63.030 99.900 ;
        RECT 63.630 98.900 64.630 99.900 ;
        RECT 64.830 98.900 65.830 99.900 ;
        RECT 66.430 98.900 67.430 99.900 ;
        RECT 68.030 98.900 69.030 99.900 ;
        RECT 80.430 100.100 81.430 101.100 ;
        RECT 82.030 100.100 83.030 101.100 ;
        RECT 83.630 100.100 84.630 101.100 ;
        RECT 84.830 100.100 85.830 101.100 ;
        RECT 86.430 100.100 87.430 101.100 ;
        RECT 88.030 100.100 89.030 101.100 ;
        RECT 103.630 103.300 104.630 104.300 ;
        RECT 103.630 101.700 104.630 102.700 ;
        RECT 105.340 102.535 105.700 102.915 ;
        RECT 105.970 102.535 106.330 102.915 ;
        RECT 106.570 102.535 106.930 102.915 ;
        RECT 105.340 101.945 105.700 102.325 ;
        RECT 105.970 101.945 106.330 102.325 ;
        RECT 106.570 101.945 106.930 102.325 ;
        RECT 63.630 97.300 64.630 98.300 ;
        RECT 64.830 97.300 65.830 98.300 ;
        RECT 63.630 95.700 64.630 96.700 ;
        RECT 64.830 95.700 65.830 96.700 ;
        RECT 80.430 98.900 81.430 99.900 ;
        RECT 82.030 98.900 83.030 99.900 ;
        RECT 83.630 98.900 84.630 99.900 ;
        RECT 84.830 98.900 85.830 99.900 ;
        RECT 86.430 98.900 87.430 99.900 ;
        RECT 88.030 98.900 89.030 99.900 ;
        RECT 100.430 100.100 101.430 101.100 ;
        RECT 102.030 100.100 103.030 101.100 ;
        RECT 103.630 100.100 104.630 101.100 ;
        RECT 83.630 97.300 84.630 98.300 ;
        RECT 84.830 97.300 85.830 98.300 ;
        RECT 83.630 95.700 84.630 96.700 ;
        RECT 84.830 95.700 85.830 96.700 ;
        RECT 100.430 98.900 101.430 99.900 ;
        RECT 102.030 98.900 103.030 99.900 ;
        RECT 103.630 98.900 104.630 99.900 ;
        RECT 103.630 97.300 104.630 98.300 ;
        RECT 103.630 95.700 104.630 96.700 ;
        RECT 105.340 96.680 105.700 97.060 ;
        RECT 105.970 96.680 106.330 97.060 ;
        RECT 106.570 96.680 106.930 97.060 ;
        RECT 105.340 96.090 105.700 96.470 ;
        RECT 105.970 96.090 106.330 96.470 ;
        RECT 106.570 96.090 106.930 96.470 ;
        RECT 2.520 86.120 2.880 86.500 ;
        RECT 3.130 86.120 3.490 86.500 ;
        RECT 3.760 86.120 4.120 86.500 ;
        RECT 2.520 85.385 2.880 85.765 ;
        RECT 3.130 85.385 3.490 85.765 ;
        RECT 3.760 85.385 4.120 85.765 ;
        RECT 2.520 84.700 2.880 85.080 ;
        RECT 3.130 84.700 3.490 85.080 ;
        RECT 3.760 84.700 4.120 85.080 ;
        RECT 2.515 83.130 2.875 83.510 ;
        RECT 3.145 83.130 3.505 83.510 ;
        RECT 3.745 83.130 4.105 83.510 ;
        RECT 4.830 83.300 5.830 84.300 ;
        RECT 2.515 82.540 2.875 82.920 ;
        RECT 3.145 82.540 3.505 82.920 ;
        RECT 3.745 82.540 4.105 82.920 ;
        RECT 4.830 81.700 5.830 82.700 ;
        RECT 4.830 80.100 5.830 81.100 ;
        RECT 6.430 80.100 7.430 81.100 ;
        RECT 8.030 80.100 9.030 81.100 ;
        RECT 23.630 83.300 24.630 84.300 ;
        RECT 24.830 83.300 25.830 84.300 ;
        RECT 23.630 81.700 24.630 82.700 ;
        RECT 24.830 81.700 25.830 82.700 ;
        RECT 4.830 78.900 5.830 79.900 ;
        RECT 6.430 78.900 7.430 79.900 ;
        RECT 8.030 78.900 9.030 79.900 ;
        RECT 20.430 80.100 21.430 81.100 ;
        RECT 22.030 80.100 23.030 81.100 ;
        RECT 23.630 80.100 24.630 81.100 ;
        RECT 24.830 80.100 25.830 81.100 ;
        RECT 26.430 80.100 27.430 81.100 ;
        RECT 28.030 80.100 29.030 81.100 ;
        RECT 43.630 83.300 44.630 84.300 ;
        RECT 44.830 83.300 45.830 84.300 ;
        RECT 43.630 81.700 44.630 82.700 ;
        RECT 44.830 81.700 45.830 82.700 ;
        RECT 2.515 77.050 2.875 77.430 ;
        RECT 3.145 77.050 3.505 77.430 ;
        RECT 3.745 77.050 4.105 77.430 ;
        RECT 4.830 77.300 5.830 78.300 ;
        RECT 2.515 76.460 2.875 76.840 ;
        RECT 3.145 76.460 3.505 76.840 ;
        RECT 3.745 76.460 4.105 76.840 ;
        RECT 4.830 75.700 5.830 76.700 ;
        RECT 20.430 78.900 21.430 79.900 ;
        RECT 22.030 78.900 23.030 79.900 ;
        RECT 23.630 78.900 24.630 79.900 ;
        RECT 24.830 78.900 25.830 79.900 ;
        RECT 26.430 78.900 27.430 79.900 ;
        RECT 28.030 78.900 29.030 79.900 ;
        RECT 40.430 80.100 41.430 81.100 ;
        RECT 42.030 80.100 43.030 81.100 ;
        RECT 43.630 80.100 44.630 81.100 ;
        RECT 44.830 80.100 45.830 81.100 ;
        RECT 46.430 80.100 47.430 81.100 ;
        RECT 48.030 80.100 49.030 81.100 ;
        RECT 63.630 83.300 64.630 84.300 ;
        RECT 64.830 83.300 65.830 84.300 ;
        RECT 63.630 81.700 64.630 82.700 ;
        RECT 64.830 81.700 65.830 82.700 ;
        RECT 2.520 74.920 2.880 75.300 ;
        RECT 3.130 74.920 3.490 75.300 ;
        RECT 3.760 74.920 4.120 75.300 ;
        RECT 2.520 74.185 2.880 74.565 ;
        RECT 3.130 74.185 3.490 74.565 ;
        RECT 3.760 74.185 4.120 74.565 ;
        RECT 2.520 73.500 2.880 73.880 ;
        RECT 3.130 73.500 3.490 73.880 ;
        RECT 3.760 73.500 4.120 73.880 ;
        RECT 23.630 77.300 24.630 78.300 ;
        RECT 24.830 77.300 25.830 78.300 ;
        RECT 23.630 75.700 24.630 76.700 ;
        RECT 24.830 75.700 25.830 76.700 ;
        RECT 40.430 78.900 41.430 79.900 ;
        RECT 42.030 78.900 43.030 79.900 ;
        RECT 43.630 78.900 44.630 79.900 ;
        RECT 44.830 78.900 45.830 79.900 ;
        RECT 46.430 78.900 47.430 79.900 ;
        RECT 48.030 78.900 49.030 79.900 ;
        RECT 60.430 80.100 61.430 81.100 ;
        RECT 62.030 80.100 63.030 81.100 ;
        RECT 63.630 80.100 64.630 81.100 ;
        RECT 64.830 80.100 65.830 81.100 ;
        RECT 66.430 80.100 67.430 81.100 ;
        RECT 68.030 80.100 69.030 81.100 ;
        RECT 83.630 83.300 84.630 84.300 ;
        RECT 84.830 83.300 85.830 84.300 ;
        RECT 83.630 81.700 84.630 82.700 ;
        RECT 84.830 81.700 85.830 82.700 ;
        RECT 43.630 77.300 44.630 78.300 ;
        RECT 44.830 77.300 45.830 78.300 ;
        RECT 43.630 75.700 44.630 76.700 ;
        RECT 44.830 75.700 45.830 76.700 ;
        RECT 60.430 78.900 61.430 79.900 ;
        RECT 62.030 78.900 63.030 79.900 ;
        RECT 63.630 78.900 64.630 79.900 ;
        RECT 64.830 78.900 65.830 79.900 ;
        RECT 66.430 78.900 67.430 79.900 ;
        RECT 68.030 78.900 69.030 79.900 ;
        RECT 80.430 80.100 81.430 81.100 ;
        RECT 82.030 80.100 83.030 81.100 ;
        RECT 83.630 80.100 84.630 81.100 ;
        RECT 84.830 80.100 85.830 81.100 ;
        RECT 86.430 80.100 87.430 81.100 ;
        RECT 88.030 80.100 89.030 81.100 ;
        RECT 103.630 83.300 104.630 84.300 ;
        RECT 105.340 82.875 105.700 83.255 ;
        RECT 105.970 82.875 106.330 83.255 ;
        RECT 106.570 82.875 106.930 83.255 ;
        RECT 103.630 81.700 104.630 82.700 ;
        RECT 105.340 82.285 105.700 82.665 ;
        RECT 105.970 82.285 106.330 82.665 ;
        RECT 106.570 82.285 106.930 82.665 ;
        RECT 63.630 77.300 64.630 78.300 ;
        RECT 64.830 77.300 65.830 78.300 ;
        RECT 63.630 75.700 64.630 76.700 ;
        RECT 64.830 75.700 65.830 76.700 ;
        RECT 80.430 78.900 81.430 79.900 ;
        RECT 82.030 78.900 83.030 79.900 ;
        RECT 83.630 78.900 84.630 79.900 ;
        RECT 84.830 78.900 85.830 79.900 ;
        RECT 86.430 78.900 87.430 79.900 ;
        RECT 88.030 78.900 89.030 79.900 ;
        RECT 100.430 80.100 101.430 81.100 ;
        RECT 102.030 80.100 103.030 81.100 ;
        RECT 103.630 80.100 104.630 81.100 ;
        RECT 83.630 77.300 84.630 78.300 ;
        RECT 84.830 77.300 85.830 78.300 ;
        RECT 83.630 75.700 84.630 76.700 ;
        RECT 84.830 75.700 85.830 76.700 ;
        RECT 100.430 78.900 101.430 79.900 ;
        RECT 102.030 78.900 103.030 79.900 ;
        RECT 103.630 78.900 104.630 79.900 ;
        RECT 103.630 77.300 104.630 78.300 ;
        RECT 105.340 76.805 105.700 77.185 ;
        RECT 105.970 76.805 106.330 77.185 ;
        RECT 106.570 76.805 106.930 77.185 ;
        RECT 103.630 75.700 104.630 76.700 ;
        RECT 105.340 76.215 105.700 76.595 ;
        RECT 105.970 76.215 106.330 76.595 ;
        RECT 106.570 76.215 106.930 76.595 ;
        RECT 2.520 66.120 2.880 66.500 ;
        RECT 3.130 66.120 3.490 66.500 ;
        RECT 3.760 66.120 4.120 66.500 ;
        RECT 2.520 65.385 2.880 65.765 ;
        RECT 3.130 65.385 3.490 65.765 ;
        RECT 3.760 65.385 4.120 65.765 ;
        RECT 2.520 64.700 2.880 65.080 ;
        RECT 3.130 64.700 3.490 65.080 ;
        RECT 3.760 64.700 4.120 65.080 ;
        RECT 4.830 63.300 5.830 64.300 ;
        RECT 2.515 62.725 2.875 63.105 ;
        RECT 3.145 62.725 3.505 63.105 ;
        RECT 3.745 62.725 4.105 63.105 ;
        RECT 2.515 62.135 2.875 62.515 ;
        RECT 3.145 62.135 3.505 62.515 ;
        RECT 3.745 62.135 4.105 62.515 ;
        RECT 4.830 61.700 5.830 62.700 ;
        RECT 4.830 60.100 5.830 61.100 ;
        RECT 6.430 60.100 7.430 61.100 ;
        RECT 8.030 60.100 9.030 61.100 ;
        RECT 23.630 63.300 24.630 64.300 ;
        RECT 24.830 63.300 25.830 64.300 ;
        RECT 23.630 61.700 24.630 62.700 ;
        RECT 24.830 61.700 25.830 62.700 ;
        RECT 4.830 58.900 5.830 59.900 ;
        RECT 6.430 58.900 7.430 59.900 ;
        RECT 8.030 58.900 9.030 59.900 ;
        RECT 20.430 60.100 21.430 61.100 ;
        RECT 22.030 60.100 23.030 61.100 ;
        RECT 23.630 60.100 24.630 61.100 ;
        RECT 24.830 60.100 25.830 61.100 ;
        RECT 26.430 60.100 27.430 61.100 ;
        RECT 28.030 60.100 29.030 61.100 ;
        RECT 43.630 63.300 44.630 64.300 ;
        RECT 44.830 63.300 45.830 64.300 ;
        RECT 43.630 61.700 44.630 62.700 ;
        RECT 44.830 61.700 45.830 62.700 ;
        RECT 2.515 57.115 2.875 57.495 ;
        RECT 3.145 57.115 3.505 57.495 ;
        RECT 3.745 57.115 4.105 57.495 ;
        RECT 4.830 57.300 5.830 58.300 ;
        RECT 2.515 56.525 2.875 56.905 ;
        RECT 3.145 56.525 3.505 56.905 ;
        RECT 3.745 56.525 4.105 56.905 ;
        RECT 4.830 55.700 5.830 56.700 ;
        RECT 20.430 58.900 21.430 59.900 ;
        RECT 22.030 58.900 23.030 59.900 ;
        RECT 23.630 58.900 24.630 59.900 ;
        RECT 24.830 58.900 25.830 59.900 ;
        RECT 26.430 58.900 27.430 59.900 ;
        RECT 28.030 58.900 29.030 59.900 ;
        RECT 40.430 60.100 41.430 61.100 ;
        RECT 42.030 60.100 43.030 61.100 ;
        RECT 43.630 60.100 44.630 61.100 ;
        RECT 44.830 60.100 45.830 61.100 ;
        RECT 46.430 60.100 47.430 61.100 ;
        RECT 48.030 60.100 49.030 61.100 ;
        RECT 63.630 63.300 64.630 64.300 ;
        RECT 64.830 63.300 65.830 64.300 ;
        RECT 63.630 61.700 64.630 62.700 ;
        RECT 64.830 61.700 65.830 62.700 ;
        RECT 2.520 54.925 2.880 55.305 ;
        RECT 3.130 54.925 3.490 55.305 ;
        RECT 3.760 54.925 4.120 55.305 ;
        RECT 2.520 54.190 2.880 54.570 ;
        RECT 3.130 54.190 3.490 54.570 ;
        RECT 3.760 54.190 4.120 54.570 ;
        RECT 2.520 53.505 2.880 53.885 ;
        RECT 3.130 53.505 3.490 53.885 ;
        RECT 3.760 53.505 4.120 53.885 ;
        RECT 23.630 57.300 24.630 58.300 ;
        RECT 24.830 57.300 25.830 58.300 ;
        RECT 23.630 55.700 24.630 56.700 ;
        RECT 24.830 55.700 25.830 56.700 ;
        RECT 40.430 58.900 41.430 59.900 ;
        RECT 42.030 58.900 43.030 59.900 ;
        RECT 43.630 58.900 44.630 59.900 ;
        RECT 44.830 58.900 45.830 59.900 ;
        RECT 46.430 58.900 47.430 59.900 ;
        RECT 48.030 58.900 49.030 59.900 ;
        RECT 60.430 60.100 61.430 61.100 ;
        RECT 62.030 60.100 63.030 61.100 ;
        RECT 63.630 60.100 64.630 61.100 ;
        RECT 64.830 60.100 65.830 61.100 ;
        RECT 66.430 60.100 67.430 61.100 ;
        RECT 68.030 60.100 69.030 61.100 ;
        RECT 83.630 63.300 84.630 64.300 ;
        RECT 84.830 63.300 85.830 64.300 ;
        RECT 83.630 61.700 84.630 62.700 ;
        RECT 84.830 61.700 85.830 62.700 ;
        RECT 43.630 57.300 44.630 58.300 ;
        RECT 44.830 57.300 45.830 58.300 ;
        RECT 43.630 55.700 44.630 56.700 ;
        RECT 44.830 55.700 45.830 56.700 ;
        RECT 60.430 58.900 61.430 59.900 ;
        RECT 62.030 58.900 63.030 59.900 ;
        RECT 63.630 58.900 64.630 59.900 ;
        RECT 64.830 58.900 65.830 59.900 ;
        RECT 66.430 58.900 67.430 59.900 ;
        RECT 68.030 58.900 69.030 59.900 ;
        RECT 80.430 60.100 81.430 61.100 ;
        RECT 82.030 60.100 83.030 61.100 ;
        RECT 83.630 60.100 84.630 61.100 ;
        RECT 84.830 60.100 85.830 61.100 ;
        RECT 86.430 60.100 87.430 61.100 ;
        RECT 88.030 60.100 89.030 61.100 ;
        RECT 103.630 63.300 104.630 64.300 ;
        RECT 103.630 61.700 104.630 62.700 ;
        RECT 105.340 62.590 105.700 62.970 ;
        RECT 105.970 62.590 106.330 62.970 ;
        RECT 106.570 62.590 106.930 62.970 ;
        RECT 105.340 62.000 105.700 62.380 ;
        RECT 105.970 62.000 106.330 62.380 ;
        RECT 106.570 62.000 106.930 62.380 ;
        RECT 63.630 57.300 64.630 58.300 ;
        RECT 64.830 57.300 65.830 58.300 ;
        RECT 63.630 55.700 64.630 56.700 ;
        RECT 64.830 55.700 65.830 56.700 ;
        RECT 80.430 58.900 81.430 59.900 ;
        RECT 82.030 58.900 83.030 59.900 ;
        RECT 83.630 58.900 84.630 59.900 ;
        RECT 84.830 58.900 85.830 59.900 ;
        RECT 86.430 58.900 87.430 59.900 ;
        RECT 88.030 58.900 89.030 59.900 ;
        RECT 100.430 60.100 101.430 61.100 ;
        RECT 102.030 60.100 103.030 61.100 ;
        RECT 103.630 60.100 104.630 61.100 ;
        RECT 83.630 57.300 84.630 58.300 ;
        RECT 84.830 57.300 85.830 58.300 ;
        RECT 83.630 55.700 84.630 56.700 ;
        RECT 84.830 55.700 85.830 56.700 ;
        RECT 100.430 58.900 101.430 59.900 ;
        RECT 102.030 58.900 103.030 59.900 ;
        RECT 103.630 58.900 104.630 59.900 ;
        RECT 103.630 57.300 104.630 58.300 ;
        RECT 105.340 56.805 105.700 57.185 ;
        RECT 105.970 56.805 106.330 57.185 ;
        RECT 106.570 56.805 106.930 57.185 ;
        RECT 103.630 55.700 104.630 56.700 ;
        RECT 105.340 56.215 105.700 56.595 ;
        RECT 105.970 56.215 106.330 56.595 ;
        RECT 106.570 56.215 106.930 56.595 ;
        RECT 2.520 46.115 2.880 46.495 ;
        RECT 3.130 46.115 3.490 46.495 ;
        RECT 3.760 46.115 4.120 46.495 ;
        RECT 2.520 45.380 2.880 45.760 ;
        RECT 3.130 45.380 3.490 45.760 ;
        RECT 3.760 45.380 4.120 45.760 ;
        RECT 2.520 44.695 2.880 45.075 ;
        RECT 3.130 44.695 3.490 45.075 ;
        RECT 3.760 44.695 4.120 45.075 ;
        RECT 4.830 43.300 5.830 44.300 ;
        RECT 2.515 42.815 2.875 43.195 ;
        RECT 3.145 42.815 3.505 43.195 ;
        RECT 3.745 42.815 4.105 43.195 ;
        RECT 2.515 42.225 2.875 42.605 ;
        RECT 3.145 42.225 3.505 42.605 ;
        RECT 3.745 42.225 4.105 42.605 ;
        RECT 4.830 41.700 5.830 42.700 ;
        RECT 4.830 40.100 5.830 41.100 ;
        RECT 6.430 40.100 7.430 41.100 ;
        RECT 8.030 40.100 9.030 41.100 ;
        RECT 23.630 43.300 24.630 44.300 ;
        RECT 24.830 43.300 25.830 44.300 ;
        RECT 23.630 41.700 24.630 42.700 ;
        RECT 24.830 41.700 25.830 42.700 ;
        RECT 4.830 38.900 5.830 39.900 ;
        RECT 6.430 38.900 7.430 39.900 ;
        RECT 8.030 38.900 9.030 39.900 ;
        RECT 20.430 40.100 21.430 41.100 ;
        RECT 22.030 40.100 23.030 41.100 ;
        RECT 23.630 40.100 24.630 41.100 ;
        RECT 24.830 40.100 25.830 41.100 ;
        RECT 26.430 40.100 27.430 41.100 ;
        RECT 28.030 40.100 29.030 41.100 ;
        RECT 43.630 43.300 44.630 44.300 ;
        RECT 44.830 43.300 45.830 44.300 ;
        RECT 43.630 41.700 44.630 42.700 ;
        RECT 44.830 41.700 45.830 42.700 ;
        RECT 2.515 37.260 2.875 37.640 ;
        RECT 3.145 37.260 3.505 37.640 ;
        RECT 3.745 37.260 4.105 37.640 ;
        RECT 4.830 37.300 5.830 38.300 ;
        RECT 2.515 36.670 2.875 37.050 ;
        RECT 3.145 36.670 3.505 37.050 ;
        RECT 3.745 36.670 4.105 37.050 ;
        RECT 4.830 35.700 5.830 36.700 ;
        RECT 20.430 38.900 21.430 39.900 ;
        RECT 22.030 38.900 23.030 39.900 ;
        RECT 23.630 38.900 24.630 39.900 ;
        RECT 24.830 38.900 25.830 39.900 ;
        RECT 26.430 38.900 27.430 39.900 ;
        RECT 28.030 38.900 29.030 39.900 ;
        RECT 40.430 40.100 41.430 41.100 ;
        RECT 42.030 40.100 43.030 41.100 ;
        RECT 43.630 40.100 44.630 41.100 ;
        RECT 44.830 40.100 45.830 41.100 ;
        RECT 46.430 40.100 47.430 41.100 ;
        RECT 48.030 40.100 49.030 41.100 ;
        RECT 63.630 43.300 64.630 44.300 ;
        RECT 64.830 43.300 65.830 44.300 ;
        RECT 63.630 41.700 64.630 42.700 ;
        RECT 64.830 41.700 65.830 42.700 ;
        RECT 2.520 34.925 2.880 35.305 ;
        RECT 3.130 34.925 3.490 35.305 ;
        RECT 3.760 34.925 4.120 35.305 ;
        RECT 2.520 34.190 2.880 34.570 ;
        RECT 3.130 34.190 3.490 34.570 ;
        RECT 3.760 34.190 4.120 34.570 ;
        RECT 2.520 33.505 2.880 33.885 ;
        RECT 3.130 33.505 3.490 33.885 ;
        RECT 3.760 33.505 4.120 33.885 ;
        RECT 23.630 37.300 24.630 38.300 ;
        RECT 24.830 37.300 25.830 38.300 ;
        RECT 23.630 35.700 24.630 36.700 ;
        RECT 24.830 35.700 25.830 36.700 ;
        RECT 40.430 38.900 41.430 39.900 ;
        RECT 42.030 38.900 43.030 39.900 ;
        RECT 43.630 38.900 44.630 39.900 ;
        RECT 44.830 38.900 45.830 39.900 ;
        RECT 46.430 38.900 47.430 39.900 ;
        RECT 48.030 38.900 49.030 39.900 ;
        RECT 60.430 40.100 61.430 41.100 ;
        RECT 62.030 40.100 63.030 41.100 ;
        RECT 63.630 40.100 64.630 41.100 ;
        RECT 64.830 40.100 65.830 41.100 ;
        RECT 66.430 40.100 67.430 41.100 ;
        RECT 68.030 40.100 69.030 41.100 ;
        RECT 83.630 43.300 84.630 44.300 ;
        RECT 84.830 43.300 85.830 44.300 ;
        RECT 83.630 41.700 84.630 42.700 ;
        RECT 84.830 41.700 85.830 42.700 ;
        RECT 43.630 37.300 44.630 38.300 ;
        RECT 44.830 37.300 45.830 38.300 ;
        RECT 43.630 35.700 44.630 36.700 ;
        RECT 44.830 35.700 45.830 36.700 ;
        RECT 60.430 38.900 61.430 39.900 ;
        RECT 62.030 38.900 63.030 39.900 ;
        RECT 63.630 38.900 64.630 39.900 ;
        RECT 64.830 38.900 65.830 39.900 ;
        RECT 66.430 38.900 67.430 39.900 ;
        RECT 68.030 38.900 69.030 39.900 ;
        RECT 80.430 40.100 81.430 41.100 ;
        RECT 82.030 40.100 83.030 41.100 ;
        RECT 83.630 40.100 84.630 41.100 ;
        RECT 84.830 40.100 85.830 41.100 ;
        RECT 86.430 40.100 87.430 41.100 ;
        RECT 88.030 40.100 89.030 41.100 ;
        RECT 103.630 43.300 104.630 44.300 ;
        RECT 103.630 41.700 104.630 42.700 ;
        RECT 105.340 42.590 105.700 42.970 ;
        RECT 105.970 42.590 106.330 42.970 ;
        RECT 106.570 42.590 106.930 42.970 ;
        RECT 105.340 42.000 105.700 42.380 ;
        RECT 105.970 42.000 106.330 42.380 ;
        RECT 106.570 42.000 106.930 42.380 ;
        RECT 63.630 37.300 64.630 38.300 ;
        RECT 64.830 37.300 65.830 38.300 ;
        RECT 63.630 35.700 64.630 36.700 ;
        RECT 64.830 35.700 65.830 36.700 ;
        RECT 80.430 38.900 81.430 39.900 ;
        RECT 82.030 38.900 83.030 39.900 ;
        RECT 83.630 38.900 84.630 39.900 ;
        RECT 84.830 38.900 85.830 39.900 ;
        RECT 86.430 38.900 87.430 39.900 ;
        RECT 88.030 38.900 89.030 39.900 ;
        RECT 100.430 40.100 101.430 41.100 ;
        RECT 102.030 40.100 103.030 41.100 ;
        RECT 103.630 40.100 104.630 41.100 ;
        RECT 83.630 37.300 84.630 38.300 ;
        RECT 84.830 37.300 85.830 38.300 ;
        RECT 83.630 35.700 84.630 36.700 ;
        RECT 84.830 35.700 85.830 36.700 ;
        RECT 100.430 38.900 101.430 39.900 ;
        RECT 102.030 38.900 103.030 39.900 ;
        RECT 103.630 38.900 104.630 39.900 ;
        RECT 103.630 37.300 104.630 38.300 ;
        RECT 105.340 36.805 105.700 37.185 ;
        RECT 105.970 36.805 106.330 37.185 ;
        RECT 106.570 36.805 106.930 37.185 ;
        RECT 103.630 35.700 104.630 36.700 ;
        RECT 105.340 36.215 105.700 36.595 ;
        RECT 105.970 36.215 106.330 36.595 ;
        RECT 106.570 36.215 106.930 36.595 ;
        RECT 2.520 26.120 2.880 26.500 ;
        RECT 3.130 26.120 3.490 26.500 ;
        RECT 3.760 26.120 4.120 26.500 ;
        RECT 2.520 25.385 2.880 25.765 ;
        RECT 3.130 25.385 3.490 25.765 ;
        RECT 3.760 25.385 4.120 25.765 ;
        RECT 2.520 24.700 2.880 25.080 ;
        RECT 3.130 24.700 3.490 25.080 ;
        RECT 3.760 24.700 4.120 25.080 ;
        RECT 2.515 23.145 2.875 23.525 ;
        RECT 3.145 23.145 3.505 23.525 ;
        RECT 3.745 23.145 4.105 23.525 ;
        RECT 4.830 23.300 5.830 24.300 ;
        RECT 2.515 22.555 2.875 22.935 ;
        RECT 3.145 22.555 3.505 22.935 ;
        RECT 3.745 22.555 4.105 22.935 ;
        RECT 4.830 21.700 5.830 22.700 ;
        RECT 4.830 20.100 5.830 21.100 ;
        RECT 6.430 20.100 7.430 21.100 ;
        RECT 8.030 20.100 9.030 21.100 ;
        RECT 23.630 23.300 24.630 24.300 ;
        RECT 24.830 23.300 25.830 24.300 ;
        RECT 23.630 21.700 24.630 22.700 ;
        RECT 24.830 21.700 25.830 22.700 ;
        RECT 4.830 18.900 5.830 19.900 ;
        RECT 6.430 18.900 7.430 19.900 ;
        RECT 8.030 18.900 9.030 19.900 ;
        RECT 20.430 20.100 21.430 21.100 ;
        RECT 22.030 20.100 23.030 21.100 ;
        RECT 23.630 20.100 24.630 21.100 ;
        RECT 24.830 20.100 25.830 21.100 ;
        RECT 26.430 20.100 27.430 21.100 ;
        RECT 28.030 20.100 29.030 21.100 ;
        RECT 43.630 23.300 44.630 24.300 ;
        RECT 44.830 23.300 45.830 24.300 ;
        RECT 43.630 21.700 44.630 22.700 ;
        RECT 44.830 21.700 45.830 22.700 ;
        RECT 2.515 17.260 2.875 17.640 ;
        RECT 3.145 17.260 3.505 17.640 ;
        RECT 3.745 17.260 4.105 17.640 ;
        RECT 4.830 17.300 5.830 18.300 ;
        RECT 2.515 16.670 2.875 17.050 ;
        RECT 3.145 16.670 3.505 17.050 ;
        RECT 3.745 16.670 4.105 17.050 ;
        RECT 4.830 15.700 5.830 16.700 ;
        RECT 20.430 18.900 21.430 19.900 ;
        RECT 22.030 18.900 23.030 19.900 ;
        RECT 23.630 18.900 24.630 19.900 ;
        RECT 24.830 18.900 25.830 19.900 ;
        RECT 26.430 18.900 27.430 19.900 ;
        RECT 28.030 18.900 29.030 19.900 ;
        RECT 40.430 20.100 41.430 21.100 ;
        RECT 42.030 20.100 43.030 21.100 ;
        RECT 43.630 20.100 44.630 21.100 ;
        RECT 44.830 20.100 45.830 21.100 ;
        RECT 46.430 20.100 47.430 21.100 ;
        RECT 48.030 20.100 49.030 21.100 ;
        RECT 63.630 23.300 64.630 24.300 ;
        RECT 64.830 23.300 65.830 24.300 ;
        RECT 63.630 21.700 64.630 22.700 ;
        RECT 64.830 21.700 65.830 22.700 ;
        RECT 2.520 14.925 2.880 15.305 ;
        RECT 3.130 14.925 3.490 15.305 ;
        RECT 3.760 14.925 4.120 15.305 ;
        RECT 2.520 14.190 2.880 14.570 ;
        RECT 3.130 14.190 3.490 14.570 ;
        RECT 3.760 14.190 4.120 14.570 ;
        RECT 2.520 13.505 2.880 13.885 ;
        RECT 3.130 13.505 3.490 13.885 ;
        RECT 3.760 13.505 4.120 13.885 ;
        RECT 23.630 17.300 24.630 18.300 ;
        RECT 24.830 17.300 25.830 18.300 ;
        RECT 23.630 15.700 24.630 16.700 ;
        RECT 24.830 15.700 25.830 16.700 ;
        RECT 40.430 18.900 41.430 19.900 ;
        RECT 42.030 18.900 43.030 19.900 ;
        RECT 43.630 18.900 44.630 19.900 ;
        RECT 44.830 18.900 45.830 19.900 ;
        RECT 46.430 18.900 47.430 19.900 ;
        RECT 48.030 18.900 49.030 19.900 ;
        RECT 60.430 20.100 61.430 21.100 ;
        RECT 62.030 20.100 63.030 21.100 ;
        RECT 63.630 20.100 64.630 21.100 ;
        RECT 64.830 20.100 65.830 21.100 ;
        RECT 66.430 20.100 67.430 21.100 ;
        RECT 68.030 20.100 69.030 21.100 ;
        RECT 83.630 23.300 84.630 24.300 ;
        RECT 84.830 23.300 85.830 24.300 ;
        RECT 83.630 21.700 84.630 22.700 ;
        RECT 84.830 21.700 85.830 22.700 ;
        RECT 43.630 17.300 44.630 18.300 ;
        RECT 44.830 17.300 45.830 18.300 ;
        RECT 43.630 15.700 44.630 16.700 ;
        RECT 44.830 15.700 45.830 16.700 ;
        RECT 60.430 18.900 61.430 19.900 ;
        RECT 62.030 18.900 63.030 19.900 ;
        RECT 63.630 18.900 64.630 19.900 ;
        RECT 64.830 18.900 65.830 19.900 ;
        RECT 66.430 18.900 67.430 19.900 ;
        RECT 68.030 18.900 69.030 19.900 ;
        RECT 80.430 20.100 81.430 21.100 ;
        RECT 82.030 20.100 83.030 21.100 ;
        RECT 83.630 20.100 84.630 21.100 ;
        RECT 84.830 20.100 85.830 21.100 ;
        RECT 86.430 20.100 87.430 21.100 ;
        RECT 88.030 20.100 89.030 21.100 ;
        RECT 103.630 23.300 104.630 24.300 ;
        RECT 103.630 21.700 104.630 22.700 ;
        RECT 105.340 22.590 105.700 22.970 ;
        RECT 105.970 22.590 106.330 22.970 ;
        RECT 106.570 22.590 106.930 22.970 ;
        RECT 105.340 22.000 105.700 22.380 ;
        RECT 105.970 22.000 106.330 22.380 ;
        RECT 106.570 22.000 106.930 22.380 ;
        RECT 63.630 17.300 64.630 18.300 ;
        RECT 64.830 17.300 65.830 18.300 ;
        RECT 63.630 15.700 64.630 16.700 ;
        RECT 64.830 15.700 65.830 16.700 ;
        RECT 80.430 18.900 81.430 19.900 ;
        RECT 82.030 18.900 83.030 19.900 ;
        RECT 83.630 18.900 84.630 19.900 ;
        RECT 84.830 18.900 85.830 19.900 ;
        RECT 86.430 18.900 87.430 19.900 ;
        RECT 88.030 18.900 89.030 19.900 ;
        RECT 100.430 20.100 101.430 21.100 ;
        RECT 102.030 20.100 103.030 21.100 ;
        RECT 103.630 20.100 104.630 21.100 ;
        RECT 83.630 17.300 84.630 18.300 ;
        RECT 84.830 17.300 85.830 18.300 ;
        RECT 83.630 15.700 84.630 16.700 ;
        RECT 84.830 15.700 85.830 16.700 ;
        RECT 100.430 18.900 101.430 19.900 ;
        RECT 102.030 18.900 103.030 19.900 ;
        RECT 103.630 18.900 104.630 19.900 ;
        RECT 103.630 17.300 104.630 18.300 ;
        RECT 105.340 16.805 105.700 17.185 ;
        RECT 105.970 16.805 106.330 17.185 ;
        RECT 106.570 16.805 106.930 17.185 ;
        RECT 103.630 15.700 104.630 16.700 ;
        RECT 105.340 16.215 105.700 16.595 ;
        RECT 105.970 16.215 106.330 16.595 ;
        RECT 106.570 16.215 106.930 16.595 ;
        RECT 2.520 6.120 2.880 6.500 ;
        RECT 3.130 6.120 3.490 6.500 ;
        RECT 3.760 6.120 4.120 6.500 ;
        RECT 2.520 5.385 2.880 5.765 ;
        RECT 3.130 5.385 3.490 5.765 ;
        RECT 3.760 5.385 4.120 5.765 ;
        RECT 2.520 4.700 2.880 5.080 ;
        RECT 3.130 4.700 3.490 5.080 ;
        RECT 3.760 4.700 4.120 5.080 ;
        RECT 2.515 3.145 2.875 3.525 ;
        RECT 3.145 3.145 3.505 3.525 ;
        RECT 3.745 3.145 4.105 3.525 ;
        RECT 4.830 3.300 5.830 4.300 ;
        RECT 2.515 2.555 2.875 2.935 ;
        RECT 3.145 2.555 3.505 2.935 ;
        RECT 3.745 2.555 4.105 2.935 ;
        RECT 4.830 1.700 5.830 2.700 ;
        RECT 4.830 0.100 5.830 1.100 ;
        RECT 6.430 0.100 7.430 1.100 ;
        RECT 8.030 0.100 9.030 1.100 ;
        RECT 23.630 3.300 24.630 4.300 ;
        RECT 24.830 3.300 25.830 4.300 ;
        RECT 23.630 1.700 24.630 2.700 ;
        RECT 24.830 1.700 25.830 2.700 ;
        RECT 20.430 0.100 21.430 1.100 ;
        RECT 22.030 0.100 23.030 1.100 ;
        RECT 23.630 0.100 24.630 1.100 ;
        RECT 24.830 0.100 25.830 1.100 ;
        RECT 26.430 0.100 27.430 1.100 ;
        RECT 28.030 0.100 29.030 1.100 ;
        RECT 43.630 3.300 44.630 4.300 ;
        RECT 44.830 3.300 45.830 4.300 ;
        RECT 43.630 1.700 44.630 2.700 ;
        RECT 44.830 1.700 45.830 2.700 ;
        RECT 40.430 0.100 41.430 1.100 ;
        RECT 42.030 0.100 43.030 1.100 ;
        RECT 43.630 0.100 44.630 1.100 ;
        RECT 44.830 0.100 45.830 1.100 ;
        RECT 46.430 0.100 47.430 1.100 ;
        RECT 48.030 0.100 49.030 1.100 ;
        RECT 63.630 3.300 64.630 4.300 ;
        RECT 64.830 3.300 65.830 4.300 ;
        RECT 63.630 1.700 64.630 2.700 ;
        RECT 64.830 1.700 65.830 2.700 ;
        RECT 60.430 0.100 61.430 1.100 ;
        RECT 62.030 0.100 63.030 1.100 ;
        RECT 63.630 0.100 64.630 1.100 ;
        RECT 64.830 0.100 65.830 1.100 ;
        RECT 66.430 0.100 67.430 1.100 ;
        RECT 68.030 0.100 69.030 1.100 ;
        RECT 83.630 3.300 84.630 4.300 ;
        RECT 84.830 3.300 85.830 4.300 ;
        RECT 83.630 1.700 84.630 2.700 ;
        RECT 84.830 1.700 85.830 2.700 ;
        RECT 80.430 0.100 81.430 1.100 ;
        RECT 82.030 0.100 83.030 1.100 ;
        RECT 83.630 0.100 84.630 1.100 ;
        RECT 84.830 0.100 85.830 1.100 ;
        RECT 86.430 0.100 87.430 1.100 ;
        RECT 88.030 0.100 89.030 1.100 ;
        RECT 103.630 3.300 104.630 4.300 ;
        RECT 103.630 1.700 104.630 2.700 ;
        RECT 105.340 2.590 105.700 2.970 ;
        RECT 105.970 2.590 106.330 2.970 ;
        RECT 106.570 2.590 106.930 2.970 ;
        RECT 105.340 2.000 105.700 2.380 ;
        RECT 105.970 2.000 106.330 2.380 ;
        RECT 106.570 2.000 106.930 2.380 ;
        RECT 100.430 0.100 101.430 1.100 ;
        RECT 102.030 0.100 103.030 1.100 ;
        RECT 103.630 0.100 104.630 1.100 ;
      LAYER met2 ;
        RECT 4.730 378.800 9.130 380.000 ;
        RECT 20.330 378.800 29.130 380.000 ;
        RECT 40.330 378.800 49.130 380.000 ;
        RECT 60.330 378.800 69.130 380.000 ;
        RECT 80.330 378.800 89.130 380.000 ;
        RECT 100.330 378.800 104.730 380.000 ;
        RECT 4.730 377.850 5.940 378.800 ;
        RECT 4.730 377.700 9.880 377.850 ;
        RECT 2.315 376.110 4.320 377.385 ;
        RECT 4.730 377.250 6.330 377.700 ;
        RECT 4.730 377.100 9.880 377.250 ;
        RECT 4.730 376.650 6.330 377.100 ;
        RECT 4.730 376.500 9.880 376.650 ;
        RECT 4.730 376.050 6.330 376.500 ;
        RECT 4.730 375.900 9.880 376.050 ;
        RECT 4.730 375.600 6.330 375.900 ;
        RECT 2.315 373.250 4.315 375.545 ;
        RECT 5.930 375.450 6.330 375.600 ;
        RECT 5.930 375.300 9.880 375.450 ;
        RECT 5.930 374.850 6.330 375.300 ;
        RECT 5.930 374.700 9.880 374.850 ;
        RECT 5.930 374.250 6.330 374.700 ;
        RECT 5.930 374.100 9.880 374.250 ;
        RECT 5.930 373.650 6.330 374.100 ;
        RECT 5.930 373.500 9.880 373.650 ;
        RECT 5.930 373.050 6.330 373.500 ;
        RECT 5.930 372.900 9.880 373.050 ;
        RECT 5.930 372.450 6.330 372.900 ;
        RECT 5.930 372.300 9.880 372.450 ;
        RECT 5.930 371.850 6.330 372.300 ;
        RECT 5.930 371.700 9.880 371.850 ;
        RECT 5.930 371.250 6.330 371.700 ;
        RECT 5.930 371.100 9.880 371.250 ;
        RECT 5.930 370.650 6.330 371.100 ;
        RECT 5.930 370.500 9.880 370.650 ;
        RECT 5.930 370.200 6.330 370.500 ;
        RECT 10.480 370.200 10.630 378.400 ;
        RECT 11.080 370.200 11.230 378.400 ;
        RECT 11.680 370.200 11.830 378.400 ;
        RECT 12.280 370.200 12.430 378.400 ;
        RECT 12.880 370.200 13.030 378.400 ;
        RECT 13.480 370.200 13.630 378.400 ;
        RECT 14.080 370.200 14.230 378.400 ;
        RECT 5.930 369.800 14.230 370.200 ;
        RECT 5.930 369.500 6.330 369.800 ;
        RECT 5.930 369.350 9.880 369.500 ;
        RECT 5.930 368.900 6.330 369.350 ;
        RECT 5.930 368.750 9.880 368.900 ;
        RECT 5.930 368.300 6.330 368.750 ;
        RECT 5.930 368.150 9.880 368.300 ;
        RECT 5.930 367.700 6.330 368.150 ;
        RECT 5.930 367.550 9.880 367.700 ;
        RECT 5.930 367.100 6.330 367.550 ;
        RECT 5.930 366.950 9.880 367.100 ;
        RECT 2.315 364.450 4.315 366.745 ;
        RECT 5.930 366.500 6.330 366.950 ;
        RECT 5.930 366.350 9.880 366.500 ;
        RECT 5.930 365.900 6.330 366.350 ;
        RECT 5.930 365.750 9.880 365.900 ;
        RECT 5.930 365.300 6.330 365.750 ;
        RECT 5.930 365.150 9.880 365.300 ;
        RECT 5.930 364.700 6.330 365.150 ;
        RECT 5.930 364.550 9.880 364.700 ;
        RECT 5.930 364.400 6.330 364.550 ;
        RECT 4.730 364.100 6.330 364.400 ;
        RECT 2.315 362.745 4.320 364.020 ;
        RECT 4.730 363.950 9.880 364.100 ;
        RECT 4.730 363.500 6.330 363.950 ;
        RECT 4.730 363.350 9.880 363.500 ;
        RECT 4.730 362.900 6.330 363.350 ;
        RECT 4.730 362.750 9.880 362.900 ;
        RECT 4.730 362.300 6.330 362.750 ;
        RECT 4.730 362.150 9.880 362.300 ;
        RECT 4.730 361.200 5.930 362.150 ;
        RECT 10.480 361.600 10.630 369.800 ;
        RECT 11.080 361.600 11.230 369.800 ;
        RECT 11.680 361.600 11.830 369.800 ;
        RECT 12.280 361.600 12.430 369.800 ;
        RECT 12.880 361.600 13.030 369.800 ;
        RECT 13.480 361.600 13.630 369.800 ;
        RECT 14.080 361.600 14.230 369.800 ;
        RECT 15.230 370.200 15.380 378.400 ;
        RECT 15.830 370.200 15.980 378.400 ;
        RECT 16.430 370.200 16.580 378.400 ;
        RECT 17.030 370.200 17.180 378.400 ;
        RECT 17.630 370.200 17.780 378.400 ;
        RECT 18.230 370.200 18.380 378.400 ;
        RECT 18.830 370.200 18.980 378.400 ;
        RECT 23.530 377.850 25.940 378.800 ;
        RECT 19.580 377.700 29.880 377.850 ;
        RECT 23.130 377.250 26.330 377.700 ;
        RECT 19.580 377.100 29.880 377.250 ;
        RECT 23.130 376.650 26.330 377.100 ;
        RECT 19.580 376.500 29.880 376.650 ;
        RECT 23.130 376.050 26.330 376.500 ;
        RECT 19.580 375.900 29.880 376.050 ;
        RECT 23.130 375.600 26.330 375.900 ;
        RECT 23.130 375.450 23.530 375.600 ;
        RECT 19.580 375.300 23.530 375.450 ;
        RECT 23.130 374.850 23.530 375.300 ;
        RECT 19.580 374.700 23.530 374.850 ;
        RECT 23.130 374.250 23.530 374.700 ;
        RECT 19.580 374.100 23.530 374.250 ;
        RECT 23.130 373.650 23.530 374.100 ;
        RECT 19.580 373.500 23.530 373.650 ;
        RECT 23.130 373.050 23.530 373.500 ;
        RECT 19.580 372.900 23.530 373.050 ;
        RECT 23.130 372.450 23.530 372.900 ;
        RECT 19.580 372.300 23.530 372.450 ;
        RECT 23.130 371.850 23.530 372.300 ;
        RECT 19.580 371.700 23.530 371.850 ;
        RECT 23.130 371.250 23.530 371.700 ;
        RECT 19.580 371.100 23.530 371.250 ;
        RECT 23.130 370.650 23.530 371.100 ;
        RECT 19.580 370.500 23.530 370.650 ;
        RECT 23.130 370.200 23.530 370.500 ;
        RECT 15.230 369.800 23.530 370.200 ;
        RECT 15.230 361.600 15.380 369.800 ;
        RECT 15.830 361.600 15.980 369.800 ;
        RECT 16.430 361.600 16.580 369.800 ;
        RECT 17.030 361.600 17.180 369.800 ;
        RECT 17.630 361.600 17.780 369.800 ;
        RECT 18.230 361.600 18.380 369.800 ;
        RECT 18.830 361.600 18.980 369.800 ;
        RECT 23.130 369.500 23.530 369.800 ;
        RECT 19.580 369.350 23.530 369.500 ;
        RECT 23.130 368.900 23.530 369.350 ;
        RECT 19.580 368.750 23.530 368.900 ;
        RECT 23.130 368.300 23.530 368.750 ;
        RECT 19.580 368.150 23.530 368.300 ;
        RECT 23.130 367.700 23.530 368.150 ;
        RECT 19.580 367.550 23.530 367.700 ;
        RECT 23.130 367.100 23.530 367.550 ;
        RECT 19.580 366.950 23.530 367.100 ;
        RECT 23.130 366.500 23.530 366.950 ;
        RECT 19.580 366.350 23.530 366.500 ;
        RECT 23.130 365.900 23.530 366.350 ;
        RECT 19.580 365.750 23.530 365.900 ;
        RECT 23.130 365.300 23.530 365.750 ;
        RECT 19.580 365.150 23.530 365.300 ;
        RECT 23.130 364.700 23.530 365.150 ;
        RECT 19.580 364.550 23.530 364.700 ;
        RECT 23.130 364.400 23.530 364.550 ;
        RECT 25.930 375.450 26.330 375.600 ;
        RECT 25.930 375.300 29.880 375.450 ;
        RECT 25.930 374.850 26.330 375.300 ;
        RECT 25.930 374.700 29.880 374.850 ;
        RECT 25.930 374.250 26.330 374.700 ;
        RECT 25.930 374.100 29.880 374.250 ;
        RECT 25.930 373.650 26.330 374.100 ;
        RECT 25.930 373.500 29.880 373.650 ;
        RECT 25.930 373.050 26.330 373.500 ;
        RECT 25.930 372.900 29.880 373.050 ;
        RECT 25.930 372.450 26.330 372.900 ;
        RECT 25.930 372.300 29.880 372.450 ;
        RECT 25.930 371.850 26.330 372.300 ;
        RECT 25.930 371.700 29.880 371.850 ;
        RECT 25.930 371.250 26.330 371.700 ;
        RECT 25.930 371.100 29.880 371.250 ;
        RECT 25.930 370.650 26.330 371.100 ;
        RECT 25.930 370.500 29.880 370.650 ;
        RECT 25.930 370.200 26.330 370.500 ;
        RECT 30.480 370.200 30.630 378.400 ;
        RECT 31.080 370.200 31.230 378.400 ;
        RECT 31.680 370.200 31.830 378.400 ;
        RECT 32.280 370.200 32.430 378.400 ;
        RECT 32.880 370.200 33.030 378.400 ;
        RECT 33.480 370.200 33.630 378.400 ;
        RECT 34.080 370.200 34.230 378.400 ;
        RECT 25.930 369.800 34.230 370.200 ;
        RECT 25.930 369.500 26.330 369.800 ;
        RECT 25.930 369.350 29.880 369.500 ;
        RECT 25.930 368.900 26.330 369.350 ;
        RECT 25.930 368.750 29.880 368.900 ;
        RECT 25.930 368.300 26.330 368.750 ;
        RECT 25.930 368.150 29.880 368.300 ;
        RECT 25.930 367.700 26.330 368.150 ;
        RECT 25.930 367.550 29.880 367.700 ;
        RECT 25.930 367.100 26.330 367.550 ;
        RECT 25.930 366.950 29.880 367.100 ;
        RECT 25.930 366.500 26.330 366.950 ;
        RECT 25.930 366.350 29.880 366.500 ;
        RECT 25.930 365.900 26.330 366.350 ;
        RECT 25.930 365.750 29.880 365.900 ;
        RECT 25.930 365.300 26.330 365.750 ;
        RECT 25.930 365.150 29.880 365.300 ;
        RECT 25.930 364.700 26.330 365.150 ;
        RECT 25.930 364.550 29.880 364.700 ;
        RECT 25.930 364.400 26.330 364.550 ;
        RECT 23.130 364.100 26.330 364.400 ;
        RECT 19.580 363.950 29.880 364.100 ;
        RECT 23.130 363.500 26.330 363.950 ;
        RECT 19.580 363.350 29.880 363.500 ;
        RECT 23.130 362.900 26.330 363.350 ;
        RECT 19.580 362.750 29.880 362.900 ;
        RECT 23.130 362.300 26.330 362.750 ;
        RECT 19.580 362.150 29.880 362.300 ;
        RECT 23.530 361.200 25.930 362.150 ;
        RECT 30.480 361.600 30.630 369.800 ;
        RECT 31.080 361.600 31.230 369.800 ;
        RECT 31.680 361.600 31.830 369.800 ;
        RECT 32.280 361.600 32.430 369.800 ;
        RECT 32.880 361.600 33.030 369.800 ;
        RECT 33.480 361.600 33.630 369.800 ;
        RECT 34.080 361.600 34.230 369.800 ;
        RECT 35.230 370.200 35.380 378.400 ;
        RECT 35.830 370.200 35.980 378.400 ;
        RECT 36.430 370.200 36.580 378.400 ;
        RECT 37.030 370.200 37.180 378.400 ;
        RECT 37.630 370.200 37.780 378.400 ;
        RECT 38.230 370.200 38.380 378.400 ;
        RECT 38.830 370.200 38.980 378.400 ;
        RECT 43.530 377.850 45.940 378.800 ;
        RECT 39.580 377.700 49.880 377.850 ;
        RECT 43.130 377.250 46.330 377.700 ;
        RECT 39.580 377.100 49.880 377.250 ;
        RECT 43.130 376.650 46.330 377.100 ;
        RECT 39.580 376.500 49.880 376.650 ;
        RECT 43.130 376.050 46.330 376.500 ;
        RECT 39.580 375.900 49.880 376.050 ;
        RECT 43.130 375.600 46.330 375.900 ;
        RECT 43.130 375.450 43.530 375.600 ;
        RECT 39.580 375.300 43.530 375.450 ;
        RECT 43.130 374.850 43.530 375.300 ;
        RECT 39.580 374.700 43.530 374.850 ;
        RECT 43.130 374.250 43.530 374.700 ;
        RECT 39.580 374.100 43.530 374.250 ;
        RECT 43.130 373.650 43.530 374.100 ;
        RECT 39.580 373.500 43.530 373.650 ;
        RECT 43.130 373.050 43.530 373.500 ;
        RECT 39.580 372.900 43.530 373.050 ;
        RECT 43.130 372.450 43.530 372.900 ;
        RECT 39.580 372.300 43.530 372.450 ;
        RECT 43.130 371.850 43.530 372.300 ;
        RECT 39.580 371.700 43.530 371.850 ;
        RECT 43.130 371.250 43.530 371.700 ;
        RECT 39.580 371.100 43.530 371.250 ;
        RECT 43.130 370.650 43.530 371.100 ;
        RECT 39.580 370.500 43.530 370.650 ;
        RECT 43.130 370.200 43.530 370.500 ;
        RECT 35.230 369.800 43.530 370.200 ;
        RECT 35.230 361.600 35.380 369.800 ;
        RECT 35.830 361.600 35.980 369.800 ;
        RECT 36.430 361.600 36.580 369.800 ;
        RECT 37.030 361.600 37.180 369.800 ;
        RECT 37.630 361.600 37.780 369.800 ;
        RECT 38.230 361.600 38.380 369.800 ;
        RECT 38.830 361.600 38.980 369.800 ;
        RECT 43.130 369.500 43.530 369.800 ;
        RECT 39.580 369.350 43.530 369.500 ;
        RECT 43.130 368.900 43.530 369.350 ;
        RECT 39.580 368.750 43.530 368.900 ;
        RECT 43.130 368.300 43.530 368.750 ;
        RECT 39.580 368.150 43.530 368.300 ;
        RECT 43.130 367.700 43.530 368.150 ;
        RECT 39.580 367.550 43.530 367.700 ;
        RECT 43.130 367.100 43.530 367.550 ;
        RECT 39.580 366.950 43.530 367.100 ;
        RECT 43.130 366.500 43.530 366.950 ;
        RECT 39.580 366.350 43.530 366.500 ;
        RECT 43.130 365.900 43.530 366.350 ;
        RECT 39.580 365.750 43.530 365.900 ;
        RECT 43.130 365.300 43.530 365.750 ;
        RECT 39.580 365.150 43.530 365.300 ;
        RECT 43.130 364.700 43.530 365.150 ;
        RECT 39.580 364.550 43.530 364.700 ;
        RECT 43.130 364.400 43.530 364.550 ;
        RECT 45.930 375.450 46.330 375.600 ;
        RECT 45.930 375.300 49.880 375.450 ;
        RECT 45.930 374.850 46.330 375.300 ;
        RECT 45.930 374.700 49.880 374.850 ;
        RECT 45.930 374.250 46.330 374.700 ;
        RECT 45.930 374.100 49.880 374.250 ;
        RECT 45.930 373.650 46.330 374.100 ;
        RECT 45.930 373.500 49.880 373.650 ;
        RECT 45.930 373.050 46.330 373.500 ;
        RECT 45.930 372.900 49.880 373.050 ;
        RECT 45.930 372.450 46.330 372.900 ;
        RECT 45.930 372.300 49.880 372.450 ;
        RECT 45.930 371.850 46.330 372.300 ;
        RECT 45.930 371.700 49.880 371.850 ;
        RECT 45.930 371.250 46.330 371.700 ;
        RECT 45.930 371.100 49.880 371.250 ;
        RECT 45.930 370.650 46.330 371.100 ;
        RECT 45.930 370.500 49.880 370.650 ;
        RECT 45.930 370.200 46.330 370.500 ;
        RECT 50.480 370.200 50.630 378.400 ;
        RECT 51.080 370.200 51.230 378.400 ;
        RECT 51.680 370.200 51.830 378.400 ;
        RECT 52.280 370.200 52.430 378.400 ;
        RECT 52.880 370.200 53.030 378.400 ;
        RECT 53.480 370.200 53.630 378.400 ;
        RECT 54.080 370.200 54.230 378.400 ;
        RECT 45.930 369.800 54.230 370.200 ;
        RECT 45.930 369.500 46.330 369.800 ;
        RECT 45.930 369.350 49.880 369.500 ;
        RECT 45.930 368.900 46.330 369.350 ;
        RECT 45.930 368.750 49.880 368.900 ;
        RECT 45.930 368.300 46.330 368.750 ;
        RECT 45.930 368.150 49.880 368.300 ;
        RECT 45.930 367.700 46.330 368.150 ;
        RECT 45.930 367.550 49.880 367.700 ;
        RECT 45.930 367.100 46.330 367.550 ;
        RECT 45.930 366.950 49.880 367.100 ;
        RECT 45.930 366.500 46.330 366.950 ;
        RECT 45.930 366.350 49.880 366.500 ;
        RECT 45.930 365.900 46.330 366.350 ;
        RECT 45.930 365.750 49.880 365.900 ;
        RECT 45.930 365.300 46.330 365.750 ;
        RECT 45.930 365.150 49.880 365.300 ;
        RECT 45.930 364.700 46.330 365.150 ;
        RECT 45.930 364.550 49.880 364.700 ;
        RECT 45.930 364.400 46.330 364.550 ;
        RECT 43.130 364.100 46.330 364.400 ;
        RECT 39.580 363.950 49.880 364.100 ;
        RECT 43.130 363.500 46.330 363.950 ;
        RECT 39.580 363.350 49.880 363.500 ;
        RECT 43.130 362.900 46.330 363.350 ;
        RECT 39.580 362.750 49.880 362.900 ;
        RECT 43.130 362.300 46.330 362.750 ;
        RECT 39.580 362.150 49.880 362.300 ;
        RECT 43.530 361.200 45.930 362.150 ;
        RECT 50.480 361.600 50.630 369.800 ;
        RECT 51.080 361.600 51.230 369.800 ;
        RECT 51.680 361.600 51.830 369.800 ;
        RECT 52.280 361.600 52.430 369.800 ;
        RECT 52.880 361.600 53.030 369.800 ;
        RECT 53.480 361.600 53.630 369.800 ;
        RECT 54.080 361.600 54.230 369.800 ;
        RECT 55.230 370.200 55.380 378.400 ;
        RECT 55.830 370.200 55.980 378.400 ;
        RECT 56.430 370.200 56.580 378.400 ;
        RECT 57.030 370.200 57.180 378.400 ;
        RECT 57.630 370.200 57.780 378.400 ;
        RECT 58.230 370.200 58.380 378.400 ;
        RECT 58.830 370.200 58.980 378.400 ;
        RECT 63.530 377.850 65.940 378.800 ;
        RECT 59.580 377.700 69.880 377.850 ;
        RECT 63.130 377.250 66.330 377.700 ;
        RECT 59.580 377.100 69.880 377.250 ;
        RECT 63.130 376.650 66.330 377.100 ;
        RECT 59.580 376.500 69.880 376.650 ;
        RECT 63.130 376.050 66.330 376.500 ;
        RECT 59.580 375.900 69.880 376.050 ;
        RECT 63.130 375.600 66.330 375.900 ;
        RECT 63.130 375.450 63.530 375.600 ;
        RECT 59.580 375.300 63.530 375.450 ;
        RECT 63.130 374.850 63.530 375.300 ;
        RECT 59.580 374.700 63.530 374.850 ;
        RECT 63.130 374.250 63.530 374.700 ;
        RECT 59.580 374.100 63.530 374.250 ;
        RECT 63.130 373.650 63.530 374.100 ;
        RECT 59.580 373.500 63.530 373.650 ;
        RECT 63.130 373.050 63.530 373.500 ;
        RECT 59.580 372.900 63.530 373.050 ;
        RECT 63.130 372.450 63.530 372.900 ;
        RECT 59.580 372.300 63.530 372.450 ;
        RECT 63.130 371.850 63.530 372.300 ;
        RECT 59.580 371.700 63.530 371.850 ;
        RECT 63.130 371.250 63.530 371.700 ;
        RECT 59.580 371.100 63.530 371.250 ;
        RECT 63.130 370.650 63.530 371.100 ;
        RECT 59.580 370.500 63.530 370.650 ;
        RECT 63.130 370.200 63.530 370.500 ;
        RECT 55.230 369.800 63.530 370.200 ;
        RECT 55.230 361.600 55.380 369.800 ;
        RECT 55.830 361.600 55.980 369.800 ;
        RECT 56.430 361.600 56.580 369.800 ;
        RECT 57.030 361.600 57.180 369.800 ;
        RECT 57.630 361.600 57.780 369.800 ;
        RECT 58.230 361.600 58.380 369.800 ;
        RECT 58.830 361.600 58.980 369.800 ;
        RECT 63.130 369.500 63.530 369.800 ;
        RECT 59.580 369.350 63.530 369.500 ;
        RECT 63.130 368.900 63.530 369.350 ;
        RECT 59.580 368.750 63.530 368.900 ;
        RECT 63.130 368.300 63.530 368.750 ;
        RECT 59.580 368.150 63.530 368.300 ;
        RECT 63.130 367.700 63.530 368.150 ;
        RECT 59.580 367.550 63.530 367.700 ;
        RECT 63.130 367.100 63.530 367.550 ;
        RECT 59.580 366.950 63.530 367.100 ;
        RECT 63.130 366.500 63.530 366.950 ;
        RECT 59.580 366.350 63.530 366.500 ;
        RECT 63.130 365.900 63.530 366.350 ;
        RECT 59.580 365.750 63.530 365.900 ;
        RECT 63.130 365.300 63.530 365.750 ;
        RECT 59.580 365.150 63.530 365.300 ;
        RECT 63.130 364.700 63.530 365.150 ;
        RECT 59.580 364.550 63.530 364.700 ;
        RECT 63.130 364.400 63.530 364.550 ;
        RECT 65.930 375.450 66.330 375.600 ;
        RECT 65.930 375.300 69.880 375.450 ;
        RECT 65.930 374.850 66.330 375.300 ;
        RECT 65.930 374.700 69.880 374.850 ;
        RECT 65.930 374.250 66.330 374.700 ;
        RECT 65.930 374.100 69.880 374.250 ;
        RECT 65.930 373.650 66.330 374.100 ;
        RECT 65.930 373.500 69.880 373.650 ;
        RECT 65.930 373.050 66.330 373.500 ;
        RECT 65.930 372.900 69.880 373.050 ;
        RECT 65.930 372.450 66.330 372.900 ;
        RECT 65.930 372.300 69.880 372.450 ;
        RECT 65.930 371.850 66.330 372.300 ;
        RECT 65.930 371.700 69.880 371.850 ;
        RECT 65.930 371.250 66.330 371.700 ;
        RECT 65.930 371.100 69.880 371.250 ;
        RECT 65.930 370.650 66.330 371.100 ;
        RECT 65.930 370.500 69.880 370.650 ;
        RECT 65.930 370.200 66.330 370.500 ;
        RECT 70.480 370.200 70.630 378.400 ;
        RECT 71.080 370.200 71.230 378.400 ;
        RECT 71.680 370.200 71.830 378.400 ;
        RECT 72.280 370.200 72.430 378.400 ;
        RECT 72.880 370.200 73.030 378.400 ;
        RECT 73.480 370.200 73.630 378.400 ;
        RECT 74.080 370.200 74.230 378.400 ;
        RECT 65.930 369.800 74.230 370.200 ;
        RECT 65.930 369.500 66.330 369.800 ;
        RECT 65.930 369.350 69.880 369.500 ;
        RECT 65.930 368.900 66.330 369.350 ;
        RECT 65.930 368.750 69.880 368.900 ;
        RECT 65.930 368.300 66.330 368.750 ;
        RECT 65.930 368.150 69.880 368.300 ;
        RECT 65.930 367.700 66.330 368.150 ;
        RECT 65.930 367.550 69.880 367.700 ;
        RECT 65.930 367.100 66.330 367.550 ;
        RECT 65.930 366.950 69.880 367.100 ;
        RECT 65.930 366.500 66.330 366.950 ;
        RECT 65.930 366.350 69.880 366.500 ;
        RECT 65.930 365.900 66.330 366.350 ;
        RECT 65.930 365.750 69.880 365.900 ;
        RECT 65.930 365.300 66.330 365.750 ;
        RECT 65.930 365.150 69.880 365.300 ;
        RECT 65.930 364.700 66.330 365.150 ;
        RECT 65.930 364.550 69.880 364.700 ;
        RECT 65.930 364.400 66.330 364.550 ;
        RECT 63.130 364.100 66.330 364.400 ;
        RECT 59.580 363.950 69.880 364.100 ;
        RECT 63.130 363.500 66.330 363.950 ;
        RECT 59.580 363.350 69.880 363.500 ;
        RECT 63.130 362.900 66.330 363.350 ;
        RECT 59.580 362.750 69.880 362.900 ;
        RECT 63.130 362.300 66.330 362.750 ;
        RECT 59.580 362.150 69.880 362.300 ;
        RECT 63.530 361.200 65.930 362.150 ;
        RECT 70.480 361.600 70.630 369.800 ;
        RECT 71.080 361.600 71.230 369.800 ;
        RECT 71.680 361.600 71.830 369.800 ;
        RECT 72.280 361.600 72.430 369.800 ;
        RECT 72.880 361.600 73.030 369.800 ;
        RECT 73.480 361.600 73.630 369.800 ;
        RECT 74.080 361.600 74.230 369.800 ;
        RECT 75.230 370.200 75.380 378.400 ;
        RECT 75.830 370.200 75.980 378.400 ;
        RECT 76.430 370.200 76.580 378.400 ;
        RECT 77.030 370.200 77.180 378.400 ;
        RECT 77.630 370.200 77.780 378.400 ;
        RECT 78.230 370.200 78.380 378.400 ;
        RECT 78.830 370.200 78.980 378.400 ;
        RECT 83.530 377.850 85.940 378.800 ;
        RECT 79.580 377.700 89.880 377.850 ;
        RECT 83.130 377.250 86.330 377.700 ;
        RECT 79.580 377.100 89.880 377.250 ;
        RECT 83.130 376.650 86.330 377.100 ;
        RECT 79.580 376.500 89.880 376.650 ;
        RECT 83.130 376.050 86.330 376.500 ;
        RECT 79.580 375.900 89.880 376.050 ;
        RECT 83.130 375.600 86.330 375.900 ;
        RECT 83.130 375.450 83.530 375.600 ;
        RECT 79.580 375.300 83.530 375.450 ;
        RECT 83.130 374.850 83.530 375.300 ;
        RECT 79.580 374.700 83.530 374.850 ;
        RECT 83.130 374.250 83.530 374.700 ;
        RECT 79.580 374.100 83.530 374.250 ;
        RECT 83.130 373.650 83.530 374.100 ;
        RECT 79.580 373.500 83.530 373.650 ;
        RECT 83.130 373.050 83.530 373.500 ;
        RECT 79.580 372.900 83.530 373.050 ;
        RECT 83.130 372.450 83.530 372.900 ;
        RECT 79.580 372.300 83.530 372.450 ;
        RECT 83.130 371.850 83.530 372.300 ;
        RECT 79.580 371.700 83.530 371.850 ;
        RECT 83.130 371.250 83.530 371.700 ;
        RECT 79.580 371.100 83.530 371.250 ;
        RECT 83.130 370.650 83.530 371.100 ;
        RECT 79.580 370.500 83.530 370.650 ;
        RECT 83.130 370.200 83.530 370.500 ;
        RECT 75.230 369.800 83.530 370.200 ;
        RECT 75.230 361.600 75.380 369.800 ;
        RECT 75.830 361.600 75.980 369.800 ;
        RECT 76.430 361.600 76.580 369.800 ;
        RECT 77.030 361.600 77.180 369.800 ;
        RECT 77.630 361.600 77.780 369.800 ;
        RECT 78.230 361.600 78.380 369.800 ;
        RECT 78.830 361.600 78.980 369.800 ;
        RECT 83.130 369.500 83.530 369.800 ;
        RECT 79.580 369.350 83.530 369.500 ;
        RECT 83.130 368.900 83.530 369.350 ;
        RECT 79.580 368.750 83.530 368.900 ;
        RECT 83.130 368.300 83.530 368.750 ;
        RECT 79.580 368.150 83.530 368.300 ;
        RECT 83.130 367.700 83.530 368.150 ;
        RECT 79.580 367.550 83.530 367.700 ;
        RECT 83.130 367.100 83.530 367.550 ;
        RECT 79.580 366.950 83.530 367.100 ;
        RECT 83.130 366.500 83.530 366.950 ;
        RECT 79.580 366.350 83.530 366.500 ;
        RECT 83.130 365.900 83.530 366.350 ;
        RECT 79.580 365.750 83.530 365.900 ;
        RECT 83.130 365.300 83.530 365.750 ;
        RECT 79.580 365.150 83.530 365.300 ;
        RECT 83.130 364.700 83.530 365.150 ;
        RECT 79.580 364.550 83.530 364.700 ;
        RECT 83.130 364.400 83.530 364.550 ;
        RECT 85.930 375.450 86.330 375.600 ;
        RECT 85.930 375.300 89.880 375.450 ;
        RECT 85.930 374.850 86.330 375.300 ;
        RECT 85.930 374.700 89.880 374.850 ;
        RECT 85.930 374.250 86.330 374.700 ;
        RECT 85.930 374.100 89.880 374.250 ;
        RECT 85.930 373.650 86.330 374.100 ;
        RECT 85.930 373.500 89.880 373.650 ;
        RECT 85.930 373.050 86.330 373.500 ;
        RECT 85.930 372.900 89.880 373.050 ;
        RECT 85.930 372.450 86.330 372.900 ;
        RECT 85.930 372.300 89.880 372.450 ;
        RECT 85.930 371.850 86.330 372.300 ;
        RECT 85.930 371.700 89.880 371.850 ;
        RECT 85.930 371.250 86.330 371.700 ;
        RECT 85.930 371.100 89.880 371.250 ;
        RECT 85.930 370.650 86.330 371.100 ;
        RECT 85.930 370.500 89.880 370.650 ;
        RECT 85.930 370.200 86.330 370.500 ;
        RECT 90.480 370.200 90.630 378.400 ;
        RECT 91.080 370.200 91.230 378.400 ;
        RECT 91.680 370.200 91.830 378.400 ;
        RECT 92.280 370.200 92.430 378.400 ;
        RECT 92.880 370.200 93.030 378.400 ;
        RECT 93.480 370.200 93.630 378.400 ;
        RECT 94.080 370.200 94.230 378.400 ;
        RECT 85.930 369.800 94.230 370.200 ;
        RECT 85.930 369.500 86.330 369.800 ;
        RECT 85.930 369.350 89.880 369.500 ;
        RECT 85.930 368.900 86.330 369.350 ;
        RECT 85.930 368.750 89.880 368.900 ;
        RECT 85.930 368.300 86.330 368.750 ;
        RECT 85.930 368.150 89.880 368.300 ;
        RECT 85.930 367.700 86.330 368.150 ;
        RECT 85.930 367.550 89.880 367.700 ;
        RECT 85.930 367.100 86.330 367.550 ;
        RECT 85.930 366.950 89.880 367.100 ;
        RECT 85.930 366.500 86.330 366.950 ;
        RECT 85.930 366.350 89.880 366.500 ;
        RECT 85.930 365.900 86.330 366.350 ;
        RECT 85.930 365.750 89.880 365.900 ;
        RECT 85.930 365.300 86.330 365.750 ;
        RECT 85.930 365.150 89.880 365.300 ;
        RECT 85.930 364.700 86.330 365.150 ;
        RECT 85.930 364.550 89.880 364.700 ;
        RECT 85.930 364.400 86.330 364.550 ;
        RECT 83.130 364.100 86.330 364.400 ;
        RECT 79.580 363.950 89.880 364.100 ;
        RECT 83.130 363.500 86.330 363.950 ;
        RECT 79.580 363.350 89.880 363.500 ;
        RECT 83.130 362.900 86.330 363.350 ;
        RECT 79.580 362.750 89.880 362.900 ;
        RECT 83.130 362.300 86.330 362.750 ;
        RECT 79.580 362.150 89.880 362.300 ;
        RECT 83.530 361.200 85.930 362.150 ;
        RECT 90.480 361.600 90.630 369.800 ;
        RECT 91.080 361.600 91.230 369.800 ;
        RECT 91.680 361.600 91.830 369.800 ;
        RECT 92.280 361.600 92.430 369.800 ;
        RECT 92.880 361.600 93.030 369.800 ;
        RECT 93.480 361.600 93.630 369.800 ;
        RECT 94.080 361.600 94.230 369.800 ;
        RECT 95.230 370.200 95.380 378.400 ;
        RECT 95.830 370.200 95.980 378.400 ;
        RECT 96.430 370.200 96.580 378.400 ;
        RECT 97.030 370.200 97.180 378.400 ;
        RECT 97.630 370.200 97.780 378.400 ;
        RECT 98.230 370.200 98.380 378.400 ;
        RECT 98.830 370.200 98.980 378.400 ;
        RECT 103.530 377.850 104.730 378.800 ;
        RECT 99.580 377.700 104.730 377.850 ;
        RECT 103.130 377.250 104.730 377.700 ;
        RECT 99.580 377.100 104.730 377.250 ;
        RECT 103.130 376.650 104.730 377.100 ;
        RECT 99.580 376.500 104.730 376.650 ;
        RECT 103.130 376.050 104.730 376.500 ;
        RECT 105.130 376.310 107.130 377.585 ;
        RECT 99.580 375.900 104.730 376.050 ;
        RECT 103.130 375.600 104.730 375.900 ;
        RECT 103.130 375.450 103.530 375.600 ;
        RECT 99.580 375.300 103.530 375.450 ;
        RECT 103.130 374.850 103.530 375.300 ;
        RECT 99.580 374.700 103.530 374.850 ;
        RECT 103.130 374.250 103.530 374.700 ;
        RECT 99.580 374.100 103.530 374.250 ;
        RECT 103.130 373.650 103.530 374.100 ;
        RECT 99.580 373.500 103.530 373.650 ;
        RECT 103.130 373.050 103.530 373.500 ;
        RECT 99.580 372.900 103.530 373.050 ;
        RECT 103.130 372.450 103.530 372.900 ;
        RECT 99.580 372.300 103.530 372.450 ;
        RECT 103.130 371.850 103.530 372.300 ;
        RECT 99.580 371.700 103.530 371.850 ;
        RECT 103.130 371.250 103.530 371.700 ;
        RECT 99.580 371.100 103.530 371.250 ;
        RECT 103.130 370.650 103.530 371.100 ;
        RECT 99.580 370.500 103.530 370.650 ;
        RECT 103.130 370.200 103.530 370.500 ;
        RECT 95.230 369.800 103.530 370.200 ;
        RECT 95.230 361.600 95.380 369.800 ;
        RECT 95.830 361.600 95.980 369.800 ;
        RECT 96.430 361.600 96.580 369.800 ;
        RECT 97.030 361.600 97.180 369.800 ;
        RECT 97.630 361.600 97.780 369.800 ;
        RECT 98.230 361.600 98.380 369.800 ;
        RECT 98.830 361.600 98.980 369.800 ;
        RECT 103.130 369.500 103.530 369.800 ;
        RECT 99.580 369.350 103.530 369.500 ;
        RECT 103.130 368.900 103.530 369.350 ;
        RECT 99.580 368.750 103.530 368.900 ;
        RECT 103.130 368.300 103.530 368.750 ;
        RECT 99.580 368.150 103.530 368.300 ;
        RECT 103.130 367.700 103.530 368.150 ;
        RECT 99.580 367.550 103.530 367.700 ;
        RECT 103.130 367.100 103.530 367.550 ;
        RECT 99.580 366.950 103.530 367.100 ;
        RECT 103.130 366.500 103.530 366.950 ;
        RECT 99.580 366.350 103.530 366.500 ;
        RECT 103.130 365.900 103.530 366.350 ;
        RECT 99.580 365.750 103.530 365.900 ;
        RECT 103.130 365.300 103.530 365.750 ;
        RECT 99.580 365.150 103.530 365.300 ;
        RECT 103.130 364.700 103.530 365.150 ;
        RECT 99.580 364.550 103.530 364.700 ;
        RECT 103.130 364.400 103.530 364.550 ;
        RECT 103.130 364.100 104.730 364.400 ;
        RECT 99.580 363.950 104.730 364.100 ;
        RECT 103.130 363.500 104.730 363.950 ;
        RECT 99.580 363.350 104.730 363.500 ;
        RECT 103.130 362.900 104.730 363.350 ;
        RECT 99.580 362.750 104.730 362.900 ;
        RECT 103.130 362.300 104.730 362.750 ;
        RECT 105.140 362.325 107.140 363.600 ;
        RECT 99.580 362.150 104.730 362.300 ;
        RECT 103.530 361.200 104.730 362.150 ;
        RECT 4.730 358.800 9.130 361.200 ;
        RECT 20.330 358.800 29.130 361.200 ;
        RECT 40.330 358.800 49.130 361.200 ;
        RECT 60.330 358.800 69.130 361.200 ;
        RECT 80.330 358.800 89.130 361.200 ;
        RECT 100.330 358.800 104.730 361.200 ;
        RECT 4.730 357.850 5.940 358.800 ;
        RECT 4.730 357.700 9.880 357.850 ;
        RECT 2.315 356.110 4.320 357.385 ;
        RECT 4.730 357.250 6.330 357.700 ;
        RECT 4.730 357.100 9.880 357.250 ;
        RECT 4.730 356.650 6.330 357.100 ;
        RECT 4.730 356.500 9.880 356.650 ;
        RECT 4.730 356.050 6.330 356.500 ;
        RECT 4.730 355.900 9.880 356.050 ;
        RECT 4.730 355.600 6.330 355.900 ;
        RECT 2.315 353.250 4.315 355.545 ;
        RECT 5.930 355.450 6.330 355.600 ;
        RECT 5.930 355.300 9.880 355.450 ;
        RECT 5.930 354.850 6.330 355.300 ;
        RECT 5.930 354.700 9.880 354.850 ;
        RECT 5.930 354.250 6.330 354.700 ;
        RECT 5.930 354.100 9.880 354.250 ;
        RECT 5.930 353.650 6.330 354.100 ;
        RECT 5.930 353.500 9.880 353.650 ;
        RECT 5.930 353.050 6.330 353.500 ;
        RECT 5.930 352.900 9.880 353.050 ;
        RECT 5.930 352.450 6.330 352.900 ;
        RECT 5.930 352.300 9.880 352.450 ;
        RECT 5.930 351.850 6.330 352.300 ;
        RECT 5.930 351.700 9.880 351.850 ;
        RECT 5.930 351.250 6.330 351.700 ;
        RECT 5.930 351.100 9.880 351.250 ;
        RECT 5.930 350.650 6.330 351.100 ;
        RECT 5.930 350.500 9.880 350.650 ;
        RECT 5.930 350.200 6.330 350.500 ;
        RECT 10.480 350.200 10.630 358.400 ;
        RECT 11.080 350.200 11.230 358.400 ;
        RECT 11.680 350.200 11.830 358.400 ;
        RECT 12.280 350.200 12.430 358.400 ;
        RECT 12.880 350.200 13.030 358.400 ;
        RECT 13.480 350.200 13.630 358.400 ;
        RECT 14.080 350.200 14.230 358.400 ;
        RECT 5.930 349.800 14.230 350.200 ;
        RECT 5.930 349.500 6.330 349.800 ;
        RECT 5.930 349.350 9.880 349.500 ;
        RECT 5.930 348.900 6.330 349.350 ;
        RECT 5.930 348.750 9.880 348.900 ;
        RECT 5.930 348.300 6.330 348.750 ;
        RECT 5.930 348.150 9.880 348.300 ;
        RECT 5.930 347.700 6.330 348.150 ;
        RECT 5.930 347.550 9.880 347.700 ;
        RECT 5.930 347.100 6.330 347.550 ;
        RECT 5.930 346.950 9.880 347.100 ;
        RECT 2.315 344.450 4.315 346.745 ;
        RECT 5.930 346.500 6.330 346.950 ;
        RECT 5.930 346.350 9.880 346.500 ;
        RECT 5.930 345.900 6.330 346.350 ;
        RECT 5.930 345.750 9.880 345.900 ;
        RECT 5.930 345.300 6.330 345.750 ;
        RECT 5.930 345.150 9.880 345.300 ;
        RECT 5.930 344.700 6.330 345.150 ;
        RECT 5.930 344.550 9.880 344.700 ;
        RECT 5.930 344.400 6.330 344.550 ;
        RECT 4.730 344.100 6.330 344.400 ;
        RECT 2.315 342.745 4.320 344.020 ;
        RECT 4.730 343.950 9.880 344.100 ;
        RECT 4.730 343.500 6.330 343.950 ;
        RECT 4.730 343.350 9.880 343.500 ;
        RECT 4.730 342.900 6.330 343.350 ;
        RECT 4.730 342.750 9.880 342.900 ;
        RECT 4.730 342.300 6.330 342.750 ;
        RECT 4.730 342.150 9.880 342.300 ;
        RECT 4.730 341.200 5.930 342.150 ;
        RECT 10.480 341.600 10.630 349.800 ;
        RECT 11.080 341.600 11.230 349.800 ;
        RECT 11.680 341.600 11.830 349.800 ;
        RECT 12.280 341.600 12.430 349.800 ;
        RECT 12.880 341.600 13.030 349.800 ;
        RECT 13.480 341.600 13.630 349.800 ;
        RECT 14.080 341.600 14.230 349.800 ;
        RECT 15.230 350.200 15.380 358.400 ;
        RECT 15.830 350.200 15.980 358.400 ;
        RECT 16.430 350.200 16.580 358.400 ;
        RECT 17.030 350.200 17.180 358.400 ;
        RECT 17.630 350.200 17.780 358.400 ;
        RECT 18.230 350.200 18.380 358.400 ;
        RECT 18.830 350.200 18.980 358.400 ;
        RECT 23.530 357.850 25.940 358.800 ;
        RECT 19.580 357.700 29.880 357.850 ;
        RECT 23.130 357.250 26.330 357.700 ;
        RECT 19.580 357.100 29.880 357.250 ;
        RECT 23.130 356.650 26.330 357.100 ;
        RECT 19.580 356.500 29.880 356.650 ;
        RECT 23.130 356.050 26.330 356.500 ;
        RECT 19.580 355.900 29.880 356.050 ;
        RECT 23.130 355.600 26.330 355.900 ;
        RECT 23.130 355.450 23.530 355.600 ;
        RECT 19.580 355.300 23.530 355.450 ;
        RECT 23.130 354.850 23.530 355.300 ;
        RECT 19.580 354.700 23.530 354.850 ;
        RECT 23.130 354.250 23.530 354.700 ;
        RECT 19.580 354.100 23.530 354.250 ;
        RECT 23.130 353.650 23.530 354.100 ;
        RECT 19.580 353.500 23.530 353.650 ;
        RECT 23.130 353.050 23.530 353.500 ;
        RECT 19.580 352.900 23.530 353.050 ;
        RECT 23.130 352.450 23.530 352.900 ;
        RECT 19.580 352.300 23.530 352.450 ;
        RECT 23.130 351.850 23.530 352.300 ;
        RECT 19.580 351.700 23.530 351.850 ;
        RECT 23.130 351.250 23.530 351.700 ;
        RECT 19.580 351.100 23.530 351.250 ;
        RECT 23.130 350.650 23.530 351.100 ;
        RECT 19.580 350.500 23.530 350.650 ;
        RECT 23.130 350.200 23.530 350.500 ;
        RECT 15.230 349.800 23.530 350.200 ;
        RECT 15.230 341.600 15.380 349.800 ;
        RECT 15.830 341.600 15.980 349.800 ;
        RECT 16.430 341.600 16.580 349.800 ;
        RECT 17.030 341.600 17.180 349.800 ;
        RECT 17.630 341.600 17.780 349.800 ;
        RECT 18.230 341.600 18.380 349.800 ;
        RECT 18.830 341.600 18.980 349.800 ;
        RECT 23.130 349.500 23.530 349.800 ;
        RECT 19.580 349.350 23.530 349.500 ;
        RECT 23.130 348.900 23.530 349.350 ;
        RECT 19.580 348.750 23.530 348.900 ;
        RECT 23.130 348.300 23.530 348.750 ;
        RECT 19.580 348.150 23.530 348.300 ;
        RECT 23.130 347.700 23.530 348.150 ;
        RECT 19.580 347.550 23.530 347.700 ;
        RECT 23.130 347.100 23.530 347.550 ;
        RECT 19.580 346.950 23.530 347.100 ;
        RECT 23.130 346.500 23.530 346.950 ;
        RECT 19.580 346.350 23.530 346.500 ;
        RECT 23.130 345.900 23.530 346.350 ;
        RECT 19.580 345.750 23.530 345.900 ;
        RECT 23.130 345.300 23.530 345.750 ;
        RECT 19.580 345.150 23.530 345.300 ;
        RECT 23.130 344.700 23.530 345.150 ;
        RECT 19.580 344.550 23.530 344.700 ;
        RECT 23.130 344.400 23.530 344.550 ;
        RECT 25.930 355.450 26.330 355.600 ;
        RECT 25.930 355.300 29.880 355.450 ;
        RECT 25.930 354.850 26.330 355.300 ;
        RECT 25.930 354.700 29.880 354.850 ;
        RECT 25.930 354.250 26.330 354.700 ;
        RECT 25.930 354.100 29.880 354.250 ;
        RECT 25.930 353.650 26.330 354.100 ;
        RECT 25.930 353.500 29.880 353.650 ;
        RECT 25.930 353.050 26.330 353.500 ;
        RECT 25.930 352.900 29.880 353.050 ;
        RECT 25.930 352.450 26.330 352.900 ;
        RECT 25.930 352.300 29.880 352.450 ;
        RECT 25.930 351.850 26.330 352.300 ;
        RECT 25.930 351.700 29.880 351.850 ;
        RECT 25.930 351.250 26.330 351.700 ;
        RECT 25.930 351.100 29.880 351.250 ;
        RECT 25.930 350.650 26.330 351.100 ;
        RECT 25.930 350.500 29.880 350.650 ;
        RECT 25.930 350.200 26.330 350.500 ;
        RECT 30.480 350.200 30.630 358.400 ;
        RECT 31.080 350.200 31.230 358.400 ;
        RECT 31.680 350.200 31.830 358.400 ;
        RECT 32.280 350.200 32.430 358.400 ;
        RECT 32.880 350.200 33.030 358.400 ;
        RECT 33.480 350.200 33.630 358.400 ;
        RECT 34.080 350.200 34.230 358.400 ;
        RECT 25.930 349.800 34.230 350.200 ;
        RECT 25.930 349.500 26.330 349.800 ;
        RECT 25.930 349.350 29.880 349.500 ;
        RECT 25.930 348.900 26.330 349.350 ;
        RECT 25.930 348.750 29.880 348.900 ;
        RECT 25.930 348.300 26.330 348.750 ;
        RECT 25.930 348.150 29.880 348.300 ;
        RECT 25.930 347.700 26.330 348.150 ;
        RECT 25.930 347.550 29.880 347.700 ;
        RECT 25.930 347.100 26.330 347.550 ;
        RECT 25.930 346.950 29.880 347.100 ;
        RECT 25.930 346.500 26.330 346.950 ;
        RECT 25.930 346.350 29.880 346.500 ;
        RECT 25.930 345.900 26.330 346.350 ;
        RECT 25.930 345.750 29.880 345.900 ;
        RECT 25.930 345.300 26.330 345.750 ;
        RECT 25.930 345.150 29.880 345.300 ;
        RECT 25.930 344.700 26.330 345.150 ;
        RECT 25.930 344.550 29.880 344.700 ;
        RECT 25.930 344.400 26.330 344.550 ;
        RECT 23.130 344.100 26.330 344.400 ;
        RECT 19.580 343.950 29.880 344.100 ;
        RECT 23.130 343.500 26.330 343.950 ;
        RECT 19.580 343.350 29.880 343.500 ;
        RECT 23.130 342.900 26.330 343.350 ;
        RECT 19.580 342.750 29.880 342.900 ;
        RECT 23.130 342.300 26.330 342.750 ;
        RECT 19.580 342.150 29.880 342.300 ;
        RECT 23.530 341.200 25.930 342.150 ;
        RECT 30.480 341.600 30.630 349.800 ;
        RECT 31.080 341.600 31.230 349.800 ;
        RECT 31.680 341.600 31.830 349.800 ;
        RECT 32.280 341.600 32.430 349.800 ;
        RECT 32.880 341.600 33.030 349.800 ;
        RECT 33.480 341.600 33.630 349.800 ;
        RECT 34.080 341.600 34.230 349.800 ;
        RECT 35.230 350.200 35.380 358.400 ;
        RECT 35.830 350.200 35.980 358.400 ;
        RECT 36.430 350.200 36.580 358.400 ;
        RECT 37.030 350.200 37.180 358.400 ;
        RECT 37.630 350.200 37.780 358.400 ;
        RECT 38.230 350.200 38.380 358.400 ;
        RECT 38.830 350.200 38.980 358.400 ;
        RECT 43.530 357.850 45.940 358.800 ;
        RECT 39.580 357.700 49.880 357.850 ;
        RECT 43.130 357.250 46.330 357.700 ;
        RECT 39.580 357.100 49.880 357.250 ;
        RECT 43.130 356.650 46.330 357.100 ;
        RECT 39.580 356.500 49.880 356.650 ;
        RECT 43.130 356.050 46.330 356.500 ;
        RECT 39.580 355.900 49.880 356.050 ;
        RECT 43.130 355.600 46.330 355.900 ;
        RECT 43.130 355.450 43.530 355.600 ;
        RECT 39.580 355.300 43.530 355.450 ;
        RECT 43.130 354.850 43.530 355.300 ;
        RECT 39.580 354.700 43.530 354.850 ;
        RECT 43.130 354.250 43.530 354.700 ;
        RECT 39.580 354.100 43.530 354.250 ;
        RECT 43.130 353.650 43.530 354.100 ;
        RECT 39.580 353.500 43.530 353.650 ;
        RECT 43.130 353.050 43.530 353.500 ;
        RECT 39.580 352.900 43.530 353.050 ;
        RECT 43.130 352.450 43.530 352.900 ;
        RECT 39.580 352.300 43.530 352.450 ;
        RECT 43.130 351.850 43.530 352.300 ;
        RECT 39.580 351.700 43.530 351.850 ;
        RECT 43.130 351.250 43.530 351.700 ;
        RECT 39.580 351.100 43.530 351.250 ;
        RECT 43.130 350.650 43.530 351.100 ;
        RECT 39.580 350.500 43.530 350.650 ;
        RECT 43.130 350.200 43.530 350.500 ;
        RECT 35.230 349.800 43.530 350.200 ;
        RECT 35.230 341.600 35.380 349.800 ;
        RECT 35.830 341.600 35.980 349.800 ;
        RECT 36.430 341.600 36.580 349.800 ;
        RECT 37.030 341.600 37.180 349.800 ;
        RECT 37.630 341.600 37.780 349.800 ;
        RECT 38.230 341.600 38.380 349.800 ;
        RECT 38.830 341.600 38.980 349.800 ;
        RECT 43.130 349.500 43.530 349.800 ;
        RECT 39.580 349.350 43.530 349.500 ;
        RECT 43.130 348.900 43.530 349.350 ;
        RECT 39.580 348.750 43.530 348.900 ;
        RECT 43.130 348.300 43.530 348.750 ;
        RECT 39.580 348.150 43.530 348.300 ;
        RECT 43.130 347.700 43.530 348.150 ;
        RECT 39.580 347.550 43.530 347.700 ;
        RECT 43.130 347.100 43.530 347.550 ;
        RECT 39.580 346.950 43.530 347.100 ;
        RECT 43.130 346.500 43.530 346.950 ;
        RECT 39.580 346.350 43.530 346.500 ;
        RECT 43.130 345.900 43.530 346.350 ;
        RECT 39.580 345.750 43.530 345.900 ;
        RECT 43.130 345.300 43.530 345.750 ;
        RECT 39.580 345.150 43.530 345.300 ;
        RECT 43.130 344.700 43.530 345.150 ;
        RECT 39.580 344.550 43.530 344.700 ;
        RECT 43.130 344.400 43.530 344.550 ;
        RECT 45.930 355.450 46.330 355.600 ;
        RECT 45.930 355.300 49.880 355.450 ;
        RECT 45.930 354.850 46.330 355.300 ;
        RECT 45.930 354.700 49.880 354.850 ;
        RECT 45.930 354.250 46.330 354.700 ;
        RECT 45.930 354.100 49.880 354.250 ;
        RECT 45.930 353.650 46.330 354.100 ;
        RECT 45.930 353.500 49.880 353.650 ;
        RECT 45.930 353.050 46.330 353.500 ;
        RECT 45.930 352.900 49.880 353.050 ;
        RECT 45.930 352.450 46.330 352.900 ;
        RECT 45.930 352.300 49.880 352.450 ;
        RECT 45.930 351.850 46.330 352.300 ;
        RECT 45.930 351.700 49.880 351.850 ;
        RECT 45.930 351.250 46.330 351.700 ;
        RECT 45.930 351.100 49.880 351.250 ;
        RECT 45.930 350.650 46.330 351.100 ;
        RECT 45.930 350.500 49.880 350.650 ;
        RECT 45.930 350.200 46.330 350.500 ;
        RECT 50.480 350.200 50.630 358.400 ;
        RECT 51.080 350.200 51.230 358.400 ;
        RECT 51.680 350.200 51.830 358.400 ;
        RECT 52.280 350.200 52.430 358.400 ;
        RECT 52.880 350.200 53.030 358.400 ;
        RECT 53.480 350.200 53.630 358.400 ;
        RECT 54.080 350.200 54.230 358.400 ;
        RECT 45.930 349.800 54.230 350.200 ;
        RECT 45.930 349.500 46.330 349.800 ;
        RECT 45.930 349.350 49.880 349.500 ;
        RECT 45.930 348.900 46.330 349.350 ;
        RECT 45.930 348.750 49.880 348.900 ;
        RECT 45.930 348.300 46.330 348.750 ;
        RECT 45.930 348.150 49.880 348.300 ;
        RECT 45.930 347.700 46.330 348.150 ;
        RECT 45.930 347.550 49.880 347.700 ;
        RECT 45.930 347.100 46.330 347.550 ;
        RECT 45.930 346.950 49.880 347.100 ;
        RECT 45.930 346.500 46.330 346.950 ;
        RECT 45.930 346.350 49.880 346.500 ;
        RECT 45.930 345.900 46.330 346.350 ;
        RECT 45.930 345.750 49.880 345.900 ;
        RECT 45.930 345.300 46.330 345.750 ;
        RECT 45.930 345.150 49.880 345.300 ;
        RECT 45.930 344.700 46.330 345.150 ;
        RECT 45.930 344.550 49.880 344.700 ;
        RECT 45.930 344.400 46.330 344.550 ;
        RECT 43.130 344.100 46.330 344.400 ;
        RECT 39.580 343.950 49.880 344.100 ;
        RECT 43.130 343.500 46.330 343.950 ;
        RECT 39.580 343.350 49.880 343.500 ;
        RECT 43.130 342.900 46.330 343.350 ;
        RECT 39.580 342.750 49.880 342.900 ;
        RECT 43.130 342.300 46.330 342.750 ;
        RECT 39.580 342.150 49.880 342.300 ;
        RECT 43.530 341.200 45.930 342.150 ;
        RECT 50.480 341.600 50.630 349.800 ;
        RECT 51.080 341.600 51.230 349.800 ;
        RECT 51.680 341.600 51.830 349.800 ;
        RECT 52.280 341.600 52.430 349.800 ;
        RECT 52.880 341.600 53.030 349.800 ;
        RECT 53.480 341.600 53.630 349.800 ;
        RECT 54.080 341.600 54.230 349.800 ;
        RECT 55.230 350.200 55.380 358.400 ;
        RECT 55.830 350.200 55.980 358.400 ;
        RECT 56.430 350.200 56.580 358.400 ;
        RECT 57.030 350.200 57.180 358.400 ;
        RECT 57.630 350.200 57.780 358.400 ;
        RECT 58.230 350.200 58.380 358.400 ;
        RECT 58.830 350.200 58.980 358.400 ;
        RECT 63.530 357.850 65.940 358.800 ;
        RECT 59.580 357.700 69.880 357.850 ;
        RECT 63.130 357.250 66.330 357.700 ;
        RECT 59.580 357.100 69.880 357.250 ;
        RECT 63.130 356.650 66.330 357.100 ;
        RECT 59.580 356.500 69.880 356.650 ;
        RECT 63.130 356.050 66.330 356.500 ;
        RECT 59.580 355.900 69.880 356.050 ;
        RECT 63.130 355.600 66.330 355.900 ;
        RECT 63.130 355.450 63.530 355.600 ;
        RECT 59.580 355.300 63.530 355.450 ;
        RECT 63.130 354.850 63.530 355.300 ;
        RECT 59.580 354.700 63.530 354.850 ;
        RECT 63.130 354.250 63.530 354.700 ;
        RECT 59.580 354.100 63.530 354.250 ;
        RECT 63.130 353.650 63.530 354.100 ;
        RECT 59.580 353.500 63.530 353.650 ;
        RECT 63.130 353.050 63.530 353.500 ;
        RECT 59.580 352.900 63.530 353.050 ;
        RECT 63.130 352.450 63.530 352.900 ;
        RECT 59.580 352.300 63.530 352.450 ;
        RECT 63.130 351.850 63.530 352.300 ;
        RECT 59.580 351.700 63.530 351.850 ;
        RECT 63.130 351.250 63.530 351.700 ;
        RECT 59.580 351.100 63.530 351.250 ;
        RECT 63.130 350.650 63.530 351.100 ;
        RECT 59.580 350.500 63.530 350.650 ;
        RECT 63.130 350.200 63.530 350.500 ;
        RECT 55.230 349.800 63.530 350.200 ;
        RECT 55.230 341.600 55.380 349.800 ;
        RECT 55.830 341.600 55.980 349.800 ;
        RECT 56.430 341.600 56.580 349.800 ;
        RECT 57.030 341.600 57.180 349.800 ;
        RECT 57.630 341.600 57.780 349.800 ;
        RECT 58.230 341.600 58.380 349.800 ;
        RECT 58.830 341.600 58.980 349.800 ;
        RECT 63.130 349.500 63.530 349.800 ;
        RECT 59.580 349.350 63.530 349.500 ;
        RECT 63.130 348.900 63.530 349.350 ;
        RECT 59.580 348.750 63.530 348.900 ;
        RECT 63.130 348.300 63.530 348.750 ;
        RECT 59.580 348.150 63.530 348.300 ;
        RECT 63.130 347.700 63.530 348.150 ;
        RECT 59.580 347.550 63.530 347.700 ;
        RECT 63.130 347.100 63.530 347.550 ;
        RECT 59.580 346.950 63.530 347.100 ;
        RECT 63.130 346.500 63.530 346.950 ;
        RECT 59.580 346.350 63.530 346.500 ;
        RECT 63.130 345.900 63.530 346.350 ;
        RECT 59.580 345.750 63.530 345.900 ;
        RECT 63.130 345.300 63.530 345.750 ;
        RECT 59.580 345.150 63.530 345.300 ;
        RECT 63.130 344.700 63.530 345.150 ;
        RECT 59.580 344.550 63.530 344.700 ;
        RECT 63.130 344.400 63.530 344.550 ;
        RECT 65.930 355.450 66.330 355.600 ;
        RECT 65.930 355.300 69.880 355.450 ;
        RECT 65.930 354.850 66.330 355.300 ;
        RECT 65.930 354.700 69.880 354.850 ;
        RECT 65.930 354.250 66.330 354.700 ;
        RECT 65.930 354.100 69.880 354.250 ;
        RECT 65.930 353.650 66.330 354.100 ;
        RECT 65.930 353.500 69.880 353.650 ;
        RECT 65.930 353.050 66.330 353.500 ;
        RECT 65.930 352.900 69.880 353.050 ;
        RECT 65.930 352.450 66.330 352.900 ;
        RECT 65.930 352.300 69.880 352.450 ;
        RECT 65.930 351.850 66.330 352.300 ;
        RECT 65.930 351.700 69.880 351.850 ;
        RECT 65.930 351.250 66.330 351.700 ;
        RECT 65.930 351.100 69.880 351.250 ;
        RECT 65.930 350.650 66.330 351.100 ;
        RECT 65.930 350.500 69.880 350.650 ;
        RECT 65.930 350.200 66.330 350.500 ;
        RECT 70.480 350.200 70.630 358.400 ;
        RECT 71.080 350.200 71.230 358.400 ;
        RECT 71.680 350.200 71.830 358.400 ;
        RECT 72.280 350.200 72.430 358.400 ;
        RECT 72.880 350.200 73.030 358.400 ;
        RECT 73.480 350.200 73.630 358.400 ;
        RECT 74.080 350.200 74.230 358.400 ;
        RECT 65.930 349.800 74.230 350.200 ;
        RECT 65.930 349.500 66.330 349.800 ;
        RECT 65.930 349.350 69.880 349.500 ;
        RECT 65.930 348.900 66.330 349.350 ;
        RECT 65.930 348.750 69.880 348.900 ;
        RECT 65.930 348.300 66.330 348.750 ;
        RECT 65.930 348.150 69.880 348.300 ;
        RECT 65.930 347.700 66.330 348.150 ;
        RECT 65.930 347.550 69.880 347.700 ;
        RECT 65.930 347.100 66.330 347.550 ;
        RECT 65.930 346.950 69.880 347.100 ;
        RECT 65.930 346.500 66.330 346.950 ;
        RECT 65.930 346.350 69.880 346.500 ;
        RECT 65.930 345.900 66.330 346.350 ;
        RECT 65.930 345.750 69.880 345.900 ;
        RECT 65.930 345.300 66.330 345.750 ;
        RECT 65.930 345.150 69.880 345.300 ;
        RECT 65.930 344.700 66.330 345.150 ;
        RECT 65.930 344.550 69.880 344.700 ;
        RECT 65.930 344.400 66.330 344.550 ;
        RECT 63.130 344.100 66.330 344.400 ;
        RECT 59.580 343.950 69.880 344.100 ;
        RECT 63.130 343.500 66.330 343.950 ;
        RECT 59.580 343.350 69.880 343.500 ;
        RECT 63.130 342.900 66.330 343.350 ;
        RECT 59.580 342.750 69.880 342.900 ;
        RECT 63.130 342.300 66.330 342.750 ;
        RECT 59.580 342.150 69.880 342.300 ;
        RECT 63.530 341.200 65.930 342.150 ;
        RECT 70.480 341.600 70.630 349.800 ;
        RECT 71.080 341.600 71.230 349.800 ;
        RECT 71.680 341.600 71.830 349.800 ;
        RECT 72.280 341.600 72.430 349.800 ;
        RECT 72.880 341.600 73.030 349.800 ;
        RECT 73.480 341.600 73.630 349.800 ;
        RECT 74.080 341.600 74.230 349.800 ;
        RECT 75.230 350.200 75.380 358.400 ;
        RECT 75.830 350.200 75.980 358.400 ;
        RECT 76.430 350.200 76.580 358.400 ;
        RECT 77.030 350.200 77.180 358.400 ;
        RECT 77.630 350.200 77.780 358.400 ;
        RECT 78.230 350.200 78.380 358.400 ;
        RECT 78.830 350.200 78.980 358.400 ;
        RECT 83.530 357.850 85.940 358.800 ;
        RECT 79.580 357.700 89.880 357.850 ;
        RECT 83.130 357.250 86.330 357.700 ;
        RECT 79.580 357.100 89.880 357.250 ;
        RECT 83.130 356.650 86.330 357.100 ;
        RECT 79.580 356.500 89.880 356.650 ;
        RECT 83.130 356.050 86.330 356.500 ;
        RECT 79.580 355.900 89.880 356.050 ;
        RECT 83.130 355.600 86.330 355.900 ;
        RECT 83.130 355.450 83.530 355.600 ;
        RECT 79.580 355.300 83.530 355.450 ;
        RECT 83.130 354.850 83.530 355.300 ;
        RECT 79.580 354.700 83.530 354.850 ;
        RECT 83.130 354.250 83.530 354.700 ;
        RECT 79.580 354.100 83.530 354.250 ;
        RECT 83.130 353.650 83.530 354.100 ;
        RECT 79.580 353.500 83.530 353.650 ;
        RECT 83.130 353.050 83.530 353.500 ;
        RECT 79.580 352.900 83.530 353.050 ;
        RECT 83.130 352.450 83.530 352.900 ;
        RECT 79.580 352.300 83.530 352.450 ;
        RECT 83.130 351.850 83.530 352.300 ;
        RECT 79.580 351.700 83.530 351.850 ;
        RECT 83.130 351.250 83.530 351.700 ;
        RECT 79.580 351.100 83.530 351.250 ;
        RECT 83.130 350.650 83.530 351.100 ;
        RECT 79.580 350.500 83.530 350.650 ;
        RECT 83.130 350.200 83.530 350.500 ;
        RECT 75.230 349.800 83.530 350.200 ;
        RECT 75.230 341.600 75.380 349.800 ;
        RECT 75.830 341.600 75.980 349.800 ;
        RECT 76.430 341.600 76.580 349.800 ;
        RECT 77.030 341.600 77.180 349.800 ;
        RECT 77.630 341.600 77.780 349.800 ;
        RECT 78.230 341.600 78.380 349.800 ;
        RECT 78.830 341.600 78.980 349.800 ;
        RECT 83.130 349.500 83.530 349.800 ;
        RECT 79.580 349.350 83.530 349.500 ;
        RECT 83.130 348.900 83.530 349.350 ;
        RECT 79.580 348.750 83.530 348.900 ;
        RECT 83.130 348.300 83.530 348.750 ;
        RECT 79.580 348.150 83.530 348.300 ;
        RECT 83.130 347.700 83.530 348.150 ;
        RECT 79.580 347.550 83.530 347.700 ;
        RECT 83.130 347.100 83.530 347.550 ;
        RECT 79.580 346.950 83.530 347.100 ;
        RECT 83.130 346.500 83.530 346.950 ;
        RECT 79.580 346.350 83.530 346.500 ;
        RECT 83.130 345.900 83.530 346.350 ;
        RECT 79.580 345.750 83.530 345.900 ;
        RECT 83.130 345.300 83.530 345.750 ;
        RECT 79.580 345.150 83.530 345.300 ;
        RECT 83.130 344.700 83.530 345.150 ;
        RECT 79.580 344.550 83.530 344.700 ;
        RECT 83.130 344.400 83.530 344.550 ;
        RECT 85.930 355.450 86.330 355.600 ;
        RECT 85.930 355.300 89.880 355.450 ;
        RECT 85.930 354.850 86.330 355.300 ;
        RECT 85.930 354.700 89.880 354.850 ;
        RECT 85.930 354.250 86.330 354.700 ;
        RECT 85.930 354.100 89.880 354.250 ;
        RECT 85.930 353.650 86.330 354.100 ;
        RECT 85.930 353.500 89.880 353.650 ;
        RECT 85.930 353.050 86.330 353.500 ;
        RECT 85.930 352.900 89.880 353.050 ;
        RECT 85.930 352.450 86.330 352.900 ;
        RECT 85.930 352.300 89.880 352.450 ;
        RECT 85.930 351.850 86.330 352.300 ;
        RECT 85.930 351.700 89.880 351.850 ;
        RECT 85.930 351.250 86.330 351.700 ;
        RECT 85.930 351.100 89.880 351.250 ;
        RECT 85.930 350.650 86.330 351.100 ;
        RECT 85.930 350.500 89.880 350.650 ;
        RECT 85.930 350.200 86.330 350.500 ;
        RECT 90.480 350.200 90.630 358.400 ;
        RECT 91.080 350.200 91.230 358.400 ;
        RECT 91.680 350.200 91.830 358.400 ;
        RECT 92.280 350.200 92.430 358.400 ;
        RECT 92.880 350.200 93.030 358.400 ;
        RECT 93.480 350.200 93.630 358.400 ;
        RECT 94.080 350.200 94.230 358.400 ;
        RECT 85.930 349.800 94.230 350.200 ;
        RECT 85.930 349.500 86.330 349.800 ;
        RECT 85.930 349.350 89.880 349.500 ;
        RECT 85.930 348.900 86.330 349.350 ;
        RECT 85.930 348.750 89.880 348.900 ;
        RECT 85.930 348.300 86.330 348.750 ;
        RECT 85.930 348.150 89.880 348.300 ;
        RECT 85.930 347.700 86.330 348.150 ;
        RECT 85.930 347.550 89.880 347.700 ;
        RECT 85.930 347.100 86.330 347.550 ;
        RECT 85.930 346.950 89.880 347.100 ;
        RECT 85.930 346.500 86.330 346.950 ;
        RECT 85.930 346.350 89.880 346.500 ;
        RECT 85.930 345.900 86.330 346.350 ;
        RECT 85.930 345.750 89.880 345.900 ;
        RECT 85.930 345.300 86.330 345.750 ;
        RECT 85.930 345.150 89.880 345.300 ;
        RECT 85.930 344.700 86.330 345.150 ;
        RECT 85.930 344.550 89.880 344.700 ;
        RECT 85.930 344.400 86.330 344.550 ;
        RECT 83.130 344.100 86.330 344.400 ;
        RECT 79.580 343.950 89.880 344.100 ;
        RECT 83.130 343.500 86.330 343.950 ;
        RECT 79.580 343.350 89.880 343.500 ;
        RECT 83.130 342.900 86.330 343.350 ;
        RECT 79.580 342.750 89.880 342.900 ;
        RECT 83.130 342.300 86.330 342.750 ;
        RECT 79.580 342.150 89.880 342.300 ;
        RECT 83.530 341.200 85.930 342.150 ;
        RECT 90.480 341.600 90.630 349.800 ;
        RECT 91.080 341.600 91.230 349.800 ;
        RECT 91.680 341.600 91.830 349.800 ;
        RECT 92.280 341.600 92.430 349.800 ;
        RECT 92.880 341.600 93.030 349.800 ;
        RECT 93.480 341.600 93.630 349.800 ;
        RECT 94.080 341.600 94.230 349.800 ;
        RECT 95.230 350.200 95.380 358.400 ;
        RECT 95.830 350.200 95.980 358.400 ;
        RECT 96.430 350.200 96.580 358.400 ;
        RECT 97.030 350.200 97.180 358.400 ;
        RECT 97.630 350.200 97.780 358.400 ;
        RECT 98.230 350.200 98.380 358.400 ;
        RECT 98.830 350.200 98.980 358.400 ;
        RECT 103.530 357.850 104.730 358.800 ;
        RECT 99.580 357.700 104.730 357.850 ;
        RECT 103.130 357.250 104.730 357.700 ;
        RECT 99.580 357.100 104.730 357.250 ;
        RECT 103.130 356.650 104.730 357.100 ;
        RECT 99.580 356.500 104.730 356.650 ;
        RECT 103.130 356.050 104.730 356.500 ;
        RECT 105.130 356.310 107.130 357.585 ;
        RECT 99.580 355.900 104.730 356.050 ;
        RECT 103.130 355.600 104.730 355.900 ;
        RECT 103.130 355.450 103.530 355.600 ;
        RECT 99.580 355.300 103.530 355.450 ;
        RECT 103.130 354.850 103.530 355.300 ;
        RECT 99.580 354.700 103.530 354.850 ;
        RECT 103.130 354.250 103.530 354.700 ;
        RECT 99.580 354.100 103.530 354.250 ;
        RECT 103.130 353.650 103.530 354.100 ;
        RECT 99.580 353.500 103.530 353.650 ;
        RECT 103.130 353.050 103.530 353.500 ;
        RECT 99.580 352.900 103.530 353.050 ;
        RECT 103.130 352.450 103.530 352.900 ;
        RECT 99.580 352.300 103.530 352.450 ;
        RECT 103.130 351.850 103.530 352.300 ;
        RECT 99.580 351.700 103.530 351.850 ;
        RECT 103.130 351.250 103.530 351.700 ;
        RECT 99.580 351.100 103.530 351.250 ;
        RECT 103.130 350.650 103.530 351.100 ;
        RECT 99.580 350.500 103.530 350.650 ;
        RECT 103.130 350.200 103.530 350.500 ;
        RECT 95.230 349.800 103.530 350.200 ;
        RECT 95.230 341.600 95.380 349.800 ;
        RECT 95.830 341.600 95.980 349.800 ;
        RECT 96.430 341.600 96.580 349.800 ;
        RECT 97.030 341.600 97.180 349.800 ;
        RECT 97.630 341.600 97.780 349.800 ;
        RECT 98.230 341.600 98.380 349.800 ;
        RECT 98.830 341.600 98.980 349.800 ;
        RECT 103.130 349.500 103.530 349.800 ;
        RECT 99.580 349.350 103.530 349.500 ;
        RECT 103.130 348.900 103.530 349.350 ;
        RECT 99.580 348.750 103.530 348.900 ;
        RECT 103.130 348.300 103.530 348.750 ;
        RECT 99.580 348.150 103.530 348.300 ;
        RECT 103.130 347.700 103.530 348.150 ;
        RECT 99.580 347.550 103.530 347.700 ;
        RECT 103.130 347.100 103.530 347.550 ;
        RECT 99.580 346.950 103.530 347.100 ;
        RECT 103.130 346.500 103.530 346.950 ;
        RECT 99.580 346.350 103.530 346.500 ;
        RECT 103.130 345.900 103.530 346.350 ;
        RECT 99.580 345.750 103.530 345.900 ;
        RECT 103.130 345.300 103.530 345.750 ;
        RECT 99.580 345.150 103.530 345.300 ;
        RECT 103.130 344.700 103.530 345.150 ;
        RECT 99.580 344.550 103.530 344.700 ;
        RECT 103.130 344.400 103.530 344.550 ;
        RECT 103.130 344.100 104.730 344.400 ;
        RECT 99.580 343.950 104.730 344.100 ;
        RECT 103.130 343.500 104.730 343.950 ;
        RECT 99.580 343.350 104.730 343.500 ;
        RECT 103.130 342.900 104.730 343.350 ;
        RECT 99.580 342.750 104.730 342.900 ;
        RECT 103.130 342.300 104.730 342.750 ;
        RECT 105.140 342.325 107.140 343.600 ;
        RECT 99.580 342.150 104.730 342.300 ;
        RECT 103.530 341.200 104.730 342.150 ;
        RECT 4.730 338.800 9.130 341.200 ;
        RECT 20.330 338.800 29.130 341.200 ;
        RECT 40.330 338.800 49.130 341.200 ;
        RECT 60.330 338.800 69.130 341.200 ;
        RECT 80.330 338.800 89.130 341.200 ;
        RECT 100.330 338.800 104.730 341.200 ;
        RECT 4.730 337.850 5.940 338.800 ;
        RECT 4.730 337.700 9.880 337.850 ;
        RECT 2.315 336.100 4.320 337.375 ;
        RECT 4.730 337.250 6.330 337.700 ;
        RECT 4.730 337.100 9.880 337.250 ;
        RECT 4.730 336.650 6.330 337.100 ;
        RECT 4.730 336.500 9.880 336.650 ;
        RECT 4.730 336.050 6.330 336.500 ;
        RECT 4.730 335.900 9.880 336.050 ;
        RECT 4.730 335.600 6.330 335.900 ;
        RECT 2.315 333.250 4.315 335.545 ;
        RECT 5.930 335.450 6.330 335.600 ;
        RECT 5.930 335.300 9.880 335.450 ;
        RECT 5.930 334.850 6.330 335.300 ;
        RECT 5.930 334.700 9.880 334.850 ;
        RECT 5.930 334.250 6.330 334.700 ;
        RECT 5.930 334.100 9.880 334.250 ;
        RECT 5.930 333.650 6.330 334.100 ;
        RECT 5.930 333.500 9.880 333.650 ;
        RECT 5.930 333.050 6.330 333.500 ;
        RECT 5.930 332.900 9.880 333.050 ;
        RECT 5.930 332.450 6.330 332.900 ;
        RECT 5.930 332.300 9.880 332.450 ;
        RECT 5.930 331.850 6.330 332.300 ;
        RECT 5.930 331.700 9.880 331.850 ;
        RECT 5.930 331.250 6.330 331.700 ;
        RECT 5.930 331.100 9.880 331.250 ;
        RECT 5.930 330.650 6.330 331.100 ;
        RECT 5.930 330.500 9.880 330.650 ;
        RECT 5.930 330.200 6.330 330.500 ;
        RECT 10.480 330.200 10.630 338.400 ;
        RECT 11.080 330.200 11.230 338.400 ;
        RECT 11.680 330.200 11.830 338.400 ;
        RECT 12.280 330.200 12.430 338.400 ;
        RECT 12.880 330.200 13.030 338.400 ;
        RECT 13.480 330.200 13.630 338.400 ;
        RECT 14.080 330.200 14.230 338.400 ;
        RECT 5.930 329.800 14.230 330.200 ;
        RECT 5.930 329.500 6.330 329.800 ;
        RECT 5.930 329.350 9.880 329.500 ;
        RECT 5.930 328.900 6.330 329.350 ;
        RECT 5.930 328.750 9.880 328.900 ;
        RECT 5.930 328.300 6.330 328.750 ;
        RECT 5.930 328.150 9.880 328.300 ;
        RECT 5.930 327.700 6.330 328.150 ;
        RECT 5.930 327.550 9.880 327.700 ;
        RECT 5.930 327.100 6.330 327.550 ;
        RECT 5.930 326.950 9.880 327.100 ;
        RECT 2.315 324.455 4.315 326.750 ;
        RECT 5.930 326.500 6.330 326.950 ;
        RECT 5.930 326.350 9.880 326.500 ;
        RECT 5.930 325.900 6.330 326.350 ;
        RECT 5.930 325.750 9.880 325.900 ;
        RECT 5.930 325.300 6.330 325.750 ;
        RECT 5.930 325.150 9.880 325.300 ;
        RECT 5.930 324.700 6.330 325.150 ;
        RECT 5.930 324.550 9.880 324.700 ;
        RECT 5.930 324.400 6.330 324.550 ;
        RECT 4.730 324.100 6.330 324.400 ;
        RECT 4.730 323.950 9.880 324.100 ;
        RECT 2.315 322.400 4.320 323.675 ;
        RECT 4.730 323.500 6.330 323.950 ;
        RECT 4.730 323.350 9.880 323.500 ;
        RECT 4.730 322.900 6.330 323.350 ;
        RECT 4.730 322.750 9.880 322.900 ;
        RECT 4.730 322.300 6.330 322.750 ;
        RECT 4.730 322.150 9.880 322.300 ;
        RECT 4.730 321.200 5.930 322.150 ;
        RECT 10.480 321.600 10.630 329.800 ;
        RECT 11.080 321.600 11.230 329.800 ;
        RECT 11.680 321.600 11.830 329.800 ;
        RECT 12.280 321.600 12.430 329.800 ;
        RECT 12.880 321.600 13.030 329.800 ;
        RECT 13.480 321.600 13.630 329.800 ;
        RECT 14.080 321.600 14.230 329.800 ;
        RECT 15.230 330.200 15.380 338.400 ;
        RECT 15.830 330.200 15.980 338.400 ;
        RECT 16.430 330.200 16.580 338.400 ;
        RECT 17.030 330.200 17.180 338.400 ;
        RECT 17.630 330.200 17.780 338.400 ;
        RECT 18.230 330.200 18.380 338.400 ;
        RECT 18.830 330.200 18.980 338.400 ;
        RECT 23.530 337.850 25.940 338.800 ;
        RECT 19.580 337.700 29.880 337.850 ;
        RECT 23.130 337.250 26.330 337.700 ;
        RECT 19.580 337.100 29.880 337.250 ;
        RECT 23.130 336.650 26.330 337.100 ;
        RECT 19.580 336.500 29.880 336.650 ;
        RECT 23.130 336.050 26.330 336.500 ;
        RECT 19.580 335.900 29.880 336.050 ;
        RECT 23.130 335.600 26.330 335.900 ;
        RECT 23.130 335.450 23.530 335.600 ;
        RECT 19.580 335.300 23.530 335.450 ;
        RECT 23.130 334.850 23.530 335.300 ;
        RECT 19.580 334.700 23.530 334.850 ;
        RECT 23.130 334.250 23.530 334.700 ;
        RECT 19.580 334.100 23.530 334.250 ;
        RECT 23.130 333.650 23.530 334.100 ;
        RECT 19.580 333.500 23.530 333.650 ;
        RECT 23.130 333.050 23.530 333.500 ;
        RECT 19.580 332.900 23.530 333.050 ;
        RECT 23.130 332.450 23.530 332.900 ;
        RECT 19.580 332.300 23.530 332.450 ;
        RECT 23.130 331.850 23.530 332.300 ;
        RECT 19.580 331.700 23.530 331.850 ;
        RECT 23.130 331.250 23.530 331.700 ;
        RECT 19.580 331.100 23.530 331.250 ;
        RECT 23.130 330.650 23.530 331.100 ;
        RECT 19.580 330.500 23.530 330.650 ;
        RECT 23.130 330.200 23.530 330.500 ;
        RECT 15.230 329.800 23.530 330.200 ;
        RECT 15.230 321.600 15.380 329.800 ;
        RECT 15.830 321.600 15.980 329.800 ;
        RECT 16.430 321.600 16.580 329.800 ;
        RECT 17.030 321.600 17.180 329.800 ;
        RECT 17.630 321.600 17.780 329.800 ;
        RECT 18.230 321.600 18.380 329.800 ;
        RECT 18.830 321.600 18.980 329.800 ;
        RECT 23.130 329.500 23.530 329.800 ;
        RECT 19.580 329.350 23.530 329.500 ;
        RECT 23.130 328.900 23.530 329.350 ;
        RECT 19.580 328.750 23.530 328.900 ;
        RECT 23.130 328.300 23.530 328.750 ;
        RECT 19.580 328.150 23.530 328.300 ;
        RECT 23.130 327.700 23.530 328.150 ;
        RECT 19.580 327.550 23.530 327.700 ;
        RECT 23.130 327.100 23.530 327.550 ;
        RECT 19.580 326.950 23.530 327.100 ;
        RECT 23.130 326.500 23.530 326.950 ;
        RECT 19.580 326.350 23.530 326.500 ;
        RECT 23.130 325.900 23.530 326.350 ;
        RECT 19.580 325.750 23.530 325.900 ;
        RECT 23.130 325.300 23.530 325.750 ;
        RECT 19.580 325.150 23.530 325.300 ;
        RECT 23.130 324.700 23.530 325.150 ;
        RECT 19.580 324.550 23.530 324.700 ;
        RECT 23.130 324.400 23.530 324.550 ;
        RECT 25.930 335.450 26.330 335.600 ;
        RECT 25.930 335.300 29.880 335.450 ;
        RECT 25.930 334.850 26.330 335.300 ;
        RECT 25.930 334.700 29.880 334.850 ;
        RECT 25.930 334.250 26.330 334.700 ;
        RECT 25.930 334.100 29.880 334.250 ;
        RECT 25.930 333.650 26.330 334.100 ;
        RECT 25.930 333.500 29.880 333.650 ;
        RECT 25.930 333.050 26.330 333.500 ;
        RECT 25.930 332.900 29.880 333.050 ;
        RECT 25.930 332.450 26.330 332.900 ;
        RECT 25.930 332.300 29.880 332.450 ;
        RECT 25.930 331.850 26.330 332.300 ;
        RECT 25.930 331.700 29.880 331.850 ;
        RECT 25.930 331.250 26.330 331.700 ;
        RECT 25.930 331.100 29.880 331.250 ;
        RECT 25.930 330.650 26.330 331.100 ;
        RECT 25.930 330.500 29.880 330.650 ;
        RECT 25.930 330.200 26.330 330.500 ;
        RECT 30.480 330.200 30.630 338.400 ;
        RECT 31.080 330.200 31.230 338.400 ;
        RECT 31.680 330.200 31.830 338.400 ;
        RECT 32.280 330.200 32.430 338.400 ;
        RECT 32.880 330.200 33.030 338.400 ;
        RECT 33.480 330.200 33.630 338.400 ;
        RECT 34.080 330.200 34.230 338.400 ;
        RECT 25.930 329.800 34.230 330.200 ;
        RECT 25.930 329.500 26.330 329.800 ;
        RECT 25.930 329.350 29.880 329.500 ;
        RECT 25.930 328.900 26.330 329.350 ;
        RECT 25.930 328.750 29.880 328.900 ;
        RECT 25.930 328.300 26.330 328.750 ;
        RECT 25.930 328.150 29.880 328.300 ;
        RECT 25.930 327.700 26.330 328.150 ;
        RECT 25.930 327.550 29.880 327.700 ;
        RECT 25.930 327.100 26.330 327.550 ;
        RECT 25.930 326.950 29.880 327.100 ;
        RECT 25.930 326.500 26.330 326.950 ;
        RECT 25.930 326.350 29.880 326.500 ;
        RECT 25.930 325.900 26.330 326.350 ;
        RECT 25.930 325.750 29.880 325.900 ;
        RECT 25.930 325.300 26.330 325.750 ;
        RECT 25.930 325.150 29.880 325.300 ;
        RECT 25.930 324.700 26.330 325.150 ;
        RECT 25.930 324.550 29.880 324.700 ;
        RECT 25.930 324.400 26.330 324.550 ;
        RECT 23.130 324.100 26.330 324.400 ;
        RECT 19.580 323.950 29.880 324.100 ;
        RECT 23.130 323.500 26.330 323.950 ;
        RECT 19.580 323.350 29.880 323.500 ;
        RECT 23.130 322.900 26.330 323.350 ;
        RECT 19.580 322.750 29.880 322.900 ;
        RECT 23.130 322.300 26.330 322.750 ;
        RECT 19.580 322.150 29.880 322.300 ;
        RECT 23.530 321.200 25.930 322.150 ;
        RECT 30.480 321.600 30.630 329.800 ;
        RECT 31.080 321.600 31.230 329.800 ;
        RECT 31.680 321.600 31.830 329.800 ;
        RECT 32.280 321.600 32.430 329.800 ;
        RECT 32.880 321.600 33.030 329.800 ;
        RECT 33.480 321.600 33.630 329.800 ;
        RECT 34.080 321.600 34.230 329.800 ;
        RECT 35.230 330.200 35.380 338.400 ;
        RECT 35.830 330.200 35.980 338.400 ;
        RECT 36.430 330.200 36.580 338.400 ;
        RECT 37.030 330.200 37.180 338.400 ;
        RECT 37.630 330.200 37.780 338.400 ;
        RECT 38.230 330.200 38.380 338.400 ;
        RECT 38.830 330.200 38.980 338.400 ;
        RECT 43.530 337.850 45.940 338.800 ;
        RECT 39.580 337.700 49.880 337.850 ;
        RECT 43.130 337.250 46.330 337.700 ;
        RECT 39.580 337.100 49.880 337.250 ;
        RECT 43.130 336.650 46.330 337.100 ;
        RECT 39.580 336.500 49.880 336.650 ;
        RECT 43.130 336.050 46.330 336.500 ;
        RECT 39.580 335.900 49.880 336.050 ;
        RECT 43.130 335.600 46.330 335.900 ;
        RECT 43.130 335.450 43.530 335.600 ;
        RECT 39.580 335.300 43.530 335.450 ;
        RECT 43.130 334.850 43.530 335.300 ;
        RECT 39.580 334.700 43.530 334.850 ;
        RECT 43.130 334.250 43.530 334.700 ;
        RECT 39.580 334.100 43.530 334.250 ;
        RECT 43.130 333.650 43.530 334.100 ;
        RECT 39.580 333.500 43.530 333.650 ;
        RECT 43.130 333.050 43.530 333.500 ;
        RECT 39.580 332.900 43.530 333.050 ;
        RECT 43.130 332.450 43.530 332.900 ;
        RECT 39.580 332.300 43.530 332.450 ;
        RECT 43.130 331.850 43.530 332.300 ;
        RECT 39.580 331.700 43.530 331.850 ;
        RECT 43.130 331.250 43.530 331.700 ;
        RECT 39.580 331.100 43.530 331.250 ;
        RECT 43.130 330.650 43.530 331.100 ;
        RECT 39.580 330.500 43.530 330.650 ;
        RECT 43.130 330.200 43.530 330.500 ;
        RECT 35.230 329.800 43.530 330.200 ;
        RECT 35.230 321.600 35.380 329.800 ;
        RECT 35.830 321.600 35.980 329.800 ;
        RECT 36.430 321.600 36.580 329.800 ;
        RECT 37.030 321.600 37.180 329.800 ;
        RECT 37.630 321.600 37.780 329.800 ;
        RECT 38.230 321.600 38.380 329.800 ;
        RECT 38.830 321.600 38.980 329.800 ;
        RECT 43.130 329.500 43.530 329.800 ;
        RECT 39.580 329.350 43.530 329.500 ;
        RECT 43.130 328.900 43.530 329.350 ;
        RECT 39.580 328.750 43.530 328.900 ;
        RECT 43.130 328.300 43.530 328.750 ;
        RECT 39.580 328.150 43.530 328.300 ;
        RECT 43.130 327.700 43.530 328.150 ;
        RECT 39.580 327.550 43.530 327.700 ;
        RECT 43.130 327.100 43.530 327.550 ;
        RECT 39.580 326.950 43.530 327.100 ;
        RECT 43.130 326.500 43.530 326.950 ;
        RECT 39.580 326.350 43.530 326.500 ;
        RECT 43.130 325.900 43.530 326.350 ;
        RECT 39.580 325.750 43.530 325.900 ;
        RECT 43.130 325.300 43.530 325.750 ;
        RECT 39.580 325.150 43.530 325.300 ;
        RECT 43.130 324.700 43.530 325.150 ;
        RECT 39.580 324.550 43.530 324.700 ;
        RECT 43.130 324.400 43.530 324.550 ;
        RECT 45.930 335.450 46.330 335.600 ;
        RECT 45.930 335.300 49.880 335.450 ;
        RECT 45.930 334.850 46.330 335.300 ;
        RECT 45.930 334.700 49.880 334.850 ;
        RECT 45.930 334.250 46.330 334.700 ;
        RECT 45.930 334.100 49.880 334.250 ;
        RECT 45.930 333.650 46.330 334.100 ;
        RECT 45.930 333.500 49.880 333.650 ;
        RECT 45.930 333.050 46.330 333.500 ;
        RECT 45.930 332.900 49.880 333.050 ;
        RECT 45.930 332.450 46.330 332.900 ;
        RECT 45.930 332.300 49.880 332.450 ;
        RECT 45.930 331.850 46.330 332.300 ;
        RECT 45.930 331.700 49.880 331.850 ;
        RECT 45.930 331.250 46.330 331.700 ;
        RECT 45.930 331.100 49.880 331.250 ;
        RECT 45.930 330.650 46.330 331.100 ;
        RECT 45.930 330.500 49.880 330.650 ;
        RECT 45.930 330.200 46.330 330.500 ;
        RECT 50.480 330.200 50.630 338.400 ;
        RECT 51.080 330.200 51.230 338.400 ;
        RECT 51.680 330.200 51.830 338.400 ;
        RECT 52.280 330.200 52.430 338.400 ;
        RECT 52.880 330.200 53.030 338.400 ;
        RECT 53.480 330.200 53.630 338.400 ;
        RECT 54.080 330.200 54.230 338.400 ;
        RECT 45.930 329.800 54.230 330.200 ;
        RECT 45.930 329.500 46.330 329.800 ;
        RECT 45.930 329.350 49.880 329.500 ;
        RECT 45.930 328.900 46.330 329.350 ;
        RECT 45.930 328.750 49.880 328.900 ;
        RECT 45.930 328.300 46.330 328.750 ;
        RECT 45.930 328.150 49.880 328.300 ;
        RECT 45.930 327.700 46.330 328.150 ;
        RECT 45.930 327.550 49.880 327.700 ;
        RECT 45.930 327.100 46.330 327.550 ;
        RECT 45.930 326.950 49.880 327.100 ;
        RECT 45.930 326.500 46.330 326.950 ;
        RECT 45.930 326.350 49.880 326.500 ;
        RECT 45.930 325.900 46.330 326.350 ;
        RECT 45.930 325.750 49.880 325.900 ;
        RECT 45.930 325.300 46.330 325.750 ;
        RECT 45.930 325.150 49.880 325.300 ;
        RECT 45.930 324.700 46.330 325.150 ;
        RECT 45.930 324.550 49.880 324.700 ;
        RECT 45.930 324.400 46.330 324.550 ;
        RECT 43.130 324.100 46.330 324.400 ;
        RECT 39.580 323.950 49.880 324.100 ;
        RECT 43.130 323.500 46.330 323.950 ;
        RECT 39.580 323.350 49.880 323.500 ;
        RECT 43.130 322.900 46.330 323.350 ;
        RECT 39.580 322.750 49.880 322.900 ;
        RECT 43.130 322.300 46.330 322.750 ;
        RECT 39.580 322.150 49.880 322.300 ;
        RECT 43.530 321.200 45.930 322.150 ;
        RECT 50.480 321.600 50.630 329.800 ;
        RECT 51.080 321.600 51.230 329.800 ;
        RECT 51.680 321.600 51.830 329.800 ;
        RECT 52.280 321.600 52.430 329.800 ;
        RECT 52.880 321.600 53.030 329.800 ;
        RECT 53.480 321.600 53.630 329.800 ;
        RECT 54.080 321.600 54.230 329.800 ;
        RECT 55.230 330.200 55.380 338.400 ;
        RECT 55.830 330.200 55.980 338.400 ;
        RECT 56.430 330.200 56.580 338.400 ;
        RECT 57.030 330.200 57.180 338.400 ;
        RECT 57.630 330.200 57.780 338.400 ;
        RECT 58.230 330.200 58.380 338.400 ;
        RECT 58.830 330.200 58.980 338.400 ;
        RECT 63.530 337.850 65.940 338.800 ;
        RECT 59.580 337.700 69.880 337.850 ;
        RECT 63.130 337.250 66.330 337.700 ;
        RECT 59.580 337.100 69.880 337.250 ;
        RECT 63.130 336.650 66.330 337.100 ;
        RECT 59.580 336.500 69.880 336.650 ;
        RECT 63.130 336.050 66.330 336.500 ;
        RECT 59.580 335.900 69.880 336.050 ;
        RECT 63.130 335.600 66.330 335.900 ;
        RECT 63.130 335.450 63.530 335.600 ;
        RECT 59.580 335.300 63.530 335.450 ;
        RECT 63.130 334.850 63.530 335.300 ;
        RECT 59.580 334.700 63.530 334.850 ;
        RECT 63.130 334.250 63.530 334.700 ;
        RECT 59.580 334.100 63.530 334.250 ;
        RECT 63.130 333.650 63.530 334.100 ;
        RECT 59.580 333.500 63.530 333.650 ;
        RECT 63.130 333.050 63.530 333.500 ;
        RECT 59.580 332.900 63.530 333.050 ;
        RECT 63.130 332.450 63.530 332.900 ;
        RECT 59.580 332.300 63.530 332.450 ;
        RECT 63.130 331.850 63.530 332.300 ;
        RECT 59.580 331.700 63.530 331.850 ;
        RECT 63.130 331.250 63.530 331.700 ;
        RECT 59.580 331.100 63.530 331.250 ;
        RECT 63.130 330.650 63.530 331.100 ;
        RECT 59.580 330.500 63.530 330.650 ;
        RECT 63.130 330.200 63.530 330.500 ;
        RECT 55.230 329.800 63.530 330.200 ;
        RECT 55.230 321.600 55.380 329.800 ;
        RECT 55.830 321.600 55.980 329.800 ;
        RECT 56.430 321.600 56.580 329.800 ;
        RECT 57.030 321.600 57.180 329.800 ;
        RECT 57.630 321.600 57.780 329.800 ;
        RECT 58.230 321.600 58.380 329.800 ;
        RECT 58.830 321.600 58.980 329.800 ;
        RECT 63.130 329.500 63.530 329.800 ;
        RECT 59.580 329.350 63.530 329.500 ;
        RECT 63.130 328.900 63.530 329.350 ;
        RECT 59.580 328.750 63.530 328.900 ;
        RECT 63.130 328.300 63.530 328.750 ;
        RECT 59.580 328.150 63.530 328.300 ;
        RECT 63.130 327.700 63.530 328.150 ;
        RECT 59.580 327.550 63.530 327.700 ;
        RECT 63.130 327.100 63.530 327.550 ;
        RECT 59.580 326.950 63.530 327.100 ;
        RECT 63.130 326.500 63.530 326.950 ;
        RECT 59.580 326.350 63.530 326.500 ;
        RECT 63.130 325.900 63.530 326.350 ;
        RECT 59.580 325.750 63.530 325.900 ;
        RECT 63.130 325.300 63.530 325.750 ;
        RECT 59.580 325.150 63.530 325.300 ;
        RECT 63.130 324.700 63.530 325.150 ;
        RECT 59.580 324.550 63.530 324.700 ;
        RECT 63.130 324.400 63.530 324.550 ;
        RECT 65.930 335.450 66.330 335.600 ;
        RECT 65.930 335.300 69.880 335.450 ;
        RECT 65.930 334.850 66.330 335.300 ;
        RECT 65.930 334.700 69.880 334.850 ;
        RECT 65.930 334.250 66.330 334.700 ;
        RECT 65.930 334.100 69.880 334.250 ;
        RECT 65.930 333.650 66.330 334.100 ;
        RECT 65.930 333.500 69.880 333.650 ;
        RECT 65.930 333.050 66.330 333.500 ;
        RECT 65.930 332.900 69.880 333.050 ;
        RECT 65.930 332.450 66.330 332.900 ;
        RECT 65.930 332.300 69.880 332.450 ;
        RECT 65.930 331.850 66.330 332.300 ;
        RECT 65.930 331.700 69.880 331.850 ;
        RECT 65.930 331.250 66.330 331.700 ;
        RECT 65.930 331.100 69.880 331.250 ;
        RECT 65.930 330.650 66.330 331.100 ;
        RECT 65.930 330.500 69.880 330.650 ;
        RECT 65.930 330.200 66.330 330.500 ;
        RECT 70.480 330.200 70.630 338.400 ;
        RECT 71.080 330.200 71.230 338.400 ;
        RECT 71.680 330.200 71.830 338.400 ;
        RECT 72.280 330.200 72.430 338.400 ;
        RECT 72.880 330.200 73.030 338.400 ;
        RECT 73.480 330.200 73.630 338.400 ;
        RECT 74.080 330.200 74.230 338.400 ;
        RECT 65.930 329.800 74.230 330.200 ;
        RECT 65.930 329.500 66.330 329.800 ;
        RECT 65.930 329.350 69.880 329.500 ;
        RECT 65.930 328.900 66.330 329.350 ;
        RECT 65.930 328.750 69.880 328.900 ;
        RECT 65.930 328.300 66.330 328.750 ;
        RECT 65.930 328.150 69.880 328.300 ;
        RECT 65.930 327.700 66.330 328.150 ;
        RECT 65.930 327.550 69.880 327.700 ;
        RECT 65.930 327.100 66.330 327.550 ;
        RECT 65.930 326.950 69.880 327.100 ;
        RECT 65.930 326.500 66.330 326.950 ;
        RECT 65.930 326.350 69.880 326.500 ;
        RECT 65.930 325.900 66.330 326.350 ;
        RECT 65.930 325.750 69.880 325.900 ;
        RECT 65.930 325.300 66.330 325.750 ;
        RECT 65.930 325.150 69.880 325.300 ;
        RECT 65.930 324.700 66.330 325.150 ;
        RECT 65.930 324.550 69.880 324.700 ;
        RECT 65.930 324.400 66.330 324.550 ;
        RECT 63.130 324.100 66.330 324.400 ;
        RECT 59.580 323.950 69.880 324.100 ;
        RECT 63.130 323.500 66.330 323.950 ;
        RECT 59.580 323.350 69.880 323.500 ;
        RECT 63.130 322.900 66.330 323.350 ;
        RECT 59.580 322.750 69.880 322.900 ;
        RECT 63.130 322.300 66.330 322.750 ;
        RECT 59.580 322.150 69.880 322.300 ;
        RECT 63.530 321.200 65.930 322.150 ;
        RECT 70.480 321.600 70.630 329.800 ;
        RECT 71.080 321.600 71.230 329.800 ;
        RECT 71.680 321.600 71.830 329.800 ;
        RECT 72.280 321.600 72.430 329.800 ;
        RECT 72.880 321.600 73.030 329.800 ;
        RECT 73.480 321.600 73.630 329.800 ;
        RECT 74.080 321.600 74.230 329.800 ;
        RECT 75.230 330.200 75.380 338.400 ;
        RECT 75.830 330.200 75.980 338.400 ;
        RECT 76.430 330.200 76.580 338.400 ;
        RECT 77.030 330.200 77.180 338.400 ;
        RECT 77.630 330.200 77.780 338.400 ;
        RECT 78.230 330.200 78.380 338.400 ;
        RECT 78.830 330.200 78.980 338.400 ;
        RECT 83.530 337.850 85.940 338.800 ;
        RECT 79.580 337.700 89.880 337.850 ;
        RECT 83.130 337.250 86.330 337.700 ;
        RECT 79.580 337.100 89.880 337.250 ;
        RECT 83.130 336.650 86.330 337.100 ;
        RECT 79.580 336.500 89.880 336.650 ;
        RECT 83.130 336.050 86.330 336.500 ;
        RECT 79.580 335.900 89.880 336.050 ;
        RECT 83.130 335.600 86.330 335.900 ;
        RECT 83.130 335.450 83.530 335.600 ;
        RECT 79.580 335.300 83.530 335.450 ;
        RECT 83.130 334.850 83.530 335.300 ;
        RECT 79.580 334.700 83.530 334.850 ;
        RECT 83.130 334.250 83.530 334.700 ;
        RECT 79.580 334.100 83.530 334.250 ;
        RECT 83.130 333.650 83.530 334.100 ;
        RECT 79.580 333.500 83.530 333.650 ;
        RECT 83.130 333.050 83.530 333.500 ;
        RECT 79.580 332.900 83.530 333.050 ;
        RECT 83.130 332.450 83.530 332.900 ;
        RECT 79.580 332.300 83.530 332.450 ;
        RECT 83.130 331.850 83.530 332.300 ;
        RECT 79.580 331.700 83.530 331.850 ;
        RECT 83.130 331.250 83.530 331.700 ;
        RECT 79.580 331.100 83.530 331.250 ;
        RECT 83.130 330.650 83.530 331.100 ;
        RECT 79.580 330.500 83.530 330.650 ;
        RECT 83.130 330.200 83.530 330.500 ;
        RECT 75.230 329.800 83.530 330.200 ;
        RECT 75.230 321.600 75.380 329.800 ;
        RECT 75.830 321.600 75.980 329.800 ;
        RECT 76.430 321.600 76.580 329.800 ;
        RECT 77.030 321.600 77.180 329.800 ;
        RECT 77.630 321.600 77.780 329.800 ;
        RECT 78.230 321.600 78.380 329.800 ;
        RECT 78.830 321.600 78.980 329.800 ;
        RECT 83.130 329.500 83.530 329.800 ;
        RECT 79.580 329.350 83.530 329.500 ;
        RECT 83.130 328.900 83.530 329.350 ;
        RECT 79.580 328.750 83.530 328.900 ;
        RECT 83.130 328.300 83.530 328.750 ;
        RECT 79.580 328.150 83.530 328.300 ;
        RECT 83.130 327.700 83.530 328.150 ;
        RECT 79.580 327.550 83.530 327.700 ;
        RECT 83.130 327.100 83.530 327.550 ;
        RECT 79.580 326.950 83.530 327.100 ;
        RECT 83.130 326.500 83.530 326.950 ;
        RECT 79.580 326.350 83.530 326.500 ;
        RECT 83.130 325.900 83.530 326.350 ;
        RECT 79.580 325.750 83.530 325.900 ;
        RECT 83.130 325.300 83.530 325.750 ;
        RECT 79.580 325.150 83.530 325.300 ;
        RECT 83.130 324.700 83.530 325.150 ;
        RECT 79.580 324.550 83.530 324.700 ;
        RECT 83.130 324.400 83.530 324.550 ;
        RECT 85.930 335.450 86.330 335.600 ;
        RECT 85.930 335.300 89.880 335.450 ;
        RECT 85.930 334.850 86.330 335.300 ;
        RECT 85.930 334.700 89.880 334.850 ;
        RECT 85.930 334.250 86.330 334.700 ;
        RECT 85.930 334.100 89.880 334.250 ;
        RECT 85.930 333.650 86.330 334.100 ;
        RECT 85.930 333.500 89.880 333.650 ;
        RECT 85.930 333.050 86.330 333.500 ;
        RECT 85.930 332.900 89.880 333.050 ;
        RECT 85.930 332.450 86.330 332.900 ;
        RECT 85.930 332.300 89.880 332.450 ;
        RECT 85.930 331.850 86.330 332.300 ;
        RECT 85.930 331.700 89.880 331.850 ;
        RECT 85.930 331.250 86.330 331.700 ;
        RECT 85.930 331.100 89.880 331.250 ;
        RECT 85.930 330.650 86.330 331.100 ;
        RECT 85.930 330.500 89.880 330.650 ;
        RECT 85.930 330.200 86.330 330.500 ;
        RECT 90.480 330.200 90.630 338.400 ;
        RECT 91.080 330.200 91.230 338.400 ;
        RECT 91.680 330.200 91.830 338.400 ;
        RECT 92.280 330.200 92.430 338.400 ;
        RECT 92.880 330.200 93.030 338.400 ;
        RECT 93.480 330.200 93.630 338.400 ;
        RECT 94.080 330.200 94.230 338.400 ;
        RECT 85.930 329.800 94.230 330.200 ;
        RECT 85.930 329.500 86.330 329.800 ;
        RECT 85.930 329.350 89.880 329.500 ;
        RECT 85.930 328.900 86.330 329.350 ;
        RECT 85.930 328.750 89.880 328.900 ;
        RECT 85.930 328.300 86.330 328.750 ;
        RECT 85.930 328.150 89.880 328.300 ;
        RECT 85.930 327.700 86.330 328.150 ;
        RECT 85.930 327.550 89.880 327.700 ;
        RECT 85.930 327.100 86.330 327.550 ;
        RECT 85.930 326.950 89.880 327.100 ;
        RECT 85.930 326.500 86.330 326.950 ;
        RECT 85.930 326.350 89.880 326.500 ;
        RECT 85.930 325.900 86.330 326.350 ;
        RECT 85.930 325.750 89.880 325.900 ;
        RECT 85.930 325.300 86.330 325.750 ;
        RECT 85.930 325.150 89.880 325.300 ;
        RECT 85.930 324.700 86.330 325.150 ;
        RECT 85.930 324.550 89.880 324.700 ;
        RECT 85.930 324.400 86.330 324.550 ;
        RECT 83.130 324.100 86.330 324.400 ;
        RECT 79.580 323.950 89.880 324.100 ;
        RECT 83.130 323.500 86.330 323.950 ;
        RECT 79.580 323.350 89.880 323.500 ;
        RECT 83.130 322.900 86.330 323.350 ;
        RECT 79.580 322.750 89.880 322.900 ;
        RECT 83.130 322.300 86.330 322.750 ;
        RECT 79.580 322.150 89.880 322.300 ;
        RECT 83.530 321.200 85.930 322.150 ;
        RECT 90.480 321.600 90.630 329.800 ;
        RECT 91.080 321.600 91.230 329.800 ;
        RECT 91.680 321.600 91.830 329.800 ;
        RECT 92.280 321.600 92.430 329.800 ;
        RECT 92.880 321.600 93.030 329.800 ;
        RECT 93.480 321.600 93.630 329.800 ;
        RECT 94.080 321.600 94.230 329.800 ;
        RECT 95.230 330.200 95.380 338.400 ;
        RECT 95.830 330.200 95.980 338.400 ;
        RECT 96.430 330.200 96.580 338.400 ;
        RECT 97.030 330.200 97.180 338.400 ;
        RECT 97.630 330.200 97.780 338.400 ;
        RECT 98.230 330.200 98.380 338.400 ;
        RECT 98.830 330.200 98.980 338.400 ;
        RECT 103.530 337.850 104.730 338.800 ;
        RECT 99.580 337.700 104.730 337.850 ;
        RECT 103.130 337.250 104.730 337.700 ;
        RECT 99.580 337.100 104.730 337.250 ;
        RECT 103.130 336.650 104.730 337.100 ;
        RECT 99.580 336.500 104.730 336.650 ;
        RECT 103.130 336.050 104.730 336.500 ;
        RECT 105.130 336.310 107.130 337.585 ;
        RECT 99.580 335.900 104.730 336.050 ;
        RECT 103.130 335.600 104.730 335.900 ;
        RECT 103.130 335.450 103.530 335.600 ;
        RECT 99.580 335.300 103.530 335.450 ;
        RECT 103.130 334.850 103.530 335.300 ;
        RECT 99.580 334.700 103.530 334.850 ;
        RECT 103.130 334.250 103.530 334.700 ;
        RECT 99.580 334.100 103.530 334.250 ;
        RECT 103.130 333.650 103.530 334.100 ;
        RECT 99.580 333.500 103.530 333.650 ;
        RECT 103.130 333.050 103.530 333.500 ;
        RECT 99.580 332.900 103.530 333.050 ;
        RECT 103.130 332.450 103.530 332.900 ;
        RECT 99.580 332.300 103.530 332.450 ;
        RECT 103.130 331.850 103.530 332.300 ;
        RECT 99.580 331.700 103.530 331.850 ;
        RECT 103.130 331.250 103.530 331.700 ;
        RECT 99.580 331.100 103.530 331.250 ;
        RECT 103.130 330.650 103.530 331.100 ;
        RECT 99.580 330.500 103.530 330.650 ;
        RECT 103.130 330.200 103.530 330.500 ;
        RECT 95.230 329.800 103.530 330.200 ;
        RECT 95.230 321.600 95.380 329.800 ;
        RECT 95.830 321.600 95.980 329.800 ;
        RECT 96.430 321.600 96.580 329.800 ;
        RECT 97.030 321.600 97.180 329.800 ;
        RECT 97.630 321.600 97.780 329.800 ;
        RECT 98.230 321.600 98.380 329.800 ;
        RECT 98.830 321.600 98.980 329.800 ;
        RECT 103.130 329.500 103.530 329.800 ;
        RECT 99.580 329.350 103.530 329.500 ;
        RECT 103.130 328.900 103.530 329.350 ;
        RECT 99.580 328.750 103.530 328.900 ;
        RECT 103.130 328.300 103.530 328.750 ;
        RECT 99.580 328.150 103.530 328.300 ;
        RECT 103.130 327.700 103.530 328.150 ;
        RECT 99.580 327.550 103.530 327.700 ;
        RECT 103.130 327.100 103.530 327.550 ;
        RECT 99.580 326.950 103.530 327.100 ;
        RECT 103.130 326.500 103.530 326.950 ;
        RECT 99.580 326.350 103.530 326.500 ;
        RECT 103.130 325.900 103.530 326.350 ;
        RECT 99.580 325.750 103.530 325.900 ;
        RECT 103.130 325.300 103.530 325.750 ;
        RECT 99.580 325.150 103.530 325.300 ;
        RECT 103.130 324.700 103.530 325.150 ;
        RECT 99.580 324.550 103.530 324.700 ;
        RECT 103.130 324.400 103.530 324.550 ;
        RECT 103.130 324.100 104.730 324.400 ;
        RECT 99.580 323.950 104.730 324.100 ;
        RECT 103.130 323.500 104.730 323.950 ;
        RECT 99.580 323.350 104.730 323.500 ;
        RECT 103.130 322.900 104.730 323.350 ;
        RECT 99.580 322.750 104.730 322.900 ;
        RECT 103.130 322.300 104.730 322.750 ;
        RECT 105.140 322.325 107.140 323.600 ;
        RECT 99.580 322.150 104.730 322.300 ;
        RECT 103.530 321.200 104.730 322.150 ;
        RECT 4.730 318.800 9.130 321.200 ;
        RECT 20.330 318.800 29.130 321.200 ;
        RECT 40.330 318.800 49.130 321.200 ;
        RECT 60.330 318.800 69.130 321.200 ;
        RECT 80.330 318.800 89.130 321.200 ;
        RECT 100.330 318.800 104.730 321.200 ;
        RECT 4.730 317.850 5.940 318.800 ;
        RECT 2.315 316.510 4.320 317.785 ;
        RECT 4.730 317.700 9.880 317.850 ;
        RECT 4.730 317.250 6.330 317.700 ;
        RECT 4.730 317.100 9.880 317.250 ;
        RECT 4.730 316.650 6.330 317.100 ;
        RECT 4.730 316.500 9.880 316.650 ;
        RECT 4.730 316.050 6.330 316.500 ;
        RECT 4.730 315.900 9.880 316.050 ;
        RECT 4.730 315.600 6.330 315.900 ;
        RECT 2.320 315.340 4.320 315.545 ;
        RECT 2.315 313.250 4.320 315.340 ;
        RECT 5.930 315.450 6.330 315.600 ;
        RECT 5.930 315.300 9.880 315.450 ;
        RECT 5.930 314.850 6.330 315.300 ;
        RECT 5.930 314.700 9.880 314.850 ;
        RECT 5.930 314.250 6.330 314.700 ;
        RECT 5.930 314.100 9.880 314.250 ;
        RECT 5.930 313.650 6.330 314.100 ;
        RECT 5.930 313.500 9.880 313.650 ;
        RECT 5.930 313.050 6.330 313.500 ;
        RECT 5.930 312.900 9.880 313.050 ;
        RECT 5.930 312.450 6.330 312.900 ;
        RECT 5.930 312.300 9.880 312.450 ;
        RECT 5.930 311.850 6.330 312.300 ;
        RECT 5.930 311.700 9.880 311.850 ;
        RECT 5.930 311.250 6.330 311.700 ;
        RECT 5.930 311.100 9.880 311.250 ;
        RECT 5.930 310.650 6.330 311.100 ;
        RECT 5.930 310.500 9.880 310.650 ;
        RECT 5.930 310.200 6.330 310.500 ;
        RECT 10.480 310.200 10.630 318.400 ;
        RECT 11.080 310.200 11.230 318.400 ;
        RECT 11.680 310.200 11.830 318.400 ;
        RECT 12.280 310.200 12.430 318.400 ;
        RECT 12.880 310.200 13.030 318.400 ;
        RECT 13.480 310.200 13.630 318.400 ;
        RECT 14.080 310.200 14.230 318.400 ;
        RECT 5.930 309.800 14.230 310.200 ;
        RECT 5.930 309.500 6.330 309.800 ;
        RECT 5.930 309.350 9.880 309.500 ;
        RECT 5.930 308.900 6.330 309.350 ;
        RECT 5.930 308.750 9.880 308.900 ;
        RECT 5.930 308.300 6.330 308.750 ;
        RECT 5.930 308.150 9.880 308.300 ;
        RECT 5.930 307.700 6.330 308.150 ;
        RECT 5.930 307.550 9.880 307.700 ;
        RECT 5.930 307.100 6.330 307.550 ;
        RECT 5.930 306.950 9.880 307.100 ;
        RECT 2.315 304.455 4.315 306.750 ;
        RECT 5.930 306.500 6.330 306.950 ;
        RECT 5.930 306.350 9.880 306.500 ;
        RECT 5.930 305.900 6.330 306.350 ;
        RECT 5.930 305.750 9.880 305.900 ;
        RECT 5.930 305.300 6.330 305.750 ;
        RECT 5.930 305.150 9.880 305.300 ;
        RECT 5.930 304.700 6.330 305.150 ;
        RECT 5.930 304.550 9.880 304.700 ;
        RECT 5.930 304.400 6.330 304.550 ;
        RECT 4.730 304.100 6.330 304.400 ;
        RECT 4.730 303.950 9.880 304.100 ;
        RECT 2.315 302.270 4.330 303.545 ;
        RECT 4.730 303.500 6.330 303.950 ;
        RECT 4.730 303.350 9.880 303.500 ;
        RECT 4.730 302.900 6.330 303.350 ;
        RECT 4.730 302.750 9.880 302.900 ;
        RECT 4.730 302.300 6.330 302.750 ;
        RECT 4.730 302.150 9.880 302.300 ;
        RECT 4.730 301.200 5.930 302.150 ;
        RECT 10.480 301.600 10.630 309.800 ;
        RECT 11.080 301.600 11.230 309.800 ;
        RECT 11.680 301.600 11.830 309.800 ;
        RECT 12.280 301.600 12.430 309.800 ;
        RECT 12.880 301.600 13.030 309.800 ;
        RECT 13.480 301.600 13.630 309.800 ;
        RECT 14.080 301.600 14.230 309.800 ;
        RECT 15.230 310.200 15.380 318.400 ;
        RECT 15.830 310.200 15.980 318.400 ;
        RECT 16.430 310.200 16.580 318.400 ;
        RECT 17.030 310.200 17.180 318.400 ;
        RECT 17.630 310.200 17.780 318.400 ;
        RECT 18.230 310.200 18.380 318.400 ;
        RECT 18.830 310.200 18.980 318.400 ;
        RECT 23.530 317.850 25.940 318.800 ;
        RECT 19.580 317.700 29.880 317.850 ;
        RECT 23.130 317.250 26.330 317.700 ;
        RECT 19.580 317.100 29.880 317.250 ;
        RECT 23.130 316.650 26.330 317.100 ;
        RECT 19.580 316.500 29.880 316.650 ;
        RECT 23.130 316.050 26.330 316.500 ;
        RECT 19.580 315.900 29.880 316.050 ;
        RECT 23.130 315.600 26.330 315.900 ;
        RECT 23.130 315.450 23.530 315.600 ;
        RECT 19.580 315.300 23.530 315.450 ;
        RECT 23.130 314.850 23.530 315.300 ;
        RECT 19.580 314.700 23.530 314.850 ;
        RECT 23.130 314.250 23.530 314.700 ;
        RECT 19.580 314.100 23.530 314.250 ;
        RECT 23.130 313.650 23.530 314.100 ;
        RECT 19.580 313.500 23.530 313.650 ;
        RECT 23.130 313.050 23.530 313.500 ;
        RECT 19.580 312.900 23.530 313.050 ;
        RECT 23.130 312.450 23.530 312.900 ;
        RECT 19.580 312.300 23.530 312.450 ;
        RECT 23.130 311.850 23.530 312.300 ;
        RECT 19.580 311.700 23.530 311.850 ;
        RECT 23.130 311.250 23.530 311.700 ;
        RECT 19.580 311.100 23.530 311.250 ;
        RECT 23.130 310.650 23.530 311.100 ;
        RECT 19.580 310.500 23.530 310.650 ;
        RECT 23.130 310.200 23.530 310.500 ;
        RECT 15.230 309.800 23.530 310.200 ;
        RECT 15.230 301.600 15.380 309.800 ;
        RECT 15.830 301.600 15.980 309.800 ;
        RECT 16.430 301.600 16.580 309.800 ;
        RECT 17.030 301.600 17.180 309.800 ;
        RECT 17.630 301.600 17.780 309.800 ;
        RECT 18.230 301.600 18.380 309.800 ;
        RECT 18.830 301.600 18.980 309.800 ;
        RECT 23.130 309.500 23.530 309.800 ;
        RECT 19.580 309.350 23.530 309.500 ;
        RECT 23.130 308.900 23.530 309.350 ;
        RECT 19.580 308.750 23.530 308.900 ;
        RECT 23.130 308.300 23.530 308.750 ;
        RECT 19.580 308.150 23.530 308.300 ;
        RECT 23.130 307.700 23.530 308.150 ;
        RECT 19.580 307.550 23.530 307.700 ;
        RECT 23.130 307.100 23.530 307.550 ;
        RECT 19.580 306.950 23.530 307.100 ;
        RECT 23.130 306.500 23.530 306.950 ;
        RECT 19.580 306.350 23.530 306.500 ;
        RECT 23.130 305.900 23.530 306.350 ;
        RECT 19.580 305.750 23.530 305.900 ;
        RECT 23.130 305.300 23.530 305.750 ;
        RECT 19.580 305.150 23.530 305.300 ;
        RECT 23.130 304.700 23.530 305.150 ;
        RECT 19.580 304.550 23.530 304.700 ;
        RECT 23.130 304.400 23.530 304.550 ;
        RECT 25.930 315.450 26.330 315.600 ;
        RECT 25.930 315.300 29.880 315.450 ;
        RECT 25.930 314.850 26.330 315.300 ;
        RECT 25.930 314.700 29.880 314.850 ;
        RECT 25.930 314.250 26.330 314.700 ;
        RECT 25.930 314.100 29.880 314.250 ;
        RECT 25.930 313.650 26.330 314.100 ;
        RECT 25.930 313.500 29.880 313.650 ;
        RECT 25.930 313.050 26.330 313.500 ;
        RECT 25.930 312.900 29.880 313.050 ;
        RECT 25.930 312.450 26.330 312.900 ;
        RECT 25.930 312.300 29.880 312.450 ;
        RECT 25.930 311.850 26.330 312.300 ;
        RECT 25.930 311.700 29.880 311.850 ;
        RECT 25.930 311.250 26.330 311.700 ;
        RECT 25.930 311.100 29.880 311.250 ;
        RECT 25.930 310.650 26.330 311.100 ;
        RECT 25.930 310.500 29.880 310.650 ;
        RECT 25.930 310.200 26.330 310.500 ;
        RECT 30.480 310.200 30.630 318.400 ;
        RECT 31.080 310.200 31.230 318.400 ;
        RECT 31.680 310.200 31.830 318.400 ;
        RECT 32.280 310.200 32.430 318.400 ;
        RECT 32.880 310.200 33.030 318.400 ;
        RECT 33.480 310.200 33.630 318.400 ;
        RECT 34.080 310.200 34.230 318.400 ;
        RECT 25.930 309.800 34.230 310.200 ;
        RECT 25.930 309.500 26.330 309.800 ;
        RECT 25.930 309.350 29.880 309.500 ;
        RECT 25.930 308.900 26.330 309.350 ;
        RECT 25.930 308.750 29.880 308.900 ;
        RECT 25.930 308.300 26.330 308.750 ;
        RECT 25.930 308.150 29.880 308.300 ;
        RECT 25.930 307.700 26.330 308.150 ;
        RECT 25.930 307.550 29.880 307.700 ;
        RECT 25.930 307.100 26.330 307.550 ;
        RECT 25.930 306.950 29.880 307.100 ;
        RECT 25.930 306.500 26.330 306.950 ;
        RECT 25.930 306.350 29.880 306.500 ;
        RECT 25.930 305.900 26.330 306.350 ;
        RECT 25.930 305.750 29.880 305.900 ;
        RECT 25.930 305.300 26.330 305.750 ;
        RECT 25.930 305.150 29.880 305.300 ;
        RECT 25.930 304.700 26.330 305.150 ;
        RECT 25.930 304.550 29.880 304.700 ;
        RECT 25.930 304.400 26.330 304.550 ;
        RECT 23.130 304.100 26.330 304.400 ;
        RECT 19.580 303.950 29.880 304.100 ;
        RECT 23.130 303.500 26.330 303.950 ;
        RECT 19.580 303.350 29.880 303.500 ;
        RECT 23.130 302.900 26.330 303.350 ;
        RECT 19.580 302.750 29.880 302.900 ;
        RECT 23.130 302.300 26.330 302.750 ;
        RECT 19.580 302.150 29.880 302.300 ;
        RECT 23.530 301.200 25.930 302.150 ;
        RECT 30.480 301.600 30.630 309.800 ;
        RECT 31.080 301.600 31.230 309.800 ;
        RECT 31.680 301.600 31.830 309.800 ;
        RECT 32.280 301.600 32.430 309.800 ;
        RECT 32.880 301.600 33.030 309.800 ;
        RECT 33.480 301.600 33.630 309.800 ;
        RECT 34.080 301.600 34.230 309.800 ;
        RECT 35.230 310.200 35.380 318.400 ;
        RECT 35.830 310.200 35.980 318.400 ;
        RECT 36.430 310.200 36.580 318.400 ;
        RECT 37.030 310.200 37.180 318.400 ;
        RECT 37.630 310.200 37.780 318.400 ;
        RECT 38.230 310.200 38.380 318.400 ;
        RECT 38.830 310.200 38.980 318.400 ;
        RECT 43.530 317.850 45.940 318.800 ;
        RECT 39.580 317.700 49.880 317.850 ;
        RECT 43.130 317.250 46.330 317.700 ;
        RECT 39.580 317.100 49.880 317.250 ;
        RECT 43.130 316.650 46.330 317.100 ;
        RECT 39.580 316.500 49.880 316.650 ;
        RECT 43.130 316.050 46.330 316.500 ;
        RECT 39.580 315.900 49.880 316.050 ;
        RECT 43.130 315.600 46.330 315.900 ;
        RECT 43.130 315.450 43.530 315.600 ;
        RECT 39.580 315.300 43.530 315.450 ;
        RECT 43.130 314.850 43.530 315.300 ;
        RECT 39.580 314.700 43.530 314.850 ;
        RECT 43.130 314.250 43.530 314.700 ;
        RECT 39.580 314.100 43.530 314.250 ;
        RECT 43.130 313.650 43.530 314.100 ;
        RECT 39.580 313.500 43.530 313.650 ;
        RECT 43.130 313.050 43.530 313.500 ;
        RECT 39.580 312.900 43.530 313.050 ;
        RECT 43.130 312.450 43.530 312.900 ;
        RECT 39.580 312.300 43.530 312.450 ;
        RECT 43.130 311.850 43.530 312.300 ;
        RECT 39.580 311.700 43.530 311.850 ;
        RECT 43.130 311.250 43.530 311.700 ;
        RECT 39.580 311.100 43.530 311.250 ;
        RECT 43.130 310.650 43.530 311.100 ;
        RECT 39.580 310.500 43.530 310.650 ;
        RECT 43.130 310.200 43.530 310.500 ;
        RECT 35.230 309.800 43.530 310.200 ;
        RECT 35.230 301.600 35.380 309.800 ;
        RECT 35.830 301.600 35.980 309.800 ;
        RECT 36.430 301.600 36.580 309.800 ;
        RECT 37.030 301.600 37.180 309.800 ;
        RECT 37.630 301.600 37.780 309.800 ;
        RECT 38.230 301.600 38.380 309.800 ;
        RECT 38.830 301.600 38.980 309.800 ;
        RECT 43.130 309.500 43.530 309.800 ;
        RECT 39.580 309.350 43.530 309.500 ;
        RECT 43.130 308.900 43.530 309.350 ;
        RECT 39.580 308.750 43.530 308.900 ;
        RECT 43.130 308.300 43.530 308.750 ;
        RECT 39.580 308.150 43.530 308.300 ;
        RECT 43.130 307.700 43.530 308.150 ;
        RECT 39.580 307.550 43.530 307.700 ;
        RECT 43.130 307.100 43.530 307.550 ;
        RECT 39.580 306.950 43.530 307.100 ;
        RECT 43.130 306.500 43.530 306.950 ;
        RECT 39.580 306.350 43.530 306.500 ;
        RECT 43.130 305.900 43.530 306.350 ;
        RECT 39.580 305.750 43.530 305.900 ;
        RECT 43.130 305.300 43.530 305.750 ;
        RECT 39.580 305.150 43.530 305.300 ;
        RECT 43.130 304.700 43.530 305.150 ;
        RECT 39.580 304.550 43.530 304.700 ;
        RECT 43.130 304.400 43.530 304.550 ;
        RECT 45.930 315.450 46.330 315.600 ;
        RECT 45.930 315.300 49.880 315.450 ;
        RECT 45.930 314.850 46.330 315.300 ;
        RECT 45.930 314.700 49.880 314.850 ;
        RECT 45.930 314.250 46.330 314.700 ;
        RECT 45.930 314.100 49.880 314.250 ;
        RECT 45.930 313.650 46.330 314.100 ;
        RECT 45.930 313.500 49.880 313.650 ;
        RECT 45.930 313.050 46.330 313.500 ;
        RECT 45.930 312.900 49.880 313.050 ;
        RECT 45.930 312.450 46.330 312.900 ;
        RECT 45.930 312.300 49.880 312.450 ;
        RECT 45.930 311.850 46.330 312.300 ;
        RECT 45.930 311.700 49.880 311.850 ;
        RECT 45.930 311.250 46.330 311.700 ;
        RECT 45.930 311.100 49.880 311.250 ;
        RECT 45.930 310.650 46.330 311.100 ;
        RECT 45.930 310.500 49.880 310.650 ;
        RECT 45.930 310.200 46.330 310.500 ;
        RECT 50.480 310.200 50.630 318.400 ;
        RECT 51.080 310.200 51.230 318.400 ;
        RECT 51.680 310.200 51.830 318.400 ;
        RECT 52.280 310.200 52.430 318.400 ;
        RECT 52.880 310.200 53.030 318.400 ;
        RECT 53.480 310.200 53.630 318.400 ;
        RECT 54.080 310.200 54.230 318.400 ;
        RECT 45.930 309.800 54.230 310.200 ;
        RECT 45.930 309.500 46.330 309.800 ;
        RECT 45.930 309.350 49.880 309.500 ;
        RECT 45.930 308.900 46.330 309.350 ;
        RECT 45.930 308.750 49.880 308.900 ;
        RECT 45.930 308.300 46.330 308.750 ;
        RECT 45.930 308.150 49.880 308.300 ;
        RECT 45.930 307.700 46.330 308.150 ;
        RECT 45.930 307.550 49.880 307.700 ;
        RECT 45.930 307.100 46.330 307.550 ;
        RECT 45.930 306.950 49.880 307.100 ;
        RECT 45.930 306.500 46.330 306.950 ;
        RECT 45.930 306.350 49.880 306.500 ;
        RECT 45.930 305.900 46.330 306.350 ;
        RECT 45.930 305.750 49.880 305.900 ;
        RECT 45.930 305.300 46.330 305.750 ;
        RECT 45.930 305.150 49.880 305.300 ;
        RECT 45.930 304.700 46.330 305.150 ;
        RECT 45.930 304.550 49.880 304.700 ;
        RECT 45.930 304.400 46.330 304.550 ;
        RECT 43.130 304.100 46.330 304.400 ;
        RECT 39.580 303.950 49.880 304.100 ;
        RECT 43.130 303.500 46.330 303.950 ;
        RECT 39.580 303.350 49.880 303.500 ;
        RECT 43.130 302.900 46.330 303.350 ;
        RECT 39.580 302.750 49.880 302.900 ;
        RECT 43.130 302.300 46.330 302.750 ;
        RECT 39.580 302.150 49.880 302.300 ;
        RECT 43.530 301.200 45.930 302.150 ;
        RECT 50.480 301.600 50.630 309.800 ;
        RECT 51.080 301.600 51.230 309.800 ;
        RECT 51.680 301.600 51.830 309.800 ;
        RECT 52.280 301.600 52.430 309.800 ;
        RECT 52.880 301.600 53.030 309.800 ;
        RECT 53.480 301.600 53.630 309.800 ;
        RECT 54.080 301.600 54.230 309.800 ;
        RECT 55.230 310.200 55.380 318.400 ;
        RECT 55.830 310.200 55.980 318.400 ;
        RECT 56.430 310.200 56.580 318.400 ;
        RECT 57.030 310.200 57.180 318.400 ;
        RECT 57.630 310.200 57.780 318.400 ;
        RECT 58.230 310.200 58.380 318.400 ;
        RECT 58.830 310.200 58.980 318.400 ;
        RECT 63.530 317.850 65.940 318.800 ;
        RECT 59.580 317.700 69.880 317.850 ;
        RECT 63.130 317.250 66.330 317.700 ;
        RECT 59.580 317.100 69.880 317.250 ;
        RECT 63.130 316.650 66.330 317.100 ;
        RECT 59.580 316.500 69.880 316.650 ;
        RECT 63.130 316.050 66.330 316.500 ;
        RECT 59.580 315.900 69.880 316.050 ;
        RECT 63.130 315.600 66.330 315.900 ;
        RECT 63.130 315.450 63.530 315.600 ;
        RECT 59.580 315.300 63.530 315.450 ;
        RECT 63.130 314.850 63.530 315.300 ;
        RECT 59.580 314.700 63.530 314.850 ;
        RECT 63.130 314.250 63.530 314.700 ;
        RECT 59.580 314.100 63.530 314.250 ;
        RECT 63.130 313.650 63.530 314.100 ;
        RECT 59.580 313.500 63.530 313.650 ;
        RECT 63.130 313.050 63.530 313.500 ;
        RECT 59.580 312.900 63.530 313.050 ;
        RECT 63.130 312.450 63.530 312.900 ;
        RECT 59.580 312.300 63.530 312.450 ;
        RECT 63.130 311.850 63.530 312.300 ;
        RECT 59.580 311.700 63.530 311.850 ;
        RECT 63.130 311.250 63.530 311.700 ;
        RECT 59.580 311.100 63.530 311.250 ;
        RECT 63.130 310.650 63.530 311.100 ;
        RECT 59.580 310.500 63.530 310.650 ;
        RECT 63.130 310.200 63.530 310.500 ;
        RECT 55.230 309.800 63.530 310.200 ;
        RECT 55.230 301.600 55.380 309.800 ;
        RECT 55.830 301.600 55.980 309.800 ;
        RECT 56.430 301.600 56.580 309.800 ;
        RECT 57.030 301.600 57.180 309.800 ;
        RECT 57.630 301.600 57.780 309.800 ;
        RECT 58.230 301.600 58.380 309.800 ;
        RECT 58.830 301.600 58.980 309.800 ;
        RECT 63.130 309.500 63.530 309.800 ;
        RECT 59.580 309.350 63.530 309.500 ;
        RECT 63.130 308.900 63.530 309.350 ;
        RECT 59.580 308.750 63.530 308.900 ;
        RECT 63.130 308.300 63.530 308.750 ;
        RECT 59.580 308.150 63.530 308.300 ;
        RECT 63.130 307.700 63.530 308.150 ;
        RECT 59.580 307.550 63.530 307.700 ;
        RECT 63.130 307.100 63.530 307.550 ;
        RECT 59.580 306.950 63.530 307.100 ;
        RECT 63.130 306.500 63.530 306.950 ;
        RECT 59.580 306.350 63.530 306.500 ;
        RECT 63.130 305.900 63.530 306.350 ;
        RECT 59.580 305.750 63.530 305.900 ;
        RECT 63.130 305.300 63.530 305.750 ;
        RECT 59.580 305.150 63.530 305.300 ;
        RECT 63.130 304.700 63.530 305.150 ;
        RECT 59.580 304.550 63.530 304.700 ;
        RECT 63.130 304.400 63.530 304.550 ;
        RECT 65.930 315.450 66.330 315.600 ;
        RECT 65.930 315.300 69.880 315.450 ;
        RECT 65.930 314.850 66.330 315.300 ;
        RECT 65.930 314.700 69.880 314.850 ;
        RECT 65.930 314.250 66.330 314.700 ;
        RECT 65.930 314.100 69.880 314.250 ;
        RECT 65.930 313.650 66.330 314.100 ;
        RECT 65.930 313.500 69.880 313.650 ;
        RECT 65.930 313.050 66.330 313.500 ;
        RECT 65.930 312.900 69.880 313.050 ;
        RECT 65.930 312.450 66.330 312.900 ;
        RECT 65.930 312.300 69.880 312.450 ;
        RECT 65.930 311.850 66.330 312.300 ;
        RECT 65.930 311.700 69.880 311.850 ;
        RECT 65.930 311.250 66.330 311.700 ;
        RECT 65.930 311.100 69.880 311.250 ;
        RECT 65.930 310.650 66.330 311.100 ;
        RECT 65.930 310.500 69.880 310.650 ;
        RECT 65.930 310.200 66.330 310.500 ;
        RECT 70.480 310.200 70.630 318.400 ;
        RECT 71.080 310.200 71.230 318.400 ;
        RECT 71.680 310.200 71.830 318.400 ;
        RECT 72.280 310.200 72.430 318.400 ;
        RECT 72.880 310.200 73.030 318.400 ;
        RECT 73.480 310.200 73.630 318.400 ;
        RECT 74.080 310.200 74.230 318.400 ;
        RECT 65.930 309.800 74.230 310.200 ;
        RECT 65.930 309.500 66.330 309.800 ;
        RECT 65.930 309.350 69.880 309.500 ;
        RECT 65.930 308.900 66.330 309.350 ;
        RECT 65.930 308.750 69.880 308.900 ;
        RECT 65.930 308.300 66.330 308.750 ;
        RECT 65.930 308.150 69.880 308.300 ;
        RECT 65.930 307.700 66.330 308.150 ;
        RECT 65.930 307.550 69.880 307.700 ;
        RECT 65.930 307.100 66.330 307.550 ;
        RECT 65.930 306.950 69.880 307.100 ;
        RECT 65.930 306.500 66.330 306.950 ;
        RECT 65.930 306.350 69.880 306.500 ;
        RECT 65.930 305.900 66.330 306.350 ;
        RECT 65.930 305.750 69.880 305.900 ;
        RECT 65.930 305.300 66.330 305.750 ;
        RECT 65.930 305.150 69.880 305.300 ;
        RECT 65.930 304.700 66.330 305.150 ;
        RECT 65.930 304.550 69.880 304.700 ;
        RECT 65.930 304.400 66.330 304.550 ;
        RECT 63.130 304.100 66.330 304.400 ;
        RECT 59.580 303.950 69.880 304.100 ;
        RECT 63.130 303.500 66.330 303.950 ;
        RECT 59.580 303.350 69.880 303.500 ;
        RECT 63.130 302.900 66.330 303.350 ;
        RECT 59.580 302.750 69.880 302.900 ;
        RECT 63.130 302.300 66.330 302.750 ;
        RECT 59.580 302.150 69.880 302.300 ;
        RECT 63.530 301.200 65.930 302.150 ;
        RECT 70.480 301.600 70.630 309.800 ;
        RECT 71.080 301.600 71.230 309.800 ;
        RECT 71.680 301.600 71.830 309.800 ;
        RECT 72.280 301.600 72.430 309.800 ;
        RECT 72.880 301.600 73.030 309.800 ;
        RECT 73.480 301.600 73.630 309.800 ;
        RECT 74.080 301.600 74.230 309.800 ;
        RECT 75.230 310.200 75.380 318.400 ;
        RECT 75.830 310.200 75.980 318.400 ;
        RECT 76.430 310.200 76.580 318.400 ;
        RECT 77.030 310.200 77.180 318.400 ;
        RECT 77.630 310.200 77.780 318.400 ;
        RECT 78.230 310.200 78.380 318.400 ;
        RECT 78.830 310.200 78.980 318.400 ;
        RECT 83.530 317.850 85.940 318.800 ;
        RECT 79.580 317.700 89.880 317.850 ;
        RECT 83.130 317.250 86.330 317.700 ;
        RECT 79.580 317.100 89.880 317.250 ;
        RECT 83.130 316.650 86.330 317.100 ;
        RECT 79.580 316.500 89.880 316.650 ;
        RECT 83.130 316.050 86.330 316.500 ;
        RECT 79.580 315.900 89.880 316.050 ;
        RECT 83.130 315.600 86.330 315.900 ;
        RECT 83.130 315.450 83.530 315.600 ;
        RECT 79.580 315.300 83.530 315.450 ;
        RECT 83.130 314.850 83.530 315.300 ;
        RECT 79.580 314.700 83.530 314.850 ;
        RECT 83.130 314.250 83.530 314.700 ;
        RECT 79.580 314.100 83.530 314.250 ;
        RECT 83.130 313.650 83.530 314.100 ;
        RECT 79.580 313.500 83.530 313.650 ;
        RECT 83.130 313.050 83.530 313.500 ;
        RECT 79.580 312.900 83.530 313.050 ;
        RECT 83.130 312.450 83.530 312.900 ;
        RECT 79.580 312.300 83.530 312.450 ;
        RECT 83.130 311.850 83.530 312.300 ;
        RECT 79.580 311.700 83.530 311.850 ;
        RECT 83.130 311.250 83.530 311.700 ;
        RECT 79.580 311.100 83.530 311.250 ;
        RECT 83.130 310.650 83.530 311.100 ;
        RECT 79.580 310.500 83.530 310.650 ;
        RECT 83.130 310.200 83.530 310.500 ;
        RECT 75.230 309.800 83.530 310.200 ;
        RECT 75.230 301.600 75.380 309.800 ;
        RECT 75.830 301.600 75.980 309.800 ;
        RECT 76.430 301.600 76.580 309.800 ;
        RECT 77.030 301.600 77.180 309.800 ;
        RECT 77.630 301.600 77.780 309.800 ;
        RECT 78.230 301.600 78.380 309.800 ;
        RECT 78.830 301.600 78.980 309.800 ;
        RECT 83.130 309.500 83.530 309.800 ;
        RECT 79.580 309.350 83.530 309.500 ;
        RECT 83.130 308.900 83.530 309.350 ;
        RECT 79.580 308.750 83.530 308.900 ;
        RECT 83.130 308.300 83.530 308.750 ;
        RECT 79.580 308.150 83.530 308.300 ;
        RECT 83.130 307.700 83.530 308.150 ;
        RECT 79.580 307.550 83.530 307.700 ;
        RECT 83.130 307.100 83.530 307.550 ;
        RECT 79.580 306.950 83.530 307.100 ;
        RECT 83.130 306.500 83.530 306.950 ;
        RECT 79.580 306.350 83.530 306.500 ;
        RECT 83.130 305.900 83.530 306.350 ;
        RECT 79.580 305.750 83.530 305.900 ;
        RECT 83.130 305.300 83.530 305.750 ;
        RECT 79.580 305.150 83.530 305.300 ;
        RECT 83.130 304.700 83.530 305.150 ;
        RECT 79.580 304.550 83.530 304.700 ;
        RECT 83.130 304.400 83.530 304.550 ;
        RECT 85.930 315.450 86.330 315.600 ;
        RECT 85.930 315.300 89.880 315.450 ;
        RECT 85.930 314.850 86.330 315.300 ;
        RECT 85.930 314.700 89.880 314.850 ;
        RECT 85.930 314.250 86.330 314.700 ;
        RECT 85.930 314.100 89.880 314.250 ;
        RECT 85.930 313.650 86.330 314.100 ;
        RECT 85.930 313.500 89.880 313.650 ;
        RECT 85.930 313.050 86.330 313.500 ;
        RECT 85.930 312.900 89.880 313.050 ;
        RECT 85.930 312.450 86.330 312.900 ;
        RECT 85.930 312.300 89.880 312.450 ;
        RECT 85.930 311.850 86.330 312.300 ;
        RECT 85.930 311.700 89.880 311.850 ;
        RECT 85.930 311.250 86.330 311.700 ;
        RECT 85.930 311.100 89.880 311.250 ;
        RECT 85.930 310.650 86.330 311.100 ;
        RECT 85.930 310.500 89.880 310.650 ;
        RECT 85.930 310.200 86.330 310.500 ;
        RECT 90.480 310.200 90.630 318.400 ;
        RECT 91.080 310.200 91.230 318.400 ;
        RECT 91.680 310.200 91.830 318.400 ;
        RECT 92.280 310.200 92.430 318.400 ;
        RECT 92.880 310.200 93.030 318.400 ;
        RECT 93.480 310.200 93.630 318.400 ;
        RECT 94.080 310.200 94.230 318.400 ;
        RECT 85.930 309.800 94.230 310.200 ;
        RECT 85.930 309.500 86.330 309.800 ;
        RECT 85.930 309.350 89.880 309.500 ;
        RECT 85.930 308.900 86.330 309.350 ;
        RECT 85.930 308.750 89.880 308.900 ;
        RECT 85.930 308.300 86.330 308.750 ;
        RECT 85.930 308.150 89.880 308.300 ;
        RECT 85.930 307.700 86.330 308.150 ;
        RECT 85.930 307.550 89.880 307.700 ;
        RECT 85.930 307.100 86.330 307.550 ;
        RECT 85.930 306.950 89.880 307.100 ;
        RECT 85.930 306.500 86.330 306.950 ;
        RECT 85.930 306.350 89.880 306.500 ;
        RECT 85.930 305.900 86.330 306.350 ;
        RECT 85.930 305.750 89.880 305.900 ;
        RECT 85.930 305.300 86.330 305.750 ;
        RECT 85.930 305.150 89.880 305.300 ;
        RECT 85.930 304.700 86.330 305.150 ;
        RECT 85.930 304.550 89.880 304.700 ;
        RECT 85.930 304.400 86.330 304.550 ;
        RECT 83.130 304.100 86.330 304.400 ;
        RECT 79.580 303.950 89.880 304.100 ;
        RECT 83.130 303.500 86.330 303.950 ;
        RECT 79.580 303.350 89.880 303.500 ;
        RECT 83.130 302.900 86.330 303.350 ;
        RECT 79.580 302.750 89.880 302.900 ;
        RECT 83.130 302.300 86.330 302.750 ;
        RECT 79.580 302.150 89.880 302.300 ;
        RECT 83.530 301.200 85.930 302.150 ;
        RECT 90.480 301.600 90.630 309.800 ;
        RECT 91.080 301.600 91.230 309.800 ;
        RECT 91.680 301.600 91.830 309.800 ;
        RECT 92.280 301.600 92.430 309.800 ;
        RECT 92.880 301.600 93.030 309.800 ;
        RECT 93.480 301.600 93.630 309.800 ;
        RECT 94.080 301.600 94.230 309.800 ;
        RECT 95.230 310.200 95.380 318.400 ;
        RECT 95.830 310.200 95.980 318.400 ;
        RECT 96.430 310.200 96.580 318.400 ;
        RECT 97.030 310.200 97.180 318.400 ;
        RECT 97.630 310.200 97.780 318.400 ;
        RECT 98.230 310.200 98.380 318.400 ;
        RECT 98.830 310.200 98.980 318.400 ;
        RECT 103.530 317.850 104.730 318.800 ;
        RECT 99.580 317.700 104.730 317.850 ;
        RECT 103.130 317.250 104.730 317.700 ;
        RECT 99.580 317.100 104.730 317.250 ;
        RECT 103.130 316.650 104.730 317.100 ;
        RECT 99.580 316.500 104.730 316.650 ;
        RECT 103.130 316.050 104.730 316.500 ;
        RECT 105.130 316.310 107.130 317.585 ;
        RECT 99.580 315.900 104.730 316.050 ;
        RECT 103.130 315.600 104.730 315.900 ;
        RECT 103.130 315.450 103.530 315.600 ;
        RECT 99.580 315.300 103.530 315.450 ;
        RECT 103.130 314.850 103.530 315.300 ;
        RECT 99.580 314.700 103.530 314.850 ;
        RECT 103.130 314.250 103.530 314.700 ;
        RECT 99.580 314.100 103.530 314.250 ;
        RECT 103.130 313.650 103.530 314.100 ;
        RECT 99.580 313.500 103.530 313.650 ;
        RECT 103.130 313.050 103.530 313.500 ;
        RECT 99.580 312.900 103.530 313.050 ;
        RECT 103.130 312.450 103.530 312.900 ;
        RECT 99.580 312.300 103.530 312.450 ;
        RECT 103.130 311.850 103.530 312.300 ;
        RECT 99.580 311.700 103.530 311.850 ;
        RECT 103.130 311.250 103.530 311.700 ;
        RECT 99.580 311.100 103.530 311.250 ;
        RECT 103.130 310.650 103.530 311.100 ;
        RECT 99.580 310.500 103.530 310.650 ;
        RECT 103.130 310.200 103.530 310.500 ;
        RECT 95.230 309.800 103.530 310.200 ;
        RECT 95.230 301.600 95.380 309.800 ;
        RECT 95.830 301.600 95.980 309.800 ;
        RECT 96.430 301.600 96.580 309.800 ;
        RECT 97.030 301.600 97.180 309.800 ;
        RECT 97.630 301.600 97.780 309.800 ;
        RECT 98.230 301.600 98.380 309.800 ;
        RECT 98.830 301.600 98.980 309.800 ;
        RECT 103.130 309.500 103.530 309.800 ;
        RECT 99.580 309.350 103.530 309.500 ;
        RECT 103.130 308.900 103.530 309.350 ;
        RECT 99.580 308.750 103.530 308.900 ;
        RECT 103.130 308.300 103.530 308.750 ;
        RECT 99.580 308.150 103.530 308.300 ;
        RECT 103.130 307.700 103.530 308.150 ;
        RECT 99.580 307.550 103.530 307.700 ;
        RECT 103.130 307.100 103.530 307.550 ;
        RECT 99.580 306.950 103.530 307.100 ;
        RECT 103.130 306.500 103.530 306.950 ;
        RECT 99.580 306.350 103.530 306.500 ;
        RECT 103.130 305.900 103.530 306.350 ;
        RECT 99.580 305.750 103.530 305.900 ;
        RECT 103.130 305.300 103.530 305.750 ;
        RECT 99.580 305.150 103.530 305.300 ;
        RECT 103.130 304.700 103.530 305.150 ;
        RECT 99.580 304.550 103.530 304.700 ;
        RECT 103.130 304.400 103.530 304.550 ;
        RECT 103.130 304.100 104.730 304.400 ;
        RECT 99.580 303.950 104.730 304.100 ;
        RECT 103.130 303.500 104.730 303.950 ;
        RECT 99.580 303.350 104.730 303.500 ;
        RECT 103.130 302.900 104.730 303.350 ;
        RECT 99.580 302.750 104.730 302.900 ;
        RECT 103.130 302.300 104.730 302.750 ;
        RECT 105.140 302.325 107.140 303.600 ;
        RECT 99.580 302.150 104.730 302.300 ;
        RECT 103.530 301.200 104.730 302.150 ;
        RECT 4.730 298.800 9.130 301.200 ;
        RECT 20.330 298.800 29.130 301.200 ;
        RECT 40.330 298.800 49.130 301.200 ;
        RECT 60.330 298.800 69.130 301.200 ;
        RECT 80.330 298.800 89.130 301.200 ;
        RECT 100.330 298.800 104.730 301.200 ;
        RECT 4.730 297.850 5.940 298.800 ;
        RECT 4.730 297.700 9.880 297.850 ;
        RECT 2.315 296.255 4.320 297.530 ;
        RECT 4.730 297.250 6.330 297.700 ;
        RECT 4.730 297.100 9.880 297.250 ;
        RECT 4.730 296.650 6.330 297.100 ;
        RECT 4.730 296.500 9.880 296.650 ;
        RECT 4.730 296.050 6.330 296.500 ;
        RECT 4.730 295.900 9.880 296.050 ;
        RECT 4.730 295.600 6.330 295.900 ;
        RECT 2.320 295.340 4.320 295.545 ;
        RECT 2.315 293.250 4.320 295.340 ;
        RECT 5.930 295.450 6.330 295.600 ;
        RECT 5.930 295.300 9.880 295.450 ;
        RECT 5.930 294.850 6.330 295.300 ;
        RECT 5.930 294.700 9.880 294.850 ;
        RECT 5.930 294.250 6.330 294.700 ;
        RECT 5.930 294.100 9.880 294.250 ;
        RECT 5.930 293.650 6.330 294.100 ;
        RECT 5.930 293.500 9.880 293.650 ;
        RECT 5.930 293.050 6.330 293.500 ;
        RECT 5.930 292.900 9.880 293.050 ;
        RECT 5.930 292.450 6.330 292.900 ;
        RECT 5.930 292.300 9.880 292.450 ;
        RECT 5.930 291.850 6.330 292.300 ;
        RECT 5.930 291.700 9.880 291.850 ;
        RECT 5.930 291.250 6.330 291.700 ;
        RECT 5.930 291.100 9.880 291.250 ;
        RECT 5.930 290.650 6.330 291.100 ;
        RECT 5.930 290.500 9.880 290.650 ;
        RECT 5.930 290.200 6.330 290.500 ;
        RECT 10.480 290.200 10.630 298.400 ;
        RECT 11.080 290.200 11.230 298.400 ;
        RECT 11.680 290.200 11.830 298.400 ;
        RECT 12.280 290.200 12.430 298.400 ;
        RECT 12.880 290.200 13.030 298.400 ;
        RECT 13.480 290.200 13.630 298.400 ;
        RECT 14.080 290.200 14.230 298.400 ;
        RECT 5.930 289.800 14.230 290.200 ;
        RECT 5.930 289.500 6.330 289.800 ;
        RECT 5.930 289.350 9.880 289.500 ;
        RECT 5.930 288.900 6.330 289.350 ;
        RECT 5.930 288.750 9.880 288.900 ;
        RECT 5.930 288.300 6.330 288.750 ;
        RECT 5.930 288.150 9.880 288.300 ;
        RECT 5.930 287.700 6.330 288.150 ;
        RECT 5.930 287.550 9.880 287.700 ;
        RECT 5.930 287.100 6.330 287.550 ;
        RECT 5.930 286.950 9.880 287.100 ;
        RECT 2.315 284.445 4.315 286.740 ;
        RECT 5.930 286.500 6.330 286.950 ;
        RECT 5.930 286.350 9.880 286.500 ;
        RECT 5.930 285.900 6.330 286.350 ;
        RECT 5.930 285.750 9.880 285.900 ;
        RECT 5.930 285.300 6.330 285.750 ;
        RECT 5.930 285.150 9.880 285.300 ;
        RECT 5.930 284.700 6.330 285.150 ;
        RECT 5.930 284.550 9.880 284.700 ;
        RECT 5.930 284.400 6.330 284.550 ;
        RECT 4.730 284.100 6.330 284.400 ;
        RECT 4.730 283.950 9.880 284.100 ;
        RECT 2.315 282.370 4.320 283.645 ;
        RECT 4.730 283.500 6.330 283.950 ;
        RECT 4.730 283.350 9.880 283.500 ;
        RECT 4.730 282.900 6.330 283.350 ;
        RECT 4.730 282.750 9.880 282.900 ;
        RECT 4.730 282.300 6.330 282.750 ;
        RECT 4.730 282.150 9.880 282.300 ;
        RECT 4.730 281.200 5.930 282.150 ;
        RECT 10.480 281.600 10.630 289.800 ;
        RECT 11.080 281.600 11.230 289.800 ;
        RECT 11.680 281.600 11.830 289.800 ;
        RECT 12.280 281.600 12.430 289.800 ;
        RECT 12.880 281.600 13.030 289.800 ;
        RECT 13.480 281.600 13.630 289.800 ;
        RECT 14.080 281.600 14.230 289.800 ;
        RECT 15.230 290.200 15.380 298.400 ;
        RECT 15.830 290.200 15.980 298.400 ;
        RECT 16.430 290.200 16.580 298.400 ;
        RECT 17.030 290.200 17.180 298.400 ;
        RECT 17.630 290.200 17.780 298.400 ;
        RECT 18.230 290.200 18.380 298.400 ;
        RECT 18.830 290.200 18.980 298.400 ;
        RECT 23.530 297.850 25.940 298.800 ;
        RECT 19.580 297.700 29.880 297.850 ;
        RECT 23.130 297.250 26.330 297.700 ;
        RECT 19.580 297.100 29.880 297.250 ;
        RECT 23.130 296.650 26.330 297.100 ;
        RECT 19.580 296.500 29.880 296.650 ;
        RECT 23.130 296.050 26.330 296.500 ;
        RECT 19.580 295.900 29.880 296.050 ;
        RECT 23.130 295.600 26.330 295.900 ;
        RECT 23.130 295.450 23.530 295.600 ;
        RECT 19.580 295.300 23.530 295.450 ;
        RECT 23.130 294.850 23.530 295.300 ;
        RECT 19.580 294.700 23.530 294.850 ;
        RECT 23.130 294.250 23.530 294.700 ;
        RECT 19.580 294.100 23.530 294.250 ;
        RECT 23.130 293.650 23.530 294.100 ;
        RECT 19.580 293.500 23.530 293.650 ;
        RECT 23.130 293.050 23.530 293.500 ;
        RECT 19.580 292.900 23.530 293.050 ;
        RECT 23.130 292.450 23.530 292.900 ;
        RECT 19.580 292.300 23.530 292.450 ;
        RECT 23.130 291.850 23.530 292.300 ;
        RECT 19.580 291.700 23.530 291.850 ;
        RECT 23.130 291.250 23.530 291.700 ;
        RECT 19.580 291.100 23.530 291.250 ;
        RECT 23.130 290.650 23.530 291.100 ;
        RECT 19.580 290.500 23.530 290.650 ;
        RECT 23.130 290.200 23.530 290.500 ;
        RECT 15.230 289.800 23.530 290.200 ;
        RECT 15.230 281.600 15.380 289.800 ;
        RECT 15.830 281.600 15.980 289.800 ;
        RECT 16.430 281.600 16.580 289.800 ;
        RECT 17.030 281.600 17.180 289.800 ;
        RECT 17.630 281.600 17.780 289.800 ;
        RECT 18.230 281.600 18.380 289.800 ;
        RECT 18.830 281.600 18.980 289.800 ;
        RECT 23.130 289.500 23.530 289.800 ;
        RECT 19.580 289.350 23.530 289.500 ;
        RECT 23.130 288.900 23.530 289.350 ;
        RECT 19.580 288.750 23.530 288.900 ;
        RECT 23.130 288.300 23.530 288.750 ;
        RECT 19.580 288.150 23.530 288.300 ;
        RECT 23.130 287.700 23.530 288.150 ;
        RECT 19.580 287.550 23.530 287.700 ;
        RECT 23.130 287.100 23.530 287.550 ;
        RECT 19.580 286.950 23.530 287.100 ;
        RECT 23.130 286.500 23.530 286.950 ;
        RECT 19.580 286.350 23.530 286.500 ;
        RECT 23.130 285.900 23.530 286.350 ;
        RECT 19.580 285.750 23.530 285.900 ;
        RECT 23.130 285.300 23.530 285.750 ;
        RECT 19.580 285.150 23.530 285.300 ;
        RECT 23.130 284.700 23.530 285.150 ;
        RECT 19.580 284.550 23.530 284.700 ;
        RECT 23.130 284.400 23.530 284.550 ;
        RECT 25.930 295.450 26.330 295.600 ;
        RECT 25.930 295.300 29.880 295.450 ;
        RECT 25.930 294.850 26.330 295.300 ;
        RECT 25.930 294.700 29.880 294.850 ;
        RECT 25.930 294.250 26.330 294.700 ;
        RECT 25.930 294.100 29.880 294.250 ;
        RECT 25.930 293.650 26.330 294.100 ;
        RECT 25.930 293.500 29.880 293.650 ;
        RECT 25.930 293.050 26.330 293.500 ;
        RECT 25.930 292.900 29.880 293.050 ;
        RECT 25.930 292.450 26.330 292.900 ;
        RECT 25.930 292.300 29.880 292.450 ;
        RECT 25.930 291.850 26.330 292.300 ;
        RECT 25.930 291.700 29.880 291.850 ;
        RECT 25.930 291.250 26.330 291.700 ;
        RECT 25.930 291.100 29.880 291.250 ;
        RECT 25.930 290.650 26.330 291.100 ;
        RECT 25.930 290.500 29.880 290.650 ;
        RECT 25.930 290.200 26.330 290.500 ;
        RECT 30.480 290.200 30.630 298.400 ;
        RECT 31.080 290.200 31.230 298.400 ;
        RECT 31.680 290.200 31.830 298.400 ;
        RECT 32.280 290.200 32.430 298.400 ;
        RECT 32.880 290.200 33.030 298.400 ;
        RECT 33.480 290.200 33.630 298.400 ;
        RECT 34.080 290.200 34.230 298.400 ;
        RECT 25.930 289.800 34.230 290.200 ;
        RECT 25.930 289.500 26.330 289.800 ;
        RECT 25.930 289.350 29.880 289.500 ;
        RECT 25.930 288.900 26.330 289.350 ;
        RECT 25.930 288.750 29.880 288.900 ;
        RECT 25.930 288.300 26.330 288.750 ;
        RECT 25.930 288.150 29.880 288.300 ;
        RECT 25.930 287.700 26.330 288.150 ;
        RECT 25.930 287.550 29.880 287.700 ;
        RECT 25.930 287.100 26.330 287.550 ;
        RECT 25.930 286.950 29.880 287.100 ;
        RECT 25.930 286.500 26.330 286.950 ;
        RECT 25.930 286.350 29.880 286.500 ;
        RECT 25.930 285.900 26.330 286.350 ;
        RECT 25.930 285.750 29.880 285.900 ;
        RECT 25.930 285.300 26.330 285.750 ;
        RECT 25.930 285.150 29.880 285.300 ;
        RECT 25.930 284.700 26.330 285.150 ;
        RECT 25.930 284.550 29.880 284.700 ;
        RECT 25.930 284.400 26.330 284.550 ;
        RECT 23.130 284.100 26.330 284.400 ;
        RECT 19.580 283.950 29.880 284.100 ;
        RECT 23.130 283.500 26.330 283.950 ;
        RECT 19.580 283.350 29.880 283.500 ;
        RECT 23.130 282.900 26.330 283.350 ;
        RECT 19.580 282.750 29.880 282.900 ;
        RECT 23.130 282.300 26.330 282.750 ;
        RECT 19.580 282.150 29.880 282.300 ;
        RECT 23.530 281.200 25.930 282.150 ;
        RECT 30.480 281.600 30.630 289.800 ;
        RECT 31.080 281.600 31.230 289.800 ;
        RECT 31.680 281.600 31.830 289.800 ;
        RECT 32.280 281.600 32.430 289.800 ;
        RECT 32.880 281.600 33.030 289.800 ;
        RECT 33.480 281.600 33.630 289.800 ;
        RECT 34.080 281.600 34.230 289.800 ;
        RECT 35.230 290.200 35.380 298.400 ;
        RECT 35.830 290.200 35.980 298.400 ;
        RECT 36.430 290.200 36.580 298.400 ;
        RECT 37.030 290.200 37.180 298.400 ;
        RECT 37.630 290.200 37.780 298.400 ;
        RECT 38.230 290.200 38.380 298.400 ;
        RECT 38.830 290.200 38.980 298.400 ;
        RECT 43.530 297.850 45.940 298.800 ;
        RECT 39.580 297.700 49.880 297.850 ;
        RECT 43.130 297.250 46.330 297.700 ;
        RECT 39.580 297.100 49.880 297.250 ;
        RECT 43.130 296.650 46.330 297.100 ;
        RECT 39.580 296.500 49.880 296.650 ;
        RECT 43.130 296.050 46.330 296.500 ;
        RECT 39.580 295.900 49.880 296.050 ;
        RECT 43.130 295.600 46.330 295.900 ;
        RECT 43.130 295.450 43.530 295.600 ;
        RECT 39.580 295.300 43.530 295.450 ;
        RECT 43.130 294.850 43.530 295.300 ;
        RECT 39.580 294.700 43.530 294.850 ;
        RECT 43.130 294.250 43.530 294.700 ;
        RECT 39.580 294.100 43.530 294.250 ;
        RECT 43.130 293.650 43.530 294.100 ;
        RECT 39.580 293.500 43.530 293.650 ;
        RECT 43.130 293.050 43.530 293.500 ;
        RECT 39.580 292.900 43.530 293.050 ;
        RECT 43.130 292.450 43.530 292.900 ;
        RECT 39.580 292.300 43.530 292.450 ;
        RECT 43.130 291.850 43.530 292.300 ;
        RECT 39.580 291.700 43.530 291.850 ;
        RECT 43.130 291.250 43.530 291.700 ;
        RECT 39.580 291.100 43.530 291.250 ;
        RECT 43.130 290.650 43.530 291.100 ;
        RECT 39.580 290.500 43.530 290.650 ;
        RECT 43.130 290.200 43.530 290.500 ;
        RECT 35.230 289.800 43.530 290.200 ;
        RECT 35.230 281.600 35.380 289.800 ;
        RECT 35.830 281.600 35.980 289.800 ;
        RECT 36.430 281.600 36.580 289.800 ;
        RECT 37.030 281.600 37.180 289.800 ;
        RECT 37.630 281.600 37.780 289.800 ;
        RECT 38.230 281.600 38.380 289.800 ;
        RECT 38.830 281.600 38.980 289.800 ;
        RECT 43.130 289.500 43.530 289.800 ;
        RECT 39.580 289.350 43.530 289.500 ;
        RECT 43.130 288.900 43.530 289.350 ;
        RECT 39.580 288.750 43.530 288.900 ;
        RECT 43.130 288.300 43.530 288.750 ;
        RECT 39.580 288.150 43.530 288.300 ;
        RECT 43.130 287.700 43.530 288.150 ;
        RECT 39.580 287.550 43.530 287.700 ;
        RECT 43.130 287.100 43.530 287.550 ;
        RECT 39.580 286.950 43.530 287.100 ;
        RECT 43.130 286.500 43.530 286.950 ;
        RECT 39.580 286.350 43.530 286.500 ;
        RECT 43.130 285.900 43.530 286.350 ;
        RECT 39.580 285.750 43.530 285.900 ;
        RECT 43.130 285.300 43.530 285.750 ;
        RECT 39.580 285.150 43.530 285.300 ;
        RECT 43.130 284.700 43.530 285.150 ;
        RECT 39.580 284.550 43.530 284.700 ;
        RECT 43.130 284.400 43.530 284.550 ;
        RECT 45.930 295.450 46.330 295.600 ;
        RECT 45.930 295.300 49.880 295.450 ;
        RECT 45.930 294.850 46.330 295.300 ;
        RECT 45.930 294.700 49.880 294.850 ;
        RECT 45.930 294.250 46.330 294.700 ;
        RECT 45.930 294.100 49.880 294.250 ;
        RECT 45.930 293.650 46.330 294.100 ;
        RECT 45.930 293.500 49.880 293.650 ;
        RECT 45.930 293.050 46.330 293.500 ;
        RECT 45.930 292.900 49.880 293.050 ;
        RECT 45.930 292.450 46.330 292.900 ;
        RECT 45.930 292.300 49.880 292.450 ;
        RECT 45.930 291.850 46.330 292.300 ;
        RECT 45.930 291.700 49.880 291.850 ;
        RECT 45.930 291.250 46.330 291.700 ;
        RECT 45.930 291.100 49.880 291.250 ;
        RECT 45.930 290.650 46.330 291.100 ;
        RECT 45.930 290.500 49.880 290.650 ;
        RECT 45.930 290.200 46.330 290.500 ;
        RECT 50.480 290.200 50.630 298.400 ;
        RECT 51.080 290.200 51.230 298.400 ;
        RECT 51.680 290.200 51.830 298.400 ;
        RECT 52.280 290.200 52.430 298.400 ;
        RECT 52.880 290.200 53.030 298.400 ;
        RECT 53.480 290.200 53.630 298.400 ;
        RECT 54.080 290.200 54.230 298.400 ;
        RECT 45.930 289.800 54.230 290.200 ;
        RECT 45.930 289.500 46.330 289.800 ;
        RECT 45.930 289.350 49.880 289.500 ;
        RECT 45.930 288.900 46.330 289.350 ;
        RECT 45.930 288.750 49.880 288.900 ;
        RECT 45.930 288.300 46.330 288.750 ;
        RECT 45.930 288.150 49.880 288.300 ;
        RECT 45.930 287.700 46.330 288.150 ;
        RECT 45.930 287.550 49.880 287.700 ;
        RECT 45.930 287.100 46.330 287.550 ;
        RECT 45.930 286.950 49.880 287.100 ;
        RECT 45.930 286.500 46.330 286.950 ;
        RECT 45.930 286.350 49.880 286.500 ;
        RECT 45.930 285.900 46.330 286.350 ;
        RECT 45.930 285.750 49.880 285.900 ;
        RECT 45.930 285.300 46.330 285.750 ;
        RECT 45.930 285.150 49.880 285.300 ;
        RECT 45.930 284.700 46.330 285.150 ;
        RECT 45.930 284.550 49.880 284.700 ;
        RECT 45.930 284.400 46.330 284.550 ;
        RECT 43.130 284.100 46.330 284.400 ;
        RECT 39.580 283.950 49.880 284.100 ;
        RECT 43.130 283.500 46.330 283.950 ;
        RECT 39.580 283.350 49.880 283.500 ;
        RECT 43.130 282.900 46.330 283.350 ;
        RECT 39.580 282.750 49.880 282.900 ;
        RECT 43.130 282.300 46.330 282.750 ;
        RECT 39.580 282.150 49.880 282.300 ;
        RECT 43.530 281.200 45.930 282.150 ;
        RECT 50.480 281.600 50.630 289.800 ;
        RECT 51.080 281.600 51.230 289.800 ;
        RECT 51.680 281.600 51.830 289.800 ;
        RECT 52.280 281.600 52.430 289.800 ;
        RECT 52.880 281.600 53.030 289.800 ;
        RECT 53.480 281.600 53.630 289.800 ;
        RECT 54.080 281.600 54.230 289.800 ;
        RECT 55.230 290.200 55.380 298.400 ;
        RECT 55.830 290.200 55.980 298.400 ;
        RECT 56.430 290.200 56.580 298.400 ;
        RECT 57.030 290.200 57.180 298.400 ;
        RECT 57.630 290.200 57.780 298.400 ;
        RECT 58.230 290.200 58.380 298.400 ;
        RECT 58.830 290.200 58.980 298.400 ;
        RECT 63.530 297.850 65.940 298.800 ;
        RECT 59.580 297.700 69.880 297.850 ;
        RECT 63.130 297.250 66.330 297.700 ;
        RECT 59.580 297.100 69.880 297.250 ;
        RECT 63.130 296.650 66.330 297.100 ;
        RECT 59.580 296.500 69.880 296.650 ;
        RECT 63.130 296.050 66.330 296.500 ;
        RECT 59.580 295.900 69.880 296.050 ;
        RECT 63.130 295.600 66.330 295.900 ;
        RECT 63.130 295.450 63.530 295.600 ;
        RECT 59.580 295.300 63.530 295.450 ;
        RECT 63.130 294.850 63.530 295.300 ;
        RECT 59.580 294.700 63.530 294.850 ;
        RECT 63.130 294.250 63.530 294.700 ;
        RECT 59.580 294.100 63.530 294.250 ;
        RECT 63.130 293.650 63.530 294.100 ;
        RECT 59.580 293.500 63.530 293.650 ;
        RECT 63.130 293.050 63.530 293.500 ;
        RECT 59.580 292.900 63.530 293.050 ;
        RECT 63.130 292.450 63.530 292.900 ;
        RECT 59.580 292.300 63.530 292.450 ;
        RECT 63.130 291.850 63.530 292.300 ;
        RECT 59.580 291.700 63.530 291.850 ;
        RECT 63.130 291.250 63.530 291.700 ;
        RECT 59.580 291.100 63.530 291.250 ;
        RECT 63.130 290.650 63.530 291.100 ;
        RECT 59.580 290.500 63.530 290.650 ;
        RECT 63.130 290.200 63.530 290.500 ;
        RECT 55.230 289.800 63.530 290.200 ;
        RECT 55.230 281.600 55.380 289.800 ;
        RECT 55.830 281.600 55.980 289.800 ;
        RECT 56.430 281.600 56.580 289.800 ;
        RECT 57.030 281.600 57.180 289.800 ;
        RECT 57.630 281.600 57.780 289.800 ;
        RECT 58.230 281.600 58.380 289.800 ;
        RECT 58.830 281.600 58.980 289.800 ;
        RECT 63.130 289.500 63.530 289.800 ;
        RECT 59.580 289.350 63.530 289.500 ;
        RECT 63.130 288.900 63.530 289.350 ;
        RECT 59.580 288.750 63.530 288.900 ;
        RECT 63.130 288.300 63.530 288.750 ;
        RECT 59.580 288.150 63.530 288.300 ;
        RECT 63.130 287.700 63.530 288.150 ;
        RECT 59.580 287.550 63.530 287.700 ;
        RECT 63.130 287.100 63.530 287.550 ;
        RECT 59.580 286.950 63.530 287.100 ;
        RECT 63.130 286.500 63.530 286.950 ;
        RECT 59.580 286.350 63.530 286.500 ;
        RECT 63.130 285.900 63.530 286.350 ;
        RECT 59.580 285.750 63.530 285.900 ;
        RECT 63.130 285.300 63.530 285.750 ;
        RECT 59.580 285.150 63.530 285.300 ;
        RECT 63.130 284.700 63.530 285.150 ;
        RECT 59.580 284.550 63.530 284.700 ;
        RECT 63.130 284.400 63.530 284.550 ;
        RECT 65.930 295.450 66.330 295.600 ;
        RECT 65.930 295.300 69.880 295.450 ;
        RECT 65.930 294.850 66.330 295.300 ;
        RECT 65.930 294.700 69.880 294.850 ;
        RECT 65.930 294.250 66.330 294.700 ;
        RECT 65.930 294.100 69.880 294.250 ;
        RECT 65.930 293.650 66.330 294.100 ;
        RECT 65.930 293.500 69.880 293.650 ;
        RECT 65.930 293.050 66.330 293.500 ;
        RECT 65.930 292.900 69.880 293.050 ;
        RECT 65.930 292.450 66.330 292.900 ;
        RECT 65.930 292.300 69.880 292.450 ;
        RECT 65.930 291.850 66.330 292.300 ;
        RECT 65.930 291.700 69.880 291.850 ;
        RECT 65.930 291.250 66.330 291.700 ;
        RECT 65.930 291.100 69.880 291.250 ;
        RECT 65.930 290.650 66.330 291.100 ;
        RECT 65.930 290.500 69.880 290.650 ;
        RECT 65.930 290.200 66.330 290.500 ;
        RECT 70.480 290.200 70.630 298.400 ;
        RECT 71.080 290.200 71.230 298.400 ;
        RECT 71.680 290.200 71.830 298.400 ;
        RECT 72.280 290.200 72.430 298.400 ;
        RECT 72.880 290.200 73.030 298.400 ;
        RECT 73.480 290.200 73.630 298.400 ;
        RECT 74.080 290.200 74.230 298.400 ;
        RECT 65.930 289.800 74.230 290.200 ;
        RECT 65.930 289.500 66.330 289.800 ;
        RECT 65.930 289.350 69.880 289.500 ;
        RECT 65.930 288.900 66.330 289.350 ;
        RECT 65.930 288.750 69.880 288.900 ;
        RECT 65.930 288.300 66.330 288.750 ;
        RECT 65.930 288.150 69.880 288.300 ;
        RECT 65.930 287.700 66.330 288.150 ;
        RECT 65.930 287.550 69.880 287.700 ;
        RECT 65.930 287.100 66.330 287.550 ;
        RECT 65.930 286.950 69.880 287.100 ;
        RECT 65.930 286.500 66.330 286.950 ;
        RECT 65.930 286.350 69.880 286.500 ;
        RECT 65.930 285.900 66.330 286.350 ;
        RECT 65.930 285.750 69.880 285.900 ;
        RECT 65.930 285.300 66.330 285.750 ;
        RECT 65.930 285.150 69.880 285.300 ;
        RECT 65.930 284.700 66.330 285.150 ;
        RECT 65.930 284.550 69.880 284.700 ;
        RECT 65.930 284.400 66.330 284.550 ;
        RECT 63.130 284.100 66.330 284.400 ;
        RECT 59.580 283.950 69.880 284.100 ;
        RECT 63.130 283.500 66.330 283.950 ;
        RECT 59.580 283.350 69.880 283.500 ;
        RECT 63.130 282.900 66.330 283.350 ;
        RECT 59.580 282.750 69.880 282.900 ;
        RECT 63.130 282.300 66.330 282.750 ;
        RECT 59.580 282.150 69.880 282.300 ;
        RECT 63.530 281.200 65.930 282.150 ;
        RECT 70.480 281.600 70.630 289.800 ;
        RECT 71.080 281.600 71.230 289.800 ;
        RECT 71.680 281.600 71.830 289.800 ;
        RECT 72.280 281.600 72.430 289.800 ;
        RECT 72.880 281.600 73.030 289.800 ;
        RECT 73.480 281.600 73.630 289.800 ;
        RECT 74.080 281.600 74.230 289.800 ;
        RECT 75.230 290.200 75.380 298.400 ;
        RECT 75.830 290.200 75.980 298.400 ;
        RECT 76.430 290.200 76.580 298.400 ;
        RECT 77.030 290.200 77.180 298.400 ;
        RECT 77.630 290.200 77.780 298.400 ;
        RECT 78.230 290.200 78.380 298.400 ;
        RECT 78.830 290.200 78.980 298.400 ;
        RECT 83.530 297.850 85.940 298.800 ;
        RECT 79.580 297.700 89.880 297.850 ;
        RECT 83.130 297.250 86.330 297.700 ;
        RECT 79.580 297.100 89.880 297.250 ;
        RECT 83.130 296.650 86.330 297.100 ;
        RECT 79.580 296.500 89.880 296.650 ;
        RECT 83.130 296.050 86.330 296.500 ;
        RECT 79.580 295.900 89.880 296.050 ;
        RECT 83.130 295.600 86.330 295.900 ;
        RECT 83.130 295.450 83.530 295.600 ;
        RECT 79.580 295.300 83.530 295.450 ;
        RECT 83.130 294.850 83.530 295.300 ;
        RECT 79.580 294.700 83.530 294.850 ;
        RECT 83.130 294.250 83.530 294.700 ;
        RECT 79.580 294.100 83.530 294.250 ;
        RECT 83.130 293.650 83.530 294.100 ;
        RECT 79.580 293.500 83.530 293.650 ;
        RECT 83.130 293.050 83.530 293.500 ;
        RECT 79.580 292.900 83.530 293.050 ;
        RECT 83.130 292.450 83.530 292.900 ;
        RECT 79.580 292.300 83.530 292.450 ;
        RECT 83.130 291.850 83.530 292.300 ;
        RECT 79.580 291.700 83.530 291.850 ;
        RECT 83.130 291.250 83.530 291.700 ;
        RECT 79.580 291.100 83.530 291.250 ;
        RECT 83.130 290.650 83.530 291.100 ;
        RECT 79.580 290.500 83.530 290.650 ;
        RECT 83.130 290.200 83.530 290.500 ;
        RECT 75.230 289.800 83.530 290.200 ;
        RECT 75.230 281.600 75.380 289.800 ;
        RECT 75.830 281.600 75.980 289.800 ;
        RECT 76.430 281.600 76.580 289.800 ;
        RECT 77.030 281.600 77.180 289.800 ;
        RECT 77.630 281.600 77.780 289.800 ;
        RECT 78.230 281.600 78.380 289.800 ;
        RECT 78.830 281.600 78.980 289.800 ;
        RECT 83.130 289.500 83.530 289.800 ;
        RECT 79.580 289.350 83.530 289.500 ;
        RECT 83.130 288.900 83.530 289.350 ;
        RECT 79.580 288.750 83.530 288.900 ;
        RECT 83.130 288.300 83.530 288.750 ;
        RECT 79.580 288.150 83.530 288.300 ;
        RECT 83.130 287.700 83.530 288.150 ;
        RECT 79.580 287.550 83.530 287.700 ;
        RECT 83.130 287.100 83.530 287.550 ;
        RECT 79.580 286.950 83.530 287.100 ;
        RECT 83.130 286.500 83.530 286.950 ;
        RECT 79.580 286.350 83.530 286.500 ;
        RECT 83.130 285.900 83.530 286.350 ;
        RECT 79.580 285.750 83.530 285.900 ;
        RECT 83.130 285.300 83.530 285.750 ;
        RECT 79.580 285.150 83.530 285.300 ;
        RECT 83.130 284.700 83.530 285.150 ;
        RECT 79.580 284.550 83.530 284.700 ;
        RECT 83.130 284.400 83.530 284.550 ;
        RECT 85.930 295.450 86.330 295.600 ;
        RECT 85.930 295.300 89.880 295.450 ;
        RECT 85.930 294.850 86.330 295.300 ;
        RECT 85.930 294.700 89.880 294.850 ;
        RECT 85.930 294.250 86.330 294.700 ;
        RECT 85.930 294.100 89.880 294.250 ;
        RECT 85.930 293.650 86.330 294.100 ;
        RECT 85.930 293.500 89.880 293.650 ;
        RECT 85.930 293.050 86.330 293.500 ;
        RECT 85.930 292.900 89.880 293.050 ;
        RECT 85.930 292.450 86.330 292.900 ;
        RECT 85.930 292.300 89.880 292.450 ;
        RECT 85.930 291.850 86.330 292.300 ;
        RECT 85.930 291.700 89.880 291.850 ;
        RECT 85.930 291.250 86.330 291.700 ;
        RECT 85.930 291.100 89.880 291.250 ;
        RECT 85.930 290.650 86.330 291.100 ;
        RECT 85.930 290.500 89.880 290.650 ;
        RECT 85.930 290.200 86.330 290.500 ;
        RECT 90.480 290.200 90.630 298.400 ;
        RECT 91.080 290.200 91.230 298.400 ;
        RECT 91.680 290.200 91.830 298.400 ;
        RECT 92.280 290.200 92.430 298.400 ;
        RECT 92.880 290.200 93.030 298.400 ;
        RECT 93.480 290.200 93.630 298.400 ;
        RECT 94.080 290.200 94.230 298.400 ;
        RECT 85.930 289.800 94.230 290.200 ;
        RECT 85.930 289.500 86.330 289.800 ;
        RECT 85.930 289.350 89.880 289.500 ;
        RECT 85.930 288.900 86.330 289.350 ;
        RECT 85.930 288.750 89.880 288.900 ;
        RECT 85.930 288.300 86.330 288.750 ;
        RECT 85.930 288.150 89.880 288.300 ;
        RECT 85.930 287.700 86.330 288.150 ;
        RECT 85.930 287.550 89.880 287.700 ;
        RECT 85.930 287.100 86.330 287.550 ;
        RECT 85.930 286.950 89.880 287.100 ;
        RECT 85.930 286.500 86.330 286.950 ;
        RECT 85.930 286.350 89.880 286.500 ;
        RECT 85.930 285.900 86.330 286.350 ;
        RECT 85.930 285.750 89.880 285.900 ;
        RECT 85.930 285.300 86.330 285.750 ;
        RECT 85.930 285.150 89.880 285.300 ;
        RECT 85.930 284.700 86.330 285.150 ;
        RECT 85.930 284.550 89.880 284.700 ;
        RECT 85.930 284.400 86.330 284.550 ;
        RECT 83.130 284.100 86.330 284.400 ;
        RECT 79.580 283.950 89.880 284.100 ;
        RECT 83.130 283.500 86.330 283.950 ;
        RECT 79.580 283.350 89.880 283.500 ;
        RECT 83.130 282.900 86.330 283.350 ;
        RECT 79.580 282.750 89.880 282.900 ;
        RECT 83.130 282.300 86.330 282.750 ;
        RECT 79.580 282.150 89.880 282.300 ;
        RECT 83.530 281.200 85.930 282.150 ;
        RECT 90.480 281.600 90.630 289.800 ;
        RECT 91.080 281.600 91.230 289.800 ;
        RECT 91.680 281.600 91.830 289.800 ;
        RECT 92.280 281.600 92.430 289.800 ;
        RECT 92.880 281.600 93.030 289.800 ;
        RECT 93.480 281.600 93.630 289.800 ;
        RECT 94.080 281.600 94.230 289.800 ;
        RECT 95.230 290.200 95.380 298.400 ;
        RECT 95.830 290.200 95.980 298.400 ;
        RECT 96.430 290.200 96.580 298.400 ;
        RECT 97.030 290.200 97.180 298.400 ;
        RECT 97.630 290.200 97.780 298.400 ;
        RECT 98.230 290.200 98.380 298.400 ;
        RECT 98.830 290.200 98.980 298.400 ;
        RECT 103.530 297.850 104.730 298.800 ;
        RECT 99.580 297.700 104.730 297.850 ;
        RECT 103.130 297.250 104.730 297.700 ;
        RECT 99.580 297.100 104.730 297.250 ;
        RECT 103.130 296.650 104.730 297.100 ;
        RECT 99.580 296.500 104.730 296.650 ;
        RECT 105.135 296.580 107.135 297.855 ;
        RECT 103.130 296.050 104.730 296.500 ;
        RECT 99.580 295.900 104.730 296.050 ;
        RECT 103.130 295.600 104.730 295.900 ;
        RECT 103.130 295.450 103.530 295.600 ;
        RECT 99.580 295.300 103.530 295.450 ;
        RECT 103.130 294.850 103.530 295.300 ;
        RECT 99.580 294.700 103.530 294.850 ;
        RECT 103.130 294.250 103.530 294.700 ;
        RECT 99.580 294.100 103.530 294.250 ;
        RECT 103.130 293.650 103.530 294.100 ;
        RECT 99.580 293.500 103.530 293.650 ;
        RECT 103.130 293.050 103.530 293.500 ;
        RECT 99.580 292.900 103.530 293.050 ;
        RECT 103.130 292.450 103.530 292.900 ;
        RECT 99.580 292.300 103.530 292.450 ;
        RECT 103.130 291.850 103.530 292.300 ;
        RECT 99.580 291.700 103.530 291.850 ;
        RECT 103.130 291.250 103.530 291.700 ;
        RECT 99.580 291.100 103.530 291.250 ;
        RECT 103.130 290.650 103.530 291.100 ;
        RECT 99.580 290.500 103.530 290.650 ;
        RECT 103.130 290.200 103.530 290.500 ;
        RECT 95.230 289.800 103.530 290.200 ;
        RECT 95.230 281.600 95.380 289.800 ;
        RECT 95.830 281.600 95.980 289.800 ;
        RECT 96.430 281.600 96.580 289.800 ;
        RECT 97.030 281.600 97.180 289.800 ;
        RECT 97.630 281.600 97.780 289.800 ;
        RECT 98.230 281.600 98.380 289.800 ;
        RECT 98.830 281.600 98.980 289.800 ;
        RECT 103.130 289.500 103.530 289.800 ;
        RECT 99.580 289.350 103.530 289.500 ;
        RECT 103.130 288.900 103.530 289.350 ;
        RECT 99.580 288.750 103.530 288.900 ;
        RECT 103.130 288.300 103.530 288.750 ;
        RECT 99.580 288.150 103.530 288.300 ;
        RECT 103.130 287.700 103.530 288.150 ;
        RECT 99.580 287.550 103.530 287.700 ;
        RECT 103.130 287.100 103.530 287.550 ;
        RECT 99.580 286.950 103.530 287.100 ;
        RECT 103.130 286.500 103.530 286.950 ;
        RECT 99.580 286.350 103.530 286.500 ;
        RECT 103.130 285.900 103.530 286.350 ;
        RECT 99.580 285.750 103.530 285.900 ;
        RECT 103.130 285.300 103.530 285.750 ;
        RECT 99.580 285.150 103.530 285.300 ;
        RECT 103.130 284.700 103.530 285.150 ;
        RECT 99.580 284.550 103.530 284.700 ;
        RECT 103.130 284.400 103.530 284.550 ;
        RECT 103.130 284.100 104.730 284.400 ;
        RECT 99.580 283.950 104.730 284.100 ;
        RECT 103.130 283.500 104.730 283.950 ;
        RECT 99.580 283.350 104.730 283.500 ;
        RECT 103.130 282.900 104.730 283.350 ;
        RECT 99.580 282.750 104.730 282.900 ;
        RECT 103.130 282.300 104.730 282.750 ;
        RECT 99.580 282.150 104.730 282.300 ;
        RECT 103.530 281.200 104.730 282.150 ;
        RECT 105.140 282.000 107.140 283.275 ;
        RECT 4.730 278.800 9.130 281.200 ;
        RECT 20.330 278.800 29.130 281.200 ;
        RECT 40.330 278.800 49.130 281.200 ;
        RECT 60.330 278.800 69.130 281.200 ;
        RECT 80.330 278.800 89.130 281.200 ;
        RECT 100.330 278.800 104.730 281.200 ;
        RECT 4.730 277.850 5.940 278.800 ;
        RECT 4.730 277.700 9.880 277.850 ;
        RECT 2.315 276.335 4.330 277.610 ;
        RECT 4.730 277.250 6.330 277.700 ;
        RECT 4.730 277.100 9.880 277.250 ;
        RECT 4.730 276.650 6.330 277.100 ;
        RECT 4.730 276.500 9.880 276.650 ;
        RECT 4.730 276.050 6.330 276.500 ;
        RECT 4.730 275.900 9.880 276.050 ;
        RECT 4.730 275.600 6.330 275.900 ;
        RECT 2.315 273.250 4.315 275.545 ;
        RECT 5.930 275.450 6.330 275.600 ;
        RECT 5.930 275.300 9.880 275.450 ;
        RECT 5.930 274.850 6.330 275.300 ;
        RECT 5.930 274.700 9.880 274.850 ;
        RECT 5.930 274.250 6.330 274.700 ;
        RECT 5.930 274.100 9.880 274.250 ;
        RECT 5.930 273.650 6.330 274.100 ;
        RECT 5.930 273.500 9.880 273.650 ;
        RECT 5.930 273.050 6.330 273.500 ;
        RECT 5.930 272.900 9.880 273.050 ;
        RECT 5.930 272.450 6.330 272.900 ;
        RECT 5.930 272.300 9.880 272.450 ;
        RECT 5.930 271.850 6.330 272.300 ;
        RECT 5.930 271.700 9.880 271.850 ;
        RECT 5.930 271.250 6.330 271.700 ;
        RECT 5.930 271.100 9.880 271.250 ;
        RECT 5.930 270.650 6.330 271.100 ;
        RECT 5.930 270.500 9.880 270.650 ;
        RECT 5.930 270.200 6.330 270.500 ;
        RECT 10.480 270.200 10.630 278.400 ;
        RECT 11.080 270.200 11.230 278.400 ;
        RECT 11.680 270.200 11.830 278.400 ;
        RECT 12.280 270.200 12.430 278.400 ;
        RECT 12.880 270.200 13.030 278.400 ;
        RECT 13.480 270.200 13.630 278.400 ;
        RECT 14.080 270.200 14.230 278.400 ;
        RECT 5.930 269.800 14.230 270.200 ;
        RECT 5.930 269.500 6.330 269.800 ;
        RECT 5.930 269.350 9.880 269.500 ;
        RECT 5.930 268.900 6.330 269.350 ;
        RECT 5.930 268.750 9.880 268.900 ;
        RECT 5.930 268.300 6.330 268.750 ;
        RECT 5.930 268.150 9.880 268.300 ;
        RECT 5.930 267.700 6.330 268.150 ;
        RECT 5.930 267.550 9.880 267.700 ;
        RECT 5.930 267.100 6.330 267.550 ;
        RECT 5.930 266.950 9.880 267.100 ;
        RECT 2.315 264.455 4.315 266.750 ;
        RECT 5.930 266.500 6.330 266.950 ;
        RECT 5.930 266.350 9.880 266.500 ;
        RECT 5.930 265.900 6.330 266.350 ;
        RECT 5.930 265.750 9.880 265.900 ;
        RECT 5.930 265.300 6.330 265.750 ;
        RECT 5.930 265.150 9.880 265.300 ;
        RECT 5.930 264.700 6.330 265.150 ;
        RECT 5.930 264.550 9.880 264.700 ;
        RECT 5.930 264.400 6.330 264.550 ;
        RECT 4.730 264.100 6.330 264.400 ;
        RECT 4.730 263.950 9.880 264.100 ;
        RECT 2.315 262.505 4.320 263.780 ;
        RECT 4.730 263.500 6.330 263.950 ;
        RECT 4.730 263.350 9.880 263.500 ;
        RECT 4.730 262.900 6.330 263.350 ;
        RECT 4.730 262.750 9.880 262.900 ;
        RECT 4.730 262.300 6.330 262.750 ;
        RECT 4.730 262.150 9.880 262.300 ;
        RECT 4.730 261.200 5.930 262.150 ;
        RECT 10.480 261.600 10.630 269.800 ;
        RECT 11.080 261.600 11.230 269.800 ;
        RECT 11.680 261.600 11.830 269.800 ;
        RECT 12.280 261.600 12.430 269.800 ;
        RECT 12.880 261.600 13.030 269.800 ;
        RECT 13.480 261.600 13.630 269.800 ;
        RECT 14.080 261.600 14.230 269.800 ;
        RECT 15.230 270.200 15.380 278.400 ;
        RECT 15.830 270.200 15.980 278.400 ;
        RECT 16.430 270.200 16.580 278.400 ;
        RECT 17.030 270.200 17.180 278.400 ;
        RECT 17.630 270.200 17.780 278.400 ;
        RECT 18.230 270.200 18.380 278.400 ;
        RECT 18.830 270.200 18.980 278.400 ;
        RECT 23.530 277.850 25.940 278.800 ;
        RECT 19.580 277.700 29.880 277.850 ;
        RECT 23.130 277.250 26.330 277.700 ;
        RECT 19.580 277.100 29.880 277.250 ;
        RECT 23.130 276.650 26.330 277.100 ;
        RECT 19.580 276.500 29.880 276.650 ;
        RECT 23.130 276.050 26.330 276.500 ;
        RECT 19.580 275.900 29.880 276.050 ;
        RECT 23.130 275.600 26.330 275.900 ;
        RECT 23.130 275.450 23.530 275.600 ;
        RECT 19.580 275.300 23.530 275.450 ;
        RECT 23.130 274.850 23.530 275.300 ;
        RECT 19.580 274.700 23.530 274.850 ;
        RECT 23.130 274.250 23.530 274.700 ;
        RECT 19.580 274.100 23.530 274.250 ;
        RECT 23.130 273.650 23.530 274.100 ;
        RECT 19.580 273.500 23.530 273.650 ;
        RECT 23.130 273.050 23.530 273.500 ;
        RECT 19.580 272.900 23.530 273.050 ;
        RECT 23.130 272.450 23.530 272.900 ;
        RECT 19.580 272.300 23.530 272.450 ;
        RECT 23.130 271.850 23.530 272.300 ;
        RECT 19.580 271.700 23.530 271.850 ;
        RECT 23.130 271.250 23.530 271.700 ;
        RECT 19.580 271.100 23.530 271.250 ;
        RECT 23.130 270.650 23.530 271.100 ;
        RECT 19.580 270.500 23.530 270.650 ;
        RECT 23.130 270.200 23.530 270.500 ;
        RECT 15.230 269.800 23.530 270.200 ;
        RECT 15.230 261.600 15.380 269.800 ;
        RECT 15.830 261.600 15.980 269.800 ;
        RECT 16.430 261.600 16.580 269.800 ;
        RECT 17.030 261.600 17.180 269.800 ;
        RECT 17.630 261.600 17.780 269.800 ;
        RECT 18.230 261.600 18.380 269.800 ;
        RECT 18.830 261.600 18.980 269.800 ;
        RECT 23.130 269.500 23.530 269.800 ;
        RECT 19.580 269.350 23.530 269.500 ;
        RECT 23.130 268.900 23.530 269.350 ;
        RECT 19.580 268.750 23.530 268.900 ;
        RECT 23.130 268.300 23.530 268.750 ;
        RECT 19.580 268.150 23.530 268.300 ;
        RECT 23.130 267.700 23.530 268.150 ;
        RECT 19.580 267.550 23.530 267.700 ;
        RECT 23.130 267.100 23.530 267.550 ;
        RECT 19.580 266.950 23.530 267.100 ;
        RECT 23.130 266.500 23.530 266.950 ;
        RECT 19.580 266.350 23.530 266.500 ;
        RECT 23.130 265.900 23.530 266.350 ;
        RECT 19.580 265.750 23.530 265.900 ;
        RECT 23.130 265.300 23.530 265.750 ;
        RECT 19.580 265.150 23.530 265.300 ;
        RECT 23.130 264.700 23.530 265.150 ;
        RECT 19.580 264.550 23.530 264.700 ;
        RECT 23.130 264.400 23.530 264.550 ;
        RECT 25.930 275.450 26.330 275.600 ;
        RECT 25.930 275.300 29.880 275.450 ;
        RECT 25.930 274.850 26.330 275.300 ;
        RECT 25.930 274.700 29.880 274.850 ;
        RECT 25.930 274.250 26.330 274.700 ;
        RECT 25.930 274.100 29.880 274.250 ;
        RECT 25.930 273.650 26.330 274.100 ;
        RECT 25.930 273.500 29.880 273.650 ;
        RECT 25.930 273.050 26.330 273.500 ;
        RECT 25.930 272.900 29.880 273.050 ;
        RECT 25.930 272.450 26.330 272.900 ;
        RECT 25.930 272.300 29.880 272.450 ;
        RECT 25.930 271.850 26.330 272.300 ;
        RECT 25.930 271.700 29.880 271.850 ;
        RECT 25.930 271.250 26.330 271.700 ;
        RECT 25.930 271.100 29.880 271.250 ;
        RECT 25.930 270.650 26.330 271.100 ;
        RECT 25.930 270.500 29.880 270.650 ;
        RECT 25.930 270.200 26.330 270.500 ;
        RECT 30.480 270.200 30.630 278.400 ;
        RECT 31.080 270.200 31.230 278.400 ;
        RECT 31.680 270.200 31.830 278.400 ;
        RECT 32.280 270.200 32.430 278.400 ;
        RECT 32.880 270.200 33.030 278.400 ;
        RECT 33.480 270.200 33.630 278.400 ;
        RECT 34.080 270.200 34.230 278.400 ;
        RECT 25.930 269.800 34.230 270.200 ;
        RECT 25.930 269.500 26.330 269.800 ;
        RECT 25.930 269.350 29.880 269.500 ;
        RECT 25.930 268.900 26.330 269.350 ;
        RECT 25.930 268.750 29.880 268.900 ;
        RECT 25.930 268.300 26.330 268.750 ;
        RECT 25.930 268.150 29.880 268.300 ;
        RECT 25.930 267.700 26.330 268.150 ;
        RECT 25.930 267.550 29.880 267.700 ;
        RECT 25.930 267.100 26.330 267.550 ;
        RECT 25.930 266.950 29.880 267.100 ;
        RECT 25.930 266.500 26.330 266.950 ;
        RECT 25.930 266.350 29.880 266.500 ;
        RECT 25.930 265.900 26.330 266.350 ;
        RECT 25.930 265.750 29.880 265.900 ;
        RECT 25.930 265.300 26.330 265.750 ;
        RECT 25.930 265.150 29.880 265.300 ;
        RECT 25.930 264.700 26.330 265.150 ;
        RECT 25.930 264.550 29.880 264.700 ;
        RECT 25.930 264.400 26.330 264.550 ;
        RECT 23.130 264.100 26.330 264.400 ;
        RECT 19.580 263.950 29.880 264.100 ;
        RECT 23.130 263.500 26.330 263.950 ;
        RECT 19.580 263.350 29.880 263.500 ;
        RECT 23.130 262.900 26.330 263.350 ;
        RECT 19.580 262.750 29.880 262.900 ;
        RECT 23.130 262.300 26.330 262.750 ;
        RECT 19.580 262.150 29.880 262.300 ;
        RECT 23.530 261.200 25.930 262.150 ;
        RECT 30.480 261.600 30.630 269.800 ;
        RECT 31.080 261.600 31.230 269.800 ;
        RECT 31.680 261.600 31.830 269.800 ;
        RECT 32.280 261.600 32.430 269.800 ;
        RECT 32.880 261.600 33.030 269.800 ;
        RECT 33.480 261.600 33.630 269.800 ;
        RECT 34.080 261.600 34.230 269.800 ;
        RECT 35.230 270.200 35.380 278.400 ;
        RECT 35.830 270.200 35.980 278.400 ;
        RECT 36.430 270.200 36.580 278.400 ;
        RECT 37.030 270.200 37.180 278.400 ;
        RECT 37.630 270.200 37.780 278.400 ;
        RECT 38.230 270.200 38.380 278.400 ;
        RECT 38.830 270.200 38.980 278.400 ;
        RECT 43.530 277.850 45.940 278.800 ;
        RECT 39.580 277.700 49.880 277.850 ;
        RECT 43.130 277.250 46.330 277.700 ;
        RECT 39.580 277.100 49.880 277.250 ;
        RECT 43.130 276.650 46.330 277.100 ;
        RECT 39.580 276.500 49.880 276.650 ;
        RECT 43.130 276.050 46.330 276.500 ;
        RECT 39.580 275.900 49.880 276.050 ;
        RECT 43.130 275.600 46.330 275.900 ;
        RECT 43.130 275.450 43.530 275.600 ;
        RECT 39.580 275.300 43.530 275.450 ;
        RECT 43.130 274.850 43.530 275.300 ;
        RECT 39.580 274.700 43.530 274.850 ;
        RECT 43.130 274.250 43.530 274.700 ;
        RECT 39.580 274.100 43.530 274.250 ;
        RECT 43.130 273.650 43.530 274.100 ;
        RECT 39.580 273.500 43.530 273.650 ;
        RECT 43.130 273.050 43.530 273.500 ;
        RECT 39.580 272.900 43.530 273.050 ;
        RECT 43.130 272.450 43.530 272.900 ;
        RECT 39.580 272.300 43.530 272.450 ;
        RECT 43.130 271.850 43.530 272.300 ;
        RECT 39.580 271.700 43.530 271.850 ;
        RECT 43.130 271.250 43.530 271.700 ;
        RECT 39.580 271.100 43.530 271.250 ;
        RECT 43.130 270.650 43.530 271.100 ;
        RECT 39.580 270.500 43.530 270.650 ;
        RECT 43.130 270.200 43.530 270.500 ;
        RECT 35.230 269.800 43.530 270.200 ;
        RECT 35.230 261.600 35.380 269.800 ;
        RECT 35.830 261.600 35.980 269.800 ;
        RECT 36.430 261.600 36.580 269.800 ;
        RECT 37.030 261.600 37.180 269.800 ;
        RECT 37.630 261.600 37.780 269.800 ;
        RECT 38.230 261.600 38.380 269.800 ;
        RECT 38.830 261.600 38.980 269.800 ;
        RECT 43.130 269.500 43.530 269.800 ;
        RECT 39.580 269.350 43.530 269.500 ;
        RECT 43.130 268.900 43.530 269.350 ;
        RECT 39.580 268.750 43.530 268.900 ;
        RECT 43.130 268.300 43.530 268.750 ;
        RECT 39.580 268.150 43.530 268.300 ;
        RECT 43.130 267.700 43.530 268.150 ;
        RECT 39.580 267.550 43.530 267.700 ;
        RECT 43.130 267.100 43.530 267.550 ;
        RECT 39.580 266.950 43.530 267.100 ;
        RECT 43.130 266.500 43.530 266.950 ;
        RECT 39.580 266.350 43.530 266.500 ;
        RECT 43.130 265.900 43.530 266.350 ;
        RECT 39.580 265.750 43.530 265.900 ;
        RECT 43.130 265.300 43.530 265.750 ;
        RECT 39.580 265.150 43.530 265.300 ;
        RECT 43.130 264.700 43.530 265.150 ;
        RECT 39.580 264.550 43.530 264.700 ;
        RECT 43.130 264.400 43.530 264.550 ;
        RECT 45.930 275.450 46.330 275.600 ;
        RECT 45.930 275.300 49.880 275.450 ;
        RECT 45.930 274.850 46.330 275.300 ;
        RECT 45.930 274.700 49.880 274.850 ;
        RECT 45.930 274.250 46.330 274.700 ;
        RECT 45.930 274.100 49.880 274.250 ;
        RECT 45.930 273.650 46.330 274.100 ;
        RECT 45.930 273.500 49.880 273.650 ;
        RECT 45.930 273.050 46.330 273.500 ;
        RECT 45.930 272.900 49.880 273.050 ;
        RECT 45.930 272.450 46.330 272.900 ;
        RECT 45.930 272.300 49.880 272.450 ;
        RECT 45.930 271.850 46.330 272.300 ;
        RECT 45.930 271.700 49.880 271.850 ;
        RECT 45.930 271.250 46.330 271.700 ;
        RECT 45.930 271.100 49.880 271.250 ;
        RECT 45.930 270.650 46.330 271.100 ;
        RECT 45.930 270.500 49.880 270.650 ;
        RECT 45.930 270.200 46.330 270.500 ;
        RECT 50.480 270.200 50.630 278.400 ;
        RECT 51.080 270.200 51.230 278.400 ;
        RECT 51.680 270.200 51.830 278.400 ;
        RECT 52.280 270.200 52.430 278.400 ;
        RECT 52.880 270.200 53.030 278.400 ;
        RECT 53.480 270.200 53.630 278.400 ;
        RECT 54.080 270.200 54.230 278.400 ;
        RECT 45.930 269.800 54.230 270.200 ;
        RECT 45.930 269.500 46.330 269.800 ;
        RECT 45.930 269.350 49.880 269.500 ;
        RECT 45.930 268.900 46.330 269.350 ;
        RECT 45.930 268.750 49.880 268.900 ;
        RECT 45.930 268.300 46.330 268.750 ;
        RECT 45.930 268.150 49.880 268.300 ;
        RECT 45.930 267.700 46.330 268.150 ;
        RECT 45.930 267.550 49.880 267.700 ;
        RECT 45.930 267.100 46.330 267.550 ;
        RECT 45.930 266.950 49.880 267.100 ;
        RECT 45.930 266.500 46.330 266.950 ;
        RECT 45.930 266.350 49.880 266.500 ;
        RECT 45.930 265.900 46.330 266.350 ;
        RECT 45.930 265.750 49.880 265.900 ;
        RECT 45.930 265.300 46.330 265.750 ;
        RECT 45.930 265.150 49.880 265.300 ;
        RECT 45.930 264.700 46.330 265.150 ;
        RECT 45.930 264.550 49.880 264.700 ;
        RECT 45.930 264.400 46.330 264.550 ;
        RECT 43.130 264.100 46.330 264.400 ;
        RECT 39.580 263.950 49.880 264.100 ;
        RECT 43.130 263.500 46.330 263.950 ;
        RECT 39.580 263.350 49.880 263.500 ;
        RECT 43.130 262.900 46.330 263.350 ;
        RECT 39.580 262.750 49.880 262.900 ;
        RECT 43.130 262.300 46.330 262.750 ;
        RECT 39.580 262.150 49.880 262.300 ;
        RECT 43.530 261.200 45.930 262.150 ;
        RECT 50.480 261.600 50.630 269.800 ;
        RECT 51.080 261.600 51.230 269.800 ;
        RECT 51.680 261.600 51.830 269.800 ;
        RECT 52.280 261.600 52.430 269.800 ;
        RECT 52.880 261.600 53.030 269.800 ;
        RECT 53.480 261.600 53.630 269.800 ;
        RECT 54.080 261.600 54.230 269.800 ;
        RECT 55.230 270.200 55.380 278.400 ;
        RECT 55.830 270.200 55.980 278.400 ;
        RECT 56.430 270.200 56.580 278.400 ;
        RECT 57.030 270.200 57.180 278.400 ;
        RECT 57.630 270.200 57.780 278.400 ;
        RECT 58.230 270.200 58.380 278.400 ;
        RECT 58.830 270.200 58.980 278.400 ;
        RECT 63.530 277.850 65.940 278.800 ;
        RECT 59.580 277.700 69.880 277.850 ;
        RECT 63.130 277.250 66.330 277.700 ;
        RECT 59.580 277.100 69.880 277.250 ;
        RECT 63.130 276.650 66.330 277.100 ;
        RECT 59.580 276.500 69.880 276.650 ;
        RECT 63.130 276.050 66.330 276.500 ;
        RECT 59.580 275.900 69.880 276.050 ;
        RECT 63.130 275.600 66.330 275.900 ;
        RECT 63.130 275.450 63.530 275.600 ;
        RECT 59.580 275.300 63.530 275.450 ;
        RECT 63.130 274.850 63.530 275.300 ;
        RECT 59.580 274.700 63.530 274.850 ;
        RECT 63.130 274.250 63.530 274.700 ;
        RECT 59.580 274.100 63.530 274.250 ;
        RECT 63.130 273.650 63.530 274.100 ;
        RECT 59.580 273.500 63.530 273.650 ;
        RECT 63.130 273.050 63.530 273.500 ;
        RECT 59.580 272.900 63.530 273.050 ;
        RECT 63.130 272.450 63.530 272.900 ;
        RECT 59.580 272.300 63.530 272.450 ;
        RECT 63.130 271.850 63.530 272.300 ;
        RECT 59.580 271.700 63.530 271.850 ;
        RECT 63.130 271.250 63.530 271.700 ;
        RECT 59.580 271.100 63.530 271.250 ;
        RECT 63.130 270.650 63.530 271.100 ;
        RECT 59.580 270.500 63.530 270.650 ;
        RECT 63.130 270.200 63.530 270.500 ;
        RECT 55.230 269.800 63.530 270.200 ;
        RECT 55.230 261.600 55.380 269.800 ;
        RECT 55.830 261.600 55.980 269.800 ;
        RECT 56.430 261.600 56.580 269.800 ;
        RECT 57.030 261.600 57.180 269.800 ;
        RECT 57.630 261.600 57.780 269.800 ;
        RECT 58.230 261.600 58.380 269.800 ;
        RECT 58.830 261.600 58.980 269.800 ;
        RECT 63.130 269.500 63.530 269.800 ;
        RECT 59.580 269.350 63.530 269.500 ;
        RECT 63.130 268.900 63.530 269.350 ;
        RECT 59.580 268.750 63.530 268.900 ;
        RECT 63.130 268.300 63.530 268.750 ;
        RECT 59.580 268.150 63.530 268.300 ;
        RECT 63.130 267.700 63.530 268.150 ;
        RECT 59.580 267.550 63.530 267.700 ;
        RECT 63.130 267.100 63.530 267.550 ;
        RECT 59.580 266.950 63.530 267.100 ;
        RECT 63.130 266.500 63.530 266.950 ;
        RECT 59.580 266.350 63.530 266.500 ;
        RECT 63.130 265.900 63.530 266.350 ;
        RECT 59.580 265.750 63.530 265.900 ;
        RECT 63.130 265.300 63.530 265.750 ;
        RECT 59.580 265.150 63.530 265.300 ;
        RECT 63.130 264.700 63.530 265.150 ;
        RECT 59.580 264.550 63.530 264.700 ;
        RECT 63.130 264.400 63.530 264.550 ;
        RECT 65.930 275.450 66.330 275.600 ;
        RECT 65.930 275.300 69.880 275.450 ;
        RECT 65.930 274.850 66.330 275.300 ;
        RECT 65.930 274.700 69.880 274.850 ;
        RECT 65.930 274.250 66.330 274.700 ;
        RECT 65.930 274.100 69.880 274.250 ;
        RECT 65.930 273.650 66.330 274.100 ;
        RECT 65.930 273.500 69.880 273.650 ;
        RECT 65.930 273.050 66.330 273.500 ;
        RECT 65.930 272.900 69.880 273.050 ;
        RECT 65.930 272.450 66.330 272.900 ;
        RECT 65.930 272.300 69.880 272.450 ;
        RECT 65.930 271.850 66.330 272.300 ;
        RECT 65.930 271.700 69.880 271.850 ;
        RECT 65.930 271.250 66.330 271.700 ;
        RECT 65.930 271.100 69.880 271.250 ;
        RECT 65.930 270.650 66.330 271.100 ;
        RECT 65.930 270.500 69.880 270.650 ;
        RECT 65.930 270.200 66.330 270.500 ;
        RECT 70.480 270.200 70.630 278.400 ;
        RECT 71.080 270.200 71.230 278.400 ;
        RECT 71.680 270.200 71.830 278.400 ;
        RECT 72.280 270.200 72.430 278.400 ;
        RECT 72.880 270.200 73.030 278.400 ;
        RECT 73.480 270.200 73.630 278.400 ;
        RECT 74.080 270.200 74.230 278.400 ;
        RECT 65.930 269.800 74.230 270.200 ;
        RECT 65.930 269.500 66.330 269.800 ;
        RECT 65.930 269.350 69.880 269.500 ;
        RECT 65.930 268.900 66.330 269.350 ;
        RECT 65.930 268.750 69.880 268.900 ;
        RECT 65.930 268.300 66.330 268.750 ;
        RECT 65.930 268.150 69.880 268.300 ;
        RECT 65.930 267.700 66.330 268.150 ;
        RECT 65.930 267.550 69.880 267.700 ;
        RECT 65.930 267.100 66.330 267.550 ;
        RECT 65.930 266.950 69.880 267.100 ;
        RECT 65.930 266.500 66.330 266.950 ;
        RECT 65.930 266.350 69.880 266.500 ;
        RECT 65.930 265.900 66.330 266.350 ;
        RECT 65.930 265.750 69.880 265.900 ;
        RECT 65.930 265.300 66.330 265.750 ;
        RECT 65.930 265.150 69.880 265.300 ;
        RECT 65.930 264.700 66.330 265.150 ;
        RECT 65.930 264.550 69.880 264.700 ;
        RECT 65.930 264.400 66.330 264.550 ;
        RECT 63.130 264.100 66.330 264.400 ;
        RECT 59.580 263.950 69.880 264.100 ;
        RECT 63.130 263.500 66.330 263.950 ;
        RECT 59.580 263.350 69.880 263.500 ;
        RECT 63.130 262.900 66.330 263.350 ;
        RECT 59.580 262.750 69.880 262.900 ;
        RECT 63.130 262.300 66.330 262.750 ;
        RECT 59.580 262.150 69.880 262.300 ;
        RECT 63.530 261.200 65.930 262.150 ;
        RECT 70.480 261.600 70.630 269.800 ;
        RECT 71.080 261.600 71.230 269.800 ;
        RECT 71.680 261.600 71.830 269.800 ;
        RECT 72.280 261.600 72.430 269.800 ;
        RECT 72.880 261.600 73.030 269.800 ;
        RECT 73.480 261.600 73.630 269.800 ;
        RECT 74.080 261.600 74.230 269.800 ;
        RECT 75.230 270.200 75.380 278.400 ;
        RECT 75.830 270.200 75.980 278.400 ;
        RECT 76.430 270.200 76.580 278.400 ;
        RECT 77.030 270.200 77.180 278.400 ;
        RECT 77.630 270.200 77.780 278.400 ;
        RECT 78.230 270.200 78.380 278.400 ;
        RECT 78.830 270.200 78.980 278.400 ;
        RECT 83.530 277.850 85.940 278.800 ;
        RECT 79.580 277.700 89.880 277.850 ;
        RECT 83.130 277.250 86.330 277.700 ;
        RECT 79.580 277.100 89.880 277.250 ;
        RECT 83.130 276.650 86.330 277.100 ;
        RECT 79.580 276.500 89.880 276.650 ;
        RECT 83.130 276.050 86.330 276.500 ;
        RECT 79.580 275.900 89.880 276.050 ;
        RECT 83.130 275.600 86.330 275.900 ;
        RECT 83.130 275.450 83.530 275.600 ;
        RECT 79.580 275.300 83.530 275.450 ;
        RECT 83.130 274.850 83.530 275.300 ;
        RECT 79.580 274.700 83.530 274.850 ;
        RECT 83.130 274.250 83.530 274.700 ;
        RECT 79.580 274.100 83.530 274.250 ;
        RECT 83.130 273.650 83.530 274.100 ;
        RECT 79.580 273.500 83.530 273.650 ;
        RECT 83.130 273.050 83.530 273.500 ;
        RECT 79.580 272.900 83.530 273.050 ;
        RECT 83.130 272.450 83.530 272.900 ;
        RECT 79.580 272.300 83.530 272.450 ;
        RECT 83.130 271.850 83.530 272.300 ;
        RECT 79.580 271.700 83.530 271.850 ;
        RECT 83.130 271.250 83.530 271.700 ;
        RECT 79.580 271.100 83.530 271.250 ;
        RECT 83.130 270.650 83.530 271.100 ;
        RECT 79.580 270.500 83.530 270.650 ;
        RECT 83.130 270.200 83.530 270.500 ;
        RECT 75.230 269.800 83.530 270.200 ;
        RECT 75.230 261.600 75.380 269.800 ;
        RECT 75.830 261.600 75.980 269.800 ;
        RECT 76.430 261.600 76.580 269.800 ;
        RECT 77.030 261.600 77.180 269.800 ;
        RECT 77.630 261.600 77.780 269.800 ;
        RECT 78.230 261.600 78.380 269.800 ;
        RECT 78.830 261.600 78.980 269.800 ;
        RECT 83.130 269.500 83.530 269.800 ;
        RECT 79.580 269.350 83.530 269.500 ;
        RECT 83.130 268.900 83.530 269.350 ;
        RECT 79.580 268.750 83.530 268.900 ;
        RECT 83.130 268.300 83.530 268.750 ;
        RECT 79.580 268.150 83.530 268.300 ;
        RECT 83.130 267.700 83.530 268.150 ;
        RECT 79.580 267.550 83.530 267.700 ;
        RECT 83.130 267.100 83.530 267.550 ;
        RECT 79.580 266.950 83.530 267.100 ;
        RECT 83.130 266.500 83.530 266.950 ;
        RECT 79.580 266.350 83.530 266.500 ;
        RECT 83.130 265.900 83.530 266.350 ;
        RECT 79.580 265.750 83.530 265.900 ;
        RECT 83.130 265.300 83.530 265.750 ;
        RECT 79.580 265.150 83.530 265.300 ;
        RECT 83.130 264.700 83.530 265.150 ;
        RECT 79.580 264.550 83.530 264.700 ;
        RECT 83.130 264.400 83.530 264.550 ;
        RECT 85.930 275.450 86.330 275.600 ;
        RECT 85.930 275.300 89.880 275.450 ;
        RECT 85.930 274.850 86.330 275.300 ;
        RECT 85.930 274.700 89.880 274.850 ;
        RECT 85.930 274.250 86.330 274.700 ;
        RECT 85.930 274.100 89.880 274.250 ;
        RECT 85.930 273.650 86.330 274.100 ;
        RECT 85.930 273.500 89.880 273.650 ;
        RECT 85.930 273.050 86.330 273.500 ;
        RECT 85.930 272.900 89.880 273.050 ;
        RECT 85.930 272.450 86.330 272.900 ;
        RECT 85.930 272.300 89.880 272.450 ;
        RECT 85.930 271.850 86.330 272.300 ;
        RECT 85.930 271.700 89.880 271.850 ;
        RECT 85.930 271.250 86.330 271.700 ;
        RECT 85.930 271.100 89.880 271.250 ;
        RECT 85.930 270.650 86.330 271.100 ;
        RECT 85.930 270.500 89.880 270.650 ;
        RECT 85.930 270.200 86.330 270.500 ;
        RECT 90.480 270.200 90.630 278.400 ;
        RECT 91.080 270.200 91.230 278.400 ;
        RECT 91.680 270.200 91.830 278.400 ;
        RECT 92.280 270.200 92.430 278.400 ;
        RECT 92.880 270.200 93.030 278.400 ;
        RECT 93.480 270.200 93.630 278.400 ;
        RECT 94.080 270.200 94.230 278.400 ;
        RECT 85.930 269.800 94.230 270.200 ;
        RECT 85.930 269.500 86.330 269.800 ;
        RECT 85.930 269.350 89.880 269.500 ;
        RECT 85.930 268.900 86.330 269.350 ;
        RECT 85.930 268.750 89.880 268.900 ;
        RECT 85.930 268.300 86.330 268.750 ;
        RECT 85.930 268.150 89.880 268.300 ;
        RECT 85.930 267.700 86.330 268.150 ;
        RECT 85.930 267.550 89.880 267.700 ;
        RECT 85.930 267.100 86.330 267.550 ;
        RECT 85.930 266.950 89.880 267.100 ;
        RECT 85.930 266.500 86.330 266.950 ;
        RECT 85.930 266.350 89.880 266.500 ;
        RECT 85.930 265.900 86.330 266.350 ;
        RECT 85.930 265.750 89.880 265.900 ;
        RECT 85.930 265.300 86.330 265.750 ;
        RECT 85.930 265.150 89.880 265.300 ;
        RECT 85.930 264.700 86.330 265.150 ;
        RECT 85.930 264.550 89.880 264.700 ;
        RECT 85.930 264.400 86.330 264.550 ;
        RECT 83.130 264.100 86.330 264.400 ;
        RECT 79.580 263.950 89.880 264.100 ;
        RECT 83.130 263.500 86.330 263.950 ;
        RECT 79.580 263.350 89.880 263.500 ;
        RECT 83.130 262.900 86.330 263.350 ;
        RECT 79.580 262.750 89.880 262.900 ;
        RECT 83.130 262.300 86.330 262.750 ;
        RECT 79.580 262.150 89.880 262.300 ;
        RECT 83.530 261.200 85.930 262.150 ;
        RECT 90.480 261.600 90.630 269.800 ;
        RECT 91.080 261.600 91.230 269.800 ;
        RECT 91.680 261.600 91.830 269.800 ;
        RECT 92.280 261.600 92.430 269.800 ;
        RECT 92.880 261.600 93.030 269.800 ;
        RECT 93.480 261.600 93.630 269.800 ;
        RECT 94.080 261.600 94.230 269.800 ;
        RECT 95.230 270.200 95.380 278.400 ;
        RECT 95.830 270.200 95.980 278.400 ;
        RECT 96.430 270.200 96.580 278.400 ;
        RECT 97.030 270.200 97.180 278.400 ;
        RECT 97.630 270.200 97.780 278.400 ;
        RECT 98.230 270.200 98.380 278.400 ;
        RECT 98.830 270.200 98.980 278.400 ;
        RECT 103.530 277.850 104.730 278.800 ;
        RECT 99.580 277.700 104.730 277.850 ;
        RECT 103.130 277.250 104.730 277.700 ;
        RECT 99.580 277.100 104.730 277.250 ;
        RECT 103.130 276.650 104.730 277.100 ;
        RECT 99.580 276.500 104.730 276.650 ;
        RECT 103.130 276.050 104.730 276.500 ;
        RECT 105.135 276.085 107.135 277.360 ;
        RECT 99.580 275.900 104.730 276.050 ;
        RECT 103.130 275.600 104.730 275.900 ;
        RECT 103.130 275.450 103.530 275.600 ;
        RECT 99.580 275.300 103.530 275.450 ;
        RECT 103.130 274.850 103.530 275.300 ;
        RECT 99.580 274.700 103.530 274.850 ;
        RECT 103.130 274.250 103.530 274.700 ;
        RECT 99.580 274.100 103.530 274.250 ;
        RECT 103.130 273.650 103.530 274.100 ;
        RECT 99.580 273.500 103.530 273.650 ;
        RECT 103.130 273.050 103.530 273.500 ;
        RECT 99.580 272.900 103.530 273.050 ;
        RECT 103.130 272.450 103.530 272.900 ;
        RECT 99.580 272.300 103.530 272.450 ;
        RECT 103.130 271.850 103.530 272.300 ;
        RECT 99.580 271.700 103.530 271.850 ;
        RECT 103.130 271.250 103.530 271.700 ;
        RECT 99.580 271.100 103.530 271.250 ;
        RECT 103.130 270.650 103.530 271.100 ;
        RECT 99.580 270.500 103.530 270.650 ;
        RECT 103.130 270.200 103.530 270.500 ;
        RECT 95.230 269.800 103.530 270.200 ;
        RECT 95.230 261.600 95.380 269.800 ;
        RECT 95.830 261.600 95.980 269.800 ;
        RECT 96.430 261.600 96.580 269.800 ;
        RECT 97.030 261.600 97.180 269.800 ;
        RECT 97.630 261.600 97.780 269.800 ;
        RECT 98.230 261.600 98.380 269.800 ;
        RECT 98.830 261.600 98.980 269.800 ;
        RECT 103.130 269.500 103.530 269.800 ;
        RECT 99.580 269.350 103.530 269.500 ;
        RECT 103.130 268.900 103.530 269.350 ;
        RECT 99.580 268.750 103.530 268.900 ;
        RECT 103.130 268.300 103.530 268.750 ;
        RECT 99.580 268.150 103.530 268.300 ;
        RECT 103.130 267.700 103.530 268.150 ;
        RECT 99.580 267.550 103.530 267.700 ;
        RECT 103.130 267.100 103.530 267.550 ;
        RECT 99.580 266.950 103.530 267.100 ;
        RECT 103.130 266.500 103.530 266.950 ;
        RECT 99.580 266.350 103.530 266.500 ;
        RECT 103.130 265.900 103.530 266.350 ;
        RECT 99.580 265.750 103.530 265.900 ;
        RECT 103.130 265.300 103.530 265.750 ;
        RECT 99.580 265.150 103.530 265.300 ;
        RECT 103.130 264.700 103.530 265.150 ;
        RECT 99.580 264.550 103.530 264.700 ;
        RECT 103.130 264.400 103.530 264.550 ;
        RECT 103.130 264.100 104.730 264.400 ;
        RECT 99.580 263.950 104.730 264.100 ;
        RECT 103.130 263.500 104.730 263.950 ;
        RECT 99.580 263.350 104.730 263.500 ;
        RECT 103.130 262.900 104.730 263.350 ;
        RECT 99.580 262.750 104.730 262.900 ;
        RECT 103.130 262.300 104.730 262.750 ;
        RECT 99.580 262.150 104.730 262.300 ;
        RECT 103.530 261.200 104.730 262.150 ;
        RECT 105.140 261.725 107.140 263.000 ;
        RECT 4.730 258.800 9.130 261.200 ;
        RECT 20.330 258.800 29.130 261.200 ;
        RECT 40.330 258.800 49.130 261.200 ;
        RECT 60.330 258.800 69.130 261.200 ;
        RECT 80.330 258.800 89.130 261.200 ;
        RECT 100.330 258.800 104.730 261.200 ;
        RECT 4.730 257.850 5.940 258.800 ;
        RECT 2.315 256.570 4.320 257.845 ;
        RECT 4.730 257.700 9.880 257.850 ;
        RECT 4.730 257.250 6.330 257.700 ;
        RECT 4.730 257.100 9.880 257.250 ;
        RECT 4.730 256.650 6.330 257.100 ;
        RECT 4.730 256.500 9.880 256.650 ;
        RECT 4.730 256.050 6.330 256.500 ;
        RECT 4.730 255.900 9.880 256.050 ;
        RECT 4.730 255.600 6.330 255.900 ;
        RECT 2.315 253.250 4.315 255.545 ;
        RECT 5.930 255.450 6.330 255.600 ;
        RECT 5.930 255.300 9.880 255.450 ;
        RECT 5.930 254.850 6.330 255.300 ;
        RECT 5.930 254.700 9.880 254.850 ;
        RECT 5.930 254.250 6.330 254.700 ;
        RECT 5.930 254.100 9.880 254.250 ;
        RECT 5.930 253.650 6.330 254.100 ;
        RECT 5.930 253.500 9.880 253.650 ;
        RECT 5.930 253.050 6.330 253.500 ;
        RECT 5.930 252.900 9.880 253.050 ;
        RECT 5.930 252.450 6.330 252.900 ;
        RECT 5.930 252.300 9.880 252.450 ;
        RECT 5.930 251.850 6.330 252.300 ;
        RECT 5.930 251.700 9.880 251.850 ;
        RECT 5.930 251.250 6.330 251.700 ;
        RECT 5.930 251.100 9.880 251.250 ;
        RECT 5.930 250.650 6.330 251.100 ;
        RECT 5.930 250.500 9.880 250.650 ;
        RECT 5.930 250.200 6.330 250.500 ;
        RECT 10.480 250.200 10.630 258.400 ;
        RECT 11.080 250.200 11.230 258.400 ;
        RECT 11.680 250.200 11.830 258.400 ;
        RECT 12.280 250.200 12.430 258.400 ;
        RECT 12.880 250.200 13.030 258.400 ;
        RECT 13.480 250.200 13.630 258.400 ;
        RECT 14.080 250.200 14.230 258.400 ;
        RECT 5.930 249.800 14.230 250.200 ;
        RECT 5.930 249.500 6.330 249.800 ;
        RECT 5.930 249.350 9.880 249.500 ;
        RECT 5.930 248.900 6.330 249.350 ;
        RECT 5.930 248.750 9.880 248.900 ;
        RECT 5.930 248.300 6.330 248.750 ;
        RECT 5.930 248.150 9.880 248.300 ;
        RECT 5.930 247.700 6.330 248.150 ;
        RECT 5.930 247.550 9.880 247.700 ;
        RECT 5.930 247.100 6.330 247.550 ;
        RECT 5.930 246.950 9.880 247.100 ;
        RECT 2.315 244.455 4.315 246.750 ;
        RECT 5.930 246.500 6.330 246.950 ;
        RECT 5.930 246.350 9.880 246.500 ;
        RECT 5.930 245.900 6.330 246.350 ;
        RECT 5.930 245.750 9.880 245.900 ;
        RECT 5.930 245.300 6.330 245.750 ;
        RECT 5.930 245.150 9.880 245.300 ;
        RECT 5.930 244.700 6.330 245.150 ;
        RECT 5.930 244.550 9.880 244.700 ;
        RECT 5.930 244.400 6.330 244.550 ;
        RECT 4.730 244.100 6.330 244.400 ;
        RECT 4.730 243.950 9.880 244.100 ;
        RECT 2.315 242.460 4.320 243.735 ;
        RECT 4.730 243.500 6.330 243.950 ;
        RECT 4.730 243.350 9.880 243.500 ;
        RECT 4.730 242.900 6.330 243.350 ;
        RECT 4.730 242.750 9.880 242.900 ;
        RECT 4.730 242.300 6.330 242.750 ;
        RECT 4.730 242.150 9.880 242.300 ;
        RECT 4.730 241.200 5.930 242.150 ;
        RECT 10.480 241.600 10.630 249.800 ;
        RECT 11.080 241.600 11.230 249.800 ;
        RECT 11.680 241.600 11.830 249.800 ;
        RECT 12.280 241.600 12.430 249.800 ;
        RECT 12.880 241.600 13.030 249.800 ;
        RECT 13.480 241.600 13.630 249.800 ;
        RECT 14.080 241.600 14.230 249.800 ;
        RECT 15.230 250.200 15.380 258.400 ;
        RECT 15.830 250.200 15.980 258.400 ;
        RECT 16.430 250.200 16.580 258.400 ;
        RECT 17.030 250.200 17.180 258.400 ;
        RECT 17.630 250.200 17.780 258.400 ;
        RECT 18.230 250.200 18.380 258.400 ;
        RECT 18.830 250.200 18.980 258.400 ;
        RECT 23.530 257.850 25.940 258.800 ;
        RECT 19.580 257.700 29.880 257.850 ;
        RECT 23.130 257.250 26.330 257.700 ;
        RECT 19.580 257.100 29.880 257.250 ;
        RECT 23.130 256.650 26.330 257.100 ;
        RECT 19.580 256.500 29.880 256.650 ;
        RECT 23.130 256.050 26.330 256.500 ;
        RECT 19.580 255.900 29.880 256.050 ;
        RECT 23.130 255.600 26.330 255.900 ;
        RECT 23.130 255.450 23.530 255.600 ;
        RECT 19.580 255.300 23.530 255.450 ;
        RECT 23.130 254.850 23.530 255.300 ;
        RECT 19.580 254.700 23.530 254.850 ;
        RECT 23.130 254.250 23.530 254.700 ;
        RECT 19.580 254.100 23.530 254.250 ;
        RECT 23.130 253.650 23.530 254.100 ;
        RECT 19.580 253.500 23.530 253.650 ;
        RECT 23.130 253.050 23.530 253.500 ;
        RECT 19.580 252.900 23.530 253.050 ;
        RECT 23.130 252.450 23.530 252.900 ;
        RECT 19.580 252.300 23.530 252.450 ;
        RECT 23.130 251.850 23.530 252.300 ;
        RECT 19.580 251.700 23.530 251.850 ;
        RECT 23.130 251.250 23.530 251.700 ;
        RECT 19.580 251.100 23.530 251.250 ;
        RECT 23.130 250.650 23.530 251.100 ;
        RECT 19.580 250.500 23.530 250.650 ;
        RECT 23.130 250.200 23.530 250.500 ;
        RECT 15.230 249.800 23.530 250.200 ;
        RECT 15.230 241.600 15.380 249.800 ;
        RECT 15.830 241.600 15.980 249.800 ;
        RECT 16.430 241.600 16.580 249.800 ;
        RECT 17.030 241.600 17.180 249.800 ;
        RECT 17.630 241.600 17.780 249.800 ;
        RECT 18.230 241.600 18.380 249.800 ;
        RECT 18.830 241.600 18.980 249.800 ;
        RECT 23.130 249.500 23.530 249.800 ;
        RECT 19.580 249.350 23.530 249.500 ;
        RECT 23.130 248.900 23.530 249.350 ;
        RECT 19.580 248.750 23.530 248.900 ;
        RECT 23.130 248.300 23.530 248.750 ;
        RECT 19.580 248.150 23.530 248.300 ;
        RECT 23.130 247.700 23.530 248.150 ;
        RECT 19.580 247.550 23.530 247.700 ;
        RECT 23.130 247.100 23.530 247.550 ;
        RECT 19.580 246.950 23.530 247.100 ;
        RECT 23.130 246.500 23.530 246.950 ;
        RECT 19.580 246.350 23.530 246.500 ;
        RECT 23.130 245.900 23.530 246.350 ;
        RECT 19.580 245.750 23.530 245.900 ;
        RECT 23.130 245.300 23.530 245.750 ;
        RECT 19.580 245.150 23.530 245.300 ;
        RECT 23.130 244.700 23.530 245.150 ;
        RECT 19.580 244.550 23.530 244.700 ;
        RECT 23.130 244.400 23.530 244.550 ;
        RECT 25.930 255.450 26.330 255.600 ;
        RECT 25.930 255.300 29.880 255.450 ;
        RECT 25.930 254.850 26.330 255.300 ;
        RECT 25.930 254.700 29.880 254.850 ;
        RECT 25.930 254.250 26.330 254.700 ;
        RECT 25.930 254.100 29.880 254.250 ;
        RECT 25.930 253.650 26.330 254.100 ;
        RECT 25.930 253.500 29.880 253.650 ;
        RECT 25.930 253.050 26.330 253.500 ;
        RECT 25.930 252.900 29.880 253.050 ;
        RECT 25.930 252.450 26.330 252.900 ;
        RECT 25.930 252.300 29.880 252.450 ;
        RECT 25.930 251.850 26.330 252.300 ;
        RECT 25.930 251.700 29.880 251.850 ;
        RECT 25.930 251.250 26.330 251.700 ;
        RECT 25.930 251.100 29.880 251.250 ;
        RECT 25.930 250.650 26.330 251.100 ;
        RECT 25.930 250.500 29.880 250.650 ;
        RECT 25.930 250.200 26.330 250.500 ;
        RECT 30.480 250.200 30.630 258.400 ;
        RECT 31.080 250.200 31.230 258.400 ;
        RECT 31.680 250.200 31.830 258.400 ;
        RECT 32.280 250.200 32.430 258.400 ;
        RECT 32.880 250.200 33.030 258.400 ;
        RECT 33.480 250.200 33.630 258.400 ;
        RECT 34.080 250.200 34.230 258.400 ;
        RECT 25.930 249.800 34.230 250.200 ;
        RECT 25.930 249.500 26.330 249.800 ;
        RECT 25.930 249.350 29.880 249.500 ;
        RECT 25.930 248.900 26.330 249.350 ;
        RECT 25.930 248.750 29.880 248.900 ;
        RECT 25.930 248.300 26.330 248.750 ;
        RECT 25.930 248.150 29.880 248.300 ;
        RECT 25.930 247.700 26.330 248.150 ;
        RECT 25.930 247.550 29.880 247.700 ;
        RECT 25.930 247.100 26.330 247.550 ;
        RECT 25.930 246.950 29.880 247.100 ;
        RECT 25.930 246.500 26.330 246.950 ;
        RECT 25.930 246.350 29.880 246.500 ;
        RECT 25.930 245.900 26.330 246.350 ;
        RECT 25.930 245.750 29.880 245.900 ;
        RECT 25.930 245.300 26.330 245.750 ;
        RECT 25.930 245.150 29.880 245.300 ;
        RECT 25.930 244.700 26.330 245.150 ;
        RECT 25.930 244.550 29.880 244.700 ;
        RECT 25.930 244.400 26.330 244.550 ;
        RECT 23.130 244.100 26.330 244.400 ;
        RECT 19.580 243.950 29.880 244.100 ;
        RECT 23.130 243.500 26.330 243.950 ;
        RECT 19.580 243.350 29.880 243.500 ;
        RECT 23.130 242.900 26.330 243.350 ;
        RECT 19.580 242.750 29.880 242.900 ;
        RECT 23.130 242.300 26.330 242.750 ;
        RECT 19.580 242.150 29.880 242.300 ;
        RECT 23.530 241.200 25.930 242.150 ;
        RECT 30.480 241.600 30.630 249.800 ;
        RECT 31.080 241.600 31.230 249.800 ;
        RECT 31.680 241.600 31.830 249.800 ;
        RECT 32.280 241.600 32.430 249.800 ;
        RECT 32.880 241.600 33.030 249.800 ;
        RECT 33.480 241.600 33.630 249.800 ;
        RECT 34.080 241.600 34.230 249.800 ;
        RECT 35.230 250.200 35.380 258.400 ;
        RECT 35.830 250.200 35.980 258.400 ;
        RECT 36.430 250.200 36.580 258.400 ;
        RECT 37.030 250.200 37.180 258.400 ;
        RECT 37.630 250.200 37.780 258.400 ;
        RECT 38.230 250.200 38.380 258.400 ;
        RECT 38.830 250.200 38.980 258.400 ;
        RECT 43.530 257.850 45.940 258.800 ;
        RECT 39.580 257.700 49.880 257.850 ;
        RECT 43.130 257.250 46.330 257.700 ;
        RECT 39.580 257.100 49.880 257.250 ;
        RECT 43.130 256.650 46.330 257.100 ;
        RECT 39.580 256.500 49.880 256.650 ;
        RECT 43.130 256.050 46.330 256.500 ;
        RECT 39.580 255.900 49.880 256.050 ;
        RECT 43.130 255.600 46.330 255.900 ;
        RECT 43.130 255.450 43.530 255.600 ;
        RECT 39.580 255.300 43.530 255.450 ;
        RECT 43.130 254.850 43.530 255.300 ;
        RECT 39.580 254.700 43.530 254.850 ;
        RECT 43.130 254.250 43.530 254.700 ;
        RECT 39.580 254.100 43.530 254.250 ;
        RECT 43.130 253.650 43.530 254.100 ;
        RECT 39.580 253.500 43.530 253.650 ;
        RECT 43.130 253.050 43.530 253.500 ;
        RECT 39.580 252.900 43.530 253.050 ;
        RECT 43.130 252.450 43.530 252.900 ;
        RECT 39.580 252.300 43.530 252.450 ;
        RECT 43.130 251.850 43.530 252.300 ;
        RECT 39.580 251.700 43.530 251.850 ;
        RECT 43.130 251.250 43.530 251.700 ;
        RECT 39.580 251.100 43.530 251.250 ;
        RECT 43.130 250.650 43.530 251.100 ;
        RECT 39.580 250.500 43.530 250.650 ;
        RECT 43.130 250.200 43.530 250.500 ;
        RECT 35.230 249.800 43.530 250.200 ;
        RECT 35.230 241.600 35.380 249.800 ;
        RECT 35.830 241.600 35.980 249.800 ;
        RECT 36.430 241.600 36.580 249.800 ;
        RECT 37.030 241.600 37.180 249.800 ;
        RECT 37.630 241.600 37.780 249.800 ;
        RECT 38.230 241.600 38.380 249.800 ;
        RECT 38.830 241.600 38.980 249.800 ;
        RECT 43.130 249.500 43.530 249.800 ;
        RECT 39.580 249.350 43.530 249.500 ;
        RECT 43.130 248.900 43.530 249.350 ;
        RECT 39.580 248.750 43.530 248.900 ;
        RECT 43.130 248.300 43.530 248.750 ;
        RECT 39.580 248.150 43.530 248.300 ;
        RECT 43.130 247.700 43.530 248.150 ;
        RECT 39.580 247.550 43.530 247.700 ;
        RECT 43.130 247.100 43.530 247.550 ;
        RECT 39.580 246.950 43.530 247.100 ;
        RECT 43.130 246.500 43.530 246.950 ;
        RECT 39.580 246.350 43.530 246.500 ;
        RECT 43.130 245.900 43.530 246.350 ;
        RECT 39.580 245.750 43.530 245.900 ;
        RECT 43.130 245.300 43.530 245.750 ;
        RECT 39.580 245.150 43.530 245.300 ;
        RECT 43.130 244.700 43.530 245.150 ;
        RECT 39.580 244.550 43.530 244.700 ;
        RECT 43.130 244.400 43.530 244.550 ;
        RECT 45.930 255.450 46.330 255.600 ;
        RECT 45.930 255.300 49.880 255.450 ;
        RECT 45.930 254.850 46.330 255.300 ;
        RECT 45.930 254.700 49.880 254.850 ;
        RECT 45.930 254.250 46.330 254.700 ;
        RECT 45.930 254.100 49.880 254.250 ;
        RECT 45.930 253.650 46.330 254.100 ;
        RECT 45.930 253.500 49.880 253.650 ;
        RECT 45.930 253.050 46.330 253.500 ;
        RECT 45.930 252.900 49.880 253.050 ;
        RECT 45.930 252.450 46.330 252.900 ;
        RECT 45.930 252.300 49.880 252.450 ;
        RECT 45.930 251.850 46.330 252.300 ;
        RECT 45.930 251.700 49.880 251.850 ;
        RECT 45.930 251.250 46.330 251.700 ;
        RECT 45.930 251.100 49.880 251.250 ;
        RECT 45.930 250.650 46.330 251.100 ;
        RECT 45.930 250.500 49.880 250.650 ;
        RECT 45.930 250.200 46.330 250.500 ;
        RECT 50.480 250.200 50.630 258.400 ;
        RECT 51.080 250.200 51.230 258.400 ;
        RECT 51.680 250.200 51.830 258.400 ;
        RECT 52.280 250.200 52.430 258.400 ;
        RECT 52.880 250.200 53.030 258.400 ;
        RECT 53.480 250.200 53.630 258.400 ;
        RECT 54.080 250.200 54.230 258.400 ;
        RECT 45.930 249.800 54.230 250.200 ;
        RECT 45.930 249.500 46.330 249.800 ;
        RECT 45.930 249.350 49.880 249.500 ;
        RECT 45.930 248.900 46.330 249.350 ;
        RECT 45.930 248.750 49.880 248.900 ;
        RECT 45.930 248.300 46.330 248.750 ;
        RECT 45.930 248.150 49.880 248.300 ;
        RECT 45.930 247.700 46.330 248.150 ;
        RECT 45.930 247.550 49.880 247.700 ;
        RECT 45.930 247.100 46.330 247.550 ;
        RECT 45.930 246.950 49.880 247.100 ;
        RECT 45.930 246.500 46.330 246.950 ;
        RECT 45.930 246.350 49.880 246.500 ;
        RECT 45.930 245.900 46.330 246.350 ;
        RECT 45.930 245.750 49.880 245.900 ;
        RECT 45.930 245.300 46.330 245.750 ;
        RECT 45.930 245.150 49.880 245.300 ;
        RECT 45.930 244.700 46.330 245.150 ;
        RECT 45.930 244.550 49.880 244.700 ;
        RECT 45.930 244.400 46.330 244.550 ;
        RECT 43.130 244.100 46.330 244.400 ;
        RECT 39.580 243.950 49.880 244.100 ;
        RECT 43.130 243.500 46.330 243.950 ;
        RECT 39.580 243.350 49.880 243.500 ;
        RECT 43.130 242.900 46.330 243.350 ;
        RECT 39.580 242.750 49.880 242.900 ;
        RECT 43.130 242.300 46.330 242.750 ;
        RECT 39.580 242.150 49.880 242.300 ;
        RECT 43.530 241.200 45.930 242.150 ;
        RECT 50.480 241.600 50.630 249.800 ;
        RECT 51.080 241.600 51.230 249.800 ;
        RECT 51.680 241.600 51.830 249.800 ;
        RECT 52.280 241.600 52.430 249.800 ;
        RECT 52.880 241.600 53.030 249.800 ;
        RECT 53.480 241.600 53.630 249.800 ;
        RECT 54.080 241.600 54.230 249.800 ;
        RECT 55.230 250.200 55.380 258.400 ;
        RECT 55.830 250.200 55.980 258.400 ;
        RECT 56.430 250.200 56.580 258.400 ;
        RECT 57.030 250.200 57.180 258.400 ;
        RECT 57.630 250.200 57.780 258.400 ;
        RECT 58.230 250.200 58.380 258.400 ;
        RECT 58.830 250.200 58.980 258.400 ;
        RECT 63.530 257.850 65.940 258.800 ;
        RECT 59.580 257.700 69.880 257.850 ;
        RECT 63.130 257.250 66.330 257.700 ;
        RECT 59.580 257.100 69.880 257.250 ;
        RECT 63.130 256.650 66.330 257.100 ;
        RECT 59.580 256.500 69.880 256.650 ;
        RECT 63.130 256.050 66.330 256.500 ;
        RECT 59.580 255.900 69.880 256.050 ;
        RECT 63.130 255.600 66.330 255.900 ;
        RECT 63.130 255.450 63.530 255.600 ;
        RECT 59.580 255.300 63.530 255.450 ;
        RECT 63.130 254.850 63.530 255.300 ;
        RECT 59.580 254.700 63.530 254.850 ;
        RECT 63.130 254.250 63.530 254.700 ;
        RECT 59.580 254.100 63.530 254.250 ;
        RECT 63.130 253.650 63.530 254.100 ;
        RECT 59.580 253.500 63.530 253.650 ;
        RECT 63.130 253.050 63.530 253.500 ;
        RECT 59.580 252.900 63.530 253.050 ;
        RECT 63.130 252.450 63.530 252.900 ;
        RECT 59.580 252.300 63.530 252.450 ;
        RECT 63.130 251.850 63.530 252.300 ;
        RECT 59.580 251.700 63.530 251.850 ;
        RECT 63.130 251.250 63.530 251.700 ;
        RECT 59.580 251.100 63.530 251.250 ;
        RECT 63.130 250.650 63.530 251.100 ;
        RECT 59.580 250.500 63.530 250.650 ;
        RECT 63.130 250.200 63.530 250.500 ;
        RECT 55.230 249.800 63.530 250.200 ;
        RECT 55.230 241.600 55.380 249.800 ;
        RECT 55.830 241.600 55.980 249.800 ;
        RECT 56.430 241.600 56.580 249.800 ;
        RECT 57.030 241.600 57.180 249.800 ;
        RECT 57.630 241.600 57.780 249.800 ;
        RECT 58.230 241.600 58.380 249.800 ;
        RECT 58.830 241.600 58.980 249.800 ;
        RECT 63.130 249.500 63.530 249.800 ;
        RECT 59.580 249.350 63.530 249.500 ;
        RECT 63.130 248.900 63.530 249.350 ;
        RECT 59.580 248.750 63.530 248.900 ;
        RECT 63.130 248.300 63.530 248.750 ;
        RECT 59.580 248.150 63.530 248.300 ;
        RECT 63.130 247.700 63.530 248.150 ;
        RECT 59.580 247.550 63.530 247.700 ;
        RECT 63.130 247.100 63.530 247.550 ;
        RECT 59.580 246.950 63.530 247.100 ;
        RECT 63.130 246.500 63.530 246.950 ;
        RECT 59.580 246.350 63.530 246.500 ;
        RECT 63.130 245.900 63.530 246.350 ;
        RECT 59.580 245.750 63.530 245.900 ;
        RECT 63.130 245.300 63.530 245.750 ;
        RECT 59.580 245.150 63.530 245.300 ;
        RECT 63.130 244.700 63.530 245.150 ;
        RECT 59.580 244.550 63.530 244.700 ;
        RECT 63.130 244.400 63.530 244.550 ;
        RECT 65.930 255.450 66.330 255.600 ;
        RECT 65.930 255.300 69.880 255.450 ;
        RECT 65.930 254.850 66.330 255.300 ;
        RECT 65.930 254.700 69.880 254.850 ;
        RECT 65.930 254.250 66.330 254.700 ;
        RECT 65.930 254.100 69.880 254.250 ;
        RECT 65.930 253.650 66.330 254.100 ;
        RECT 65.930 253.500 69.880 253.650 ;
        RECT 65.930 253.050 66.330 253.500 ;
        RECT 65.930 252.900 69.880 253.050 ;
        RECT 65.930 252.450 66.330 252.900 ;
        RECT 65.930 252.300 69.880 252.450 ;
        RECT 65.930 251.850 66.330 252.300 ;
        RECT 65.930 251.700 69.880 251.850 ;
        RECT 65.930 251.250 66.330 251.700 ;
        RECT 65.930 251.100 69.880 251.250 ;
        RECT 65.930 250.650 66.330 251.100 ;
        RECT 65.930 250.500 69.880 250.650 ;
        RECT 65.930 250.200 66.330 250.500 ;
        RECT 70.480 250.200 70.630 258.400 ;
        RECT 71.080 250.200 71.230 258.400 ;
        RECT 71.680 250.200 71.830 258.400 ;
        RECT 72.280 250.200 72.430 258.400 ;
        RECT 72.880 250.200 73.030 258.400 ;
        RECT 73.480 250.200 73.630 258.400 ;
        RECT 74.080 250.200 74.230 258.400 ;
        RECT 65.930 249.800 74.230 250.200 ;
        RECT 65.930 249.500 66.330 249.800 ;
        RECT 65.930 249.350 69.880 249.500 ;
        RECT 65.930 248.900 66.330 249.350 ;
        RECT 65.930 248.750 69.880 248.900 ;
        RECT 65.930 248.300 66.330 248.750 ;
        RECT 65.930 248.150 69.880 248.300 ;
        RECT 65.930 247.700 66.330 248.150 ;
        RECT 65.930 247.550 69.880 247.700 ;
        RECT 65.930 247.100 66.330 247.550 ;
        RECT 65.930 246.950 69.880 247.100 ;
        RECT 65.930 246.500 66.330 246.950 ;
        RECT 65.930 246.350 69.880 246.500 ;
        RECT 65.930 245.900 66.330 246.350 ;
        RECT 65.930 245.750 69.880 245.900 ;
        RECT 65.930 245.300 66.330 245.750 ;
        RECT 65.930 245.150 69.880 245.300 ;
        RECT 65.930 244.700 66.330 245.150 ;
        RECT 65.930 244.550 69.880 244.700 ;
        RECT 65.930 244.400 66.330 244.550 ;
        RECT 63.130 244.100 66.330 244.400 ;
        RECT 59.580 243.950 69.880 244.100 ;
        RECT 63.130 243.500 66.330 243.950 ;
        RECT 59.580 243.350 69.880 243.500 ;
        RECT 63.130 242.900 66.330 243.350 ;
        RECT 59.580 242.750 69.880 242.900 ;
        RECT 63.130 242.300 66.330 242.750 ;
        RECT 59.580 242.150 69.880 242.300 ;
        RECT 63.530 241.200 65.930 242.150 ;
        RECT 70.480 241.600 70.630 249.800 ;
        RECT 71.080 241.600 71.230 249.800 ;
        RECT 71.680 241.600 71.830 249.800 ;
        RECT 72.280 241.600 72.430 249.800 ;
        RECT 72.880 241.600 73.030 249.800 ;
        RECT 73.480 241.600 73.630 249.800 ;
        RECT 74.080 241.600 74.230 249.800 ;
        RECT 75.230 250.200 75.380 258.400 ;
        RECT 75.830 250.200 75.980 258.400 ;
        RECT 76.430 250.200 76.580 258.400 ;
        RECT 77.030 250.200 77.180 258.400 ;
        RECT 77.630 250.200 77.780 258.400 ;
        RECT 78.230 250.200 78.380 258.400 ;
        RECT 78.830 250.200 78.980 258.400 ;
        RECT 83.530 257.850 85.940 258.800 ;
        RECT 79.580 257.700 89.880 257.850 ;
        RECT 83.130 257.250 86.330 257.700 ;
        RECT 79.580 257.100 89.880 257.250 ;
        RECT 83.130 256.650 86.330 257.100 ;
        RECT 79.580 256.500 89.880 256.650 ;
        RECT 83.130 256.050 86.330 256.500 ;
        RECT 79.580 255.900 89.880 256.050 ;
        RECT 83.130 255.600 86.330 255.900 ;
        RECT 83.130 255.450 83.530 255.600 ;
        RECT 79.580 255.300 83.530 255.450 ;
        RECT 83.130 254.850 83.530 255.300 ;
        RECT 79.580 254.700 83.530 254.850 ;
        RECT 83.130 254.250 83.530 254.700 ;
        RECT 79.580 254.100 83.530 254.250 ;
        RECT 83.130 253.650 83.530 254.100 ;
        RECT 79.580 253.500 83.530 253.650 ;
        RECT 83.130 253.050 83.530 253.500 ;
        RECT 79.580 252.900 83.530 253.050 ;
        RECT 83.130 252.450 83.530 252.900 ;
        RECT 79.580 252.300 83.530 252.450 ;
        RECT 83.130 251.850 83.530 252.300 ;
        RECT 79.580 251.700 83.530 251.850 ;
        RECT 83.130 251.250 83.530 251.700 ;
        RECT 79.580 251.100 83.530 251.250 ;
        RECT 83.130 250.650 83.530 251.100 ;
        RECT 79.580 250.500 83.530 250.650 ;
        RECT 83.130 250.200 83.530 250.500 ;
        RECT 75.230 249.800 83.530 250.200 ;
        RECT 75.230 241.600 75.380 249.800 ;
        RECT 75.830 241.600 75.980 249.800 ;
        RECT 76.430 241.600 76.580 249.800 ;
        RECT 77.030 241.600 77.180 249.800 ;
        RECT 77.630 241.600 77.780 249.800 ;
        RECT 78.230 241.600 78.380 249.800 ;
        RECT 78.830 241.600 78.980 249.800 ;
        RECT 83.130 249.500 83.530 249.800 ;
        RECT 79.580 249.350 83.530 249.500 ;
        RECT 83.130 248.900 83.530 249.350 ;
        RECT 79.580 248.750 83.530 248.900 ;
        RECT 83.130 248.300 83.530 248.750 ;
        RECT 79.580 248.150 83.530 248.300 ;
        RECT 83.130 247.700 83.530 248.150 ;
        RECT 79.580 247.550 83.530 247.700 ;
        RECT 83.130 247.100 83.530 247.550 ;
        RECT 79.580 246.950 83.530 247.100 ;
        RECT 83.130 246.500 83.530 246.950 ;
        RECT 79.580 246.350 83.530 246.500 ;
        RECT 83.130 245.900 83.530 246.350 ;
        RECT 79.580 245.750 83.530 245.900 ;
        RECT 83.130 245.300 83.530 245.750 ;
        RECT 79.580 245.150 83.530 245.300 ;
        RECT 83.130 244.700 83.530 245.150 ;
        RECT 79.580 244.550 83.530 244.700 ;
        RECT 83.130 244.400 83.530 244.550 ;
        RECT 85.930 255.450 86.330 255.600 ;
        RECT 85.930 255.300 89.880 255.450 ;
        RECT 85.930 254.850 86.330 255.300 ;
        RECT 85.930 254.700 89.880 254.850 ;
        RECT 85.930 254.250 86.330 254.700 ;
        RECT 85.930 254.100 89.880 254.250 ;
        RECT 85.930 253.650 86.330 254.100 ;
        RECT 85.930 253.500 89.880 253.650 ;
        RECT 85.930 253.050 86.330 253.500 ;
        RECT 85.930 252.900 89.880 253.050 ;
        RECT 85.930 252.450 86.330 252.900 ;
        RECT 85.930 252.300 89.880 252.450 ;
        RECT 85.930 251.850 86.330 252.300 ;
        RECT 85.930 251.700 89.880 251.850 ;
        RECT 85.930 251.250 86.330 251.700 ;
        RECT 85.930 251.100 89.880 251.250 ;
        RECT 85.930 250.650 86.330 251.100 ;
        RECT 85.930 250.500 89.880 250.650 ;
        RECT 85.930 250.200 86.330 250.500 ;
        RECT 90.480 250.200 90.630 258.400 ;
        RECT 91.080 250.200 91.230 258.400 ;
        RECT 91.680 250.200 91.830 258.400 ;
        RECT 92.280 250.200 92.430 258.400 ;
        RECT 92.880 250.200 93.030 258.400 ;
        RECT 93.480 250.200 93.630 258.400 ;
        RECT 94.080 250.200 94.230 258.400 ;
        RECT 85.930 249.800 94.230 250.200 ;
        RECT 85.930 249.500 86.330 249.800 ;
        RECT 85.930 249.350 89.880 249.500 ;
        RECT 85.930 248.900 86.330 249.350 ;
        RECT 85.930 248.750 89.880 248.900 ;
        RECT 85.930 248.300 86.330 248.750 ;
        RECT 85.930 248.150 89.880 248.300 ;
        RECT 85.930 247.700 86.330 248.150 ;
        RECT 85.930 247.550 89.880 247.700 ;
        RECT 85.930 247.100 86.330 247.550 ;
        RECT 85.930 246.950 89.880 247.100 ;
        RECT 85.930 246.500 86.330 246.950 ;
        RECT 85.930 246.350 89.880 246.500 ;
        RECT 85.930 245.900 86.330 246.350 ;
        RECT 85.930 245.750 89.880 245.900 ;
        RECT 85.930 245.300 86.330 245.750 ;
        RECT 85.930 245.150 89.880 245.300 ;
        RECT 85.930 244.700 86.330 245.150 ;
        RECT 85.930 244.550 89.880 244.700 ;
        RECT 85.930 244.400 86.330 244.550 ;
        RECT 83.130 244.100 86.330 244.400 ;
        RECT 79.580 243.950 89.880 244.100 ;
        RECT 83.130 243.500 86.330 243.950 ;
        RECT 79.580 243.350 89.880 243.500 ;
        RECT 83.130 242.900 86.330 243.350 ;
        RECT 79.580 242.750 89.880 242.900 ;
        RECT 83.130 242.300 86.330 242.750 ;
        RECT 79.580 242.150 89.880 242.300 ;
        RECT 83.530 241.200 85.930 242.150 ;
        RECT 90.480 241.600 90.630 249.800 ;
        RECT 91.080 241.600 91.230 249.800 ;
        RECT 91.680 241.600 91.830 249.800 ;
        RECT 92.280 241.600 92.430 249.800 ;
        RECT 92.880 241.600 93.030 249.800 ;
        RECT 93.480 241.600 93.630 249.800 ;
        RECT 94.080 241.600 94.230 249.800 ;
        RECT 95.230 250.200 95.380 258.400 ;
        RECT 95.830 250.200 95.980 258.400 ;
        RECT 96.430 250.200 96.580 258.400 ;
        RECT 97.030 250.200 97.180 258.400 ;
        RECT 97.630 250.200 97.780 258.400 ;
        RECT 98.230 250.200 98.380 258.400 ;
        RECT 98.830 250.200 98.980 258.400 ;
        RECT 103.530 257.850 104.730 258.800 ;
        RECT 99.580 257.700 104.730 257.850 ;
        RECT 103.130 257.250 104.730 257.700 ;
        RECT 99.580 257.100 104.730 257.250 ;
        RECT 103.130 256.650 104.730 257.100 ;
        RECT 99.580 256.500 104.730 256.650 ;
        RECT 103.130 256.050 104.730 256.500 ;
        RECT 105.140 256.050 107.140 257.325 ;
        RECT 99.580 255.900 104.730 256.050 ;
        RECT 103.130 255.600 104.730 255.900 ;
        RECT 103.130 255.450 103.530 255.600 ;
        RECT 99.580 255.300 103.530 255.450 ;
        RECT 103.130 254.850 103.530 255.300 ;
        RECT 99.580 254.700 103.530 254.850 ;
        RECT 103.130 254.250 103.530 254.700 ;
        RECT 99.580 254.100 103.530 254.250 ;
        RECT 103.130 253.650 103.530 254.100 ;
        RECT 99.580 253.500 103.530 253.650 ;
        RECT 103.130 253.050 103.530 253.500 ;
        RECT 99.580 252.900 103.530 253.050 ;
        RECT 103.130 252.450 103.530 252.900 ;
        RECT 99.580 252.300 103.530 252.450 ;
        RECT 103.130 251.850 103.530 252.300 ;
        RECT 99.580 251.700 103.530 251.850 ;
        RECT 103.130 251.250 103.530 251.700 ;
        RECT 99.580 251.100 103.530 251.250 ;
        RECT 103.130 250.650 103.530 251.100 ;
        RECT 99.580 250.500 103.530 250.650 ;
        RECT 103.130 250.200 103.530 250.500 ;
        RECT 95.230 249.800 103.530 250.200 ;
        RECT 95.230 241.600 95.380 249.800 ;
        RECT 95.830 241.600 95.980 249.800 ;
        RECT 96.430 241.600 96.580 249.800 ;
        RECT 97.030 241.600 97.180 249.800 ;
        RECT 97.630 241.600 97.780 249.800 ;
        RECT 98.230 241.600 98.380 249.800 ;
        RECT 98.830 241.600 98.980 249.800 ;
        RECT 103.130 249.500 103.530 249.800 ;
        RECT 99.580 249.350 103.530 249.500 ;
        RECT 103.130 248.900 103.530 249.350 ;
        RECT 99.580 248.750 103.530 248.900 ;
        RECT 103.130 248.300 103.530 248.750 ;
        RECT 99.580 248.150 103.530 248.300 ;
        RECT 103.130 247.700 103.530 248.150 ;
        RECT 99.580 247.550 103.530 247.700 ;
        RECT 103.130 247.100 103.530 247.550 ;
        RECT 99.580 246.950 103.530 247.100 ;
        RECT 103.130 246.500 103.530 246.950 ;
        RECT 99.580 246.350 103.530 246.500 ;
        RECT 103.130 245.900 103.530 246.350 ;
        RECT 99.580 245.750 103.530 245.900 ;
        RECT 103.130 245.300 103.530 245.750 ;
        RECT 99.580 245.150 103.530 245.300 ;
        RECT 103.130 244.700 103.530 245.150 ;
        RECT 99.580 244.550 103.530 244.700 ;
        RECT 103.130 244.400 103.530 244.550 ;
        RECT 103.130 244.100 104.730 244.400 ;
        RECT 99.580 243.950 104.730 244.100 ;
        RECT 103.130 243.500 104.730 243.950 ;
        RECT 99.580 243.350 104.730 243.500 ;
        RECT 103.130 242.900 104.730 243.350 ;
        RECT 99.580 242.750 104.730 242.900 ;
        RECT 103.130 242.300 104.730 242.750 ;
        RECT 99.580 242.150 104.730 242.300 ;
        RECT 105.140 242.255 107.140 243.530 ;
        RECT 103.530 241.200 104.730 242.150 ;
        RECT 4.730 238.800 9.130 241.200 ;
        RECT 20.330 238.800 29.130 241.200 ;
        RECT 40.330 238.800 49.130 241.200 ;
        RECT 60.330 238.800 69.130 241.200 ;
        RECT 80.330 238.800 89.130 241.200 ;
        RECT 100.330 238.800 104.730 241.200 ;
        RECT 2.315 236.695 4.320 237.970 ;
        RECT 4.730 237.850 5.940 238.800 ;
        RECT 4.730 237.700 9.880 237.850 ;
        RECT 4.730 237.250 6.330 237.700 ;
        RECT 4.730 237.100 9.880 237.250 ;
        RECT 4.730 236.650 6.330 237.100 ;
        RECT 4.730 236.500 9.880 236.650 ;
        RECT 4.730 236.050 6.330 236.500 ;
        RECT 4.730 235.900 9.880 236.050 ;
        RECT 4.730 235.600 6.330 235.900 ;
        RECT 2.315 233.250 4.315 235.545 ;
        RECT 5.930 235.450 6.330 235.600 ;
        RECT 5.930 235.300 9.880 235.450 ;
        RECT 5.930 234.850 6.330 235.300 ;
        RECT 5.930 234.700 9.880 234.850 ;
        RECT 5.930 234.250 6.330 234.700 ;
        RECT 5.930 234.100 9.880 234.250 ;
        RECT 5.930 233.650 6.330 234.100 ;
        RECT 5.930 233.500 9.880 233.650 ;
        RECT 5.930 233.050 6.330 233.500 ;
        RECT 5.930 232.900 9.880 233.050 ;
        RECT 5.930 232.450 6.330 232.900 ;
        RECT 5.930 232.300 9.880 232.450 ;
        RECT 5.930 231.850 6.330 232.300 ;
        RECT 5.930 231.700 9.880 231.850 ;
        RECT 5.930 231.250 6.330 231.700 ;
        RECT 5.930 231.100 9.880 231.250 ;
        RECT 5.930 230.650 6.330 231.100 ;
        RECT 5.930 230.500 9.880 230.650 ;
        RECT 5.930 230.200 6.330 230.500 ;
        RECT 10.480 230.200 10.630 238.400 ;
        RECT 11.080 230.200 11.230 238.400 ;
        RECT 11.680 230.200 11.830 238.400 ;
        RECT 12.280 230.200 12.430 238.400 ;
        RECT 12.880 230.200 13.030 238.400 ;
        RECT 13.480 230.200 13.630 238.400 ;
        RECT 14.080 230.200 14.230 238.400 ;
        RECT 5.930 229.800 14.230 230.200 ;
        RECT 5.930 229.500 6.330 229.800 ;
        RECT 5.930 229.350 9.880 229.500 ;
        RECT 5.930 228.900 6.330 229.350 ;
        RECT 5.930 228.750 9.880 228.900 ;
        RECT 5.930 228.300 6.330 228.750 ;
        RECT 5.930 228.150 9.880 228.300 ;
        RECT 5.930 227.700 6.330 228.150 ;
        RECT 5.930 227.550 9.880 227.700 ;
        RECT 5.930 227.100 6.330 227.550 ;
        RECT 5.930 226.950 9.880 227.100 ;
        RECT 2.315 224.455 4.315 226.750 ;
        RECT 5.930 226.500 6.330 226.950 ;
        RECT 5.930 226.350 9.880 226.500 ;
        RECT 5.930 225.900 6.330 226.350 ;
        RECT 5.930 225.750 9.880 225.900 ;
        RECT 5.930 225.300 6.330 225.750 ;
        RECT 5.930 225.150 9.880 225.300 ;
        RECT 5.930 224.700 6.330 225.150 ;
        RECT 5.930 224.550 9.880 224.700 ;
        RECT 2.315 224.450 4.180 224.455 ;
        RECT 5.930 224.400 6.330 224.550 ;
        RECT 4.730 224.100 6.330 224.400 ;
        RECT 4.730 223.950 9.880 224.100 ;
        RECT 4.730 223.500 6.330 223.950 ;
        RECT 4.730 223.350 9.880 223.500 ;
        RECT 4.730 222.900 6.330 223.350 ;
        RECT 4.730 222.750 9.880 222.900 ;
        RECT 2.315 221.395 4.315 222.670 ;
        RECT 4.730 222.300 6.330 222.750 ;
        RECT 4.730 222.150 9.880 222.300 ;
        RECT 4.730 221.200 5.930 222.150 ;
        RECT 10.480 221.600 10.630 229.800 ;
        RECT 11.080 221.600 11.230 229.800 ;
        RECT 11.680 221.600 11.830 229.800 ;
        RECT 12.280 221.600 12.430 229.800 ;
        RECT 12.880 221.600 13.030 229.800 ;
        RECT 13.480 221.600 13.630 229.800 ;
        RECT 14.080 221.600 14.230 229.800 ;
        RECT 15.230 230.200 15.380 238.400 ;
        RECT 15.830 230.200 15.980 238.400 ;
        RECT 16.430 230.200 16.580 238.400 ;
        RECT 17.030 230.200 17.180 238.400 ;
        RECT 17.630 230.200 17.780 238.400 ;
        RECT 18.230 230.200 18.380 238.400 ;
        RECT 18.830 230.200 18.980 238.400 ;
        RECT 23.530 237.850 25.940 238.800 ;
        RECT 19.580 237.700 29.880 237.850 ;
        RECT 23.130 237.250 26.330 237.700 ;
        RECT 19.580 237.100 29.880 237.250 ;
        RECT 23.130 236.650 26.330 237.100 ;
        RECT 19.580 236.500 29.880 236.650 ;
        RECT 23.130 236.050 26.330 236.500 ;
        RECT 19.580 235.900 29.880 236.050 ;
        RECT 23.130 235.600 26.330 235.900 ;
        RECT 23.130 235.450 23.530 235.600 ;
        RECT 19.580 235.300 23.530 235.450 ;
        RECT 23.130 234.850 23.530 235.300 ;
        RECT 19.580 234.700 23.530 234.850 ;
        RECT 23.130 234.250 23.530 234.700 ;
        RECT 19.580 234.100 23.530 234.250 ;
        RECT 23.130 233.650 23.530 234.100 ;
        RECT 19.580 233.500 23.530 233.650 ;
        RECT 23.130 233.050 23.530 233.500 ;
        RECT 19.580 232.900 23.530 233.050 ;
        RECT 23.130 232.450 23.530 232.900 ;
        RECT 19.580 232.300 23.530 232.450 ;
        RECT 23.130 231.850 23.530 232.300 ;
        RECT 19.580 231.700 23.530 231.850 ;
        RECT 23.130 231.250 23.530 231.700 ;
        RECT 19.580 231.100 23.530 231.250 ;
        RECT 23.130 230.650 23.530 231.100 ;
        RECT 19.580 230.500 23.530 230.650 ;
        RECT 23.130 230.200 23.530 230.500 ;
        RECT 15.230 229.800 23.530 230.200 ;
        RECT 15.230 221.600 15.380 229.800 ;
        RECT 15.830 221.600 15.980 229.800 ;
        RECT 16.430 221.600 16.580 229.800 ;
        RECT 17.030 221.600 17.180 229.800 ;
        RECT 17.630 221.600 17.780 229.800 ;
        RECT 18.230 221.600 18.380 229.800 ;
        RECT 18.830 221.600 18.980 229.800 ;
        RECT 23.130 229.500 23.530 229.800 ;
        RECT 19.580 229.350 23.530 229.500 ;
        RECT 23.130 228.900 23.530 229.350 ;
        RECT 19.580 228.750 23.530 228.900 ;
        RECT 23.130 228.300 23.530 228.750 ;
        RECT 19.580 228.150 23.530 228.300 ;
        RECT 23.130 227.700 23.530 228.150 ;
        RECT 19.580 227.550 23.530 227.700 ;
        RECT 23.130 227.100 23.530 227.550 ;
        RECT 19.580 226.950 23.530 227.100 ;
        RECT 23.130 226.500 23.530 226.950 ;
        RECT 19.580 226.350 23.530 226.500 ;
        RECT 23.130 225.900 23.530 226.350 ;
        RECT 19.580 225.750 23.530 225.900 ;
        RECT 23.130 225.300 23.530 225.750 ;
        RECT 19.580 225.150 23.530 225.300 ;
        RECT 23.130 224.700 23.530 225.150 ;
        RECT 19.580 224.550 23.530 224.700 ;
        RECT 23.130 224.400 23.530 224.550 ;
        RECT 25.930 235.450 26.330 235.600 ;
        RECT 25.930 235.300 29.880 235.450 ;
        RECT 25.930 234.850 26.330 235.300 ;
        RECT 25.930 234.700 29.880 234.850 ;
        RECT 25.930 234.250 26.330 234.700 ;
        RECT 25.930 234.100 29.880 234.250 ;
        RECT 25.930 233.650 26.330 234.100 ;
        RECT 25.930 233.500 29.880 233.650 ;
        RECT 25.930 233.050 26.330 233.500 ;
        RECT 25.930 232.900 29.880 233.050 ;
        RECT 25.930 232.450 26.330 232.900 ;
        RECT 25.930 232.300 29.880 232.450 ;
        RECT 25.930 231.850 26.330 232.300 ;
        RECT 25.930 231.700 29.880 231.850 ;
        RECT 25.930 231.250 26.330 231.700 ;
        RECT 25.930 231.100 29.880 231.250 ;
        RECT 25.930 230.650 26.330 231.100 ;
        RECT 25.930 230.500 29.880 230.650 ;
        RECT 25.930 230.200 26.330 230.500 ;
        RECT 30.480 230.200 30.630 238.400 ;
        RECT 31.080 230.200 31.230 238.400 ;
        RECT 31.680 230.200 31.830 238.400 ;
        RECT 32.280 230.200 32.430 238.400 ;
        RECT 32.880 230.200 33.030 238.400 ;
        RECT 33.480 230.200 33.630 238.400 ;
        RECT 34.080 230.200 34.230 238.400 ;
        RECT 25.930 229.800 34.230 230.200 ;
        RECT 25.930 229.500 26.330 229.800 ;
        RECT 25.930 229.350 29.880 229.500 ;
        RECT 25.930 228.900 26.330 229.350 ;
        RECT 25.930 228.750 29.880 228.900 ;
        RECT 25.930 228.300 26.330 228.750 ;
        RECT 25.930 228.150 29.880 228.300 ;
        RECT 25.930 227.700 26.330 228.150 ;
        RECT 25.930 227.550 29.880 227.700 ;
        RECT 25.930 227.100 26.330 227.550 ;
        RECT 25.930 226.950 29.880 227.100 ;
        RECT 25.930 226.500 26.330 226.950 ;
        RECT 25.930 226.350 29.880 226.500 ;
        RECT 25.930 225.900 26.330 226.350 ;
        RECT 25.930 225.750 29.880 225.900 ;
        RECT 25.930 225.300 26.330 225.750 ;
        RECT 25.930 225.150 29.880 225.300 ;
        RECT 25.930 224.700 26.330 225.150 ;
        RECT 25.930 224.550 29.880 224.700 ;
        RECT 25.930 224.400 26.330 224.550 ;
        RECT 23.130 224.100 26.330 224.400 ;
        RECT 19.580 223.950 29.880 224.100 ;
        RECT 23.130 223.500 26.330 223.950 ;
        RECT 19.580 223.350 29.880 223.500 ;
        RECT 23.130 222.900 26.330 223.350 ;
        RECT 19.580 222.750 29.880 222.900 ;
        RECT 23.130 222.300 26.330 222.750 ;
        RECT 19.580 222.150 29.880 222.300 ;
        RECT 23.530 221.200 25.930 222.150 ;
        RECT 30.480 221.600 30.630 229.800 ;
        RECT 31.080 221.600 31.230 229.800 ;
        RECT 31.680 221.600 31.830 229.800 ;
        RECT 32.280 221.600 32.430 229.800 ;
        RECT 32.880 221.600 33.030 229.800 ;
        RECT 33.480 221.600 33.630 229.800 ;
        RECT 34.080 221.600 34.230 229.800 ;
        RECT 35.230 230.200 35.380 238.400 ;
        RECT 35.830 230.200 35.980 238.400 ;
        RECT 36.430 230.200 36.580 238.400 ;
        RECT 37.030 230.200 37.180 238.400 ;
        RECT 37.630 230.200 37.780 238.400 ;
        RECT 38.230 230.200 38.380 238.400 ;
        RECT 38.830 230.200 38.980 238.400 ;
        RECT 43.530 237.850 45.940 238.800 ;
        RECT 39.580 237.700 49.880 237.850 ;
        RECT 43.130 237.250 46.330 237.700 ;
        RECT 39.580 237.100 49.880 237.250 ;
        RECT 43.130 236.650 46.330 237.100 ;
        RECT 39.580 236.500 49.880 236.650 ;
        RECT 43.130 236.050 46.330 236.500 ;
        RECT 39.580 235.900 49.880 236.050 ;
        RECT 43.130 235.600 46.330 235.900 ;
        RECT 43.130 235.450 43.530 235.600 ;
        RECT 39.580 235.300 43.530 235.450 ;
        RECT 43.130 234.850 43.530 235.300 ;
        RECT 39.580 234.700 43.530 234.850 ;
        RECT 43.130 234.250 43.530 234.700 ;
        RECT 39.580 234.100 43.530 234.250 ;
        RECT 43.130 233.650 43.530 234.100 ;
        RECT 39.580 233.500 43.530 233.650 ;
        RECT 43.130 233.050 43.530 233.500 ;
        RECT 39.580 232.900 43.530 233.050 ;
        RECT 43.130 232.450 43.530 232.900 ;
        RECT 39.580 232.300 43.530 232.450 ;
        RECT 43.130 231.850 43.530 232.300 ;
        RECT 39.580 231.700 43.530 231.850 ;
        RECT 43.130 231.250 43.530 231.700 ;
        RECT 39.580 231.100 43.530 231.250 ;
        RECT 43.130 230.650 43.530 231.100 ;
        RECT 39.580 230.500 43.530 230.650 ;
        RECT 43.130 230.200 43.530 230.500 ;
        RECT 35.230 229.800 43.530 230.200 ;
        RECT 35.230 221.600 35.380 229.800 ;
        RECT 35.830 221.600 35.980 229.800 ;
        RECT 36.430 221.600 36.580 229.800 ;
        RECT 37.030 221.600 37.180 229.800 ;
        RECT 37.630 221.600 37.780 229.800 ;
        RECT 38.230 221.600 38.380 229.800 ;
        RECT 38.830 221.600 38.980 229.800 ;
        RECT 43.130 229.500 43.530 229.800 ;
        RECT 39.580 229.350 43.530 229.500 ;
        RECT 43.130 228.900 43.530 229.350 ;
        RECT 39.580 228.750 43.530 228.900 ;
        RECT 43.130 228.300 43.530 228.750 ;
        RECT 39.580 228.150 43.530 228.300 ;
        RECT 43.130 227.700 43.530 228.150 ;
        RECT 39.580 227.550 43.530 227.700 ;
        RECT 43.130 227.100 43.530 227.550 ;
        RECT 39.580 226.950 43.530 227.100 ;
        RECT 43.130 226.500 43.530 226.950 ;
        RECT 39.580 226.350 43.530 226.500 ;
        RECT 43.130 225.900 43.530 226.350 ;
        RECT 39.580 225.750 43.530 225.900 ;
        RECT 43.130 225.300 43.530 225.750 ;
        RECT 39.580 225.150 43.530 225.300 ;
        RECT 43.130 224.700 43.530 225.150 ;
        RECT 39.580 224.550 43.530 224.700 ;
        RECT 43.130 224.400 43.530 224.550 ;
        RECT 45.930 235.450 46.330 235.600 ;
        RECT 45.930 235.300 49.880 235.450 ;
        RECT 45.930 234.850 46.330 235.300 ;
        RECT 45.930 234.700 49.880 234.850 ;
        RECT 45.930 234.250 46.330 234.700 ;
        RECT 45.930 234.100 49.880 234.250 ;
        RECT 45.930 233.650 46.330 234.100 ;
        RECT 45.930 233.500 49.880 233.650 ;
        RECT 45.930 233.050 46.330 233.500 ;
        RECT 45.930 232.900 49.880 233.050 ;
        RECT 45.930 232.450 46.330 232.900 ;
        RECT 45.930 232.300 49.880 232.450 ;
        RECT 45.930 231.850 46.330 232.300 ;
        RECT 45.930 231.700 49.880 231.850 ;
        RECT 45.930 231.250 46.330 231.700 ;
        RECT 45.930 231.100 49.880 231.250 ;
        RECT 45.930 230.650 46.330 231.100 ;
        RECT 45.930 230.500 49.880 230.650 ;
        RECT 45.930 230.200 46.330 230.500 ;
        RECT 50.480 230.200 50.630 238.400 ;
        RECT 51.080 230.200 51.230 238.400 ;
        RECT 51.680 230.200 51.830 238.400 ;
        RECT 52.280 230.200 52.430 238.400 ;
        RECT 52.880 230.200 53.030 238.400 ;
        RECT 53.480 230.200 53.630 238.400 ;
        RECT 54.080 230.200 54.230 238.400 ;
        RECT 45.930 229.800 54.230 230.200 ;
        RECT 45.930 229.500 46.330 229.800 ;
        RECT 45.930 229.350 49.880 229.500 ;
        RECT 45.930 228.900 46.330 229.350 ;
        RECT 45.930 228.750 49.880 228.900 ;
        RECT 45.930 228.300 46.330 228.750 ;
        RECT 45.930 228.150 49.880 228.300 ;
        RECT 45.930 227.700 46.330 228.150 ;
        RECT 45.930 227.550 49.880 227.700 ;
        RECT 45.930 227.100 46.330 227.550 ;
        RECT 45.930 226.950 49.880 227.100 ;
        RECT 45.930 226.500 46.330 226.950 ;
        RECT 45.930 226.350 49.880 226.500 ;
        RECT 45.930 225.900 46.330 226.350 ;
        RECT 45.930 225.750 49.880 225.900 ;
        RECT 45.930 225.300 46.330 225.750 ;
        RECT 45.930 225.150 49.880 225.300 ;
        RECT 45.930 224.700 46.330 225.150 ;
        RECT 45.930 224.550 49.880 224.700 ;
        RECT 45.930 224.400 46.330 224.550 ;
        RECT 43.130 224.100 46.330 224.400 ;
        RECT 39.580 223.950 49.880 224.100 ;
        RECT 43.130 223.500 46.330 223.950 ;
        RECT 39.580 223.350 49.880 223.500 ;
        RECT 43.130 222.900 46.330 223.350 ;
        RECT 39.580 222.750 49.880 222.900 ;
        RECT 43.130 222.300 46.330 222.750 ;
        RECT 39.580 222.150 49.880 222.300 ;
        RECT 43.530 221.200 45.930 222.150 ;
        RECT 50.480 221.600 50.630 229.800 ;
        RECT 51.080 221.600 51.230 229.800 ;
        RECT 51.680 221.600 51.830 229.800 ;
        RECT 52.280 221.600 52.430 229.800 ;
        RECT 52.880 221.600 53.030 229.800 ;
        RECT 53.480 221.600 53.630 229.800 ;
        RECT 54.080 221.600 54.230 229.800 ;
        RECT 55.230 230.200 55.380 238.400 ;
        RECT 55.830 230.200 55.980 238.400 ;
        RECT 56.430 230.200 56.580 238.400 ;
        RECT 57.030 230.200 57.180 238.400 ;
        RECT 57.630 230.200 57.780 238.400 ;
        RECT 58.230 230.200 58.380 238.400 ;
        RECT 58.830 230.200 58.980 238.400 ;
        RECT 63.530 237.850 65.940 238.800 ;
        RECT 59.580 237.700 69.880 237.850 ;
        RECT 63.130 237.250 66.330 237.700 ;
        RECT 59.580 237.100 69.880 237.250 ;
        RECT 63.130 236.650 66.330 237.100 ;
        RECT 59.580 236.500 69.880 236.650 ;
        RECT 63.130 236.050 66.330 236.500 ;
        RECT 59.580 235.900 69.880 236.050 ;
        RECT 63.130 235.600 66.330 235.900 ;
        RECT 63.130 235.450 63.530 235.600 ;
        RECT 59.580 235.300 63.530 235.450 ;
        RECT 63.130 234.850 63.530 235.300 ;
        RECT 59.580 234.700 63.530 234.850 ;
        RECT 63.130 234.250 63.530 234.700 ;
        RECT 59.580 234.100 63.530 234.250 ;
        RECT 63.130 233.650 63.530 234.100 ;
        RECT 59.580 233.500 63.530 233.650 ;
        RECT 63.130 233.050 63.530 233.500 ;
        RECT 59.580 232.900 63.530 233.050 ;
        RECT 63.130 232.450 63.530 232.900 ;
        RECT 59.580 232.300 63.530 232.450 ;
        RECT 63.130 231.850 63.530 232.300 ;
        RECT 59.580 231.700 63.530 231.850 ;
        RECT 63.130 231.250 63.530 231.700 ;
        RECT 59.580 231.100 63.530 231.250 ;
        RECT 63.130 230.650 63.530 231.100 ;
        RECT 59.580 230.500 63.530 230.650 ;
        RECT 63.130 230.200 63.530 230.500 ;
        RECT 55.230 229.800 63.530 230.200 ;
        RECT 55.230 221.600 55.380 229.800 ;
        RECT 55.830 221.600 55.980 229.800 ;
        RECT 56.430 221.600 56.580 229.800 ;
        RECT 57.030 221.600 57.180 229.800 ;
        RECT 57.630 221.600 57.780 229.800 ;
        RECT 58.230 221.600 58.380 229.800 ;
        RECT 58.830 221.600 58.980 229.800 ;
        RECT 63.130 229.500 63.530 229.800 ;
        RECT 59.580 229.350 63.530 229.500 ;
        RECT 63.130 228.900 63.530 229.350 ;
        RECT 59.580 228.750 63.530 228.900 ;
        RECT 63.130 228.300 63.530 228.750 ;
        RECT 59.580 228.150 63.530 228.300 ;
        RECT 63.130 227.700 63.530 228.150 ;
        RECT 59.580 227.550 63.530 227.700 ;
        RECT 63.130 227.100 63.530 227.550 ;
        RECT 59.580 226.950 63.530 227.100 ;
        RECT 63.130 226.500 63.530 226.950 ;
        RECT 59.580 226.350 63.530 226.500 ;
        RECT 63.130 225.900 63.530 226.350 ;
        RECT 59.580 225.750 63.530 225.900 ;
        RECT 63.130 225.300 63.530 225.750 ;
        RECT 59.580 225.150 63.530 225.300 ;
        RECT 63.130 224.700 63.530 225.150 ;
        RECT 59.580 224.550 63.530 224.700 ;
        RECT 63.130 224.400 63.530 224.550 ;
        RECT 65.930 235.450 66.330 235.600 ;
        RECT 65.930 235.300 69.880 235.450 ;
        RECT 65.930 234.850 66.330 235.300 ;
        RECT 65.930 234.700 69.880 234.850 ;
        RECT 65.930 234.250 66.330 234.700 ;
        RECT 65.930 234.100 69.880 234.250 ;
        RECT 65.930 233.650 66.330 234.100 ;
        RECT 65.930 233.500 69.880 233.650 ;
        RECT 65.930 233.050 66.330 233.500 ;
        RECT 65.930 232.900 69.880 233.050 ;
        RECT 65.930 232.450 66.330 232.900 ;
        RECT 65.930 232.300 69.880 232.450 ;
        RECT 65.930 231.850 66.330 232.300 ;
        RECT 65.930 231.700 69.880 231.850 ;
        RECT 65.930 231.250 66.330 231.700 ;
        RECT 65.930 231.100 69.880 231.250 ;
        RECT 65.930 230.650 66.330 231.100 ;
        RECT 65.930 230.500 69.880 230.650 ;
        RECT 65.930 230.200 66.330 230.500 ;
        RECT 70.480 230.200 70.630 238.400 ;
        RECT 71.080 230.200 71.230 238.400 ;
        RECT 71.680 230.200 71.830 238.400 ;
        RECT 72.280 230.200 72.430 238.400 ;
        RECT 72.880 230.200 73.030 238.400 ;
        RECT 73.480 230.200 73.630 238.400 ;
        RECT 74.080 230.200 74.230 238.400 ;
        RECT 65.930 229.800 74.230 230.200 ;
        RECT 65.930 229.500 66.330 229.800 ;
        RECT 65.930 229.350 69.880 229.500 ;
        RECT 65.930 228.900 66.330 229.350 ;
        RECT 65.930 228.750 69.880 228.900 ;
        RECT 65.930 228.300 66.330 228.750 ;
        RECT 65.930 228.150 69.880 228.300 ;
        RECT 65.930 227.700 66.330 228.150 ;
        RECT 65.930 227.550 69.880 227.700 ;
        RECT 65.930 227.100 66.330 227.550 ;
        RECT 65.930 226.950 69.880 227.100 ;
        RECT 65.930 226.500 66.330 226.950 ;
        RECT 65.930 226.350 69.880 226.500 ;
        RECT 65.930 225.900 66.330 226.350 ;
        RECT 65.930 225.750 69.880 225.900 ;
        RECT 65.930 225.300 66.330 225.750 ;
        RECT 65.930 225.150 69.880 225.300 ;
        RECT 65.930 224.700 66.330 225.150 ;
        RECT 65.930 224.550 69.880 224.700 ;
        RECT 65.930 224.400 66.330 224.550 ;
        RECT 63.130 224.100 66.330 224.400 ;
        RECT 59.580 223.950 69.880 224.100 ;
        RECT 63.130 223.500 66.330 223.950 ;
        RECT 59.580 223.350 69.880 223.500 ;
        RECT 63.130 222.900 66.330 223.350 ;
        RECT 59.580 222.750 69.880 222.900 ;
        RECT 63.130 222.300 66.330 222.750 ;
        RECT 59.580 222.150 69.880 222.300 ;
        RECT 63.530 221.200 65.930 222.150 ;
        RECT 70.480 221.600 70.630 229.800 ;
        RECT 71.080 221.600 71.230 229.800 ;
        RECT 71.680 221.600 71.830 229.800 ;
        RECT 72.280 221.600 72.430 229.800 ;
        RECT 72.880 221.600 73.030 229.800 ;
        RECT 73.480 221.600 73.630 229.800 ;
        RECT 74.080 221.600 74.230 229.800 ;
        RECT 75.230 230.200 75.380 238.400 ;
        RECT 75.830 230.200 75.980 238.400 ;
        RECT 76.430 230.200 76.580 238.400 ;
        RECT 77.030 230.200 77.180 238.400 ;
        RECT 77.630 230.200 77.780 238.400 ;
        RECT 78.230 230.200 78.380 238.400 ;
        RECT 78.830 230.200 78.980 238.400 ;
        RECT 83.530 237.850 85.940 238.800 ;
        RECT 79.580 237.700 89.880 237.850 ;
        RECT 83.130 237.250 86.330 237.700 ;
        RECT 79.580 237.100 89.880 237.250 ;
        RECT 83.130 236.650 86.330 237.100 ;
        RECT 79.580 236.500 89.880 236.650 ;
        RECT 83.130 236.050 86.330 236.500 ;
        RECT 79.580 235.900 89.880 236.050 ;
        RECT 83.130 235.600 86.330 235.900 ;
        RECT 83.130 235.450 83.530 235.600 ;
        RECT 79.580 235.300 83.530 235.450 ;
        RECT 83.130 234.850 83.530 235.300 ;
        RECT 79.580 234.700 83.530 234.850 ;
        RECT 83.130 234.250 83.530 234.700 ;
        RECT 79.580 234.100 83.530 234.250 ;
        RECT 83.130 233.650 83.530 234.100 ;
        RECT 79.580 233.500 83.530 233.650 ;
        RECT 83.130 233.050 83.530 233.500 ;
        RECT 79.580 232.900 83.530 233.050 ;
        RECT 83.130 232.450 83.530 232.900 ;
        RECT 79.580 232.300 83.530 232.450 ;
        RECT 83.130 231.850 83.530 232.300 ;
        RECT 79.580 231.700 83.530 231.850 ;
        RECT 83.130 231.250 83.530 231.700 ;
        RECT 79.580 231.100 83.530 231.250 ;
        RECT 83.130 230.650 83.530 231.100 ;
        RECT 79.580 230.500 83.530 230.650 ;
        RECT 83.130 230.200 83.530 230.500 ;
        RECT 75.230 229.800 83.530 230.200 ;
        RECT 75.230 221.600 75.380 229.800 ;
        RECT 75.830 221.600 75.980 229.800 ;
        RECT 76.430 221.600 76.580 229.800 ;
        RECT 77.030 221.600 77.180 229.800 ;
        RECT 77.630 221.600 77.780 229.800 ;
        RECT 78.230 221.600 78.380 229.800 ;
        RECT 78.830 221.600 78.980 229.800 ;
        RECT 83.130 229.500 83.530 229.800 ;
        RECT 79.580 229.350 83.530 229.500 ;
        RECT 83.130 228.900 83.530 229.350 ;
        RECT 79.580 228.750 83.530 228.900 ;
        RECT 83.130 228.300 83.530 228.750 ;
        RECT 79.580 228.150 83.530 228.300 ;
        RECT 83.130 227.700 83.530 228.150 ;
        RECT 79.580 227.550 83.530 227.700 ;
        RECT 83.130 227.100 83.530 227.550 ;
        RECT 79.580 226.950 83.530 227.100 ;
        RECT 83.130 226.500 83.530 226.950 ;
        RECT 79.580 226.350 83.530 226.500 ;
        RECT 83.130 225.900 83.530 226.350 ;
        RECT 79.580 225.750 83.530 225.900 ;
        RECT 83.130 225.300 83.530 225.750 ;
        RECT 79.580 225.150 83.530 225.300 ;
        RECT 83.130 224.700 83.530 225.150 ;
        RECT 79.580 224.550 83.530 224.700 ;
        RECT 83.130 224.400 83.530 224.550 ;
        RECT 85.930 235.450 86.330 235.600 ;
        RECT 85.930 235.300 89.880 235.450 ;
        RECT 85.930 234.850 86.330 235.300 ;
        RECT 85.930 234.700 89.880 234.850 ;
        RECT 85.930 234.250 86.330 234.700 ;
        RECT 85.930 234.100 89.880 234.250 ;
        RECT 85.930 233.650 86.330 234.100 ;
        RECT 85.930 233.500 89.880 233.650 ;
        RECT 85.930 233.050 86.330 233.500 ;
        RECT 85.930 232.900 89.880 233.050 ;
        RECT 85.930 232.450 86.330 232.900 ;
        RECT 85.930 232.300 89.880 232.450 ;
        RECT 85.930 231.850 86.330 232.300 ;
        RECT 85.930 231.700 89.880 231.850 ;
        RECT 85.930 231.250 86.330 231.700 ;
        RECT 85.930 231.100 89.880 231.250 ;
        RECT 85.930 230.650 86.330 231.100 ;
        RECT 85.930 230.500 89.880 230.650 ;
        RECT 85.930 230.200 86.330 230.500 ;
        RECT 90.480 230.200 90.630 238.400 ;
        RECT 91.080 230.200 91.230 238.400 ;
        RECT 91.680 230.200 91.830 238.400 ;
        RECT 92.280 230.200 92.430 238.400 ;
        RECT 92.880 230.200 93.030 238.400 ;
        RECT 93.480 230.200 93.630 238.400 ;
        RECT 94.080 230.200 94.230 238.400 ;
        RECT 85.930 229.800 94.230 230.200 ;
        RECT 85.930 229.500 86.330 229.800 ;
        RECT 85.930 229.350 89.880 229.500 ;
        RECT 85.930 228.900 86.330 229.350 ;
        RECT 85.930 228.750 89.880 228.900 ;
        RECT 85.930 228.300 86.330 228.750 ;
        RECT 85.930 228.150 89.880 228.300 ;
        RECT 85.930 227.700 86.330 228.150 ;
        RECT 85.930 227.550 89.880 227.700 ;
        RECT 85.930 227.100 86.330 227.550 ;
        RECT 85.930 226.950 89.880 227.100 ;
        RECT 85.930 226.500 86.330 226.950 ;
        RECT 85.930 226.350 89.880 226.500 ;
        RECT 85.930 225.900 86.330 226.350 ;
        RECT 85.930 225.750 89.880 225.900 ;
        RECT 85.930 225.300 86.330 225.750 ;
        RECT 85.930 225.150 89.880 225.300 ;
        RECT 85.930 224.700 86.330 225.150 ;
        RECT 85.930 224.550 89.880 224.700 ;
        RECT 85.930 224.400 86.330 224.550 ;
        RECT 83.130 224.100 86.330 224.400 ;
        RECT 79.580 223.950 89.880 224.100 ;
        RECT 83.130 223.500 86.330 223.950 ;
        RECT 79.580 223.350 89.880 223.500 ;
        RECT 83.130 222.900 86.330 223.350 ;
        RECT 79.580 222.750 89.880 222.900 ;
        RECT 83.130 222.300 86.330 222.750 ;
        RECT 79.580 222.150 89.880 222.300 ;
        RECT 83.530 221.200 85.930 222.150 ;
        RECT 90.480 221.600 90.630 229.800 ;
        RECT 91.080 221.600 91.230 229.800 ;
        RECT 91.680 221.600 91.830 229.800 ;
        RECT 92.280 221.600 92.430 229.800 ;
        RECT 92.880 221.600 93.030 229.800 ;
        RECT 93.480 221.600 93.630 229.800 ;
        RECT 94.080 221.600 94.230 229.800 ;
        RECT 95.230 230.200 95.380 238.400 ;
        RECT 95.830 230.200 95.980 238.400 ;
        RECT 96.430 230.200 96.580 238.400 ;
        RECT 97.030 230.200 97.180 238.400 ;
        RECT 97.630 230.200 97.780 238.400 ;
        RECT 98.230 230.200 98.380 238.400 ;
        RECT 98.830 230.200 98.980 238.400 ;
        RECT 103.530 237.850 104.730 238.800 ;
        RECT 99.580 237.700 104.730 237.850 ;
        RECT 103.130 237.250 104.730 237.700 ;
        RECT 99.580 237.100 104.730 237.250 ;
        RECT 103.130 236.650 104.730 237.100 ;
        RECT 99.580 236.500 104.730 236.650 ;
        RECT 103.130 236.050 104.730 236.500 ;
        RECT 105.140 236.490 107.140 237.765 ;
        RECT 99.580 235.900 104.730 236.050 ;
        RECT 103.130 235.600 104.730 235.900 ;
        RECT 103.130 235.450 103.530 235.600 ;
        RECT 99.580 235.300 103.530 235.450 ;
        RECT 103.130 234.850 103.530 235.300 ;
        RECT 99.580 234.700 103.530 234.850 ;
        RECT 103.130 234.250 103.530 234.700 ;
        RECT 99.580 234.100 103.530 234.250 ;
        RECT 103.130 233.650 103.530 234.100 ;
        RECT 99.580 233.500 103.530 233.650 ;
        RECT 103.130 233.050 103.530 233.500 ;
        RECT 99.580 232.900 103.530 233.050 ;
        RECT 103.130 232.450 103.530 232.900 ;
        RECT 99.580 232.300 103.530 232.450 ;
        RECT 103.130 231.850 103.530 232.300 ;
        RECT 99.580 231.700 103.530 231.850 ;
        RECT 103.130 231.250 103.530 231.700 ;
        RECT 99.580 231.100 103.530 231.250 ;
        RECT 103.130 230.650 103.530 231.100 ;
        RECT 99.580 230.500 103.530 230.650 ;
        RECT 103.130 230.200 103.530 230.500 ;
        RECT 95.230 229.800 103.530 230.200 ;
        RECT 95.230 221.600 95.380 229.800 ;
        RECT 95.830 221.600 95.980 229.800 ;
        RECT 96.430 221.600 96.580 229.800 ;
        RECT 97.030 221.600 97.180 229.800 ;
        RECT 97.630 221.600 97.780 229.800 ;
        RECT 98.230 221.600 98.380 229.800 ;
        RECT 98.830 221.600 98.980 229.800 ;
        RECT 103.130 229.500 103.530 229.800 ;
        RECT 99.580 229.350 103.530 229.500 ;
        RECT 103.130 228.900 103.530 229.350 ;
        RECT 99.580 228.750 103.530 228.900 ;
        RECT 103.130 228.300 103.530 228.750 ;
        RECT 99.580 228.150 103.530 228.300 ;
        RECT 103.130 227.700 103.530 228.150 ;
        RECT 99.580 227.550 103.530 227.700 ;
        RECT 103.130 227.100 103.530 227.550 ;
        RECT 99.580 226.950 103.530 227.100 ;
        RECT 103.130 226.500 103.530 226.950 ;
        RECT 99.580 226.350 103.530 226.500 ;
        RECT 103.130 225.900 103.530 226.350 ;
        RECT 99.580 225.750 103.530 225.900 ;
        RECT 103.130 225.300 103.530 225.750 ;
        RECT 99.580 225.150 103.530 225.300 ;
        RECT 103.130 224.700 103.530 225.150 ;
        RECT 99.580 224.550 103.530 224.700 ;
        RECT 103.130 224.400 103.530 224.550 ;
        RECT 103.130 224.100 104.730 224.400 ;
        RECT 99.580 223.950 104.730 224.100 ;
        RECT 103.130 223.500 104.730 223.950 ;
        RECT 99.580 223.350 104.730 223.500 ;
        RECT 103.130 222.900 104.730 223.350 ;
        RECT 99.580 222.750 104.730 222.900 ;
        RECT 103.130 222.300 104.730 222.750 ;
        RECT 99.580 222.150 104.730 222.300 ;
        RECT 103.530 221.200 104.730 222.150 ;
        RECT 4.730 220.000 9.130 221.200 ;
        RECT 20.330 220.000 29.130 221.200 ;
        RECT 40.330 220.000 49.130 221.200 ;
        RECT 60.330 220.000 69.130 221.200 ;
        RECT 80.330 220.000 89.130 221.200 ;
        RECT 100.330 220.000 104.730 221.200 ;
        RECT 105.140 220.910 107.140 222.185 ;
        RECT 2.315 195.215 4.025 195.695 ;
        RECT 2.315 189.775 4.025 190.255 ;
        RECT 2.315 184.335 4.025 184.815 ;
        RECT 42.635 181.460 47.035 182.660 ;
        RECT 58.235 181.460 67.035 182.660 ;
        RECT 78.235 181.460 87.035 182.660 ;
        RECT 98.235 181.460 102.635 182.660 ;
        RECT 42.635 180.510 43.845 181.460 ;
        RECT 42.635 180.360 47.785 180.510 ;
        RECT 42.635 179.910 44.235 180.360 ;
        RECT 42.635 179.760 47.785 179.910 ;
        RECT 42.635 179.310 44.235 179.760 ;
        RECT 42.635 179.160 47.785 179.310 ;
        RECT 42.635 178.710 44.235 179.160 ;
        RECT 42.635 178.560 47.785 178.710 ;
        RECT 42.635 178.260 44.235 178.560 ;
        RECT 43.835 178.110 44.235 178.260 ;
        RECT 43.835 177.960 47.785 178.110 ;
        RECT 43.835 177.510 44.235 177.960 ;
        RECT 43.835 177.360 47.785 177.510 ;
        RECT 43.835 176.910 44.235 177.360 ;
        RECT 43.835 176.760 47.785 176.910 ;
        RECT 43.835 176.310 44.235 176.760 ;
        RECT 43.835 176.160 47.785 176.310 ;
        RECT 43.835 175.710 44.235 176.160 ;
        RECT 43.835 175.560 47.785 175.710 ;
        RECT 43.835 175.110 44.235 175.560 ;
        RECT 43.835 174.960 47.785 175.110 ;
        RECT 43.835 174.510 44.235 174.960 ;
        RECT 43.835 174.360 47.785 174.510 ;
        RECT 43.835 173.910 44.235 174.360 ;
        RECT 43.835 173.760 47.785 173.910 ;
        RECT 43.835 173.310 44.235 173.760 ;
        RECT 43.835 173.160 47.785 173.310 ;
        RECT 43.835 172.860 44.235 173.160 ;
        RECT 48.385 172.860 48.535 181.060 ;
        RECT 48.985 172.860 49.135 181.060 ;
        RECT 49.585 172.860 49.735 181.060 ;
        RECT 50.185 172.860 50.335 181.060 ;
        RECT 50.785 172.860 50.935 181.060 ;
        RECT 51.385 172.860 51.535 181.060 ;
        RECT 51.985 172.860 52.135 181.060 ;
        RECT 43.835 172.460 52.135 172.860 ;
        RECT 43.835 172.160 44.235 172.460 ;
        RECT 43.835 172.010 47.785 172.160 ;
        RECT 43.835 171.560 44.235 172.010 ;
        RECT 43.835 171.410 47.785 171.560 ;
        RECT 43.835 170.960 44.235 171.410 ;
        RECT 43.835 170.810 47.785 170.960 ;
        RECT 43.835 170.360 44.235 170.810 ;
        RECT 43.835 170.210 47.785 170.360 ;
        RECT 43.835 169.760 44.235 170.210 ;
        RECT 43.835 169.610 47.785 169.760 ;
        RECT 43.835 169.160 44.235 169.610 ;
        RECT 43.835 169.010 47.785 169.160 ;
        RECT 43.835 168.560 44.235 169.010 ;
        RECT 43.835 168.410 47.785 168.560 ;
        RECT 43.835 167.960 44.235 168.410 ;
        RECT 43.835 167.810 47.785 167.960 ;
        RECT 43.835 167.360 44.235 167.810 ;
        RECT 43.835 167.210 47.785 167.360 ;
        RECT 43.835 167.060 44.235 167.210 ;
        RECT 42.635 166.760 44.235 167.060 ;
        RECT 42.635 166.610 47.785 166.760 ;
        RECT 42.635 166.160 44.235 166.610 ;
        RECT 42.635 166.010 47.785 166.160 ;
        RECT 42.635 165.560 44.235 166.010 ;
        RECT 42.635 165.410 47.785 165.560 ;
        RECT 42.635 164.960 44.235 165.410 ;
        RECT 42.635 164.810 47.785 164.960 ;
        RECT 42.635 163.860 43.835 164.810 ;
        RECT 48.385 164.260 48.535 172.460 ;
        RECT 48.985 164.260 49.135 172.460 ;
        RECT 49.585 164.260 49.735 172.460 ;
        RECT 50.185 164.260 50.335 172.460 ;
        RECT 50.785 164.260 50.935 172.460 ;
        RECT 51.385 164.260 51.535 172.460 ;
        RECT 51.985 164.260 52.135 172.460 ;
        RECT 53.135 172.860 53.285 181.060 ;
        RECT 53.735 172.860 53.885 181.060 ;
        RECT 54.335 172.860 54.485 181.060 ;
        RECT 54.935 172.860 55.085 181.060 ;
        RECT 55.535 172.860 55.685 181.060 ;
        RECT 56.135 172.860 56.285 181.060 ;
        RECT 56.735 172.860 56.885 181.060 ;
        RECT 61.435 180.510 63.845 181.460 ;
        RECT 57.485 180.360 67.785 180.510 ;
        RECT 61.035 179.910 64.235 180.360 ;
        RECT 57.485 179.760 67.785 179.910 ;
        RECT 61.035 179.310 64.235 179.760 ;
        RECT 57.485 179.160 67.785 179.310 ;
        RECT 61.035 178.710 64.235 179.160 ;
        RECT 57.485 178.560 67.785 178.710 ;
        RECT 61.035 178.260 64.235 178.560 ;
        RECT 61.035 178.110 61.435 178.260 ;
        RECT 57.485 177.960 61.435 178.110 ;
        RECT 61.035 177.510 61.435 177.960 ;
        RECT 57.485 177.360 61.435 177.510 ;
        RECT 61.035 176.910 61.435 177.360 ;
        RECT 57.485 176.760 61.435 176.910 ;
        RECT 61.035 176.310 61.435 176.760 ;
        RECT 57.485 176.160 61.435 176.310 ;
        RECT 61.035 175.710 61.435 176.160 ;
        RECT 57.485 175.560 61.435 175.710 ;
        RECT 61.035 175.110 61.435 175.560 ;
        RECT 57.485 174.960 61.435 175.110 ;
        RECT 61.035 174.510 61.435 174.960 ;
        RECT 57.485 174.360 61.435 174.510 ;
        RECT 61.035 173.910 61.435 174.360 ;
        RECT 57.485 173.760 61.435 173.910 ;
        RECT 61.035 173.310 61.435 173.760 ;
        RECT 57.485 173.160 61.435 173.310 ;
        RECT 61.035 172.860 61.435 173.160 ;
        RECT 53.135 172.460 61.435 172.860 ;
        RECT 53.135 164.260 53.285 172.460 ;
        RECT 53.735 164.260 53.885 172.460 ;
        RECT 54.335 164.260 54.485 172.460 ;
        RECT 54.935 164.260 55.085 172.460 ;
        RECT 55.535 164.260 55.685 172.460 ;
        RECT 56.135 164.260 56.285 172.460 ;
        RECT 56.735 164.260 56.885 172.460 ;
        RECT 61.035 172.160 61.435 172.460 ;
        RECT 57.485 172.010 61.435 172.160 ;
        RECT 61.035 171.560 61.435 172.010 ;
        RECT 57.485 171.410 61.435 171.560 ;
        RECT 61.035 170.960 61.435 171.410 ;
        RECT 57.485 170.810 61.435 170.960 ;
        RECT 61.035 170.360 61.435 170.810 ;
        RECT 57.485 170.210 61.435 170.360 ;
        RECT 61.035 169.760 61.435 170.210 ;
        RECT 57.485 169.610 61.435 169.760 ;
        RECT 61.035 169.160 61.435 169.610 ;
        RECT 57.485 169.010 61.435 169.160 ;
        RECT 61.035 168.560 61.435 169.010 ;
        RECT 57.485 168.410 61.435 168.560 ;
        RECT 61.035 167.960 61.435 168.410 ;
        RECT 57.485 167.810 61.435 167.960 ;
        RECT 61.035 167.360 61.435 167.810 ;
        RECT 57.485 167.210 61.435 167.360 ;
        RECT 61.035 167.060 61.435 167.210 ;
        RECT 63.835 178.110 64.235 178.260 ;
        RECT 63.835 177.960 67.785 178.110 ;
        RECT 63.835 177.510 64.235 177.960 ;
        RECT 63.835 177.360 67.785 177.510 ;
        RECT 63.835 176.910 64.235 177.360 ;
        RECT 63.835 176.760 67.785 176.910 ;
        RECT 63.835 176.310 64.235 176.760 ;
        RECT 63.835 176.160 67.785 176.310 ;
        RECT 63.835 175.710 64.235 176.160 ;
        RECT 63.835 175.560 67.785 175.710 ;
        RECT 63.835 175.110 64.235 175.560 ;
        RECT 63.835 174.960 67.785 175.110 ;
        RECT 63.835 174.510 64.235 174.960 ;
        RECT 63.835 174.360 67.785 174.510 ;
        RECT 63.835 173.910 64.235 174.360 ;
        RECT 63.835 173.760 67.785 173.910 ;
        RECT 63.835 173.310 64.235 173.760 ;
        RECT 63.835 173.160 67.785 173.310 ;
        RECT 63.835 172.860 64.235 173.160 ;
        RECT 68.385 172.860 68.535 181.060 ;
        RECT 68.985 172.860 69.135 181.060 ;
        RECT 69.585 172.860 69.735 181.060 ;
        RECT 70.185 172.860 70.335 181.060 ;
        RECT 70.785 172.860 70.935 181.060 ;
        RECT 71.385 172.860 71.535 181.060 ;
        RECT 71.985 172.860 72.135 181.060 ;
        RECT 63.835 172.460 72.135 172.860 ;
        RECT 63.835 172.160 64.235 172.460 ;
        RECT 63.835 172.010 67.785 172.160 ;
        RECT 63.835 171.560 64.235 172.010 ;
        RECT 63.835 171.410 67.785 171.560 ;
        RECT 63.835 170.960 64.235 171.410 ;
        RECT 63.835 170.810 67.785 170.960 ;
        RECT 63.835 170.360 64.235 170.810 ;
        RECT 63.835 170.210 67.785 170.360 ;
        RECT 63.835 169.760 64.235 170.210 ;
        RECT 63.835 169.610 67.785 169.760 ;
        RECT 63.835 169.160 64.235 169.610 ;
        RECT 63.835 169.010 67.785 169.160 ;
        RECT 63.835 168.560 64.235 169.010 ;
        RECT 63.835 168.410 67.785 168.560 ;
        RECT 63.835 167.960 64.235 168.410 ;
        RECT 63.835 167.810 67.785 167.960 ;
        RECT 63.835 167.360 64.235 167.810 ;
        RECT 63.835 167.210 67.785 167.360 ;
        RECT 63.835 167.060 64.235 167.210 ;
        RECT 61.035 166.760 64.235 167.060 ;
        RECT 57.485 166.610 67.785 166.760 ;
        RECT 61.035 166.160 64.235 166.610 ;
        RECT 57.485 166.010 67.785 166.160 ;
        RECT 61.035 165.560 64.235 166.010 ;
        RECT 57.485 165.410 67.785 165.560 ;
        RECT 61.035 164.960 64.235 165.410 ;
        RECT 57.485 164.810 67.785 164.960 ;
        RECT 61.435 163.860 63.835 164.810 ;
        RECT 68.385 164.260 68.535 172.460 ;
        RECT 68.985 164.260 69.135 172.460 ;
        RECT 69.585 164.260 69.735 172.460 ;
        RECT 70.185 164.260 70.335 172.460 ;
        RECT 70.785 164.260 70.935 172.460 ;
        RECT 71.385 164.260 71.535 172.460 ;
        RECT 71.985 164.260 72.135 172.460 ;
        RECT 73.135 172.860 73.285 181.060 ;
        RECT 73.735 172.860 73.885 181.060 ;
        RECT 74.335 172.860 74.485 181.060 ;
        RECT 74.935 172.860 75.085 181.060 ;
        RECT 75.535 172.860 75.685 181.060 ;
        RECT 76.135 172.860 76.285 181.060 ;
        RECT 76.735 172.860 76.885 181.060 ;
        RECT 81.435 180.510 83.845 181.460 ;
        RECT 77.485 180.360 87.785 180.510 ;
        RECT 81.035 179.910 84.235 180.360 ;
        RECT 77.485 179.760 87.785 179.910 ;
        RECT 81.035 179.310 84.235 179.760 ;
        RECT 77.485 179.160 87.785 179.310 ;
        RECT 81.035 178.710 84.235 179.160 ;
        RECT 77.485 178.560 87.785 178.710 ;
        RECT 81.035 178.260 84.235 178.560 ;
        RECT 81.035 178.110 81.435 178.260 ;
        RECT 77.485 177.960 81.435 178.110 ;
        RECT 81.035 177.510 81.435 177.960 ;
        RECT 77.485 177.360 81.435 177.510 ;
        RECT 81.035 176.910 81.435 177.360 ;
        RECT 77.485 176.760 81.435 176.910 ;
        RECT 81.035 176.310 81.435 176.760 ;
        RECT 77.485 176.160 81.435 176.310 ;
        RECT 81.035 175.710 81.435 176.160 ;
        RECT 77.485 175.560 81.435 175.710 ;
        RECT 81.035 175.110 81.435 175.560 ;
        RECT 77.485 174.960 81.435 175.110 ;
        RECT 81.035 174.510 81.435 174.960 ;
        RECT 77.485 174.360 81.435 174.510 ;
        RECT 81.035 173.910 81.435 174.360 ;
        RECT 77.485 173.760 81.435 173.910 ;
        RECT 81.035 173.310 81.435 173.760 ;
        RECT 77.485 173.160 81.435 173.310 ;
        RECT 81.035 172.860 81.435 173.160 ;
        RECT 73.135 172.460 81.435 172.860 ;
        RECT 73.135 164.260 73.285 172.460 ;
        RECT 73.735 164.260 73.885 172.460 ;
        RECT 74.335 164.260 74.485 172.460 ;
        RECT 74.935 164.260 75.085 172.460 ;
        RECT 75.535 164.260 75.685 172.460 ;
        RECT 76.135 164.260 76.285 172.460 ;
        RECT 76.735 164.260 76.885 172.460 ;
        RECT 81.035 172.160 81.435 172.460 ;
        RECT 77.485 172.010 81.435 172.160 ;
        RECT 81.035 171.560 81.435 172.010 ;
        RECT 77.485 171.410 81.435 171.560 ;
        RECT 81.035 170.960 81.435 171.410 ;
        RECT 77.485 170.810 81.435 170.960 ;
        RECT 81.035 170.360 81.435 170.810 ;
        RECT 77.485 170.210 81.435 170.360 ;
        RECT 81.035 169.760 81.435 170.210 ;
        RECT 77.485 169.610 81.435 169.760 ;
        RECT 81.035 169.160 81.435 169.610 ;
        RECT 77.485 169.010 81.435 169.160 ;
        RECT 81.035 168.560 81.435 169.010 ;
        RECT 77.485 168.410 81.435 168.560 ;
        RECT 81.035 167.960 81.435 168.410 ;
        RECT 77.485 167.810 81.435 167.960 ;
        RECT 81.035 167.360 81.435 167.810 ;
        RECT 77.485 167.210 81.435 167.360 ;
        RECT 81.035 167.060 81.435 167.210 ;
        RECT 83.835 178.110 84.235 178.260 ;
        RECT 83.835 177.960 87.785 178.110 ;
        RECT 83.835 177.510 84.235 177.960 ;
        RECT 83.835 177.360 87.785 177.510 ;
        RECT 83.835 176.910 84.235 177.360 ;
        RECT 83.835 176.760 87.785 176.910 ;
        RECT 83.835 176.310 84.235 176.760 ;
        RECT 83.835 176.160 87.785 176.310 ;
        RECT 83.835 175.710 84.235 176.160 ;
        RECT 83.835 175.560 87.785 175.710 ;
        RECT 83.835 175.110 84.235 175.560 ;
        RECT 83.835 174.960 87.785 175.110 ;
        RECT 83.835 174.510 84.235 174.960 ;
        RECT 83.835 174.360 87.785 174.510 ;
        RECT 83.835 173.910 84.235 174.360 ;
        RECT 83.835 173.760 87.785 173.910 ;
        RECT 83.835 173.310 84.235 173.760 ;
        RECT 83.835 173.160 87.785 173.310 ;
        RECT 83.835 172.860 84.235 173.160 ;
        RECT 88.385 172.860 88.535 181.060 ;
        RECT 88.985 172.860 89.135 181.060 ;
        RECT 89.585 172.860 89.735 181.060 ;
        RECT 90.185 172.860 90.335 181.060 ;
        RECT 90.785 172.860 90.935 181.060 ;
        RECT 91.385 172.860 91.535 181.060 ;
        RECT 91.985 172.860 92.135 181.060 ;
        RECT 83.835 172.460 92.135 172.860 ;
        RECT 83.835 172.160 84.235 172.460 ;
        RECT 83.835 172.010 87.785 172.160 ;
        RECT 83.835 171.560 84.235 172.010 ;
        RECT 83.835 171.410 87.785 171.560 ;
        RECT 83.835 170.960 84.235 171.410 ;
        RECT 83.835 170.810 87.785 170.960 ;
        RECT 83.835 170.360 84.235 170.810 ;
        RECT 83.835 170.210 87.785 170.360 ;
        RECT 83.835 169.760 84.235 170.210 ;
        RECT 83.835 169.610 87.785 169.760 ;
        RECT 83.835 169.160 84.235 169.610 ;
        RECT 83.835 169.010 87.785 169.160 ;
        RECT 83.835 168.560 84.235 169.010 ;
        RECT 83.835 168.410 87.785 168.560 ;
        RECT 83.835 167.960 84.235 168.410 ;
        RECT 83.835 167.810 87.785 167.960 ;
        RECT 83.835 167.360 84.235 167.810 ;
        RECT 83.835 167.210 87.785 167.360 ;
        RECT 83.835 167.060 84.235 167.210 ;
        RECT 81.035 166.760 84.235 167.060 ;
        RECT 77.485 166.610 87.785 166.760 ;
        RECT 81.035 166.160 84.235 166.610 ;
        RECT 77.485 166.010 87.785 166.160 ;
        RECT 81.035 165.560 84.235 166.010 ;
        RECT 77.485 165.410 87.785 165.560 ;
        RECT 81.035 164.960 84.235 165.410 ;
        RECT 77.485 164.810 87.785 164.960 ;
        RECT 81.435 163.860 83.835 164.810 ;
        RECT 88.385 164.260 88.535 172.460 ;
        RECT 88.985 164.260 89.135 172.460 ;
        RECT 89.585 164.260 89.735 172.460 ;
        RECT 90.185 164.260 90.335 172.460 ;
        RECT 90.785 164.260 90.935 172.460 ;
        RECT 91.385 164.260 91.535 172.460 ;
        RECT 91.985 164.260 92.135 172.460 ;
        RECT 93.135 172.860 93.285 181.060 ;
        RECT 93.735 172.860 93.885 181.060 ;
        RECT 94.335 172.860 94.485 181.060 ;
        RECT 94.935 172.860 95.085 181.060 ;
        RECT 95.535 172.860 95.685 181.060 ;
        RECT 96.135 172.860 96.285 181.060 ;
        RECT 96.735 172.860 96.885 181.060 ;
        RECT 101.435 180.510 102.635 181.460 ;
        RECT 97.485 180.360 102.635 180.510 ;
        RECT 101.035 179.910 102.635 180.360 ;
        RECT 97.485 179.760 102.635 179.910 ;
        RECT 101.035 179.310 102.635 179.760 ;
        RECT 105.140 179.715 107.140 180.990 ;
        RECT 97.485 179.160 102.635 179.310 ;
        RECT 101.035 178.710 102.635 179.160 ;
        RECT 97.485 178.560 102.635 178.710 ;
        RECT 101.035 178.260 102.635 178.560 ;
        RECT 101.035 178.110 101.435 178.260 ;
        RECT 97.485 177.960 101.435 178.110 ;
        RECT 101.035 177.510 101.435 177.960 ;
        RECT 97.485 177.360 101.435 177.510 ;
        RECT 101.035 176.910 101.435 177.360 ;
        RECT 97.485 176.760 101.435 176.910 ;
        RECT 101.035 176.310 101.435 176.760 ;
        RECT 97.485 176.160 101.435 176.310 ;
        RECT 101.035 175.710 101.435 176.160 ;
        RECT 105.140 175.915 107.140 178.210 ;
        RECT 105.140 175.910 107.005 175.915 ;
        RECT 97.485 175.560 101.435 175.710 ;
        RECT 101.035 175.110 101.435 175.560 ;
        RECT 97.485 174.960 101.435 175.110 ;
        RECT 101.035 174.510 101.435 174.960 ;
        RECT 97.485 174.360 101.435 174.510 ;
        RECT 101.035 173.910 101.435 174.360 ;
        RECT 97.485 173.760 101.435 173.910 ;
        RECT 101.035 173.310 101.435 173.760 ;
        RECT 97.485 173.160 101.435 173.310 ;
        RECT 101.035 172.860 101.435 173.160 ;
        RECT 93.135 172.460 101.435 172.860 ;
        RECT 93.135 164.260 93.285 172.460 ;
        RECT 93.735 164.260 93.885 172.460 ;
        RECT 94.335 164.260 94.485 172.460 ;
        RECT 94.935 164.260 95.085 172.460 ;
        RECT 95.535 164.260 95.685 172.460 ;
        RECT 96.135 164.260 96.285 172.460 ;
        RECT 96.735 164.260 96.885 172.460 ;
        RECT 101.035 172.160 101.435 172.460 ;
        RECT 97.485 172.010 101.435 172.160 ;
        RECT 101.035 171.560 101.435 172.010 ;
        RECT 97.485 171.410 101.435 171.560 ;
        RECT 101.035 170.960 101.435 171.410 ;
        RECT 97.485 170.810 101.435 170.960 ;
        RECT 101.035 170.360 101.435 170.810 ;
        RECT 97.485 170.210 101.435 170.360 ;
        RECT 101.035 169.760 101.435 170.210 ;
        RECT 97.485 169.610 101.435 169.760 ;
        RECT 101.035 169.160 101.435 169.610 ;
        RECT 97.485 169.010 101.435 169.160 ;
        RECT 101.035 168.560 101.435 169.010 ;
        RECT 97.485 168.410 101.435 168.560 ;
        RECT 101.035 167.960 101.435 168.410 ;
        RECT 97.485 167.810 101.435 167.960 ;
        RECT 101.035 167.360 101.435 167.810 ;
        RECT 97.485 167.210 101.435 167.360 ;
        RECT 101.035 167.060 101.435 167.210 ;
        RECT 105.140 167.115 107.140 169.410 ;
        RECT 105.140 167.110 107.005 167.115 ;
        RECT 101.035 166.760 102.635 167.060 ;
        RECT 97.485 166.610 102.635 166.760 ;
        RECT 101.035 166.160 102.635 166.610 ;
        RECT 97.485 166.010 102.635 166.160 ;
        RECT 101.035 165.560 102.635 166.010 ;
        RECT 97.485 165.410 102.635 165.560 ;
        RECT 101.035 164.960 102.635 165.410 ;
        RECT 97.485 164.810 102.635 164.960 ;
        RECT 101.435 163.860 102.635 164.810 ;
        RECT 105.135 164.440 107.135 165.715 ;
        RECT 42.635 162.660 47.035 163.860 ;
        RECT 58.235 162.660 67.035 163.860 ;
        RECT 78.235 162.660 87.035 163.860 ;
        RECT 98.235 162.660 102.635 163.860 ;
        RECT 2.315 160.360 4.330 161.800 ;
        RECT 105.125 160.360 107.140 161.800 ;
        RECT 4.730 158.800 9.130 160.000 ;
        RECT 20.330 158.800 29.130 160.000 ;
        RECT 40.330 158.800 49.130 160.000 ;
        RECT 60.330 158.800 69.130 160.000 ;
        RECT 80.330 158.800 89.130 160.000 ;
        RECT 100.330 158.800 104.730 160.000 ;
        RECT 4.730 157.850 5.940 158.800 ;
        RECT 2.315 156.450 4.315 157.725 ;
        RECT 4.730 157.700 9.880 157.850 ;
        RECT 4.730 157.250 6.330 157.700 ;
        RECT 4.730 157.100 9.880 157.250 ;
        RECT 4.730 156.650 6.330 157.100 ;
        RECT 4.730 156.500 9.880 156.650 ;
        RECT 4.730 156.050 6.330 156.500 ;
        RECT 4.730 155.900 9.880 156.050 ;
        RECT 4.730 155.600 6.330 155.900 ;
        RECT 2.315 153.255 4.315 155.555 ;
        RECT 5.930 155.450 6.330 155.600 ;
        RECT 5.930 155.300 9.880 155.450 ;
        RECT 5.930 154.850 6.330 155.300 ;
        RECT 5.930 154.700 9.880 154.850 ;
        RECT 5.930 154.250 6.330 154.700 ;
        RECT 5.930 154.100 9.880 154.250 ;
        RECT 5.930 153.650 6.330 154.100 ;
        RECT 5.930 153.500 9.880 153.650 ;
        RECT 5.930 153.050 6.330 153.500 ;
        RECT 5.930 152.900 9.880 153.050 ;
        RECT 5.930 152.450 6.330 152.900 ;
        RECT 5.930 152.300 9.880 152.450 ;
        RECT 5.930 151.850 6.330 152.300 ;
        RECT 5.930 151.700 9.880 151.850 ;
        RECT 5.930 151.250 6.330 151.700 ;
        RECT 5.930 151.100 9.880 151.250 ;
        RECT 5.930 150.650 6.330 151.100 ;
        RECT 5.930 150.500 9.880 150.650 ;
        RECT 5.930 150.200 6.330 150.500 ;
        RECT 10.480 150.200 10.630 158.400 ;
        RECT 11.080 150.200 11.230 158.400 ;
        RECT 11.680 150.200 11.830 158.400 ;
        RECT 12.280 150.200 12.430 158.400 ;
        RECT 12.880 150.200 13.030 158.400 ;
        RECT 13.480 150.200 13.630 158.400 ;
        RECT 14.080 150.200 14.230 158.400 ;
        RECT 5.930 149.800 14.230 150.200 ;
        RECT 5.930 149.500 6.330 149.800 ;
        RECT 5.930 149.350 9.880 149.500 ;
        RECT 5.930 148.900 6.330 149.350 ;
        RECT 5.930 148.750 9.880 148.900 ;
        RECT 5.930 148.300 6.330 148.750 ;
        RECT 5.930 148.150 9.880 148.300 ;
        RECT 5.930 147.700 6.330 148.150 ;
        RECT 5.930 147.550 9.880 147.700 ;
        RECT 5.930 147.100 6.330 147.550 ;
        RECT 5.930 146.950 9.880 147.100 ;
        RECT 2.315 144.450 4.315 146.745 ;
        RECT 5.930 146.500 6.330 146.950 ;
        RECT 5.930 146.350 9.880 146.500 ;
        RECT 5.930 145.900 6.330 146.350 ;
        RECT 5.930 145.750 9.880 145.900 ;
        RECT 5.930 145.300 6.330 145.750 ;
        RECT 5.930 145.150 9.880 145.300 ;
        RECT 5.930 144.700 6.330 145.150 ;
        RECT 5.930 144.550 9.880 144.700 ;
        RECT 5.930 144.400 6.330 144.550 ;
        RECT 4.730 144.100 6.330 144.400 ;
        RECT 4.730 143.950 9.880 144.100 ;
        RECT 4.730 143.500 6.330 143.950 ;
        RECT 4.730 143.350 9.880 143.500 ;
        RECT 2.315 141.890 4.315 143.165 ;
        RECT 4.730 142.900 6.330 143.350 ;
        RECT 4.730 142.750 9.880 142.900 ;
        RECT 4.730 142.300 6.330 142.750 ;
        RECT 4.730 142.150 9.880 142.300 ;
        RECT 4.730 141.200 5.930 142.150 ;
        RECT 10.480 141.600 10.630 149.800 ;
        RECT 11.080 141.600 11.230 149.800 ;
        RECT 11.680 141.600 11.830 149.800 ;
        RECT 12.280 141.600 12.430 149.800 ;
        RECT 12.880 141.600 13.030 149.800 ;
        RECT 13.480 141.600 13.630 149.800 ;
        RECT 14.080 141.600 14.230 149.800 ;
        RECT 15.230 150.200 15.380 158.400 ;
        RECT 15.830 150.200 15.980 158.400 ;
        RECT 16.430 150.200 16.580 158.400 ;
        RECT 17.030 150.200 17.180 158.400 ;
        RECT 17.630 150.200 17.780 158.400 ;
        RECT 18.230 150.200 18.380 158.400 ;
        RECT 18.830 150.200 18.980 158.400 ;
        RECT 23.530 157.850 25.940 158.800 ;
        RECT 19.580 157.700 29.880 157.850 ;
        RECT 23.130 157.250 26.330 157.700 ;
        RECT 19.580 157.100 29.880 157.250 ;
        RECT 23.130 156.650 26.330 157.100 ;
        RECT 19.580 156.500 29.880 156.650 ;
        RECT 23.130 156.050 26.330 156.500 ;
        RECT 19.580 155.900 29.880 156.050 ;
        RECT 23.130 155.600 26.330 155.900 ;
        RECT 23.130 155.450 23.530 155.600 ;
        RECT 19.580 155.300 23.530 155.450 ;
        RECT 23.130 154.850 23.530 155.300 ;
        RECT 19.580 154.700 23.530 154.850 ;
        RECT 23.130 154.250 23.530 154.700 ;
        RECT 19.580 154.100 23.530 154.250 ;
        RECT 23.130 153.650 23.530 154.100 ;
        RECT 19.580 153.500 23.530 153.650 ;
        RECT 23.130 153.050 23.530 153.500 ;
        RECT 19.580 152.900 23.530 153.050 ;
        RECT 23.130 152.450 23.530 152.900 ;
        RECT 19.580 152.300 23.530 152.450 ;
        RECT 23.130 151.850 23.530 152.300 ;
        RECT 19.580 151.700 23.530 151.850 ;
        RECT 23.130 151.250 23.530 151.700 ;
        RECT 19.580 151.100 23.530 151.250 ;
        RECT 23.130 150.650 23.530 151.100 ;
        RECT 19.580 150.500 23.530 150.650 ;
        RECT 23.130 150.200 23.530 150.500 ;
        RECT 15.230 149.800 23.530 150.200 ;
        RECT 15.230 141.600 15.380 149.800 ;
        RECT 15.830 141.600 15.980 149.800 ;
        RECT 16.430 141.600 16.580 149.800 ;
        RECT 17.030 141.600 17.180 149.800 ;
        RECT 17.630 141.600 17.780 149.800 ;
        RECT 18.230 141.600 18.380 149.800 ;
        RECT 18.830 141.600 18.980 149.800 ;
        RECT 23.130 149.500 23.530 149.800 ;
        RECT 19.580 149.350 23.530 149.500 ;
        RECT 23.130 148.900 23.530 149.350 ;
        RECT 19.580 148.750 23.530 148.900 ;
        RECT 23.130 148.300 23.530 148.750 ;
        RECT 19.580 148.150 23.530 148.300 ;
        RECT 23.130 147.700 23.530 148.150 ;
        RECT 19.580 147.550 23.530 147.700 ;
        RECT 23.130 147.100 23.530 147.550 ;
        RECT 19.580 146.950 23.530 147.100 ;
        RECT 23.130 146.500 23.530 146.950 ;
        RECT 19.580 146.350 23.530 146.500 ;
        RECT 23.130 145.900 23.530 146.350 ;
        RECT 19.580 145.750 23.530 145.900 ;
        RECT 23.130 145.300 23.530 145.750 ;
        RECT 19.580 145.150 23.530 145.300 ;
        RECT 23.130 144.700 23.530 145.150 ;
        RECT 19.580 144.550 23.530 144.700 ;
        RECT 23.130 144.400 23.530 144.550 ;
        RECT 25.930 155.450 26.330 155.600 ;
        RECT 25.930 155.300 29.880 155.450 ;
        RECT 25.930 154.850 26.330 155.300 ;
        RECT 25.930 154.700 29.880 154.850 ;
        RECT 25.930 154.250 26.330 154.700 ;
        RECT 25.930 154.100 29.880 154.250 ;
        RECT 25.930 153.650 26.330 154.100 ;
        RECT 25.930 153.500 29.880 153.650 ;
        RECT 25.930 153.050 26.330 153.500 ;
        RECT 25.930 152.900 29.880 153.050 ;
        RECT 25.930 152.450 26.330 152.900 ;
        RECT 25.930 152.300 29.880 152.450 ;
        RECT 25.930 151.850 26.330 152.300 ;
        RECT 25.930 151.700 29.880 151.850 ;
        RECT 25.930 151.250 26.330 151.700 ;
        RECT 25.930 151.100 29.880 151.250 ;
        RECT 25.930 150.650 26.330 151.100 ;
        RECT 25.930 150.500 29.880 150.650 ;
        RECT 25.930 150.200 26.330 150.500 ;
        RECT 30.480 150.200 30.630 158.400 ;
        RECT 31.080 150.200 31.230 158.400 ;
        RECT 31.680 150.200 31.830 158.400 ;
        RECT 32.280 150.200 32.430 158.400 ;
        RECT 32.880 150.200 33.030 158.400 ;
        RECT 33.480 150.200 33.630 158.400 ;
        RECT 34.080 150.200 34.230 158.400 ;
        RECT 25.930 149.800 34.230 150.200 ;
        RECT 25.930 149.500 26.330 149.800 ;
        RECT 25.930 149.350 29.880 149.500 ;
        RECT 25.930 148.900 26.330 149.350 ;
        RECT 25.930 148.750 29.880 148.900 ;
        RECT 25.930 148.300 26.330 148.750 ;
        RECT 25.930 148.150 29.880 148.300 ;
        RECT 25.930 147.700 26.330 148.150 ;
        RECT 25.930 147.550 29.880 147.700 ;
        RECT 25.930 147.100 26.330 147.550 ;
        RECT 25.930 146.950 29.880 147.100 ;
        RECT 25.930 146.500 26.330 146.950 ;
        RECT 25.930 146.350 29.880 146.500 ;
        RECT 25.930 145.900 26.330 146.350 ;
        RECT 25.930 145.750 29.880 145.900 ;
        RECT 25.930 145.300 26.330 145.750 ;
        RECT 25.930 145.150 29.880 145.300 ;
        RECT 25.930 144.700 26.330 145.150 ;
        RECT 25.930 144.550 29.880 144.700 ;
        RECT 25.930 144.400 26.330 144.550 ;
        RECT 23.130 144.100 26.330 144.400 ;
        RECT 19.580 143.950 29.880 144.100 ;
        RECT 23.130 143.500 26.330 143.950 ;
        RECT 19.580 143.350 29.880 143.500 ;
        RECT 23.130 142.900 26.330 143.350 ;
        RECT 19.580 142.750 29.880 142.900 ;
        RECT 23.130 142.300 26.330 142.750 ;
        RECT 19.580 142.150 29.880 142.300 ;
        RECT 23.530 141.200 25.930 142.150 ;
        RECT 30.480 141.600 30.630 149.800 ;
        RECT 31.080 141.600 31.230 149.800 ;
        RECT 31.680 141.600 31.830 149.800 ;
        RECT 32.280 141.600 32.430 149.800 ;
        RECT 32.880 141.600 33.030 149.800 ;
        RECT 33.480 141.600 33.630 149.800 ;
        RECT 34.080 141.600 34.230 149.800 ;
        RECT 35.230 150.200 35.380 158.400 ;
        RECT 35.830 150.200 35.980 158.400 ;
        RECT 36.430 150.200 36.580 158.400 ;
        RECT 37.030 150.200 37.180 158.400 ;
        RECT 37.630 150.200 37.780 158.400 ;
        RECT 38.230 150.200 38.380 158.400 ;
        RECT 38.830 150.200 38.980 158.400 ;
        RECT 43.530 157.850 45.940 158.800 ;
        RECT 39.580 157.700 49.880 157.850 ;
        RECT 43.130 157.250 46.330 157.700 ;
        RECT 39.580 157.100 49.880 157.250 ;
        RECT 43.130 156.650 46.330 157.100 ;
        RECT 39.580 156.500 49.880 156.650 ;
        RECT 43.130 156.050 46.330 156.500 ;
        RECT 39.580 155.900 49.880 156.050 ;
        RECT 43.130 155.600 46.330 155.900 ;
        RECT 43.130 155.450 43.530 155.600 ;
        RECT 39.580 155.300 43.530 155.450 ;
        RECT 43.130 154.850 43.530 155.300 ;
        RECT 39.580 154.700 43.530 154.850 ;
        RECT 43.130 154.250 43.530 154.700 ;
        RECT 39.580 154.100 43.530 154.250 ;
        RECT 43.130 153.650 43.530 154.100 ;
        RECT 39.580 153.500 43.530 153.650 ;
        RECT 43.130 153.050 43.530 153.500 ;
        RECT 39.580 152.900 43.530 153.050 ;
        RECT 43.130 152.450 43.530 152.900 ;
        RECT 39.580 152.300 43.530 152.450 ;
        RECT 43.130 151.850 43.530 152.300 ;
        RECT 39.580 151.700 43.530 151.850 ;
        RECT 43.130 151.250 43.530 151.700 ;
        RECT 39.580 151.100 43.530 151.250 ;
        RECT 43.130 150.650 43.530 151.100 ;
        RECT 39.580 150.500 43.530 150.650 ;
        RECT 43.130 150.200 43.530 150.500 ;
        RECT 35.230 149.800 43.530 150.200 ;
        RECT 35.230 141.600 35.380 149.800 ;
        RECT 35.830 141.600 35.980 149.800 ;
        RECT 36.430 141.600 36.580 149.800 ;
        RECT 37.030 141.600 37.180 149.800 ;
        RECT 37.630 141.600 37.780 149.800 ;
        RECT 38.230 141.600 38.380 149.800 ;
        RECT 38.830 141.600 38.980 149.800 ;
        RECT 43.130 149.500 43.530 149.800 ;
        RECT 39.580 149.350 43.530 149.500 ;
        RECT 43.130 148.900 43.530 149.350 ;
        RECT 39.580 148.750 43.530 148.900 ;
        RECT 43.130 148.300 43.530 148.750 ;
        RECT 39.580 148.150 43.530 148.300 ;
        RECT 43.130 147.700 43.530 148.150 ;
        RECT 39.580 147.550 43.530 147.700 ;
        RECT 43.130 147.100 43.530 147.550 ;
        RECT 39.580 146.950 43.530 147.100 ;
        RECT 43.130 146.500 43.530 146.950 ;
        RECT 39.580 146.350 43.530 146.500 ;
        RECT 43.130 145.900 43.530 146.350 ;
        RECT 39.580 145.750 43.530 145.900 ;
        RECT 43.130 145.300 43.530 145.750 ;
        RECT 39.580 145.150 43.530 145.300 ;
        RECT 43.130 144.700 43.530 145.150 ;
        RECT 39.580 144.550 43.530 144.700 ;
        RECT 43.130 144.400 43.530 144.550 ;
        RECT 45.930 155.450 46.330 155.600 ;
        RECT 45.930 155.300 49.880 155.450 ;
        RECT 45.930 154.850 46.330 155.300 ;
        RECT 45.930 154.700 49.880 154.850 ;
        RECT 45.930 154.250 46.330 154.700 ;
        RECT 45.930 154.100 49.880 154.250 ;
        RECT 45.930 153.650 46.330 154.100 ;
        RECT 45.930 153.500 49.880 153.650 ;
        RECT 45.930 153.050 46.330 153.500 ;
        RECT 45.930 152.900 49.880 153.050 ;
        RECT 45.930 152.450 46.330 152.900 ;
        RECT 45.930 152.300 49.880 152.450 ;
        RECT 45.930 151.850 46.330 152.300 ;
        RECT 45.930 151.700 49.880 151.850 ;
        RECT 45.930 151.250 46.330 151.700 ;
        RECT 45.930 151.100 49.880 151.250 ;
        RECT 45.930 150.650 46.330 151.100 ;
        RECT 45.930 150.500 49.880 150.650 ;
        RECT 45.930 150.200 46.330 150.500 ;
        RECT 50.480 150.200 50.630 158.400 ;
        RECT 51.080 150.200 51.230 158.400 ;
        RECT 51.680 150.200 51.830 158.400 ;
        RECT 52.280 150.200 52.430 158.400 ;
        RECT 52.880 150.200 53.030 158.400 ;
        RECT 53.480 150.200 53.630 158.400 ;
        RECT 54.080 150.200 54.230 158.400 ;
        RECT 45.930 149.800 54.230 150.200 ;
        RECT 45.930 149.500 46.330 149.800 ;
        RECT 45.930 149.350 49.880 149.500 ;
        RECT 45.930 148.900 46.330 149.350 ;
        RECT 45.930 148.750 49.880 148.900 ;
        RECT 45.930 148.300 46.330 148.750 ;
        RECT 45.930 148.150 49.880 148.300 ;
        RECT 45.930 147.700 46.330 148.150 ;
        RECT 45.930 147.550 49.880 147.700 ;
        RECT 45.930 147.100 46.330 147.550 ;
        RECT 45.930 146.950 49.880 147.100 ;
        RECT 45.930 146.500 46.330 146.950 ;
        RECT 45.930 146.350 49.880 146.500 ;
        RECT 45.930 145.900 46.330 146.350 ;
        RECT 45.930 145.750 49.880 145.900 ;
        RECT 45.930 145.300 46.330 145.750 ;
        RECT 45.930 145.150 49.880 145.300 ;
        RECT 45.930 144.700 46.330 145.150 ;
        RECT 45.930 144.550 49.880 144.700 ;
        RECT 45.930 144.400 46.330 144.550 ;
        RECT 43.130 144.100 46.330 144.400 ;
        RECT 39.580 143.950 49.880 144.100 ;
        RECT 43.130 143.500 46.330 143.950 ;
        RECT 39.580 143.350 49.880 143.500 ;
        RECT 43.130 142.900 46.330 143.350 ;
        RECT 39.580 142.750 49.880 142.900 ;
        RECT 43.130 142.300 46.330 142.750 ;
        RECT 39.580 142.150 49.880 142.300 ;
        RECT 43.530 141.200 45.930 142.150 ;
        RECT 50.480 141.600 50.630 149.800 ;
        RECT 51.080 141.600 51.230 149.800 ;
        RECT 51.680 141.600 51.830 149.800 ;
        RECT 52.280 141.600 52.430 149.800 ;
        RECT 52.880 141.600 53.030 149.800 ;
        RECT 53.480 141.600 53.630 149.800 ;
        RECT 54.080 141.600 54.230 149.800 ;
        RECT 55.230 150.200 55.380 158.400 ;
        RECT 55.830 150.200 55.980 158.400 ;
        RECT 56.430 150.200 56.580 158.400 ;
        RECT 57.030 150.200 57.180 158.400 ;
        RECT 57.630 150.200 57.780 158.400 ;
        RECT 58.230 150.200 58.380 158.400 ;
        RECT 58.830 150.200 58.980 158.400 ;
        RECT 63.530 157.850 65.940 158.800 ;
        RECT 59.580 157.700 69.880 157.850 ;
        RECT 63.130 157.250 66.330 157.700 ;
        RECT 59.580 157.100 69.880 157.250 ;
        RECT 63.130 156.650 66.330 157.100 ;
        RECT 59.580 156.500 69.880 156.650 ;
        RECT 63.130 156.050 66.330 156.500 ;
        RECT 59.580 155.900 69.880 156.050 ;
        RECT 63.130 155.600 66.330 155.900 ;
        RECT 63.130 155.450 63.530 155.600 ;
        RECT 59.580 155.300 63.530 155.450 ;
        RECT 63.130 154.850 63.530 155.300 ;
        RECT 59.580 154.700 63.530 154.850 ;
        RECT 63.130 154.250 63.530 154.700 ;
        RECT 59.580 154.100 63.530 154.250 ;
        RECT 63.130 153.650 63.530 154.100 ;
        RECT 59.580 153.500 63.530 153.650 ;
        RECT 63.130 153.050 63.530 153.500 ;
        RECT 59.580 152.900 63.530 153.050 ;
        RECT 63.130 152.450 63.530 152.900 ;
        RECT 59.580 152.300 63.530 152.450 ;
        RECT 63.130 151.850 63.530 152.300 ;
        RECT 59.580 151.700 63.530 151.850 ;
        RECT 63.130 151.250 63.530 151.700 ;
        RECT 59.580 151.100 63.530 151.250 ;
        RECT 63.130 150.650 63.530 151.100 ;
        RECT 59.580 150.500 63.530 150.650 ;
        RECT 63.130 150.200 63.530 150.500 ;
        RECT 55.230 149.800 63.530 150.200 ;
        RECT 55.230 141.600 55.380 149.800 ;
        RECT 55.830 141.600 55.980 149.800 ;
        RECT 56.430 141.600 56.580 149.800 ;
        RECT 57.030 141.600 57.180 149.800 ;
        RECT 57.630 141.600 57.780 149.800 ;
        RECT 58.230 141.600 58.380 149.800 ;
        RECT 58.830 141.600 58.980 149.800 ;
        RECT 63.130 149.500 63.530 149.800 ;
        RECT 59.580 149.350 63.530 149.500 ;
        RECT 63.130 148.900 63.530 149.350 ;
        RECT 59.580 148.750 63.530 148.900 ;
        RECT 63.130 148.300 63.530 148.750 ;
        RECT 59.580 148.150 63.530 148.300 ;
        RECT 63.130 147.700 63.530 148.150 ;
        RECT 59.580 147.550 63.530 147.700 ;
        RECT 63.130 147.100 63.530 147.550 ;
        RECT 59.580 146.950 63.530 147.100 ;
        RECT 63.130 146.500 63.530 146.950 ;
        RECT 59.580 146.350 63.530 146.500 ;
        RECT 63.130 145.900 63.530 146.350 ;
        RECT 59.580 145.750 63.530 145.900 ;
        RECT 63.130 145.300 63.530 145.750 ;
        RECT 59.580 145.150 63.530 145.300 ;
        RECT 63.130 144.700 63.530 145.150 ;
        RECT 59.580 144.550 63.530 144.700 ;
        RECT 63.130 144.400 63.530 144.550 ;
        RECT 65.930 155.450 66.330 155.600 ;
        RECT 65.930 155.300 69.880 155.450 ;
        RECT 65.930 154.850 66.330 155.300 ;
        RECT 65.930 154.700 69.880 154.850 ;
        RECT 65.930 154.250 66.330 154.700 ;
        RECT 65.930 154.100 69.880 154.250 ;
        RECT 65.930 153.650 66.330 154.100 ;
        RECT 65.930 153.500 69.880 153.650 ;
        RECT 65.930 153.050 66.330 153.500 ;
        RECT 65.930 152.900 69.880 153.050 ;
        RECT 65.930 152.450 66.330 152.900 ;
        RECT 65.930 152.300 69.880 152.450 ;
        RECT 65.930 151.850 66.330 152.300 ;
        RECT 65.930 151.700 69.880 151.850 ;
        RECT 65.930 151.250 66.330 151.700 ;
        RECT 65.930 151.100 69.880 151.250 ;
        RECT 65.930 150.650 66.330 151.100 ;
        RECT 65.930 150.500 69.880 150.650 ;
        RECT 65.930 150.200 66.330 150.500 ;
        RECT 70.480 150.200 70.630 158.400 ;
        RECT 71.080 150.200 71.230 158.400 ;
        RECT 71.680 150.200 71.830 158.400 ;
        RECT 72.280 150.200 72.430 158.400 ;
        RECT 72.880 150.200 73.030 158.400 ;
        RECT 73.480 150.200 73.630 158.400 ;
        RECT 74.080 150.200 74.230 158.400 ;
        RECT 65.930 149.800 74.230 150.200 ;
        RECT 65.930 149.500 66.330 149.800 ;
        RECT 65.930 149.350 69.880 149.500 ;
        RECT 65.930 148.900 66.330 149.350 ;
        RECT 65.930 148.750 69.880 148.900 ;
        RECT 65.930 148.300 66.330 148.750 ;
        RECT 65.930 148.150 69.880 148.300 ;
        RECT 65.930 147.700 66.330 148.150 ;
        RECT 65.930 147.550 69.880 147.700 ;
        RECT 65.930 147.100 66.330 147.550 ;
        RECT 65.930 146.950 69.880 147.100 ;
        RECT 65.930 146.500 66.330 146.950 ;
        RECT 65.930 146.350 69.880 146.500 ;
        RECT 65.930 145.900 66.330 146.350 ;
        RECT 65.930 145.750 69.880 145.900 ;
        RECT 65.930 145.300 66.330 145.750 ;
        RECT 65.930 145.150 69.880 145.300 ;
        RECT 65.930 144.700 66.330 145.150 ;
        RECT 65.930 144.550 69.880 144.700 ;
        RECT 65.930 144.400 66.330 144.550 ;
        RECT 63.130 144.100 66.330 144.400 ;
        RECT 59.580 143.950 69.880 144.100 ;
        RECT 63.130 143.500 66.330 143.950 ;
        RECT 59.580 143.350 69.880 143.500 ;
        RECT 63.130 142.900 66.330 143.350 ;
        RECT 59.580 142.750 69.880 142.900 ;
        RECT 63.130 142.300 66.330 142.750 ;
        RECT 59.580 142.150 69.880 142.300 ;
        RECT 63.530 141.200 65.930 142.150 ;
        RECT 70.480 141.600 70.630 149.800 ;
        RECT 71.080 141.600 71.230 149.800 ;
        RECT 71.680 141.600 71.830 149.800 ;
        RECT 72.280 141.600 72.430 149.800 ;
        RECT 72.880 141.600 73.030 149.800 ;
        RECT 73.480 141.600 73.630 149.800 ;
        RECT 74.080 141.600 74.230 149.800 ;
        RECT 75.230 150.200 75.380 158.400 ;
        RECT 75.830 150.200 75.980 158.400 ;
        RECT 76.430 150.200 76.580 158.400 ;
        RECT 77.030 150.200 77.180 158.400 ;
        RECT 77.630 150.200 77.780 158.400 ;
        RECT 78.230 150.200 78.380 158.400 ;
        RECT 78.830 150.200 78.980 158.400 ;
        RECT 83.530 157.850 85.940 158.800 ;
        RECT 79.580 157.700 89.880 157.850 ;
        RECT 83.130 157.250 86.330 157.700 ;
        RECT 79.580 157.100 89.880 157.250 ;
        RECT 83.130 156.650 86.330 157.100 ;
        RECT 79.580 156.500 89.880 156.650 ;
        RECT 83.130 156.050 86.330 156.500 ;
        RECT 79.580 155.900 89.880 156.050 ;
        RECT 83.130 155.600 86.330 155.900 ;
        RECT 83.130 155.450 83.530 155.600 ;
        RECT 79.580 155.300 83.530 155.450 ;
        RECT 83.130 154.850 83.530 155.300 ;
        RECT 79.580 154.700 83.530 154.850 ;
        RECT 83.130 154.250 83.530 154.700 ;
        RECT 79.580 154.100 83.530 154.250 ;
        RECT 83.130 153.650 83.530 154.100 ;
        RECT 79.580 153.500 83.530 153.650 ;
        RECT 83.130 153.050 83.530 153.500 ;
        RECT 79.580 152.900 83.530 153.050 ;
        RECT 83.130 152.450 83.530 152.900 ;
        RECT 79.580 152.300 83.530 152.450 ;
        RECT 83.130 151.850 83.530 152.300 ;
        RECT 79.580 151.700 83.530 151.850 ;
        RECT 83.130 151.250 83.530 151.700 ;
        RECT 79.580 151.100 83.530 151.250 ;
        RECT 83.130 150.650 83.530 151.100 ;
        RECT 79.580 150.500 83.530 150.650 ;
        RECT 83.130 150.200 83.530 150.500 ;
        RECT 75.230 149.800 83.530 150.200 ;
        RECT 75.230 141.600 75.380 149.800 ;
        RECT 75.830 141.600 75.980 149.800 ;
        RECT 76.430 141.600 76.580 149.800 ;
        RECT 77.030 141.600 77.180 149.800 ;
        RECT 77.630 141.600 77.780 149.800 ;
        RECT 78.230 141.600 78.380 149.800 ;
        RECT 78.830 141.600 78.980 149.800 ;
        RECT 83.130 149.500 83.530 149.800 ;
        RECT 79.580 149.350 83.530 149.500 ;
        RECT 83.130 148.900 83.530 149.350 ;
        RECT 79.580 148.750 83.530 148.900 ;
        RECT 83.130 148.300 83.530 148.750 ;
        RECT 79.580 148.150 83.530 148.300 ;
        RECT 83.130 147.700 83.530 148.150 ;
        RECT 79.580 147.550 83.530 147.700 ;
        RECT 83.130 147.100 83.530 147.550 ;
        RECT 79.580 146.950 83.530 147.100 ;
        RECT 83.130 146.500 83.530 146.950 ;
        RECT 79.580 146.350 83.530 146.500 ;
        RECT 83.130 145.900 83.530 146.350 ;
        RECT 79.580 145.750 83.530 145.900 ;
        RECT 83.130 145.300 83.530 145.750 ;
        RECT 79.580 145.150 83.530 145.300 ;
        RECT 83.130 144.700 83.530 145.150 ;
        RECT 79.580 144.550 83.530 144.700 ;
        RECT 83.130 144.400 83.530 144.550 ;
        RECT 85.930 155.450 86.330 155.600 ;
        RECT 85.930 155.300 89.880 155.450 ;
        RECT 85.930 154.850 86.330 155.300 ;
        RECT 85.930 154.700 89.880 154.850 ;
        RECT 85.930 154.250 86.330 154.700 ;
        RECT 85.930 154.100 89.880 154.250 ;
        RECT 85.930 153.650 86.330 154.100 ;
        RECT 85.930 153.500 89.880 153.650 ;
        RECT 85.930 153.050 86.330 153.500 ;
        RECT 85.930 152.900 89.880 153.050 ;
        RECT 85.930 152.450 86.330 152.900 ;
        RECT 85.930 152.300 89.880 152.450 ;
        RECT 85.930 151.850 86.330 152.300 ;
        RECT 85.930 151.700 89.880 151.850 ;
        RECT 85.930 151.250 86.330 151.700 ;
        RECT 85.930 151.100 89.880 151.250 ;
        RECT 85.930 150.650 86.330 151.100 ;
        RECT 85.930 150.500 89.880 150.650 ;
        RECT 85.930 150.200 86.330 150.500 ;
        RECT 90.480 150.200 90.630 158.400 ;
        RECT 91.080 150.200 91.230 158.400 ;
        RECT 91.680 150.200 91.830 158.400 ;
        RECT 92.280 150.200 92.430 158.400 ;
        RECT 92.880 150.200 93.030 158.400 ;
        RECT 93.480 150.200 93.630 158.400 ;
        RECT 94.080 150.200 94.230 158.400 ;
        RECT 85.930 149.800 94.230 150.200 ;
        RECT 85.930 149.500 86.330 149.800 ;
        RECT 85.930 149.350 89.880 149.500 ;
        RECT 85.930 148.900 86.330 149.350 ;
        RECT 85.930 148.750 89.880 148.900 ;
        RECT 85.930 148.300 86.330 148.750 ;
        RECT 85.930 148.150 89.880 148.300 ;
        RECT 85.930 147.700 86.330 148.150 ;
        RECT 85.930 147.550 89.880 147.700 ;
        RECT 85.930 147.100 86.330 147.550 ;
        RECT 85.930 146.950 89.880 147.100 ;
        RECT 85.930 146.500 86.330 146.950 ;
        RECT 85.930 146.350 89.880 146.500 ;
        RECT 85.930 145.900 86.330 146.350 ;
        RECT 85.930 145.750 89.880 145.900 ;
        RECT 85.930 145.300 86.330 145.750 ;
        RECT 85.930 145.150 89.880 145.300 ;
        RECT 85.930 144.700 86.330 145.150 ;
        RECT 85.930 144.550 89.880 144.700 ;
        RECT 85.930 144.400 86.330 144.550 ;
        RECT 83.130 144.100 86.330 144.400 ;
        RECT 79.580 143.950 89.880 144.100 ;
        RECT 83.130 143.500 86.330 143.950 ;
        RECT 79.580 143.350 89.880 143.500 ;
        RECT 83.130 142.900 86.330 143.350 ;
        RECT 79.580 142.750 89.880 142.900 ;
        RECT 83.130 142.300 86.330 142.750 ;
        RECT 79.580 142.150 89.880 142.300 ;
        RECT 83.530 141.200 85.930 142.150 ;
        RECT 90.480 141.600 90.630 149.800 ;
        RECT 91.080 141.600 91.230 149.800 ;
        RECT 91.680 141.600 91.830 149.800 ;
        RECT 92.280 141.600 92.430 149.800 ;
        RECT 92.880 141.600 93.030 149.800 ;
        RECT 93.480 141.600 93.630 149.800 ;
        RECT 94.080 141.600 94.230 149.800 ;
        RECT 95.230 150.200 95.380 158.400 ;
        RECT 95.830 150.200 95.980 158.400 ;
        RECT 96.430 150.200 96.580 158.400 ;
        RECT 97.030 150.200 97.180 158.400 ;
        RECT 97.630 150.200 97.780 158.400 ;
        RECT 98.230 150.200 98.380 158.400 ;
        RECT 98.830 150.200 98.980 158.400 ;
        RECT 103.530 157.850 104.730 158.800 ;
        RECT 99.580 157.700 104.730 157.850 ;
        RECT 103.130 157.250 104.730 157.700 ;
        RECT 99.580 157.100 104.730 157.250 ;
        RECT 103.130 156.650 104.730 157.100 ;
        RECT 99.580 156.500 104.730 156.650 ;
        RECT 103.130 156.050 104.730 156.500 ;
        RECT 105.140 156.450 107.140 157.725 ;
        RECT 99.580 155.900 104.730 156.050 ;
        RECT 103.130 155.600 104.730 155.900 ;
        RECT 103.130 155.450 103.530 155.600 ;
        RECT 99.580 155.300 103.530 155.450 ;
        RECT 103.130 154.850 103.530 155.300 ;
        RECT 99.580 154.700 103.530 154.850 ;
        RECT 103.130 154.250 103.530 154.700 ;
        RECT 99.580 154.100 103.530 154.250 ;
        RECT 103.130 153.650 103.530 154.100 ;
        RECT 99.580 153.500 103.530 153.650 ;
        RECT 103.130 153.050 103.530 153.500 ;
        RECT 99.580 152.900 103.530 153.050 ;
        RECT 103.130 152.450 103.530 152.900 ;
        RECT 99.580 152.300 103.530 152.450 ;
        RECT 103.130 151.850 103.530 152.300 ;
        RECT 99.580 151.700 103.530 151.850 ;
        RECT 103.130 151.250 103.530 151.700 ;
        RECT 99.580 151.100 103.530 151.250 ;
        RECT 103.130 150.650 103.530 151.100 ;
        RECT 99.580 150.500 103.530 150.650 ;
        RECT 103.130 150.200 103.530 150.500 ;
        RECT 95.230 149.800 103.530 150.200 ;
        RECT 95.230 141.600 95.380 149.800 ;
        RECT 95.830 141.600 95.980 149.800 ;
        RECT 96.430 141.600 96.580 149.800 ;
        RECT 97.030 141.600 97.180 149.800 ;
        RECT 97.630 141.600 97.780 149.800 ;
        RECT 98.230 141.600 98.380 149.800 ;
        RECT 98.830 141.600 98.980 149.800 ;
        RECT 103.130 149.500 103.530 149.800 ;
        RECT 99.580 149.350 103.530 149.500 ;
        RECT 103.130 148.900 103.530 149.350 ;
        RECT 99.580 148.750 103.530 148.900 ;
        RECT 103.130 148.300 103.530 148.750 ;
        RECT 99.580 148.150 103.530 148.300 ;
        RECT 103.130 147.700 103.530 148.150 ;
        RECT 99.580 147.550 103.530 147.700 ;
        RECT 103.130 147.100 103.530 147.550 ;
        RECT 99.580 146.950 103.530 147.100 ;
        RECT 103.130 146.500 103.530 146.950 ;
        RECT 99.580 146.350 103.530 146.500 ;
        RECT 103.130 145.900 103.530 146.350 ;
        RECT 99.580 145.750 103.530 145.900 ;
        RECT 103.130 145.300 103.530 145.750 ;
        RECT 99.580 145.150 103.530 145.300 ;
        RECT 103.130 144.700 103.530 145.150 ;
        RECT 99.580 144.550 103.530 144.700 ;
        RECT 103.130 144.400 103.530 144.550 ;
        RECT 103.130 144.100 104.730 144.400 ;
        RECT 99.580 143.950 104.730 144.100 ;
        RECT 103.130 143.500 104.730 143.950 ;
        RECT 99.580 143.350 104.730 143.500 ;
        RECT 103.130 142.900 104.730 143.350 ;
        RECT 99.580 142.750 104.730 142.900 ;
        RECT 103.130 142.300 104.730 142.750 ;
        RECT 99.580 142.150 104.730 142.300 ;
        RECT 103.530 141.200 104.730 142.150 ;
        RECT 105.140 141.645 107.140 142.920 ;
        RECT 4.730 138.800 9.130 141.200 ;
        RECT 20.330 138.800 29.130 141.200 ;
        RECT 40.330 138.800 49.130 141.200 ;
        RECT 60.330 138.800 69.130 141.200 ;
        RECT 80.330 138.800 89.130 141.200 ;
        RECT 100.330 138.800 104.730 141.200 ;
        RECT 2.315 136.870 4.315 138.145 ;
        RECT 4.730 137.850 5.940 138.800 ;
        RECT 4.730 137.700 9.880 137.850 ;
        RECT 4.730 137.250 6.330 137.700 ;
        RECT 4.730 137.100 9.880 137.250 ;
        RECT 4.730 136.650 6.330 137.100 ;
        RECT 4.730 136.500 9.880 136.650 ;
        RECT 4.730 136.050 6.330 136.500 ;
        RECT 4.730 135.900 9.880 136.050 ;
        RECT 4.730 135.600 6.330 135.900 ;
        RECT 2.315 133.250 4.315 135.545 ;
        RECT 5.930 135.450 6.330 135.600 ;
        RECT 5.930 135.300 9.880 135.450 ;
        RECT 5.930 134.850 6.330 135.300 ;
        RECT 5.930 134.700 9.880 134.850 ;
        RECT 5.930 134.250 6.330 134.700 ;
        RECT 5.930 134.100 9.880 134.250 ;
        RECT 5.930 133.650 6.330 134.100 ;
        RECT 5.930 133.500 9.880 133.650 ;
        RECT 5.930 133.050 6.330 133.500 ;
        RECT 5.930 132.900 9.880 133.050 ;
        RECT 5.930 132.450 6.330 132.900 ;
        RECT 5.930 132.300 9.880 132.450 ;
        RECT 5.930 131.850 6.330 132.300 ;
        RECT 5.930 131.700 9.880 131.850 ;
        RECT 5.930 131.250 6.330 131.700 ;
        RECT 5.930 131.100 9.880 131.250 ;
        RECT 5.930 130.650 6.330 131.100 ;
        RECT 5.930 130.500 9.880 130.650 ;
        RECT 5.930 130.200 6.330 130.500 ;
        RECT 10.480 130.200 10.630 138.400 ;
        RECT 11.080 130.200 11.230 138.400 ;
        RECT 11.680 130.200 11.830 138.400 ;
        RECT 12.280 130.200 12.430 138.400 ;
        RECT 12.880 130.200 13.030 138.400 ;
        RECT 13.480 130.200 13.630 138.400 ;
        RECT 14.080 130.200 14.230 138.400 ;
        RECT 5.930 129.800 14.230 130.200 ;
        RECT 5.930 129.500 6.330 129.800 ;
        RECT 5.930 129.350 9.880 129.500 ;
        RECT 5.930 128.900 6.330 129.350 ;
        RECT 5.930 128.750 9.880 128.900 ;
        RECT 5.930 128.300 6.330 128.750 ;
        RECT 5.930 128.150 9.880 128.300 ;
        RECT 5.930 127.700 6.330 128.150 ;
        RECT 5.930 127.550 9.880 127.700 ;
        RECT 5.930 127.100 6.330 127.550 ;
        RECT 5.930 126.950 9.880 127.100 ;
        RECT 2.315 124.450 4.315 126.745 ;
        RECT 5.930 126.500 6.330 126.950 ;
        RECT 5.930 126.350 9.880 126.500 ;
        RECT 5.930 125.900 6.330 126.350 ;
        RECT 5.930 125.750 9.880 125.900 ;
        RECT 5.930 125.300 6.330 125.750 ;
        RECT 5.930 125.150 9.880 125.300 ;
        RECT 5.930 124.700 6.330 125.150 ;
        RECT 5.930 124.550 9.880 124.700 ;
        RECT 5.930 124.400 6.330 124.550 ;
        RECT 4.730 124.100 6.330 124.400 ;
        RECT 4.730 123.950 9.880 124.100 ;
        RECT 4.730 123.500 6.330 123.950 ;
        RECT 4.730 123.350 9.880 123.500 ;
        RECT 2.315 121.980 4.320 123.255 ;
        RECT 4.730 122.900 6.330 123.350 ;
        RECT 4.730 122.750 9.880 122.900 ;
        RECT 4.730 122.300 6.330 122.750 ;
        RECT 4.730 122.150 9.880 122.300 ;
        RECT 4.730 121.200 5.930 122.150 ;
        RECT 10.480 121.600 10.630 129.800 ;
        RECT 11.080 121.600 11.230 129.800 ;
        RECT 11.680 121.600 11.830 129.800 ;
        RECT 12.280 121.600 12.430 129.800 ;
        RECT 12.880 121.600 13.030 129.800 ;
        RECT 13.480 121.600 13.630 129.800 ;
        RECT 14.080 121.600 14.230 129.800 ;
        RECT 15.230 130.200 15.380 138.400 ;
        RECT 15.830 130.200 15.980 138.400 ;
        RECT 16.430 130.200 16.580 138.400 ;
        RECT 17.030 130.200 17.180 138.400 ;
        RECT 17.630 130.200 17.780 138.400 ;
        RECT 18.230 130.200 18.380 138.400 ;
        RECT 18.830 130.200 18.980 138.400 ;
        RECT 23.530 137.850 25.940 138.800 ;
        RECT 19.580 137.700 29.880 137.850 ;
        RECT 23.130 137.250 26.330 137.700 ;
        RECT 19.580 137.100 29.880 137.250 ;
        RECT 23.130 136.650 26.330 137.100 ;
        RECT 19.580 136.500 29.880 136.650 ;
        RECT 23.130 136.050 26.330 136.500 ;
        RECT 19.580 135.900 29.880 136.050 ;
        RECT 23.130 135.600 26.330 135.900 ;
        RECT 23.130 135.450 23.530 135.600 ;
        RECT 19.580 135.300 23.530 135.450 ;
        RECT 23.130 134.850 23.530 135.300 ;
        RECT 19.580 134.700 23.530 134.850 ;
        RECT 23.130 134.250 23.530 134.700 ;
        RECT 19.580 134.100 23.530 134.250 ;
        RECT 23.130 133.650 23.530 134.100 ;
        RECT 19.580 133.500 23.530 133.650 ;
        RECT 23.130 133.050 23.530 133.500 ;
        RECT 19.580 132.900 23.530 133.050 ;
        RECT 23.130 132.450 23.530 132.900 ;
        RECT 19.580 132.300 23.530 132.450 ;
        RECT 23.130 131.850 23.530 132.300 ;
        RECT 19.580 131.700 23.530 131.850 ;
        RECT 23.130 131.250 23.530 131.700 ;
        RECT 19.580 131.100 23.530 131.250 ;
        RECT 23.130 130.650 23.530 131.100 ;
        RECT 19.580 130.500 23.530 130.650 ;
        RECT 23.130 130.200 23.530 130.500 ;
        RECT 15.230 129.800 23.530 130.200 ;
        RECT 15.230 121.600 15.380 129.800 ;
        RECT 15.830 121.600 15.980 129.800 ;
        RECT 16.430 121.600 16.580 129.800 ;
        RECT 17.030 121.600 17.180 129.800 ;
        RECT 17.630 121.600 17.780 129.800 ;
        RECT 18.230 121.600 18.380 129.800 ;
        RECT 18.830 121.600 18.980 129.800 ;
        RECT 23.130 129.500 23.530 129.800 ;
        RECT 19.580 129.350 23.530 129.500 ;
        RECT 23.130 128.900 23.530 129.350 ;
        RECT 19.580 128.750 23.530 128.900 ;
        RECT 23.130 128.300 23.530 128.750 ;
        RECT 19.580 128.150 23.530 128.300 ;
        RECT 23.130 127.700 23.530 128.150 ;
        RECT 19.580 127.550 23.530 127.700 ;
        RECT 23.130 127.100 23.530 127.550 ;
        RECT 19.580 126.950 23.530 127.100 ;
        RECT 23.130 126.500 23.530 126.950 ;
        RECT 19.580 126.350 23.530 126.500 ;
        RECT 23.130 125.900 23.530 126.350 ;
        RECT 19.580 125.750 23.530 125.900 ;
        RECT 23.130 125.300 23.530 125.750 ;
        RECT 19.580 125.150 23.530 125.300 ;
        RECT 23.130 124.700 23.530 125.150 ;
        RECT 19.580 124.550 23.530 124.700 ;
        RECT 23.130 124.400 23.530 124.550 ;
        RECT 25.930 135.450 26.330 135.600 ;
        RECT 25.930 135.300 29.880 135.450 ;
        RECT 25.930 134.850 26.330 135.300 ;
        RECT 25.930 134.700 29.880 134.850 ;
        RECT 25.930 134.250 26.330 134.700 ;
        RECT 25.930 134.100 29.880 134.250 ;
        RECT 25.930 133.650 26.330 134.100 ;
        RECT 25.930 133.500 29.880 133.650 ;
        RECT 25.930 133.050 26.330 133.500 ;
        RECT 25.930 132.900 29.880 133.050 ;
        RECT 25.930 132.450 26.330 132.900 ;
        RECT 25.930 132.300 29.880 132.450 ;
        RECT 25.930 131.850 26.330 132.300 ;
        RECT 25.930 131.700 29.880 131.850 ;
        RECT 25.930 131.250 26.330 131.700 ;
        RECT 25.930 131.100 29.880 131.250 ;
        RECT 25.930 130.650 26.330 131.100 ;
        RECT 25.930 130.500 29.880 130.650 ;
        RECT 25.930 130.200 26.330 130.500 ;
        RECT 30.480 130.200 30.630 138.400 ;
        RECT 31.080 130.200 31.230 138.400 ;
        RECT 31.680 130.200 31.830 138.400 ;
        RECT 32.280 130.200 32.430 138.400 ;
        RECT 32.880 130.200 33.030 138.400 ;
        RECT 33.480 130.200 33.630 138.400 ;
        RECT 34.080 130.200 34.230 138.400 ;
        RECT 25.930 129.800 34.230 130.200 ;
        RECT 25.930 129.500 26.330 129.800 ;
        RECT 25.930 129.350 29.880 129.500 ;
        RECT 25.930 128.900 26.330 129.350 ;
        RECT 25.930 128.750 29.880 128.900 ;
        RECT 25.930 128.300 26.330 128.750 ;
        RECT 25.930 128.150 29.880 128.300 ;
        RECT 25.930 127.700 26.330 128.150 ;
        RECT 25.930 127.550 29.880 127.700 ;
        RECT 25.930 127.100 26.330 127.550 ;
        RECT 25.930 126.950 29.880 127.100 ;
        RECT 25.930 126.500 26.330 126.950 ;
        RECT 25.930 126.350 29.880 126.500 ;
        RECT 25.930 125.900 26.330 126.350 ;
        RECT 25.930 125.750 29.880 125.900 ;
        RECT 25.930 125.300 26.330 125.750 ;
        RECT 25.930 125.150 29.880 125.300 ;
        RECT 25.930 124.700 26.330 125.150 ;
        RECT 25.930 124.550 29.880 124.700 ;
        RECT 25.930 124.400 26.330 124.550 ;
        RECT 23.130 124.100 26.330 124.400 ;
        RECT 19.580 123.950 29.880 124.100 ;
        RECT 23.130 123.500 26.330 123.950 ;
        RECT 19.580 123.350 29.880 123.500 ;
        RECT 23.130 122.900 26.330 123.350 ;
        RECT 19.580 122.750 29.880 122.900 ;
        RECT 23.130 122.300 26.330 122.750 ;
        RECT 19.580 122.150 29.880 122.300 ;
        RECT 23.530 121.200 25.930 122.150 ;
        RECT 30.480 121.600 30.630 129.800 ;
        RECT 31.080 121.600 31.230 129.800 ;
        RECT 31.680 121.600 31.830 129.800 ;
        RECT 32.280 121.600 32.430 129.800 ;
        RECT 32.880 121.600 33.030 129.800 ;
        RECT 33.480 121.600 33.630 129.800 ;
        RECT 34.080 121.600 34.230 129.800 ;
        RECT 35.230 130.200 35.380 138.400 ;
        RECT 35.830 130.200 35.980 138.400 ;
        RECT 36.430 130.200 36.580 138.400 ;
        RECT 37.030 130.200 37.180 138.400 ;
        RECT 37.630 130.200 37.780 138.400 ;
        RECT 38.230 130.200 38.380 138.400 ;
        RECT 38.830 130.200 38.980 138.400 ;
        RECT 43.530 137.850 45.940 138.800 ;
        RECT 39.580 137.700 49.880 137.850 ;
        RECT 43.130 137.250 46.330 137.700 ;
        RECT 39.580 137.100 49.880 137.250 ;
        RECT 43.130 136.650 46.330 137.100 ;
        RECT 39.580 136.500 49.880 136.650 ;
        RECT 43.130 136.050 46.330 136.500 ;
        RECT 39.580 135.900 49.880 136.050 ;
        RECT 43.130 135.600 46.330 135.900 ;
        RECT 43.130 135.450 43.530 135.600 ;
        RECT 39.580 135.300 43.530 135.450 ;
        RECT 43.130 134.850 43.530 135.300 ;
        RECT 39.580 134.700 43.530 134.850 ;
        RECT 43.130 134.250 43.530 134.700 ;
        RECT 39.580 134.100 43.530 134.250 ;
        RECT 43.130 133.650 43.530 134.100 ;
        RECT 39.580 133.500 43.530 133.650 ;
        RECT 43.130 133.050 43.530 133.500 ;
        RECT 39.580 132.900 43.530 133.050 ;
        RECT 43.130 132.450 43.530 132.900 ;
        RECT 39.580 132.300 43.530 132.450 ;
        RECT 43.130 131.850 43.530 132.300 ;
        RECT 39.580 131.700 43.530 131.850 ;
        RECT 43.130 131.250 43.530 131.700 ;
        RECT 39.580 131.100 43.530 131.250 ;
        RECT 43.130 130.650 43.530 131.100 ;
        RECT 39.580 130.500 43.530 130.650 ;
        RECT 43.130 130.200 43.530 130.500 ;
        RECT 35.230 129.800 43.530 130.200 ;
        RECT 35.230 121.600 35.380 129.800 ;
        RECT 35.830 121.600 35.980 129.800 ;
        RECT 36.430 121.600 36.580 129.800 ;
        RECT 37.030 121.600 37.180 129.800 ;
        RECT 37.630 121.600 37.780 129.800 ;
        RECT 38.230 121.600 38.380 129.800 ;
        RECT 38.830 121.600 38.980 129.800 ;
        RECT 43.130 129.500 43.530 129.800 ;
        RECT 39.580 129.350 43.530 129.500 ;
        RECT 43.130 128.900 43.530 129.350 ;
        RECT 39.580 128.750 43.530 128.900 ;
        RECT 43.130 128.300 43.530 128.750 ;
        RECT 39.580 128.150 43.530 128.300 ;
        RECT 43.130 127.700 43.530 128.150 ;
        RECT 39.580 127.550 43.530 127.700 ;
        RECT 43.130 127.100 43.530 127.550 ;
        RECT 39.580 126.950 43.530 127.100 ;
        RECT 43.130 126.500 43.530 126.950 ;
        RECT 39.580 126.350 43.530 126.500 ;
        RECT 43.130 125.900 43.530 126.350 ;
        RECT 39.580 125.750 43.530 125.900 ;
        RECT 43.130 125.300 43.530 125.750 ;
        RECT 39.580 125.150 43.530 125.300 ;
        RECT 43.130 124.700 43.530 125.150 ;
        RECT 39.580 124.550 43.530 124.700 ;
        RECT 43.130 124.400 43.530 124.550 ;
        RECT 45.930 135.450 46.330 135.600 ;
        RECT 45.930 135.300 49.880 135.450 ;
        RECT 45.930 134.850 46.330 135.300 ;
        RECT 45.930 134.700 49.880 134.850 ;
        RECT 45.930 134.250 46.330 134.700 ;
        RECT 45.930 134.100 49.880 134.250 ;
        RECT 45.930 133.650 46.330 134.100 ;
        RECT 45.930 133.500 49.880 133.650 ;
        RECT 45.930 133.050 46.330 133.500 ;
        RECT 45.930 132.900 49.880 133.050 ;
        RECT 45.930 132.450 46.330 132.900 ;
        RECT 45.930 132.300 49.880 132.450 ;
        RECT 45.930 131.850 46.330 132.300 ;
        RECT 45.930 131.700 49.880 131.850 ;
        RECT 45.930 131.250 46.330 131.700 ;
        RECT 45.930 131.100 49.880 131.250 ;
        RECT 45.930 130.650 46.330 131.100 ;
        RECT 45.930 130.500 49.880 130.650 ;
        RECT 45.930 130.200 46.330 130.500 ;
        RECT 50.480 130.200 50.630 138.400 ;
        RECT 51.080 130.200 51.230 138.400 ;
        RECT 51.680 130.200 51.830 138.400 ;
        RECT 52.280 130.200 52.430 138.400 ;
        RECT 52.880 130.200 53.030 138.400 ;
        RECT 53.480 130.200 53.630 138.400 ;
        RECT 54.080 130.200 54.230 138.400 ;
        RECT 45.930 129.800 54.230 130.200 ;
        RECT 45.930 129.500 46.330 129.800 ;
        RECT 45.930 129.350 49.880 129.500 ;
        RECT 45.930 128.900 46.330 129.350 ;
        RECT 45.930 128.750 49.880 128.900 ;
        RECT 45.930 128.300 46.330 128.750 ;
        RECT 45.930 128.150 49.880 128.300 ;
        RECT 45.930 127.700 46.330 128.150 ;
        RECT 45.930 127.550 49.880 127.700 ;
        RECT 45.930 127.100 46.330 127.550 ;
        RECT 45.930 126.950 49.880 127.100 ;
        RECT 45.930 126.500 46.330 126.950 ;
        RECT 45.930 126.350 49.880 126.500 ;
        RECT 45.930 125.900 46.330 126.350 ;
        RECT 45.930 125.750 49.880 125.900 ;
        RECT 45.930 125.300 46.330 125.750 ;
        RECT 45.930 125.150 49.880 125.300 ;
        RECT 45.930 124.700 46.330 125.150 ;
        RECT 45.930 124.550 49.880 124.700 ;
        RECT 45.930 124.400 46.330 124.550 ;
        RECT 43.130 124.100 46.330 124.400 ;
        RECT 39.580 123.950 49.880 124.100 ;
        RECT 43.130 123.500 46.330 123.950 ;
        RECT 39.580 123.350 49.880 123.500 ;
        RECT 43.130 122.900 46.330 123.350 ;
        RECT 39.580 122.750 49.880 122.900 ;
        RECT 43.130 122.300 46.330 122.750 ;
        RECT 39.580 122.150 49.880 122.300 ;
        RECT 43.530 121.200 45.930 122.150 ;
        RECT 50.480 121.600 50.630 129.800 ;
        RECT 51.080 121.600 51.230 129.800 ;
        RECT 51.680 121.600 51.830 129.800 ;
        RECT 52.280 121.600 52.430 129.800 ;
        RECT 52.880 121.600 53.030 129.800 ;
        RECT 53.480 121.600 53.630 129.800 ;
        RECT 54.080 121.600 54.230 129.800 ;
        RECT 55.230 130.200 55.380 138.400 ;
        RECT 55.830 130.200 55.980 138.400 ;
        RECT 56.430 130.200 56.580 138.400 ;
        RECT 57.030 130.200 57.180 138.400 ;
        RECT 57.630 130.200 57.780 138.400 ;
        RECT 58.230 130.200 58.380 138.400 ;
        RECT 58.830 130.200 58.980 138.400 ;
        RECT 63.530 137.850 65.940 138.800 ;
        RECT 59.580 137.700 69.880 137.850 ;
        RECT 63.130 137.250 66.330 137.700 ;
        RECT 59.580 137.100 69.880 137.250 ;
        RECT 63.130 136.650 66.330 137.100 ;
        RECT 59.580 136.500 69.880 136.650 ;
        RECT 63.130 136.050 66.330 136.500 ;
        RECT 59.580 135.900 69.880 136.050 ;
        RECT 63.130 135.600 66.330 135.900 ;
        RECT 63.130 135.450 63.530 135.600 ;
        RECT 59.580 135.300 63.530 135.450 ;
        RECT 63.130 134.850 63.530 135.300 ;
        RECT 59.580 134.700 63.530 134.850 ;
        RECT 63.130 134.250 63.530 134.700 ;
        RECT 59.580 134.100 63.530 134.250 ;
        RECT 63.130 133.650 63.530 134.100 ;
        RECT 59.580 133.500 63.530 133.650 ;
        RECT 63.130 133.050 63.530 133.500 ;
        RECT 59.580 132.900 63.530 133.050 ;
        RECT 63.130 132.450 63.530 132.900 ;
        RECT 59.580 132.300 63.530 132.450 ;
        RECT 63.130 131.850 63.530 132.300 ;
        RECT 59.580 131.700 63.530 131.850 ;
        RECT 63.130 131.250 63.530 131.700 ;
        RECT 59.580 131.100 63.530 131.250 ;
        RECT 63.130 130.650 63.530 131.100 ;
        RECT 59.580 130.500 63.530 130.650 ;
        RECT 63.130 130.200 63.530 130.500 ;
        RECT 55.230 129.800 63.530 130.200 ;
        RECT 55.230 121.600 55.380 129.800 ;
        RECT 55.830 121.600 55.980 129.800 ;
        RECT 56.430 121.600 56.580 129.800 ;
        RECT 57.030 121.600 57.180 129.800 ;
        RECT 57.630 121.600 57.780 129.800 ;
        RECT 58.230 121.600 58.380 129.800 ;
        RECT 58.830 121.600 58.980 129.800 ;
        RECT 63.130 129.500 63.530 129.800 ;
        RECT 59.580 129.350 63.530 129.500 ;
        RECT 63.130 128.900 63.530 129.350 ;
        RECT 59.580 128.750 63.530 128.900 ;
        RECT 63.130 128.300 63.530 128.750 ;
        RECT 59.580 128.150 63.530 128.300 ;
        RECT 63.130 127.700 63.530 128.150 ;
        RECT 59.580 127.550 63.530 127.700 ;
        RECT 63.130 127.100 63.530 127.550 ;
        RECT 59.580 126.950 63.530 127.100 ;
        RECT 63.130 126.500 63.530 126.950 ;
        RECT 59.580 126.350 63.530 126.500 ;
        RECT 63.130 125.900 63.530 126.350 ;
        RECT 59.580 125.750 63.530 125.900 ;
        RECT 63.130 125.300 63.530 125.750 ;
        RECT 59.580 125.150 63.530 125.300 ;
        RECT 63.130 124.700 63.530 125.150 ;
        RECT 59.580 124.550 63.530 124.700 ;
        RECT 63.130 124.400 63.530 124.550 ;
        RECT 65.930 135.450 66.330 135.600 ;
        RECT 65.930 135.300 69.880 135.450 ;
        RECT 65.930 134.850 66.330 135.300 ;
        RECT 65.930 134.700 69.880 134.850 ;
        RECT 65.930 134.250 66.330 134.700 ;
        RECT 65.930 134.100 69.880 134.250 ;
        RECT 65.930 133.650 66.330 134.100 ;
        RECT 65.930 133.500 69.880 133.650 ;
        RECT 65.930 133.050 66.330 133.500 ;
        RECT 65.930 132.900 69.880 133.050 ;
        RECT 65.930 132.450 66.330 132.900 ;
        RECT 65.930 132.300 69.880 132.450 ;
        RECT 65.930 131.850 66.330 132.300 ;
        RECT 65.930 131.700 69.880 131.850 ;
        RECT 65.930 131.250 66.330 131.700 ;
        RECT 65.930 131.100 69.880 131.250 ;
        RECT 65.930 130.650 66.330 131.100 ;
        RECT 65.930 130.500 69.880 130.650 ;
        RECT 65.930 130.200 66.330 130.500 ;
        RECT 70.480 130.200 70.630 138.400 ;
        RECT 71.080 130.200 71.230 138.400 ;
        RECT 71.680 130.200 71.830 138.400 ;
        RECT 72.280 130.200 72.430 138.400 ;
        RECT 72.880 130.200 73.030 138.400 ;
        RECT 73.480 130.200 73.630 138.400 ;
        RECT 74.080 130.200 74.230 138.400 ;
        RECT 65.930 129.800 74.230 130.200 ;
        RECT 65.930 129.500 66.330 129.800 ;
        RECT 65.930 129.350 69.880 129.500 ;
        RECT 65.930 128.900 66.330 129.350 ;
        RECT 65.930 128.750 69.880 128.900 ;
        RECT 65.930 128.300 66.330 128.750 ;
        RECT 65.930 128.150 69.880 128.300 ;
        RECT 65.930 127.700 66.330 128.150 ;
        RECT 65.930 127.550 69.880 127.700 ;
        RECT 65.930 127.100 66.330 127.550 ;
        RECT 65.930 126.950 69.880 127.100 ;
        RECT 65.930 126.500 66.330 126.950 ;
        RECT 65.930 126.350 69.880 126.500 ;
        RECT 65.930 125.900 66.330 126.350 ;
        RECT 65.930 125.750 69.880 125.900 ;
        RECT 65.930 125.300 66.330 125.750 ;
        RECT 65.930 125.150 69.880 125.300 ;
        RECT 65.930 124.700 66.330 125.150 ;
        RECT 65.930 124.550 69.880 124.700 ;
        RECT 65.930 124.400 66.330 124.550 ;
        RECT 63.130 124.100 66.330 124.400 ;
        RECT 59.580 123.950 69.880 124.100 ;
        RECT 63.130 123.500 66.330 123.950 ;
        RECT 59.580 123.350 69.880 123.500 ;
        RECT 63.130 122.900 66.330 123.350 ;
        RECT 59.580 122.750 69.880 122.900 ;
        RECT 63.130 122.300 66.330 122.750 ;
        RECT 59.580 122.150 69.880 122.300 ;
        RECT 63.530 121.200 65.930 122.150 ;
        RECT 70.480 121.600 70.630 129.800 ;
        RECT 71.080 121.600 71.230 129.800 ;
        RECT 71.680 121.600 71.830 129.800 ;
        RECT 72.280 121.600 72.430 129.800 ;
        RECT 72.880 121.600 73.030 129.800 ;
        RECT 73.480 121.600 73.630 129.800 ;
        RECT 74.080 121.600 74.230 129.800 ;
        RECT 75.230 130.200 75.380 138.400 ;
        RECT 75.830 130.200 75.980 138.400 ;
        RECT 76.430 130.200 76.580 138.400 ;
        RECT 77.030 130.200 77.180 138.400 ;
        RECT 77.630 130.200 77.780 138.400 ;
        RECT 78.230 130.200 78.380 138.400 ;
        RECT 78.830 130.200 78.980 138.400 ;
        RECT 83.530 137.850 85.940 138.800 ;
        RECT 79.580 137.700 89.880 137.850 ;
        RECT 83.130 137.250 86.330 137.700 ;
        RECT 79.580 137.100 89.880 137.250 ;
        RECT 83.130 136.650 86.330 137.100 ;
        RECT 79.580 136.500 89.880 136.650 ;
        RECT 83.130 136.050 86.330 136.500 ;
        RECT 79.580 135.900 89.880 136.050 ;
        RECT 83.130 135.600 86.330 135.900 ;
        RECT 83.130 135.450 83.530 135.600 ;
        RECT 79.580 135.300 83.530 135.450 ;
        RECT 83.130 134.850 83.530 135.300 ;
        RECT 79.580 134.700 83.530 134.850 ;
        RECT 83.130 134.250 83.530 134.700 ;
        RECT 79.580 134.100 83.530 134.250 ;
        RECT 83.130 133.650 83.530 134.100 ;
        RECT 79.580 133.500 83.530 133.650 ;
        RECT 83.130 133.050 83.530 133.500 ;
        RECT 79.580 132.900 83.530 133.050 ;
        RECT 83.130 132.450 83.530 132.900 ;
        RECT 79.580 132.300 83.530 132.450 ;
        RECT 83.130 131.850 83.530 132.300 ;
        RECT 79.580 131.700 83.530 131.850 ;
        RECT 83.130 131.250 83.530 131.700 ;
        RECT 79.580 131.100 83.530 131.250 ;
        RECT 83.130 130.650 83.530 131.100 ;
        RECT 79.580 130.500 83.530 130.650 ;
        RECT 83.130 130.200 83.530 130.500 ;
        RECT 75.230 129.800 83.530 130.200 ;
        RECT 75.230 121.600 75.380 129.800 ;
        RECT 75.830 121.600 75.980 129.800 ;
        RECT 76.430 121.600 76.580 129.800 ;
        RECT 77.030 121.600 77.180 129.800 ;
        RECT 77.630 121.600 77.780 129.800 ;
        RECT 78.230 121.600 78.380 129.800 ;
        RECT 78.830 121.600 78.980 129.800 ;
        RECT 83.130 129.500 83.530 129.800 ;
        RECT 79.580 129.350 83.530 129.500 ;
        RECT 83.130 128.900 83.530 129.350 ;
        RECT 79.580 128.750 83.530 128.900 ;
        RECT 83.130 128.300 83.530 128.750 ;
        RECT 79.580 128.150 83.530 128.300 ;
        RECT 83.130 127.700 83.530 128.150 ;
        RECT 79.580 127.550 83.530 127.700 ;
        RECT 83.130 127.100 83.530 127.550 ;
        RECT 79.580 126.950 83.530 127.100 ;
        RECT 83.130 126.500 83.530 126.950 ;
        RECT 79.580 126.350 83.530 126.500 ;
        RECT 83.130 125.900 83.530 126.350 ;
        RECT 79.580 125.750 83.530 125.900 ;
        RECT 83.130 125.300 83.530 125.750 ;
        RECT 79.580 125.150 83.530 125.300 ;
        RECT 83.130 124.700 83.530 125.150 ;
        RECT 79.580 124.550 83.530 124.700 ;
        RECT 83.130 124.400 83.530 124.550 ;
        RECT 85.930 135.450 86.330 135.600 ;
        RECT 85.930 135.300 89.880 135.450 ;
        RECT 85.930 134.850 86.330 135.300 ;
        RECT 85.930 134.700 89.880 134.850 ;
        RECT 85.930 134.250 86.330 134.700 ;
        RECT 85.930 134.100 89.880 134.250 ;
        RECT 85.930 133.650 86.330 134.100 ;
        RECT 85.930 133.500 89.880 133.650 ;
        RECT 85.930 133.050 86.330 133.500 ;
        RECT 85.930 132.900 89.880 133.050 ;
        RECT 85.930 132.450 86.330 132.900 ;
        RECT 85.930 132.300 89.880 132.450 ;
        RECT 85.930 131.850 86.330 132.300 ;
        RECT 85.930 131.700 89.880 131.850 ;
        RECT 85.930 131.250 86.330 131.700 ;
        RECT 85.930 131.100 89.880 131.250 ;
        RECT 85.930 130.650 86.330 131.100 ;
        RECT 85.930 130.500 89.880 130.650 ;
        RECT 85.930 130.200 86.330 130.500 ;
        RECT 90.480 130.200 90.630 138.400 ;
        RECT 91.080 130.200 91.230 138.400 ;
        RECT 91.680 130.200 91.830 138.400 ;
        RECT 92.280 130.200 92.430 138.400 ;
        RECT 92.880 130.200 93.030 138.400 ;
        RECT 93.480 130.200 93.630 138.400 ;
        RECT 94.080 130.200 94.230 138.400 ;
        RECT 85.930 129.800 94.230 130.200 ;
        RECT 85.930 129.500 86.330 129.800 ;
        RECT 85.930 129.350 89.880 129.500 ;
        RECT 85.930 128.900 86.330 129.350 ;
        RECT 85.930 128.750 89.880 128.900 ;
        RECT 85.930 128.300 86.330 128.750 ;
        RECT 85.930 128.150 89.880 128.300 ;
        RECT 85.930 127.700 86.330 128.150 ;
        RECT 85.930 127.550 89.880 127.700 ;
        RECT 85.930 127.100 86.330 127.550 ;
        RECT 85.930 126.950 89.880 127.100 ;
        RECT 85.930 126.500 86.330 126.950 ;
        RECT 85.930 126.350 89.880 126.500 ;
        RECT 85.930 125.900 86.330 126.350 ;
        RECT 85.930 125.750 89.880 125.900 ;
        RECT 85.930 125.300 86.330 125.750 ;
        RECT 85.930 125.150 89.880 125.300 ;
        RECT 85.930 124.700 86.330 125.150 ;
        RECT 85.930 124.550 89.880 124.700 ;
        RECT 85.930 124.400 86.330 124.550 ;
        RECT 83.130 124.100 86.330 124.400 ;
        RECT 79.580 123.950 89.880 124.100 ;
        RECT 83.130 123.500 86.330 123.950 ;
        RECT 79.580 123.350 89.880 123.500 ;
        RECT 83.130 122.900 86.330 123.350 ;
        RECT 79.580 122.750 89.880 122.900 ;
        RECT 83.130 122.300 86.330 122.750 ;
        RECT 79.580 122.150 89.880 122.300 ;
        RECT 83.530 121.200 85.930 122.150 ;
        RECT 90.480 121.600 90.630 129.800 ;
        RECT 91.080 121.600 91.230 129.800 ;
        RECT 91.680 121.600 91.830 129.800 ;
        RECT 92.280 121.600 92.430 129.800 ;
        RECT 92.880 121.600 93.030 129.800 ;
        RECT 93.480 121.600 93.630 129.800 ;
        RECT 94.080 121.600 94.230 129.800 ;
        RECT 95.230 130.200 95.380 138.400 ;
        RECT 95.830 130.200 95.980 138.400 ;
        RECT 96.430 130.200 96.580 138.400 ;
        RECT 97.030 130.200 97.180 138.400 ;
        RECT 97.630 130.200 97.780 138.400 ;
        RECT 98.230 130.200 98.380 138.400 ;
        RECT 98.830 130.200 98.980 138.400 ;
        RECT 103.530 137.850 104.730 138.800 ;
        RECT 99.580 137.700 104.730 137.850 ;
        RECT 103.130 137.250 104.730 137.700 ;
        RECT 99.580 137.100 104.730 137.250 ;
        RECT 103.130 136.650 104.730 137.100 ;
        RECT 99.580 136.500 104.730 136.650 ;
        RECT 103.130 136.050 104.730 136.500 ;
        RECT 105.135 136.060 107.135 137.335 ;
        RECT 99.580 135.900 104.730 136.050 ;
        RECT 103.130 135.600 104.730 135.900 ;
        RECT 103.130 135.450 103.530 135.600 ;
        RECT 99.580 135.300 103.530 135.450 ;
        RECT 103.130 134.850 103.530 135.300 ;
        RECT 99.580 134.700 103.530 134.850 ;
        RECT 103.130 134.250 103.530 134.700 ;
        RECT 99.580 134.100 103.530 134.250 ;
        RECT 103.130 133.650 103.530 134.100 ;
        RECT 99.580 133.500 103.530 133.650 ;
        RECT 103.130 133.050 103.530 133.500 ;
        RECT 99.580 132.900 103.530 133.050 ;
        RECT 103.130 132.450 103.530 132.900 ;
        RECT 99.580 132.300 103.530 132.450 ;
        RECT 103.130 131.850 103.530 132.300 ;
        RECT 99.580 131.700 103.530 131.850 ;
        RECT 103.130 131.250 103.530 131.700 ;
        RECT 99.580 131.100 103.530 131.250 ;
        RECT 103.130 130.650 103.530 131.100 ;
        RECT 99.580 130.500 103.530 130.650 ;
        RECT 103.130 130.200 103.530 130.500 ;
        RECT 95.230 129.800 103.530 130.200 ;
        RECT 95.230 121.600 95.380 129.800 ;
        RECT 95.830 121.600 95.980 129.800 ;
        RECT 96.430 121.600 96.580 129.800 ;
        RECT 97.030 121.600 97.180 129.800 ;
        RECT 97.630 121.600 97.780 129.800 ;
        RECT 98.230 121.600 98.380 129.800 ;
        RECT 98.830 121.600 98.980 129.800 ;
        RECT 103.130 129.500 103.530 129.800 ;
        RECT 99.580 129.350 103.530 129.500 ;
        RECT 103.130 128.900 103.530 129.350 ;
        RECT 99.580 128.750 103.530 128.900 ;
        RECT 103.130 128.300 103.530 128.750 ;
        RECT 99.580 128.150 103.530 128.300 ;
        RECT 103.130 127.700 103.530 128.150 ;
        RECT 99.580 127.550 103.530 127.700 ;
        RECT 103.130 127.100 103.530 127.550 ;
        RECT 99.580 126.950 103.530 127.100 ;
        RECT 103.130 126.500 103.530 126.950 ;
        RECT 99.580 126.350 103.530 126.500 ;
        RECT 103.130 125.900 103.530 126.350 ;
        RECT 99.580 125.750 103.530 125.900 ;
        RECT 103.130 125.300 103.530 125.750 ;
        RECT 99.580 125.150 103.530 125.300 ;
        RECT 103.130 124.700 103.530 125.150 ;
        RECT 99.580 124.550 103.530 124.700 ;
        RECT 103.130 124.400 103.530 124.550 ;
        RECT 103.130 124.100 104.730 124.400 ;
        RECT 99.580 123.950 104.730 124.100 ;
        RECT 103.130 123.500 104.730 123.950 ;
        RECT 99.580 123.350 104.730 123.500 ;
        RECT 103.130 122.900 104.730 123.350 ;
        RECT 99.580 122.750 104.730 122.900 ;
        RECT 103.130 122.300 104.730 122.750 ;
        RECT 99.580 122.150 104.730 122.300 ;
        RECT 103.530 121.200 104.730 122.150 ;
        RECT 105.140 121.845 107.140 123.120 ;
        RECT 4.730 118.800 9.130 121.200 ;
        RECT 20.330 118.800 29.130 121.200 ;
        RECT 40.330 118.800 49.130 121.200 ;
        RECT 60.330 118.800 69.130 121.200 ;
        RECT 80.330 118.800 89.130 121.200 ;
        RECT 100.330 118.800 104.730 121.200 ;
        RECT 4.730 117.850 5.940 118.800 ;
        RECT 2.315 116.570 4.320 117.845 ;
        RECT 4.730 117.700 9.880 117.850 ;
        RECT 4.730 117.250 6.330 117.700 ;
        RECT 4.730 117.100 9.880 117.250 ;
        RECT 4.730 116.650 6.330 117.100 ;
        RECT 4.730 116.500 9.880 116.650 ;
        RECT 4.730 116.050 6.330 116.500 ;
        RECT 4.730 115.900 9.880 116.050 ;
        RECT 4.730 115.600 6.330 115.900 ;
        RECT 2.315 113.250 4.315 115.545 ;
        RECT 5.930 115.450 6.330 115.600 ;
        RECT 5.930 115.300 9.880 115.450 ;
        RECT 5.930 114.850 6.330 115.300 ;
        RECT 5.930 114.700 9.880 114.850 ;
        RECT 5.930 114.250 6.330 114.700 ;
        RECT 5.930 114.100 9.880 114.250 ;
        RECT 5.930 113.650 6.330 114.100 ;
        RECT 5.930 113.500 9.880 113.650 ;
        RECT 5.930 113.050 6.330 113.500 ;
        RECT 5.930 112.900 9.880 113.050 ;
        RECT 5.930 112.450 6.330 112.900 ;
        RECT 5.930 112.300 9.880 112.450 ;
        RECT 5.930 111.850 6.330 112.300 ;
        RECT 5.930 111.700 9.880 111.850 ;
        RECT 5.930 111.250 6.330 111.700 ;
        RECT 5.930 111.100 9.880 111.250 ;
        RECT 5.930 110.650 6.330 111.100 ;
        RECT 5.930 110.500 9.880 110.650 ;
        RECT 5.930 110.200 6.330 110.500 ;
        RECT 10.480 110.200 10.630 118.400 ;
        RECT 11.080 110.200 11.230 118.400 ;
        RECT 11.680 110.200 11.830 118.400 ;
        RECT 12.280 110.200 12.430 118.400 ;
        RECT 12.880 110.200 13.030 118.400 ;
        RECT 13.480 110.200 13.630 118.400 ;
        RECT 14.080 110.200 14.230 118.400 ;
        RECT 5.930 109.800 14.230 110.200 ;
        RECT 5.930 109.500 6.330 109.800 ;
        RECT 5.930 109.350 9.880 109.500 ;
        RECT 5.930 108.900 6.330 109.350 ;
        RECT 5.930 108.750 9.880 108.900 ;
        RECT 5.930 108.300 6.330 108.750 ;
        RECT 5.930 108.150 9.880 108.300 ;
        RECT 5.930 107.700 6.330 108.150 ;
        RECT 5.930 107.550 9.880 107.700 ;
        RECT 5.930 107.100 6.330 107.550 ;
        RECT 5.930 106.950 9.880 107.100 ;
        RECT 2.315 104.455 4.315 106.750 ;
        RECT 5.930 106.500 6.330 106.950 ;
        RECT 5.930 106.350 9.880 106.500 ;
        RECT 5.930 105.900 6.330 106.350 ;
        RECT 5.930 105.750 9.880 105.900 ;
        RECT 5.930 105.300 6.330 105.750 ;
        RECT 5.930 105.150 9.880 105.300 ;
        RECT 5.930 104.700 6.330 105.150 ;
        RECT 5.930 104.550 9.880 104.700 ;
        RECT 5.930 104.400 6.330 104.550 ;
        RECT 4.730 104.100 6.330 104.400 ;
        RECT 4.730 103.950 9.880 104.100 ;
        RECT 4.730 103.500 6.330 103.950 ;
        RECT 2.315 102.195 4.320 103.470 ;
        RECT 4.730 103.350 9.880 103.500 ;
        RECT 4.730 102.900 6.330 103.350 ;
        RECT 4.730 102.750 9.880 102.900 ;
        RECT 4.730 102.300 6.330 102.750 ;
        RECT 4.730 102.150 9.880 102.300 ;
        RECT 4.730 101.200 5.930 102.150 ;
        RECT 10.480 101.600 10.630 109.800 ;
        RECT 11.080 101.600 11.230 109.800 ;
        RECT 11.680 101.600 11.830 109.800 ;
        RECT 12.280 101.600 12.430 109.800 ;
        RECT 12.880 101.600 13.030 109.800 ;
        RECT 13.480 101.600 13.630 109.800 ;
        RECT 14.080 101.600 14.230 109.800 ;
        RECT 15.230 110.200 15.380 118.400 ;
        RECT 15.830 110.200 15.980 118.400 ;
        RECT 16.430 110.200 16.580 118.400 ;
        RECT 17.030 110.200 17.180 118.400 ;
        RECT 17.630 110.200 17.780 118.400 ;
        RECT 18.230 110.200 18.380 118.400 ;
        RECT 18.830 110.200 18.980 118.400 ;
        RECT 23.530 117.850 25.940 118.800 ;
        RECT 19.580 117.700 29.880 117.850 ;
        RECT 23.130 117.250 26.330 117.700 ;
        RECT 19.580 117.100 29.880 117.250 ;
        RECT 23.130 116.650 26.330 117.100 ;
        RECT 19.580 116.500 29.880 116.650 ;
        RECT 23.130 116.050 26.330 116.500 ;
        RECT 19.580 115.900 29.880 116.050 ;
        RECT 23.130 115.600 26.330 115.900 ;
        RECT 23.130 115.450 23.530 115.600 ;
        RECT 19.580 115.300 23.530 115.450 ;
        RECT 23.130 114.850 23.530 115.300 ;
        RECT 19.580 114.700 23.530 114.850 ;
        RECT 23.130 114.250 23.530 114.700 ;
        RECT 19.580 114.100 23.530 114.250 ;
        RECT 23.130 113.650 23.530 114.100 ;
        RECT 19.580 113.500 23.530 113.650 ;
        RECT 23.130 113.050 23.530 113.500 ;
        RECT 19.580 112.900 23.530 113.050 ;
        RECT 23.130 112.450 23.530 112.900 ;
        RECT 19.580 112.300 23.530 112.450 ;
        RECT 23.130 111.850 23.530 112.300 ;
        RECT 19.580 111.700 23.530 111.850 ;
        RECT 23.130 111.250 23.530 111.700 ;
        RECT 19.580 111.100 23.530 111.250 ;
        RECT 23.130 110.650 23.530 111.100 ;
        RECT 19.580 110.500 23.530 110.650 ;
        RECT 23.130 110.200 23.530 110.500 ;
        RECT 15.230 109.800 23.530 110.200 ;
        RECT 15.230 101.600 15.380 109.800 ;
        RECT 15.830 101.600 15.980 109.800 ;
        RECT 16.430 101.600 16.580 109.800 ;
        RECT 17.030 101.600 17.180 109.800 ;
        RECT 17.630 101.600 17.780 109.800 ;
        RECT 18.230 101.600 18.380 109.800 ;
        RECT 18.830 101.600 18.980 109.800 ;
        RECT 23.130 109.500 23.530 109.800 ;
        RECT 19.580 109.350 23.530 109.500 ;
        RECT 23.130 108.900 23.530 109.350 ;
        RECT 19.580 108.750 23.530 108.900 ;
        RECT 23.130 108.300 23.530 108.750 ;
        RECT 19.580 108.150 23.530 108.300 ;
        RECT 23.130 107.700 23.530 108.150 ;
        RECT 19.580 107.550 23.530 107.700 ;
        RECT 23.130 107.100 23.530 107.550 ;
        RECT 19.580 106.950 23.530 107.100 ;
        RECT 23.130 106.500 23.530 106.950 ;
        RECT 19.580 106.350 23.530 106.500 ;
        RECT 23.130 105.900 23.530 106.350 ;
        RECT 19.580 105.750 23.530 105.900 ;
        RECT 23.130 105.300 23.530 105.750 ;
        RECT 19.580 105.150 23.530 105.300 ;
        RECT 23.130 104.700 23.530 105.150 ;
        RECT 19.580 104.550 23.530 104.700 ;
        RECT 23.130 104.400 23.530 104.550 ;
        RECT 25.930 115.450 26.330 115.600 ;
        RECT 25.930 115.300 29.880 115.450 ;
        RECT 25.930 114.850 26.330 115.300 ;
        RECT 25.930 114.700 29.880 114.850 ;
        RECT 25.930 114.250 26.330 114.700 ;
        RECT 25.930 114.100 29.880 114.250 ;
        RECT 25.930 113.650 26.330 114.100 ;
        RECT 25.930 113.500 29.880 113.650 ;
        RECT 25.930 113.050 26.330 113.500 ;
        RECT 25.930 112.900 29.880 113.050 ;
        RECT 25.930 112.450 26.330 112.900 ;
        RECT 25.930 112.300 29.880 112.450 ;
        RECT 25.930 111.850 26.330 112.300 ;
        RECT 25.930 111.700 29.880 111.850 ;
        RECT 25.930 111.250 26.330 111.700 ;
        RECT 25.930 111.100 29.880 111.250 ;
        RECT 25.930 110.650 26.330 111.100 ;
        RECT 25.930 110.500 29.880 110.650 ;
        RECT 25.930 110.200 26.330 110.500 ;
        RECT 30.480 110.200 30.630 118.400 ;
        RECT 31.080 110.200 31.230 118.400 ;
        RECT 31.680 110.200 31.830 118.400 ;
        RECT 32.280 110.200 32.430 118.400 ;
        RECT 32.880 110.200 33.030 118.400 ;
        RECT 33.480 110.200 33.630 118.400 ;
        RECT 34.080 110.200 34.230 118.400 ;
        RECT 25.930 109.800 34.230 110.200 ;
        RECT 25.930 109.500 26.330 109.800 ;
        RECT 25.930 109.350 29.880 109.500 ;
        RECT 25.930 108.900 26.330 109.350 ;
        RECT 25.930 108.750 29.880 108.900 ;
        RECT 25.930 108.300 26.330 108.750 ;
        RECT 25.930 108.150 29.880 108.300 ;
        RECT 25.930 107.700 26.330 108.150 ;
        RECT 25.930 107.550 29.880 107.700 ;
        RECT 25.930 107.100 26.330 107.550 ;
        RECT 25.930 106.950 29.880 107.100 ;
        RECT 25.930 106.500 26.330 106.950 ;
        RECT 25.930 106.350 29.880 106.500 ;
        RECT 25.930 105.900 26.330 106.350 ;
        RECT 25.930 105.750 29.880 105.900 ;
        RECT 25.930 105.300 26.330 105.750 ;
        RECT 25.930 105.150 29.880 105.300 ;
        RECT 25.930 104.700 26.330 105.150 ;
        RECT 25.930 104.550 29.880 104.700 ;
        RECT 25.930 104.400 26.330 104.550 ;
        RECT 23.130 104.100 26.330 104.400 ;
        RECT 19.580 103.950 29.880 104.100 ;
        RECT 23.130 103.500 26.330 103.950 ;
        RECT 19.580 103.350 29.880 103.500 ;
        RECT 23.130 102.900 26.330 103.350 ;
        RECT 19.580 102.750 29.880 102.900 ;
        RECT 23.130 102.300 26.330 102.750 ;
        RECT 19.580 102.150 29.880 102.300 ;
        RECT 23.530 101.200 25.930 102.150 ;
        RECT 30.480 101.600 30.630 109.800 ;
        RECT 31.080 101.600 31.230 109.800 ;
        RECT 31.680 101.600 31.830 109.800 ;
        RECT 32.280 101.600 32.430 109.800 ;
        RECT 32.880 101.600 33.030 109.800 ;
        RECT 33.480 101.600 33.630 109.800 ;
        RECT 34.080 101.600 34.230 109.800 ;
        RECT 35.230 110.200 35.380 118.400 ;
        RECT 35.830 110.200 35.980 118.400 ;
        RECT 36.430 110.200 36.580 118.400 ;
        RECT 37.030 110.200 37.180 118.400 ;
        RECT 37.630 110.200 37.780 118.400 ;
        RECT 38.230 110.200 38.380 118.400 ;
        RECT 38.830 110.200 38.980 118.400 ;
        RECT 43.530 117.850 45.940 118.800 ;
        RECT 39.580 117.700 49.880 117.850 ;
        RECT 43.130 117.250 46.330 117.700 ;
        RECT 39.580 117.100 49.880 117.250 ;
        RECT 43.130 116.650 46.330 117.100 ;
        RECT 39.580 116.500 49.880 116.650 ;
        RECT 43.130 116.050 46.330 116.500 ;
        RECT 39.580 115.900 49.880 116.050 ;
        RECT 43.130 115.600 46.330 115.900 ;
        RECT 43.130 115.450 43.530 115.600 ;
        RECT 39.580 115.300 43.530 115.450 ;
        RECT 43.130 114.850 43.530 115.300 ;
        RECT 39.580 114.700 43.530 114.850 ;
        RECT 43.130 114.250 43.530 114.700 ;
        RECT 39.580 114.100 43.530 114.250 ;
        RECT 43.130 113.650 43.530 114.100 ;
        RECT 39.580 113.500 43.530 113.650 ;
        RECT 43.130 113.050 43.530 113.500 ;
        RECT 39.580 112.900 43.530 113.050 ;
        RECT 43.130 112.450 43.530 112.900 ;
        RECT 39.580 112.300 43.530 112.450 ;
        RECT 43.130 111.850 43.530 112.300 ;
        RECT 39.580 111.700 43.530 111.850 ;
        RECT 43.130 111.250 43.530 111.700 ;
        RECT 39.580 111.100 43.530 111.250 ;
        RECT 43.130 110.650 43.530 111.100 ;
        RECT 39.580 110.500 43.530 110.650 ;
        RECT 43.130 110.200 43.530 110.500 ;
        RECT 35.230 109.800 43.530 110.200 ;
        RECT 35.230 101.600 35.380 109.800 ;
        RECT 35.830 101.600 35.980 109.800 ;
        RECT 36.430 101.600 36.580 109.800 ;
        RECT 37.030 101.600 37.180 109.800 ;
        RECT 37.630 101.600 37.780 109.800 ;
        RECT 38.230 101.600 38.380 109.800 ;
        RECT 38.830 101.600 38.980 109.800 ;
        RECT 43.130 109.500 43.530 109.800 ;
        RECT 39.580 109.350 43.530 109.500 ;
        RECT 43.130 108.900 43.530 109.350 ;
        RECT 39.580 108.750 43.530 108.900 ;
        RECT 43.130 108.300 43.530 108.750 ;
        RECT 39.580 108.150 43.530 108.300 ;
        RECT 43.130 107.700 43.530 108.150 ;
        RECT 39.580 107.550 43.530 107.700 ;
        RECT 43.130 107.100 43.530 107.550 ;
        RECT 39.580 106.950 43.530 107.100 ;
        RECT 43.130 106.500 43.530 106.950 ;
        RECT 39.580 106.350 43.530 106.500 ;
        RECT 43.130 105.900 43.530 106.350 ;
        RECT 39.580 105.750 43.530 105.900 ;
        RECT 43.130 105.300 43.530 105.750 ;
        RECT 39.580 105.150 43.530 105.300 ;
        RECT 43.130 104.700 43.530 105.150 ;
        RECT 39.580 104.550 43.530 104.700 ;
        RECT 43.130 104.400 43.530 104.550 ;
        RECT 45.930 115.450 46.330 115.600 ;
        RECT 45.930 115.300 49.880 115.450 ;
        RECT 45.930 114.850 46.330 115.300 ;
        RECT 45.930 114.700 49.880 114.850 ;
        RECT 45.930 114.250 46.330 114.700 ;
        RECT 45.930 114.100 49.880 114.250 ;
        RECT 45.930 113.650 46.330 114.100 ;
        RECT 45.930 113.500 49.880 113.650 ;
        RECT 45.930 113.050 46.330 113.500 ;
        RECT 45.930 112.900 49.880 113.050 ;
        RECT 45.930 112.450 46.330 112.900 ;
        RECT 45.930 112.300 49.880 112.450 ;
        RECT 45.930 111.850 46.330 112.300 ;
        RECT 45.930 111.700 49.880 111.850 ;
        RECT 45.930 111.250 46.330 111.700 ;
        RECT 45.930 111.100 49.880 111.250 ;
        RECT 45.930 110.650 46.330 111.100 ;
        RECT 45.930 110.500 49.880 110.650 ;
        RECT 45.930 110.200 46.330 110.500 ;
        RECT 50.480 110.200 50.630 118.400 ;
        RECT 51.080 110.200 51.230 118.400 ;
        RECT 51.680 110.200 51.830 118.400 ;
        RECT 52.280 110.200 52.430 118.400 ;
        RECT 52.880 110.200 53.030 118.400 ;
        RECT 53.480 110.200 53.630 118.400 ;
        RECT 54.080 110.200 54.230 118.400 ;
        RECT 45.930 109.800 54.230 110.200 ;
        RECT 45.930 109.500 46.330 109.800 ;
        RECT 45.930 109.350 49.880 109.500 ;
        RECT 45.930 108.900 46.330 109.350 ;
        RECT 45.930 108.750 49.880 108.900 ;
        RECT 45.930 108.300 46.330 108.750 ;
        RECT 45.930 108.150 49.880 108.300 ;
        RECT 45.930 107.700 46.330 108.150 ;
        RECT 45.930 107.550 49.880 107.700 ;
        RECT 45.930 107.100 46.330 107.550 ;
        RECT 45.930 106.950 49.880 107.100 ;
        RECT 45.930 106.500 46.330 106.950 ;
        RECT 45.930 106.350 49.880 106.500 ;
        RECT 45.930 105.900 46.330 106.350 ;
        RECT 45.930 105.750 49.880 105.900 ;
        RECT 45.930 105.300 46.330 105.750 ;
        RECT 45.930 105.150 49.880 105.300 ;
        RECT 45.930 104.700 46.330 105.150 ;
        RECT 45.930 104.550 49.880 104.700 ;
        RECT 45.930 104.400 46.330 104.550 ;
        RECT 43.130 104.100 46.330 104.400 ;
        RECT 39.580 103.950 49.880 104.100 ;
        RECT 43.130 103.500 46.330 103.950 ;
        RECT 39.580 103.350 49.880 103.500 ;
        RECT 43.130 102.900 46.330 103.350 ;
        RECT 39.580 102.750 49.880 102.900 ;
        RECT 43.130 102.300 46.330 102.750 ;
        RECT 39.580 102.150 49.880 102.300 ;
        RECT 43.530 101.200 45.930 102.150 ;
        RECT 50.480 101.600 50.630 109.800 ;
        RECT 51.080 101.600 51.230 109.800 ;
        RECT 51.680 101.600 51.830 109.800 ;
        RECT 52.280 101.600 52.430 109.800 ;
        RECT 52.880 101.600 53.030 109.800 ;
        RECT 53.480 101.600 53.630 109.800 ;
        RECT 54.080 101.600 54.230 109.800 ;
        RECT 55.230 110.200 55.380 118.400 ;
        RECT 55.830 110.200 55.980 118.400 ;
        RECT 56.430 110.200 56.580 118.400 ;
        RECT 57.030 110.200 57.180 118.400 ;
        RECT 57.630 110.200 57.780 118.400 ;
        RECT 58.230 110.200 58.380 118.400 ;
        RECT 58.830 110.200 58.980 118.400 ;
        RECT 63.530 117.850 65.940 118.800 ;
        RECT 59.580 117.700 69.880 117.850 ;
        RECT 63.130 117.250 66.330 117.700 ;
        RECT 59.580 117.100 69.880 117.250 ;
        RECT 63.130 116.650 66.330 117.100 ;
        RECT 59.580 116.500 69.880 116.650 ;
        RECT 63.130 116.050 66.330 116.500 ;
        RECT 59.580 115.900 69.880 116.050 ;
        RECT 63.130 115.600 66.330 115.900 ;
        RECT 63.130 115.450 63.530 115.600 ;
        RECT 59.580 115.300 63.530 115.450 ;
        RECT 63.130 114.850 63.530 115.300 ;
        RECT 59.580 114.700 63.530 114.850 ;
        RECT 63.130 114.250 63.530 114.700 ;
        RECT 59.580 114.100 63.530 114.250 ;
        RECT 63.130 113.650 63.530 114.100 ;
        RECT 59.580 113.500 63.530 113.650 ;
        RECT 63.130 113.050 63.530 113.500 ;
        RECT 59.580 112.900 63.530 113.050 ;
        RECT 63.130 112.450 63.530 112.900 ;
        RECT 59.580 112.300 63.530 112.450 ;
        RECT 63.130 111.850 63.530 112.300 ;
        RECT 59.580 111.700 63.530 111.850 ;
        RECT 63.130 111.250 63.530 111.700 ;
        RECT 59.580 111.100 63.530 111.250 ;
        RECT 63.130 110.650 63.530 111.100 ;
        RECT 59.580 110.500 63.530 110.650 ;
        RECT 63.130 110.200 63.530 110.500 ;
        RECT 55.230 109.800 63.530 110.200 ;
        RECT 55.230 101.600 55.380 109.800 ;
        RECT 55.830 101.600 55.980 109.800 ;
        RECT 56.430 101.600 56.580 109.800 ;
        RECT 57.030 101.600 57.180 109.800 ;
        RECT 57.630 101.600 57.780 109.800 ;
        RECT 58.230 101.600 58.380 109.800 ;
        RECT 58.830 101.600 58.980 109.800 ;
        RECT 63.130 109.500 63.530 109.800 ;
        RECT 59.580 109.350 63.530 109.500 ;
        RECT 63.130 108.900 63.530 109.350 ;
        RECT 59.580 108.750 63.530 108.900 ;
        RECT 63.130 108.300 63.530 108.750 ;
        RECT 59.580 108.150 63.530 108.300 ;
        RECT 63.130 107.700 63.530 108.150 ;
        RECT 59.580 107.550 63.530 107.700 ;
        RECT 63.130 107.100 63.530 107.550 ;
        RECT 59.580 106.950 63.530 107.100 ;
        RECT 63.130 106.500 63.530 106.950 ;
        RECT 59.580 106.350 63.530 106.500 ;
        RECT 63.130 105.900 63.530 106.350 ;
        RECT 59.580 105.750 63.530 105.900 ;
        RECT 63.130 105.300 63.530 105.750 ;
        RECT 59.580 105.150 63.530 105.300 ;
        RECT 63.130 104.700 63.530 105.150 ;
        RECT 59.580 104.550 63.530 104.700 ;
        RECT 63.130 104.400 63.530 104.550 ;
        RECT 65.930 115.450 66.330 115.600 ;
        RECT 65.930 115.300 69.880 115.450 ;
        RECT 65.930 114.850 66.330 115.300 ;
        RECT 65.930 114.700 69.880 114.850 ;
        RECT 65.930 114.250 66.330 114.700 ;
        RECT 65.930 114.100 69.880 114.250 ;
        RECT 65.930 113.650 66.330 114.100 ;
        RECT 65.930 113.500 69.880 113.650 ;
        RECT 65.930 113.050 66.330 113.500 ;
        RECT 65.930 112.900 69.880 113.050 ;
        RECT 65.930 112.450 66.330 112.900 ;
        RECT 65.930 112.300 69.880 112.450 ;
        RECT 65.930 111.850 66.330 112.300 ;
        RECT 65.930 111.700 69.880 111.850 ;
        RECT 65.930 111.250 66.330 111.700 ;
        RECT 65.930 111.100 69.880 111.250 ;
        RECT 65.930 110.650 66.330 111.100 ;
        RECT 65.930 110.500 69.880 110.650 ;
        RECT 65.930 110.200 66.330 110.500 ;
        RECT 70.480 110.200 70.630 118.400 ;
        RECT 71.080 110.200 71.230 118.400 ;
        RECT 71.680 110.200 71.830 118.400 ;
        RECT 72.280 110.200 72.430 118.400 ;
        RECT 72.880 110.200 73.030 118.400 ;
        RECT 73.480 110.200 73.630 118.400 ;
        RECT 74.080 110.200 74.230 118.400 ;
        RECT 65.930 109.800 74.230 110.200 ;
        RECT 65.930 109.500 66.330 109.800 ;
        RECT 65.930 109.350 69.880 109.500 ;
        RECT 65.930 108.900 66.330 109.350 ;
        RECT 65.930 108.750 69.880 108.900 ;
        RECT 65.930 108.300 66.330 108.750 ;
        RECT 65.930 108.150 69.880 108.300 ;
        RECT 65.930 107.700 66.330 108.150 ;
        RECT 65.930 107.550 69.880 107.700 ;
        RECT 65.930 107.100 66.330 107.550 ;
        RECT 65.930 106.950 69.880 107.100 ;
        RECT 65.930 106.500 66.330 106.950 ;
        RECT 65.930 106.350 69.880 106.500 ;
        RECT 65.930 105.900 66.330 106.350 ;
        RECT 65.930 105.750 69.880 105.900 ;
        RECT 65.930 105.300 66.330 105.750 ;
        RECT 65.930 105.150 69.880 105.300 ;
        RECT 65.930 104.700 66.330 105.150 ;
        RECT 65.930 104.550 69.880 104.700 ;
        RECT 65.930 104.400 66.330 104.550 ;
        RECT 63.130 104.100 66.330 104.400 ;
        RECT 59.580 103.950 69.880 104.100 ;
        RECT 63.130 103.500 66.330 103.950 ;
        RECT 59.580 103.350 69.880 103.500 ;
        RECT 63.130 102.900 66.330 103.350 ;
        RECT 59.580 102.750 69.880 102.900 ;
        RECT 63.130 102.300 66.330 102.750 ;
        RECT 59.580 102.150 69.880 102.300 ;
        RECT 63.530 101.200 65.930 102.150 ;
        RECT 70.480 101.600 70.630 109.800 ;
        RECT 71.080 101.600 71.230 109.800 ;
        RECT 71.680 101.600 71.830 109.800 ;
        RECT 72.280 101.600 72.430 109.800 ;
        RECT 72.880 101.600 73.030 109.800 ;
        RECT 73.480 101.600 73.630 109.800 ;
        RECT 74.080 101.600 74.230 109.800 ;
        RECT 75.230 110.200 75.380 118.400 ;
        RECT 75.830 110.200 75.980 118.400 ;
        RECT 76.430 110.200 76.580 118.400 ;
        RECT 77.030 110.200 77.180 118.400 ;
        RECT 77.630 110.200 77.780 118.400 ;
        RECT 78.230 110.200 78.380 118.400 ;
        RECT 78.830 110.200 78.980 118.400 ;
        RECT 83.530 117.850 85.940 118.800 ;
        RECT 79.580 117.700 89.880 117.850 ;
        RECT 83.130 117.250 86.330 117.700 ;
        RECT 79.580 117.100 89.880 117.250 ;
        RECT 83.130 116.650 86.330 117.100 ;
        RECT 79.580 116.500 89.880 116.650 ;
        RECT 83.130 116.050 86.330 116.500 ;
        RECT 79.580 115.900 89.880 116.050 ;
        RECT 83.130 115.600 86.330 115.900 ;
        RECT 83.130 115.450 83.530 115.600 ;
        RECT 79.580 115.300 83.530 115.450 ;
        RECT 83.130 114.850 83.530 115.300 ;
        RECT 79.580 114.700 83.530 114.850 ;
        RECT 83.130 114.250 83.530 114.700 ;
        RECT 79.580 114.100 83.530 114.250 ;
        RECT 83.130 113.650 83.530 114.100 ;
        RECT 79.580 113.500 83.530 113.650 ;
        RECT 83.130 113.050 83.530 113.500 ;
        RECT 79.580 112.900 83.530 113.050 ;
        RECT 83.130 112.450 83.530 112.900 ;
        RECT 79.580 112.300 83.530 112.450 ;
        RECT 83.130 111.850 83.530 112.300 ;
        RECT 79.580 111.700 83.530 111.850 ;
        RECT 83.130 111.250 83.530 111.700 ;
        RECT 79.580 111.100 83.530 111.250 ;
        RECT 83.130 110.650 83.530 111.100 ;
        RECT 79.580 110.500 83.530 110.650 ;
        RECT 83.130 110.200 83.530 110.500 ;
        RECT 75.230 109.800 83.530 110.200 ;
        RECT 75.230 101.600 75.380 109.800 ;
        RECT 75.830 101.600 75.980 109.800 ;
        RECT 76.430 101.600 76.580 109.800 ;
        RECT 77.030 101.600 77.180 109.800 ;
        RECT 77.630 101.600 77.780 109.800 ;
        RECT 78.230 101.600 78.380 109.800 ;
        RECT 78.830 101.600 78.980 109.800 ;
        RECT 83.130 109.500 83.530 109.800 ;
        RECT 79.580 109.350 83.530 109.500 ;
        RECT 83.130 108.900 83.530 109.350 ;
        RECT 79.580 108.750 83.530 108.900 ;
        RECT 83.130 108.300 83.530 108.750 ;
        RECT 79.580 108.150 83.530 108.300 ;
        RECT 83.130 107.700 83.530 108.150 ;
        RECT 79.580 107.550 83.530 107.700 ;
        RECT 83.130 107.100 83.530 107.550 ;
        RECT 79.580 106.950 83.530 107.100 ;
        RECT 83.130 106.500 83.530 106.950 ;
        RECT 79.580 106.350 83.530 106.500 ;
        RECT 83.130 105.900 83.530 106.350 ;
        RECT 79.580 105.750 83.530 105.900 ;
        RECT 83.130 105.300 83.530 105.750 ;
        RECT 79.580 105.150 83.530 105.300 ;
        RECT 83.130 104.700 83.530 105.150 ;
        RECT 79.580 104.550 83.530 104.700 ;
        RECT 83.130 104.400 83.530 104.550 ;
        RECT 85.930 115.450 86.330 115.600 ;
        RECT 85.930 115.300 89.880 115.450 ;
        RECT 85.930 114.850 86.330 115.300 ;
        RECT 85.930 114.700 89.880 114.850 ;
        RECT 85.930 114.250 86.330 114.700 ;
        RECT 85.930 114.100 89.880 114.250 ;
        RECT 85.930 113.650 86.330 114.100 ;
        RECT 85.930 113.500 89.880 113.650 ;
        RECT 85.930 113.050 86.330 113.500 ;
        RECT 85.930 112.900 89.880 113.050 ;
        RECT 85.930 112.450 86.330 112.900 ;
        RECT 85.930 112.300 89.880 112.450 ;
        RECT 85.930 111.850 86.330 112.300 ;
        RECT 85.930 111.700 89.880 111.850 ;
        RECT 85.930 111.250 86.330 111.700 ;
        RECT 85.930 111.100 89.880 111.250 ;
        RECT 85.930 110.650 86.330 111.100 ;
        RECT 85.930 110.500 89.880 110.650 ;
        RECT 85.930 110.200 86.330 110.500 ;
        RECT 90.480 110.200 90.630 118.400 ;
        RECT 91.080 110.200 91.230 118.400 ;
        RECT 91.680 110.200 91.830 118.400 ;
        RECT 92.280 110.200 92.430 118.400 ;
        RECT 92.880 110.200 93.030 118.400 ;
        RECT 93.480 110.200 93.630 118.400 ;
        RECT 94.080 110.200 94.230 118.400 ;
        RECT 85.930 109.800 94.230 110.200 ;
        RECT 85.930 109.500 86.330 109.800 ;
        RECT 85.930 109.350 89.880 109.500 ;
        RECT 85.930 108.900 86.330 109.350 ;
        RECT 85.930 108.750 89.880 108.900 ;
        RECT 85.930 108.300 86.330 108.750 ;
        RECT 85.930 108.150 89.880 108.300 ;
        RECT 85.930 107.700 86.330 108.150 ;
        RECT 85.930 107.550 89.880 107.700 ;
        RECT 85.930 107.100 86.330 107.550 ;
        RECT 85.930 106.950 89.880 107.100 ;
        RECT 85.930 106.500 86.330 106.950 ;
        RECT 85.930 106.350 89.880 106.500 ;
        RECT 85.930 105.900 86.330 106.350 ;
        RECT 85.930 105.750 89.880 105.900 ;
        RECT 85.930 105.300 86.330 105.750 ;
        RECT 85.930 105.150 89.880 105.300 ;
        RECT 85.930 104.700 86.330 105.150 ;
        RECT 85.930 104.550 89.880 104.700 ;
        RECT 85.930 104.400 86.330 104.550 ;
        RECT 83.130 104.100 86.330 104.400 ;
        RECT 79.580 103.950 89.880 104.100 ;
        RECT 83.130 103.500 86.330 103.950 ;
        RECT 79.580 103.350 89.880 103.500 ;
        RECT 83.130 102.900 86.330 103.350 ;
        RECT 79.580 102.750 89.880 102.900 ;
        RECT 83.130 102.300 86.330 102.750 ;
        RECT 79.580 102.150 89.880 102.300 ;
        RECT 83.530 101.200 85.930 102.150 ;
        RECT 90.480 101.600 90.630 109.800 ;
        RECT 91.080 101.600 91.230 109.800 ;
        RECT 91.680 101.600 91.830 109.800 ;
        RECT 92.280 101.600 92.430 109.800 ;
        RECT 92.880 101.600 93.030 109.800 ;
        RECT 93.480 101.600 93.630 109.800 ;
        RECT 94.080 101.600 94.230 109.800 ;
        RECT 95.230 110.200 95.380 118.400 ;
        RECT 95.830 110.200 95.980 118.400 ;
        RECT 96.430 110.200 96.580 118.400 ;
        RECT 97.030 110.200 97.180 118.400 ;
        RECT 97.630 110.200 97.780 118.400 ;
        RECT 98.230 110.200 98.380 118.400 ;
        RECT 98.830 110.200 98.980 118.400 ;
        RECT 103.530 117.850 104.730 118.800 ;
        RECT 99.580 117.700 104.730 117.850 ;
        RECT 103.130 117.250 104.730 117.700 ;
        RECT 99.580 117.100 104.730 117.250 ;
        RECT 103.130 116.650 104.730 117.100 ;
        RECT 99.580 116.500 104.730 116.650 ;
        RECT 103.130 116.050 104.730 116.500 ;
        RECT 99.580 115.900 104.730 116.050 ;
        RECT 105.140 115.970 107.140 117.245 ;
        RECT 103.130 115.600 104.730 115.900 ;
        RECT 103.130 115.450 103.530 115.600 ;
        RECT 99.580 115.300 103.530 115.450 ;
        RECT 103.130 114.850 103.530 115.300 ;
        RECT 99.580 114.700 103.530 114.850 ;
        RECT 103.130 114.250 103.530 114.700 ;
        RECT 99.580 114.100 103.530 114.250 ;
        RECT 103.130 113.650 103.530 114.100 ;
        RECT 99.580 113.500 103.530 113.650 ;
        RECT 103.130 113.050 103.530 113.500 ;
        RECT 99.580 112.900 103.530 113.050 ;
        RECT 103.130 112.450 103.530 112.900 ;
        RECT 99.580 112.300 103.530 112.450 ;
        RECT 103.130 111.850 103.530 112.300 ;
        RECT 99.580 111.700 103.530 111.850 ;
        RECT 103.130 111.250 103.530 111.700 ;
        RECT 99.580 111.100 103.530 111.250 ;
        RECT 103.130 110.650 103.530 111.100 ;
        RECT 99.580 110.500 103.530 110.650 ;
        RECT 103.130 110.200 103.530 110.500 ;
        RECT 95.230 109.800 103.530 110.200 ;
        RECT 95.230 101.600 95.380 109.800 ;
        RECT 95.830 101.600 95.980 109.800 ;
        RECT 96.430 101.600 96.580 109.800 ;
        RECT 97.030 101.600 97.180 109.800 ;
        RECT 97.630 101.600 97.780 109.800 ;
        RECT 98.230 101.600 98.380 109.800 ;
        RECT 98.830 101.600 98.980 109.800 ;
        RECT 103.130 109.500 103.530 109.800 ;
        RECT 99.580 109.350 103.530 109.500 ;
        RECT 103.130 108.900 103.530 109.350 ;
        RECT 99.580 108.750 103.530 108.900 ;
        RECT 103.130 108.300 103.530 108.750 ;
        RECT 99.580 108.150 103.530 108.300 ;
        RECT 103.130 107.700 103.530 108.150 ;
        RECT 99.580 107.550 103.530 107.700 ;
        RECT 103.130 107.100 103.530 107.550 ;
        RECT 99.580 106.950 103.530 107.100 ;
        RECT 103.130 106.500 103.530 106.950 ;
        RECT 99.580 106.350 103.530 106.500 ;
        RECT 103.130 105.900 103.530 106.350 ;
        RECT 99.580 105.750 103.530 105.900 ;
        RECT 103.130 105.300 103.530 105.750 ;
        RECT 99.580 105.150 103.530 105.300 ;
        RECT 103.130 104.700 103.530 105.150 ;
        RECT 99.580 104.550 103.530 104.700 ;
        RECT 103.130 104.400 103.530 104.550 ;
        RECT 103.130 104.100 104.730 104.400 ;
        RECT 99.580 103.950 104.730 104.100 ;
        RECT 103.130 103.500 104.730 103.950 ;
        RECT 99.580 103.350 104.730 103.500 ;
        RECT 103.130 102.900 104.730 103.350 ;
        RECT 99.580 102.750 104.730 102.900 ;
        RECT 103.130 102.300 104.730 102.750 ;
        RECT 99.580 102.150 104.730 102.300 ;
        RECT 103.530 101.200 104.730 102.150 ;
        RECT 105.135 101.765 107.135 103.040 ;
        RECT 4.730 98.800 9.130 101.200 ;
        RECT 20.330 98.800 29.130 101.200 ;
        RECT 40.330 98.800 49.130 101.200 ;
        RECT 60.330 98.800 69.130 101.200 ;
        RECT 80.330 98.800 89.130 101.200 ;
        RECT 100.330 98.800 104.730 101.200 ;
        RECT 2.315 96.690 4.320 97.965 ;
        RECT 4.730 97.850 5.940 98.800 ;
        RECT 4.730 97.700 9.880 97.850 ;
        RECT 4.730 97.250 6.330 97.700 ;
        RECT 4.730 97.100 9.880 97.250 ;
        RECT 4.730 96.650 6.330 97.100 ;
        RECT 4.730 96.500 9.880 96.650 ;
        RECT 4.730 96.050 6.330 96.500 ;
        RECT 4.730 95.900 9.880 96.050 ;
        RECT 4.730 95.600 6.330 95.900 ;
        RECT 2.315 93.250 4.315 95.545 ;
        RECT 5.930 95.450 6.330 95.600 ;
        RECT 5.930 95.300 9.880 95.450 ;
        RECT 5.930 94.850 6.330 95.300 ;
        RECT 5.930 94.700 9.880 94.850 ;
        RECT 5.930 94.250 6.330 94.700 ;
        RECT 5.930 94.100 9.880 94.250 ;
        RECT 5.930 93.650 6.330 94.100 ;
        RECT 5.930 93.500 9.880 93.650 ;
        RECT 5.930 93.050 6.330 93.500 ;
        RECT 5.930 92.900 9.880 93.050 ;
        RECT 5.930 92.450 6.330 92.900 ;
        RECT 5.930 92.300 9.880 92.450 ;
        RECT 5.930 91.850 6.330 92.300 ;
        RECT 5.930 91.700 9.880 91.850 ;
        RECT 5.930 91.250 6.330 91.700 ;
        RECT 5.930 91.100 9.880 91.250 ;
        RECT 5.930 90.650 6.330 91.100 ;
        RECT 5.930 90.500 9.880 90.650 ;
        RECT 5.930 90.200 6.330 90.500 ;
        RECT 10.480 90.200 10.630 98.400 ;
        RECT 11.080 90.200 11.230 98.400 ;
        RECT 11.680 90.200 11.830 98.400 ;
        RECT 12.280 90.200 12.430 98.400 ;
        RECT 12.880 90.200 13.030 98.400 ;
        RECT 13.480 90.200 13.630 98.400 ;
        RECT 14.080 90.200 14.230 98.400 ;
        RECT 5.930 89.800 14.230 90.200 ;
        RECT 5.930 89.500 6.330 89.800 ;
        RECT 5.930 89.350 9.880 89.500 ;
        RECT 5.930 88.900 6.330 89.350 ;
        RECT 5.930 88.750 9.880 88.900 ;
        RECT 5.930 88.300 6.330 88.750 ;
        RECT 5.930 88.150 9.880 88.300 ;
        RECT 5.930 87.700 6.330 88.150 ;
        RECT 5.930 87.550 9.880 87.700 ;
        RECT 5.930 87.100 6.330 87.550 ;
        RECT 5.930 86.950 9.880 87.100 ;
        RECT 2.315 84.450 4.315 86.745 ;
        RECT 5.930 86.500 6.330 86.950 ;
        RECT 5.930 86.350 9.880 86.500 ;
        RECT 5.930 85.900 6.330 86.350 ;
        RECT 5.930 85.750 9.880 85.900 ;
        RECT 5.930 85.300 6.330 85.750 ;
        RECT 5.930 85.150 9.880 85.300 ;
        RECT 5.930 84.700 6.330 85.150 ;
        RECT 5.930 84.550 9.880 84.700 ;
        RECT 5.930 84.400 6.330 84.550 ;
        RECT 4.730 84.100 6.330 84.400 ;
        RECT 4.730 83.950 9.880 84.100 ;
        RECT 2.315 82.360 4.325 83.635 ;
        RECT 4.730 83.500 6.330 83.950 ;
        RECT 4.730 83.350 9.880 83.500 ;
        RECT 4.730 82.900 6.330 83.350 ;
        RECT 4.730 82.750 9.880 82.900 ;
        RECT 4.730 82.300 6.330 82.750 ;
        RECT 4.730 82.150 9.880 82.300 ;
        RECT 4.730 81.200 5.930 82.150 ;
        RECT 10.480 81.600 10.630 89.800 ;
        RECT 11.080 81.600 11.230 89.800 ;
        RECT 11.680 81.600 11.830 89.800 ;
        RECT 12.280 81.600 12.430 89.800 ;
        RECT 12.880 81.600 13.030 89.800 ;
        RECT 13.480 81.600 13.630 89.800 ;
        RECT 14.080 81.600 14.230 89.800 ;
        RECT 15.230 90.200 15.380 98.400 ;
        RECT 15.830 90.200 15.980 98.400 ;
        RECT 16.430 90.200 16.580 98.400 ;
        RECT 17.030 90.200 17.180 98.400 ;
        RECT 17.630 90.200 17.780 98.400 ;
        RECT 18.230 90.200 18.380 98.400 ;
        RECT 18.830 90.200 18.980 98.400 ;
        RECT 23.530 97.850 25.940 98.800 ;
        RECT 19.580 97.700 29.880 97.850 ;
        RECT 23.130 97.250 26.330 97.700 ;
        RECT 19.580 97.100 29.880 97.250 ;
        RECT 23.130 96.650 26.330 97.100 ;
        RECT 19.580 96.500 29.880 96.650 ;
        RECT 23.130 96.050 26.330 96.500 ;
        RECT 19.580 95.900 29.880 96.050 ;
        RECT 23.130 95.600 26.330 95.900 ;
        RECT 23.130 95.450 23.530 95.600 ;
        RECT 19.580 95.300 23.530 95.450 ;
        RECT 23.130 94.850 23.530 95.300 ;
        RECT 19.580 94.700 23.530 94.850 ;
        RECT 23.130 94.250 23.530 94.700 ;
        RECT 19.580 94.100 23.530 94.250 ;
        RECT 23.130 93.650 23.530 94.100 ;
        RECT 19.580 93.500 23.530 93.650 ;
        RECT 23.130 93.050 23.530 93.500 ;
        RECT 19.580 92.900 23.530 93.050 ;
        RECT 23.130 92.450 23.530 92.900 ;
        RECT 19.580 92.300 23.530 92.450 ;
        RECT 23.130 91.850 23.530 92.300 ;
        RECT 19.580 91.700 23.530 91.850 ;
        RECT 23.130 91.250 23.530 91.700 ;
        RECT 19.580 91.100 23.530 91.250 ;
        RECT 23.130 90.650 23.530 91.100 ;
        RECT 19.580 90.500 23.530 90.650 ;
        RECT 23.130 90.200 23.530 90.500 ;
        RECT 15.230 89.800 23.530 90.200 ;
        RECT 15.230 81.600 15.380 89.800 ;
        RECT 15.830 81.600 15.980 89.800 ;
        RECT 16.430 81.600 16.580 89.800 ;
        RECT 17.030 81.600 17.180 89.800 ;
        RECT 17.630 81.600 17.780 89.800 ;
        RECT 18.230 81.600 18.380 89.800 ;
        RECT 18.830 81.600 18.980 89.800 ;
        RECT 23.130 89.500 23.530 89.800 ;
        RECT 19.580 89.350 23.530 89.500 ;
        RECT 23.130 88.900 23.530 89.350 ;
        RECT 19.580 88.750 23.530 88.900 ;
        RECT 23.130 88.300 23.530 88.750 ;
        RECT 19.580 88.150 23.530 88.300 ;
        RECT 23.130 87.700 23.530 88.150 ;
        RECT 19.580 87.550 23.530 87.700 ;
        RECT 23.130 87.100 23.530 87.550 ;
        RECT 19.580 86.950 23.530 87.100 ;
        RECT 23.130 86.500 23.530 86.950 ;
        RECT 19.580 86.350 23.530 86.500 ;
        RECT 23.130 85.900 23.530 86.350 ;
        RECT 19.580 85.750 23.530 85.900 ;
        RECT 23.130 85.300 23.530 85.750 ;
        RECT 19.580 85.150 23.530 85.300 ;
        RECT 23.130 84.700 23.530 85.150 ;
        RECT 19.580 84.550 23.530 84.700 ;
        RECT 23.130 84.400 23.530 84.550 ;
        RECT 25.930 95.450 26.330 95.600 ;
        RECT 25.930 95.300 29.880 95.450 ;
        RECT 25.930 94.850 26.330 95.300 ;
        RECT 25.930 94.700 29.880 94.850 ;
        RECT 25.930 94.250 26.330 94.700 ;
        RECT 25.930 94.100 29.880 94.250 ;
        RECT 25.930 93.650 26.330 94.100 ;
        RECT 25.930 93.500 29.880 93.650 ;
        RECT 25.930 93.050 26.330 93.500 ;
        RECT 25.930 92.900 29.880 93.050 ;
        RECT 25.930 92.450 26.330 92.900 ;
        RECT 25.930 92.300 29.880 92.450 ;
        RECT 25.930 91.850 26.330 92.300 ;
        RECT 25.930 91.700 29.880 91.850 ;
        RECT 25.930 91.250 26.330 91.700 ;
        RECT 25.930 91.100 29.880 91.250 ;
        RECT 25.930 90.650 26.330 91.100 ;
        RECT 25.930 90.500 29.880 90.650 ;
        RECT 25.930 90.200 26.330 90.500 ;
        RECT 30.480 90.200 30.630 98.400 ;
        RECT 31.080 90.200 31.230 98.400 ;
        RECT 31.680 90.200 31.830 98.400 ;
        RECT 32.280 90.200 32.430 98.400 ;
        RECT 32.880 90.200 33.030 98.400 ;
        RECT 33.480 90.200 33.630 98.400 ;
        RECT 34.080 90.200 34.230 98.400 ;
        RECT 25.930 89.800 34.230 90.200 ;
        RECT 25.930 89.500 26.330 89.800 ;
        RECT 25.930 89.350 29.880 89.500 ;
        RECT 25.930 88.900 26.330 89.350 ;
        RECT 25.930 88.750 29.880 88.900 ;
        RECT 25.930 88.300 26.330 88.750 ;
        RECT 25.930 88.150 29.880 88.300 ;
        RECT 25.930 87.700 26.330 88.150 ;
        RECT 25.930 87.550 29.880 87.700 ;
        RECT 25.930 87.100 26.330 87.550 ;
        RECT 25.930 86.950 29.880 87.100 ;
        RECT 25.930 86.500 26.330 86.950 ;
        RECT 25.930 86.350 29.880 86.500 ;
        RECT 25.930 85.900 26.330 86.350 ;
        RECT 25.930 85.750 29.880 85.900 ;
        RECT 25.930 85.300 26.330 85.750 ;
        RECT 25.930 85.150 29.880 85.300 ;
        RECT 25.930 84.700 26.330 85.150 ;
        RECT 25.930 84.550 29.880 84.700 ;
        RECT 25.930 84.400 26.330 84.550 ;
        RECT 23.130 84.100 26.330 84.400 ;
        RECT 19.580 83.950 29.880 84.100 ;
        RECT 23.130 83.500 26.330 83.950 ;
        RECT 19.580 83.350 29.880 83.500 ;
        RECT 23.130 82.900 26.330 83.350 ;
        RECT 19.580 82.750 29.880 82.900 ;
        RECT 23.130 82.300 26.330 82.750 ;
        RECT 19.580 82.150 29.880 82.300 ;
        RECT 23.530 81.200 25.930 82.150 ;
        RECT 30.480 81.600 30.630 89.800 ;
        RECT 31.080 81.600 31.230 89.800 ;
        RECT 31.680 81.600 31.830 89.800 ;
        RECT 32.280 81.600 32.430 89.800 ;
        RECT 32.880 81.600 33.030 89.800 ;
        RECT 33.480 81.600 33.630 89.800 ;
        RECT 34.080 81.600 34.230 89.800 ;
        RECT 35.230 90.200 35.380 98.400 ;
        RECT 35.830 90.200 35.980 98.400 ;
        RECT 36.430 90.200 36.580 98.400 ;
        RECT 37.030 90.200 37.180 98.400 ;
        RECT 37.630 90.200 37.780 98.400 ;
        RECT 38.230 90.200 38.380 98.400 ;
        RECT 38.830 90.200 38.980 98.400 ;
        RECT 43.530 97.850 45.940 98.800 ;
        RECT 39.580 97.700 49.880 97.850 ;
        RECT 43.130 97.250 46.330 97.700 ;
        RECT 39.580 97.100 49.880 97.250 ;
        RECT 43.130 96.650 46.330 97.100 ;
        RECT 39.580 96.500 49.880 96.650 ;
        RECT 43.130 96.050 46.330 96.500 ;
        RECT 39.580 95.900 49.880 96.050 ;
        RECT 43.130 95.600 46.330 95.900 ;
        RECT 43.130 95.450 43.530 95.600 ;
        RECT 39.580 95.300 43.530 95.450 ;
        RECT 43.130 94.850 43.530 95.300 ;
        RECT 39.580 94.700 43.530 94.850 ;
        RECT 43.130 94.250 43.530 94.700 ;
        RECT 39.580 94.100 43.530 94.250 ;
        RECT 43.130 93.650 43.530 94.100 ;
        RECT 39.580 93.500 43.530 93.650 ;
        RECT 43.130 93.050 43.530 93.500 ;
        RECT 39.580 92.900 43.530 93.050 ;
        RECT 43.130 92.450 43.530 92.900 ;
        RECT 39.580 92.300 43.530 92.450 ;
        RECT 43.130 91.850 43.530 92.300 ;
        RECT 39.580 91.700 43.530 91.850 ;
        RECT 43.130 91.250 43.530 91.700 ;
        RECT 39.580 91.100 43.530 91.250 ;
        RECT 43.130 90.650 43.530 91.100 ;
        RECT 39.580 90.500 43.530 90.650 ;
        RECT 43.130 90.200 43.530 90.500 ;
        RECT 35.230 89.800 43.530 90.200 ;
        RECT 35.230 81.600 35.380 89.800 ;
        RECT 35.830 81.600 35.980 89.800 ;
        RECT 36.430 81.600 36.580 89.800 ;
        RECT 37.030 81.600 37.180 89.800 ;
        RECT 37.630 81.600 37.780 89.800 ;
        RECT 38.230 81.600 38.380 89.800 ;
        RECT 38.830 81.600 38.980 89.800 ;
        RECT 43.130 89.500 43.530 89.800 ;
        RECT 39.580 89.350 43.530 89.500 ;
        RECT 43.130 88.900 43.530 89.350 ;
        RECT 39.580 88.750 43.530 88.900 ;
        RECT 43.130 88.300 43.530 88.750 ;
        RECT 39.580 88.150 43.530 88.300 ;
        RECT 43.130 87.700 43.530 88.150 ;
        RECT 39.580 87.550 43.530 87.700 ;
        RECT 43.130 87.100 43.530 87.550 ;
        RECT 39.580 86.950 43.530 87.100 ;
        RECT 43.130 86.500 43.530 86.950 ;
        RECT 39.580 86.350 43.530 86.500 ;
        RECT 43.130 85.900 43.530 86.350 ;
        RECT 39.580 85.750 43.530 85.900 ;
        RECT 43.130 85.300 43.530 85.750 ;
        RECT 39.580 85.150 43.530 85.300 ;
        RECT 43.130 84.700 43.530 85.150 ;
        RECT 39.580 84.550 43.530 84.700 ;
        RECT 43.130 84.400 43.530 84.550 ;
        RECT 45.930 95.450 46.330 95.600 ;
        RECT 45.930 95.300 49.880 95.450 ;
        RECT 45.930 94.850 46.330 95.300 ;
        RECT 45.930 94.700 49.880 94.850 ;
        RECT 45.930 94.250 46.330 94.700 ;
        RECT 45.930 94.100 49.880 94.250 ;
        RECT 45.930 93.650 46.330 94.100 ;
        RECT 45.930 93.500 49.880 93.650 ;
        RECT 45.930 93.050 46.330 93.500 ;
        RECT 45.930 92.900 49.880 93.050 ;
        RECT 45.930 92.450 46.330 92.900 ;
        RECT 45.930 92.300 49.880 92.450 ;
        RECT 45.930 91.850 46.330 92.300 ;
        RECT 45.930 91.700 49.880 91.850 ;
        RECT 45.930 91.250 46.330 91.700 ;
        RECT 45.930 91.100 49.880 91.250 ;
        RECT 45.930 90.650 46.330 91.100 ;
        RECT 45.930 90.500 49.880 90.650 ;
        RECT 45.930 90.200 46.330 90.500 ;
        RECT 50.480 90.200 50.630 98.400 ;
        RECT 51.080 90.200 51.230 98.400 ;
        RECT 51.680 90.200 51.830 98.400 ;
        RECT 52.280 90.200 52.430 98.400 ;
        RECT 52.880 90.200 53.030 98.400 ;
        RECT 53.480 90.200 53.630 98.400 ;
        RECT 54.080 90.200 54.230 98.400 ;
        RECT 45.930 89.800 54.230 90.200 ;
        RECT 45.930 89.500 46.330 89.800 ;
        RECT 45.930 89.350 49.880 89.500 ;
        RECT 45.930 88.900 46.330 89.350 ;
        RECT 45.930 88.750 49.880 88.900 ;
        RECT 45.930 88.300 46.330 88.750 ;
        RECT 45.930 88.150 49.880 88.300 ;
        RECT 45.930 87.700 46.330 88.150 ;
        RECT 45.930 87.550 49.880 87.700 ;
        RECT 45.930 87.100 46.330 87.550 ;
        RECT 45.930 86.950 49.880 87.100 ;
        RECT 45.930 86.500 46.330 86.950 ;
        RECT 45.930 86.350 49.880 86.500 ;
        RECT 45.930 85.900 46.330 86.350 ;
        RECT 45.930 85.750 49.880 85.900 ;
        RECT 45.930 85.300 46.330 85.750 ;
        RECT 45.930 85.150 49.880 85.300 ;
        RECT 45.930 84.700 46.330 85.150 ;
        RECT 45.930 84.550 49.880 84.700 ;
        RECT 45.930 84.400 46.330 84.550 ;
        RECT 43.130 84.100 46.330 84.400 ;
        RECT 39.580 83.950 49.880 84.100 ;
        RECT 43.130 83.500 46.330 83.950 ;
        RECT 39.580 83.350 49.880 83.500 ;
        RECT 43.130 82.900 46.330 83.350 ;
        RECT 39.580 82.750 49.880 82.900 ;
        RECT 43.130 82.300 46.330 82.750 ;
        RECT 39.580 82.150 49.880 82.300 ;
        RECT 43.530 81.200 45.930 82.150 ;
        RECT 50.480 81.600 50.630 89.800 ;
        RECT 51.080 81.600 51.230 89.800 ;
        RECT 51.680 81.600 51.830 89.800 ;
        RECT 52.280 81.600 52.430 89.800 ;
        RECT 52.880 81.600 53.030 89.800 ;
        RECT 53.480 81.600 53.630 89.800 ;
        RECT 54.080 81.600 54.230 89.800 ;
        RECT 55.230 90.200 55.380 98.400 ;
        RECT 55.830 90.200 55.980 98.400 ;
        RECT 56.430 90.200 56.580 98.400 ;
        RECT 57.030 90.200 57.180 98.400 ;
        RECT 57.630 90.200 57.780 98.400 ;
        RECT 58.230 90.200 58.380 98.400 ;
        RECT 58.830 90.200 58.980 98.400 ;
        RECT 63.530 97.850 65.940 98.800 ;
        RECT 59.580 97.700 69.880 97.850 ;
        RECT 63.130 97.250 66.330 97.700 ;
        RECT 59.580 97.100 69.880 97.250 ;
        RECT 63.130 96.650 66.330 97.100 ;
        RECT 59.580 96.500 69.880 96.650 ;
        RECT 63.130 96.050 66.330 96.500 ;
        RECT 59.580 95.900 69.880 96.050 ;
        RECT 63.130 95.600 66.330 95.900 ;
        RECT 63.130 95.450 63.530 95.600 ;
        RECT 59.580 95.300 63.530 95.450 ;
        RECT 63.130 94.850 63.530 95.300 ;
        RECT 59.580 94.700 63.530 94.850 ;
        RECT 63.130 94.250 63.530 94.700 ;
        RECT 59.580 94.100 63.530 94.250 ;
        RECT 63.130 93.650 63.530 94.100 ;
        RECT 59.580 93.500 63.530 93.650 ;
        RECT 63.130 93.050 63.530 93.500 ;
        RECT 59.580 92.900 63.530 93.050 ;
        RECT 63.130 92.450 63.530 92.900 ;
        RECT 59.580 92.300 63.530 92.450 ;
        RECT 63.130 91.850 63.530 92.300 ;
        RECT 59.580 91.700 63.530 91.850 ;
        RECT 63.130 91.250 63.530 91.700 ;
        RECT 59.580 91.100 63.530 91.250 ;
        RECT 63.130 90.650 63.530 91.100 ;
        RECT 59.580 90.500 63.530 90.650 ;
        RECT 63.130 90.200 63.530 90.500 ;
        RECT 55.230 89.800 63.530 90.200 ;
        RECT 55.230 81.600 55.380 89.800 ;
        RECT 55.830 81.600 55.980 89.800 ;
        RECT 56.430 81.600 56.580 89.800 ;
        RECT 57.030 81.600 57.180 89.800 ;
        RECT 57.630 81.600 57.780 89.800 ;
        RECT 58.230 81.600 58.380 89.800 ;
        RECT 58.830 81.600 58.980 89.800 ;
        RECT 63.130 89.500 63.530 89.800 ;
        RECT 59.580 89.350 63.530 89.500 ;
        RECT 63.130 88.900 63.530 89.350 ;
        RECT 59.580 88.750 63.530 88.900 ;
        RECT 63.130 88.300 63.530 88.750 ;
        RECT 59.580 88.150 63.530 88.300 ;
        RECT 63.130 87.700 63.530 88.150 ;
        RECT 59.580 87.550 63.530 87.700 ;
        RECT 63.130 87.100 63.530 87.550 ;
        RECT 59.580 86.950 63.530 87.100 ;
        RECT 63.130 86.500 63.530 86.950 ;
        RECT 59.580 86.350 63.530 86.500 ;
        RECT 63.130 85.900 63.530 86.350 ;
        RECT 59.580 85.750 63.530 85.900 ;
        RECT 63.130 85.300 63.530 85.750 ;
        RECT 59.580 85.150 63.530 85.300 ;
        RECT 63.130 84.700 63.530 85.150 ;
        RECT 59.580 84.550 63.530 84.700 ;
        RECT 63.130 84.400 63.530 84.550 ;
        RECT 65.930 95.450 66.330 95.600 ;
        RECT 65.930 95.300 69.880 95.450 ;
        RECT 65.930 94.850 66.330 95.300 ;
        RECT 65.930 94.700 69.880 94.850 ;
        RECT 65.930 94.250 66.330 94.700 ;
        RECT 65.930 94.100 69.880 94.250 ;
        RECT 65.930 93.650 66.330 94.100 ;
        RECT 65.930 93.500 69.880 93.650 ;
        RECT 65.930 93.050 66.330 93.500 ;
        RECT 65.930 92.900 69.880 93.050 ;
        RECT 65.930 92.450 66.330 92.900 ;
        RECT 65.930 92.300 69.880 92.450 ;
        RECT 65.930 91.850 66.330 92.300 ;
        RECT 65.930 91.700 69.880 91.850 ;
        RECT 65.930 91.250 66.330 91.700 ;
        RECT 65.930 91.100 69.880 91.250 ;
        RECT 65.930 90.650 66.330 91.100 ;
        RECT 65.930 90.500 69.880 90.650 ;
        RECT 65.930 90.200 66.330 90.500 ;
        RECT 70.480 90.200 70.630 98.400 ;
        RECT 71.080 90.200 71.230 98.400 ;
        RECT 71.680 90.200 71.830 98.400 ;
        RECT 72.280 90.200 72.430 98.400 ;
        RECT 72.880 90.200 73.030 98.400 ;
        RECT 73.480 90.200 73.630 98.400 ;
        RECT 74.080 90.200 74.230 98.400 ;
        RECT 65.930 89.800 74.230 90.200 ;
        RECT 65.930 89.500 66.330 89.800 ;
        RECT 65.930 89.350 69.880 89.500 ;
        RECT 65.930 88.900 66.330 89.350 ;
        RECT 65.930 88.750 69.880 88.900 ;
        RECT 65.930 88.300 66.330 88.750 ;
        RECT 65.930 88.150 69.880 88.300 ;
        RECT 65.930 87.700 66.330 88.150 ;
        RECT 65.930 87.550 69.880 87.700 ;
        RECT 65.930 87.100 66.330 87.550 ;
        RECT 65.930 86.950 69.880 87.100 ;
        RECT 65.930 86.500 66.330 86.950 ;
        RECT 65.930 86.350 69.880 86.500 ;
        RECT 65.930 85.900 66.330 86.350 ;
        RECT 65.930 85.750 69.880 85.900 ;
        RECT 65.930 85.300 66.330 85.750 ;
        RECT 65.930 85.150 69.880 85.300 ;
        RECT 65.930 84.700 66.330 85.150 ;
        RECT 65.930 84.550 69.880 84.700 ;
        RECT 65.930 84.400 66.330 84.550 ;
        RECT 63.130 84.100 66.330 84.400 ;
        RECT 59.580 83.950 69.880 84.100 ;
        RECT 63.130 83.500 66.330 83.950 ;
        RECT 59.580 83.350 69.880 83.500 ;
        RECT 63.130 82.900 66.330 83.350 ;
        RECT 59.580 82.750 69.880 82.900 ;
        RECT 63.130 82.300 66.330 82.750 ;
        RECT 59.580 82.150 69.880 82.300 ;
        RECT 63.530 81.200 65.930 82.150 ;
        RECT 70.480 81.600 70.630 89.800 ;
        RECT 71.080 81.600 71.230 89.800 ;
        RECT 71.680 81.600 71.830 89.800 ;
        RECT 72.280 81.600 72.430 89.800 ;
        RECT 72.880 81.600 73.030 89.800 ;
        RECT 73.480 81.600 73.630 89.800 ;
        RECT 74.080 81.600 74.230 89.800 ;
        RECT 75.230 90.200 75.380 98.400 ;
        RECT 75.830 90.200 75.980 98.400 ;
        RECT 76.430 90.200 76.580 98.400 ;
        RECT 77.030 90.200 77.180 98.400 ;
        RECT 77.630 90.200 77.780 98.400 ;
        RECT 78.230 90.200 78.380 98.400 ;
        RECT 78.830 90.200 78.980 98.400 ;
        RECT 83.530 97.850 85.940 98.800 ;
        RECT 79.580 97.700 89.880 97.850 ;
        RECT 83.130 97.250 86.330 97.700 ;
        RECT 79.580 97.100 89.880 97.250 ;
        RECT 83.130 96.650 86.330 97.100 ;
        RECT 79.580 96.500 89.880 96.650 ;
        RECT 83.130 96.050 86.330 96.500 ;
        RECT 79.580 95.900 89.880 96.050 ;
        RECT 83.130 95.600 86.330 95.900 ;
        RECT 83.130 95.450 83.530 95.600 ;
        RECT 79.580 95.300 83.530 95.450 ;
        RECT 83.130 94.850 83.530 95.300 ;
        RECT 79.580 94.700 83.530 94.850 ;
        RECT 83.130 94.250 83.530 94.700 ;
        RECT 79.580 94.100 83.530 94.250 ;
        RECT 83.130 93.650 83.530 94.100 ;
        RECT 79.580 93.500 83.530 93.650 ;
        RECT 83.130 93.050 83.530 93.500 ;
        RECT 79.580 92.900 83.530 93.050 ;
        RECT 83.130 92.450 83.530 92.900 ;
        RECT 79.580 92.300 83.530 92.450 ;
        RECT 83.130 91.850 83.530 92.300 ;
        RECT 79.580 91.700 83.530 91.850 ;
        RECT 83.130 91.250 83.530 91.700 ;
        RECT 79.580 91.100 83.530 91.250 ;
        RECT 83.130 90.650 83.530 91.100 ;
        RECT 79.580 90.500 83.530 90.650 ;
        RECT 83.130 90.200 83.530 90.500 ;
        RECT 75.230 89.800 83.530 90.200 ;
        RECT 75.230 81.600 75.380 89.800 ;
        RECT 75.830 81.600 75.980 89.800 ;
        RECT 76.430 81.600 76.580 89.800 ;
        RECT 77.030 81.600 77.180 89.800 ;
        RECT 77.630 81.600 77.780 89.800 ;
        RECT 78.230 81.600 78.380 89.800 ;
        RECT 78.830 81.600 78.980 89.800 ;
        RECT 83.130 89.500 83.530 89.800 ;
        RECT 79.580 89.350 83.530 89.500 ;
        RECT 83.130 88.900 83.530 89.350 ;
        RECT 79.580 88.750 83.530 88.900 ;
        RECT 83.130 88.300 83.530 88.750 ;
        RECT 79.580 88.150 83.530 88.300 ;
        RECT 83.130 87.700 83.530 88.150 ;
        RECT 79.580 87.550 83.530 87.700 ;
        RECT 83.130 87.100 83.530 87.550 ;
        RECT 79.580 86.950 83.530 87.100 ;
        RECT 83.130 86.500 83.530 86.950 ;
        RECT 79.580 86.350 83.530 86.500 ;
        RECT 83.130 85.900 83.530 86.350 ;
        RECT 79.580 85.750 83.530 85.900 ;
        RECT 83.130 85.300 83.530 85.750 ;
        RECT 79.580 85.150 83.530 85.300 ;
        RECT 83.130 84.700 83.530 85.150 ;
        RECT 79.580 84.550 83.530 84.700 ;
        RECT 83.130 84.400 83.530 84.550 ;
        RECT 85.930 95.450 86.330 95.600 ;
        RECT 85.930 95.300 89.880 95.450 ;
        RECT 85.930 94.850 86.330 95.300 ;
        RECT 85.930 94.700 89.880 94.850 ;
        RECT 85.930 94.250 86.330 94.700 ;
        RECT 85.930 94.100 89.880 94.250 ;
        RECT 85.930 93.650 86.330 94.100 ;
        RECT 85.930 93.500 89.880 93.650 ;
        RECT 85.930 93.050 86.330 93.500 ;
        RECT 85.930 92.900 89.880 93.050 ;
        RECT 85.930 92.450 86.330 92.900 ;
        RECT 85.930 92.300 89.880 92.450 ;
        RECT 85.930 91.850 86.330 92.300 ;
        RECT 85.930 91.700 89.880 91.850 ;
        RECT 85.930 91.250 86.330 91.700 ;
        RECT 85.930 91.100 89.880 91.250 ;
        RECT 85.930 90.650 86.330 91.100 ;
        RECT 85.930 90.500 89.880 90.650 ;
        RECT 85.930 90.200 86.330 90.500 ;
        RECT 90.480 90.200 90.630 98.400 ;
        RECT 91.080 90.200 91.230 98.400 ;
        RECT 91.680 90.200 91.830 98.400 ;
        RECT 92.280 90.200 92.430 98.400 ;
        RECT 92.880 90.200 93.030 98.400 ;
        RECT 93.480 90.200 93.630 98.400 ;
        RECT 94.080 90.200 94.230 98.400 ;
        RECT 85.930 89.800 94.230 90.200 ;
        RECT 85.930 89.500 86.330 89.800 ;
        RECT 85.930 89.350 89.880 89.500 ;
        RECT 85.930 88.900 86.330 89.350 ;
        RECT 85.930 88.750 89.880 88.900 ;
        RECT 85.930 88.300 86.330 88.750 ;
        RECT 85.930 88.150 89.880 88.300 ;
        RECT 85.930 87.700 86.330 88.150 ;
        RECT 85.930 87.550 89.880 87.700 ;
        RECT 85.930 87.100 86.330 87.550 ;
        RECT 85.930 86.950 89.880 87.100 ;
        RECT 85.930 86.500 86.330 86.950 ;
        RECT 85.930 86.350 89.880 86.500 ;
        RECT 85.930 85.900 86.330 86.350 ;
        RECT 85.930 85.750 89.880 85.900 ;
        RECT 85.930 85.300 86.330 85.750 ;
        RECT 85.930 85.150 89.880 85.300 ;
        RECT 85.930 84.700 86.330 85.150 ;
        RECT 85.930 84.550 89.880 84.700 ;
        RECT 85.930 84.400 86.330 84.550 ;
        RECT 83.130 84.100 86.330 84.400 ;
        RECT 79.580 83.950 89.880 84.100 ;
        RECT 83.130 83.500 86.330 83.950 ;
        RECT 79.580 83.350 89.880 83.500 ;
        RECT 83.130 82.900 86.330 83.350 ;
        RECT 79.580 82.750 89.880 82.900 ;
        RECT 83.130 82.300 86.330 82.750 ;
        RECT 79.580 82.150 89.880 82.300 ;
        RECT 83.530 81.200 85.930 82.150 ;
        RECT 90.480 81.600 90.630 89.800 ;
        RECT 91.080 81.600 91.230 89.800 ;
        RECT 91.680 81.600 91.830 89.800 ;
        RECT 92.280 81.600 92.430 89.800 ;
        RECT 92.880 81.600 93.030 89.800 ;
        RECT 93.480 81.600 93.630 89.800 ;
        RECT 94.080 81.600 94.230 89.800 ;
        RECT 95.230 90.200 95.380 98.400 ;
        RECT 95.830 90.200 95.980 98.400 ;
        RECT 96.430 90.200 96.580 98.400 ;
        RECT 97.030 90.200 97.180 98.400 ;
        RECT 97.630 90.200 97.780 98.400 ;
        RECT 98.230 90.200 98.380 98.400 ;
        RECT 98.830 90.200 98.980 98.400 ;
        RECT 103.530 97.850 104.730 98.800 ;
        RECT 99.580 97.700 104.730 97.850 ;
        RECT 103.130 97.250 104.730 97.700 ;
        RECT 99.580 97.100 104.730 97.250 ;
        RECT 103.130 96.650 104.730 97.100 ;
        RECT 99.580 96.500 104.730 96.650 ;
        RECT 103.130 96.050 104.730 96.500 ;
        RECT 99.580 95.900 104.730 96.050 ;
        RECT 105.135 95.910 107.135 97.185 ;
        RECT 103.130 95.600 104.730 95.900 ;
        RECT 103.130 95.450 103.530 95.600 ;
        RECT 99.580 95.300 103.530 95.450 ;
        RECT 103.130 94.850 103.530 95.300 ;
        RECT 99.580 94.700 103.530 94.850 ;
        RECT 103.130 94.250 103.530 94.700 ;
        RECT 99.580 94.100 103.530 94.250 ;
        RECT 103.130 93.650 103.530 94.100 ;
        RECT 99.580 93.500 103.530 93.650 ;
        RECT 103.130 93.050 103.530 93.500 ;
        RECT 99.580 92.900 103.530 93.050 ;
        RECT 103.130 92.450 103.530 92.900 ;
        RECT 99.580 92.300 103.530 92.450 ;
        RECT 103.130 91.850 103.530 92.300 ;
        RECT 99.580 91.700 103.530 91.850 ;
        RECT 103.130 91.250 103.530 91.700 ;
        RECT 99.580 91.100 103.530 91.250 ;
        RECT 103.130 90.650 103.530 91.100 ;
        RECT 99.580 90.500 103.530 90.650 ;
        RECT 103.130 90.200 103.530 90.500 ;
        RECT 95.230 89.800 103.530 90.200 ;
        RECT 95.230 81.600 95.380 89.800 ;
        RECT 95.830 81.600 95.980 89.800 ;
        RECT 96.430 81.600 96.580 89.800 ;
        RECT 97.030 81.600 97.180 89.800 ;
        RECT 97.630 81.600 97.780 89.800 ;
        RECT 98.230 81.600 98.380 89.800 ;
        RECT 98.830 81.600 98.980 89.800 ;
        RECT 103.130 89.500 103.530 89.800 ;
        RECT 99.580 89.350 103.530 89.500 ;
        RECT 103.130 88.900 103.530 89.350 ;
        RECT 99.580 88.750 103.530 88.900 ;
        RECT 103.130 88.300 103.530 88.750 ;
        RECT 99.580 88.150 103.530 88.300 ;
        RECT 103.130 87.700 103.530 88.150 ;
        RECT 99.580 87.550 103.530 87.700 ;
        RECT 103.130 87.100 103.530 87.550 ;
        RECT 99.580 86.950 103.530 87.100 ;
        RECT 103.130 86.500 103.530 86.950 ;
        RECT 99.580 86.350 103.530 86.500 ;
        RECT 103.130 85.900 103.530 86.350 ;
        RECT 99.580 85.750 103.530 85.900 ;
        RECT 103.130 85.300 103.530 85.750 ;
        RECT 99.580 85.150 103.530 85.300 ;
        RECT 103.130 84.700 103.530 85.150 ;
        RECT 99.580 84.550 103.530 84.700 ;
        RECT 103.130 84.400 103.530 84.550 ;
        RECT 103.130 84.100 104.730 84.400 ;
        RECT 99.580 83.950 104.730 84.100 ;
        RECT 103.130 83.500 104.730 83.950 ;
        RECT 99.580 83.350 104.730 83.500 ;
        RECT 103.130 82.900 104.730 83.350 ;
        RECT 99.580 82.750 104.730 82.900 ;
        RECT 103.130 82.300 104.730 82.750 ;
        RECT 99.580 82.150 104.730 82.300 ;
        RECT 103.530 81.200 104.730 82.150 ;
        RECT 105.135 82.105 107.135 83.380 ;
        RECT 4.730 78.800 9.130 81.200 ;
        RECT 20.330 78.800 29.130 81.200 ;
        RECT 40.330 78.800 49.130 81.200 ;
        RECT 60.330 78.800 69.130 81.200 ;
        RECT 80.330 78.800 89.130 81.200 ;
        RECT 100.330 78.800 104.730 81.200 ;
        RECT 4.730 77.850 5.940 78.800 ;
        RECT 4.730 77.700 9.880 77.850 ;
        RECT 2.315 76.280 4.330 77.555 ;
        RECT 4.730 77.250 6.330 77.700 ;
        RECT 4.730 77.100 9.880 77.250 ;
        RECT 4.730 76.650 6.330 77.100 ;
        RECT 4.730 76.500 9.880 76.650 ;
        RECT 4.730 76.050 6.330 76.500 ;
        RECT 4.730 75.900 9.880 76.050 ;
        RECT 4.730 75.600 6.330 75.900 ;
        RECT 2.315 73.250 4.315 75.545 ;
        RECT 5.930 75.450 6.330 75.600 ;
        RECT 5.930 75.300 9.880 75.450 ;
        RECT 5.930 74.850 6.330 75.300 ;
        RECT 5.930 74.700 9.880 74.850 ;
        RECT 5.930 74.250 6.330 74.700 ;
        RECT 5.930 74.100 9.880 74.250 ;
        RECT 5.930 73.650 6.330 74.100 ;
        RECT 5.930 73.500 9.880 73.650 ;
        RECT 5.930 73.050 6.330 73.500 ;
        RECT 5.930 72.900 9.880 73.050 ;
        RECT 5.930 72.450 6.330 72.900 ;
        RECT 5.930 72.300 9.880 72.450 ;
        RECT 5.930 71.850 6.330 72.300 ;
        RECT 5.930 71.700 9.880 71.850 ;
        RECT 5.930 71.250 6.330 71.700 ;
        RECT 5.930 71.100 9.880 71.250 ;
        RECT 5.930 70.650 6.330 71.100 ;
        RECT 5.930 70.500 9.880 70.650 ;
        RECT 5.930 70.200 6.330 70.500 ;
        RECT 10.480 70.200 10.630 78.400 ;
        RECT 11.080 70.200 11.230 78.400 ;
        RECT 11.680 70.200 11.830 78.400 ;
        RECT 12.280 70.200 12.430 78.400 ;
        RECT 12.880 70.200 13.030 78.400 ;
        RECT 13.480 70.200 13.630 78.400 ;
        RECT 14.080 70.200 14.230 78.400 ;
        RECT 5.930 69.800 14.230 70.200 ;
        RECT 5.930 69.500 6.330 69.800 ;
        RECT 5.930 69.350 9.880 69.500 ;
        RECT 5.930 68.900 6.330 69.350 ;
        RECT 5.930 68.750 9.880 68.900 ;
        RECT 5.930 68.300 6.330 68.750 ;
        RECT 5.930 68.150 9.880 68.300 ;
        RECT 5.930 67.700 6.330 68.150 ;
        RECT 5.930 67.550 9.880 67.700 ;
        RECT 5.930 67.100 6.330 67.550 ;
        RECT 5.930 66.950 9.880 67.100 ;
        RECT 2.315 64.450 4.315 66.745 ;
        RECT 5.930 66.500 6.330 66.950 ;
        RECT 5.930 66.350 9.880 66.500 ;
        RECT 5.930 65.900 6.330 66.350 ;
        RECT 5.930 65.750 9.880 65.900 ;
        RECT 5.930 65.300 6.330 65.750 ;
        RECT 5.930 65.150 9.880 65.300 ;
        RECT 5.930 64.700 6.330 65.150 ;
        RECT 5.930 64.550 9.880 64.700 ;
        RECT 5.930 64.400 6.330 64.550 ;
        RECT 4.730 64.100 6.330 64.400 ;
        RECT 4.730 63.950 9.880 64.100 ;
        RECT 4.730 63.500 6.330 63.950 ;
        RECT 4.730 63.350 9.880 63.500 ;
        RECT 2.315 61.955 4.320 63.230 ;
        RECT 4.730 62.900 6.330 63.350 ;
        RECT 4.730 62.750 9.880 62.900 ;
        RECT 4.730 62.300 6.330 62.750 ;
        RECT 4.730 62.150 9.880 62.300 ;
        RECT 4.730 61.200 5.930 62.150 ;
        RECT 10.480 61.600 10.630 69.800 ;
        RECT 11.080 61.600 11.230 69.800 ;
        RECT 11.680 61.600 11.830 69.800 ;
        RECT 12.280 61.600 12.430 69.800 ;
        RECT 12.880 61.600 13.030 69.800 ;
        RECT 13.480 61.600 13.630 69.800 ;
        RECT 14.080 61.600 14.230 69.800 ;
        RECT 15.230 70.200 15.380 78.400 ;
        RECT 15.830 70.200 15.980 78.400 ;
        RECT 16.430 70.200 16.580 78.400 ;
        RECT 17.030 70.200 17.180 78.400 ;
        RECT 17.630 70.200 17.780 78.400 ;
        RECT 18.230 70.200 18.380 78.400 ;
        RECT 18.830 70.200 18.980 78.400 ;
        RECT 23.530 77.850 25.940 78.800 ;
        RECT 19.580 77.700 29.880 77.850 ;
        RECT 23.130 77.250 26.330 77.700 ;
        RECT 19.580 77.100 29.880 77.250 ;
        RECT 23.130 76.650 26.330 77.100 ;
        RECT 19.580 76.500 29.880 76.650 ;
        RECT 23.130 76.050 26.330 76.500 ;
        RECT 19.580 75.900 29.880 76.050 ;
        RECT 23.130 75.600 26.330 75.900 ;
        RECT 23.130 75.450 23.530 75.600 ;
        RECT 19.580 75.300 23.530 75.450 ;
        RECT 23.130 74.850 23.530 75.300 ;
        RECT 19.580 74.700 23.530 74.850 ;
        RECT 23.130 74.250 23.530 74.700 ;
        RECT 19.580 74.100 23.530 74.250 ;
        RECT 23.130 73.650 23.530 74.100 ;
        RECT 19.580 73.500 23.530 73.650 ;
        RECT 23.130 73.050 23.530 73.500 ;
        RECT 19.580 72.900 23.530 73.050 ;
        RECT 23.130 72.450 23.530 72.900 ;
        RECT 19.580 72.300 23.530 72.450 ;
        RECT 23.130 71.850 23.530 72.300 ;
        RECT 19.580 71.700 23.530 71.850 ;
        RECT 23.130 71.250 23.530 71.700 ;
        RECT 19.580 71.100 23.530 71.250 ;
        RECT 23.130 70.650 23.530 71.100 ;
        RECT 19.580 70.500 23.530 70.650 ;
        RECT 23.130 70.200 23.530 70.500 ;
        RECT 15.230 69.800 23.530 70.200 ;
        RECT 15.230 61.600 15.380 69.800 ;
        RECT 15.830 61.600 15.980 69.800 ;
        RECT 16.430 61.600 16.580 69.800 ;
        RECT 17.030 61.600 17.180 69.800 ;
        RECT 17.630 61.600 17.780 69.800 ;
        RECT 18.230 61.600 18.380 69.800 ;
        RECT 18.830 61.600 18.980 69.800 ;
        RECT 23.130 69.500 23.530 69.800 ;
        RECT 19.580 69.350 23.530 69.500 ;
        RECT 23.130 68.900 23.530 69.350 ;
        RECT 19.580 68.750 23.530 68.900 ;
        RECT 23.130 68.300 23.530 68.750 ;
        RECT 19.580 68.150 23.530 68.300 ;
        RECT 23.130 67.700 23.530 68.150 ;
        RECT 19.580 67.550 23.530 67.700 ;
        RECT 23.130 67.100 23.530 67.550 ;
        RECT 19.580 66.950 23.530 67.100 ;
        RECT 23.130 66.500 23.530 66.950 ;
        RECT 19.580 66.350 23.530 66.500 ;
        RECT 23.130 65.900 23.530 66.350 ;
        RECT 19.580 65.750 23.530 65.900 ;
        RECT 23.130 65.300 23.530 65.750 ;
        RECT 19.580 65.150 23.530 65.300 ;
        RECT 23.130 64.700 23.530 65.150 ;
        RECT 19.580 64.550 23.530 64.700 ;
        RECT 23.130 64.400 23.530 64.550 ;
        RECT 25.930 75.450 26.330 75.600 ;
        RECT 25.930 75.300 29.880 75.450 ;
        RECT 25.930 74.850 26.330 75.300 ;
        RECT 25.930 74.700 29.880 74.850 ;
        RECT 25.930 74.250 26.330 74.700 ;
        RECT 25.930 74.100 29.880 74.250 ;
        RECT 25.930 73.650 26.330 74.100 ;
        RECT 25.930 73.500 29.880 73.650 ;
        RECT 25.930 73.050 26.330 73.500 ;
        RECT 25.930 72.900 29.880 73.050 ;
        RECT 25.930 72.450 26.330 72.900 ;
        RECT 25.930 72.300 29.880 72.450 ;
        RECT 25.930 71.850 26.330 72.300 ;
        RECT 25.930 71.700 29.880 71.850 ;
        RECT 25.930 71.250 26.330 71.700 ;
        RECT 25.930 71.100 29.880 71.250 ;
        RECT 25.930 70.650 26.330 71.100 ;
        RECT 25.930 70.500 29.880 70.650 ;
        RECT 25.930 70.200 26.330 70.500 ;
        RECT 30.480 70.200 30.630 78.400 ;
        RECT 31.080 70.200 31.230 78.400 ;
        RECT 31.680 70.200 31.830 78.400 ;
        RECT 32.280 70.200 32.430 78.400 ;
        RECT 32.880 70.200 33.030 78.400 ;
        RECT 33.480 70.200 33.630 78.400 ;
        RECT 34.080 70.200 34.230 78.400 ;
        RECT 25.930 69.800 34.230 70.200 ;
        RECT 25.930 69.500 26.330 69.800 ;
        RECT 25.930 69.350 29.880 69.500 ;
        RECT 25.930 68.900 26.330 69.350 ;
        RECT 25.930 68.750 29.880 68.900 ;
        RECT 25.930 68.300 26.330 68.750 ;
        RECT 25.930 68.150 29.880 68.300 ;
        RECT 25.930 67.700 26.330 68.150 ;
        RECT 25.930 67.550 29.880 67.700 ;
        RECT 25.930 67.100 26.330 67.550 ;
        RECT 25.930 66.950 29.880 67.100 ;
        RECT 25.930 66.500 26.330 66.950 ;
        RECT 25.930 66.350 29.880 66.500 ;
        RECT 25.930 65.900 26.330 66.350 ;
        RECT 25.930 65.750 29.880 65.900 ;
        RECT 25.930 65.300 26.330 65.750 ;
        RECT 25.930 65.150 29.880 65.300 ;
        RECT 25.930 64.700 26.330 65.150 ;
        RECT 25.930 64.550 29.880 64.700 ;
        RECT 25.930 64.400 26.330 64.550 ;
        RECT 23.130 64.100 26.330 64.400 ;
        RECT 19.580 63.950 29.880 64.100 ;
        RECT 23.130 63.500 26.330 63.950 ;
        RECT 19.580 63.350 29.880 63.500 ;
        RECT 23.130 62.900 26.330 63.350 ;
        RECT 19.580 62.750 29.880 62.900 ;
        RECT 23.130 62.300 26.330 62.750 ;
        RECT 19.580 62.150 29.880 62.300 ;
        RECT 23.530 61.200 25.930 62.150 ;
        RECT 30.480 61.600 30.630 69.800 ;
        RECT 31.080 61.600 31.230 69.800 ;
        RECT 31.680 61.600 31.830 69.800 ;
        RECT 32.280 61.600 32.430 69.800 ;
        RECT 32.880 61.600 33.030 69.800 ;
        RECT 33.480 61.600 33.630 69.800 ;
        RECT 34.080 61.600 34.230 69.800 ;
        RECT 35.230 70.200 35.380 78.400 ;
        RECT 35.830 70.200 35.980 78.400 ;
        RECT 36.430 70.200 36.580 78.400 ;
        RECT 37.030 70.200 37.180 78.400 ;
        RECT 37.630 70.200 37.780 78.400 ;
        RECT 38.230 70.200 38.380 78.400 ;
        RECT 38.830 70.200 38.980 78.400 ;
        RECT 43.530 77.850 45.940 78.800 ;
        RECT 39.580 77.700 49.880 77.850 ;
        RECT 43.130 77.250 46.330 77.700 ;
        RECT 39.580 77.100 49.880 77.250 ;
        RECT 43.130 76.650 46.330 77.100 ;
        RECT 39.580 76.500 49.880 76.650 ;
        RECT 43.130 76.050 46.330 76.500 ;
        RECT 39.580 75.900 49.880 76.050 ;
        RECT 43.130 75.600 46.330 75.900 ;
        RECT 43.130 75.450 43.530 75.600 ;
        RECT 39.580 75.300 43.530 75.450 ;
        RECT 43.130 74.850 43.530 75.300 ;
        RECT 39.580 74.700 43.530 74.850 ;
        RECT 43.130 74.250 43.530 74.700 ;
        RECT 39.580 74.100 43.530 74.250 ;
        RECT 43.130 73.650 43.530 74.100 ;
        RECT 39.580 73.500 43.530 73.650 ;
        RECT 43.130 73.050 43.530 73.500 ;
        RECT 39.580 72.900 43.530 73.050 ;
        RECT 43.130 72.450 43.530 72.900 ;
        RECT 39.580 72.300 43.530 72.450 ;
        RECT 43.130 71.850 43.530 72.300 ;
        RECT 39.580 71.700 43.530 71.850 ;
        RECT 43.130 71.250 43.530 71.700 ;
        RECT 39.580 71.100 43.530 71.250 ;
        RECT 43.130 70.650 43.530 71.100 ;
        RECT 39.580 70.500 43.530 70.650 ;
        RECT 43.130 70.200 43.530 70.500 ;
        RECT 35.230 69.800 43.530 70.200 ;
        RECT 35.230 61.600 35.380 69.800 ;
        RECT 35.830 61.600 35.980 69.800 ;
        RECT 36.430 61.600 36.580 69.800 ;
        RECT 37.030 61.600 37.180 69.800 ;
        RECT 37.630 61.600 37.780 69.800 ;
        RECT 38.230 61.600 38.380 69.800 ;
        RECT 38.830 61.600 38.980 69.800 ;
        RECT 43.130 69.500 43.530 69.800 ;
        RECT 39.580 69.350 43.530 69.500 ;
        RECT 43.130 68.900 43.530 69.350 ;
        RECT 39.580 68.750 43.530 68.900 ;
        RECT 43.130 68.300 43.530 68.750 ;
        RECT 39.580 68.150 43.530 68.300 ;
        RECT 43.130 67.700 43.530 68.150 ;
        RECT 39.580 67.550 43.530 67.700 ;
        RECT 43.130 67.100 43.530 67.550 ;
        RECT 39.580 66.950 43.530 67.100 ;
        RECT 43.130 66.500 43.530 66.950 ;
        RECT 39.580 66.350 43.530 66.500 ;
        RECT 43.130 65.900 43.530 66.350 ;
        RECT 39.580 65.750 43.530 65.900 ;
        RECT 43.130 65.300 43.530 65.750 ;
        RECT 39.580 65.150 43.530 65.300 ;
        RECT 43.130 64.700 43.530 65.150 ;
        RECT 39.580 64.550 43.530 64.700 ;
        RECT 43.130 64.400 43.530 64.550 ;
        RECT 45.930 75.450 46.330 75.600 ;
        RECT 45.930 75.300 49.880 75.450 ;
        RECT 45.930 74.850 46.330 75.300 ;
        RECT 45.930 74.700 49.880 74.850 ;
        RECT 45.930 74.250 46.330 74.700 ;
        RECT 45.930 74.100 49.880 74.250 ;
        RECT 45.930 73.650 46.330 74.100 ;
        RECT 45.930 73.500 49.880 73.650 ;
        RECT 45.930 73.050 46.330 73.500 ;
        RECT 45.930 72.900 49.880 73.050 ;
        RECT 45.930 72.450 46.330 72.900 ;
        RECT 45.930 72.300 49.880 72.450 ;
        RECT 45.930 71.850 46.330 72.300 ;
        RECT 45.930 71.700 49.880 71.850 ;
        RECT 45.930 71.250 46.330 71.700 ;
        RECT 45.930 71.100 49.880 71.250 ;
        RECT 45.930 70.650 46.330 71.100 ;
        RECT 45.930 70.500 49.880 70.650 ;
        RECT 45.930 70.200 46.330 70.500 ;
        RECT 50.480 70.200 50.630 78.400 ;
        RECT 51.080 70.200 51.230 78.400 ;
        RECT 51.680 70.200 51.830 78.400 ;
        RECT 52.280 70.200 52.430 78.400 ;
        RECT 52.880 70.200 53.030 78.400 ;
        RECT 53.480 70.200 53.630 78.400 ;
        RECT 54.080 70.200 54.230 78.400 ;
        RECT 45.930 69.800 54.230 70.200 ;
        RECT 45.930 69.500 46.330 69.800 ;
        RECT 45.930 69.350 49.880 69.500 ;
        RECT 45.930 68.900 46.330 69.350 ;
        RECT 45.930 68.750 49.880 68.900 ;
        RECT 45.930 68.300 46.330 68.750 ;
        RECT 45.930 68.150 49.880 68.300 ;
        RECT 45.930 67.700 46.330 68.150 ;
        RECT 45.930 67.550 49.880 67.700 ;
        RECT 45.930 67.100 46.330 67.550 ;
        RECT 45.930 66.950 49.880 67.100 ;
        RECT 45.930 66.500 46.330 66.950 ;
        RECT 45.930 66.350 49.880 66.500 ;
        RECT 45.930 65.900 46.330 66.350 ;
        RECT 45.930 65.750 49.880 65.900 ;
        RECT 45.930 65.300 46.330 65.750 ;
        RECT 45.930 65.150 49.880 65.300 ;
        RECT 45.930 64.700 46.330 65.150 ;
        RECT 45.930 64.550 49.880 64.700 ;
        RECT 45.930 64.400 46.330 64.550 ;
        RECT 43.130 64.100 46.330 64.400 ;
        RECT 39.580 63.950 49.880 64.100 ;
        RECT 43.130 63.500 46.330 63.950 ;
        RECT 39.580 63.350 49.880 63.500 ;
        RECT 43.130 62.900 46.330 63.350 ;
        RECT 39.580 62.750 49.880 62.900 ;
        RECT 43.130 62.300 46.330 62.750 ;
        RECT 39.580 62.150 49.880 62.300 ;
        RECT 43.530 61.200 45.930 62.150 ;
        RECT 50.480 61.600 50.630 69.800 ;
        RECT 51.080 61.600 51.230 69.800 ;
        RECT 51.680 61.600 51.830 69.800 ;
        RECT 52.280 61.600 52.430 69.800 ;
        RECT 52.880 61.600 53.030 69.800 ;
        RECT 53.480 61.600 53.630 69.800 ;
        RECT 54.080 61.600 54.230 69.800 ;
        RECT 55.230 70.200 55.380 78.400 ;
        RECT 55.830 70.200 55.980 78.400 ;
        RECT 56.430 70.200 56.580 78.400 ;
        RECT 57.030 70.200 57.180 78.400 ;
        RECT 57.630 70.200 57.780 78.400 ;
        RECT 58.230 70.200 58.380 78.400 ;
        RECT 58.830 70.200 58.980 78.400 ;
        RECT 63.530 77.850 65.940 78.800 ;
        RECT 59.580 77.700 69.880 77.850 ;
        RECT 63.130 77.250 66.330 77.700 ;
        RECT 59.580 77.100 69.880 77.250 ;
        RECT 63.130 76.650 66.330 77.100 ;
        RECT 59.580 76.500 69.880 76.650 ;
        RECT 63.130 76.050 66.330 76.500 ;
        RECT 59.580 75.900 69.880 76.050 ;
        RECT 63.130 75.600 66.330 75.900 ;
        RECT 63.130 75.450 63.530 75.600 ;
        RECT 59.580 75.300 63.530 75.450 ;
        RECT 63.130 74.850 63.530 75.300 ;
        RECT 59.580 74.700 63.530 74.850 ;
        RECT 63.130 74.250 63.530 74.700 ;
        RECT 59.580 74.100 63.530 74.250 ;
        RECT 63.130 73.650 63.530 74.100 ;
        RECT 59.580 73.500 63.530 73.650 ;
        RECT 63.130 73.050 63.530 73.500 ;
        RECT 59.580 72.900 63.530 73.050 ;
        RECT 63.130 72.450 63.530 72.900 ;
        RECT 59.580 72.300 63.530 72.450 ;
        RECT 63.130 71.850 63.530 72.300 ;
        RECT 59.580 71.700 63.530 71.850 ;
        RECT 63.130 71.250 63.530 71.700 ;
        RECT 59.580 71.100 63.530 71.250 ;
        RECT 63.130 70.650 63.530 71.100 ;
        RECT 59.580 70.500 63.530 70.650 ;
        RECT 63.130 70.200 63.530 70.500 ;
        RECT 55.230 69.800 63.530 70.200 ;
        RECT 55.230 61.600 55.380 69.800 ;
        RECT 55.830 61.600 55.980 69.800 ;
        RECT 56.430 61.600 56.580 69.800 ;
        RECT 57.030 61.600 57.180 69.800 ;
        RECT 57.630 61.600 57.780 69.800 ;
        RECT 58.230 61.600 58.380 69.800 ;
        RECT 58.830 61.600 58.980 69.800 ;
        RECT 63.130 69.500 63.530 69.800 ;
        RECT 59.580 69.350 63.530 69.500 ;
        RECT 63.130 68.900 63.530 69.350 ;
        RECT 59.580 68.750 63.530 68.900 ;
        RECT 63.130 68.300 63.530 68.750 ;
        RECT 59.580 68.150 63.530 68.300 ;
        RECT 63.130 67.700 63.530 68.150 ;
        RECT 59.580 67.550 63.530 67.700 ;
        RECT 63.130 67.100 63.530 67.550 ;
        RECT 59.580 66.950 63.530 67.100 ;
        RECT 63.130 66.500 63.530 66.950 ;
        RECT 59.580 66.350 63.530 66.500 ;
        RECT 63.130 65.900 63.530 66.350 ;
        RECT 59.580 65.750 63.530 65.900 ;
        RECT 63.130 65.300 63.530 65.750 ;
        RECT 59.580 65.150 63.530 65.300 ;
        RECT 63.130 64.700 63.530 65.150 ;
        RECT 59.580 64.550 63.530 64.700 ;
        RECT 63.130 64.400 63.530 64.550 ;
        RECT 65.930 75.450 66.330 75.600 ;
        RECT 65.930 75.300 69.880 75.450 ;
        RECT 65.930 74.850 66.330 75.300 ;
        RECT 65.930 74.700 69.880 74.850 ;
        RECT 65.930 74.250 66.330 74.700 ;
        RECT 65.930 74.100 69.880 74.250 ;
        RECT 65.930 73.650 66.330 74.100 ;
        RECT 65.930 73.500 69.880 73.650 ;
        RECT 65.930 73.050 66.330 73.500 ;
        RECT 65.930 72.900 69.880 73.050 ;
        RECT 65.930 72.450 66.330 72.900 ;
        RECT 65.930 72.300 69.880 72.450 ;
        RECT 65.930 71.850 66.330 72.300 ;
        RECT 65.930 71.700 69.880 71.850 ;
        RECT 65.930 71.250 66.330 71.700 ;
        RECT 65.930 71.100 69.880 71.250 ;
        RECT 65.930 70.650 66.330 71.100 ;
        RECT 65.930 70.500 69.880 70.650 ;
        RECT 65.930 70.200 66.330 70.500 ;
        RECT 70.480 70.200 70.630 78.400 ;
        RECT 71.080 70.200 71.230 78.400 ;
        RECT 71.680 70.200 71.830 78.400 ;
        RECT 72.280 70.200 72.430 78.400 ;
        RECT 72.880 70.200 73.030 78.400 ;
        RECT 73.480 70.200 73.630 78.400 ;
        RECT 74.080 70.200 74.230 78.400 ;
        RECT 65.930 69.800 74.230 70.200 ;
        RECT 65.930 69.500 66.330 69.800 ;
        RECT 65.930 69.350 69.880 69.500 ;
        RECT 65.930 68.900 66.330 69.350 ;
        RECT 65.930 68.750 69.880 68.900 ;
        RECT 65.930 68.300 66.330 68.750 ;
        RECT 65.930 68.150 69.880 68.300 ;
        RECT 65.930 67.700 66.330 68.150 ;
        RECT 65.930 67.550 69.880 67.700 ;
        RECT 65.930 67.100 66.330 67.550 ;
        RECT 65.930 66.950 69.880 67.100 ;
        RECT 65.930 66.500 66.330 66.950 ;
        RECT 65.930 66.350 69.880 66.500 ;
        RECT 65.930 65.900 66.330 66.350 ;
        RECT 65.930 65.750 69.880 65.900 ;
        RECT 65.930 65.300 66.330 65.750 ;
        RECT 65.930 65.150 69.880 65.300 ;
        RECT 65.930 64.700 66.330 65.150 ;
        RECT 65.930 64.550 69.880 64.700 ;
        RECT 65.930 64.400 66.330 64.550 ;
        RECT 63.130 64.100 66.330 64.400 ;
        RECT 59.580 63.950 69.880 64.100 ;
        RECT 63.130 63.500 66.330 63.950 ;
        RECT 59.580 63.350 69.880 63.500 ;
        RECT 63.130 62.900 66.330 63.350 ;
        RECT 59.580 62.750 69.880 62.900 ;
        RECT 63.130 62.300 66.330 62.750 ;
        RECT 59.580 62.150 69.880 62.300 ;
        RECT 63.530 61.200 65.930 62.150 ;
        RECT 70.480 61.600 70.630 69.800 ;
        RECT 71.080 61.600 71.230 69.800 ;
        RECT 71.680 61.600 71.830 69.800 ;
        RECT 72.280 61.600 72.430 69.800 ;
        RECT 72.880 61.600 73.030 69.800 ;
        RECT 73.480 61.600 73.630 69.800 ;
        RECT 74.080 61.600 74.230 69.800 ;
        RECT 75.230 70.200 75.380 78.400 ;
        RECT 75.830 70.200 75.980 78.400 ;
        RECT 76.430 70.200 76.580 78.400 ;
        RECT 77.030 70.200 77.180 78.400 ;
        RECT 77.630 70.200 77.780 78.400 ;
        RECT 78.230 70.200 78.380 78.400 ;
        RECT 78.830 70.200 78.980 78.400 ;
        RECT 83.530 77.850 85.940 78.800 ;
        RECT 79.580 77.700 89.880 77.850 ;
        RECT 83.130 77.250 86.330 77.700 ;
        RECT 79.580 77.100 89.880 77.250 ;
        RECT 83.130 76.650 86.330 77.100 ;
        RECT 79.580 76.500 89.880 76.650 ;
        RECT 83.130 76.050 86.330 76.500 ;
        RECT 79.580 75.900 89.880 76.050 ;
        RECT 83.130 75.600 86.330 75.900 ;
        RECT 83.130 75.450 83.530 75.600 ;
        RECT 79.580 75.300 83.530 75.450 ;
        RECT 83.130 74.850 83.530 75.300 ;
        RECT 79.580 74.700 83.530 74.850 ;
        RECT 83.130 74.250 83.530 74.700 ;
        RECT 79.580 74.100 83.530 74.250 ;
        RECT 83.130 73.650 83.530 74.100 ;
        RECT 79.580 73.500 83.530 73.650 ;
        RECT 83.130 73.050 83.530 73.500 ;
        RECT 79.580 72.900 83.530 73.050 ;
        RECT 83.130 72.450 83.530 72.900 ;
        RECT 79.580 72.300 83.530 72.450 ;
        RECT 83.130 71.850 83.530 72.300 ;
        RECT 79.580 71.700 83.530 71.850 ;
        RECT 83.130 71.250 83.530 71.700 ;
        RECT 79.580 71.100 83.530 71.250 ;
        RECT 83.130 70.650 83.530 71.100 ;
        RECT 79.580 70.500 83.530 70.650 ;
        RECT 83.130 70.200 83.530 70.500 ;
        RECT 75.230 69.800 83.530 70.200 ;
        RECT 75.230 61.600 75.380 69.800 ;
        RECT 75.830 61.600 75.980 69.800 ;
        RECT 76.430 61.600 76.580 69.800 ;
        RECT 77.030 61.600 77.180 69.800 ;
        RECT 77.630 61.600 77.780 69.800 ;
        RECT 78.230 61.600 78.380 69.800 ;
        RECT 78.830 61.600 78.980 69.800 ;
        RECT 83.130 69.500 83.530 69.800 ;
        RECT 79.580 69.350 83.530 69.500 ;
        RECT 83.130 68.900 83.530 69.350 ;
        RECT 79.580 68.750 83.530 68.900 ;
        RECT 83.130 68.300 83.530 68.750 ;
        RECT 79.580 68.150 83.530 68.300 ;
        RECT 83.130 67.700 83.530 68.150 ;
        RECT 79.580 67.550 83.530 67.700 ;
        RECT 83.130 67.100 83.530 67.550 ;
        RECT 79.580 66.950 83.530 67.100 ;
        RECT 83.130 66.500 83.530 66.950 ;
        RECT 79.580 66.350 83.530 66.500 ;
        RECT 83.130 65.900 83.530 66.350 ;
        RECT 79.580 65.750 83.530 65.900 ;
        RECT 83.130 65.300 83.530 65.750 ;
        RECT 79.580 65.150 83.530 65.300 ;
        RECT 83.130 64.700 83.530 65.150 ;
        RECT 79.580 64.550 83.530 64.700 ;
        RECT 83.130 64.400 83.530 64.550 ;
        RECT 85.930 75.450 86.330 75.600 ;
        RECT 85.930 75.300 89.880 75.450 ;
        RECT 85.930 74.850 86.330 75.300 ;
        RECT 85.930 74.700 89.880 74.850 ;
        RECT 85.930 74.250 86.330 74.700 ;
        RECT 85.930 74.100 89.880 74.250 ;
        RECT 85.930 73.650 86.330 74.100 ;
        RECT 85.930 73.500 89.880 73.650 ;
        RECT 85.930 73.050 86.330 73.500 ;
        RECT 85.930 72.900 89.880 73.050 ;
        RECT 85.930 72.450 86.330 72.900 ;
        RECT 85.930 72.300 89.880 72.450 ;
        RECT 85.930 71.850 86.330 72.300 ;
        RECT 85.930 71.700 89.880 71.850 ;
        RECT 85.930 71.250 86.330 71.700 ;
        RECT 85.930 71.100 89.880 71.250 ;
        RECT 85.930 70.650 86.330 71.100 ;
        RECT 85.930 70.500 89.880 70.650 ;
        RECT 85.930 70.200 86.330 70.500 ;
        RECT 90.480 70.200 90.630 78.400 ;
        RECT 91.080 70.200 91.230 78.400 ;
        RECT 91.680 70.200 91.830 78.400 ;
        RECT 92.280 70.200 92.430 78.400 ;
        RECT 92.880 70.200 93.030 78.400 ;
        RECT 93.480 70.200 93.630 78.400 ;
        RECT 94.080 70.200 94.230 78.400 ;
        RECT 85.930 69.800 94.230 70.200 ;
        RECT 85.930 69.500 86.330 69.800 ;
        RECT 85.930 69.350 89.880 69.500 ;
        RECT 85.930 68.900 86.330 69.350 ;
        RECT 85.930 68.750 89.880 68.900 ;
        RECT 85.930 68.300 86.330 68.750 ;
        RECT 85.930 68.150 89.880 68.300 ;
        RECT 85.930 67.700 86.330 68.150 ;
        RECT 85.930 67.550 89.880 67.700 ;
        RECT 85.930 67.100 86.330 67.550 ;
        RECT 85.930 66.950 89.880 67.100 ;
        RECT 85.930 66.500 86.330 66.950 ;
        RECT 85.930 66.350 89.880 66.500 ;
        RECT 85.930 65.900 86.330 66.350 ;
        RECT 85.930 65.750 89.880 65.900 ;
        RECT 85.930 65.300 86.330 65.750 ;
        RECT 85.930 65.150 89.880 65.300 ;
        RECT 85.930 64.700 86.330 65.150 ;
        RECT 85.930 64.550 89.880 64.700 ;
        RECT 85.930 64.400 86.330 64.550 ;
        RECT 83.130 64.100 86.330 64.400 ;
        RECT 79.580 63.950 89.880 64.100 ;
        RECT 83.130 63.500 86.330 63.950 ;
        RECT 79.580 63.350 89.880 63.500 ;
        RECT 83.130 62.900 86.330 63.350 ;
        RECT 79.580 62.750 89.880 62.900 ;
        RECT 83.130 62.300 86.330 62.750 ;
        RECT 79.580 62.150 89.880 62.300 ;
        RECT 83.530 61.200 85.930 62.150 ;
        RECT 90.480 61.600 90.630 69.800 ;
        RECT 91.080 61.600 91.230 69.800 ;
        RECT 91.680 61.600 91.830 69.800 ;
        RECT 92.280 61.600 92.430 69.800 ;
        RECT 92.880 61.600 93.030 69.800 ;
        RECT 93.480 61.600 93.630 69.800 ;
        RECT 94.080 61.600 94.230 69.800 ;
        RECT 95.230 70.200 95.380 78.400 ;
        RECT 95.830 70.200 95.980 78.400 ;
        RECT 96.430 70.200 96.580 78.400 ;
        RECT 97.030 70.200 97.180 78.400 ;
        RECT 97.630 70.200 97.780 78.400 ;
        RECT 98.230 70.200 98.380 78.400 ;
        RECT 98.830 70.200 98.980 78.400 ;
        RECT 103.530 77.850 104.730 78.800 ;
        RECT 99.580 77.700 104.730 77.850 ;
        RECT 103.130 77.250 104.730 77.700 ;
        RECT 99.580 77.100 104.730 77.250 ;
        RECT 103.130 76.650 104.730 77.100 ;
        RECT 99.580 76.500 104.730 76.650 ;
        RECT 103.130 76.050 104.730 76.500 ;
        RECT 99.580 75.900 104.730 76.050 ;
        RECT 105.135 76.035 107.135 77.310 ;
        RECT 103.130 75.600 104.730 75.900 ;
        RECT 103.130 75.450 103.530 75.600 ;
        RECT 99.580 75.300 103.530 75.450 ;
        RECT 103.130 74.850 103.530 75.300 ;
        RECT 99.580 74.700 103.530 74.850 ;
        RECT 103.130 74.250 103.530 74.700 ;
        RECT 99.580 74.100 103.530 74.250 ;
        RECT 103.130 73.650 103.530 74.100 ;
        RECT 99.580 73.500 103.530 73.650 ;
        RECT 103.130 73.050 103.530 73.500 ;
        RECT 99.580 72.900 103.530 73.050 ;
        RECT 103.130 72.450 103.530 72.900 ;
        RECT 99.580 72.300 103.530 72.450 ;
        RECT 103.130 71.850 103.530 72.300 ;
        RECT 99.580 71.700 103.530 71.850 ;
        RECT 103.130 71.250 103.530 71.700 ;
        RECT 99.580 71.100 103.530 71.250 ;
        RECT 103.130 70.650 103.530 71.100 ;
        RECT 99.580 70.500 103.530 70.650 ;
        RECT 103.130 70.200 103.530 70.500 ;
        RECT 95.230 69.800 103.530 70.200 ;
        RECT 95.230 61.600 95.380 69.800 ;
        RECT 95.830 61.600 95.980 69.800 ;
        RECT 96.430 61.600 96.580 69.800 ;
        RECT 97.030 61.600 97.180 69.800 ;
        RECT 97.630 61.600 97.780 69.800 ;
        RECT 98.230 61.600 98.380 69.800 ;
        RECT 98.830 61.600 98.980 69.800 ;
        RECT 103.130 69.500 103.530 69.800 ;
        RECT 99.580 69.350 103.530 69.500 ;
        RECT 103.130 68.900 103.530 69.350 ;
        RECT 99.580 68.750 103.530 68.900 ;
        RECT 103.130 68.300 103.530 68.750 ;
        RECT 99.580 68.150 103.530 68.300 ;
        RECT 103.130 67.700 103.530 68.150 ;
        RECT 99.580 67.550 103.530 67.700 ;
        RECT 103.130 67.100 103.530 67.550 ;
        RECT 99.580 66.950 103.530 67.100 ;
        RECT 103.130 66.500 103.530 66.950 ;
        RECT 99.580 66.350 103.530 66.500 ;
        RECT 103.130 65.900 103.530 66.350 ;
        RECT 99.580 65.750 103.530 65.900 ;
        RECT 103.130 65.300 103.530 65.750 ;
        RECT 99.580 65.150 103.530 65.300 ;
        RECT 103.130 64.700 103.530 65.150 ;
        RECT 99.580 64.550 103.530 64.700 ;
        RECT 103.130 64.400 103.530 64.550 ;
        RECT 103.130 64.100 104.730 64.400 ;
        RECT 99.580 63.950 104.730 64.100 ;
        RECT 103.130 63.500 104.730 63.950 ;
        RECT 99.580 63.350 104.730 63.500 ;
        RECT 103.130 62.900 104.730 63.350 ;
        RECT 99.580 62.750 104.730 62.900 ;
        RECT 103.130 62.300 104.730 62.750 ;
        RECT 99.580 62.150 104.730 62.300 ;
        RECT 103.530 61.200 104.730 62.150 ;
        RECT 105.140 61.820 107.140 63.095 ;
        RECT 4.730 58.800 9.130 61.200 ;
        RECT 20.330 58.800 29.130 61.200 ;
        RECT 40.330 58.800 49.130 61.200 ;
        RECT 60.330 58.800 69.130 61.200 ;
        RECT 80.330 58.800 89.130 61.200 ;
        RECT 100.330 58.800 104.730 61.200 ;
        RECT 4.730 57.850 5.940 58.800 ;
        RECT 4.730 57.700 9.880 57.850 ;
        RECT 2.315 56.345 4.320 57.620 ;
        RECT 4.730 57.250 6.330 57.700 ;
        RECT 4.730 57.100 9.880 57.250 ;
        RECT 4.730 56.650 6.330 57.100 ;
        RECT 4.730 56.500 9.880 56.650 ;
        RECT 4.730 56.050 6.330 56.500 ;
        RECT 4.730 55.900 9.880 56.050 ;
        RECT 4.730 55.600 6.330 55.900 ;
        RECT 2.315 53.255 4.315 55.550 ;
        RECT 5.930 55.450 6.330 55.600 ;
        RECT 5.930 55.300 9.880 55.450 ;
        RECT 5.930 54.850 6.330 55.300 ;
        RECT 5.930 54.700 9.880 54.850 ;
        RECT 5.930 54.250 6.330 54.700 ;
        RECT 5.930 54.100 9.880 54.250 ;
        RECT 5.930 53.650 6.330 54.100 ;
        RECT 5.930 53.500 9.880 53.650 ;
        RECT 5.930 53.050 6.330 53.500 ;
        RECT 5.930 52.900 9.880 53.050 ;
        RECT 5.930 52.450 6.330 52.900 ;
        RECT 5.930 52.300 9.880 52.450 ;
        RECT 5.930 51.850 6.330 52.300 ;
        RECT 5.930 51.700 9.880 51.850 ;
        RECT 5.930 51.250 6.330 51.700 ;
        RECT 5.930 51.100 9.880 51.250 ;
        RECT 5.930 50.650 6.330 51.100 ;
        RECT 5.930 50.500 9.880 50.650 ;
        RECT 5.930 50.200 6.330 50.500 ;
        RECT 10.480 50.200 10.630 58.400 ;
        RECT 11.080 50.200 11.230 58.400 ;
        RECT 11.680 50.200 11.830 58.400 ;
        RECT 12.280 50.200 12.430 58.400 ;
        RECT 12.880 50.200 13.030 58.400 ;
        RECT 13.480 50.200 13.630 58.400 ;
        RECT 14.080 50.200 14.230 58.400 ;
        RECT 5.930 49.800 14.230 50.200 ;
        RECT 5.930 49.500 6.330 49.800 ;
        RECT 5.930 49.350 9.880 49.500 ;
        RECT 5.930 48.900 6.330 49.350 ;
        RECT 5.930 48.750 9.880 48.900 ;
        RECT 5.930 48.300 6.330 48.750 ;
        RECT 5.930 48.150 9.880 48.300 ;
        RECT 5.930 47.700 6.330 48.150 ;
        RECT 5.930 47.550 9.880 47.700 ;
        RECT 5.930 47.100 6.330 47.550 ;
        RECT 5.930 46.950 9.880 47.100 ;
        RECT 2.315 44.445 4.315 46.740 ;
        RECT 5.930 46.500 6.330 46.950 ;
        RECT 5.930 46.350 9.880 46.500 ;
        RECT 5.930 45.900 6.330 46.350 ;
        RECT 5.930 45.750 9.880 45.900 ;
        RECT 5.930 45.300 6.330 45.750 ;
        RECT 5.930 45.150 9.880 45.300 ;
        RECT 5.930 44.700 6.330 45.150 ;
        RECT 5.930 44.550 9.880 44.700 ;
        RECT 5.930 44.400 6.330 44.550 ;
        RECT 4.730 44.100 6.330 44.400 ;
        RECT 4.730 43.950 9.880 44.100 ;
        RECT 4.730 43.500 6.330 43.950 ;
        RECT 4.730 43.350 9.880 43.500 ;
        RECT 2.315 42.045 4.315 43.320 ;
        RECT 4.730 42.900 6.330 43.350 ;
        RECT 4.730 42.750 9.880 42.900 ;
        RECT 4.730 42.300 6.330 42.750 ;
        RECT 4.730 42.150 9.880 42.300 ;
        RECT 4.730 41.200 5.930 42.150 ;
        RECT 10.480 41.600 10.630 49.800 ;
        RECT 11.080 41.600 11.230 49.800 ;
        RECT 11.680 41.600 11.830 49.800 ;
        RECT 12.280 41.600 12.430 49.800 ;
        RECT 12.880 41.600 13.030 49.800 ;
        RECT 13.480 41.600 13.630 49.800 ;
        RECT 14.080 41.600 14.230 49.800 ;
        RECT 15.230 50.200 15.380 58.400 ;
        RECT 15.830 50.200 15.980 58.400 ;
        RECT 16.430 50.200 16.580 58.400 ;
        RECT 17.030 50.200 17.180 58.400 ;
        RECT 17.630 50.200 17.780 58.400 ;
        RECT 18.230 50.200 18.380 58.400 ;
        RECT 18.830 50.200 18.980 58.400 ;
        RECT 23.530 57.850 25.940 58.800 ;
        RECT 19.580 57.700 29.880 57.850 ;
        RECT 23.130 57.250 26.330 57.700 ;
        RECT 19.580 57.100 29.880 57.250 ;
        RECT 23.130 56.650 26.330 57.100 ;
        RECT 19.580 56.500 29.880 56.650 ;
        RECT 23.130 56.050 26.330 56.500 ;
        RECT 19.580 55.900 29.880 56.050 ;
        RECT 23.130 55.600 26.330 55.900 ;
        RECT 23.130 55.450 23.530 55.600 ;
        RECT 19.580 55.300 23.530 55.450 ;
        RECT 23.130 54.850 23.530 55.300 ;
        RECT 19.580 54.700 23.530 54.850 ;
        RECT 23.130 54.250 23.530 54.700 ;
        RECT 19.580 54.100 23.530 54.250 ;
        RECT 23.130 53.650 23.530 54.100 ;
        RECT 19.580 53.500 23.530 53.650 ;
        RECT 23.130 53.050 23.530 53.500 ;
        RECT 19.580 52.900 23.530 53.050 ;
        RECT 23.130 52.450 23.530 52.900 ;
        RECT 19.580 52.300 23.530 52.450 ;
        RECT 23.130 51.850 23.530 52.300 ;
        RECT 19.580 51.700 23.530 51.850 ;
        RECT 23.130 51.250 23.530 51.700 ;
        RECT 19.580 51.100 23.530 51.250 ;
        RECT 23.130 50.650 23.530 51.100 ;
        RECT 19.580 50.500 23.530 50.650 ;
        RECT 23.130 50.200 23.530 50.500 ;
        RECT 15.230 49.800 23.530 50.200 ;
        RECT 15.230 41.600 15.380 49.800 ;
        RECT 15.830 41.600 15.980 49.800 ;
        RECT 16.430 41.600 16.580 49.800 ;
        RECT 17.030 41.600 17.180 49.800 ;
        RECT 17.630 41.600 17.780 49.800 ;
        RECT 18.230 41.600 18.380 49.800 ;
        RECT 18.830 41.600 18.980 49.800 ;
        RECT 23.130 49.500 23.530 49.800 ;
        RECT 19.580 49.350 23.530 49.500 ;
        RECT 23.130 48.900 23.530 49.350 ;
        RECT 19.580 48.750 23.530 48.900 ;
        RECT 23.130 48.300 23.530 48.750 ;
        RECT 19.580 48.150 23.530 48.300 ;
        RECT 23.130 47.700 23.530 48.150 ;
        RECT 19.580 47.550 23.530 47.700 ;
        RECT 23.130 47.100 23.530 47.550 ;
        RECT 19.580 46.950 23.530 47.100 ;
        RECT 23.130 46.500 23.530 46.950 ;
        RECT 19.580 46.350 23.530 46.500 ;
        RECT 23.130 45.900 23.530 46.350 ;
        RECT 19.580 45.750 23.530 45.900 ;
        RECT 23.130 45.300 23.530 45.750 ;
        RECT 19.580 45.150 23.530 45.300 ;
        RECT 23.130 44.700 23.530 45.150 ;
        RECT 19.580 44.550 23.530 44.700 ;
        RECT 23.130 44.400 23.530 44.550 ;
        RECT 25.930 55.450 26.330 55.600 ;
        RECT 25.930 55.300 29.880 55.450 ;
        RECT 25.930 54.850 26.330 55.300 ;
        RECT 25.930 54.700 29.880 54.850 ;
        RECT 25.930 54.250 26.330 54.700 ;
        RECT 25.930 54.100 29.880 54.250 ;
        RECT 25.930 53.650 26.330 54.100 ;
        RECT 25.930 53.500 29.880 53.650 ;
        RECT 25.930 53.050 26.330 53.500 ;
        RECT 25.930 52.900 29.880 53.050 ;
        RECT 25.930 52.450 26.330 52.900 ;
        RECT 25.930 52.300 29.880 52.450 ;
        RECT 25.930 51.850 26.330 52.300 ;
        RECT 25.930 51.700 29.880 51.850 ;
        RECT 25.930 51.250 26.330 51.700 ;
        RECT 25.930 51.100 29.880 51.250 ;
        RECT 25.930 50.650 26.330 51.100 ;
        RECT 25.930 50.500 29.880 50.650 ;
        RECT 25.930 50.200 26.330 50.500 ;
        RECT 30.480 50.200 30.630 58.400 ;
        RECT 31.080 50.200 31.230 58.400 ;
        RECT 31.680 50.200 31.830 58.400 ;
        RECT 32.280 50.200 32.430 58.400 ;
        RECT 32.880 50.200 33.030 58.400 ;
        RECT 33.480 50.200 33.630 58.400 ;
        RECT 34.080 50.200 34.230 58.400 ;
        RECT 25.930 49.800 34.230 50.200 ;
        RECT 25.930 49.500 26.330 49.800 ;
        RECT 25.930 49.350 29.880 49.500 ;
        RECT 25.930 48.900 26.330 49.350 ;
        RECT 25.930 48.750 29.880 48.900 ;
        RECT 25.930 48.300 26.330 48.750 ;
        RECT 25.930 48.150 29.880 48.300 ;
        RECT 25.930 47.700 26.330 48.150 ;
        RECT 25.930 47.550 29.880 47.700 ;
        RECT 25.930 47.100 26.330 47.550 ;
        RECT 25.930 46.950 29.880 47.100 ;
        RECT 25.930 46.500 26.330 46.950 ;
        RECT 25.930 46.350 29.880 46.500 ;
        RECT 25.930 45.900 26.330 46.350 ;
        RECT 25.930 45.750 29.880 45.900 ;
        RECT 25.930 45.300 26.330 45.750 ;
        RECT 25.930 45.150 29.880 45.300 ;
        RECT 25.930 44.700 26.330 45.150 ;
        RECT 25.930 44.550 29.880 44.700 ;
        RECT 25.930 44.400 26.330 44.550 ;
        RECT 23.130 44.100 26.330 44.400 ;
        RECT 19.580 43.950 29.880 44.100 ;
        RECT 23.130 43.500 26.330 43.950 ;
        RECT 19.580 43.350 29.880 43.500 ;
        RECT 23.130 42.900 26.330 43.350 ;
        RECT 19.580 42.750 29.880 42.900 ;
        RECT 23.130 42.300 26.330 42.750 ;
        RECT 19.580 42.150 29.880 42.300 ;
        RECT 23.530 41.200 25.930 42.150 ;
        RECT 30.480 41.600 30.630 49.800 ;
        RECT 31.080 41.600 31.230 49.800 ;
        RECT 31.680 41.600 31.830 49.800 ;
        RECT 32.280 41.600 32.430 49.800 ;
        RECT 32.880 41.600 33.030 49.800 ;
        RECT 33.480 41.600 33.630 49.800 ;
        RECT 34.080 41.600 34.230 49.800 ;
        RECT 35.230 50.200 35.380 58.400 ;
        RECT 35.830 50.200 35.980 58.400 ;
        RECT 36.430 50.200 36.580 58.400 ;
        RECT 37.030 50.200 37.180 58.400 ;
        RECT 37.630 50.200 37.780 58.400 ;
        RECT 38.230 50.200 38.380 58.400 ;
        RECT 38.830 50.200 38.980 58.400 ;
        RECT 43.530 57.850 45.940 58.800 ;
        RECT 39.580 57.700 49.880 57.850 ;
        RECT 43.130 57.250 46.330 57.700 ;
        RECT 39.580 57.100 49.880 57.250 ;
        RECT 43.130 56.650 46.330 57.100 ;
        RECT 39.580 56.500 49.880 56.650 ;
        RECT 43.130 56.050 46.330 56.500 ;
        RECT 39.580 55.900 49.880 56.050 ;
        RECT 43.130 55.600 46.330 55.900 ;
        RECT 43.130 55.450 43.530 55.600 ;
        RECT 39.580 55.300 43.530 55.450 ;
        RECT 43.130 54.850 43.530 55.300 ;
        RECT 39.580 54.700 43.530 54.850 ;
        RECT 43.130 54.250 43.530 54.700 ;
        RECT 39.580 54.100 43.530 54.250 ;
        RECT 43.130 53.650 43.530 54.100 ;
        RECT 39.580 53.500 43.530 53.650 ;
        RECT 43.130 53.050 43.530 53.500 ;
        RECT 39.580 52.900 43.530 53.050 ;
        RECT 43.130 52.450 43.530 52.900 ;
        RECT 39.580 52.300 43.530 52.450 ;
        RECT 43.130 51.850 43.530 52.300 ;
        RECT 39.580 51.700 43.530 51.850 ;
        RECT 43.130 51.250 43.530 51.700 ;
        RECT 39.580 51.100 43.530 51.250 ;
        RECT 43.130 50.650 43.530 51.100 ;
        RECT 39.580 50.500 43.530 50.650 ;
        RECT 43.130 50.200 43.530 50.500 ;
        RECT 35.230 49.800 43.530 50.200 ;
        RECT 35.230 41.600 35.380 49.800 ;
        RECT 35.830 41.600 35.980 49.800 ;
        RECT 36.430 41.600 36.580 49.800 ;
        RECT 37.030 41.600 37.180 49.800 ;
        RECT 37.630 41.600 37.780 49.800 ;
        RECT 38.230 41.600 38.380 49.800 ;
        RECT 38.830 41.600 38.980 49.800 ;
        RECT 43.130 49.500 43.530 49.800 ;
        RECT 39.580 49.350 43.530 49.500 ;
        RECT 43.130 48.900 43.530 49.350 ;
        RECT 39.580 48.750 43.530 48.900 ;
        RECT 43.130 48.300 43.530 48.750 ;
        RECT 39.580 48.150 43.530 48.300 ;
        RECT 43.130 47.700 43.530 48.150 ;
        RECT 39.580 47.550 43.530 47.700 ;
        RECT 43.130 47.100 43.530 47.550 ;
        RECT 39.580 46.950 43.530 47.100 ;
        RECT 43.130 46.500 43.530 46.950 ;
        RECT 39.580 46.350 43.530 46.500 ;
        RECT 43.130 45.900 43.530 46.350 ;
        RECT 39.580 45.750 43.530 45.900 ;
        RECT 43.130 45.300 43.530 45.750 ;
        RECT 39.580 45.150 43.530 45.300 ;
        RECT 43.130 44.700 43.530 45.150 ;
        RECT 39.580 44.550 43.530 44.700 ;
        RECT 43.130 44.400 43.530 44.550 ;
        RECT 45.930 55.450 46.330 55.600 ;
        RECT 45.930 55.300 49.880 55.450 ;
        RECT 45.930 54.850 46.330 55.300 ;
        RECT 45.930 54.700 49.880 54.850 ;
        RECT 45.930 54.250 46.330 54.700 ;
        RECT 45.930 54.100 49.880 54.250 ;
        RECT 45.930 53.650 46.330 54.100 ;
        RECT 45.930 53.500 49.880 53.650 ;
        RECT 45.930 53.050 46.330 53.500 ;
        RECT 45.930 52.900 49.880 53.050 ;
        RECT 45.930 52.450 46.330 52.900 ;
        RECT 45.930 52.300 49.880 52.450 ;
        RECT 45.930 51.850 46.330 52.300 ;
        RECT 45.930 51.700 49.880 51.850 ;
        RECT 45.930 51.250 46.330 51.700 ;
        RECT 45.930 51.100 49.880 51.250 ;
        RECT 45.930 50.650 46.330 51.100 ;
        RECT 45.930 50.500 49.880 50.650 ;
        RECT 45.930 50.200 46.330 50.500 ;
        RECT 50.480 50.200 50.630 58.400 ;
        RECT 51.080 50.200 51.230 58.400 ;
        RECT 51.680 50.200 51.830 58.400 ;
        RECT 52.280 50.200 52.430 58.400 ;
        RECT 52.880 50.200 53.030 58.400 ;
        RECT 53.480 50.200 53.630 58.400 ;
        RECT 54.080 50.200 54.230 58.400 ;
        RECT 45.930 49.800 54.230 50.200 ;
        RECT 45.930 49.500 46.330 49.800 ;
        RECT 45.930 49.350 49.880 49.500 ;
        RECT 45.930 48.900 46.330 49.350 ;
        RECT 45.930 48.750 49.880 48.900 ;
        RECT 45.930 48.300 46.330 48.750 ;
        RECT 45.930 48.150 49.880 48.300 ;
        RECT 45.930 47.700 46.330 48.150 ;
        RECT 45.930 47.550 49.880 47.700 ;
        RECT 45.930 47.100 46.330 47.550 ;
        RECT 45.930 46.950 49.880 47.100 ;
        RECT 45.930 46.500 46.330 46.950 ;
        RECT 45.930 46.350 49.880 46.500 ;
        RECT 45.930 45.900 46.330 46.350 ;
        RECT 45.930 45.750 49.880 45.900 ;
        RECT 45.930 45.300 46.330 45.750 ;
        RECT 45.930 45.150 49.880 45.300 ;
        RECT 45.930 44.700 46.330 45.150 ;
        RECT 45.930 44.550 49.880 44.700 ;
        RECT 45.930 44.400 46.330 44.550 ;
        RECT 43.130 44.100 46.330 44.400 ;
        RECT 39.580 43.950 49.880 44.100 ;
        RECT 43.130 43.500 46.330 43.950 ;
        RECT 39.580 43.350 49.880 43.500 ;
        RECT 43.130 42.900 46.330 43.350 ;
        RECT 39.580 42.750 49.880 42.900 ;
        RECT 43.130 42.300 46.330 42.750 ;
        RECT 39.580 42.150 49.880 42.300 ;
        RECT 43.530 41.200 45.930 42.150 ;
        RECT 50.480 41.600 50.630 49.800 ;
        RECT 51.080 41.600 51.230 49.800 ;
        RECT 51.680 41.600 51.830 49.800 ;
        RECT 52.280 41.600 52.430 49.800 ;
        RECT 52.880 41.600 53.030 49.800 ;
        RECT 53.480 41.600 53.630 49.800 ;
        RECT 54.080 41.600 54.230 49.800 ;
        RECT 55.230 50.200 55.380 58.400 ;
        RECT 55.830 50.200 55.980 58.400 ;
        RECT 56.430 50.200 56.580 58.400 ;
        RECT 57.030 50.200 57.180 58.400 ;
        RECT 57.630 50.200 57.780 58.400 ;
        RECT 58.230 50.200 58.380 58.400 ;
        RECT 58.830 50.200 58.980 58.400 ;
        RECT 63.530 57.850 65.940 58.800 ;
        RECT 59.580 57.700 69.880 57.850 ;
        RECT 63.130 57.250 66.330 57.700 ;
        RECT 59.580 57.100 69.880 57.250 ;
        RECT 63.130 56.650 66.330 57.100 ;
        RECT 59.580 56.500 69.880 56.650 ;
        RECT 63.130 56.050 66.330 56.500 ;
        RECT 59.580 55.900 69.880 56.050 ;
        RECT 63.130 55.600 66.330 55.900 ;
        RECT 63.130 55.450 63.530 55.600 ;
        RECT 59.580 55.300 63.530 55.450 ;
        RECT 63.130 54.850 63.530 55.300 ;
        RECT 59.580 54.700 63.530 54.850 ;
        RECT 63.130 54.250 63.530 54.700 ;
        RECT 59.580 54.100 63.530 54.250 ;
        RECT 63.130 53.650 63.530 54.100 ;
        RECT 59.580 53.500 63.530 53.650 ;
        RECT 63.130 53.050 63.530 53.500 ;
        RECT 59.580 52.900 63.530 53.050 ;
        RECT 63.130 52.450 63.530 52.900 ;
        RECT 59.580 52.300 63.530 52.450 ;
        RECT 63.130 51.850 63.530 52.300 ;
        RECT 59.580 51.700 63.530 51.850 ;
        RECT 63.130 51.250 63.530 51.700 ;
        RECT 59.580 51.100 63.530 51.250 ;
        RECT 63.130 50.650 63.530 51.100 ;
        RECT 59.580 50.500 63.530 50.650 ;
        RECT 63.130 50.200 63.530 50.500 ;
        RECT 55.230 49.800 63.530 50.200 ;
        RECT 55.230 41.600 55.380 49.800 ;
        RECT 55.830 41.600 55.980 49.800 ;
        RECT 56.430 41.600 56.580 49.800 ;
        RECT 57.030 41.600 57.180 49.800 ;
        RECT 57.630 41.600 57.780 49.800 ;
        RECT 58.230 41.600 58.380 49.800 ;
        RECT 58.830 41.600 58.980 49.800 ;
        RECT 63.130 49.500 63.530 49.800 ;
        RECT 59.580 49.350 63.530 49.500 ;
        RECT 63.130 48.900 63.530 49.350 ;
        RECT 59.580 48.750 63.530 48.900 ;
        RECT 63.130 48.300 63.530 48.750 ;
        RECT 59.580 48.150 63.530 48.300 ;
        RECT 63.130 47.700 63.530 48.150 ;
        RECT 59.580 47.550 63.530 47.700 ;
        RECT 63.130 47.100 63.530 47.550 ;
        RECT 59.580 46.950 63.530 47.100 ;
        RECT 63.130 46.500 63.530 46.950 ;
        RECT 59.580 46.350 63.530 46.500 ;
        RECT 63.130 45.900 63.530 46.350 ;
        RECT 59.580 45.750 63.530 45.900 ;
        RECT 63.130 45.300 63.530 45.750 ;
        RECT 59.580 45.150 63.530 45.300 ;
        RECT 63.130 44.700 63.530 45.150 ;
        RECT 59.580 44.550 63.530 44.700 ;
        RECT 63.130 44.400 63.530 44.550 ;
        RECT 65.930 55.450 66.330 55.600 ;
        RECT 65.930 55.300 69.880 55.450 ;
        RECT 65.930 54.850 66.330 55.300 ;
        RECT 65.930 54.700 69.880 54.850 ;
        RECT 65.930 54.250 66.330 54.700 ;
        RECT 65.930 54.100 69.880 54.250 ;
        RECT 65.930 53.650 66.330 54.100 ;
        RECT 65.930 53.500 69.880 53.650 ;
        RECT 65.930 53.050 66.330 53.500 ;
        RECT 65.930 52.900 69.880 53.050 ;
        RECT 65.930 52.450 66.330 52.900 ;
        RECT 65.930 52.300 69.880 52.450 ;
        RECT 65.930 51.850 66.330 52.300 ;
        RECT 65.930 51.700 69.880 51.850 ;
        RECT 65.930 51.250 66.330 51.700 ;
        RECT 65.930 51.100 69.880 51.250 ;
        RECT 65.930 50.650 66.330 51.100 ;
        RECT 65.930 50.500 69.880 50.650 ;
        RECT 65.930 50.200 66.330 50.500 ;
        RECT 70.480 50.200 70.630 58.400 ;
        RECT 71.080 50.200 71.230 58.400 ;
        RECT 71.680 50.200 71.830 58.400 ;
        RECT 72.280 50.200 72.430 58.400 ;
        RECT 72.880 50.200 73.030 58.400 ;
        RECT 73.480 50.200 73.630 58.400 ;
        RECT 74.080 50.200 74.230 58.400 ;
        RECT 65.930 49.800 74.230 50.200 ;
        RECT 65.930 49.500 66.330 49.800 ;
        RECT 65.930 49.350 69.880 49.500 ;
        RECT 65.930 48.900 66.330 49.350 ;
        RECT 65.930 48.750 69.880 48.900 ;
        RECT 65.930 48.300 66.330 48.750 ;
        RECT 65.930 48.150 69.880 48.300 ;
        RECT 65.930 47.700 66.330 48.150 ;
        RECT 65.930 47.550 69.880 47.700 ;
        RECT 65.930 47.100 66.330 47.550 ;
        RECT 65.930 46.950 69.880 47.100 ;
        RECT 65.930 46.500 66.330 46.950 ;
        RECT 65.930 46.350 69.880 46.500 ;
        RECT 65.930 45.900 66.330 46.350 ;
        RECT 65.930 45.750 69.880 45.900 ;
        RECT 65.930 45.300 66.330 45.750 ;
        RECT 65.930 45.150 69.880 45.300 ;
        RECT 65.930 44.700 66.330 45.150 ;
        RECT 65.930 44.550 69.880 44.700 ;
        RECT 65.930 44.400 66.330 44.550 ;
        RECT 63.130 44.100 66.330 44.400 ;
        RECT 59.580 43.950 69.880 44.100 ;
        RECT 63.130 43.500 66.330 43.950 ;
        RECT 59.580 43.350 69.880 43.500 ;
        RECT 63.130 42.900 66.330 43.350 ;
        RECT 59.580 42.750 69.880 42.900 ;
        RECT 63.130 42.300 66.330 42.750 ;
        RECT 59.580 42.150 69.880 42.300 ;
        RECT 63.530 41.200 65.930 42.150 ;
        RECT 70.480 41.600 70.630 49.800 ;
        RECT 71.080 41.600 71.230 49.800 ;
        RECT 71.680 41.600 71.830 49.800 ;
        RECT 72.280 41.600 72.430 49.800 ;
        RECT 72.880 41.600 73.030 49.800 ;
        RECT 73.480 41.600 73.630 49.800 ;
        RECT 74.080 41.600 74.230 49.800 ;
        RECT 75.230 50.200 75.380 58.400 ;
        RECT 75.830 50.200 75.980 58.400 ;
        RECT 76.430 50.200 76.580 58.400 ;
        RECT 77.030 50.200 77.180 58.400 ;
        RECT 77.630 50.200 77.780 58.400 ;
        RECT 78.230 50.200 78.380 58.400 ;
        RECT 78.830 50.200 78.980 58.400 ;
        RECT 83.530 57.850 85.940 58.800 ;
        RECT 79.580 57.700 89.880 57.850 ;
        RECT 83.130 57.250 86.330 57.700 ;
        RECT 79.580 57.100 89.880 57.250 ;
        RECT 83.130 56.650 86.330 57.100 ;
        RECT 79.580 56.500 89.880 56.650 ;
        RECT 83.130 56.050 86.330 56.500 ;
        RECT 79.580 55.900 89.880 56.050 ;
        RECT 83.130 55.600 86.330 55.900 ;
        RECT 83.130 55.450 83.530 55.600 ;
        RECT 79.580 55.300 83.530 55.450 ;
        RECT 83.130 54.850 83.530 55.300 ;
        RECT 79.580 54.700 83.530 54.850 ;
        RECT 83.130 54.250 83.530 54.700 ;
        RECT 79.580 54.100 83.530 54.250 ;
        RECT 83.130 53.650 83.530 54.100 ;
        RECT 79.580 53.500 83.530 53.650 ;
        RECT 83.130 53.050 83.530 53.500 ;
        RECT 79.580 52.900 83.530 53.050 ;
        RECT 83.130 52.450 83.530 52.900 ;
        RECT 79.580 52.300 83.530 52.450 ;
        RECT 83.130 51.850 83.530 52.300 ;
        RECT 79.580 51.700 83.530 51.850 ;
        RECT 83.130 51.250 83.530 51.700 ;
        RECT 79.580 51.100 83.530 51.250 ;
        RECT 83.130 50.650 83.530 51.100 ;
        RECT 79.580 50.500 83.530 50.650 ;
        RECT 83.130 50.200 83.530 50.500 ;
        RECT 75.230 49.800 83.530 50.200 ;
        RECT 75.230 41.600 75.380 49.800 ;
        RECT 75.830 41.600 75.980 49.800 ;
        RECT 76.430 41.600 76.580 49.800 ;
        RECT 77.030 41.600 77.180 49.800 ;
        RECT 77.630 41.600 77.780 49.800 ;
        RECT 78.230 41.600 78.380 49.800 ;
        RECT 78.830 41.600 78.980 49.800 ;
        RECT 83.130 49.500 83.530 49.800 ;
        RECT 79.580 49.350 83.530 49.500 ;
        RECT 83.130 48.900 83.530 49.350 ;
        RECT 79.580 48.750 83.530 48.900 ;
        RECT 83.130 48.300 83.530 48.750 ;
        RECT 79.580 48.150 83.530 48.300 ;
        RECT 83.130 47.700 83.530 48.150 ;
        RECT 79.580 47.550 83.530 47.700 ;
        RECT 83.130 47.100 83.530 47.550 ;
        RECT 79.580 46.950 83.530 47.100 ;
        RECT 83.130 46.500 83.530 46.950 ;
        RECT 79.580 46.350 83.530 46.500 ;
        RECT 83.130 45.900 83.530 46.350 ;
        RECT 79.580 45.750 83.530 45.900 ;
        RECT 83.130 45.300 83.530 45.750 ;
        RECT 79.580 45.150 83.530 45.300 ;
        RECT 83.130 44.700 83.530 45.150 ;
        RECT 79.580 44.550 83.530 44.700 ;
        RECT 83.130 44.400 83.530 44.550 ;
        RECT 85.930 55.450 86.330 55.600 ;
        RECT 85.930 55.300 89.880 55.450 ;
        RECT 85.930 54.850 86.330 55.300 ;
        RECT 85.930 54.700 89.880 54.850 ;
        RECT 85.930 54.250 86.330 54.700 ;
        RECT 85.930 54.100 89.880 54.250 ;
        RECT 85.930 53.650 86.330 54.100 ;
        RECT 85.930 53.500 89.880 53.650 ;
        RECT 85.930 53.050 86.330 53.500 ;
        RECT 85.930 52.900 89.880 53.050 ;
        RECT 85.930 52.450 86.330 52.900 ;
        RECT 85.930 52.300 89.880 52.450 ;
        RECT 85.930 51.850 86.330 52.300 ;
        RECT 85.930 51.700 89.880 51.850 ;
        RECT 85.930 51.250 86.330 51.700 ;
        RECT 85.930 51.100 89.880 51.250 ;
        RECT 85.930 50.650 86.330 51.100 ;
        RECT 85.930 50.500 89.880 50.650 ;
        RECT 85.930 50.200 86.330 50.500 ;
        RECT 90.480 50.200 90.630 58.400 ;
        RECT 91.080 50.200 91.230 58.400 ;
        RECT 91.680 50.200 91.830 58.400 ;
        RECT 92.280 50.200 92.430 58.400 ;
        RECT 92.880 50.200 93.030 58.400 ;
        RECT 93.480 50.200 93.630 58.400 ;
        RECT 94.080 50.200 94.230 58.400 ;
        RECT 85.930 49.800 94.230 50.200 ;
        RECT 85.930 49.500 86.330 49.800 ;
        RECT 85.930 49.350 89.880 49.500 ;
        RECT 85.930 48.900 86.330 49.350 ;
        RECT 85.930 48.750 89.880 48.900 ;
        RECT 85.930 48.300 86.330 48.750 ;
        RECT 85.930 48.150 89.880 48.300 ;
        RECT 85.930 47.700 86.330 48.150 ;
        RECT 85.930 47.550 89.880 47.700 ;
        RECT 85.930 47.100 86.330 47.550 ;
        RECT 85.930 46.950 89.880 47.100 ;
        RECT 85.930 46.500 86.330 46.950 ;
        RECT 85.930 46.350 89.880 46.500 ;
        RECT 85.930 45.900 86.330 46.350 ;
        RECT 85.930 45.750 89.880 45.900 ;
        RECT 85.930 45.300 86.330 45.750 ;
        RECT 85.930 45.150 89.880 45.300 ;
        RECT 85.930 44.700 86.330 45.150 ;
        RECT 85.930 44.550 89.880 44.700 ;
        RECT 85.930 44.400 86.330 44.550 ;
        RECT 83.130 44.100 86.330 44.400 ;
        RECT 79.580 43.950 89.880 44.100 ;
        RECT 83.130 43.500 86.330 43.950 ;
        RECT 79.580 43.350 89.880 43.500 ;
        RECT 83.130 42.900 86.330 43.350 ;
        RECT 79.580 42.750 89.880 42.900 ;
        RECT 83.130 42.300 86.330 42.750 ;
        RECT 79.580 42.150 89.880 42.300 ;
        RECT 83.530 41.200 85.930 42.150 ;
        RECT 90.480 41.600 90.630 49.800 ;
        RECT 91.080 41.600 91.230 49.800 ;
        RECT 91.680 41.600 91.830 49.800 ;
        RECT 92.280 41.600 92.430 49.800 ;
        RECT 92.880 41.600 93.030 49.800 ;
        RECT 93.480 41.600 93.630 49.800 ;
        RECT 94.080 41.600 94.230 49.800 ;
        RECT 95.230 50.200 95.380 58.400 ;
        RECT 95.830 50.200 95.980 58.400 ;
        RECT 96.430 50.200 96.580 58.400 ;
        RECT 97.030 50.200 97.180 58.400 ;
        RECT 97.630 50.200 97.780 58.400 ;
        RECT 98.230 50.200 98.380 58.400 ;
        RECT 98.830 50.200 98.980 58.400 ;
        RECT 103.530 57.850 104.730 58.800 ;
        RECT 99.580 57.700 104.730 57.850 ;
        RECT 103.130 57.250 104.730 57.700 ;
        RECT 99.580 57.100 104.730 57.250 ;
        RECT 103.130 56.650 104.730 57.100 ;
        RECT 99.580 56.500 104.730 56.650 ;
        RECT 103.130 56.050 104.730 56.500 ;
        RECT 99.580 55.900 104.730 56.050 ;
        RECT 105.135 56.035 107.135 57.310 ;
        RECT 103.130 55.600 104.730 55.900 ;
        RECT 103.130 55.450 103.530 55.600 ;
        RECT 99.580 55.300 103.530 55.450 ;
        RECT 103.130 54.850 103.530 55.300 ;
        RECT 99.580 54.700 103.530 54.850 ;
        RECT 103.130 54.250 103.530 54.700 ;
        RECT 99.580 54.100 103.530 54.250 ;
        RECT 103.130 53.650 103.530 54.100 ;
        RECT 99.580 53.500 103.530 53.650 ;
        RECT 103.130 53.050 103.530 53.500 ;
        RECT 99.580 52.900 103.530 53.050 ;
        RECT 103.130 52.450 103.530 52.900 ;
        RECT 99.580 52.300 103.530 52.450 ;
        RECT 103.130 51.850 103.530 52.300 ;
        RECT 99.580 51.700 103.530 51.850 ;
        RECT 103.130 51.250 103.530 51.700 ;
        RECT 99.580 51.100 103.530 51.250 ;
        RECT 103.130 50.650 103.530 51.100 ;
        RECT 99.580 50.500 103.530 50.650 ;
        RECT 103.130 50.200 103.530 50.500 ;
        RECT 95.230 49.800 103.530 50.200 ;
        RECT 95.230 41.600 95.380 49.800 ;
        RECT 95.830 41.600 95.980 49.800 ;
        RECT 96.430 41.600 96.580 49.800 ;
        RECT 97.030 41.600 97.180 49.800 ;
        RECT 97.630 41.600 97.780 49.800 ;
        RECT 98.230 41.600 98.380 49.800 ;
        RECT 98.830 41.600 98.980 49.800 ;
        RECT 103.130 49.500 103.530 49.800 ;
        RECT 99.580 49.350 103.530 49.500 ;
        RECT 103.130 48.900 103.530 49.350 ;
        RECT 99.580 48.750 103.530 48.900 ;
        RECT 103.130 48.300 103.530 48.750 ;
        RECT 99.580 48.150 103.530 48.300 ;
        RECT 103.130 47.700 103.530 48.150 ;
        RECT 99.580 47.550 103.530 47.700 ;
        RECT 103.130 47.100 103.530 47.550 ;
        RECT 99.580 46.950 103.530 47.100 ;
        RECT 103.130 46.500 103.530 46.950 ;
        RECT 99.580 46.350 103.530 46.500 ;
        RECT 103.130 45.900 103.530 46.350 ;
        RECT 99.580 45.750 103.530 45.900 ;
        RECT 103.130 45.300 103.530 45.750 ;
        RECT 99.580 45.150 103.530 45.300 ;
        RECT 103.130 44.700 103.530 45.150 ;
        RECT 99.580 44.550 103.530 44.700 ;
        RECT 103.130 44.400 103.530 44.550 ;
        RECT 103.130 44.100 104.730 44.400 ;
        RECT 99.580 43.950 104.730 44.100 ;
        RECT 103.130 43.500 104.730 43.950 ;
        RECT 99.580 43.350 104.730 43.500 ;
        RECT 103.130 42.900 104.730 43.350 ;
        RECT 99.580 42.750 104.730 42.900 ;
        RECT 103.130 42.300 104.730 42.750 ;
        RECT 99.580 42.150 104.730 42.300 ;
        RECT 103.530 41.200 104.730 42.150 ;
        RECT 105.140 41.820 107.140 43.095 ;
        RECT 4.730 38.800 9.130 41.200 ;
        RECT 20.330 38.800 29.130 41.200 ;
        RECT 40.330 38.800 49.130 41.200 ;
        RECT 60.330 38.800 69.130 41.200 ;
        RECT 80.330 38.800 89.130 41.200 ;
        RECT 100.330 38.800 104.730 41.200 ;
        RECT 4.730 37.850 5.940 38.800 ;
        RECT 2.315 36.490 4.315 37.765 ;
        RECT 4.730 37.700 9.880 37.850 ;
        RECT 4.730 37.250 6.330 37.700 ;
        RECT 4.730 37.100 9.880 37.250 ;
        RECT 4.730 36.650 6.330 37.100 ;
        RECT 4.730 36.500 9.880 36.650 ;
        RECT 4.730 36.050 6.330 36.500 ;
        RECT 4.730 35.900 9.880 36.050 ;
        RECT 4.730 35.600 6.330 35.900 ;
        RECT 2.315 33.255 4.315 35.550 ;
        RECT 5.930 35.450 6.330 35.600 ;
        RECT 5.930 35.300 9.880 35.450 ;
        RECT 5.930 34.850 6.330 35.300 ;
        RECT 5.930 34.700 9.880 34.850 ;
        RECT 5.930 34.250 6.330 34.700 ;
        RECT 5.930 34.100 9.880 34.250 ;
        RECT 5.930 33.650 6.330 34.100 ;
        RECT 5.930 33.500 9.880 33.650 ;
        RECT 5.930 33.050 6.330 33.500 ;
        RECT 5.930 32.900 9.880 33.050 ;
        RECT 5.930 32.450 6.330 32.900 ;
        RECT 5.930 32.300 9.880 32.450 ;
        RECT 5.930 31.850 6.330 32.300 ;
        RECT 5.930 31.700 9.880 31.850 ;
        RECT 5.930 31.250 6.330 31.700 ;
        RECT 5.930 31.100 9.880 31.250 ;
        RECT 5.930 30.650 6.330 31.100 ;
        RECT 5.930 30.500 9.880 30.650 ;
        RECT 5.930 30.200 6.330 30.500 ;
        RECT 10.480 30.200 10.630 38.400 ;
        RECT 11.080 30.200 11.230 38.400 ;
        RECT 11.680 30.200 11.830 38.400 ;
        RECT 12.280 30.200 12.430 38.400 ;
        RECT 12.880 30.200 13.030 38.400 ;
        RECT 13.480 30.200 13.630 38.400 ;
        RECT 14.080 30.200 14.230 38.400 ;
        RECT 5.930 29.800 14.230 30.200 ;
        RECT 5.930 29.500 6.330 29.800 ;
        RECT 5.930 29.350 9.880 29.500 ;
        RECT 5.930 28.900 6.330 29.350 ;
        RECT 5.930 28.750 9.880 28.900 ;
        RECT 5.930 28.300 6.330 28.750 ;
        RECT 5.930 28.150 9.880 28.300 ;
        RECT 5.930 27.700 6.330 28.150 ;
        RECT 5.930 27.550 9.880 27.700 ;
        RECT 5.930 27.100 6.330 27.550 ;
        RECT 5.930 26.950 9.880 27.100 ;
        RECT 2.315 24.450 4.315 26.745 ;
        RECT 5.930 26.500 6.330 26.950 ;
        RECT 5.930 26.350 9.880 26.500 ;
        RECT 5.930 25.900 6.330 26.350 ;
        RECT 5.930 25.750 9.880 25.900 ;
        RECT 5.930 25.300 6.330 25.750 ;
        RECT 5.930 25.150 9.880 25.300 ;
        RECT 5.930 24.700 6.330 25.150 ;
        RECT 5.930 24.550 9.880 24.700 ;
        RECT 5.930 24.400 6.330 24.550 ;
        RECT 4.730 24.100 6.330 24.400 ;
        RECT 4.730 23.950 9.880 24.100 ;
        RECT 2.315 22.375 4.325 23.650 ;
        RECT 4.730 23.500 6.330 23.950 ;
        RECT 4.730 23.350 9.880 23.500 ;
        RECT 4.730 22.900 6.330 23.350 ;
        RECT 4.730 22.750 9.880 22.900 ;
        RECT 4.730 22.300 6.330 22.750 ;
        RECT 4.730 22.150 9.880 22.300 ;
        RECT 4.730 21.200 5.930 22.150 ;
        RECT 10.480 21.600 10.630 29.800 ;
        RECT 11.080 21.600 11.230 29.800 ;
        RECT 11.680 21.600 11.830 29.800 ;
        RECT 12.280 21.600 12.430 29.800 ;
        RECT 12.880 21.600 13.030 29.800 ;
        RECT 13.480 21.600 13.630 29.800 ;
        RECT 14.080 21.600 14.230 29.800 ;
        RECT 15.230 30.200 15.380 38.400 ;
        RECT 15.830 30.200 15.980 38.400 ;
        RECT 16.430 30.200 16.580 38.400 ;
        RECT 17.030 30.200 17.180 38.400 ;
        RECT 17.630 30.200 17.780 38.400 ;
        RECT 18.230 30.200 18.380 38.400 ;
        RECT 18.830 30.200 18.980 38.400 ;
        RECT 23.530 37.850 25.940 38.800 ;
        RECT 19.580 37.700 29.880 37.850 ;
        RECT 23.130 37.250 26.330 37.700 ;
        RECT 19.580 37.100 29.880 37.250 ;
        RECT 23.130 36.650 26.330 37.100 ;
        RECT 19.580 36.500 29.880 36.650 ;
        RECT 23.130 36.050 26.330 36.500 ;
        RECT 19.580 35.900 29.880 36.050 ;
        RECT 23.130 35.600 26.330 35.900 ;
        RECT 23.130 35.450 23.530 35.600 ;
        RECT 19.580 35.300 23.530 35.450 ;
        RECT 23.130 34.850 23.530 35.300 ;
        RECT 19.580 34.700 23.530 34.850 ;
        RECT 23.130 34.250 23.530 34.700 ;
        RECT 19.580 34.100 23.530 34.250 ;
        RECT 23.130 33.650 23.530 34.100 ;
        RECT 19.580 33.500 23.530 33.650 ;
        RECT 23.130 33.050 23.530 33.500 ;
        RECT 19.580 32.900 23.530 33.050 ;
        RECT 23.130 32.450 23.530 32.900 ;
        RECT 19.580 32.300 23.530 32.450 ;
        RECT 23.130 31.850 23.530 32.300 ;
        RECT 19.580 31.700 23.530 31.850 ;
        RECT 23.130 31.250 23.530 31.700 ;
        RECT 19.580 31.100 23.530 31.250 ;
        RECT 23.130 30.650 23.530 31.100 ;
        RECT 19.580 30.500 23.530 30.650 ;
        RECT 23.130 30.200 23.530 30.500 ;
        RECT 15.230 29.800 23.530 30.200 ;
        RECT 15.230 21.600 15.380 29.800 ;
        RECT 15.830 21.600 15.980 29.800 ;
        RECT 16.430 21.600 16.580 29.800 ;
        RECT 17.030 21.600 17.180 29.800 ;
        RECT 17.630 21.600 17.780 29.800 ;
        RECT 18.230 21.600 18.380 29.800 ;
        RECT 18.830 21.600 18.980 29.800 ;
        RECT 23.130 29.500 23.530 29.800 ;
        RECT 19.580 29.350 23.530 29.500 ;
        RECT 23.130 28.900 23.530 29.350 ;
        RECT 19.580 28.750 23.530 28.900 ;
        RECT 23.130 28.300 23.530 28.750 ;
        RECT 19.580 28.150 23.530 28.300 ;
        RECT 23.130 27.700 23.530 28.150 ;
        RECT 19.580 27.550 23.530 27.700 ;
        RECT 23.130 27.100 23.530 27.550 ;
        RECT 19.580 26.950 23.530 27.100 ;
        RECT 23.130 26.500 23.530 26.950 ;
        RECT 19.580 26.350 23.530 26.500 ;
        RECT 23.130 25.900 23.530 26.350 ;
        RECT 19.580 25.750 23.530 25.900 ;
        RECT 23.130 25.300 23.530 25.750 ;
        RECT 19.580 25.150 23.530 25.300 ;
        RECT 23.130 24.700 23.530 25.150 ;
        RECT 19.580 24.550 23.530 24.700 ;
        RECT 23.130 24.400 23.530 24.550 ;
        RECT 25.930 35.450 26.330 35.600 ;
        RECT 25.930 35.300 29.880 35.450 ;
        RECT 25.930 34.850 26.330 35.300 ;
        RECT 25.930 34.700 29.880 34.850 ;
        RECT 25.930 34.250 26.330 34.700 ;
        RECT 25.930 34.100 29.880 34.250 ;
        RECT 25.930 33.650 26.330 34.100 ;
        RECT 25.930 33.500 29.880 33.650 ;
        RECT 25.930 33.050 26.330 33.500 ;
        RECT 25.930 32.900 29.880 33.050 ;
        RECT 25.930 32.450 26.330 32.900 ;
        RECT 25.930 32.300 29.880 32.450 ;
        RECT 25.930 31.850 26.330 32.300 ;
        RECT 25.930 31.700 29.880 31.850 ;
        RECT 25.930 31.250 26.330 31.700 ;
        RECT 25.930 31.100 29.880 31.250 ;
        RECT 25.930 30.650 26.330 31.100 ;
        RECT 25.930 30.500 29.880 30.650 ;
        RECT 25.930 30.200 26.330 30.500 ;
        RECT 30.480 30.200 30.630 38.400 ;
        RECT 31.080 30.200 31.230 38.400 ;
        RECT 31.680 30.200 31.830 38.400 ;
        RECT 32.280 30.200 32.430 38.400 ;
        RECT 32.880 30.200 33.030 38.400 ;
        RECT 33.480 30.200 33.630 38.400 ;
        RECT 34.080 30.200 34.230 38.400 ;
        RECT 25.930 29.800 34.230 30.200 ;
        RECT 25.930 29.500 26.330 29.800 ;
        RECT 25.930 29.350 29.880 29.500 ;
        RECT 25.930 28.900 26.330 29.350 ;
        RECT 25.930 28.750 29.880 28.900 ;
        RECT 25.930 28.300 26.330 28.750 ;
        RECT 25.930 28.150 29.880 28.300 ;
        RECT 25.930 27.700 26.330 28.150 ;
        RECT 25.930 27.550 29.880 27.700 ;
        RECT 25.930 27.100 26.330 27.550 ;
        RECT 25.930 26.950 29.880 27.100 ;
        RECT 25.930 26.500 26.330 26.950 ;
        RECT 25.930 26.350 29.880 26.500 ;
        RECT 25.930 25.900 26.330 26.350 ;
        RECT 25.930 25.750 29.880 25.900 ;
        RECT 25.930 25.300 26.330 25.750 ;
        RECT 25.930 25.150 29.880 25.300 ;
        RECT 25.930 24.700 26.330 25.150 ;
        RECT 25.930 24.550 29.880 24.700 ;
        RECT 25.930 24.400 26.330 24.550 ;
        RECT 23.130 24.100 26.330 24.400 ;
        RECT 19.580 23.950 29.880 24.100 ;
        RECT 23.130 23.500 26.330 23.950 ;
        RECT 19.580 23.350 29.880 23.500 ;
        RECT 23.130 22.900 26.330 23.350 ;
        RECT 19.580 22.750 29.880 22.900 ;
        RECT 23.130 22.300 26.330 22.750 ;
        RECT 19.580 22.150 29.880 22.300 ;
        RECT 23.530 21.200 25.930 22.150 ;
        RECT 30.480 21.600 30.630 29.800 ;
        RECT 31.080 21.600 31.230 29.800 ;
        RECT 31.680 21.600 31.830 29.800 ;
        RECT 32.280 21.600 32.430 29.800 ;
        RECT 32.880 21.600 33.030 29.800 ;
        RECT 33.480 21.600 33.630 29.800 ;
        RECT 34.080 21.600 34.230 29.800 ;
        RECT 35.230 30.200 35.380 38.400 ;
        RECT 35.830 30.200 35.980 38.400 ;
        RECT 36.430 30.200 36.580 38.400 ;
        RECT 37.030 30.200 37.180 38.400 ;
        RECT 37.630 30.200 37.780 38.400 ;
        RECT 38.230 30.200 38.380 38.400 ;
        RECT 38.830 30.200 38.980 38.400 ;
        RECT 43.530 37.850 45.940 38.800 ;
        RECT 39.580 37.700 49.880 37.850 ;
        RECT 43.130 37.250 46.330 37.700 ;
        RECT 39.580 37.100 49.880 37.250 ;
        RECT 43.130 36.650 46.330 37.100 ;
        RECT 39.580 36.500 49.880 36.650 ;
        RECT 43.130 36.050 46.330 36.500 ;
        RECT 39.580 35.900 49.880 36.050 ;
        RECT 43.130 35.600 46.330 35.900 ;
        RECT 43.130 35.450 43.530 35.600 ;
        RECT 39.580 35.300 43.530 35.450 ;
        RECT 43.130 34.850 43.530 35.300 ;
        RECT 39.580 34.700 43.530 34.850 ;
        RECT 43.130 34.250 43.530 34.700 ;
        RECT 39.580 34.100 43.530 34.250 ;
        RECT 43.130 33.650 43.530 34.100 ;
        RECT 39.580 33.500 43.530 33.650 ;
        RECT 43.130 33.050 43.530 33.500 ;
        RECT 39.580 32.900 43.530 33.050 ;
        RECT 43.130 32.450 43.530 32.900 ;
        RECT 39.580 32.300 43.530 32.450 ;
        RECT 43.130 31.850 43.530 32.300 ;
        RECT 39.580 31.700 43.530 31.850 ;
        RECT 43.130 31.250 43.530 31.700 ;
        RECT 39.580 31.100 43.530 31.250 ;
        RECT 43.130 30.650 43.530 31.100 ;
        RECT 39.580 30.500 43.530 30.650 ;
        RECT 43.130 30.200 43.530 30.500 ;
        RECT 35.230 29.800 43.530 30.200 ;
        RECT 35.230 21.600 35.380 29.800 ;
        RECT 35.830 21.600 35.980 29.800 ;
        RECT 36.430 21.600 36.580 29.800 ;
        RECT 37.030 21.600 37.180 29.800 ;
        RECT 37.630 21.600 37.780 29.800 ;
        RECT 38.230 21.600 38.380 29.800 ;
        RECT 38.830 21.600 38.980 29.800 ;
        RECT 43.130 29.500 43.530 29.800 ;
        RECT 39.580 29.350 43.530 29.500 ;
        RECT 43.130 28.900 43.530 29.350 ;
        RECT 39.580 28.750 43.530 28.900 ;
        RECT 43.130 28.300 43.530 28.750 ;
        RECT 39.580 28.150 43.530 28.300 ;
        RECT 43.130 27.700 43.530 28.150 ;
        RECT 39.580 27.550 43.530 27.700 ;
        RECT 43.130 27.100 43.530 27.550 ;
        RECT 39.580 26.950 43.530 27.100 ;
        RECT 43.130 26.500 43.530 26.950 ;
        RECT 39.580 26.350 43.530 26.500 ;
        RECT 43.130 25.900 43.530 26.350 ;
        RECT 39.580 25.750 43.530 25.900 ;
        RECT 43.130 25.300 43.530 25.750 ;
        RECT 39.580 25.150 43.530 25.300 ;
        RECT 43.130 24.700 43.530 25.150 ;
        RECT 39.580 24.550 43.530 24.700 ;
        RECT 43.130 24.400 43.530 24.550 ;
        RECT 45.930 35.450 46.330 35.600 ;
        RECT 45.930 35.300 49.880 35.450 ;
        RECT 45.930 34.850 46.330 35.300 ;
        RECT 45.930 34.700 49.880 34.850 ;
        RECT 45.930 34.250 46.330 34.700 ;
        RECT 45.930 34.100 49.880 34.250 ;
        RECT 45.930 33.650 46.330 34.100 ;
        RECT 45.930 33.500 49.880 33.650 ;
        RECT 45.930 33.050 46.330 33.500 ;
        RECT 45.930 32.900 49.880 33.050 ;
        RECT 45.930 32.450 46.330 32.900 ;
        RECT 45.930 32.300 49.880 32.450 ;
        RECT 45.930 31.850 46.330 32.300 ;
        RECT 45.930 31.700 49.880 31.850 ;
        RECT 45.930 31.250 46.330 31.700 ;
        RECT 45.930 31.100 49.880 31.250 ;
        RECT 45.930 30.650 46.330 31.100 ;
        RECT 45.930 30.500 49.880 30.650 ;
        RECT 45.930 30.200 46.330 30.500 ;
        RECT 50.480 30.200 50.630 38.400 ;
        RECT 51.080 30.200 51.230 38.400 ;
        RECT 51.680 30.200 51.830 38.400 ;
        RECT 52.280 30.200 52.430 38.400 ;
        RECT 52.880 30.200 53.030 38.400 ;
        RECT 53.480 30.200 53.630 38.400 ;
        RECT 54.080 30.200 54.230 38.400 ;
        RECT 45.930 29.800 54.230 30.200 ;
        RECT 45.930 29.500 46.330 29.800 ;
        RECT 45.930 29.350 49.880 29.500 ;
        RECT 45.930 28.900 46.330 29.350 ;
        RECT 45.930 28.750 49.880 28.900 ;
        RECT 45.930 28.300 46.330 28.750 ;
        RECT 45.930 28.150 49.880 28.300 ;
        RECT 45.930 27.700 46.330 28.150 ;
        RECT 45.930 27.550 49.880 27.700 ;
        RECT 45.930 27.100 46.330 27.550 ;
        RECT 45.930 26.950 49.880 27.100 ;
        RECT 45.930 26.500 46.330 26.950 ;
        RECT 45.930 26.350 49.880 26.500 ;
        RECT 45.930 25.900 46.330 26.350 ;
        RECT 45.930 25.750 49.880 25.900 ;
        RECT 45.930 25.300 46.330 25.750 ;
        RECT 45.930 25.150 49.880 25.300 ;
        RECT 45.930 24.700 46.330 25.150 ;
        RECT 45.930 24.550 49.880 24.700 ;
        RECT 45.930 24.400 46.330 24.550 ;
        RECT 43.130 24.100 46.330 24.400 ;
        RECT 39.580 23.950 49.880 24.100 ;
        RECT 43.130 23.500 46.330 23.950 ;
        RECT 39.580 23.350 49.880 23.500 ;
        RECT 43.130 22.900 46.330 23.350 ;
        RECT 39.580 22.750 49.880 22.900 ;
        RECT 43.130 22.300 46.330 22.750 ;
        RECT 39.580 22.150 49.880 22.300 ;
        RECT 43.530 21.200 45.930 22.150 ;
        RECT 50.480 21.600 50.630 29.800 ;
        RECT 51.080 21.600 51.230 29.800 ;
        RECT 51.680 21.600 51.830 29.800 ;
        RECT 52.280 21.600 52.430 29.800 ;
        RECT 52.880 21.600 53.030 29.800 ;
        RECT 53.480 21.600 53.630 29.800 ;
        RECT 54.080 21.600 54.230 29.800 ;
        RECT 55.230 30.200 55.380 38.400 ;
        RECT 55.830 30.200 55.980 38.400 ;
        RECT 56.430 30.200 56.580 38.400 ;
        RECT 57.030 30.200 57.180 38.400 ;
        RECT 57.630 30.200 57.780 38.400 ;
        RECT 58.230 30.200 58.380 38.400 ;
        RECT 58.830 30.200 58.980 38.400 ;
        RECT 63.530 37.850 65.940 38.800 ;
        RECT 59.580 37.700 69.880 37.850 ;
        RECT 63.130 37.250 66.330 37.700 ;
        RECT 59.580 37.100 69.880 37.250 ;
        RECT 63.130 36.650 66.330 37.100 ;
        RECT 59.580 36.500 69.880 36.650 ;
        RECT 63.130 36.050 66.330 36.500 ;
        RECT 59.580 35.900 69.880 36.050 ;
        RECT 63.130 35.600 66.330 35.900 ;
        RECT 63.130 35.450 63.530 35.600 ;
        RECT 59.580 35.300 63.530 35.450 ;
        RECT 63.130 34.850 63.530 35.300 ;
        RECT 59.580 34.700 63.530 34.850 ;
        RECT 63.130 34.250 63.530 34.700 ;
        RECT 59.580 34.100 63.530 34.250 ;
        RECT 63.130 33.650 63.530 34.100 ;
        RECT 59.580 33.500 63.530 33.650 ;
        RECT 63.130 33.050 63.530 33.500 ;
        RECT 59.580 32.900 63.530 33.050 ;
        RECT 63.130 32.450 63.530 32.900 ;
        RECT 59.580 32.300 63.530 32.450 ;
        RECT 63.130 31.850 63.530 32.300 ;
        RECT 59.580 31.700 63.530 31.850 ;
        RECT 63.130 31.250 63.530 31.700 ;
        RECT 59.580 31.100 63.530 31.250 ;
        RECT 63.130 30.650 63.530 31.100 ;
        RECT 59.580 30.500 63.530 30.650 ;
        RECT 63.130 30.200 63.530 30.500 ;
        RECT 55.230 29.800 63.530 30.200 ;
        RECT 55.230 21.600 55.380 29.800 ;
        RECT 55.830 21.600 55.980 29.800 ;
        RECT 56.430 21.600 56.580 29.800 ;
        RECT 57.030 21.600 57.180 29.800 ;
        RECT 57.630 21.600 57.780 29.800 ;
        RECT 58.230 21.600 58.380 29.800 ;
        RECT 58.830 21.600 58.980 29.800 ;
        RECT 63.130 29.500 63.530 29.800 ;
        RECT 59.580 29.350 63.530 29.500 ;
        RECT 63.130 28.900 63.530 29.350 ;
        RECT 59.580 28.750 63.530 28.900 ;
        RECT 63.130 28.300 63.530 28.750 ;
        RECT 59.580 28.150 63.530 28.300 ;
        RECT 63.130 27.700 63.530 28.150 ;
        RECT 59.580 27.550 63.530 27.700 ;
        RECT 63.130 27.100 63.530 27.550 ;
        RECT 59.580 26.950 63.530 27.100 ;
        RECT 63.130 26.500 63.530 26.950 ;
        RECT 59.580 26.350 63.530 26.500 ;
        RECT 63.130 25.900 63.530 26.350 ;
        RECT 59.580 25.750 63.530 25.900 ;
        RECT 63.130 25.300 63.530 25.750 ;
        RECT 59.580 25.150 63.530 25.300 ;
        RECT 63.130 24.700 63.530 25.150 ;
        RECT 59.580 24.550 63.530 24.700 ;
        RECT 63.130 24.400 63.530 24.550 ;
        RECT 65.930 35.450 66.330 35.600 ;
        RECT 65.930 35.300 69.880 35.450 ;
        RECT 65.930 34.850 66.330 35.300 ;
        RECT 65.930 34.700 69.880 34.850 ;
        RECT 65.930 34.250 66.330 34.700 ;
        RECT 65.930 34.100 69.880 34.250 ;
        RECT 65.930 33.650 66.330 34.100 ;
        RECT 65.930 33.500 69.880 33.650 ;
        RECT 65.930 33.050 66.330 33.500 ;
        RECT 65.930 32.900 69.880 33.050 ;
        RECT 65.930 32.450 66.330 32.900 ;
        RECT 65.930 32.300 69.880 32.450 ;
        RECT 65.930 31.850 66.330 32.300 ;
        RECT 65.930 31.700 69.880 31.850 ;
        RECT 65.930 31.250 66.330 31.700 ;
        RECT 65.930 31.100 69.880 31.250 ;
        RECT 65.930 30.650 66.330 31.100 ;
        RECT 65.930 30.500 69.880 30.650 ;
        RECT 65.930 30.200 66.330 30.500 ;
        RECT 70.480 30.200 70.630 38.400 ;
        RECT 71.080 30.200 71.230 38.400 ;
        RECT 71.680 30.200 71.830 38.400 ;
        RECT 72.280 30.200 72.430 38.400 ;
        RECT 72.880 30.200 73.030 38.400 ;
        RECT 73.480 30.200 73.630 38.400 ;
        RECT 74.080 30.200 74.230 38.400 ;
        RECT 65.930 29.800 74.230 30.200 ;
        RECT 65.930 29.500 66.330 29.800 ;
        RECT 65.930 29.350 69.880 29.500 ;
        RECT 65.930 28.900 66.330 29.350 ;
        RECT 65.930 28.750 69.880 28.900 ;
        RECT 65.930 28.300 66.330 28.750 ;
        RECT 65.930 28.150 69.880 28.300 ;
        RECT 65.930 27.700 66.330 28.150 ;
        RECT 65.930 27.550 69.880 27.700 ;
        RECT 65.930 27.100 66.330 27.550 ;
        RECT 65.930 26.950 69.880 27.100 ;
        RECT 65.930 26.500 66.330 26.950 ;
        RECT 65.930 26.350 69.880 26.500 ;
        RECT 65.930 25.900 66.330 26.350 ;
        RECT 65.930 25.750 69.880 25.900 ;
        RECT 65.930 25.300 66.330 25.750 ;
        RECT 65.930 25.150 69.880 25.300 ;
        RECT 65.930 24.700 66.330 25.150 ;
        RECT 65.930 24.550 69.880 24.700 ;
        RECT 65.930 24.400 66.330 24.550 ;
        RECT 63.130 24.100 66.330 24.400 ;
        RECT 59.580 23.950 69.880 24.100 ;
        RECT 63.130 23.500 66.330 23.950 ;
        RECT 59.580 23.350 69.880 23.500 ;
        RECT 63.130 22.900 66.330 23.350 ;
        RECT 59.580 22.750 69.880 22.900 ;
        RECT 63.130 22.300 66.330 22.750 ;
        RECT 59.580 22.150 69.880 22.300 ;
        RECT 63.530 21.200 65.930 22.150 ;
        RECT 70.480 21.600 70.630 29.800 ;
        RECT 71.080 21.600 71.230 29.800 ;
        RECT 71.680 21.600 71.830 29.800 ;
        RECT 72.280 21.600 72.430 29.800 ;
        RECT 72.880 21.600 73.030 29.800 ;
        RECT 73.480 21.600 73.630 29.800 ;
        RECT 74.080 21.600 74.230 29.800 ;
        RECT 75.230 30.200 75.380 38.400 ;
        RECT 75.830 30.200 75.980 38.400 ;
        RECT 76.430 30.200 76.580 38.400 ;
        RECT 77.030 30.200 77.180 38.400 ;
        RECT 77.630 30.200 77.780 38.400 ;
        RECT 78.230 30.200 78.380 38.400 ;
        RECT 78.830 30.200 78.980 38.400 ;
        RECT 83.530 37.850 85.940 38.800 ;
        RECT 79.580 37.700 89.880 37.850 ;
        RECT 83.130 37.250 86.330 37.700 ;
        RECT 79.580 37.100 89.880 37.250 ;
        RECT 83.130 36.650 86.330 37.100 ;
        RECT 79.580 36.500 89.880 36.650 ;
        RECT 83.130 36.050 86.330 36.500 ;
        RECT 79.580 35.900 89.880 36.050 ;
        RECT 83.130 35.600 86.330 35.900 ;
        RECT 83.130 35.450 83.530 35.600 ;
        RECT 79.580 35.300 83.530 35.450 ;
        RECT 83.130 34.850 83.530 35.300 ;
        RECT 79.580 34.700 83.530 34.850 ;
        RECT 83.130 34.250 83.530 34.700 ;
        RECT 79.580 34.100 83.530 34.250 ;
        RECT 83.130 33.650 83.530 34.100 ;
        RECT 79.580 33.500 83.530 33.650 ;
        RECT 83.130 33.050 83.530 33.500 ;
        RECT 79.580 32.900 83.530 33.050 ;
        RECT 83.130 32.450 83.530 32.900 ;
        RECT 79.580 32.300 83.530 32.450 ;
        RECT 83.130 31.850 83.530 32.300 ;
        RECT 79.580 31.700 83.530 31.850 ;
        RECT 83.130 31.250 83.530 31.700 ;
        RECT 79.580 31.100 83.530 31.250 ;
        RECT 83.130 30.650 83.530 31.100 ;
        RECT 79.580 30.500 83.530 30.650 ;
        RECT 83.130 30.200 83.530 30.500 ;
        RECT 75.230 29.800 83.530 30.200 ;
        RECT 75.230 21.600 75.380 29.800 ;
        RECT 75.830 21.600 75.980 29.800 ;
        RECT 76.430 21.600 76.580 29.800 ;
        RECT 77.030 21.600 77.180 29.800 ;
        RECT 77.630 21.600 77.780 29.800 ;
        RECT 78.230 21.600 78.380 29.800 ;
        RECT 78.830 21.600 78.980 29.800 ;
        RECT 83.130 29.500 83.530 29.800 ;
        RECT 79.580 29.350 83.530 29.500 ;
        RECT 83.130 28.900 83.530 29.350 ;
        RECT 79.580 28.750 83.530 28.900 ;
        RECT 83.130 28.300 83.530 28.750 ;
        RECT 79.580 28.150 83.530 28.300 ;
        RECT 83.130 27.700 83.530 28.150 ;
        RECT 79.580 27.550 83.530 27.700 ;
        RECT 83.130 27.100 83.530 27.550 ;
        RECT 79.580 26.950 83.530 27.100 ;
        RECT 83.130 26.500 83.530 26.950 ;
        RECT 79.580 26.350 83.530 26.500 ;
        RECT 83.130 25.900 83.530 26.350 ;
        RECT 79.580 25.750 83.530 25.900 ;
        RECT 83.130 25.300 83.530 25.750 ;
        RECT 79.580 25.150 83.530 25.300 ;
        RECT 83.130 24.700 83.530 25.150 ;
        RECT 79.580 24.550 83.530 24.700 ;
        RECT 83.130 24.400 83.530 24.550 ;
        RECT 85.930 35.450 86.330 35.600 ;
        RECT 85.930 35.300 89.880 35.450 ;
        RECT 85.930 34.850 86.330 35.300 ;
        RECT 85.930 34.700 89.880 34.850 ;
        RECT 85.930 34.250 86.330 34.700 ;
        RECT 85.930 34.100 89.880 34.250 ;
        RECT 85.930 33.650 86.330 34.100 ;
        RECT 85.930 33.500 89.880 33.650 ;
        RECT 85.930 33.050 86.330 33.500 ;
        RECT 85.930 32.900 89.880 33.050 ;
        RECT 85.930 32.450 86.330 32.900 ;
        RECT 85.930 32.300 89.880 32.450 ;
        RECT 85.930 31.850 86.330 32.300 ;
        RECT 85.930 31.700 89.880 31.850 ;
        RECT 85.930 31.250 86.330 31.700 ;
        RECT 85.930 31.100 89.880 31.250 ;
        RECT 85.930 30.650 86.330 31.100 ;
        RECT 85.930 30.500 89.880 30.650 ;
        RECT 85.930 30.200 86.330 30.500 ;
        RECT 90.480 30.200 90.630 38.400 ;
        RECT 91.080 30.200 91.230 38.400 ;
        RECT 91.680 30.200 91.830 38.400 ;
        RECT 92.280 30.200 92.430 38.400 ;
        RECT 92.880 30.200 93.030 38.400 ;
        RECT 93.480 30.200 93.630 38.400 ;
        RECT 94.080 30.200 94.230 38.400 ;
        RECT 85.930 29.800 94.230 30.200 ;
        RECT 85.930 29.500 86.330 29.800 ;
        RECT 85.930 29.350 89.880 29.500 ;
        RECT 85.930 28.900 86.330 29.350 ;
        RECT 85.930 28.750 89.880 28.900 ;
        RECT 85.930 28.300 86.330 28.750 ;
        RECT 85.930 28.150 89.880 28.300 ;
        RECT 85.930 27.700 86.330 28.150 ;
        RECT 85.930 27.550 89.880 27.700 ;
        RECT 85.930 27.100 86.330 27.550 ;
        RECT 85.930 26.950 89.880 27.100 ;
        RECT 85.930 26.500 86.330 26.950 ;
        RECT 85.930 26.350 89.880 26.500 ;
        RECT 85.930 25.900 86.330 26.350 ;
        RECT 85.930 25.750 89.880 25.900 ;
        RECT 85.930 25.300 86.330 25.750 ;
        RECT 85.930 25.150 89.880 25.300 ;
        RECT 85.930 24.700 86.330 25.150 ;
        RECT 85.930 24.550 89.880 24.700 ;
        RECT 85.930 24.400 86.330 24.550 ;
        RECT 83.130 24.100 86.330 24.400 ;
        RECT 79.580 23.950 89.880 24.100 ;
        RECT 83.130 23.500 86.330 23.950 ;
        RECT 79.580 23.350 89.880 23.500 ;
        RECT 83.130 22.900 86.330 23.350 ;
        RECT 79.580 22.750 89.880 22.900 ;
        RECT 83.130 22.300 86.330 22.750 ;
        RECT 79.580 22.150 89.880 22.300 ;
        RECT 83.530 21.200 85.930 22.150 ;
        RECT 90.480 21.600 90.630 29.800 ;
        RECT 91.080 21.600 91.230 29.800 ;
        RECT 91.680 21.600 91.830 29.800 ;
        RECT 92.280 21.600 92.430 29.800 ;
        RECT 92.880 21.600 93.030 29.800 ;
        RECT 93.480 21.600 93.630 29.800 ;
        RECT 94.080 21.600 94.230 29.800 ;
        RECT 95.230 30.200 95.380 38.400 ;
        RECT 95.830 30.200 95.980 38.400 ;
        RECT 96.430 30.200 96.580 38.400 ;
        RECT 97.030 30.200 97.180 38.400 ;
        RECT 97.630 30.200 97.780 38.400 ;
        RECT 98.230 30.200 98.380 38.400 ;
        RECT 98.830 30.200 98.980 38.400 ;
        RECT 103.530 37.850 104.730 38.800 ;
        RECT 99.580 37.700 104.730 37.850 ;
        RECT 103.130 37.250 104.730 37.700 ;
        RECT 99.580 37.100 104.730 37.250 ;
        RECT 103.130 36.650 104.730 37.100 ;
        RECT 99.580 36.500 104.730 36.650 ;
        RECT 103.130 36.050 104.730 36.500 ;
        RECT 99.580 35.900 104.730 36.050 ;
        RECT 105.135 36.035 107.135 37.310 ;
        RECT 103.130 35.600 104.730 35.900 ;
        RECT 103.130 35.450 103.530 35.600 ;
        RECT 99.580 35.300 103.530 35.450 ;
        RECT 103.130 34.850 103.530 35.300 ;
        RECT 99.580 34.700 103.530 34.850 ;
        RECT 103.130 34.250 103.530 34.700 ;
        RECT 99.580 34.100 103.530 34.250 ;
        RECT 103.130 33.650 103.530 34.100 ;
        RECT 99.580 33.500 103.530 33.650 ;
        RECT 103.130 33.050 103.530 33.500 ;
        RECT 99.580 32.900 103.530 33.050 ;
        RECT 103.130 32.450 103.530 32.900 ;
        RECT 99.580 32.300 103.530 32.450 ;
        RECT 103.130 31.850 103.530 32.300 ;
        RECT 99.580 31.700 103.530 31.850 ;
        RECT 103.130 31.250 103.530 31.700 ;
        RECT 99.580 31.100 103.530 31.250 ;
        RECT 103.130 30.650 103.530 31.100 ;
        RECT 99.580 30.500 103.530 30.650 ;
        RECT 103.130 30.200 103.530 30.500 ;
        RECT 95.230 29.800 103.530 30.200 ;
        RECT 95.230 21.600 95.380 29.800 ;
        RECT 95.830 21.600 95.980 29.800 ;
        RECT 96.430 21.600 96.580 29.800 ;
        RECT 97.030 21.600 97.180 29.800 ;
        RECT 97.630 21.600 97.780 29.800 ;
        RECT 98.230 21.600 98.380 29.800 ;
        RECT 98.830 21.600 98.980 29.800 ;
        RECT 103.130 29.500 103.530 29.800 ;
        RECT 99.580 29.350 103.530 29.500 ;
        RECT 103.130 28.900 103.530 29.350 ;
        RECT 99.580 28.750 103.530 28.900 ;
        RECT 103.130 28.300 103.530 28.750 ;
        RECT 99.580 28.150 103.530 28.300 ;
        RECT 103.130 27.700 103.530 28.150 ;
        RECT 99.580 27.550 103.530 27.700 ;
        RECT 103.130 27.100 103.530 27.550 ;
        RECT 99.580 26.950 103.530 27.100 ;
        RECT 103.130 26.500 103.530 26.950 ;
        RECT 99.580 26.350 103.530 26.500 ;
        RECT 103.130 25.900 103.530 26.350 ;
        RECT 99.580 25.750 103.530 25.900 ;
        RECT 103.130 25.300 103.530 25.750 ;
        RECT 99.580 25.150 103.530 25.300 ;
        RECT 103.130 24.700 103.530 25.150 ;
        RECT 99.580 24.550 103.530 24.700 ;
        RECT 103.130 24.400 103.530 24.550 ;
        RECT 103.130 24.100 104.730 24.400 ;
        RECT 99.580 23.950 104.730 24.100 ;
        RECT 103.130 23.500 104.730 23.950 ;
        RECT 99.580 23.350 104.730 23.500 ;
        RECT 103.130 22.900 104.730 23.350 ;
        RECT 99.580 22.750 104.730 22.900 ;
        RECT 103.130 22.300 104.730 22.750 ;
        RECT 99.580 22.150 104.730 22.300 ;
        RECT 103.530 21.200 104.730 22.150 ;
        RECT 105.140 21.820 107.140 23.095 ;
        RECT 4.730 18.800 9.130 21.200 ;
        RECT 20.330 18.800 29.130 21.200 ;
        RECT 40.330 18.800 49.130 21.200 ;
        RECT 60.330 18.800 69.130 21.200 ;
        RECT 80.330 18.800 89.130 21.200 ;
        RECT 100.330 18.800 104.730 21.200 ;
        RECT 4.730 17.850 5.940 18.800 ;
        RECT 2.315 16.490 4.315 17.765 ;
        RECT 4.730 17.700 9.880 17.850 ;
        RECT 4.730 17.250 6.330 17.700 ;
        RECT 4.730 17.100 9.880 17.250 ;
        RECT 4.730 16.650 6.330 17.100 ;
        RECT 4.730 16.500 9.880 16.650 ;
        RECT 4.730 16.050 6.330 16.500 ;
        RECT 4.730 15.900 9.880 16.050 ;
        RECT 4.730 15.600 6.330 15.900 ;
        RECT 2.315 13.255 4.315 15.550 ;
        RECT 5.930 15.450 6.330 15.600 ;
        RECT 5.930 15.300 9.880 15.450 ;
        RECT 5.930 14.850 6.330 15.300 ;
        RECT 5.930 14.700 9.880 14.850 ;
        RECT 5.930 14.250 6.330 14.700 ;
        RECT 5.930 14.100 9.880 14.250 ;
        RECT 5.930 13.650 6.330 14.100 ;
        RECT 5.930 13.500 9.880 13.650 ;
        RECT 5.930 13.050 6.330 13.500 ;
        RECT 5.930 12.900 9.880 13.050 ;
        RECT 5.930 12.450 6.330 12.900 ;
        RECT 5.930 12.300 9.880 12.450 ;
        RECT 5.930 11.850 6.330 12.300 ;
        RECT 5.930 11.700 9.880 11.850 ;
        RECT 5.930 11.250 6.330 11.700 ;
        RECT 5.930 11.100 9.880 11.250 ;
        RECT 5.930 10.650 6.330 11.100 ;
        RECT 5.930 10.500 9.880 10.650 ;
        RECT 5.930 10.200 6.330 10.500 ;
        RECT 10.480 10.200 10.630 18.400 ;
        RECT 11.080 10.200 11.230 18.400 ;
        RECT 11.680 10.200 11.830 18.400 ;
        RECT 12.280 10.200 12.430 18.400 ;
        RECT 12.880 10.200 13.030 18.400 ;
        RECT 13.480 10.200 13.630 18.400 ;
        RECT 14.080 10.200 14.230 18.400 ;
        RECT 5.930 9.800 14.230 10.200 ;
        RECT 5.930 9.500 6.330 9.800 ;
        RECT 5.930 9.350 9.880 9.500 ;
        RECT 5.930 8.900 6.330 9.350 ;
        RECT 5.930 8.750 9.880 8.900 ;
        RECT 5.930 8.300 6.330 8.750 ;
        RECT 5.930 8.150 9.880 8.300 ;
        RECT 5.930 7.700 6.330 8.150 ;
        RECT 5.930 7.550 9.880 7.700 ;
        RECT 5.930 7.100 6.330 7.550 ;
        RECT 5.930 6.950 9.880 7.100 ;
        RECT 2.315 4.450 4.315 6.745 ;
        RECT 5.930 6.500 6.330 6.950 ;
        RECT 5.930 6.350 9.880 6.500 ;
        RECT 5.930 5.900 6.330 6.350 ;
        RECT 5.930 5.750 9.880 5.900 ;
        RECT 5.930 5.300 6.330 5.750 ;
        RECT 5.930 5.150 9.880 5.300 ;
        RECT 5.930 4.700 6.330 5.150 ;
        RECT 5.930 4.550 9.880 4.700 ;
        RECT 5.930 4.400 6.330 4.550 ;
        RECT 4.730 4.100 6.330 4.400 ;
        RECT 4.730 3.950 9.880 4.100 ;
        RECT 2.315 2.375 4.325 3.650 ;
        RECT 4.730 3.500 6.330 3.950 ;
        RECT 4.730 3.350 9.880 3.500 ;
        RECT 4.730 2.900 6.330 3.350 ;
        RECT 4.730 2.750 9.880 2.900 ;
        RECT 4.730 2.300 6.330 2.750 ;
        RECT 4.730 2.150 9.880 2.300 ;
        RECT 4.730 1.200 5.930 2.150 ;
        RECT 10.480 1.600 10.630 9.800 ;
        RECT 11.080 1.600 11.230 9.800 ;
        RECT 11.680 1.600 11.830 9.800 ;
        RECT 12.280 1.600 12.430 9.800 ;
        RECT 12.880 1.600 13.030 9.800 ;
        RECT 13.480 1.600 13.630 9.800 ;
        RECT 14.080 1.600 14.230 9.800 ;
        RECT 15.230 10.200 15.380 18.400 ;
        RECT 15.830 10.200 15.980 18.400 ;
        RECT 16.430 10.200 16.580 18.400 ;
        RECT 17.030 10.200 17.180 18.400 ;
        RECT 17.630 10.200 17.780 18.400 ;
        RECT 18.230 10.200 18.380 18.400 ;
        RECT 18.830 10.200 18.980 18.400 ;
        RECT 23.530 17.850 25.940 18.800 ;
        RECT 19.580 17.700 29.880 17.850 ;
        RECT 23.130 17.250 26.330 17.700 ;
        RECT 19.580 17.100 29.880 17.250 ;
        RECT 23.130 16.650 26.330 17.100 ;
        RECT 19.580 16.500 29.880 16.650 ;
        RECT 23.130 16.050 26.330 16.500 ;
        RECT 19.580 15.900 29.880 16.050 ;
        RECT 23.130 15.600 26.330 15.900 ;
        RECT 23.130 15.450 23.530 15.600 ;
        RECT 19.580 15.300 23.530 15.450 ;
        RECT 23.130 14.850 23.530 15.300 ;
        RECT 19.580 14.700 23.530 14.850 ;
        RECT 23.130 14.250 23.530 14.700 ;
        RECT 19.580 14.100 23.530 14.250 ;
        RECT 23.130 13.650 23.530 14.100 ;
        RECT 19.580 13.500 23.530 13.650 ;
        RECT 23.130 13.050 23.530 13.500 ;
        RECT 19.580 12.900 23.530 13.050 ;
        RECT 23.130 12.450 23.530 12.900 ;
        RECT 19.580 12.300 23.530 12.450 ;
        RECT 23.130 11.850 23.530 12.300 ;
        RECT 19.580 11.700 23.530 11.850 ;
        RECT 23.130 11.250 23.530 11.700 ;
        RECT 19.580 11.100 23.530 11.250 ;
        RECT 23.130 10.650 23.530 11.100 ;
        RECT 19.580 10.500 23.530 10.650 ;
        RECT 23.130 10.200 23.530 10.500 ;
        RECT 15.230 9.800 23.530 10.200 ;
        RECT 15.230 1.600 15.380 9.800 ;
        RECT 15.830 1.600 15.980 9.800 ;
        RECT 16.430 1.600 16.580 9.800 ;
        RECT 17.030 1.600 17.180 9.800 ;
        RECT 17.630 1.600 17.780 9.800 ;
        RECT 18.230 1.600 18.380 9.800 ;
        RECT 18.830 1.600 18.980 9.800 ;
        RECT 23.130 9.500 23.530 9.800 ;
        RECT 19.580 9.350 23.530 9.500 ;
        RECT 23.130 8.900 23.530 9.350 ;
        RECT 19.580 8.750 23.530 8.900 ;
        RECT 23.130 8.300 23.530 8.750 ;
        RECT 19.580 8.150 23.530 8.300 ;
        RECT 23.130 7.700 23.530 8.150 ;
        RECT 19.580 7.550 23.530 7.700 ;
        RECT 23.130 7.100 23.530 7.550 ;
        RECT 19.580 6.950 23.530 7.100 ;
        RECT 23.130 6.500 23.530 6.950 ;
        RECT 19.580 6.350 23.530 6.500 ;
        RECT 23.130 5.900 23.530 6.350 ;
        RECT 19.580 5.750 23.530 5.900 ;
        RECT 23.130 5.300 23.530 5.750 ;
        RECT 19.580 5.150 23.530 5.300 ;
        RECT 23.130 4.700 23.530 5.150 ;
        RECT 19.580 4.550 23.530 4.700 ;
        RECT 23.130 4.400 23.530 4.550 ;
        RECT 25.930 15.450 26.330 15.600 ;
        RECT 25.930 15.300 29.880 15.450 ;
        RECT 25.930 14.850 26.330 15.300 ;
        RECT 25.930 14.700 29.880 14.850 ;
        RECT 25.930 14.250 26.330 14.700 ;
        RECT 25.930 14.100 29.880 14.250 ;
        RECT 25.930 13.650 26.330 14.100 ;
        RECT 25.930 13.500 29.880 13.650 ;
        RECT 25.930 13.050 26.330 13.500 ;
        RECT 25.930 12.900 29.880 13.050 ;
        RECT 25.930 12.450 26.330 12.900 ;
        RECT 25.930 12.300 29.880 12.450 ;
        RECT 25.930 11.850 26.330 12.300 ;
        RECT 25.930 11.700 29.880 11.850 ;
        RECT 25.930 11.250 26.330 11.700 ;
        RECT 25.930 11.100 29.880 11.250 ;
        RECT 25.930 10.650 26.330 11.100 ;
        RECT 25.930 10.500 29.880 10.650 ;
        RECT 25.930 10.200 26.330 10.500 ;
        RECT 30.480 10.200 30.630 18.400 ;
        RECT 31.080 10.200 31.230 18.400 ;
        RECT 31.680 10.200 31.830 18.400 ;
        RECT 32.280 10.200 32.430 18.400 ;
        RECT 32.880 10.200 33.030 18.400 ;
        RECT 33.480 10.200 33.630 18.400 ;
        RECT 34.080 10.200 34.230 18.400 ;
        RECT 25.930 9.800 34.230 10.200 ;
        RECT 25.930 9.500 26.330 9.800 ;
        RECT 25.930 9.350 29.880 9.500 ;
        RECT 25.930 8.900 26.330 9.350 ;
        RECT 25.930 8.750 29.880 8.900 ;
        RECT 25.930 8.300 26.330 8.750 ;
        RECT 25.930 8.150 29.880 8.300 ;
        RECT 25.930 7.700 26.330 8.150 ;
        RECT 25.930 7.550 29.880 7.700 ;
        RECT 25.930 7.100 26.330 7.550 ;
        RECT 25.930 6.950 29.880 7.100 ;
        RECT 25.930 6.500 26.330 6.950 ;
        RECT 25.930 6.350 29.880 6.500 ;
        RECT 25.930 5.900 26.330 6.350 ;
        RECT 25.930 5.750 29.880 5.900 ;
        RECT 25.930 5.300 26.330 5.750 ;
        RECT 25.930 5.150 29.880 5.300 ;
        RECT 25.930 4.700 26.330 5.150 ;
        RECT 25.930 4.550 29.880 4.700 ;
        RECT 25.930 4.400 26.330 4.550 ;
        RECT 23.130 4.100 26.330 4.400 ;
        RECT 19.580 3.950 29.880 4.100 ;
        RECT 23.130 3.500 26.330 3.950 ;
        RECT 19.580 3.350 29.880 3.500 ;
        RECT 23.130 2.900 26.330 3.350 ;
        RECT 19.580 2.750 29.880 2.900 ;
        RECT 23.130 2.300 26.330 2.750 ;
        RECT 19.580 2.150 29.880 2.300 ;
        RECT 23.530 1.200 25.930 2.150 ;
        RECT 30.480 1.600 30.630 9.800 ;
        RECT 31.080 1.600 31.230 9.800 ;
        RECT 31.680 1.600 31.830 9.800 ;
        RECT 32.280 1.600 32.430 9.800 ;
        RECT 32.880 1.600 33.030 9.800 ;
        RECT 33.480 1.600 33.630 9.800 ;
        RECT 34.080 1.600 34.230 9.800 ;
        RECT 35.230 10.200 35.380 18.400 ;
        RECT 35.830 10.200 35.980 18.400 ;
        RECT 36.430 10.200 36.580 18.400 ;
        RECT 37.030 10.200 37.180 18.400 ;
        RECT 37.630 10.200 37.780 18.400 ;
        RECT 38.230 10.200 38.380 18.400 ;
        RECT 38.830 10.200 38.980 18.400 ;
        RECT 43.530 17.850 45.940 18.800 ;
        RECT 39.580 17.700 49.880 17.850 ;
        RECT 43.130 17.250 46.330 17.700 ;
        RECT 39.580 17.100 49.880 17.250 ;
        RECT 43.130 16.650 46.330 17.100 ;
        RECT 39.580 16.500 49.880 16.650 ;
        RECT 43.130 16.050 46.330 16.500 ;
        RECT 39.580 15.900 49.880 16.050 ;
        RECT 43.130 15.600 46.330 15.900 ;
        RECT 43.130 15.450 43.530 15.600 ;
        RECT 39.580 15.300 43.530 15.450 ;
        RECT 43.130 14.850 43.530 15.300 ;
        RECT 39.580 14.700 43.530 14.850 ;
        RECT 43.130 14.250 43.530 14.700 ;
        RECT 39.580 14.100 43.530 14.250 ;
        RECT 43.130 13.650 43.530 14.100 ;
        RECT 39.580 13.500 43.530 13.650 ;
        RECT 43.130 13.050 43.530 13.500 ;
        RECT 39.580 12.900 43.530 13.050 ;
        RECT 43.130 12.450 43.530 12.900 ;
        RECT 39.580 12.300 43.530 12.450 ;
        RECT 43.130 11.850 43.530 12.300 ;
        RECT 39.580 11.700 43.530 11.850 ;
        RECT 43.130 11.250 43.530 11.700 ;
        RECT 39.580 11.100 43.530 11.250 ;
        RECT 43.130 10.650 43.530 11.100 ;
        RECT 39.580 10.500 43.530 10.650 ;
        RECT 43.130 10.200 43.530 10.500 ;
        RECT 35.230 9.800 43.530 10.200 ;
        RECT 35.230 1.600 35.380 9.800 ;
        RECT 35.830 1.600 35.980 9.800 ;
        RECT 36.430 1.600 36.580 9.800 ;
        RECT 37.030 1.600 37.180 9.800 ;
        RECT 37.630 1.600 37.780 9.800 ;
        RECT 38.230 1.600 38.380 9.800 ;
        RECT 38.830 1.600 38.980 9.800 ;
        RECT 43.130 9.500 43.530 9.800 ;
        RECT 39.580 9.350 43.530 9.500 ;
        RECT 43.130 8.900 43.530 9.350 ;
        RECT 39.580 8.750 43.530 8.900 ;
        RECT 43.130 8.300 43.530 8.750 ;
        RECT 39.580 8.150 43.530 8.300 ;
        RECT 43.130 7.700 43.530 8.150 ;
        RECT 39.580 7.550 43.530 7.700 ;
        RECT 43.130 7.100 43.530 7.550 ;
        RECT 39.580 6.950 43.530 7.100 ;
        RECT 43.130 6.500 43.530 6.950 ;
        RECT 39.580 6.350 43.530 6.500 ;
        RECT 43.130 5.900 43.530 6.350 ;
        RECT 39.580 5.750 43.530 5.900 ;
        RECT 43.130 5.300 43.530 5.750 ;
        RECT 39.580 5.150 43.530 5.300 ;
        RECT 43.130 4.700 43.530 5.150 ;
        RECT 39.580 4.550 43.530 4.700 ;
        RECT 43.130 4.400 43.530 4.550 ;
        RECT 45.930 15.450 46.330 15.600 ;
        RECT 45.930 15.300 49.880 15.450 ;
        RECT 45.930 14.850 46.330 15.300 ;
        RECT 45.930 14.700 49.880 14.850 ;
        RECT 45.930 14.250 46.330 14.700 ;
        RECT 45.930 14.100 49.880 14.250 ;
        RECT 45.930 13.650 46.330 14.100 ;
        RECT 45.930 13.500 49.880 13.650 ;
        RECT 45.930 13.050 46.330 13.500 ;
        RECT 45.930 12.900 49.880 13.050 ;
        RECT 45.930 12.450 46.330 12.900 ;
        RECT 45.930 12.300 49.880 12.450 ;
        RECT 45.930 11.850 46.330 12.300 ;
        RECT 45.930 11.700 49.880 11.850 ;
        RECT 45.930 11.250 46.330 11.700 ;
        RECT 45.930 11.100 49.880 11.250 ;
        RECT 45.930 10.650 46.330 11.100 ;
        RECT 45.930 10.500 49.880 10.650 ;
        RECT 45.930 10.200 46.330 10.500 ;
        RECT 50.480 10.200 50.630 18.400 ;
        RECT 51.080 10.200 51.230 18.400 ;
        RECT 51.680 10.200 51.830 18.400 ;
        RECT 52.280 10.200 52.430 18.400 ;
        RECT 52.880 10.200 53.030 18.400 ;
        RECT 53.480 10.200 53.630 18.400 ;
        RECT 54.080 10.200 54.230 18.400 ;
        RECT 45.930 9.800 54.230 10.200 ;
        RECT 45.930 9.500 46.330 9.800 ;
        RECT 45.930 9.350 49.880 9.500 ;
        RECT 45.930 8.900 46.330 9.350 ;
        RECT 45.930 8.750 49.880 8.900 ;
        RECT 45.930 8.300 46.330 8.750 ;
        RECT 45.930 8.150 49.880 8.300 ;
        RECT 45.930 7.700 46.330 8.150 ;
        RECT 45.930 7.550 49.880 7.700 ;
        RECT 45.930 7.100 46.330 7.550 ;
        RECT 45.930 6.950 49.880 7.100 ;
        RECT 45.930 6.500 46.330 6.950 ;
        RECT 45.930 6.350 49.880 6.500 ;
        RECT 45.930 5.900 46.330 6.350 ;
        RECT 45.930 5.750 49.880 5.900 ;
        RECT 45.930 5.300 46.330 5.750 ;
        RECT 45.930 5.150 49.880 5.300 ;
        RECT 45.930 4.700 46.330 5.150 ;
        RECT 45.930 4.550 49.880 4.700 ;
        RECT 45.930 4.400 46.330 4.550 ;
        RECT 43.130 4.100 46.330 4.400 ;
        RECT 39.580 3.950 49.880 4.100 ;
        RECT 43.130 3.500 46.330 3.950 ;
        RECT 39.580 3.350 49.880 3.500 ;
        RECT 43.130 2.900 46.330 3.350 ;
        RECT 39.580 2.750 49.880 2.900 ;
        RECT 43.130 2.300 46.330 2.750 ;
        RECT 39.580 2.150 49.880 2.300 ;
        RECT 43.530 1.200 45.930 2.150 ;
        RECT 50.480 1.600 50.630 9.800 ;
        RECT 51.080 1.600 51.230 9.800 ;
        RECT 51.680 1.600 51.830 9.800 ;
        RECT 52.280 1.600 52.430 9.800 ;
        RECT 52.880 1.600 53.030 9.800 ;
        RECT 53.480 1.600 53.630 9.800 ;
        RECT 54.080 1.600 54.230 9.800 ;
        RECT 55.230 10.200 55.380 18.400 ;
        RECT 55.830 10.200 55.980 18.400 ;
        RECT 56.430 10.200 56.580 18.400 ;
        RECT 57.030 10.200 57.180 18.400 ;
        RECT 57.630 10.200 57.780 18.400 ;
        RECT 58.230 10.200 58.380 18.400 ;
        RECT 58.830 10.200 58.980 18.400 ;
        RECT 63.530 17.850 65.940 18.800 ;
        RECT 59.580 17.700 69.880 17.850 ;
        RECT 63.130 17.250 66.330 17.700 ;
        RECT 59.580 17.100 69.880 17.250 ;
        RECT 63.130 16.650 66.330 17.100 ;
        RECT 59.580 16.500 69.880 16.650 ;
        RECT 63.130 16.050 66.330 16.500 ;
        RECT 59.580 15.900 69.880 16.050 ;
        RECT 63.130 15.600 66.330 15.900 ;
        RECT 63.130 15.450 63.530 15.600 ;
        RECT 59.580 15.300 63.530 15.450 ;
        RECT 63.130 14.850 63.530 15.300 ;
        RECT 59.580 14.700 63.530 14.850 ;
        RECT 63.130 14.250 63.530 14.700 ;
        RECT 59.580 14.100 63.530 14.250 ;
        RECT 63.130 13.650 63.530 14.100 ;
        RECT 59.580 13.500 63.530 13.650 ;
        RECT 63.130 13.050 63.530 13.500 ;
        RECT 59.580 12.900 63.530 13.050 ;
        RECT 63.130 12.450 63.530 12.900 ;
        RECT 59.580 12.300 63.530 12.450 ;
        RECT 63.130 11.850 63.530 12.300 ;
        RECT 59.580 11.700 63.530 11.850 ;
        RECT 63.130 11.250 63.530 11.700 ;
        RECT 59.580 11.100 63.530 11.250 ;
        RECT 63.130 10.650 63.530 11.100 ;
        RECT 59.580 10.500 63.530 10.650 ;
        RECT 63.130 10.200 63.530 10.500 ;
        RECT 55.230 9.800 63.530 10.200 ;
        RECT 55.230 1.600 55.380 9.800 ;
        RECT 55.830 1.600 55.980 9.800 ;
        RECT 56.430 1.600 56.580 9.800 ;
        RECT 57.030 1.600 57.180 9.800 ;
        RECT 57.630 1.600 57.780 9.800 ;
        RECT 58.230 1.600 58.380 9.800 ;
        RECT 58.830 1.600 58.980 9.800 ;
        RECT 63.130 9.500 63.530 9.800 ;
        RECT 59.580 9.350 63.530 9.500 ;
        RECT 63.130 8.900 63.530 9.350 ;
        RECT 59.580 8.750 63.530 8.900 ;
        RECT 63.130 8.300 63.530 8.750 ;
        RECT 59.580 8.150 63.530 8.300 ;
        RECT 63.130 7.700 63.530 8.150 ;
        RECT 59.580 7.550 63.530 7.700 ;
        RECT 63.130 7.100 63.530 7.550 ;
        RECT 59.580 6.950 63.530 7.100 ;
        RECT 63.130 6.500 63.530 6.950 ;
        RECT 59.580 6.350 63.530 6.500 ;
        RECT 63.130 5.900 63.530 6.350 ;
        RECT 59.580 5.750 63.530 5.900 ;
        RECT 63.130 5.300 63.530 5.750 ;
        RECT 59.580 5.150 63.530 5.300 ;
        RECT 63.130 4.700 63.530 5.150 ;
        RECT 59.580 4.550 63.530 4.700 ;
        RECT 63.130 4.400 63.530 4.550 ;
        RECT 65.930 15.450 66.330 15.600 ;
        RECT 65.930 15.300 69.880 15.450 ;
        RECT 65.930 14.850 66.330 15.300 ;
        RECT 65.930 14.700 69.880 14.850 ;
        RECT 65.930 14.250 66.330 14.700 ;
        RECT 65.930 14.100 69.880 14.250 ;
        RECT 65.930 13.650 66.330 14.100 ;
        RECT 65.930 13.500 69.880 13.650 ;
        RECT 65.930 13.050 66.330 13.500 ;
        RECT 65.930 12.900 69.880 13.050 ;
        RECT 65.930 12.450 66.330 12.900 ;
        RECT 65.930 12.300 69.880 12.450 ;
        RECT 65.930 11.850 66.330 12.300 ;
        RECT 65.930 11.700 69.880 11.850 ;
        RECT 65.930 11.250 66.330 11.700 ;
        RECT 65.930 11.100 69.880 11.250 ;
        RECT 65.930 10.650 66.330 11.100 ;
        RECT 65.930 10.500 69.880 10.650 ;
        RECT 65.930 10.200 66.330 10.500 ;
        RECT 70.480 10.200 70.630 18.400 ;
        RECT 71.080 10.200 71.230 18.400 ;
        RECT 71.680 10.200 71.830 18.400 ;
        RECT 72.280 10.200 72.430 18.400 ;
        RECT 72.880 10.200 73.030 18.400 ;
        RECT 73.480 10.200 73.630 18.400 ;
        RECT 74.080 10.200 74.230 18.400 ;
        RECT 65.930 9.800 74.230 10.200 ;
        RECT 65.930 9.500 66.330 9.800 ;
        RECT 65.930 9.350 69.880 9.500 ;
        RECT 65.930 8.900 66.330 9.350 ;
        RECT 65.930 8.750 69.880 8.900 ;
        RECT 65.930 8.300 66.330 8.750 ;
        RECT 65.930 8.150 69.880 8.300 ;
        RECT 65.930 7.700 66.330 8.150 ;
        RECT 65.930 7.550 69.880 7.700 ;
        RECT 65.930 7.100 66.330 7.550 ;
        RECT 65.930 6.950 69.880 7.100 ;
        RECT 65.930 6.500 66.330 6.950 ;
        RECT 65.930 6.350 69.880 6.500 ;
        RECT 65.930 5.900 66.330 6.350 ;
        RECT 65.930 5.750 69.880 5.900 ;
        RECT 65.930 5.300 66.330 5.750 ;
        RECT 65.930 5.150 69.880 5.300 ;
        RECT 65.930 4.700 66.330 5.150 ;
        RECT 65.930 4.550 69.880 4.700 ;
        RECT 65.930 4.400 66.330 4.550 ;
        RECT 63.130 4.100 66.330 4.400 ;
        RECT 59.580 3.950 69.880 4.100 ;
        RECT 63.130 3.500 66.330 3.950 ;
        RECT 59.580 3.350 69.880 3.500 ;
        RECT 63.130 2.900 66.330 3.350 ;
        RECT 59.580 2.750 69.880 2.900 ;
        RECT 63.130 2.300 66.330 2.750 ;
        RECT 59.580 2.150 69.880 2.300 ;
        RECT 63.530 1.200 65.930 2.150 ;
        RECT 70.480 1.600 70.630 9.800 ;
        RECT 71.080 1.600 71.230 9.800 ;
        RECT 71.680 1.600 71.830 9.800 ;
        RECT 72.280 1.600 72.430 9.800 ;
        RECT 72.880 1.600 73.030 9.800 ;
        RECT 73.480 1.600 73.630 9.800 ;
        RECT 74.080 1.600 74.230 9.800 ;
        RECT 75.230 10.200 75.380 18.400 ;
        RECT 75.830 10.200 75.980 18.400 ;
        RECT 76.430 10.200 76.580 18.400 ;
        RECT 77.030 10.200 77.180 18.400 ;
        RECT 77.630 10.200 77.780 18.400 ;
        RECT 78.230 10.200 78.380 18.400 ;
        RECT 78.830 10.200 78.980 18.400 ;
        RECT 83.530 17.850 85.940 18.800 ;
        RECT 79.580 17.700 89.880 17.850 ;
        RECT 83.130 17.250 86.330 17.700 ;
        RECT 79.580 17.100 89.880 17.250 ;
        RECT 83.130 16.650 86.330 17.100 ;
        RECT 79.580 16.500 89.880 16.650 ;
        RECT 83.130 16.050 86.330 16.500 ;
        RECT 79.580 15.900 89.880 16.050 ;
        RECT 83.130 15.600 86.330 15.900 ;
        RECT 83.130 15.450 83.530 15.600 ;
        RECT 79.580 15.300 83.530 15.450 ;
        RECT 83.130 14.850 83.530 15.300 ;
        RECT 79.580 14.700 83.530 14.850 ;
        RECT 83.130 14.250 83.530 14.700 ;
        RECT 79.580 14.100 83.530 14.250 ;
        RECT 83.130 13.650 83.530 14.100 ;
        RECT 79.580 13.500 83.530 13.650 ;
        RECT 83.130 13.050 83.530 13.500 ;
        RECT 79.580 12.900 83.530 13.050 ;
        RECT 83.130 12.450 83.530 12.900 ;
        RECT 79.580 12.300 83.530 12.450 ;
        RECT 83.130 11.850 83.530 12.300 ;
        RECT 79.580 11.700 83.530 11.850 ;
        RECT 83.130 11.250 83.530 11.700 ;
        RECT 79.580 11.100 83.530 11.250 ;
        RECT 83.130 10.650 83.530 11.100 ;
        RECT 79.580 10.500 83.530 10.650 ;
        RECT 83.130 10.200 83.530 10.500 ;
        RECT 75.230 9.800 83.530 10.200 ;
        RECT 75.230 1.600 75.380 9.800 ;
        RECT 75.830 1.600 75.980 9.800 ;
        RECT 76.430 1.600 76.580 9.800 ;
        RECT 77.030 1.600 77.180 9.800 ;
        RECT 77.630 1.600 77.780 9.800 ;
        RECT 78.230 1.600 78.380 9.800 ;
        RECT 78.830 1.600 78.980 9.800 ;
        RECT 83.130 9.500 83.530 9.800 ;
        RECT 79.580 9.350 83.530 9.500 ;
        RECT 83.130 8.900 83.530 9.350 ;
        RECT 79.580 8.750 83.530 8.900 ;
        RECT 83.130 8.300 83.530 8.750 ;
        RECT 79.580 8.150 83.530 8.300 ;
        RECT 83.130 7.700 83.530 8.150 ;
        RECT 79.580 7.550 83.530 7.700 ;
        RECT 83.130 7.100 83.530 7.550 ;
        RECT 79.580 6.950 83.530 7.100 ;
        RECT 83.130 6.500 83.530 6.950 ;
        RECT 79.580 6.350 83.530 6.500 ;
        RECT 83.130 5.900 83.530 6.350 ;
        RECT 79.580 5.750 83.530 5.900 ;
        RECT 83.130 5.300 83.530 5.750 ;
        RECT 79.580 5.150 83.530 5.300 ;
        RECT 83.130 4.700 83.530 5.150 ;
        RECT 79.580 4.550 83.530 4.700 ;
        RECT 83.130 4.400 83.530 4.550 ;
        RECT 85.930 15.450 86.330 15.600 ;
        RECT 85.930 15.300 89.880 15.450 ;
        RECT 85.930 14.850 86.330 15.300 ;
        RECT 85.930 14.700 89.880 14.850 ;
        RECT 85.930 14.250 86.330 14.700 ;
        RECT 85.930 14.100 89.880 14.250 ;
        RECT 85.930 13.650 86.330 14.100 ;
        RECT 85.930 13.500 89.880 13.650 ;
        RECT 85.930 13.050 86.330 13.500 ;
        RECT 85.930 12.900 89.880 13.050 ;
        RECT 85.930 12.450 86.330 12.900 ;
        RECT 85.930 12.300 89.880 12.450 ;
        RECT 85.930 11.850 86.330 12.300 ;
        RECT 85.930 11.700 89.880 11.850 ;
        RECT 85.930 11.250 86.330 11.700 ;
        RECT 85.930 11.100 89.880 11.250 ;
        RECT 85.930 10.650 86.330 11.100 ;
        RECT 85.930 10.500 89.880 10.650 ;
        RECT 85.930 10.200 86.330 10.500 ;
        RECT 90.480 10.200 90.630 18.400 ;
        RECT 91.080 10.200 91.230 18.400 ;
        RECT 91.680 10.200 91.830 18.400 ;
        RECT 92.280 10.200 92.430 18.400 ;
        RECT 92.880 10.200 93.030 18.400 ;
        RECT 93.480 10.200 93.630 18.400 ;
        RECT 94.080 10.200 94.230 18.400 ;
        RECT 85.930 9.800 94.230 10.200 ;
        RECT 85.930 9.500 86.330 9.800 ;
        RECT 85.930 9.350 89.880 9.500 ;
        RECT 85.930 8.900 86.330 9.350 ;
        RECT 85.930 8.750 89.880 8.900 ;
        RECT 85.930 8.300 86.330 8.750 ;
        RECT 85.930 8.150 89.880 8.300 ;
        RECT 85.930 7.700 86.330 8.150 ;
        RECT 85.930 7.550 89.880 7.700 ;
        RECT 85.930 7.100 86.330 7.550 ;
        RECT 85.930 6.950 89.880 7.100 ;
        RECT 85.930 6.500 86.330 6.950 ;
        RECT 85.930 6.350 89.880 6.500 ;
        RECT 85.930 5.900 86.330 6.350 ;
        RECT 85.930 5.750 89.880 5.900 ;
        RECT 85.930 5.300 86.330 5.750 ;
        RECT 85.930 5.150 89.880 5.300 ;
        RECT 85.930 4.700 86.330 5.150 ;
        RECT 85.930 4.550 89.880 4.700 ;
        RECT 85.930 4.400 86.330 4.550 ;
        RECT 83.130 4.100 86.330 4.400 ;
        RECT 79.580 3.950 89.880 4.100 ;
        RECT 83.130 3.500 86.330 3.950 ;
        RECT 79.580 3.350 89.880 3.500 ;
        RECT 83.130 2.900 86.330 3.350 ;
        RECT 79.580 2.750 89.880 2.900 ;
        RECT 83.130 2.300 86.330 2.750 ;
        RECT 79.580 2.150 89.880 2.300 ;
        RECT 83.530 1.200 85.930 2.150 ;
        RECT 90.480 1.600 90.630 9.800 ;
        RECT 91.080 1.600 91.230 9.800 ;
        RECT 91.680 1.600 91.830 9.800 ;
        RECT 92.280 1.600 92.430 9.800 ;
        RECT 92.880 1.600 93.030 9.800 ;
        RECT 93.480 1.600 93.630 9.800 ;
        RECT 94.080 1.600 94.230 9.800 ;
        RECT 95.230 10.200 95.380 18.400 ;
        RECT 95.830 10.200 95.980 18.400 ;
        RECT 96.430 10.200 96.580 18.400 ;
        RECT 97.030 10.200 97.180 18.400 ;
        RECT 97.630 10.200 97.780 18.400 ;
        RECT 98.230 10.200 98.380 18.400 ;
        RECT 98.830 10.200 98.980 18.400 ;
        RECT 103.530 17.850 104.730 18.800 ;
        RECT 99.580 17.700 104.730 17.850 ;
        RECT 103.130 17.250 104.730 17.700 ;
        RECT 99.580 17.100 104.730 17.250 ;
        RECT 103.130 16.650 104.730 17.100 ;
        RECT 99.580 16.500 104.730 16.650 ;
        RECT 103.130 16.050 104.730 16.500 ;
        RECT 99.580 15.900 104.730 16.050 ;
        RECT 105.135 16.035 107.135 17.310 ;
        RECT 103.130 15.600 104.730 15.900 ;
        RECT 103.130 15.450 103.530 15.600 ;
        RECT 99.580 15.300 103.530 15.450 ;
        RECT 103.130 14.850 103.530 15.300 ;
        RECT 99.580 14.700 103.530 14.850 ;
        RECT 103.130 14.250 103.530 14.700 ;
        RECT 99.580 14.100 103.530 14.250 ;
        RECT 103.130 13.650 103.530 14.100 ;
        RECT 99.580 13.500 103.530 13.650 ;
        RECT 103.130 13.050 103.530 13.500 ;
        RECT 99.580 12.900 103.530 13.050 ;
        RECT 103.130 12.450 103.530 12.900 ;
        RECT 99.580 12.300 103.530 12.450 ;
        RECT 103.130 11.850 103.530 12.300 ;
        RECT 99.580 11.700 103.530 11.850 ;
        RECT 103.130 11.250 103.530 11.700 ;
        RECT 99.580 11.100 103.530 11.250 ;
        RECT 103.130 10.650 103.530 11.100 ;
        RECT 99.580 10.500 103.530 10.650 ;
        RECT 103.130 10.200 103.530 10.500 ;
        RECT 95.230 9.800 103.530 10.200 ;
        RECT 95.230 1.600 95.380 9.800 ;
        RECT 95.830 1.600 95.980 9.800 ;
        RECT 96.430 1.600 96.580 9.800 ;
        RECT 97.030 1.600 97.180 9.800 ;
        RECT 97.630 1.600 97.780 9.800 ;
        RECT 98.230 1.600 98.380 9.800 ;
        RECT 98.830 1.600 98.980 9.800 ;
        RECT 103.130 9.500 103.530 9.800 ;
        RECT 99.580 9.350 103.530 9.500 ;
        RECT 103.130 8.900 103.530 9.350 ;
        RECT 99.580 8.750 103.530 8.900 ;
        RECT 103.130 8.300 103.530 8.750 ;
        RECT 99.580 8.150 103.530 8.300 ;
        RECT 103.130 7.700 103.530 8.150 ;
        RECT 99.580 7.550 103.530 7.700 ;
        RECT 103.130 7.100 103.530 7.550 ;
        RECT 99.580 6.950 103.530 7.100 ;
        RECT 103.130 6.500 103.530 6.950 ;
        RECT 99.580 6.350 103.530 6.500 ;
        RECT 103.130 5.900 103.530 6.350 ;
        RECT 99.580 5.750 103.530 5.900 ;
        RECT 103.130 5.300 103.530 5.750 ;
        RECT 99.580 5.150 103.530 5.300 ;
        RECT 103.130 4.700 103.530 5.150 ;
        RECT 99.580 4.550 103.530 4.700 ;
        RECT 103.130 4.400 103.530 4.550 ;
        RECT 103.130 4.100 104.730 4.400 ;
        RECT 99.580 3.950 104.730 4.100 ;
        RECT 103.130 3.500 104.730 3.950 ;
        RECT 99.580 3.350 104.730 3.500 ;
        RECT 103.130 2.900 104.730 3.350 ;
        RECT 99.580 2.750 104.730 2.900 ;
        RECT 103.130 2.300 104.730 2.750 ;
        RECT 99.580 2.150 104.730 2.300 ;
        RECT 103.530 1.200 104.730 2.150 ;
        RECT 105.140 1.820 107.140 3.095 ;
        RECT 4.730 0.000 9.130 1.200 ;
        RECT 20.330 0.000 29.130 1.200 ;
        RECT 40.330 0.000 49.130 1.200 ;
        RECT 60.330 0.000 69.130 1.200 ;
        RECT 80.330 0.000 89.130 1.200 ;
        RECT 100.330 0.000 104.730 1.200 ;
      LAYER via2 ;
        RECT 2.515 376.880 2.875 377.260 ;
        RECT 3.145 376.880 3.505 377.260 ;
        RECT 3.745 376.880 4.105 377.260 ;
        RECT 2.515 376.290 2.875 376.670 ;
        RECT 3.145 376.290 3.505 376.670 ;
        RECT 3.745 376.290 4.105 376.670 ;
        RECT 2.520 374.920 2.880 375.300 ;
        RECT 3.130 374.920 3.490 375.300 ;
        RECT 3.760 374.920 4.120 375.300 ;
        RECT 2.520 374.185 2.880 374.565 ;
        RECT 3.130 374.185 3.490 374.565 ;
        RECT 3.760 374.185 4.120 374.565 ;
        RECT 2.520 373.500 2.880 373.880 ;
        RECT 3.130 373.500 3.490 373.880 ;
        RECT 3.760 373.500 4.120 373.880 ;
        RECT 2.520 366.120 2.880 366.500 ;
        RECT 3.130 366.120 3.490 366.500 ;
        RECT 3.760 366.120 4.120 366.500 ;
        RECT 2.520 365.385 2.880 365.765 ;
        RECT 3.130 365.385 3.490 365.765 ;
        RECT 3.760 365.385 4.120 365.765 ;
        RECT 2.520 364.700 2.880 365.080 ;
        RECT 3.130 364.700 3.490 365.080 ;
        RECT 3.760 364.700 4.120 365.080 ;
        RECT 2.515 363.515 2.875 363.895 ;
        RECT 3.145 363.515 3.505 363.895 ;
        RECT 3.745 363.515 4.105 363.895 ;
        RECT 2.515 362.925 2.875 363.305 ;
        RECT 3.145 362.925 3.505 363.305 ;
        RECT 3.745 362.925 4.105 363.305 ;
        RECT 105.340 377.080 105.700 377.460 ;
        RECT 105.970 377.080 106.330 377.460 ;
        RECT 106.570 377.080 106.930 377.460 ;
        RECT 105.340 376.490 105.700 376.870 ;
        RECT 105.970 376.490 106.330 376.870 ;
        RECT 106.570 376.490 106.930 376.870 ;
        RECT 105.340 363.095 105.700 363.475 ;
        RECT 105.970 363.095 106.330 363.475 ;
        RECT 106.570 363.095 106.930 363.475 ;
        RECT 105.340 362.505 105.700 362.885 ;
        RECT 105.970 362.505 106.330 362.885 ;
        RECT 106.570 362.505 106.930 362.885 ;
        RECT 2.515 356.880 2.875 357.260 ;
        RECT 3.145 356.880 3.505 357.260 ;
        RECT 3.745 356.880 4.105 357.260 ;
        RECT 2.515 356.290 2.875 356.670 ;
        RECT 3.145 356.290 3.505 356.670 ;
        RECT 3.745 356.290 4.105 356.670 ;
        RECT 2.520 354.920 2.880 355.300 ;
        RECT 3.130 354.920 3.490 355.300 ;
        RECT 3.760 354.920 4.120 355.300 ;
        RECT 2.520 354.185 2.880 354.565 ;
        RECT 3.130 354.185 3.490 354.565 ;
        RECT 3.760 354.185 4.120 354.565 ;
        RECT 2.520 353.500 2.880 353.880 ;
        RECT 3.130 353.500 3.490 353.880 ;
        RECT 3.760 353.500 4.120 353.880 ;
        RECT 2.520 346.120 2.880 346.500 ;
        RECT 3.130 346.120 3.490 346.500 ;
        RECT 3.760 346.120 4.120 346.500 ;
        RECT 2.520 345.385 2.880 345.765 ;
        RECT 3.130 345.385 3.490 345.765 ;
        RECT 3.760 345.385 4.120 345.765 ;
        RECT 2.520 344.700 2.880 345.080 ;
        RECT 3.130 344.700 3.490 345.080 ;
        RECT 3.760 344.700 4.120 345.080 ;
        RECT 2.515 343.515 2.875 343.895 ;
        RECT 3.145 343.515 3.505 343.895 ;
        RECT 3.745 343.515 4.105 343.895 ;
        RECT 2.515 342.925 2.875 343.305 ;
        RECT 3.145 342.925 3.505 343.305 ;
        RECT 3.745 342.925 4.105 343.305 ;
        RECT 105.340 357.080 105.700 357.460 ;
        RECT 105.970 357.080 106.330 357.460 ;
        RECT 106.570 357.080 106.930 357.460 ;
        RECT 105.340 356.490 105.700 356.870 ;
        RECT 105.970 356.490 106.330 356.870 ;
        RECT 106.570 356.490 106.930 356.870 ;
        RECT 105.340 343.095 105.700 343.475 ;
        RECT 105.970 343.095 106.330 343.475 ;
        RECT 106.570 343.095 106.930 343.475 ;
        RECT 105.340 342.505 105.700 342.885 ;
        RECT 105.970 342.505 106.330 342.885 ;
        RECT 106.570 342.505 106.930 342.885 ;
        RECT 2.515 336.870 2.875 337.250 ;
        RECT 3.145 336.870 3.505 337.250 ;
        RECT 3.745 336.870 4.105 337.250 ;
        RECT 2.515 336.280 2.875 336.660 ;
        RECT 3.145 336.280 3.505 336.660 ;
        RECT 3.745 336.280 4.105 336.660 ;
        RECT 2.520 334.920 2.880 335.300 ;
        RECT 3.130 334.920 3.490 335.300 ;
        RECT 3.760 334.920 4.120 335.300 ;
        RECT 2.520 334.185 2.880 334.565 ;
        RECT 3.130 334.185 3.490 334.565 ;
        RECT 3.760 334.185 4.120 334.565 ;
        RECT 2.520 333.500 2.880 333.880 ;
        RECT 3.130 333.500 3.490 333.880 ;
        RECT 3.760 333.500 4.120 333.880 ;
        RECT 2.520 326.125 2.880 326.505 ;
        RECT 3.130 326.125 3.490 326.505 ;
        RECT 3.760 326.125 4.120 326.505 ;
        RECT 2.520 325.390 2.880 325.770 ;
        RECT 3.130 325.390 3.490 325.770 ;
        RECT 3.760 325.390 4.120 325.770 ;
        RECT 2.520 324.705 2.880 325.085 ;
        RECT 3.130 324.705 3.490 325.085 ;
        RECT 3.760 324.705 4.120 325.085 ;
        RECT 2.515 323.170 2.875 323.550 ;
        RECT 3.145 323.170 3.505 323.550 ;
        RECT 3.745 323.170 4.105 323.550 ;
        RECT 2.515 322.580 2.875 322.960 ;
        RECT 3.145 322.580 3.505 322.960 ;
        RECT 3.745 322.580 4.105 322.960 ;
        RECT 105.340 337.080 105.700 337.460 ;
        RECT 105.970 337.080 106.330 337.460 ;
        RECT 106.570 337.080 106.930 337.460 ;
        RECT 105.340 336.490 105.700 336.870 ;
        RECT 105.970 336.490 106.330 336.870 ;
        RECT 106.570 336.490 106.930 336.870 ;
        RECT 105.340 323.095 105.700 323.475 ;
        RECT 105.970 323.095 106.330 323.475 ;
        RECT 106.570 323.095 106.930 323.475 ;
        RECT 105.340 322.505 105.700 322.885 ;
        RECT 105.970 322.505 106.330 322.885 ;
        RECT 106.570 322.505 106.930 322.885 ;
        RECT 2.515 317.280 2.875 317.660 ;
        RECT 3.145 317.280 3.505 317.660 ;
        RECT 3.745 317.280 4.105 317.660 ;
        RECT 2.515 316.690 2.875 317.070 ;
        RECT 3.145 316.690 3.505 317.070 ;
        RECT 3.745 316.690 4.105 317.070 ;
        RECT 2.520 314.920 2.880 315.300 ;
        RECT 3.130 314.920 3.490 315.300 ;
        RECT 3.760 314.920 4.120 315.300 ;
        RECT 2.520 314.185 2.880 314.565 ;
        RECT 3.130 314.185 3.490 314.565 ;
        RECT 3.760 314.185 4.120 314.565 ;
        RECT 2.520 313.500 2.880 313.880 ;
        RECT 3.130 313.500 3.490 313.880 ;
        RECT 3.760 313.500 4.120 313.880 ;
        RECT 2.520 306.125 2.880 306.505 ;
        RECT 3.130 306.125 3.490 306.505 ;
        RECT 3.760 306.125 4.120 306.505 ;
        RECT 2.520 305.390 2.880 305.770 ;
        RECT 3.130 305.390 3.490 305.770 ;
        RECT 3.760 305.390 4.120 305.770 ;
        RECT 2.520 304.705 2.880 305.085 ;
        RECT 3.130 304.705 3.490 305.085 ;
        RECT 3.760 304.705 4.120 305.085 ;
        RECT 2.515 303.040 2.875 303.420 ;
        RECT 3.145 303.040 3.505 303.420 ;
        RECT 3.745 303.040 4.105 303.420 ;
        RECT 2.515 302.450 2.875 302.830 ;
        RECT 3.145 302.450 3.505 302.830 ;
        RECT 3.745 302.450 4.105 302.830 ;
        RECT 105.340 317.080 105.700 317.460 ;
        RECT 105.970 317.080 106.330 317.460 ;
        RECT 106.570 317.080 106.930 317.460 ;
        RECT 105.340 316.490 105.700 316.870 ;
        RECT 105.970 316.490 106.330 316.870 ;
        RECT 106.570 316.490 106.930 316.870 ;
        RECT 105.340 303.095 105.700 303.475 ;
        RECT 105.970 303.095 106.330 303.475 ;
        RECT 106.570 303.095 106.930 303.475 ;
        RECT 105.340 302.505 105.700 302.885 ;
        RECT 105.970 302.505 106.330 302.885 ;
        RECT 106.570 302.505 106.930 302.885 ;
        RECT 2.515 297.025 2.875 297.405 ;
        RECT 3.145 297.025 3.505 297.405 ;
        RECT 3.745 297.025 4.105 297.405 ;
        RECT 2.515 296.435 2.875 296.815 ;
        RECT 3.145 296.435 3.505 296.815 ;
        RECT 3.745 296.435 4.105 296.815 ;
        RECT 2.520 294.920 2.880 295.300 ;
        RECT 3.130 294.920 3.490 295.300 ;
        RECT 3.760 294.920 4.120 295.300 ;
        RECT 2.520 294.185 2.880 294.565 ;
        RECT 3.130 294.185 3.490 294.565 ;
        RECT 3.760 294.185 4.120 294.565 ;
        RECT 2.520 293.500 2.880 293.880 ;
        RECT 3.130 293.500 3.490 293.880 ;
        RECT 3.760 293.500 4.120 293.880 ;
        RECT 2.520 286.115 2.880 286.495 ;
        RECT 3.130 286.115 3.490 286.495 ;
        RECT 3.760 286.115 4.120 286.495 ;
        RECT 2.520 285.380 2.880 285.760 ;
        RECT 3.130 285.380 3.490 285.760 ;
        RECT 3.760 285.380 4.120 285.760 ;
        RECT 2.520 284.695 2.880 285.075 ;
        RECT 3.130 284.695 3.490 285.075 ;
        RECT 3.760 284.695 4.120 285.075 ;
        RECT 2.515 283.140 2.875 283.520 ;
        RECT 3.145 283.140 3.505 283.520 ;
        RECT 3.745 283.140 4.105 283.520 ;
        RECT 2.515 282.550 2.875 282.930 ;
        RECT 3.145 282.550 3.505 282.930 ;
        RECT 3.745 282.550 4.105 282.930 ;
        RECT 105.340 297.350 105.700 297.730 ;
        RECT 105.970 297.350 106.330 297.730 ;
        RECT 106.570 297.350 106.930 297.730 ;
        RECT 105.340 296.760 105.700 297.140 ;
        RECT 105.970 296.760 106.330 297.140 ;
        RECT 106.570 296.760 106.930 297.140 ;
        RECT 105.340 282.770 105.700 283.150 ;
        RECT 105.970 282.770 106.330 283.150 ;
        RECT 106.570 282.770 106.930 283.150 ;
        RECT 105.340 282.180 105.700 282.560 ;
        RECT 105.970 282.180 106.330 282.560 ;
        RECT 106.570 282.180 106.930 282.560 ;
        RECT 2.515 277.105 2.875 277.485 ;
        RECT 3.145 277.105 3.505 277.485 ;
        RECT 3.745 277.105 4.105 277.485 ;
        RECT 2.515 276.515 2.875 276.895 ;
        RECT 3.145 276.515 3.505 276.895 ;
        RECT 3.745 276.515 4.105 276.895 ;
        RECT 2.520 274.920 2.880 275.300 ;
        RECT 3.130 274.920 3.490 275.300 ;
        RECT 3.760 274.920 4.120 275.300 ;
        RECT 2.520 274.185 2.880 274.565 ;
        RECT 3.130 274.185 3.490 274.565 ;
        RECT 3.760 274.185 4.120 274.565 ;
        RECT 2.520 273.500 2.880 273.880 ;
        RECT 3.130 273.500 3.490 273.880 ;
        RECT 3.760 273.500 4.120 273.880 ;
        RECT 2.520 266.125 2.880 266.505 ;
        RECT 3.130 266.125 3.490 266.505 ;
        RECT 3.760 266.125 4.120 266.505 ;
        RECT 2.520 265.390 2.880 265.770 ;
        RECT 3.130 265.390 3.490 265.770 ;
        RECT 3.760 265.390 4.120 265.770 ;
        RECT 2.520 264.705 2.880 265.085 ;
        RECT 3.130 264.705 3.490 265.085 ;
        RECT 3.760 264.705 4.120 265.085 ;
        RECT 2.515 263.275 2.875 263.655 ;
        RECT 3.145 263.275 3.505 263.655 ;
        RECT 3.745 263.275 4.105 263.655 ;
        RECT 2.515 262.685 2.875 263.065 ;
        RECT 3.145 262.685 3.505 263.065 ;
        RECT 3.745 262.685 4.105 263.065 ;
        RECT 105.340 276.855 105.700 277.235 ;
        RECT 105.970 276.855 106.330 277.235 ;
        RECT 106.570 276.855 106.930 277.235 ;
        RECT 105.340 276.265 105.700 276.645 ;
        RECT 105.970 276.265 106.330 276.645 ;
        RECT 106.570 276.265 106.930 276.645 ;
        RECT 105.340 262.495 105.700 262.875 ;
        RECT 105.970 262.495 106.330 262.875 ;
        RECT 106.570 262.495 106.930 262.875 ;
        RECT 105.340 261.905 105.700 262.285 ;
        RECT 105.970 261.905 106.330 262.285 ;
        RECT 106.570 261.905 106.930 262.285 ;
        RECT 2.515 257.340 2.875 257.720 ;
        RECT 3.145 257.340 3.505 257.720 ;
        RECT 3.745 257.340 4.105 257.720 ;
        RECT 2.515 256.750 2.875 257.130 ;
        RECT 3.145 256.750 3.505 257.130 ;
        RECT 3.745 256.750 4.105 257.130 ;
        RECT 2.520 254.920 2.880 255.300 ;
        RECT 3.130 254.920 3.490 255.300 ;
        RECT 3.760 254.920 4.120 255.300 ;
        RECT 2.520 254.185 2.880 254.565 ;
        RECT 3.130 254.185 3.490 254.565 ;
        RECT 3.760 254.185 4.120 254.565 ;
        RECT 2.520 253.500 2.880 253.880 ;
        RECT 3.130 253.500 3.490 253.880 ;
        RECT 3.760 253.500 4.120 253.880 ;
        RECT 2.520 246.125 2.880 246.505 ;
        RECT 3.130 246.125 3.490 246.505 ;
        RECT 3.760 246.125 4.120 246.505 ;
        RECT 2.520 245.390 2.880 245.770 ;
        RECT 3.130 245.390 3.490 245.770 ;
        RECT 3.760 245.390 4.120 245.770 ;
        RECT 2.520 244.705 2.880 245.085 ;
        RECT 3.130 244.705 3.490 245.085 ;
        RECT 3.760 244.705 4.120 245.085 ;
        RECT 2.515 243.230 2.875 243.610 ;
        RECT 3.145 243.230 3.505 243.610 ;
        RECT 3.745 243.230 4.105 243.610 ;
        RECT 2.515 242.640 2.875 243.020 ;
        RECT 3.145 242.640 3.505 243.020 ;
        RECT 3.745 242.640 4.105 243.020 ;
        RECT 105.340 256.820 105.700 257.200 ;
        RECT 105.970 256.820 106.330 257.200 ;
        RECT 106.570 256.820 106.930 257.200 ;
        RECT 105.340 256.230 105.700 256.610 ;
        RECT 105.970 256.230 106.330 256.610 ;
        RECT 106.570 256.230 106.930 256.610 ;
        RECT 105.340 243.025 105.700 243.405 ;
        RECT 105.970 243.025 106.330 243.405 ;
        RECT 106.570 243.025 106.930 243.405 ;
        RECT 105.340 242.435 105.700 242.815 ;
        RECT 105.970 242.435 106.330 242.815 ;
        RECT 106.570 242.435 106.930 242.815 ;
        RECT 2.515 237.465 2.875 237.845 ;
        RECT 3.145 237.465 3.505 237.845 ;
        RECT 3.745 237.465 4.105 237.845 ;
        RECT 2.515 236.875 2.875 237.255 ;
        RECT 3.145 236.875 3.505 237.255 ;
        RECT 3.745 236.875 4.105 237.255 ;
        RECT 2.520 234.920 2.880 235.300 ;
        RECT 3.130 234.920 3.490 235.300 ;
        RECT 3.760 234.920 4.120 235.300 ;
        RECT 2.520 234.185 2.880 234.565 ;
        RECT 3.130 234.185 3.490 234.565 ;
        RECT 3.760 234.185 4.120 234.565 ;
        RECT 2.520 233.500 2.880 233.880 ;
        RECT 3.130 233.500 3.490 233.880 ;
        RECT 3.760 233.500 4.120 233.880 ;
        RECT 2.520 226.120 2.880 226.500 ;
        RECT 3.130 226.120 3.490 226.500 ;
        RECT 3.760 226.120 4.120 226.500 ;
        RECT 2.520 225.385 2.880 225.765 ;
        RECT 3.130 225.385 3.490 225.765 ;
        RECT 3.760 225.385 4.120 225.765 ;
        RECT 2.520 224.700 2.880 225.080 ;
        RECT 3.130 224.700 3.490 225.080 ;
        RECT 3.760 224.700 4.120 225.080 ;
        RECT 2.515 222.165 2.875 222.545 ;
        RECT 3.145 222.165 3.505 222.545 ;
        RECT 3.745 222.165 4.105 222.545 ;
        RECT 2.515 221.575 2.875 221.955 ;
        RECT 3.145 221.575 3.505 221.955 ;
        RECT 3.745 221.575 4.105 221.955 ;
        RECT 105.340 237.260 105.700 237.640 ;
        RECT 105.970 237.260 106.330 237.640 ;
        RECT 106.570 237.260 106.930 237.640 ;
        RECT 105.340 236.670 105.700 237.050 ;
        RECT 105.970 236.670 106.330 237.050 ;
        RECT 106.570 236.670 106.930 237.050 ;
        RECT 105.340 221.680 105.700 222.060 ;
        RECT 105.970 221.680 106.330 222.060 ;
        RECT 106.570 221.680 106.930 222.060 ;
        RECT 105.340 221.090 105.700 221.470 ;
        RECT 105.970 221.090 106.330 221.470 ;
        RECT 106.570 221.090 106.930 221.470 ;
        RECT 2.395 195.260 2.805 195.650 ;
        RECT 2.965 195.260 3.375 195.650 ;
        RECT 3.535 195.260 3.945 195.650 ;
        RECT 2.395 189.820 2.805 190.210 ;
        RECT 2.965 189.820 3.375 190.210 ;
        RECT 3.535 189.820 3.945 190.210 ;
        RECT 2.395 184.380 2.805 184.770 ;
        RECT 2.965 184.380 3.375 184.770 ;
        RECT 3.535 184.380 3.945 184.770 ;
        RECT 105.305 180.460 105.705 180.860 ;
        RECT 105.930 180.460 106.330 180.860 ;
        RECT 106.555 180.460 106.955 180.860 ;
        RECT 105.300 179.860 105.700 180.260 ;
        RECT 105.925 179.860 106.325 180.260 ;
        RECT 106.550 179.860 106.950 180.260 ;
        RECT 105.345 177.580 105.705 177.960 ;
        RECT 105.955 177.580 106.315 177.960 ;
        RECT 106.585 177.580 106.945 177.960 ;
        RECT 105.345 176.845 105.705 177.225 ;
        RECT 105.955 176.845 106.315 177.225 ;
        RECT 106.585 176.845 106.945 177.225 ;
        RECT 105.345 176.160 105.705 176.540 ;
        RECT 105.955 176.160 106.315 176.540 ;
        RECT 106.585 176.160 106.945 176.540 ;
        RECT 105.345 168.780 105.705 169.160 ;
        RECT 105.955 168.780 106.315 169.160 ;
        RECT 106.585 168.780 106.945 169.160 ;
        RECT 105.345 168.045 105.705 168.425 ;
        RECT 105.955 168.045 106.315 168.425 ;
        RECT 106.585 168.045 106.945 168.425 ;
        RECT 105.345 167.360 105.705 167.740 ;
        RECT 105.955 167.360 106.315 167.740 ;
        RECT 106.585 167.360 106.945 167.740 ;
        RECT 105.300 165.185 105.700 165.585 ;
        RECT 105.925 165.185 106.325 165.585 ;
        RECT 106.550 165.185 106.950 165.585 ;
        RECT 105.295 164.585 105.695 164.985 ;
        RECT 105.920 164.585 106.320 164.985 ;
        RECT 106.545 164.585 106.945 164.985 ;
        RECT 2.515 161.130 2.875 161.510 ;
        RECT 3.145 161.130 3.505 161.510 ;
        RECT 3.745 161.130 4.105 161.510 ;
        RECT 2.515 160.540 2.875 160.920 ;
        RECT 3.145 160.540 3.505 160.920 ;
        RECT 3.745 160.540 4.105 160.920 ;
        RECT 105.340 161.130 105.700 161.510 ;
        RECT 105.970 161.130 106.330 161.510 ;
        RECT 106.570 161.130 106.930 161.510 ;
        RECT 105.340 160.540 105.700 160.920 ;
        RECT 105.970 160.540 106.330 160.920 ;
        RECT 106.570 160.540 106.930 160.920 ;
        RECT 2.515 157.220 2.875 157.600 ;
        RECT 3.145 157.220 3.505 157.600 ;
        RECT 3.745 157.220 4.105 157.600 ;
        RECT 2.515 156.630 2.875 157.010 ;
        RECT 3.145 156.630 3.505 157.010 ;
        RECT 3.745 156.630 4.105 157.010 ;
        RECT 2.520 154.925 2.880 155.305 ;
        RECT 3.130 154.925 3.490 155.305 ;
        RECT 3.760 154.925 4.120 155.305 ;
        RECT 2.520 154.190 2.880 154.570 ;
        RECT 3.130 154.190 3.490 154.570 ;
        RECT 3.760 154.190 4.120 154.570 ;
        RECT 2.520 153.505 2.880 153.885 ;
        RECT 3.130 153.505 3.490 153.885 ;
        RECT 3.760 153.505 4.120 153.885 ;
        RECT 2.520 146.090 2.880 146.470 ;
        RECT 3.130 146.090 3.490 146.470 ;
        RECT 3.760 146.090 4.120 146.470 ;
        RECT 2.520 145.355 2.880 145.735 ;
        RECT 3.130 145.355 3.490 145.735 ;
        RECT 3.760 145.355 4.120 145.735 ;
        RECT 2.520 144.670 2.880 145.050 ;
        RECT 3.130 144.670 3.490 145.050 ;
        RECT 3.760 144.670 4.120 145.050 ;
        RECT 2.515 142.660 2.875 143.040 ;
        RECT 3.145 142.660 3.505 143.040 ;
        RECT 3.745 142.660 4.105 143.040 ;
        RECT 2.515 142.070 2.875 142.450 ;
        RECT 3.145 142.070 3.505 142.450 ;
        RECT 3.745 142.070 4.105 142.450 ;
        RECT 105.340 157.220 105.700 157.600 ;
        RECT 105.970 157.220 106.330 157.600 ;
        RECT 106.570 157.220 106.930 157.600 ;
        RECT 105.340 156.630 105.700 157.010 ;
        RECT 105.970 156.630 106.330 157.010 ;
        RECT 106.570 156.630 106.930 157.010 ;
        RECT 105.340 142.415 105.700 142.795 ;
        RECT 105.970 142.415 106.330 142.795 ;
        RECT 106.570 142.415 106.930 142.795 ;
        RECT 105.340 141.825 105.700 142.205 ;
        RECT 105.970 141.825 106.330 142.205 ;
        RECT 106.570 141.825 106.930 142.205 ;
        RECT 2.515 137.640 2.875 138.020 ;
        RECT 3.145 137.640 3.505 138.020 ;
        RECT 3.745 137.640 4.105 138.020 ;
        RECT 2.515 137.050 2.875 137.430 ;
        RECT 3.145 137.050 3.505 137.430 ;
        RECT 3.745 137.050 4.105 137.430 ;
        RECT 2.520 134.920 2.880 135.300 ;
        RECT 3.130 134.920 3.490 135.300 ;
        RECT 3.760 134.920 4.120 135.300 ;
        RECT 2.520 134.185 2.880 134.565 ;
        RECT 3.130 134.185 3.490 134.565 ;
        RECT 3.760 134.185 4.120 134.565 ;
        RECT 2.520 133.500 2.880 133.880 ;
        RECT 3.130 133.500 3.490 133.880 ;
        RECT 3.760 133.500 4.120 133.880 ;
        RECT 2.520 126.120 2.880 126.500 ;
        RECT 3.130 126.120 3.490 126.500 ;
        RECT 3.760 126.120 4.120 126.500 ;
        RECT 2.520 125.385 2.880 125.765 ;
        RECT 3.130 125.385 3.490 125.765 ;
        RECT 3.760 125.385 4.120 125.765 ;
        RECT 2.520 124.700 2.880 125.080 ;
        RECT 3.130 124.700 3.490 125.080 ;
        RECT 3.760 124.700 4.120 125.080 ;
        RECT 2.515 122.750 2.875 123.130 ;
        RECT 3.145 122.750 3.505 123.130 ;
        RECT 3.745 122.750 4.105 123.130 ;
        RECT 2.515 122.160 2.875 122.540 ;
        RECT 3.145 122.160 3.505 122.540 ;
        RECT 3.745 122.160 4.105 122.540 ;
        RECT 105.340 136.830 105.700 137.210 ;
        RECT 105.970 136.830 106.330 137.210 ;
        RECT 106.570 136.830 106.930 137.210 ;
        RECT 105.340 136.240 105.700 136.620 ;
        RECT 105.970 136.240 106.330 136.620 ;
        RECT 106.570 136.240 106.930 136.620 ;
        RECT 105.340 122.615 105.700 122.995 ;
        RECT 105.970 122.615 106.330 122.995 ;
        RECT 106.570 122.615 106.930 122.995 ;
        RECT 105.340 122.025 105.700 122.405 ;
        RECT 105.970 122.025 106.330 122.405 ;
        RECT 106.570 122.025 106.930 122.405 ;
        RECT 2.515 117.340 2.875 117.720 ;
        RECT 3.145 117.340 3.505 117.720 ;
        RECT 3.745 117.340 4.105 117.720 ;
        RECT 2.515 116.750 2.875 117.130 ;
        RECT 3.145 116.750 3.505 117.130 ;
        RECT 3.745 116.750 4.105 117.130 ;
        RECT 2.520 114.920 2.880 115.300 ;
        RECT 3.130 114.920 3.490 115.300 ;
        RECT 3.760 114.920 4.120 115.300 ;
        RECT 2.520 114.185 2.880 114.565 ;
        RECT 3.130 114.185 3.490 114.565 ;
        RECT 3.760 114.185 4.120 114.565 ;
        RECT 2.520 113.500 2.880 113.880 ;
        RECT 3.130 113.500 3.490 113.880 ;
        RECT 3.760 113.500 4.120 113.880 ;
        RECT 2.520 106.125 2.880 106.505 ;
        RECT 3.130 106.125 3.490 106.505 ;
        RECT 3.760 106.125 4.120 106.505 ;
        RECT 2.520 105.390 2.880 105.770 ;
        RECT 3.130 105.390 3.490 105.770 ;
        RECT 3.760 105.390 4.120 105.770 ;
        RECT 2.520 104.705 2.880 105.085 ;
        RECT 3.130 104.705 3.490 105.085 ;
        RECT 3.760 104.705 4.120 105.085 ;
        RECT 2.515 102.965 2.875 103.345 ;
        RECT 3.145 102.965 3.505 103.345 ;
        RECT 3.745 102.965 4.105 103.345 ;
        RECT 2.515 102.375 2.875 102.755 ;
        RECT 3.145 102.375 3.505 102.755 ;
        RECT 3.745 102.375 4.105 102.755 ;
        RECT 105.340 116.740 105.700 117.120 ;
        RECT 105.970 116.740 106.330 117.120 ;
        RECT 106.570 116.740 106.930 117.120 ;
        RECT 105.340 116.150 105.700 116.530 ;
        RECT 105.970 116.150 106.330 116.530 ;
        RECT 106.570 116.150 106.930 116.530 ;
        RECT 105.340 102.535 105.700 102.915 ;
        RECT 105.970 102.535 106.330 102.915 ;
        RECT 106.570 102.535 106.930 102.915 ;
        RECT 105.340 101.945 105.700 102.325 ;
        RECT 105.970 101.945 106.330 102.325 ;
        RECT 106.570 101.945 106.930 102.325 ;
        RECT 2.515 97.460 2.875 97.840 ;
        RECT 3.145 97.460 3.505 97.840 ;
        RECT 3.745 97.460 4.105 97.840 ;
        RECT 2.515 96.870 2.875 97.250 ;
        RECT 3.145 96.870 3.505 97.250 ;
        RECT 3.745 96.870 4.105 97.250 ;
        RECT 2.520 94.920 2.880 95.300 ;
        RECT 3.130 94.920 3.490 95.300 ;
        RECT 3.760 94.920 4.120 95.300 ;
        RECT 2.520 94.185 2.880 94.565 ;
        RECT 3.130 94.185 3.490 94.565 ;
        RECT 3.760 94.185 4.120 94.565 ;
        RECT 2.520 93.500 2.880 93.880 ;
        RECT 3.130 93.500 3.490 93.880 ;
        RECT 3.760 93.500 4.120 93.880 ;
        RECT 2.520 86.120 2.880 86.500 ;
        RECT 3.130 86.120 3.490 86.500 ;
        RECT 3.760 86.120 4.120 86.500 ;
        RECT 2.520 85.385 2.880 85.765 ;
        RECT 3.130 85.385 3.490 85.765 ;
        RECT 3.760 85.385 4.120 85.765 ;
        RECT 2.520 84.700 2.880 85.080 ;
        RECT 3.130 84.700 3.490 85.080 ;
        RECT 3.760 84.700 4.120 85.080 ;
        RECT 2.515 83.130 2.875 83.510 ;
        RECT 3.145 83.130 3.505 83.510 ;
        RECT 3.745 83.130 4.105 83.510 ;
        RECT 2.515 82.540 2.875 82.920 ;
        RECT 3.145 82.540 3.505 82.920 ;
        RECT 3.745 82.540 4.105 82.920 ;
        RECT 105.340 96.680 105.700 97.060 ;
        RECT 105.970 96.680 106.330 97.060 ;
        RECT 106.570 96.680 106.930 97.060 ;
        RECT 105.340 96.090 105.700 96.470 ;
        RECT 105.970 96.090 106.330 96.470 ;
        RECT 106.570 96.090 106.930 96.470 ;
        RECT 105.340 82.875 105.700 83.255 ;
        RECT 105.970 82.875 106.330 83.255 ;
        RECT 106.570 82.875 106.930 83.255 ;
        RECT 105.340 82.285 105.700 82.665 ;
        RECT 105.970 82.285 106.330 82.665 ;
        RECT 106.570 82.285 106.930 82.665 ;
        RECT 2.515 77.050 2.875 77.430 ;
        RECT 3.145 77.050 3.505 77.430 ;
        RECT 3.745 77.050 4.105 77.430 ;
        RECT 2.515 76.460 2.875 76.840 ;
        RECT 3.145 76.460 3.505 76.840 ;
        RECT 3.745 76.460 4.105 76.840 ;
        RECT 2.520 74.920 2.880 75.300 ;
        RECT 3.130 74.920 3.490 75.300 ;
        RECT 3.760 74.920 4.120 75.300 ;
        RECT 2.520 74.185 2.880 74.565 ;
        RECT 3.130 74.185 3.490 74.565 ;
        RECT 3.760 74.185 4.120 74.565 ;
        RECT 2.520 73.500 2.880 73.880 ;
        RECT 3.130 73.500 3.490 73.880 ;
        RECT 3.760 73.500 4.120 73.880 ;
        RECT 2.520 66.120 2.880 66.500 ;
        RECT 3.130 66.120 3.490 66.500 ;
        RECT 3.760 66.120 4.120 66.500 ;
        RECT 2.520 65.385 2.880 65.765 ;
        RECT 3.130 65.385 3.490 65.765 ;
        RECT 3.760 65.385 4.120 65.765 ;
        RECT 2.520 64.700 2.880 65.080 ;
        RECT 3.130 64.700 3.490 65.080 ;
        RECT 3.760 64.700 4.120 65.080 ;
        RECT 2.515 62.725 2.875 63.105 ;
        RECT 3.145 62.725 3.505 63.105 ;
        RECT 3.745 62.725 4.105 63.105 ;
        RECT 2.515 62.135 2.875 62.515 ;
        RECT 3.145 62.135 3.505 62.515 ;
        RECT 3.745 62.135 4.105 62.515 ;
        RECT 105.340 76.805 105.700 77.185 ;
        RECT 105.970 76.805 106.330 77.185 ;
        RECT 106.570 76.805 106.930 77.185 ;
        RECT 105.340 76.215 105.700 76.595 ;
        RECT 105.970 76.215 106.330 76.595 ;
        RECT 106.570 76.215 106.930 76.595 ;
        RECT 105.340 62.590 105.700 62.970 ;
        RECT 105.970 62.590 106.330 62.970 ;
        RECT 106.570 62.590 106.930 62.970 ;
        RECT 105.340 62.000 105.700 62.380 ;
        RECT 105.970 62.000 106.330 62.380 ;
        RECT 106.570 62.000 106.930 62.380 ;
        RECT 2.515 57.115 2.875 57.495 ;
        RECT 3.145 57.115 3.505 57.495 ;
        RECT 3.745 57.115 4.105 57.495 ;
        RECT 2.515 56.525 2.875 56.905 ;
        RECT 3.145 56.525 3.505 56.905 ;
        RECT 3.745 56.525 4.105 56.905 ;
        RECT 2.520 54.925 2.880 55.305 ;
        RECT 3.130 54.925 3.490 55.305 ;
        RECT 3.760 54.925 4.120 55.305 ;
        RECT 2.520 54.190 2.880 54.570 ;
        RECT 3.130 54.190 3.490 54.570 ;
        RECT 3.760 54.190 4.120 54.570 ;
        RECT 2.520 53.505 2.880 53.885 ;
        RECT 3.130 53.505 3.490 53.885 ;
        RECT 3.760 53.505 4.120 53.885 ;
        RECT 2.520 46.115 2.880 46.495 ;
        RECT 3.130 46.115 3.490 46.495 ;
        RECT 3.760 46.115 4.120 46.495 ;
        RECT 2.520 45.380 2.880 45.760 ;
        RECT 3.130 45.380 3.490 45.760 ;
        RECT 3.760 45.380 4.120 45.760 ;
        RECT 2.520 44.695 2.880 45.075 ;
        RECT 3.130 44.695 3.490 45.075 ;
        RECT 3.760 44.695 4.120 45.075 ;
        RECT 2.515 42.815 2.875 43.195 ;
        RECT 3.145 42.815 3.505 43.195 ;
        RECT 3.745 42.815 4.105 43.195 ;
        RECT 2.515 42.225 2.875 42.605 ;
        RECT 3.145 42.225 3.505 42.605 ;
        RECT 3.745 42.225 4.105 42.605 ;
        RECT 105.340 56.805 105.700 57.185 ;
        RECT 105.970 56.805 106.330 57.185 ;
        RECT 106.570 56.805 106.930 57.185 ;
        RECT 105.340 56.215 105.700 56.595 ;
        RECT 105.970 56.215 106.330 56.595 ;
        RECT 106.570 56.215 106.930 56.595 ;
        RECT 105.340 42.590 105.700 42.970 ;
        RECT 105.970 42.590 106.330 42.970 ;
        RECT 106.570 42.590 106.930 42.970 ;
        RECT 105.340 42.000 105.700 42.380 ;
        RECT 105.970 42.000 106.330 42.380 ;
        RECT 106.570 42.000 106.930 42.380 ;
        RECT 2.515 37.260 2.875 37.640 ;
        RECT 3.145 37.260 3.505 37.640 ;
        RECT 3.745 37.260 4.105 37.640 ;
        RECT 2.515 36.670 2.875 37.050 ;
        RECT 3.145 36.670 3.505 37.050 ;
        RECT 3.745 36.670 4.105 37.050 ;
        RECT 2.520 34.925 2.880 35.305 ;
        RECT 3.130 34.925 3.490 35.305 ;
        RECT 3.760 34.925 4.120 35.305 ;
        RECT 2.520 34.190 2.880 34.570 ;
        RECT 3.130 34.190 3.490 34.570 ;
        RECT 3.760 34.190 4.120 34.570 ;
        RECT 2.520 33.505 2.880 33.885 ;
        RECT 3.130 33.505 3.490 33.885 ;
        RECT 3.760 33.505 4.120 33.885 ;
        RECT 2.520 26.120 2.880 26.500 ;
        RECT 3.130 26.120 3.490 26.500 ;
        RECT 3.760 26.120 4.120 26.500 ;
        RECT 2.520 25.385 2.880 25.765 ;
        RECT 3.130 25.385 3.490 25.765 ;
        RECT 3.760 25.385 4.120 25.765 ;
        RECT 2.520 24.700 2.880 25.080 ;
        RECT 3.130 24.700 3.490 25.080 ;
        RECT 3.760 24.700 4.120 25.080 ;
        RECT 2.515 23.145 2.875 23.525 ;
        RECT 3.145 23.145 3.505 23.525 ;
        RECT 3.745 23.145 4.105 23.525 ;
        RECT 2.515 22.555 2.875 22.935 ;
        RECT 3.145 22.555 3.505 22.935 ;
        RECT 3.745 22.555 4.105 22.935 ;
        RECT 105.340 36.805 105.700 37.185 ;
        RECT 105.970 36.805 106.330 37.185 ;
        RECT 106.570 36.805 106.930 37.185 ;
        RECT 105.340 36.215 105.700 36.595 ;
        RECT 105.970 36.215 106.330 36.595 ;
        RECT 106.570 36.215 106.930 36.595 ;
        RECT 105.340 22.590 105.700 22.970 ;
        RECT 105.970 22.590 106.330 22.970 ;
        RECT 106.570 22.590 106.930 22.970 ;
        RECT 105.340 22.000 105.700 22.380 ;
        RECT 105.970 22.000 106.330 22.380 ;
        RECT 106.570 22.000 106.930 22.380 ;
        RECT 2.515 17.260 2.875 17.640 ;
        RECT 3.145 17.260 3.505 17.640 ;
        RECT 3.745 17.260 4.105 17.640 ;
        RECT 2.515 16.670 2.875 17.050 ;
        RECT 3.145 16.670 3.505 17.050 ;
        RECT 3.745 16.670 4.105 17.050 ;
        RECT 2.520 14.925 2.880 15.305 ;
        RECT 3.130 14.925 3.490 15.305 ;
        RECT 3.760 14.925 4.120 15.305 ;
        RECT 2.520 14.190 2.880 14.570 ;
        RECT 3.130 14.190 3.490 14.570 ;
        RECT 3.760 14.190 4.120 14.570 ;
        RECT 2.520 13.505 2.880 13.885 ;
        RECT 3.130 13.505 3.490 13.885 ;
        RECT 3.760 13.505 4.120 13.885 ;
        RECT 2.520 6.120 2.880 6.500 ;
        RECT 3.130 6.120 3.490 6.500 ;
        RECT 3.760 6.120 4.120 6.500 ;
        RECT 2.520 5.385 2.880 5.765 ;
        RECT 3.130 5.385 3.490 5.765 ;
        RECT 3.760 5.385 4.120 5.765 ;
        RECT 2.520 4.700 2.880 5.080 ;
        RECT 3.130 4.700 3.490 5.080 ;
        RECT 3.760 4.700 4.120 5.080 ;
        RECT 2.515 3.145 2.875 3.525 ;
        RECT 3.145 3.145 3.505 3.525 ;
        RECT 3.745 3.145 4.105 3.525 ;
        RECT 2.515 2.555 2.875 2.935 ;
        RECT 3.145 2.555 3.505 2.935 ;
        RECT 3.745 2.555 4.105 2.935 ;
        RECT 105.340 16.805 105.700 17.185 ;
        RECT 105.970 16.805 106.330 17.185 ;
        RECT 106.570 16.805 106.930 17.185 ;
        RECT 105.340 16.215 105.700 16.595 ;
        RECT 105.970 16.215 106.330 16.595 ;
        RECT 106.570 16.215 106.930 16.595 ;
        RECT 105.340 2.590 105.700 2.970 ;
        RECT 105.970 2.590 106.330 2.970 ;
        RECT 106.570 2.590 106.930 2.970 ;
        RECT 105.340 2.000 105.700 2.380 ;
        RECT 105.970 2.000 106.330 2.380 ;
        RECT 106.570 2.000 106.930 2.380 ;
      LAYER met3 ;
        RECT 2.315 376.110 4.320 377.385 ;
        RECT 105.130 376.310 107.130 377.585 ;
        RECT 2.315 373.250 4.315 375.545 ;
        RECT 2.315 364.450 4.315 366.745 ;
        RECT 2.315 362.745 4.320 364.020 ;
        RECT 105.140 362.325 107.140 363.600 ;
        RECT 2.315 356.110 4.320 357.385 ;
        RECT 105.130 356.310 107.130 357.585 ;
        RECT 2.315 353.250 4.315 355.545 ;
        RECT 2.315 344.450 4.315 346.745 ;
        RECT 2.315 342.745 4.320 344.020 ;
        RECT 105.140 342.325 107.140 343.600 ;
        RECT 2.315 336.100 4.320 337.375 ;
        RECT 105.130 336.310 107.130 337.585 ;
        RECT 2.315 333.250 4.315 335.545 ;
        RECT 2.315 324.455 4.315 326.750 ;
        RECT 2.315 322.400 4.320 323.675 ;
        RECT 105.140 322.325 107.140 323.600 ;
        RECT 2.315 316.510 4.320 317.785 ;
        RECT 105.130 316.310 107.130 317.585 ;
        RECT 2.320 315.340 4.320 315.545 ;
        RECT 2.315 313.250 4.320 315.340 ;
        RECT 2.315 304.455 4.315 306.750 ;
        RECT 2.315 302.270 4.330 303.545 ;
        RECT 105.140 302.325 107.140 303.600 ;
        RECT 2.315 296.255 4.320 297.530 ;
        RECT 105.135 296.580 107.135 297.855 ;
        RECT 2.320 295.340 4.320 295.545 ;
        RECT 2.315 293.250 4.320 295.340 ;
        RECT 2.315 284.445 4.315 286.740 ;
        RECT 2.315 282.370 4.320 283.645 ;
        RECT 105.140 282.000 107.140 283.275 ;
        RECT 2.315 276.335 4.330 277.610 ;
        RECT 105.135 276.085 107.135 277.360 ;
        RECT 2.315 273.250 4.315 275.545 ;
        RECT 2.315 264.455 4.315 266.750 ;
        RECT 2.315 262.505 4.320 263.780 ;
        RECT 105.140 261.725 107.140 263.000 ;
        RECT 2.315 256.570 4.320 257.845 ;
        RECT 105.140 256.050 107.140 257.325 ;
        RECT 2.315 253.250 4.315 255.545 ;
        RECT 2.315 244.455 4.315 246.750 ;
        RECT 2.315 242.460 4.320 243.735 ;
        RECT 105.140 242.255 107.140 243.530 ;
        RECT 2.315 236.695 4.320 237.970 ;
        RECT 105.140 236.490 107.140 237.765 ;
        RECT 2.315 233.250 4.315 235.545 ;
        RECT 2.315 224.455 4.315 226.750 ;
        RECT 2.315 224.450 4.180 224.455 ;
        RECT 2.315 221.395 4.315 222.670 ;
        RECT 105.140 220.910 107.140 222.185 ;
        RECT 2.315 195.215 4.025 195.695 ;
        RECT 2.315 189.775 4.025 190.255 ;
        RECT 2.315 184.335 4.025 184.815 ;
        RECT 42.635 181.410 47.035 182.660 ;
        RECT 58.235 181.410 67.035 182.660 ;
        RECT 78.235 181.410 87.035 182.660 ;
        RECT 98.235 181.410 102.635 182.660 ;
        RECT 42.635 178.260 102.635 181.410 ;
        RECT 105.140 179.715 107.140 180.990 ;
        RECT 43.885 167.060 61.385 178.260 ;
        RECT 63.885 167.060 81.385 178.260 ;
        RECT 83.885 167.060 101.385 178.260 ;
        RECT 105.140 175.915 107.140 178.210 ;
        RECT 105.140 175.910 107.005 175.915 ;
        RECT 105.140 167.115 107.140 169.410 ;
        RECT 105.140 167.110 107.005 167.115 ;
        RECT 42.635 163.910 102.635 167.060 ;
        RECT 105.135 164.440 107.135 165.715 ;
        RECT 42.635 162.660 47.035 163.910 ;
        RECT 58.235 162.660 67.035 163.910 ;
        RECT 78.235 162.660 87.035 163.910 ;
        RECT 98.235 162.660 102.635 163.910 ;
        RECT 2.315 160.360 4.330 161.800 ;
        RECT 105.125 160.360 107.140 161.800 ;
        RECT 4.730 158.750 9.130 160.000 ;
        RECT 20.330 158.750 29.130 160.000 ;
        RECT 40.330 158.750 49.130 160.000 ;
        RECT 60.330 158.750 69.130 160.000 ;
        RECT 80.330 158.750 89.130 160.000 ;
        RECT 100.330 158.750 104.730 160.000 ;
        RECT 2.315 156.450 4.315 157.725 ;
        RECT 4.730 155.600 104.730 158.750 ;
        RECT 105.140 156.450 107.140 157.725 ;
        RECT 2.315 153.255 4.315 155.555 ;
        RECT 2.315 144.450 4.315 146.745 ;
        RECT 5.980 144.400 23.480 155.600 ;
        RECT 25.980 144.400 43.480 155.600 ;
        RECT 45.980 144.400 63.480 155.600 ;
        RECT 65.980 144.400 83.480 155.600 ;
        RECT 85.980 144.400 103.480 155.600 ;
        RECT 2.315 141.890 4.315 143.165 ;
        RECT 4.730 141.250 104.730 144.400 ;
        RECT 105.140 141.645 107.140 142.920 ;
        RECT 4.730 138.750 9.130 141.250 ;
        RECT 20.330 138.750 29.130 141.250 ;
        RECT 40.330 138.750 49.130 141.250 ;
        RECT 60.330 138.750 69.130 141.250 ;
        RECT 80.330 138.750 89.130 141.250 ;
        RECT 100.330 138.750 104.730 141.250 ;
        RECT 2.315 136.870 4.315 138.145 ;
        RECT 4.730 135.600 104.730 138.750 ;
        RECT 105.135 136.060 107.135 137.335 ;
        RECT 2.315 133.250 4.315 135.545 ;
        RECT 2.315 124.450 4.315 126.745 ;
        RECT 5.980 124.400 23.480 135.600 ;
        RECT 25.980 124.400 43.480 135.600 ;
        RECT 45.980 124.400 63.480 135.600 ;
        RECT 65.980 124.400 83.480 135.600 ;
        RECT 85.980 124.400 103.480 135.600 ;
        RECT 2.315 121.980 4.320 123.255 ;
        RECT 4.730 121.250 104.730 124.400 ;
        RECT 105.140 121.845 107.140 123.120 ;
        RECT 4.730 118.750 9.130 121.250 ;
        RECT 20.330 118.750 29.130 121.250 ;
        RECT 40.330 118.750 49.130 121.250 ;
        RECT 60.330 118.750 69.130 121.250 ;
        RECT 80.330 118.750 89.130 121.250 ;
        RECT 100.330 118.750 104.730 121.250 ;
        RECT 2.315 116.570 4.320 117.845 ;
        RECT 4.730 115.600 104.730 118.750 ;
        RECT 105.140 115.970 107.140 117.245 ;
        RECT 2.315 113.250 4.315 115.545 ;
        RECT 2.315 104.455 4.315 106.750 ;
        RECT 5.980 104.400 23.480 115.600 ;
        RECT 25.980 104.400 43.480 115.600 ;
        RECT 45.980 104.400 63.480 115.600 ;
        RECT 65.980 104.400 83.480 115.600 ;
        RECT 85.980 104.400 103.480 115.600 ;
        RECT 2.315 102.195 4.320 103.470 ;
        RECT 4.730 101.250 104.730 104.400 ;
        RECT 105.135 101.765 107.135 103.040 ;
        RECT 4.730 98.750 9.130 101.250 ;
        RECT 20.330 98.750 29.130 101.250 ;
        RECT 40.330 98.750 49.130 101.250 ;
        RECT 60.330 98.750 69.130 101.250 ;
        RECT 80.330 98.750 89.130 101.250 ;
        RECT 100.330 98.750 104.730 101.250 ;
        RECT 2.315 96.690 4.320 97.965 ;
        RECT 4.730 95.600 104.730 98.750 ;
        RECT 105.135 95.910 107.135 97.185 ;
        RECT 2.315 93.250 4.315 95.545 ;
        RECT 2.315 84.450 4.315 86.745 ;
        RECT 5.980 84.400 23.480 95.600 ;
        RECT 25.980 84.400 43.480 95.600 ;
        RECT 45.980 84.400 63.480 95.600 ;
        RECT 65.980 84.400 83.480 95.600 ;
        RECT 85.980 84.400 103.480 95.600 ;
        RECT 2.315 82.360 4.325 83.635 ;
        RECT 4.730 81.250 104.730 84.400 ;
        RECT 105.135 82.105 107.135 83.380 ;
        RECT 4.730 78.750 9.130 81.250 ;
        RECT 20.330 78.750 29.130 81.250 ;
        RECT 40.330 78.750 49.130 81.250 ;
        RECT 60.330 78.750 69.130 81.250 ;
        RECT 80.330 78.750 89.130 81.250 ;
        RECT 100.330 78.750 104.730 81.250 ;
        RECT 2.315 76.280 4.330 77.555 ;
        RECT 4.730 75.600 104.730 78.750 ;
        RECT 105.135 76.035 107.135 77.310 ;
        RECT 2.315 73.250 4.315 75.545 ;
        RECT 2.315 64.450 4.315 66.745 ;
        RECT 5.980 64.400 23.480 75.600 ;
        RECT 25.980 64.400 43.480 75.600 ;
        RECT 45.980 64.400 63.480 75.600 ;
        RECT 65.980 64.400 83.480 75.600 ;
        RECT 85.980 64.400 103.480 75.600 ;
        RECT 2.315 61.955 4.320 63.230 ;
        RECT 4.730 61.250 104.730 64.400 ;
        RECT 105.140 61.820 107.140 63.095 ;
        RECT 4.730 58.750 9.130 61.250 ;
        RECT 20.330 58.750 29.130 61.250 ;
        RECT 40.330 58.750 49.130 61.250 ;
        RECT 60.330 58.750 69.130 61.250 ;
        RECT 80.330 58.750 89.130 61.250 ;
        RECT 100.330 58.750 104.730 61.250 ;
        RECT 2.315 56.345 4.320 57.620 ;
        RECT 4.730 55.600 104.730 58.750 ;
        RECT 105.135 56.035 107.135 57.310 ;
        RECT 2.315 53.255 4.315 55.550 ;
        RECT 2.315 44.445 4.315 46.740 ;
        RECT 5.980 44.400 23.480 55.600 ;
        RECT 25.980 44.400 43.480 55.600 ;
        RECT 45.980 44.400 63.480 55.600 ;
        RECT 65.980 44.400 83.480 55.600 ;
        RECT 85.980 44.400 103.480 55.600 ;
        RECT 2.315 42.045 4.315 43.320 ;
        RECT 4.730 41.250 104.730 44.400 ;
        RECT 105.140 41.820 107.140 43.095 ;
        RECT 4.730 38.750 9.130 41.250 ;
        RECT 20.330 38.750 29.130 41.250 ;
        RECT 40.330 38.750 49.130 41.250 ;
        RECT 60.330 38.750 69.130 41.250 ;
        RECT 80.330 38.750 89.130 41.250 ;
        RECT 100.330 38.750 104.730 41.250 ;
        RECT 2.315 36.490 4.315 37.765 ;
        RECT 4.730 35.600 104.730 38.750 ;
        RECT 105.135 36.035 107.135 37.310 ;
        RECT 2.315 33.255 4.315 35.550 ;
        RECT 2.315 24.450 4.315 26.745 ;
        RECT 5.980 24.400 23.480 35.600 ;
        RECT 25.980 24.400 43.480 35.600 ;
        RECT 45.980 24.400 63.480 35.600 ;
        RECT 65.980 24.400 83.480 35.600 ;
        RECT 85.980 24.400 103.480 35.600 ;
        RECT 2.315 22.375 4.325 23.650 ;
        RECT 4.730 21.250 104.730 24.400 ;
        RECT 105.140 21.820 107.140 23.095 ;
        RECT 4.730 18.750 9.130 21.250 ;
        RECT 20.330 18.750 29.130 21.250 ;
        RECT 40.330 18.750 49.130 21.250 ;
        RECT 60.330 18.750 69.130 21.250 ;
        RECT 80.330 18.750 89.130 21.250 ;
        RECT 100.330 18.750 104.730 21.250 ;
        RECT 2.315 16.490 4.315 17.765 ;
        RECT 4.730 15.600 104.730 18.750 ;
        RECT 105.135 16.035 107.135 17.310 ;
        RECT 2.315 13.255 4.315 15.550 ;
        RECT 2.315 4.450 4.315 6.745 ;
        RECT 5.980 4.400 23.480 15.600 ;
        RECT 25.980 4.400 43.480 15.600 ;
        RECT 45.980 4.400 63.480 15.600 ;
        RECT 65.980 4.400 83.480 15.600 ;
        RECT 85.980 4.400 103.480 15.600 ;
        RECT 2.315 2.375 4.325 3.650 ;
        RECT 4.730 1.250 104.730 4.400 ;
        RECT 105.140 1.820 107.140 3.095 ;
        RECT 4.730 0.000 9.130 1.250 ;
        RECT 20.330 0.000 29.130 1.250 ;
        RECT 40.330 0.000 49.130 1.250 ;
        RECT 60.330 0.000 69.130 1.250 ;
        RECT 80.330 0.000 89.130 1.250 ;
        RECT 100.330 0.000 104.730 1.250 ;
      LAYER via3 ;
        RECT 2.515 376.880 2.875 377.260 ;
        RECT 3.145 376.880 3.505 377.260 ;
        RECT 3.745 376.880 4.105 377.260 ;
        RECT 2.515 376.290 2.875 376.670 ;
        RECT 3.145 376.290 3.505 376.670 ;
        RECT 3.745 376.290 4.105 376.670 ;
        RECT 105.340 377.080 105.700 377.460 ;
        RECT 105.970 377.080 106.330 377.460 ;
        RECT 106.570 377.080 106.930 377.460 ;
        RECT 105.340 376.490 105.700 376.870 ;
        RECT 105.970 376.490 106.330 376.870 ;
        RECT 106.570 376.490 106.930 376.870 ;
        RECT 2.520 374.920 2.880 375.300 ;
        RECT 3.130 374.920 3.490 375.300 ;
        RECT 3.760 374.920 4.120 375.300 ;
        RECT 2.520 374.185 2.880 374.565 ;
        RECT 3.130 374.185 3.490 374.565 ;
        RECT 3.760 374.185 4.120 374.565 ;
        RECT 2.520 373.500 2.880 373.880 ;
        RECT 3.130 373.500 3.490 373.880 ;
        RECT 3.760 373.500 4.120 373.880 ;
        RECT 2.520 366.120 2.880 366.500 ;
        RECT 3.130 366.120 3.490 366.500 ;
        RECT 3.760 366.120 4.120 366.500 ;
        RECT 2.520 365.385 2.880 365.765 ;
        RECT 3.130 365.385 3.490 365.765 ;
        RECT 3.760 365.385 4.120 365.765 ;
        RECT 2.520 364.700 2.880 365.080 ;
        RECT 3.130 364.700 3.490 365.080 ;
        RECT 3.760 364.700 4.120 365.080 ;
        RECT 2.515 363.515 2.875 363.895 ;
        RECT 3.145 363.515 3.505 363.895 ;
        RECT 3.745 363.515 4.105 363.895 ;
        RECT 2.515 362.925 2.875 363.305 ;
        RECT 3.145 362.925 3.505 363.305 ;
        RECT 3.745 362.925 4.105 363.305 ;
        RECT 105.340 363.095 105.700 363.475 ;
        RECT 105.970 363.095 106.330 363.475 ;
        RECT 106.570 363.095 106.930 363.475 ;
        RECT 105.340 362.505 105.700 362.885 ;
        RECT 105.970 362.505 106.330 362.885 ;
        RECT 106.570 362.505 106.930 362.885 ;
        RECT 2.515 356.880 2.875 357.260 ;
        RECT 3.145 356.880 3.505 357.260 ;
        RECT 3.745 356.880 4.105 357.260 ;
        RECT 2.515 356.290 2.875 356.670 ;
        RECT 3.145 356.290 3.505 356.670 ;
        RECT 3.745 356.290 4.105 356.670 ;
        RECT 105.340 357.080 105.700 357.460 ;
        RECT 105.970 357.080 106.330 357.460 ;
        RECT 106.570 357.080 106.930 357.460 ;
        RECT 105.340 356.490 105.700 356.870 ;
        RECT 105.970 356.490 106.330 356.870 ;
        RECT 106.570 356.490 106.930 356.870 ;
        RECT 2.520 354.920 2.880 355.300 ;
        RECT 3.130 354.920 3.490 355.300 ;
        RECT 3.760 354.920 4.120 355.300 ;
        RECT 2.520 354.185 2.880 354.565 ;
        RECT 3.130 354.185 3.490 354.565 ;
        RECT 3.760 354.185 4.120 354.565 ;
        RECT 2.520 353.500 2.880 353.880 ;
        RECT 3.130 353.500 3.490 353.880 ;
        RECT 3.760 353.500 4.120 353.880 ;
        RECT 2.520 346.120 2.880 346.500 ;
        RECT 3.130 346.120 3.490 346.500 ;
        RECT 3.760 346.120 4.120 346.500 ;
        RECT 2.520 345.385 2.880 345.765 ;
        RECT 3.130 345.385 3.490 345.765 ;
        RECT 3.760 345.385 4.120 345.765 ;
        RECT 2.520 344.700 2.880 345.080 ;
        RECT 3.130 344.700 3.490 345.080 ;
        RECT 3.760 344.700 4.120 345.080 ;
        RECT 2.515 343.515 2.875 343.895 ;
        RECT 3.145 343.515 3.505 343.895 ;
        RECT 3.745 343.515 4.105 343.895 ;
        RECT 2.515 342.925 2.875 343.305 ;
        RECT 3.145 342.925 3.505 343.305 ;
        RECT 3.745 342.925 4.105 343.305 ;
        RECT 105.340 343.095 105.700 343.475 ;
        RECT 105.970 343.095 106.330 343.475 ;
        RECT 106.570 343.095 106.930 343.475 ;
        RECT 105.340 342.505 105.700 342.885 ;
        RECT 105.970 342.505 106.330 342.885 ;
        RECT 106.570 342.505 106.930 342.885 ;
        RECT 2.515 336.870 2.875 337.250 ;
        RECT 3.145 336.870 3.505 337.250 ;
        RECT 3.745 336.870 4.105 337.250 ;
        RECT 2.515 336.280 2.875 336.660 ;
        RECT 3.145 336.280 3.505 336.660 ;
        RECT 3.745 336.280 4.105 336.660 ;
        RECT 105.340 337.080 105.700 337.460 ;
        RECT 105.970 337.080 106.330 337.460 ;
        RECT 106.570 337.080 106.930 337.460 ;
        RECT 105.340 336.490 105.700 336.870 ;
        RECT 105.970 336.490 106.330 336.870 ;
        RECT 106.570 336.490 106.930 336.870 ;
        RECT 2.520 334.920 2.880 335.300 ;
        RECT 3.130 334.920 3.490 335.300 ;
        RECT 3.760 334.920 4.120 335.300 ;
        RECT 2.520 334.185 2.880 334.565 ;
        RECT 3.130 334.185 3.490 334.565 ;
        RECT 3.760 334.185 4.120 334.565 ;
        RECT 2.520 333.500 2.880 333.880 ;
        RECT 3.130 333.500 3.490 333.880 ;
        RECT 3.760 333.500 4.120 333.880 ;
        RECT 2.520 326.125 2.880 326.505 ;
        RECT 3.130 326.125 3.490 326.505 ;
        RECT 3.760 326.125 4.120 326.505 ;
        RECT 2.520 325.390 2.880 325.770 ;
        RECT 3.130 325.390 3.490 325.770 ;
        RECT 3.760 325.390 4.120 325.770 ;
        RECT 2.520 324.705 2.880 325.085 ;
        RECT 3.130 324.705 3.490 325.085 ;
        RECT 3.760 324.705 4.120 325.085 ;
        RECT 2.515 323.170 2.875 323.550 ;
        RECT 3.145 323.170 3.505 323.550 ;
        RECT 3.745 323.170 4.105 323.550 ;
        RECT 2.515 322.580 2.875 322.960 ;
        RECT 3.145 322.580 3.505 322.960 ;
        RECT 3.745 322.580 4.105 322.960 ;
        RECT 105.340 323.095 105.700 323.475 ;
        RECT 105.970 323.095 106.330 323.475 ;
        RECT 106.570 323.095 106.930 323.475 ;
        RECT 105.340 322.505 105.700 322.885 ;
        RECT 105.970 322.505 106.330 322.885 ;
        RECT 106.570 322.505 106.930 322.885 ;
        RECT 2.515 317.280 2.875 317.660 ;
        RECT 3.145 317.280 3.505 317.660 ;
        RECT 3.745 317.280 4.105 317.660 ;
        RECT 2.515 316.690 2.875 317.070 ;
        RECT 3.145 316.690 3.505 317.070 ;
        RECT 3.745 316.690 4.105 317.070 ;
        RECT 105.340 317.080 105.700 317.460 ;
        RECT 105.970 317.080 106.330 317.460 ;
        RECT 106.570 317.080 106.930 317.460 ;
        RECT 105.340 316.490 105.700 316.870 ;
        RECT 105.970 316.490 106.330 316.870 ;
        RECT 106.570 316.490 106.930 316.870 ;
        RECT 2.520 314.920 2.880 315.300 ;
        RECT 3.130 314.920 3.490 315.300 ;
        RECT 3.760 314.920 4.120 315.300 ;
        RECT 2.520 314.185 2.880 314.565 ;
        RECT 3.130 314.185 3.490 314.565 ;
        RECT 3.760 314.185 4.120 314.565 ;
        RECT 2.520 313.500 2.880 313.880 ;
        RECT 3.130 313.500 3.490 313.880 ;
        RECT 3.760 313.500 4.120 313.880 ;
        RECT 2.520 306.125 2.880 306.505 ;
        RECT 3.130 306.125 3.490 306.505 ;
        RECT 3.760 306.125 4.120 306.505 ;
        RECT 2.520 305.390 2.880 305.770 ;
        RECT 3.130 305.390 3.490 305.770 ;
        RECT 3.760 305.390 4.120 305.770 ;
        RECT 2.520 304.705 2.880 305.085 ;
        RECT 3.130 304.705 3.490 305.085 ;
        RECT 3.760 304.705 4.120 305.085 ;
        RECT 2.515 303.040 2.875 303.420 ;
        RECT 3.145 303.040 3.505 303.420 ;
        RECT 3.745 303.040 4.105 303.420 ;
        RECT 2.515 302.450 2.875 302.830 ;
        RECT 3.145 302.450 3.505 302.830 ;
        RECT 3.745 302.450 4.105 302.830 ;
        RECT 105.340 303.095 105.700 303.475 ;
        RECT 105.970 303.095 106.330 303.475 ;
        RECT 106.570 303.095 106.930 303.475 ;
        RECT 105.340 302.505 105.700 302.885 ;
        RECT 105.970 302.505 106.330 302.885 ;
        RECT 106.570 302.505 106.930 302.885 ;
        RECT 2.515 297.025 2.875 297.405 ;
        RECT 3.145 297.025 3.505 297.405 ;
        RECT 3.745 297.025 4.105 297.405 ;
        RECT 2.515 296.435 2.875 296.815 ;
        RECT 3.145 296.435 3.505 296.815 ;
        RECT 3.745 296.435 4.105 296.815 ;
        RECT 105.340 297.350 105.700 297.730 ;
        RECT 105.970 297.350 106.330 297.730 ;
        RECT 106.570 297.350 106.930 297.730 ;
        RECT 105.340 296.760 105.700 297.140 ;
        RECT 105.970 296.760 106.330 297.140 ;
        RECT 106.570 296.760 106.930 297.140 ;
        RECT 2.520 294.920 2.880 295.300 ;
        RECT 3.130 294.920 3.490 295.300 ;
        RECT 3.760 294.920 4.120 295.300 ;
        RECT 2.520 294.185 2.880 294.565 ;
        RECT 3.130 294.185 3.490 294.565 ;
        RECT 3.760 294.185 4.120 294.565 ;
        RECT 2.520 293.500 2.880 293.880 ;
        RECT 3.130 293.500 3.490 293.880 ;
        RECT 3.760 293.500 4.120 293.880 ;
        RECT 2.520 286.115 2.880 286.495 ;
        RECT 3.130 286.115 3.490 286.495 ;
        RECT 3.760 286.115 4.120 286.495 ;
        RECT 2.520 285.380 2.880 285.760 ;
        RECT 3.130 285.380 3.490 285.760 ;
        RECT 3.760 285.380 4.120 285.760 ;
        RECT 2.520 284.695 2.880 285.075 ;
        RECT 3.130 284.695 3.490 285.075 ;
        RECT 3.760 284.695 4.120 285.075 ;
        RECT 2.515 283.140 2.875 283.520 ;
        RECT 3.145 283.140 3.505 283.520 ;
        RECT 3.745 283.140 4.105 283.520 ;
        RECT 2.515 282.550 2.875 282.930 ;
        RECT 3.145 282.550 3.505 282.930 ;
        RECT 3.745 282.550 4.105 282.930 ;
        RECT 105.340 282.770 105.700 283.150 ;
        RECT 105.970 282.770 106.330 283.150 ;
        RECT 106.570 282.770 106.930 283.150 ;
        RECT 105.340 282.180 105.700 282.560 ;
        RECT 105.970 282.180 106.330 282.560 ;
        RECT 106.570 282.180 106.930 282.560 ;
        RECT 2.515 277.105 2.875 277.485 ;
        RECT 3.145 277.105 3.505 277.485 ;
        RECT 3.745 277.105 4.105 277.485 ;
        RECT 2.515 276.515 2.875 276.895 ;
        RECT 3.145 276.515 3.505 276.895 ;
        RECT 3.745 276.515 4.105 276.895 ;
        RECT 105.340 276.855 105.700 277.235 ;
        RECT 105.970 276.855 106.330 277.235 ;
        RECT 106.570 276.855 106.930 277.235 ;
        RECT 105.340 276.265 105.700 276.645 ;
        RECT 105.970 276.265 106.330 276.645 ;
        RECT 106.570 276.265 106.930 276.645 ;
        RECT 2.520 274.920 2.880 275.300 ;
        RECT 3.130 274.920 3.490 275.300 ;
        RECT 3.760 274.920 4.120 275.300 ;
        RECT 2.520 274.185 2.880 274.565 ;
        RECT 3.130 274.185 3.490 274.565 ;
        RECT 3.760 274.185 4.120 274.565 ;
        RECT 2.520 273.500 2.880 273.880 ;
        RECT 3.130 273.500 3.490 273.880 ;
        RECT 3.760 273.500 4.120 273.880 ;
        RECT 2.520 266.125 2.880 266.505 ;
        RECT 3.130 266.125 3.490 266.505 ;
        RECT 3.760 266.125 4.120 266.505 ;
        RECT 2.520 265.390 2.880 265.770 ;
        RECT 3.130 265.390 3.490 265.770 ;
        RECT 3.760 265.390 4.120 265.770 ;
        RECT 2.520 264.705 2.880 265.085 ;
        RECT 3.130 264.705 3.490 265.085 ;
        RECT 3.760 264.705 4.120 265.085 ;
        RECT 2.515 263.275 2.875 263.655 ;
        RECT 3.145 263.275 3.505 263.655 ;
        RECT 3.745 263.275 4.105 263.655 ;
        RECT 2.515 262.685 2.875 263.065 ;
        RECT 3.145 262.685 3.505 263.065 ;
        RECT 3.745 262.685 4.105 263.065 ;
        RECT 105.340 262.495 105.700 262.875 ;
        RECT 105.970 262.495 106.330 262.875 ;
        RECT 106.570 262.495 106.930 262.875 ;
        RECT 105.340 261.905 105.700 262.285 ;
        RECT 105.970 261.905 106.330 262.285 ;
        RECT 106.570 261.905 106.930 262.285 ;
        RECT 2.515 257.340 2.875 257.720 ;
        RECT 3.145 257.340 3.505 257.720 ;
        RECT 3.745 257.340 4.105 257.720 ;
        RECT 2.515 256.750 2.875 257.130 ;
        RECT 3.145 256.750 3.505 257.130 ;
        RECT 3.745 256.750 4.105 257.130 ;
        RECT 105.340 256.820 105.700 257.200 ;
        RECT 105.970 256.820 106.330 257.200 ;
        RECT 106.570 256.820 106.930 257.200 ;
        RECT 105.340 256.230 105.700 256.610 ;
        RECT 105.970 256.230 106.330 256.610 ;
        RECT 106.570 256.230 106.930 256.610 ;
        RECT 2.520 254.920 2.880 255.300 ;
        RECT 3.130 254.920 3.490 255.300 ;
        RECT 3.760 254.920 4.120 255.300 ;
        RECT 2.520 254.185 2.880 254.565 ;
        RECT 3.130 254.185 3.490 254.565 ;
        RECT 3.760 254.185 4.120 254.565 ;
        RECT 2.520 253.500 2.880 253.880 ;
        RECT 3.130 253.500 3.490 253.880 ;
        RECT 3.760 253.500 4.120 253.880 ;
        RECT 2.520 246.125 2.880 246.505 ;
        RECT 3.130 246.125 3.490 246.505 ;
        RECT 3.760 246.125 4.120 246.505 ;
        RECT 2.520 245.390 2.880 245.770 ;
        RECT 3.130 245.390 3.490 245.770 ;
        RECT 3.760 245.390 4.120 245.770 ;
        RECT 2.520 244.705 2.880 245.085 ;
        RECT 3.130 244.705 3.490 245.085 ;
        RECT 3.760 244.705 4.120 245.085 ;
        RECT 2.515 243.230 2.875 243.610 ;
        RECT 3.145 243.230 3.505 243.610 ;
        RECT 3.745 243.230 4.105 243.610 ;
        RECT 2.515 242.640 2.875 243.020 ;
        RECT 3.145 242.640 3.505 243.020 ;
        RECT 3.745 242.640 4.105 243.020 ;
        RECT 105.340 243.025 105.700 243.405 ;
        RECT 105.970 243.025 106.330 243.405 ;
        RECT 106.570 243.025 106.930 243.405 ;
        RECT 105.340 242.435 105.700 242.815 ;
        RECT 105.970 242.435 106.330 242.815 ;
        RECT 106.570 242.435 106.930 242.815 ;
        RECT 2.515 237.465 2.875 237.845 ;
        RECT 3.145 237.465 3.505 237.845 ;
        RECT 3.745 237.465 4.105 237.845 ;
        RECT 2.515 236.875 2.875 237.255 ;
        RECT 3.145 236.875 3.505 237.255 ;
        RECT 3.745 236.875 4.105 237.255 ;
        RECT 105.340 237.260 105.700 237.640 ;
        RECT 105.970 237.260 106.330 237.640 ;
        RECT 106.570 237.260 106.930 237.640 ;
        RECT 105.340 236.670 105.700 237.050 ;
        RECT 105.970 236.670 106.330 237.050 ;
        RECT 106.570 236.670 106.930 237.050 ;
        RECT 2.520 234.920 2.880 235.300 ;
        RECT 3.130 234.920 3.490 235.300 ;
        RECT 3.760 234.920 4.120 235.300 ;
        RECT 2.520 234.185 2.880 234.565 ;
        RECT 3.130 234.185 3.490 234.565 ;
        RECT 3.760 234.185 4.120 234.565 ;
        RECT 2.520 233.500 2.880 233.880 ;
        RECT 3.130 233.500 3.490 233.880 ;
        RECT 3.760 233.500 4.120 233.880 ;
        RECT 2.520 226.120 2.880 226.500 ;
        RECT 3.130 226.120 3.490 226.500 ;
        RECT 3.760 226.120 4.120 226.500 ;
        RECT 2.520 225.385 2.880 225.765 ;
        RECT 3.130 225.385 3.490 225.765 ;
        RECT 3.760 225.385 4.120 225.765 ;
        RECT 2.520 224.700 2.880 225.080 ;
        RECT 3.130 224.700 3.490 225.080 ;
        RECT 3.760 224.700 4.120 225.080 ;
        RECT 2.515 222.165 2.875 222.545 ;
        RECT 3.145 222.165 3.505 222.545 ;
        RECT 3.745 222.165 4.105 222.545 ;
        RECT 2.515 221.575 2.875 221.955 ;
        RECT 3.145 221.575 3.505 221.955 ;
        RECT 3.745 221.575 4.105 221.955 ;
        RECT 105.340 221.680 105.700 222.060 ;
        RECT 105.970 221.680 106.330 222.060 ;
        RECT 106.570 221.680 106.930 222.060 ;
        RECT 105.340 221.090 105.700 221.470 ;
        RECT 105.970 221.090 106.330 221.470 ;
        RECT 106.570 221.090 106.930 221.470 ;
        RECT 2.390 195.255 2.810 195.655 ;
        RECT 2.960 195.255 3.380 195.655 ;
        RECT 3.530 195.255 3.950 195.655 ;
        RECT 2.390 189.815 2.810 190.215 ;
        RECT 2.960 189.815 3.380 190.215 ;
        RECT 3.530 189.815 3.950 190.215 ;
        RECT 2.390 184.375 2.810 184.775 ;
        RECT 2.960 184.375 3.380 184.775 ;
        RECT 3.530 184.375 3.950 184.775 ;
        RECT 42.735 181.710 43.585 182.560 ;
        RECT 43.685 181.710 44.535 182.560 ;
        RECT 45.135 181.710 45.985 182.560 ;
        RECT 46.085 181.710 46.935 182.560 ;
        RECT 42.735 180.760 43.585 181.610 ;
        RECT 58.335 181.710 59.185 182.560 ;
        RECT 59.285 181.710 60.135 182.560 ;
        RECT 60.735 181.710 61.585 182.560 ;
        RECT 61.685 181.710 62.535 182.560 ;
        RECT 62.735 181.710 63.585 182.560 ;
        RECT 63.685 181.710 64.535 182.560 ;
        RECT 65.135 181.710 65.985 182.560 ;
        RECT 66.085 181.710 66.935 182.560 ;
        RECT 61.685 180.760 62.535 181.610 ;
        RECT 62.735 180.760 63.585 181.610 ;
        RECT 78.335 181.710 79.185 182.560 ;
        RECT 79.285 181.710 80.135 182.560 ;
        RECT 80.735 181.710 81.585 182.560 ;
        RECT 81.685 181.710 82.535 182.560 ;
        RECT 82.735 181.710 83.585 182.560 ;
        RECT 83.685 181.710 84.535 182.560 ;
        RECT 85.135 181.710 85.985 182.560 ;
        RECT 86.085 181.710 86.935 182.560 ;
        RECT 81.685 180.760 82.535 181.610 ;
        RECT 82.735 180.760 83.585 181.610 ;
        RECT 98.335 181.710 99.185 182.560 ;
        RECT 99.285 181.710 100.135 182.560 ;
        RECT 100.735 181.710 101.585 182.560 ;
        RECT 101.685 181.710 102.535 182.560 ;
        RECT 101.685 180.760 102.535 181.610 ;
        RECT 42.735 179.310 43.585 180.160 ;
        RECT 61.685 179.310 62.535 180.160 ;
        RECT 62.735 179.310 63.585 180.160 ;
        RECT 81.685 179.310 82.535 180.160 ;
        RECT 82.735 179.310 83.585 180.160 ;
        RECT 101.685 179.310 102.535 180.160 ;
        RECT 105.305 180.460 105.705 180.860 ;
        RECT 105.930 180.460 106.330 180.860 ;
        RECT 106.555 180.460 106.955 180.860 ;
        RECT 105.300 179.860 105.700 180.260 ;
        RECT 105.925 179.860 106.325 180.260 ;
        RECT 106.550 179.860 106.950 180.260 ;
        RECT 42.735 178.360 43.585 179.210 ;
        RECT 61.685 178.360 62.535 179.210 ;
        RECT 62.735 178.360 63.585 179.210 ;
        RECT 81.685 178.360 82.535 179.210 ;
        RECT 82.735 178.360 83.585 179.210 ;
        RECT 101.685 178.360 102.535 179.210 ;
        RECT 105.345 177.580 105.705 177.960 ;
        RECT 105.955 177.580 106.315 177.960 ;
        RECT 106.585 177.580 106.945 177.960 ;
        RECT 105.345 176.845 105.705 177.225 ;
        RECT 105.955 176.845 106.315 177.225 ;
        RECT 106.585 176.845 106.945 177.225 ;
        RECT 105.345 176.160 105.705 176.540 ;
        RECT 105.955 176.160 106.315 176.540 ;
        RECT 106.585 176.160 106.945 176.540 ;
        RECT 105.345 168.780 105.705 169.160 ;
        RECT 105.955 168.780 106.315 169.160 ;
        RECT 106.585 168.780 106.945 169.160 ;
        RECT 105.345 168.045 105.705 168.425 ;
        RECT 105.955 168.045 106.315 168.425 ;
        RECT 106.585 168.045 106.945 168.425 ;
        RECT 105.345 167.360 105.705 167.740 ;
        RECT 105.955 167.360 106.315 167.740 ;
        RECT 106.585 167.360 106.945 167.740 ;
        RECT 42.735 166.110 43.585 166.960 ;
        RECT 61.685 166.110 62.535 166.960 ;
        RECT 62.735 166.110 63.585 166.960 ;
        RECT 81.685 166.110 82.535 166.960 ;
        RECT 82.735 166.110 83.585 166.960 ;
        RECT 101.685 166.110 102.535 166.960 ;
        RECT 42.735 165.160 43.585 166.010 ;
        RECT 61.685 165.160 62.535 166.010 ;
        RECT 62.735 165.160 63.585 166.010 ;
        RECT 81.685 165.160 82.535 166.010 ;
        RECT 82.735 165.160 83.585 166.010 ;
        RECT 101.685 165.160 102.535 166.010 ;
        RECT 42.735 163.710 43.585 164.560 ;
        RECT 42.735 162.760 43.585 163.610 ;
        RECT 43.685 162.760 44.535 163.610 ;
        RECT 45.135 162.760 45.985 163.610 ;
        RECT 46.085 162.760 46.935 163.610 ;
        RECT 61.685 163.710 62.535 164.560 ;
        RECT 62.735 163.710 63.585 164.560 ;
        RECT 58.335 162.760 59.185 163.610 ;
        RECT 59.285 162.760 60.135 163.610 ;
        RECT 60.735 162.760 61.585 163.610 ;
        RECT 61.685 162.760 62.535 163.610 ;
        RECT 62.735 162.760 63.585 163.610 ;
        RECT 63.685 162.760 64.535 163.610 ;
        RECT 65.135 162.760 65.985 163.610 ;
        RECT 66.085 162.760 66.935 163.610 ;
        RECT 81.685 163.710 82.535 164.560 ;
        RECT 82.735 163.710 83.585 164.560 ;
        RECT 78.335 162.760 79.185 163.610 ;
        RECT 79.285 162.760 80.135 163.610 ;
        RECT 80.735 162.760 81.585 163.610 ;
        RECT 81.685 162.760 82.535 163.610 ;
        RECT 82.735 162.760 83.585 163.610 ;
        RECT 83.685 162.760 84.535 163.610 ;
        RECT 85.135 162.760 85.985 163.610 ;
        RECT 86.085 162.760 86.935 163.610 ;
        RECT 101.685 163.710 102.535 164.560 ;
        RECT 105.300 165.185 105.700 165.585 ;
        RECT 105.925 165.185 106.325 165.585 ;
        RECT 106.550 165.185 106.950 165.585 ;
        RECT 105.295 164.585 105.695 164.985 ;
        RECT 105.920 164.585 106.320 164.985 ;
        RECT 106.545 164.585 106.945 164.985 ;
        RECT 98.335 162.760 99.185 163.610 ;
        RECT 99.285 162.760 100.135 163.610 ;
        RECT 100.735 162.760 101.585 163.610 ;
        RECT 101.685 162.760 102.535 163.610 ;
        RECT 2.515 161.130 2.875 161.510 ;
        RECT 3.145 161.130 3.505 161.510 ;
        RECT 3.745 161.130 4.105 161.510 ;
        RECT 2.515 160.540 2.875 160.920 ;
        RECT 3.145 160.540 3.505 160.920 ;
        RECT 3.745 160.540 4.105 160.920 ;
        RECT 105.340 161.130 105.700 161.510 ;
        RECT 105.970 161.130 106.330 161.510 ;
        RECT 106.570 161.130 106.930 161.510 ;
        RECT 105.340 160.540 105.700 160.920 ;
        RECT 105.970 160.540 106.330 160.920 ;
        RECT 106.570 160.540 106.930 160.920 ;
        RECT 4.830 159.050 5.680 159.900 ;
        RECT 5.780 159.050 6.630 159.900 ;
        RECT 7.230 159.050 8.080 159.900 ;
        RECT 8.180 159.050 9.030 159.900 ;
        RECT 4.830 158.100 5.680 158.950 ;
        RECT 20.430 159.050 21.280 159.900 ;
        RECT 21.380 159.050 22.230 159.900 ;
        RECT 22.830 159.050 23.680 159.900 ;
        RECT 23.780 159.050 24.630 159.900 ;
        RECT 24.830 159.050 25.680 159.900 ;
        RECT 25.780 159.050 26.630 159.900 ;
        RECT 27.230 159.050 28.080 159.900 ;
        RECT 28.180 159.050 29.030 159.900 ;
        RECT 23.780 158.100 24.630 158.950 ;
        RECT 24.830 158.100 25.680 158.950 ;
        RECT 40.430 159.050 41.280 159.900 ;
        RECT 41.380 159.050 42.230 159.900 ;
        RECT 42.830 159.050 43.680 159.900 ;
        RECT 43.780 159.050 44.630 159.900 ;
        RECT 44.830 159.050 45.680 159.900 ;
        RECT 45.780 159.050 46.630 159.900 ;
        RECT 47.230 159.050 48.080 159.900 ;
        RECT 48.180 159.050 49.030 159.900 ;
        RECT 43.780 158.100 44.630 158.950 ;
        RECT 44.830 158.100 45.680 158.950 ;
        RECT 60.430 159.050 61.280 159.900 ;
        RECT 61.380 159.050 62.230 159.900 ;
        RECT 62.830 159.050 63.680 159.900 ;
        RECT 63.780 159.050 64.630 159.900 ;
        RECT 64.830 159.050 65.680 159.900 ;
        RECT 65.780 159.050 66.630 159.900 ;
        RECT 67.230 159.050 68.080 159.900 ;
        RECT 68.180 159.050 69.030 159.900 ;
        RECT 63.780 158.100 64.630 158.950 ;
        RECT 64.830 158.100 65.680 158.950 ;
        RECT 80.430 159.050 81.280 159.900 ;
        RECT 81.380 159.050 82.230 159.900 ;
        RECT 82.830 159.050 83.680 159.900 ;
        RECT 83.780 159.050 84.630 159.900 ;
        RECT 84.830 159.050 85.680 159.900 ;
        RECT 85.780 159.050 86.630 159.900 ;
        RECT 87.230 159.050 88.080 159.900 ;
        RECT 88.180 159.050 89.030 159.900 ;
        RECT 83.780 158.100 84.630 158.950 ;
        RECT 84.830 158.100 85.680 158.950 ;
        RECT 100.430 159.050 101.280 159.900 ;
        RECT 101.380 159.050 102.230 159.900 ;
        RECT 102.830 159.050 103.680 159.900 ;
        RECT 103.780 159.050 104.630 159.900 ;
        RECT 103.780 158.100 104.630 158.950 ;
        RECT 2.515 157.220 2.875 157.600 ;
        RECT 3.145 157.220 3.505 157.600 ;
        RECT 3.745 157.220 4.105 157.600 ;
        RECT 2.515 156.630 2.875 157.010 ;
        RECT 3.145 156.630 3.505 157.010 ;
        RECT 3.745 156.630 4.105 157.010 ;
        RECT 4.830 156.650 5.680 157.500 ;
        RECT 23.780 156.650 24.630 157.500 ;
        RECT 24.830 156.650 25.680 157.500 ;
        RECT 43.780 156.650 44.630 157.500 ;
        RECT 44.830 156.650 45.680 157.500 ;
        RECT 63.780 156.650 64.630 157.500 ;
        RECT 64.830 156.650 65.680 157.500 ;
        RECT 83.780 156.650 84.630 157.500 ;
        RECT 84.830 156.650 85.680 157.500 ;
        RECT 103.780 156.650 104.630 157.500 ;
        RECT 4.830 155.700 5.680 156.550 ;
        RECT 23.780 155.700 24.630 156.550 ;
        RECT 24.830 155.700 25.680 156.550 ;
        RECT 43.780 155.700 44.630 156.550 ;
        RECT 44.830 155.700 45.680 156.550 ;
        RECT 63.780 155.700 64.630 156.550 ;
        RECT 64.830 155.700 65.680 156.550 ;
        RECT 83.780 155.700 84.630 156.550 ;
        RECT 84.830 155.700 85.680 156.550 ;
        RECT 103.780 155.700 104.630 156.550 ;
        RECT 105.340 157.220 105.700 157.600 ;
        RECT 105.970 157.220 106.330 157.600 ;
        RECT 106.570 157.220 106.930 157.600 ;
        RECT 105.340 156.630 105.700 157.010 ;
        RECT 105.970 156.630 106.330 157.010 ;
        RECT 106.570 156.630 106.930 157.010 ;
        RECT 2.520 154.925 2.880 155.305 ;
        RECT 3.130 154.925 3.490 155.305 ;
        RECT 3.760 154.925 4.120 155.305 ;
        RECT 2.520 154.190 2.880 154.570 ;
        RECT 3.130 154.190 3.490 154.570 ;
        RECT 3.760 154.190 4.120 154.570 ;
        RECT 2.520 153.505 2.880 153.885 ;
        RECT 3.130 153.505 3.490 153.885 ;
        RECT 3.760 153.505 4.120 153.885 ;
        RECT 2.520 146.090 2.880 146.470 ;
        RECT 3.130 146.090 3.490 146.470 ;
        RECT 3.760 146.090 4.120 146.470 ;
        RECT 2.520 145.355 2.880 145.735 ;
        RECT 3.130 145.355 3.490 145.735 ;
        RECT 3.760 145.355 4.120 145.735 ;
        RECT 2.520 144.670 2.880 145.050 ;
        RECT 3.130 144.670 3.490 145.050 ;
        RECT 3.760 144.670 4.120 145.050 ;
        RECT 4.830 143.450 5.680 144.300 ;
        RECT 23.780 143.450 24.630 144.300 ;
        RECT 24.830 143.450 25.680 144.300 ;
        RECT 43.780 143.450 44.630 144.300 ;
        RECT 44.830 143.450 45.680 144.300 ;
        RECT 63.780 143.450 64.630 144.300 ;
        RECT 64.830 143.450 65.680 144.300 ;
        RECT 83.780 143.450 84.630 144.300 ;
        RECT 84.830 143.450 85.680 144.300 ;
        RECT 103.780 143.450 104.630 144.300 ;
        RECT 2.515 142.660 2.875 143.040 ;
        RECT 3.145 142.660 3.505 143.040 ;
        RECT 3.745 142.660 4.105 143.040 ;
        RECT 2.515 142.070 2.875 142.450 ;
        RECT 3.145 142.070 3.505 142.450 ;
        RECT 3.745 142.070 4.105 142.450 ;
        RECT 4.830 142.500 5.680 143.350 ;
        RECT 23.780 142.500 24.630 143.350 ;
        RECT 24.830 142.500 25.680 143.350 ;
        RECT 43.780 142.500 44.630 143.350 ;
        RECT 44.830 142.500 45.680 143.350 ;
        RECT 63.780 142.500 64.630 143.350 ;
        RECT 64.830 142.500 65.680 143.350 ;
        RECT 83.780 142.500 84.630 143.350 ;
        RECT 84.830 142.500 85.680 143.350 ;
        RECT 103.780 142.500 104.630 143.350 ;
        RECT 4.830 141.050 5.680 141.900 ;
        RECT 4.830 140.100 5.680 140.950 ;
        RECT 5.780 140.100 6.630 140.950 ;
        RECT 7.230 140.100 8.080 140.950 ;
        RECT 8.180 140.100 9.030 140.950 ;
        RECT 4.830 139.050 5.680 139.900 ;
        RECT 5.780 139.050 6.630 139.900 ;
        RECT 7.230 139.050 8.080 139.900 ;
        RECT 8.180 139.050 9.030 139.900 ;
        RECT 2.515 137.640 2.875 138.020 ;
        RECT 3.145 137.640 3.505 138.020 ;
        RECT 3.745 137.640 4.105 138.020 ;
        RECT 2.515 137.050 2.875 137.430 ;
        RECT 3.145 137.050 3.505 137.430 ;
        RECT 3.745 137.050 4.105 137.430 ;
        RECT 4.830 138.100 5.680 138.950 ;
        RECT 23.780 141.050 24.630 141.900 ;
        RECT 24.830 141.050 25.680 141.900 ;
        RECT 20.430 140.100 21.280 140.950 ;
        RECT 21.380 140.100 22.230 140.950 ;
        RECT 22.830 140.100 23.680 140.950 ;
        RECT 23.780 140.100 24.630 140.950 ;
        RECT 24.830 140.100 25.680 140.950 ;
        RECT 25.780 140.100 26.630 140.950 ;
        RECT 27.230 140.100 28.080 140.950 ;
        RECT 28.180 140.100 29.030 140.950 ;
        RECT 20.430 139.050 21.280 139.900 ;
        RECT 21.380 139.050 22.230 139.900 ;
        RECT 22.830 139.050 23.680 139.900 ;
        RECT 23.780 139.050 24.630 139.900 ;
        RECT 24.830 139.050 25.680 139.900 ;
        RECT 25.780 139.050 26.630 139.900 ;
        RECT 27.230 139.050 28.080 139.900 ;
        RECT 28.180 139.050 29.030 139.900 ;
        RECT 23.780 138.100 24.630 138.950 ;
        RECT 24.830 138.100 25.680 138.950 ;
        RECT 43.780 141.050 44.630 141.900 ;
        RECT 44.830 141.050 45.680 141.900 ;
        RECT 40.430 140.100 41.280 140.950 ;
        RECT 41.380 140.100 42.230 140.950 ;
        RECT 42.830 140.100 43.680 140.950 ;
        RECT 43.780 140.100 44.630 140.950 ;
        RECT 44.830 140.100 45.680 140.950 ;
        RECT 45.780 140.100 46.630 140.950 ;
        RECT 47.230 140.100 48.080 140.950 ;
        RECT 48.180 140.100 49.030 140.950 ;
        RECT 40.430 139.050 41.280 139.900 ;
        RECT 41.380 139.050 42.230 139.900 ;
        RECT 42.830 139.050 43.680 139.900 ;
        RECT 43.780 139.050 44.630 139.900 ;
        RECT 44.830 139.050 45.680 139.900 ;
        RECT 45.780 139.050 46.630 139.900 ;
        RECT 47.230 139.050 48.080 139.900 ;
        RECT 48.180 139.050 49.030 139.900 ;
        RECT 43.780 138.100 44.630 138.950 ;
        RECT 44.830 138.100 45.680 138.950 ;
        RECT 63.780 141.050 64.630 141.900 ;
        RECT 64.830 141.050 65.680 141.900 ;
        RECT 60.430 140.100 61.280 140.950 ;
        RECT 61.380 140.100 62.230 140.950 ;
        RECT 62.830 140.100 63.680 140.950 ;
        RECT 63.780 140.100 64.630 140.950 ;
        RECT 64.830 140.100 65.680 140.950 ;
        RECT 65.780 140.100 66.630 140.950 ;
        RECT 67.230 140.100 68.080 140.950 ;
        RECT 68.180 140.100 69.030 140.950 ;
        RECT 60.430 139.050 61.280 139.900 ;
        RECT 61.380 139.050 62.230 139.900 ;
        RECT 62.830 139.050 63.680 139.900 ;
        RECT 63.780 139.050 64.630 139.900 ;
        RECT 64.830 139.050 65.680 139.900 ;
        RECT 65.780 139.050 66.630 139.900 ;
        RECT 67.230 139.050 68.080 139.900 ;
        RECT 68.180 139.050 69.030 139.900 ;
        RECT 63.780 138.100 64.630 138.950 ;
        RECT 64.830 138.100 65.680 138.950 ;
        RECT 83.780 141.050 84.630 141.900 ;
        RECT 84.830 141.050 85.680 141.900 ;
        RECT 80.430 140.100 81.280 140.950 ;
        RECT 81.380 140.100 82.230 140.950 ;
        RECT 82.830 140.100 83.680 140.950 ;
        RECT 83.780 140.100 84.630 140.950 ;
        RECT 84.830 140.100 85.680 140.950 ;
        RECT 85.780 140.100 86.630 140.950 ;
        RECT 87.230 140.100 88.080 140.950 ;
        RECT 88.180 140.100 89.030 140.950 ;
        RECT 80.430 139.050 81.280 139.900 ;
        RECT 81.380 139.050 82.230 139.900 ;
        RECT 82.830 139.050 83.680 139.900 ;
        RECT 83.780 139.050 84.630 139.900 ;
        RECT 84.830 139.050 85.680 139.900 ;
        RECT 85.780 139.050 86.630 139.900 ;
        RECT 87.230 139.050 88.080 139.900 ;
        RECT 88.180 139.050 89.030 139.900 ;
        RECT 83.780 138.100 84.630 138.950 ;
        RECT 84.830 138.100 85.680 138.950 ;
        RECT 103.780 141.050 104.630 141.900 ;
        RECT 105.340 142.415 105.700 142.795 ;
        RECT 105.970 142.415 106.330 142.795 ;
        RECT 106.570 142.415 106.930 142.795 ;
        RECT 105.340 141.825 105.700 142.205 ;
        RECT 105.970 141.825 106.330 142.205 ;
        RECT 106.570 141.825 106.930 142.205 ;
        RECT 100.430 140.100 101.280 140.950 ;
        RECT 101.380 140.100 102.230 140.950 ;
        RECT 102.830 140.100 103.680 140.950 ;
        RECT 103.780 140.100 104.630 140.950 ;
        RECT 100.430 139.050 101.280 139.900 ;
        RECT 101.380 139.050 102.230 139.900 ;
        RECT 102.830 139.050 103.680 139.900 ;
        RECT 103.780 139.050 104.630 139.900 ;
        RECT 103.780 138.100 104.630 138.950 ;
        RECT 4.830 136.650 5.680 137.500 ;
        RECT 23.780 136.650 24.630 137.500 ;
        RECT 24.830 136.650 25.680 137.500 ;
        RECT 43.780 136.650 44.630 137.500 ;
        RECT 44.830 136.650 45.680 137.500 ;
        RECT 63.780 136.650 64.630 137.500 ;
        RECT 64.830 136.650 65.680 137.500 ;
        RECT 83.780 136.650 84.630 137.500 ;
        RECT 84.830 136.650 85.680 137.500 ;
        RECT 103.780 136.650 104.630 137.500 ;
        RECT 4.830 135.700 5.680 136.550 ;
        RECT 23.780 135.700 24.630 136.550 ;
        RECT 24.830 135.700 25.680 136.550 ;
        RECT 43.780 135.700 44.630 136.550 ;
        RECT 44.830 135.700 45.680 136.550 ;
        RECT 63.780 135.700 64.630 136.550 ;
        RECT 64.830 135.700 65.680 136.550 ;
        RECT 83.780 135.700 84.630 136.550 ;
        RECT 84.830 135.700 85.680 136.550 ;
        RECT 103.780 135.700 104.630 136.550 ;
        RECT 105.340 136.830 105.700 137.210 ;
        RECT 105.970 136.830 106.330 137.210 ;
        RECT 106.570 136.830 106.930 137.210 ;
        RECT 105.340 136.240 105.700 136.620 ;
        RECT 105.970 136.240 106.330 136.620 ;
        RECT 106.570 136.240 106.930 136.620 ;
        RECT 2.520 134.920 2.880 135.300 ;
        RECT 3.130 134.920 3.490 135.300 ;
        RECT 3.760 134.920 4.120 135.300 ;
        RECT 2.520 134.185 2.880 134.565 ;
        RECT 3.130 134.185 3.490 134.565 ;
        RECT 3.760 134.185 4.120 134.565 ;
        RECT 2.520 133.500 2.880 133.880 ;
        RECT 3.130 133.500 3.490 133.880 ;
        RECT 3.760 133.500 4.120 133.880 ;
        RECT 2.520 126.120 2.880 126.500 ;
        RECT 3.130 126.120 3.490 126.500 ;
        RECT 3.760 126.120 4.120 126.500 ;
        RECT 2.520 125.385 2.880 125.765 ;
        RECT 3.130 125.385 3.490 125.765 ;
        RECT 3.760 125.385 4.120 125.765 ;
        RECT 2.520 124.700 2.880 125.080 ;
        RECT 3.130 124.700 3.490 125.080 ;
        RECT 3.760 124.700 4.120 125.080 ;
        RECT 4.830 123.450 5.680 124.300 ;
        RECT 23.780 123.450 24.630 124.300 ;
        RECT 24.830 123.450 25.680 124.300 ;
        RECT 43.780 123.450 44.630 124.300 ;
        RECT 44.830 123.450 45.680 124.300 ;
        RECT 63.780 123.450 64.630 124.300 ;
        RECT 64.830 123.450 65.680 124.300 ;
        RECT 83.780 123.450 84.630 124.300 ;
        RECT 84.830 123.450 85.680 124.300 ;
        RECT 103.780 123.450 104.630 124.300 ;
        RECT 2.515 122.750 2.875 123.130 ;
        RECT 3.145 122.750 3.505 123.130 ;
        RECT 3.745 122.750 4.105 123.130 ;
        RECT 2.515 122.160 2.875 122.540 ;
        RECT 3.145 122.160 3.505 122.540 ;
        RECT 3.745 122.160 4.105 122.540 ;
        RECT 4.830 122.500 5.680 123.350 ;
        RECT 23.780 122.500 24.630 123.350 ;
        RECT 24.830 122.500 25.680 123.350 ;
        RECT 43.780 122.500 44.630 123.350 ;
        RECT 44.830 122.500 45.680 123.350 ;
        RECT 63.780 122.500 64.630 123.350 ;
        RECT 64.830 122.500 65.680 123.350 ;
        RECT 83.780 122.500 84.630 123.350 ;
        RECT 84.830 122.500 85.680 123.350 ;
        RECT 103.780 122.500 104.630 123.350 ;
        RECT 4.830 121.050 5.680 121.900 ;
        RECT 4.830 120.100 5.680 120.950 ;
        RECT 5.780 120.100 6.630 120.950 ;
        RECT 7.230 120.100 8.080 120.950 ;
        RECT 8.180 120.100 9.030 120.950 ;
        RECT 4.830 119.050 5.680 119.900 ;
        RECT 5.780 119.050 6.630 119.900 ;
        RECT 7.230 119.050 8.080 119.900 ;
        RECT 8.180 119.050 9.030 119.900 ;
        RECT 4.830 118.100 5.680 118.950 ;
        RECT 23.780 121.050 24.630 121.900 ;
        RECT 24.830 121.050 25.680 121.900 ;
        RECT 20.430 120.100 21.280 120.950 ;
        RECT 21.380 120.100 22.230 120.950 ;
        RECT 22.830 120.100 23.680 120.950 ;
        RECT 23.780 120.100 24.630 120.950 ;
        RECT 24.830 120.100 25.680 120.950 ;
        RECT 25.780 120.100 26.630 120.950 ;
        RECT 27.230 120.100 28.080 120.950 ;
        RECT 28.180 120.100 29.030 120.950 ;
        RECT 20.430 119.050 21.280 119.900 ;
        RECT 21.380 119.050 22.230 119.900 ;
        RECT 22.830 119.050 23.680 119.900 ;
        RECT 23.780 119.050 24.630 119.900 ;
        RECT 24.830 119.050 25.680 119.900 ;
        RECT 25.780 119.050 26.630 119.900 ;
        RECT 27.230 119.050 28.080 119.900 ;
        RECT 28.180 119.050 29.030 119.900 ;
        RECT 23.780 118.100 24.630 118.950 ;
        RECT 24.830 118.100 25.680 118.950 ;
        RECT 43.780 121.050 44.630 121.900 ;
        RECT 44.830 121.050 45.680 121.900 ;
        RECT 40.430 120.100 41.280 120.950 ;
        RECT 41.380 120.100 42.230 120.950 ;
        RECT 42.830 120.100 43.680 120.950 ;
        RECT 43.780 120.100 44.630 120.950 ;
        RECT 44.830 120.100 45.680 120.950 ;
        RECT 45.780 120.100 46.630 120.950 ;
        RECT 47.230 120.100 48.080 120.950 ;
        RECT 48.180 120.100 49.030 120.950 ;
        RECT 40.430 119.050 41.280 119.900 ;
        RECT 41.380 119.050 42.230 119.900 ;
        RECT 42.830 119.050 43.680 119.900 ;
        RECT 43.780 119.050 44.630 119.900 ;
        RECT 44.830 119.050 45.680 119.900 ;
        RECT 45.780 119.050 46.630 119.900 ;
        RECT 47.230 119.050 48.080 119.900 ;
        RECT 48.180 119.050 49.030 119.900 ;
        RECT 43.780 118.100 44.630 118.950 ;
        RECT 44.830 118.100 45.680 118.950 ;
        RECT 63.780 121.050 64.630 121.900 ;
        RECT 64.830 121.050 65.680 121.900 ;
        RECT 60.430 120.100 61.280 120.950 ;
        RECT 61.380 120.100 62.230 120.950 ;
        RECT 62.830 120.100 63.680 120.950 ;
        RECT 63.780 120.100 64.630 120.950 ;
        RECT 64.830 120.100 65.680 120.950 ;
        RECT 65.780 120.100 66.630 120.950 ;
        RECT 67.230 120.100 68.080 120.950 ;
        RECT 68.180 120.100 69.030 120.950 ;
        RECT 60.430 119.050 61.280 119.900 ;
        RECT 61.380 119.050 62.230 119.900 ;
        RECT 62.830 119.050 63.680 119.900 ;
        RECT 63.780 119.050 64.630 119.900 ;
        RECT 64.830 119.050 65.680 119.900 ;
        RECT 65.780 119.050 66.630 119.900 ;
        RECT 67.230 119.050 68.080 119.900 ;
        RECT 68.180 119.050 69.030 119.900 ;
        RECT 63.780 118.100 64.630 118.950 ;
        RECT 64.830 118.100 65.680 118.950 ;
        RECT 83.780 121.050 84.630 121.900 ;
        RECT 84.830 121.050 85.680 121.900 ;
        RECT 80.430 120.100 81.280 120.950 ;
        RECT 81.380 120.100 82.230 120.950 ;
        RECT 82.830 120.100 83.680 120.950 ;
        RECT 83.780 120.100 84.630 120.950 ;
        RECT 84.830 120.100 85.680 120.950 ;
        RECT 85.780 120.100 86.630 120.950 ;
        RECT 87.230 120.100 88.080 120.950 ;
        RECT 88.180 120.100 89.030 120.950 ;
        RECT 80.430 119.050 81.280 119.900 ;
        RECT 81.380 119.050 82.230 119.900 ;
        RECT 82.830 119.050 83.680 119.900 ;
        RECT 83.780 119.050 84.630 119.900 ;
        RECT 84.830 119.050 85.680 119.900 ;
        RECT 85.780 119.050 86.630 119.900 ;
        RECT 87.230 119.050 88.080 119.900 ;
        RECT 88.180 119.050 89.030 119.900 ;
        RECT 83.780 118.100 84.630 118.950 ;
        RECT 84.830 118.100 85.680 118.950 ;
        RECT 103.780 121.050 104.630 121.900 ;
        RECT 105.340 122.615 105.700 122.995 ;
        RECT 105.970 122.615 106.330 122.995 ;
        RECT 106.570 122.615 106.930 122.995 ;
        RECT 105.340 122.025 105.700 122.405 ;
        RECT 105.970 122.025 106.330 122.405 ;
        RECT 106.570 122.025 106.930 122.405 ;
        RECT 100.430 120.100 101.280 120.950 ;
        RECT 101.380 120.100 102.230 120.950 ;
        RECT 102.830 120.100 103.680 120.950 ;
        RECT 103.780 120.100 104.630 120.950 ;
        RECT 100.430 119.050 101.280 119.900 ;
        RECT 101.380 119.050 102.230 119.900 ;
        RECT 102.830 119.050 103.680 119.900 ;
        RECT 103.780 119.050 104.630 119.900 ;
        RECT 103.780 118.100 104.630 118.950 ;
        RECT 2.515 117.340 2.875 117.720 ;
        RECT 3.145 117.340 3.505 117.720 ;
        RECT 3.745 117.340 4.105 117.720 ;
        RECT 2.515 116.750 2.875 117.130 ;
        RECT 3.145 116.750 3.505 117.130 ;
        RECT 3.745 116.750 4.105 117.130 ;
        RECT 4.830 116.650 5.680 117.500 ;
        RECT 23.780 116.650 24.630 117.500 ;
        RECT 24.830 116.650 25.680 117.500 ;
        RECT 43.780 116.650 44.630 117.500 ;
        RECT 44.830 116.650 45.680 117.500 ;
        RECT 63.780 116.650 64.630 117.500 ;
        RECT 64.830 116.650 65.680 117.500 ;
        RECT 83.780 116.650 84.630 117.500 ;
        RECT 84.830 116.650 85.680 117.500 ;
        RECT 103.780 116.650 104.630 117.500 ;
        RECT 4.830 115.700 5.680 116.550 ;
        RECT 23.780 115.700 24.630 116.550 ;
        RECT 24.830 115.700 25.680 116.550 ;
        RECT 43.780 115.700 44.630 116.550 ;
        RECT 44.830 115.700 45.680 116.550 ;
        RECT 63.780 115.700 64.630 116.550 ;
        RECT 64.830 115.700 65.680 116.550 ;
        RECT 83.780 115.700 84.630 116.550 ;
        RECT 84.830 115.700 85.680 116.550 ;
        RECT 103.780 115.700 104.630 116.550 ;
        RECT 105.340 116.740 105.700 117.120 ;
        RECT 105.970 116.740 106.330 117.120 ;
        RECT 106.570 116.740 106.930 117.120 ;
        RECT 105.340 116.150 105.700 116.530 ;
        RECT 105.970 116.150 106.330 116.530 ;
        RECT 106.570 116.150 106.930 116.530 ;
        RECT 2.520 114.920 2.880 115.300 ;
        RECT 3.130 114.920 3.490 115.300 ;
        RECT 3.760 114.920 4.120 115.300 ;
        RECT 2.520 114.185 2.880 114.565 ;
        RECT 3.130 114.185 3.490 114.565 ;
        RECT 3.760 114.185 4.120 114.565 ;
        RECT 2.520 113.500 2.880 113.880 ;
        RECT 3.130 113.500 3.490 113.880 ;
        RECT 3.760 113.500 4.120 113.880 ;
        RECT 2.520 106.125 2.880 106.505 ;
        RECT 3.130 106.125 3.490 106.505 ;
        RECT 3.760 106.125 4.120 106.505 ;
        RECT 2.520 105.390 2.880 105.770 ;
        RECT 3.130 105.390 3.490 105.770 ;
        RECT 3.760 105.390 4.120 105.770 ;
        RECT 2.520 104.705 2.880 105.085 ;
        RECT 3.130 104.705 3.490 105.085 ;
        RECT 3.760 104.705 4.120 105.085 ;
        RECT 2.515 102.965 2.875 103.345 ;
        RECT 3.145 102.965 3.505 103.345 ;
        RECT 3.745 102.965 4.105 103.345 ;
        RECT 2.515 102.375 2.875 102.755 ;
        RECT 3.145 102.375 3.505 102.755 ;
        RECT 3.745 102.375 4.105 102.755 ;
        RECT 4.830 103.450 5.680 104.300 ;
        RECT 23.780 103.450 24.630 104.300 ;
        RECT 24.830 103.450 25.680 104.300 ;
        RECT 43.780 103.450 44.630 104.300 ;
        RECT 44.830 103.450 45.680 104.300 ;
        RECT 63.780 103.450 64.630 104.300 ;
        RECT 64.830 103.450 65.680 104.300 ;
        RECT 83.780 103.450 84.630 104.300 ;
        RECT 84.830 103.450 85.680 104.300 ;
        RECT 103.780 103.450 104.630 104.300 ;
        RECT 4.830 102.500 5.680 103.350 ;
        RECT 23.780 102.500 24.630 103.350 ;
        RECT 24.830 102.500 25.680 103.350 ;
        RECT 43.780 102.500 44.630 103.350 ;
        RECT 44.830 102.500 45.680 103.350 ;
        RECT 63.780 102.500 64.630 103.350 ;
        RECT 64.830 102.500 65.680 103.350 ;
        RECT 83.780 102.500 84.630 103.350 ;
        RECT 84.830 102.500 85.680 103.350 ;
        RECT 103.780 102.500 104.630 103.350 ;
        RECT 4.830 101.050 5.680 101.900 ;
        RECT 4.830 100.100 5.680 100.950 ;
        RECT 5.780 100.100 6.630 100.950 ;
        RECT 7.230 100.100 8.080 100.950 ;
        RECT 8.180 100.100 9.030 100.950 ;
        RECT 4.830 99.050 5.680 99.900 ;
        RECT 5.780 99.050 6.630 99.900 ;
        RECT 7.230 99.050 8.080 99.900 ;
        RECT 8.180 99.050 9.030 99.900 ;
        RECT 4.830 98.100 5.680 98.950 ;
        RECT 23.780 101.050 24.630 101.900 ;
        RECT 24.830 101.050 25.680 101.900 ;
        RECT 20.430 100.100 21.280 100.950 ;
        RECT 21.380 100.100 22.230 100.950 ;
        RECT 22.830 100.100 23.680 100.950 ;
        RECT 23.780 100.100 24.630 100.950 ;
        RECT 24.830 100.100 25.680 100.950 ;
        RECT 25.780 100.100 26.630 100.950 ;
        RECT 27.230 100.100 28.080 100.950 ;
        RECT 28.180 100.100 29.030 100.950 ;
        RECT 20.430 99.050 21.280 99.900 ;
        RECT 21.380 99.050 22.230 99.900 ;
        RECT 22.830 99.050 23.680 99.900 ;
        RECT 23.780 99.050 24.630 99.900 ;
        RECT 24.830 99.050 25.680 99.900 ;
        RECT 25.780 99.050 26.630 99.900 ;
        RECT 27.230 99.050 28.080 99.900 ;
        RECT 28.180 99.050 29.030 99.900 ;
        RECT 23.780 98.100 24.630 98.950 ;
        RECT 24.830 98.100 25.680 98.950 ;
        RECT 43.780 101.050 44.630 101.900 ;
        RECT 44.830 101.050 45.680 101.900 ;
        RECT 40.430 100.100 41.280 100.950 ;
        RECT 41.380 100.100 42.230 100.950 ;
        RECT 42.830 100.100 43.680 100.950 ;
        RECT 43.780 100.100 44.630 100.950 ;
        RECT 44.830 100.100 45.680 100.950 ;
        RECT 45.780 100.100 46.630 100.950 ;
        RECT 47.230 100.100 48.080 100.950 ;
        RECT 48.180 100.100 49.030 100.950 ;
        RECT 40.430 99.050 41.280 99.900 ;
        RECT 41.380 99.050 42.230 99.900 ;
        RECT 42.830 99.050 43.680 99.900 ;
        RECT 43.780 99.050 44.630 99.900 ;
        RECT 44.830 99.050 45.680 99.900 ;
        RECT 45.780 99.050 46.630 99.900 ;
        RECT 47.230 99.050 48.080 99.900 ;
        RECT 48.180 99.050 49.030 99.900 ;
        RECT 43.780 98.100 44.630 98.950 ;
        RECT 44.830 98.100 45.680 98.950 ;
        RECT 63.780 101.050 64.630 101.900 ;
        RECT 64.830 101.050 65.680 101.900 ;
        RECT 60.430 100.100 61.280 100.950 ;
        RECT 61.380 100.100 62.230 100.950 ;
        RECT 62.830 100.100 63.680 100.950 ;
        RECT 63.780 100.100 64.630 100.950 ;
        RECT 64.830 100.100 65.680 100.950 ;
        RECT 65.780 100.100 66.630 100.950 ;
        RECT 67.230 100.100 68.080 100.950 ;
        RECT 68.180 100.100 69.030 100.950 ;
        RECT 60.430 99.050 61.280 99.900 ;
        RECT 61.380 99.050 62.230 99.900 ;
        RECT 62.830 99.050 63.680 99.900 ;
        RECT 63.780 99.050 64.630 99.900 ;
        RECT 64.830 99.050 65.680 99.900 ;
        RECT 65.780 99.050 66.630 99.900 ;
        RECT 67.230 99.050 68.080 99.900 ;
        RECT 68.180 99.050 69.030 99.900 ;
        RECT 63.780 98.100 64.630 98.950 ;
        RECT 64.830 98.100 65.680 98.950 ;
        RECT 83.780 101.050 84.630 101.900 ;
        RECT 84.830 101.050 85.680 101.900 ;
        RECT 80.430 100.100 81.280 100.950 ;
        RECT 81.380 100.100 82.230 100.950 ;
        RECT 82.830 100.100 83.680 100.950 ;
        RECT 83.780 100.100 84.630 100.950 ;
        RECT 84.830 100.100 85.680 100.950 ;
        RECT 85.780 100.100 86.630 100.950 ;
        RECT 87.230 100.100 88.080 100.950 ;
        RECT 88.180 100.100 89.030 100.950 ;
        RECT 80.430 99.050 81.280 99.900 ;
        RECT 81.380 99.050 82.230 99.900 ;
        RECT 82.830 99.050 83.680 99.900 ;
        RECT 83.780 99.050 84.630 99.900 ;
        RECT 84.830 99.050 85.680 99.900 ;
        RECT 85.780 99.050 86.630 99.900 ;
        RECT 87.230 99.050 88.080 99.900 ;
        RECT 88.180 99.050 89.030 99.900 ;
        RECT 83.780 98.100 84.630 98.950 ;
        RECT 84.830 98.100 85.680 98.950 ;
        RECT 103.780 101.050 104.630 101.900 ;
        RECT 105.340 102.535 105.700 102.915 ;
        RECT 105.970 102.535 106.330 102.915 ;
        RECT 106.570 102.535 106.930 102.915 ;
        RECT 105.340 101.945 105.700 102.325 ;
        RECT 105.970 101.945 106.330 102.325 ;
        RECT 106.570 101.945 106.930 102.325 ;
        RECT 100.430 100.100 101.280 100.950 ;
        RECT 101.380 100.100 102.230 100.950 ;
        RECT 102.830 100.100 103.680 100.950 ;
        RECT 103.780 100.100 104.630 100.950 ;
        RECT 100.430 99.050 101.280 99.900 ;
        RECT 101.380 99.050 102.230 99.900 ;
        RECT 102.830 99.050 103.680 99.900 ;
        RECT 103.780 99.050 104.630 99.900 ;
        RECT 103.780 98.100 104.630 98.950 ;
        RECT 2.515 97.460 2.875 97.840 ;
        RECT 3.145 97.460 3.505 97.840 ;
        RECT 3.745 97.460 4.105 97.840 ;
        RECT 2.515 96.870 2.875 97.250 ;
        RECT 3.145 96.870 3.505 97.250 ;
        RECT 3.745 96.870 4.105 97.250 ;
        RECT 4.830 96.650 5.680 97.500 ;
        RECT 23.780 96.650 24.630 97.500 ;
        RECT 24.830 96.650 25.680 97.500 ;
        RECT 43.780 96.650 44.630 97.500 ;
        RECT 44.830 96.650 45.680 97.500 ;
        RECT 63.780 96.650 64.630 97.500 ;
        RECT 64.830 96.650 65.680 97.500 ;
        RECT 83.780 96.650 84.630 97.500 ;
        RECT 84.830 96.650 85.680 97.500 ;
        RECT 103.780 96.650 104.630 97.500 ;
        RECT 4.830 95.700 5.680 96.550 ;
        RECT 23.780 95.700 24.630 96.550 ;
        RECT 24.830 95.700 25.680 96.550 ;
        RECT 43.780 95.700 44.630 96.550 ;
        RECT 44.830 95.700 45.680 96.550 ;
        RECT 63.780 95.700 64.630 96.550 ;
        RECT 64.830 95.700 65.680 96.550 ;
        RECT 83.780 95.700 84.630 96.550 ;
        RECT 84.830 95.700 85.680 96.550 ;
        RECT 103.780 95.700 104.630 96.550 ;
        RECT 105.340 96.680 105.700 97.060 ;
        RECT 105.970 96.680 106.330 97.060 ;
        RECT 106.570 96.680 106.930 97.060 ;
        RECT 105.340 96.090 105.700 96.470 ;
        RECT 105.970 96.090 106.330 96.470 ;
        RECT 106.570 96.090 106.930 96.470 ;
        RECT 2.520 94.920 2.880 95.300 ;
        RECT 3.130 94.920 3.490 95.300 ;
        RECT 3.760 94.920 4.120 95.300 ;
        RECT 2.520 94.185 2.880 94.565 ;
        RECT 3.130 94.185 3.490 94.565 ;
        RECT 3.760 94.185 4.120 94.565 ;
        RECT 2.520 93.500 2.880 93.880 ;
        RECT 3.130 93.500 3.490 93.880 ;
        RECT 3.760 93.500 4.120 93.880 ;
        RECT 2.520 86.120 2.880 86.500 ;
        RECT 3.130 86.120 3.490 86.500 ;
        RECT 3.760 86.120 4.120 86.500 ;
        RECT 2.520 85.385 2.880 85.765 ;
        RECT 3.130 85.385 3.490 85.765 ;
        RECT 3.760 85.385 4.120 85.765 ;
        RECT 2.520 84.700 2.880 85.080 ;
        RECT 3.130 84.700 3.490 85.080 ;
        RECT 3.760 84.700 4.120 85.080 ;
        RECT 2.515 83.130 2.875 83.510 ;
        RECT 3.145 83.130 3.505 83.510 ;
        RECT 3.745 83.130 4.105 83.510 ;
        RECT 2.515 82.540 2.875 82.920 ;
        RECT 3.145 82.540 3.505 82.920 ;
        RECT 3.745 82.540 4.105 82.920 ;
        RECT 4.830 83.450 5.680 84.300 ;
        RECT 23.780 83.450 24.630 84.300 ;
        RECT 24.830 83.450 25.680 84.300 ;
        RECT 43.780 83.450 44.630 84.300 ;
        RECT 44.830 83.450 45.680 84.300 ;
        RECT 63.780 83.450 64.630 84.300 ;
        RECT 64.830 83.450 65.680 84.300 ;
        RECT 83.780 83.450 84.630 84.300 ;
        RECT 84.830 83.450 85.680 84.300 ;
        RECT 103.780 83.450 104.630 84.300 ;
        RECT 4.830 82.500 5.680 83.350 ;
        RECT 23.780 82.500 24.630 83.350 ;
        RECT 24.830 82.500 25.680 83.350 ;
        RECT 43.780 82.500 44.630 83.350 ;
        RECT 44.830 82.500 45.680 83.350 ;
        RECT 63.780 82.500 64.630 83.350 ;
        RECT 64.830 82.500 65.680 83.350 ;
        RECT 83.780 82.500 84.630 83.350 ;
        RECT 84.830 82.500 85.680 83.350 ;
        RECT 103.780 82.500 104.630 83.350 ;
        RECT 105.340 82.875 105.700 83.255 ;
        RECT 105.970 82.875 106.330 83.255 ;
        RECT 106.570 82.875 106.930 83.255 ;
        RECT 105.340 82.285 105.700 82.665 ;
        RECT 105.970 82.285 106.330 82.665 ;
        RECT 106.570 82.285 106.930 82.665 ;
        RECT 4.830 81.050 5.680 81.900 ;
        RECT 4.830 80.100 5.680 80.950 ;
        RECT 5.780 80.100 6.630 80.950 ;
        RECT 7.230 80.100 8.080 80.950 ;
        RECT 8.180 80.100 9.030 80.950 ;
        RECT 4.830 79.050 5.680 79.900 ;
        RECT 5.780 79.050 6.630 79.900 ;
        RECT 7.230 79.050 8.080 79.900 ;
        RECT 8.180 79.050 9.030 79.900 ;
        RECT 4.830 78.100 5.680 78.950 ;
        RECT 23.780 81.050 24.630 81.900 ;
        RECT 24.830 81.050 25.680 81.900 ;
        RECT 20.430 80.100 21.280 80.950 ;
        RECT 21.380 80.100 22.230 80.950 ;
        RECT 22.830 80.100 23.680 80.950 ;
        RECT 23.780 80.100 24.630 80.950 ;
        RECT 24.830 80.100 25.680 80.950 ;
        RECT 25.780 80.100 26.630 80.950 ;
        RECT 27.230 80.100 28.080 80.950 ;
        RECT 28.180 80.100 29.030 80.950 ;
        RECT 20.430 79.050 21.280 79.900 ;
        RECT 21.380 79.050 22.230 79.900 ;
        RECT 22.830 79.050 23.680 79.900 ;
        RECT 23.780 79.050 24.630 79.900 ;
        RECT 24.830 79.050 25.680 79.900 ;
        RECT 25.780 79.050 26.630 79.900 ;
        RECT 27.230 79.050 28.080 79.900 ;
        RECT 28.180 79.050 29.030 79.900 ;
        RECT 23.780 78.100 24.630 78.950 ;
        RECT 24.830 78.100 25.680 78.950 ;
        RECT 43.780 81.050 44.630 81.900 ;
        RECT 44.830 81.050 45.680 81.900 ;
        RECT 40.430 80.100 41.280 80.950 ;
        RECT 41.380 80.100 42.230 80.950 ;
        RECT 42.830 80.100 43.680 80.950 ;
        RECT 43.780 80.100 44.630 80.950 ;
        RECT 44.830 80.100 45.680 80.950 ;
        RECT 45.780 80.100 46.630 80.950 ;
        RECT 47.230 80.100 48.080 80.950 ;
        RECT 48.180 80.100 49.030 80.950 ;
        RECT 40.430 79.050 41.280 79.900 ;
        RECT 41.380 79.050 42.230 79.900 ;
        RECT 42.830 79.050 43.680 79.900 ;
        RECT 43.780 79.050 44.630 79.900 ;
        RECT 44.830 79.050 45.680 79.900 ;
        RECT 45.780 79.050 46.630 79.900 ;
        RECT 47.230 79.050 48.080 79.900 ;
        RECT 48.180 79.050 49.030 79.900 ;
        RECT 43.780 78.100 44.630 78.950 ;
        RECT 44.830 78.100 45.680 78.950 ;
        RECT 63.780 81.050 64.630 81.900 ;
        RECT 64.830 81.050 65.680 81.900 ;
        RECT 60.430 80.100 61.280 80.950 ;
        RECT 61.380 80.100 62.230 80.950 ;
        RECT 62.830 80.100 63.680 80.950 ;
        RECT 63.780 80.100 64.630 80.950 ;
        RECT 64.830 80.100 65.680 80.950 ;
        RECT 65.780 80.100 66.630 80.950 ;
        RECT 67.230 80.100 68.080 80.950 ;
        RECT 68.180 80.100 69.030 80.950 ;
        RECT 60.430 79.050 61.280 79.900 ;
        RECT 61.380 79.050 62.230 79.900 ;
        RECT 62.830 79.050 63.680 79.900 ;
        RECT 63.780 79.050 64.630 79.900 ;
        RECT 64.830 79.050 65.680 79.900 ;
        RECT 65.780 79.050 66.630 79.900 ;
        RECT 67.230 79.050 68.080 79.900 ;
        RECT 68.180 79.050 69.030 79.900 ;
        RECT 63.780 78.100 64.630 78.950 ;
        RECT 64.830 78.100 65.680 78.950 ;
        RECT 83.780 81.050 84.630 81.900 ;
        RECT 84.830 81.050 85.680 81.900 ;
        RECT 80.430 80.100 81.280 80.950 ;
        RECT 81.380 80.100 82.230 80.950 ;
        RECT 82.830 80.100 83.680 80.950 ;
        RECT 83.780 80.100 84.630 80.950 ;
        RECT 84.830 80.100 85.680 80.950 ;
        RECT 85.780 80.100 86.630 80.950 ;
        RECT 87.230 80.100 88.080 80.950 ;
        RECT 88.180 80.100 89.030 80.950 ;
        RECT 80.430 79.050 81.280 79.900 ;
        RECT 81.380 79.050 82.230 79.900 ;
        RECT 82.830 79.050 83.680 79.900 ;
        RECT 83.780 79.050 84.630 79.900 ;
        RECT 84.830 79.050 85.680 79.900 ;
        RECT 85.780 79.050 86.630 79.900 ;
        RECT 87.230 79.050 88.080 79.900 ;
        RECT 88.180 79.050 89.030 79.900 ;
        RECT 83.780 78.100 84.630 78.950 ;
        RECT 84.830 78.100 85.680 78.950 ;
        RECT 103.780 81.050 104.630 81.900 ;
        RECT 100.430 80.100 101.280 80.950 ;
        RECT 101.380 80.100 102.230 80.950 ;
        RECT 102.830 80.100 103.680 80.950 ;
        RECT 103.780 80.100 104.630 80.950 ;
        RECT 100.430 79.050 101.280 79.900 ;
        RECT 101.380 79.050 102.230 79.900 ;
        RECT 102.830 79.050 103.680 79.900 ;
        RECT 103.780 79.050 104.630 79.900 ;
        RECT 103.780 78.100 104.630 78.950 ;
        RECT 2.515 77.050 2.875 77.430 ;
        RECT 3.145 77.050 3.505 77.430 ;
        RECT 3.745 77.050 4.105 77.430 ;
        RECT 2.515 76.460 2.875 76.840 ;
        RECT 3.145 76.460 3.505 76.840 ;
        RECT 3.745 76.460 4.105 76.840 ;
        RECT 4.830 76.650 5.680 77.500 ;
        RECT 23.780 76.650 24.630 77.500 ;
        RECT 24.830 76.650 25.680 77.500 ;
        RECT 43.780 76.650 44.630 77.500 ;
        RECT 44.830 76.650 45.680 77.500 ;
        RECT 63.780 76.650 64.630 77.500 ;
        RECT 64.830 76.650 65.680 77.500 ;
        RECT 83.780 76.650 84.630 77.500 ;
        RECT 84.830 76.650 85.680 77.500 ;
        RECT 103.780 76.650 104.630 77.500 ;
        RECT 4.830 75.700 5.680 76.550 ;
        RECT 23.780 75.700 24.630 76.550 ;
        RECT 24.830 75.700 25.680 76.550 ;
        RECT 43.780 75.700 44.630 76.550 ;
        RECT 44.830 75.700 45.680 76.550 ;
        RECT 63.780 75.700 64.630 76.550 ;
        RECT 64.830 75.700 65.680 76.550 ;
        RECT 83.780 75.700 84.630 76.550 ;
        RECT 84.830 75.700 85.680 76.550 ;
        RECT 103.780 75.700 104.630 76.550 ;
        RECT 105.340 76.805 105.700 77.185 ;
        RECT 105.970 76.805 106.330 77.185 ;
        RECT 106.570 76.805 106.930 77.185 ;
        RECT 105.340 76.215 105.700 76.595 ;
        RECT 105.970 76.215 106.330 76.595 ;
        RECT 106.570 76.215 106.930 76.595 ;
        RECT 2.520 74.920 2.880 75.300 ;
        RECT 3.130 74.920 3.490 75.300 ;
        RECT 3.760 74.920 4.120 75.300 ;
        RECT 2.520 74.185 2.880 74.565 ;
        RECT 3.130 74.185 3.490 74.565 ;
        RECT 3.760 74.185 4.120 74.565 ;
        RECT 2.520 73.500 2.880 73.880 ;
        RECT 3.130 73.500 3.490 73.880 ;
        RECT 3.760 73.500 4.120 73.880 ;
        RECT 2.520 66.120 2.880 66.500 ;
        RECT 3.130 66.120 3.490 66.500 ;
        RECT 3.760 66.120 4.120 66.500 ;
        RECT 2.520 65.385 2.880 65.765 ;
        RECT 3.130 65.385 3.490 65.765 ;
        RECT 3.760 65.385 4.120 65.765 ;
        RECT 2.520 64.700 2.880 65.080 ;
        RECT 3.130 64.700 3.490 65.080 ;
        RECT 3.760 64.700 4.120 65.080 ;
        RECT 4.830 63.450 5.680 64.300 ;
        RECT 23.780 63.450 24.630 64.300 ;
        RECT 24.830 63.450 25.680 64.300 ;
        RECT 43.780 63.450 44.630 64.300 ;
        RECT 44.830 63.450 45.680 64.300 ;
        RECT 63.780 63.450 64.630 64.300 ;
        RECT 64.830 63.450 65.680 64.300 ;
        RECT 83.780 63.450 84.630 64.300 ;
        RECT 84.830 63.450 85.680 64.300 ;
        RECT 103.780 63.450 104.630 64.300 ;
        RECT 2.515 62.725 2.875 63.105 ;
        RECT 3.145 62.725 3.505 63.105 ;
        RECT 3.745 62.725 4.105 63.105 ;
        RECT 2.515 62.135 2.875 62.515 ;
        RECT 3.145 62.135 3.505 62.515 ;
        RECT 3.745 62.135 4.105 62.515 ;
        RECT 4.830 62.500 5.680 63.350 ;
        RECT 23.780 62.500 24.630 63.350 ;
        RECT 24.830 62.500 25.680 63.350 ;
        RECT 43.780 62.500 44.630 63.350 ;
        RECT 44.830 62.500 45.680 63.350 ;
        RECT 63.780 62.500 64.630 63.350 ;
        RECT 64.830 62.500 65.680 63.350 ;
        RECT 83.780 62.500 84.630 63.350 ;
        RECT 84.830 62.500 85.680 63.350 ;
        RECT 103.780 62.500 104.630 63.350 ;
        RECT 4.830 61.050 5.680 61.900 ;
        RECT 4.830 60.100 5.680 60.950 ;
        RECT 5.780 60.100 6.630 60.950 ;
        RECT 7.230 60.100 8.080 60.950 ;
        RECT 8.180 60.100 9.030 60.950 ;
        RECT 4.830 59.050 5.680 59.900 ;
        RECT 5.780 59.050 6.630 59.900 ;
        RECT 7.230 59.050 8.080 59.900 ;
        RECT 8.180 59.050 9.030 59.900 ;
        RECT 4.830 58.100 5.680 58.950 ;
        RECT 23.780 61.050 24.630 61.900 ;
        RECT 24.830 61.050 25.680 61.900 ;
        RECT 20.430 60.100 21.280 60.950 ;
        RECT 21.380 60.100 22.230 60.950 ;
        RECT 22.830 60.100 23.680 60.950 ;
        RECT 23.780 60.100 24.630 60.950 ;
        RECT 24.830 60.100 25.680 60.950 ;
        RECT 25.780 60.100 26.630 60.950 ;
        RECT 27.230 60.100 28.080 60.950 ;
        RECT 28.180 60.100 29.030 60.950 ;
        RECT 20.430 59.050 21.280 59.900 ;
        RECT 21.380 59.050 22.230 59.900 ;
        RECT 22.830 59.050 23.680 59.900 ;
        RECT 23.780 59.050 24.630 59.900 ;
        RECT 24.830 59.050 25.680 59.900 ;
        RECT 25.780 59.050 26.630 59.900 ;
        RECT 27.230 59.050 28.080 59.900 ;
        RECT 28.180 59.050 29.030 59.900 ;
        RECT 23.780 58.100 24.630 58.950 ;
        RECT 24.830 58.100 25.680 58.950 ;
        RECT 43.780 61.050 44.630 61.900 ;
        RECT 44.830 61.050 45.680 61.900 ;
        RECT 40.430 60.100 41.280 60.950 ;
        RECT 41.380 60.100 42.230 60.950 ;
        RECT 42.830 60.100 43.680 60.950 ;
        RECT 43.780 60.100 44.630 60.950 ;
        RECT 44.830 60.100 45.680 60.950 ;
        RECT 45.780 60.100 46.630 60.950 ;
        RECT 47.230 60.100 48.080 60.950 ;
        RECT 48.180 60.100 49.030 60.950 ;
        RECT 40.430 59.050 41.280 59.900 ;
        RECT 41.380 59.050 42.230 59.900 ;
        RECT 42.830 59.050 43.680 59.900 ;
        RECT 43.780 59.050 44.630 59.900 ;
        RECT 44.830 59.050 45.680 59.900 ;
        RECT 45.780 59.050 46.630 59.900 ;
        RECT 47.230 59.050 48.080 59.900 ;
        RECT 48.180 59.050 49.030 59.900 ;
        RECT 43.780 58.100 44.630 58.950 ;
        RECT 44.830 58.100 45.680 58.950 ;
        RECT 63.780 61.050 64.630 61.900 ;
        RECT 64.830 61.050 65.680 61.900 ;
        RECT 60.430 60.100 61.280 60.950 ;
        RECT 61.380 60.100 62.230 60.950 ;
        RECT 62.830 60.100 63.680 60.950 ;
        RECT 63.780 60.100 64.630 60.950 ;
        RECT 64.830 60.100 65.680 60.950 ;
        RECT 65.780 60.100 66.630 60.950 ;
        RECT 67.230 60.100 68.080 60.950 ;
        RECT 68.180 60.100 69.030 60.950 ;
        RECT 60.430 59.050 61.280 59.900 ;
        RECT 61.380 59.050 62.230 59.900 ;
        RECT 62.830 59.050 63.680 59.900 ;
        RECT 63.780 59.050 64.630 59.900 ;
        RECT 64.830 59.050 65.680 59.900 ;
        RECT 65.780 59.050 66.630 59.900 ;
        RECT 67.230 59.050 68.080 59.900 ;
        RECT 68.180 59.050 69.030 59.900 ;
        RECT 63.780 58.100 64.630 58.950 ;
        RECT 64.830 58.100 65.680 58.950 ;
        RECT 83.780 61.050 84.630 61.900 ;
        RECT 84.830 61.050 85.680 61.900 ;
        RECT 80.430 60.100 81.280 60.950 ;
        RECT 81.380 60.100 82.230 60.950 ;
        RECT 82.830 60.100 83.680 60.950 ;
        RECT 83.780 60.100 84.630 60.950 ;
        RECT 84.830 60.100 85.680 60.950 ;
        RECT 85.780 60.100 86.630 60.950 ;
        RECT 87.230 60.100 88.080 60.950 ;
        RECT 88.180 60.100 89.030 60.950 ;
        RECT 80.430 59.050 81.280 59.900 ;
        RECT 81.380 59.050 82.230 59.900 ;
        RECT 82.830 59.050 83.680 59.900 ;
        RECT 83.780 59.050 84.630 59.900 ;
        RECT 84.830 59.050 85.680 59.900 ;
        RECT 85.780 59.050 86.630 59.900 ;
        RECT 87.230 59.050 88.080 59.900 ;
        RECT 88.180 59.050 89.030 59.900 ;
        RECT 83.780 58.100 84.630 58.950 ;
        RECT 84.830 58.100 85.680 58.950 ;
        RECT 103.780 61.050 104.630 61.900 ;
        RECT 105.340 62.590 105.700 62.970 ;
        RECT 105.970 62.590 106.330 62.970 ;
        RECT 106.570 62.590 106.930 62.970 ;
        RECT 105.340 62.000 105.700 62.380 ;
        RECT 105.970 62.000 106.330 62.380 ;
        RECT 106.570 62.000 106.930 62.380 ;
        RECT 100.430 60.100 101.280 60.950 ;
        RECT 101.380 60.100 102.230 60.950 ;
        RECT 102.830 60.100 103.680 60.950 ;
        RECT 103.780 60.100 104.630 60.950 ;
        RECT 100.430 59.050 101.280 59.900 ;
        RECT 101.380 59.050 102.230 59.900 ;
        RECT 102.830 59.050 103.680 59.900 ;
        RECT 103.780 59.050 104.630 59.900 ;
        RECT 103.780 58.100 104.630 58.950 ;
        RECT 2.515 57.115 2.875 57.495 ;
        RECT 3.145 57.115 3.505 57.495 ;
        RECT 3.745 57.115 4.105 57.495 ;
        RECT 2.515 56.525 2.875 56.905 ;
        RECT 3.145 56.525 3.505 56.905 ;
        RECT 3.745 56.525 4.105 56.905 ;
        RECT 4.830 56.650 5.680 57.500 ;
        RECT 23.780 56.650 24.630 57.500 ;
        RECT 24.830 56.650 25.680 57.500 ;
        RECT 43.780 56.650 44.630 57.500 ;
        RECT 44.830 56.650 45.680 57.500 ;
        RECT 63.780 56.650 64.630 57.500 ;
        RECT 64.830 56.650 65.680 57.500 ;
        RECT 83.780 56.650 84.630 57.500 ;
        RECT 84.830 56.650 85.680 57.500 ;
        RECT 103.780 56.650 104.630 57.500 ;
        RECT 4.830 55.700 5.680 56.550 ;
        RECT 23.780 55.700 24.630 56.550 ;
        RECT 24.830 55.700 25.680 56.550 ;
        RECT 43.780 55.700 44.630 56.550 ;
        RECT 44.830 55.700 45.680 56.550 ;
        RECT 63.780 55.700 64.630 56.550 ;
        RECT 64.830 55.700 65.680 56.550 ;
        RECT 83.780 55.700 84.630 56.550 ;
        RECT 84.830 55.700 85.680 56.550 ;
        RECT 103.780 55.700 104.630 56.550 ;
        RECT 105.340 56.805 105.700 57.185 ;
        RECT 105.970 56.805 106.330 57.185 ;
        RECT 106.570 56.805 106.930 57.185 ;
        RECT 105.340 56.215 105.700 56.595 ;
        RECT 105.970 56.215 106.330 56.595 ;
        RECT 106.570 56.215 106.930 56.595 ;
        RECT 2.520 54.925 2.880 55.305 ;
        RECT 3.130 54.925 3.490 55.305 ;
        RECT 3.760 54.925 4.120 55.305 ;
        RECT 2.520 54.190 2.880 54.570 ;
        RECT 3.130 54.190 3.490 54.570 ;
        RECT 3.760 54.190 4.120 54.570 ;
        RECT 2.520 53.505 2.880 53.885 ;
        RECT 3.130 53.505 3.490 53.885 ;
        RECT 3.760 53.505 4.120 53.885 ;
        RECT 2.520 46.115 2.880 46.495 ;
        RECT 3.130 46.115 3.490 46.495 ;
        RECT 3.760 46.115 4.120 46.495 ;
        RECT 2.520 45.380 2.880 45.760 ;
        RECT 3.130 45.380 3.490 45.760 ;
        RECT 3.760 45.380 4.120 45.760 ;
        RECT 2.520 44.695 2.880 45.075 ;
        RECT 3.130 44.695 3.490 45.075 ;
        RECT 3.760 44.695 4.120 45.075 ;
        RECT 4.830 43.450 5.680 44.300 ;
        RECT 23.780 43.450 24.630 44.300 ;
        RECT 24.830 43.450 25.680 44.300 ;
        RECT 43.780 43.450 44.630 44.300 ;
        RECT 44.830 43.450 45.680 44.300 ;
        RECT 63.780 43.450 64.630 44.300 ;
        RECT 64.830 43.450 65.680 44.300 ;
        RECT 83.780 43.450 84.630 44.300 ;
        RECT 84.830 43.450 85.680 44.300 ;
        RECT 103.780 43.450 104.630 44.300 ;
        RECT 2.515 42.815 2.875 43.195 ;
        RECT 3.145 42.815 3.505 43.195 ;
        RECT 3.745 42.815 4.105 43.195 ;
        RECT 2.515 42.225 2.875 42.605 ;
        RECT 3.145 42.225 3.505 42.605 ;
        RECT 3.745 42.225 4.105 42.605 ;
        RECT 4.830 42.500 5.680 43.350 ;
        RECT 23.780 42.500 24.630 43.350 ;
        RECT 24.830 42.500 25.680 43.350 ;
        RECT 43.780 42.500 44.630 43.350 ;
        RECT 44.830 42.500 45.680 43.350 ;
        RECT 63.780 42.500 64.630 43.350 ;
        RECT 64.830 42.500 65.680 43.350 ;
        RECT 83.780 42.500 84.630 43.350 ;
        RECT 84.830 42.500 85.680 43.350 ;
        RECT 103.780 42.500 104.630 43.350 ;
        RECT 4.830 41.050 5.680 41.900 ;
        RECT 4.830 40.100 5.680 40.950 ;
        RECT 5.780 40.100 6.630 40.950 ;
        RECT 7.230 40.100 8.080 40.950 ;
        RECT 8.180 40.100 9.030 40.950 ;
        RECT 4.830 39.050 5.680 39.900 ;
        RECT 5.780 39.050 6.630 39.900 ;
        RECT 7.230 39.050 8.080 39.900 ;
        RECT 8.180 39.050 9.030 39.900 ;
        RECT 4.830 38.100 5.680 38.950 ;
        RECT 23.780 41.050 24.630 41.900 ;
        RECT 24.830 41.050 25.680 41.900 ;
        RECT 20.430 40.100 21.280 40.950 ;
        RECT 21.380 40.100 22.230 40.950 ;
        RECT 22.830 40.100 23.680 40.950 ;
        RECT 23.780 40.100 24.630 40.950 ;
        RECT 24.830 40.100 25.680 40.950 ;
        RECT 25.780 40.100 26.630 40.950 ;
        RECT 27.230 40.100 28.080 40.950 ;
        RECT 28.180 40.100 29.030 40.950 ;
        RECT 20.430 39.050 21.280 39.900 ;
        RECT 21.380 39.050 22.230 39.900 ;
        RECT 22.830 39.050 23.680 39.900 ;
        RECT 23.780 39.050 24.630 39.900 ;
        RECT 24.830 39.050 25.680 39.900 ;
        RECT 25.780 39.050 26.630 39.900 ;
        RECT 27.230 39.050 28.080 39.900 ;
        RECT 28.180 39.050 29.030 39.900 ;
        RECT 23.780 38.100 24.630 38.950 ;
        RECT 24.830 38.100 25.680 38.950 ;
        RECT 43.780 41.050 44.630 41.900 ;
        RECT 44.830 41.050 45.680 41.900 ;
        RECT 40.430 40.100 41.280 40.950 ;
        RECT 41.380 40.100 42.230 40.950 ;
        RECT 42.830 40.100 43.680 40.950 ;
        RECT 43.780 40.100 44.630 40.950 ;
        RECT 44.830 40.100 45.680 40.950 ;
        RECT 45.780 40.100 46.630 40.950 ;
        RECT 47.230 40.100 48.080 40.950 ;
        RECT 48.180 40.100 49.030 40.950 ;
        RECT 40.430 39.050 41.280 39.900 ;
        RECT 41.380 39.050 42.230 39.900 ;
        RECT 42.830 39.050 43.680 39.900 ;
        RECT 43.780 39.050 44.630 39.900 ;
        RECT 44.830 39.050 45.680 39.900 ;
        RECT 45.780 39.050 46.630 39.900 ;
        RECT 47.230 39.050 48.080 39.900 ;
        RECT 48.180 39.050 49.030 39.900 ;
        RECT 43.780 38.100 44.630 38.950 ;
        RECT 44.830 38.100 45.680 38.950 ;
        RECT 63.780 41.050 64.630 41.900 ;
        RECT 64.830 41.050 65.680 41.900 ;
        RECT 60.430 40.100 61.280 40.950 ;
        RECT 61.380 40.100 62.230 40.950 ;
        RECT 62.830 40.100 63.680 40.950 ;
        RECT 63.780 40.100 64.630 40.950 ;
        RECT 64.830 40.100 65.680 40.950 ;
        RECT 65.780 40.100 66.630 40.950 ;
        RECT 67.230 40.100 68.080 40.950 ;
        RECT 68.180 40.100 69.030 40.950 ;
        RECT 60.430 39.050 61.280 39.900 ;
        RECT 61.380 39.050 62.230 39.900 ;
        RECT 62.830 39.050 63.680 39.900 ;
        RECT 63.780 39.050 64.630 39.900 ;
        RECT 64.830 39.050 65.680 39.900 ;
        RECT 65.780 39.050 66.630 39.900 ;
        RECT 67.230 39.050 68.080 39.900 ;
        RECT 68.180 39.050 69.030 39.900 ;
        RECT 63.780 38.100 64.630 38.950 ;
        RECT 64.830 38.100 65.680 38.950 ;
        RECT 83.780 41.050 84.630 41.900 ;
        RECT 84.830 41.050 85.680 41.900 ;
        RECT 80.430 40.100 81.280 40.950 ;
        RECT 81.380 40.100 82.230 40.950 ;
        RECT 82.830 40.100 83.680 40.950 ;
        RECT 83.780 40.100 84.630 40.950 ;
        RECT 84.830 40.100 85.680 40.950 ;
        RECT 85.780 40.100 86.630 40.950 ;
        RECT 87.230 40.100 88.080 40.950 ;
        RECT 88.180 40.100 89.030 40.950 ;
        RECT 80.430 39.050 81.280 39.900 ;
        RECT 81.380 39.050 82.230 39.900 ;
        RECT 82.830 39.050 83.680 39.900 ;
        RECT 83.780 39.050 84.630 39.900 ;
        RECT 84.830 39.050 85.680 39.900 ;
        RECT 85.780 39.050 86.630 39.900 ;
        RECT 87.230 39.050 88.080 39.900 ;
        RECT 88.180 39.050 89.030 39.900 ;
        RECT 83.780 38.100 84.630 38.950 ;
        RECT 84.830 38.100 85.680 38.950 ;
        RECT 103.780 41.050 104.630 41.900 ;
        RECT 105.340 42.590 105.700 42.970 ;
        RECT 105.970 42.590 106.330 42.970 ;
        RECT 106.570 42.590 106.930 42.970 ;
        RECT 105.340 42.000 105.700 42.380 ;
        RECT 105.970 42.000 106.330 42.380 ;
        RECT 106.570 42.000 106.930 42.380 ;
        RECT 100.430 40.100 101.280 40.950 ;
        RECT 101.380 40.100 102.230 40.950 ;
        RECT 102.830 40.100 103.680 40.950 ;
        RECT 103.780 40.100 104.630 40.950 ;
        RECT 100.430 39.050 101.280 39.900 ;
        RECT 101.380 39.050 102.230 39.900 ;
        RECT 102.830 39.050 103.680 39.900 ;
        RECT 103.780 39.050 104.630 39.900 ;
        RECT 103.780 38.100 104.630 38.950 ;
        RECT 2.515 37.260 2.875 37.640 ;
        RECT 3.145 37.260 3.505 37.640 ;
        RECT 3.745 37.260 4.105 37.640 ;
        RECT 2.515 36.670 2.875 37.050 ;
        RECT 3.145 36.670 3.505 37.050 ;
        RECT 3.745 36.670 4.105 37.050 ;
        RECT 4.830 36.650 5.680 37.500 ;
        RECT 23.780 36.650 24.630 37.500 ;
        RECT 24.830 36.650 25.680 37.500 ;
        RECT 43.780 36.650 44.630 37.500 ;
        RECT 44.830 36.650 45.680 37.500 ;
        RECT 63.780 36.650 64.630 37.500 ;
        RECT 64.830 36.650 65.680 37.500 ;
        RECT 83.780 36.650 84.630 37.500 ;
        RECT 84.830 36.650 85.680 37.500 ;
        RECT 103.780 36.650 104.630 37.500 ;
        RECT 4.830 35.700 5.680 36.550 ;
        RECT 23.780 35.700 24.630 36.550 ;
        RECT 24.830 35.700 25.680 36.550 ;
        RECT 43.780 35.700 44.630 36.550 ;
        RECT 44.830 35.700 45.680 36.550 ;
        RECT 63.780 35.700 64.630 36.550 ;
        RECT 64.830 35.700 65.680 36.550 ;
        RECT 83.780 35.700 84.630 36.550 ;
        RECT 84.830 35.700 85.680 36.550 ;
        RECT 103.780 35.700 104.630 36.550 ;
        RECT 105.340 36.805 105.700 37.185 ;
        RECT 105.970 36.805 106.330 37.185 ;
        RECT 106.570 36.805 106.930 37.185 ;
        RECT 105.340 36.215 105.700 36.595 ;
        RECT 105.970 36.215 106.330 36.595 ;
        RECT 106.570 36.215 106.930 36.595 ;
        RECT 2.520 34.925 2.880 35.305 ;
        RECT 3.130 34.925 3.490 35.305 ;
        RECT 3.760 34.925 4.120 35.305 ;
        RECT 2.520 34.190 2.880 34.570 ;
        RECT 3.130 34.190 3.490 34.570 ;
        RECT 3.760 34.190 4.120 34.570 ;
        RECT 2.520 33.505 2.880 33.885 ;
        RECT 3.130 33.505 3.490 33.885 ;
        RECT 3.760 33.505 4.120 33.885 ;
        RECT 2.520 26.120 2.880 26.500 ;
        RECT 3.130 26.120 3.490 26.500 ;
        RECT 3.760 26.120 4.120 26.500 ;
        RECT 2.520 25.385 2.880 25.765 ;
        RECT 3.130 25.385 3.490 25.765 ;
        RECT 3.760 25.385 4.120 25.765 ;
        RECT 2.520 24.700 2.880 25.080 ;
        RECT 3.130 24.700 3.490 25.080 ;
        RECT 3.760 24.700 4.120 25.080 ;
        RECT 2.515 23.145 2.875 23.525 ;
        RECT 3.145 23.145 3.505 23.525 ;
        RECT 3.745 23.145 4.105 23.525 ;
        RECT 2.515 22.555 2.875 22.935 ;
        RECT 3.145 22.555 3.505 22.935 ;
        RECT 3.745 22.555 4.105 22.935 ;
        RECT 4.830 23.450 5.680 24.300 ;
        RECT 23.780 23.450 24.630 24.300 ;
        RECT 24.830 23.450 25.680 24.300 ;
        RECT 43.780 23.450 44.630 24.300 ;
        RECT 44.830 23.450 45.680 24.300 ;
        RECT 63.780 23.450 64.630 24.300 ;
        RECT 64.830 23.450 65.680 24.300 ;
        RECT 83.780 23.450 84.630 24.300 ;
        RECT 84.830 23.450 85.680 24.300 ;
        RECT 103.780 23.450 104.630 24.300 ;
        RECT 4.830 22.500 5.680 23.350 ;
        RECT 23.780 22.500 24.630 23.350 ;
        RECT 24.830 22.500 25.680 23.350 ;
        RECT 43.780 22.500 44.630 23.350 ;
        RECT 44.830 22.500 45.680 23.350 ;
        RECT 63.780 22.500 64.630 23.350 ;
        RECT 64.830 22.500 65.680 23.350 ;
        RECT 83.780 22.500 84.630 23.350 ;
        RECT 84.830 22.500 85.680 23.350 ;
        RECT 103.780 22.500 104.630 23.350 ;
        RECT 4.830 21.050 5.680 21.900 ;
        RECT 4.830 20.100 5.680 20.950 ;
        RECT 5.780 20.100 6.630 20.950 ;
        RECT 7.230 20.100 8.080 20.950 ;
        RECT 8.180 20.100 9.030 20.950 ;
        RECT 4.830 19.050 5.680 19.900 ;
        RECT 5.780 19.050 6.630 19.900 ;
        RECT 7.230 19.050 8.080 19.900 ;
        RECT 8.180 19.050 9.030 19.900 ;
        RECT 4.830 18.100 5.680 18.950 ;
        RECT 23.780 21.050 24.630 21.900 ;
        RECT 24.830 21.050 25.680 21.900 ;
        RECT 20.430 20.100 21.280 20.950 ;
        RECT 21.380 20.100 22.230 20.950 ;
        RECT 22.830 20.100 23.680 20.950 ;
        RECT 23.780 20.100 24.630 20.950 ;
        RECT 24.830 20.100 25.680 20.950 ;
        RECT 25.780 20.100 26.630 20.950 ;
        RECT 27.230 20.100 28.080 20.950 ;
        RECT 28.180 20.100 29.030 20.950 ;
        RECT 20.430 19.050 21.280 19.900 ;
        RECT 21.380 19.050 22.230 19.900 ;
        RECT 22.830 19.050 23.680 19.900 ;
        RECT 23.780 19.050 24.630 19.900 ;
        RECT 24.830 19.050 25.680 19.900 ;
        RECT 25.780 19.050 26.630 19.900 ;
        RECT 27.230 19.050 28.080 19.900 ;
        RECT 28.180 19.050 29.030 19.900 ;
        RECT 23.780 18.100 24.630 18.950 ;
        RECT 24.830 18.100 25.680 18.950 ;
        RECT 43.780 21.050 44.630 21.900 ;
        RECT 44.830 21.050 45.680 21.900 ;
        RECT 40.430 20.100 41.280 20.950 ;
        RECT 41.380 20.100 42.230 20.950 ;
        RECT 42.830 20.100 43.680 20.950 ;
        RECT 43.780 20.100 44.630 20.950 ;
        RECT 44.830 20.100 45.680 20.950 ;
        RECT 45.780 20.100 46.630 20.950 ;
        RECT 47.230 20.100 48.080 20.950 ;
        RECT 48.180 20.100 49.030 20.950 ;
        RECT 40.430 19.050 41.280 19.900 ;
        RECT 41.380 19.050 42.230 19.900 ;
        RECT 42.830 19.050 43.680 19.900 ;
        RECT 43.780 19.050 44.630 19.900 ;
        RECT 44.830 19.050 45.680 19.900 ;
        RECT 45.780 19.050 46.630 19.900 ;
        RECT 47.230 19.050 48.080 19.900 ;
        RECT 48.180 19.050 49.030 19.900 ;
        RECT 43.780 18.100 44.630 18.950 ;
        RECT 44.830 18.100 45.680 18.950 ;
        RECT 63.780 21.050 64.630 21.900 ;
        RECT 64.830 21.050 65.680 21.900 ;
        RECT 60.430 20.100 61.280 20.950 ;
        RECT 61.380 20.100 62.230 20.950 ;
        RECT 62.830 20.100 63.680 20.950 ;
        RECT 63.780 20.100 64.630 20.950 ;
        RECT 64.830 20.100 65.680 20.950 ;
        RECT 65.780 20.100 66.630 20.950 ;
        RECT 67.230 20.100 68.080 20.950 ;
        RECT 68.180 20.100 69.030 20.950 ;
        RECT 60.430 19.050 61.280 19.900 ;
        RECT 61.380 19.050 62.230 19.900 ;
        RECT 62.830 19.050 63.680 19.900 ;
        RECT 63.780 19.050 64.630 19.900 ;
        RECT 64.830 19.050 65.680 19.900 ;
        RECT 65.780 19.050 66.630 19.900 ;
        RECT 67.230 19.050 68.080 19.900 ;
        RECT 68.180 19.050 69.030 19.900 ;
        RECT 63.780 18.100 64.630 18.950 ;
        RECT 64.830 18.100 65.680 18.950 ;
        RECT 83.780 21.050 84.630 21.900 ;
        RECT 84.830 21.050 85.680 21.900 ;
        RECT 80.430 20.100 81.280 20.950 ;
        RECT 81.380 20.100 82.230 20.950 ;
        RECT 82.830 20.100 83.680 20.950 ;
        RECT 83.780 20.100 84.630 20.950 ;
        RECT 84.830 20.100 85.680 20.950 ;
        RECT 85.780 20.100 86.630 20.950 ;
        RECT 87.230 20.100 88.080 20.950 ;
        RECT 88.180 20.100 89.030 20.950 ;
        RECT 80.430 19.050 81.280 19.900 ;
        RECT 81.380 19.050 82.230 19.900 ;
        RECT 82.830 19.050 83.680 19.900 ;
        RECT 83.780 19.050 84.630 19.900 ;
        RECT 84.830 19.050 85.680 19.900 ;
        RECT 85.780 19.050 86.630 19.900 ;
        RECT 87.230 19.050 88.080 19.900 ;
        RECT 88.180 19.050 89.030 19.900 ;
        RECT 83.780 18.100 84.630 18.950 ;
        RECT 84.830 18.100 85.680 18.950 ;
        RECT 103.780 21.050 104.630 21.900 ;
        RECT 105.340 22.590 105.700 22.970 ;
        RECT 105.970 22.590 106.330 22.970 ;
        RECT 106.570 22.590 106.930 22.970 ;
        RECT 105.340 22.000 105.700 22.380 ;
        RECT 105.970 22.000 106.330 22.380 ;
        RECT 106.570 22.000 106.930 22.380 ;
        RECT 100.430 20.100 101.280 20.950 ;
        RECT 101.380 20.100 102.230 20.950 ;
        RECT 102.830 20.100 103.680 20.950 ;
        RECT 103.780 20.100 104.630 20.950 ;
        RECT 100.430 19.050 101.280 19.900 ;
        RECT 101.380 19.050 102.230 19.900 ;
        RECT 102.830 19.050 103.680 19.900 ;
        RECT 103.780 19.050 104.630 19.900 ;
        RECT 103.780 18.100 104.630 18.950 ;
        RECT 2.515 17.260 2.875 17.640 ;
        RECT 3.145 17.260 3.505 17.640 ;
        RECT 3.745 17.260 4.105 17.640 ;
        RECT 2.515 16.670 2.875 17.050 ;
        RECT 3.145 16.670 3.505 17.050 ;
        RECT 3.745 16.670 4.105 17.050 ;
        RECT 4.830 16.650 5.680 17.500 ;
        RECT 23.780 16.650 24.630 17.500 ;
        RECT 24.830 16.650 25.680 17.500 ;
        RECT 43.780 16.650 44.630 17.500 ;
        RECT 44.830 16.650 45.680 17.500 ;
        RECT 63.780 16.650 64.630 17.500 ;
        RECT 64.830 16.650 65.680 17.500 ;
        RECT 83.780 16.650 84.630 17.500 ;
        RECT 84.830 16.650 85.680 17.500 ;
        RECT 103.780 16.650 104.630 17.500 ;
        RECT 4.830 15.700 5.680 16.550 ;
        RECT 23.780 15.700 24.630 16.550 ;
        RECT 24.830 15.700 25.680 16.550 ;
        RECT 43.780 15.700 44.630 16.550 ;
        RECT 44.830 15.700 45.680 16.550 ;
        RECT 63.780 15.700 64.630 16.550 ;
        RECT 64.830 15.700 65.680 16.550 ;
        RECT 83.780 15.700 84.630 16.550 ;
        RECT 84.830 15.700 85.680 16.550 ;
        RECT 103.780 15.700 104.630 16.550 ;
        RECT 105.340 16.805 105.700 17.185 ;
        RECT 105.970 16.805 106.330 17.185 ;
        RECT 106.570 16.805 106.930 17.185 ;
        RECT 105.340 16.215 105.700 16.595 ;
        RECT 105.970 16.215 106.330 16.595 ;
        RECT 106.570 16.215 106.930 16.595 ;
        RECT 2.520 14.925 2.880 15.305 ;
        RECT 3.130 14.925 3.490 15.305 ;
        RECT 3.760 14.925 4.120 15.305 ;
        RECT 2.520 14.190 2.880 14.570 ;
        RECT 3.130 14.190 3.490 14.570 ;
        RECT 3.760 14.190 4.120 14.570 ;
        RECT 2.520 13.505 2.880 13.885 ;
        RECT 3.130 13.505 3.490 13.885 ;
        RECT 3.760 13.505 4.120 13.885 ;
        RECT 2.520 6.120 2.880 6.500 ;
        RECT 3.130 6.120 3.490 6.500 ;
        RECT 3.760 6.120 4.120 6.500 ;
        RECT 2.520 5.385 2.880 5.765 ;
        RECT 3.130 5.385 3.490 5.765 ;
        RECT 3.760 5.385 4.120 5.765 ;
        RECT 2.520 4.700 2.880 5.080 ;
        RECT 3.130 4.700 3.490 5.080 ;
        RECT 3.760 4.700 4.120 5.080 ;
        RECT 2.515 3.145 2.875 3.525 ;
        RECT 3.145 3.145 3.505 3.525 ;
        RECT 3.745 3.145 4.105 3.525 ;
        RECT 2.515 2.555 2.875 2.935 ;
        RECT 3.145 2.555 3.505 2.935 ;
        RECT 3.745 2.555 4.105 2.935 ;
        RECT 4.830 3.450 5.680 4.300 ;
        RECT 23.780 3.450 24.630 4.300 ;
        RECT 24.830 3.450 25.680 4.300 ;
        RECT 43.780 3.450 44.630 4.300 ;
        RECT 44.830 3.450 45.680 4.300 ;
        RECT 63.780 3.450 64.630 4.300 ;
        RECT 64.830 3.450 65.680 4.300 ;
        RECT 83.780 3.450 84.630 4.300 ;
        RECT 84.830 3.450 85.680 4.300 ;
        RECT 103.780 3.450 104.630 4.300 ;
        RECT 4.830 2.500 5.680 3.350 ;
        RECT 23.780 2.500 24.630 3.350 ;
        RECT 24.830 2.500 25.680 3.350 ;
        RECT 43.780 2.500 44.630 3.350 ;
        RECT 44.830 2.500 45.680 3.350 ;
        RECT 63.780 2.500 64.630 3.350 ;
        RECT 64.830 2.500 65.680 3.350 ;
        RECT 83.780 2.500 84.630 3.350 ;
        RECT 84.830 2.500 85.680 3.350 ;
        RECT 103.780 2.500 104.630 3.350 ;
        RECT 4.830 1.050 5.680 1.900 ;
        RECT 4.830 0.100 5.680 0.950 ;
        RECT 5.780 0.100 6.630 0.950 ;
        RECT 7.230 0.100 8.080 0.950 ;
        RECT 8.180 0.100 9.030 0.950 ;
        RECT 23.780 1.050 24.630 1.900 ;
        RECT 24.830 1.050 25.680 1.900 ;
        RECT 20.430 0.100 21.280 0.950 ;
        RECT 21.380 0.100 22.230 0.950 ;
        RECT 22.830 0.100 23.680 0.950 ;
        RECT 23.780 0.100 24.630 0.950 ;
        RECT 24.830 0.100 25.680 0.950 ;
        RECT 25.780 0.100 26.630 0.950 ;
        RECT 27.230 0.100 28.080 0.950 ;
        RECT 28.180 0.100 29.030 0.950 ;
        RECT 43.780 1.050 44.630 1.900 ;
        RECT 44.830 1.050 45.680 1.900 ;
        RECT 40.430 0.100 41.280 0.950 ;
        RECT 41.380 0.100 42.230 0.950 ;
        RECT 42.830 0.100 43.680 0.950 ;
        RECT 43.780 0.100 44.630 0.950 ;
        RECT 44.830 0.100 45.680 0.950 ;
        RECT 45.780 0.100 46.630 0.950 ;
        RECT 47.230 0.100 48.080 0.950 ;
        RECT 48.180 0.100 49.030 0.950 ;
        RECT 63.780 1.050 64.630 1.900 ;
        RECT 64.830 1.050 65.680 1.900 ;
        RECT 60.430 0.100 61.280 0.950 ;
        RECT 61.380 0.100 62.230 0.950 ;
        RECT 62.830 0.100 63.680 0.950 ;
        RECT 63.780 0.100 64.630 0.950 ;
        RECT 64.830 0.100 65.680 0.950 ;
        RECT 65.780 0.100 66.630 0.950 ;
        RECT 67.230 0.100 68.080 0.950 ;
        RECT 68.180 0.100 69.030 0.950 ;
        RECT 83.780 1.050 84.630 1.900 ;
        RECT 84.830 1.050 85.680 1.900 ;
        RECT 80.430 0.100 81.280 0.950 ;
        RECT 81.380 0.100 82.230 0.950 ;
        RECT 82.830 0.100 83.680 0.950 ;
        RECT 83.780 0.100 84.630 0.950 ;
        RECT 84.830 0.100 85.680 0.950 ;
        RECT 85.780 0.100 86.630 0.950 ;
        RECT 87.230 0.100 88.080 0.950 ;
        RECT 88.180 0.100 89.030 0.950 ;
        RECT 103.780 1.050 104.630 1.900 ;
        RECT 105.340 2.590 105.700 2.970 ;
        RECT 105.970 2.590 106.330 2.970 ;
        RECT 106.570 2.590 106.930 2.970 ;
        RECT 105.340 2.000 105.700 2.380 ;
        RECT 105.970 2.000 106.330 2.380 ;
        RECT 106.570 2.000 106.930 2.380 ;
        RECT 100.430 0.100 101.280 0.950 ;
        RECT 101.380 0.100 102.230 0.950 ;
        RECT 102.830 0.100 103.680 0.950 ;
        RECT 103.780 0.100 104.630 0.950 ;
      LAYER met4 ;
        RECT 2.315 377.385 4.315 380.000 ;
        RECT 105.140 377.585 107.140 380.000 ;
        RECT 2.315 376.110 4.320 377.385 ;
        RECT 105.130 376.310 107.140 377.585 ;
        RECT 2.315 364.020 4.315 376.110 ;
        RECT 2.315 362.745 4.320 364.020 ;
        RECT 2.315 357.385 4.315 362.745 ;
        RECT 105.140 357.585 107.140 376.310 ;
        RECT 2.315 356.110 4.320 357.385 ;
        RECT 105.130 356.310 107.140 357.585 ;
        RECT 2.315 344.020 4.315 356.110 ;
        RECT 2.315 342.745 4.320 344.020 ;
        RECT 2.315 337.375 4.315 342.745 ;
        RECT 105.140 337.585 107.140 356.310 ;
        RECT 2.315 336.100 4.320 337.375 ;
        RECT 105.130 336.310 107.140 337.585 ;
        RECT 2.315 323.675 4.315 336.100 ;
        RECT 2.315 322.400 4.320 323.675 ;
        RECT 2.315 317.785 4.315 322.400 ;
        RECT 2.315 316.510 4.320 317.785 ;
        RECT 105.140 317.585 107.140 336.310 ;
        RECT 2.315 315.545 4.315 316.510 ;
        RECT 105.130 316.310 107.140 317.585 ;
        RECT 2.315 313.250 4.320 315.545 ;
        RECT 2.315 303.545 4.315 313.250 ;
        RECT 2.315 302.270 4.330 303.545 ;
        RECT 2.315 297.530 4.315 302.270 ;
        RECT 105.140 297.855 107.140 316.310 ;
        RECT 2.315 296.255 4.320 297.530 ;
        RECT 105.135 296.580 107.140 297.855 ;
        RECT 2.315 295.545 4.315 296.255 ;
        RECT 2.315 293.250 4.320 295.545 ;
        RECT 2.315 283.645 4.315 293.250 ;
        RECT 2.315 282.370 4.320 283.645 ;
        RECT 2.315 277.610 4.315 282.370 ;
        RECT 2.315 276.335 4.330 277.610 ;
        RECT 105.140 277.360 107.140 296.580 ;
        RECT 2.315 263.780 4.315 276.335 ;
        RECT 105.135 276.085 107.140 277.360 ;
        RECT 2.315 262.505 4.320 263.780 ;
        RECT 2.315 257.845 4.315 262.505 ;
        RECT 2.315 256.570 4.320 257.845 ;
        RECT 2.315 243.735 4.315 256.570 ;
        RECT 2.315 242.460 4.320 243.735 ;
        RECT 2.315 237.970 4.315 242.460 ;
        RECT 2.315 236.695 4.320 237.970 ;
        RECT 2.315 161.800 4.315 236.695 ;
        RECT 42.635 181.610 47.035 182.660 ;
        RECT 58.235 181.610 67.035 182.660 ;
        RECT 78.235 181.610 87.035 182.660 ;
        RECT 98.235 181.610 102.635 182.660 ;
        RECT 42.635 178.260 43.685 181.610 ;
        RECT 61.585 178.260 63.685 181.610 ;
        RECT 81.585 178.260 83.685 181.610 ;
        RECT 101.585 180.990 102.635 181.610 ;
        RECT 105.140 180.990 107.140 276.085 ;
        RECT 101.585 179.715 107.140 180.990 ;
        RECT 101.585 178.260 102.635 179.715 ;
        RECT 42.635 163.710 43.685 167.060 ;
        RECT 61.585 163.710 63.685 167.060 ;
        RECT 81.585 163.710 83.685 167.060 ;
        RECT 101.585 165.715 102.635 167.060 ;
        RECT 105.140 165.715 107.140 179.715 ;
        RECT 101.585 164.440 107.140 165.715 ;
        RECT 101.585 163.710 102.635 164.440 ;
        RECT 42.635 162.660 47.035 163.710 ;
        RECT 58.235 162.660 67.035 163.710 ;
        RECT 78.235 162.660 87.035 163.710 ;
        RECT 98.235 162.660 102.635 163.710 ;
        RECT 105.140 161.800 107.140 164.440 ;
        RECT 2.315 160.360 4.330 161.800 ;
        RECT 105.125 160.360 107.140 161.800 ;
        RECT 2.315 160.000 4.315 160.360 ;
        RECT 2.315 158.950 9.130 160.000 ;
        RECT 20.330 158.950 29.130 160.000 ;
        RECT 40.330 158.950 49.130 160.000 ;
        RECT 60.330 158.950 69.130 160.000 ;
        RECT 80.330 158.950 89.130 160.000 ;
        RECT 100.330 158.950 104.730 160.000 ;
        RECT 2.315 158.800 5.780 158.950 ;
        RECT 2.315 141.190 4.315 158.800 ;
        RECT 4.730 155.600 5.780 158.800 ;
        RECT 23.680 155.600 25.780 158.950 ;
        RECT 43.680 155.600 45.780 158.950 ;
        RECT 63.680 155.600 65.780 158.950 ;
        RECT 83.680 155.600 85.780 158.950 ;
        RECT 103.680 155.600 104.730 158.950 ;
        RECT 4.730 141.190 5.780 144.400 ;
        RECT 2.315 141.050 5.780 141.190 ;
        RECT 23.680 141.050 25.780 144.400 ;
        RECT 43.680 141.050 45.780 144.400 ;
        RECT 63.680 141.050 65.780 144.400 ;
        RECT 83.680 141.050 85.780 144.400 ;
        RECT 103.680 141.160 104.730 144.400 ;
        RECT 105.140 141.160 107.140 160.360 ;
        RECT 103.680 141.050 107.140 141.160 ;
        RECT 2.315 141.045 9.130 141.050 ;
        RECT 2.310 139.895 9.130 141.045 ;
        RECT 2.315 138.950 9.130 139.895 ;
        RECT 20.330 138.950 29.130 141.050 ;
        RECT 40.330 138.950 49.130 141.050 ;
        RECT 60.330 138.950 69.130 141.050 ;
        RECT 80.330 138.950 89.130 141.050 ;
        RECT 100.330 138.950 107.140 141.050 ;
        RECT 2.315 138.800 5.780 138.950 ;
        RECT 2.315 123.255 4.315 138.800 ;
        RECT 4.730 135.600 5.780 138.800 ;
        RECT 23.680 135.600 25.780 138.950 ;
        RECT 43.680 135.600 45.780 138.950 ;
        RECT 63.680 135.600 65.780 138.950 ;
        RECT 83.680 135.600 85.780 138.950 ;
        RECT 103.680 138.830 107.140 138.950 ;
        RECT 103.680 135.600 104.730 138.830 ;
        RECT 105.140 137.335 107.140 138.830 ;
        RECT 105.135 136.060 107.140 137.335 ;
        RECT 2.315 121.980 4.320 123.255 ;
        RECT 2.315 121.195 4.315 121.980 ;
        RECT 4.730 121.195 5.780 124.400 ;
        RECT 2.315 121.050 5.780 121.195 ;
        RECT 23.680 121.050 25.780 124.400 ;
        RECT 43.680 121.050 45.780 124.400 ;
        RECT 63.680 121.050 65.780 124.400 ;
        RECT 83.680 121.050 85.780 124.400 ;
        RECT 103.680 121.160 104.730 124.400 ;
        RECT 105.140 121.160 107.140 136.060 ;
        RECT 103.680 121.050 107.140 121.160 ;
        RECT 2.315 118.950 9.130 121.050 ;
        RECT 20.330 118.950 29.130 121.050 ;
        RECT 40.330 118.950 49.130 121.050 ;
        RECT 60.330 118.950 69.130 121.050 ;
        RECT 80.330 118.950 89.130 121.050 ;
        RECT 100.330 118.950 107.140 121.050 ;
        RECT 2.315 118.795 5.780 118.950 ;
        RECT 2.315 117.845 4.315 118.795 ;
        RECT 2.315 116.570 4.320 117.845 ;
        RECT 2.315 103.470 4.315 116.570 ;
        RECT 4.730 115.600 5.780 118.795 ;
        RECT 23.680 115.600 25.780 118.950 ;
        RECT 43.680 115.600 45.780 118.950 ;
        RECT 63.680 115.600 65.780 118.950 ;
        RECT 83.680 115.600 85.780 118.950 ;
        RECT 103.680 118.835 107.140 118.950 ;
        RECT 103.680 115.600 104.730 118.835 ;
        RECT 2.315 102.195 4.320 103.470 ;
        RECT 2.315 101.200 4.315 102.195 ;
        RECT 4.730 101.200 5.780 104.400 ;
        RECT 2.315 101.050 5.780 101.200 ;
        RECT 23.680 101.050 25.780 104.400 ;
        RECT 43.680 101.050 45.780 104.400 ;
        RECT 63.680 101.050 65.780 104.400 ;
        RECT 83.680 101.050 85.780 104.400 ;
        RECT 103.680 101.165 104.730 104.400 ;
        RECT 105.140 103.040 107.140 118.835 ;
        RECT 105.135 101.765 107.140 103.040 ;
        RECT 105.140 101.165 107.140 101.765 ;
        RECT 103.680 101.050 107.140 101.165 ;
        RECT 2.315 98.950 9.130 101.050 ;
        RECT 20.330 98.950 29.130 101.050 ;
        RECT 40.330 98.950 49.130 101.050 ;
        RECT 60.330 98.950 69.130 101.050 ;
        RECT 80.330 98.950 89.130 101.050 ;
        RECT 100.330 98.950 107.140 101.050 ;
        RECT 2.315 98.800 5.780 98.950 ;
        RECT 2.315 97.965 4.315 98.800 ;
        RECT 2.315 96.690 4.320 97.965 ;
        RECT 2.315 83.635 4.315 96.690 ;
        RECT 4.730 95.600 5.780 98.800 ;
        RECT 23.680 95.600 25.780 98.950 ;
        RECT 43.680 95.600 45.780 98.950 ;
        RECT 63.680 95.600 65.780 98.950 ;
        RECT 83.680 95.600 85.780 98.950 ;
        RECT 103.680 98.840 107.140 98.950 ;
        RECT 103.680 95.600 104.730 98.840 ;
        RECT 105.140 97.185 107.140 98.840 ;
        RECT 105.135 95.910 107.140 97.185 ;
        RECT 2.315 82.360 4.325 83.635 ;
        RECT 2.315 81.195 4.315 82.360 ;
        RECT 4.730 81.195 5.780 84.400 ;
        RECT 2.315 81.050 5.780 81.195 ;
        RECT 23.680 81.050 25.780 84.400 ;
        RECT 43.680 81.050 45.780 84.400 ;
        RECT 63.680 81.050 65.780 84.400 ;
        RECT 83.680 81.050 85.780 84.400 ;
        RECT 103.680 81.160 104.730 84.400 ;
        RECT 105.140 83.380 107.140 95.910 ;
        RECT 105.135 82.105 107.140 83.380 ;
        RECT 105.140 81.160 107.140 82.105 ;
        RECT 103.680 81.050 107.140 81.160 ;
        RECT 2.315 78.950 9.130 81.050 ;
        RECT 20.330 78.950 29.130 81.050 ;
        RECT 40.330 78.950 49.130 81.050 ;
        RECT 60.330 78.950 69.130 81.050 ;
        RECT 80.330 78.950 89.130 81.050 ;
        RECT 100.330 78.950 107.140 81.050 ;
        RECT 2.315 78.795 5.780 78.950 ;
        RECT 2.315 77.555 4.315 78.795 ;
        RECT 2.315 76.280 4.330 77.555 ;
        RECT 2.315 63.230 4.315 76.280 ;
        RECT 4.730 75.600 5.780 78.795 ;
        RECT 23.680 75.600 25.780 78.950 ;
        RECT 43.680 75.600 45.780 78.950 ;
        RECT 63.680 75.600 65.780 78.950 ;
        RECT 83.680 75.600 85.780 78.950 ;
        RECT 103.680 78.830 107.140 78.950 ;
        RECT 103.680 75.600 104.730 78.830 ;
        RECT 105.140 77.310 107.140 78.830 ;
        RECT 105.135 76.035 107.140 77.310 ;
        RECT 2.315 61.955 4.320 63.230 ;
        RECT 2.315 61.190 4.315 61.955 ;
        RECT 4.730 61.190 5.780 64.400 ;
        RECT 2.315 61.050 5.780 61.190 ;
        RECT 23.680 61.050 25.780 64.400 ;
        RECT 43.680 61.050 45.780 64.400 ;
        RECT 63.680 61.050 65.780 64.400 ;
        RECT 83.680 61.050 85.780 64.400 ;
        RECT 103.680 61.165 104.730 64.400 ;
        RECT 105.140 61.165 107.140 76.035 ;
        RECT 103.680 61.050 107.140 61.165 ;
        RECT 2.315 58.950 9.130 61.050 ;
        RECT 20.330 58.950 29.130 61.050 ;
        RECT 40.330 58.950 49.130 61.050 ;
        RECT 60.330 58.950 69.130 61.050 ;
        RECT 80.330 58.950 89.130 61.050 ;
        RECT 100.330 58.950 107.140 61.050 ;
        RECT 2.315 58.790 5.780 58.950 ;
        RECT 2.315 57.620 4.315 58.790 ;
        RECT 2.315 56.345 4.320 57.620 ;
        RECT 2.315 41.190 4.315 56.345 ;
        RECT 4.730 55.600 5.780 58.790 ;
        RECT 23.680 55.600 25.780 58.950 ;
        RECT 43.680 55.600 45.780 58.950 ;
        RECT 63.680 55.600 65.780 58.950 ;
        RECT 83.680 55.600 85.780 58.950 ;
        RECT 103.680 58.830 107.140 58.950 ;
        RECT 103.680 55.600 104.730 58.830 ;
        RECT 105.140 57.310 107.140 58.830 ;
        RECT 105.135 56.035 107.140 57.310 ;
        RECT 4.730 41.190 5.780 44.400 ;
        RECT 2.315 41.050 5.780 41.190 ;
        RECT 23.680 41.050 25.780 44.400 ;
        RECT 43.680 41.050 45.780 44.400 ;
        RECT 63.680 41.050 65.780 44.400 ;
        RECT 83.680 41.050 85.780 44.400 ;
        RECT 103.680 41.165 104.730 44.400 ;
        RECT 105.140 41.165 107.140 56.035 ;
        RECT 103.680 41.050 107.140 41.165 ;
        RECT 2.315 38.950 9.130 41.050 ;
        RECT 20.330 38.950 29.130 41.050 ;
        RECT 40.330 38.950 49.130 41.050 ;
        RECT 60.330 38.950 69.130 41.050 ;
        RECT 80.330 38.950 89.130 41.050 ;
        RECT 100.330 38.950 107.140 41.050 ;
        RECT 2.315 38.800 5.780 38.950 ;
        RECT 2.315 23.650 4.315 38.800 ;
        RECT 4.730 35.600 5.780 38.800 ;
        RECT 23.680 35.600 25.780 38.950 ;
        RECT 43.680 35.600 45.780 38.950 ;
        RECT 63.680 35.600 65.780 38.950 ;
        RECT 83.680 35.600 85.780 38.950 ;
        RECT 103.680 38.830 107.140 38.950 ;
        RECT 103.680 35.600 104.730 38.830 ;
        RECT 105.140 37.310 107.140 38.830 ;
        RECT 105.135 36.035 107.140 37.310 ;
        RECT 2.315 22.375 4.325 23.650 ;
        RECT 2.315 21.195 4.315 22.375 ;
        RECT 4.730 21.195 5.780 24.400 ;
        RECT 2.315 21.050 5.780 21.195 ;
        RECT 23.680 21.050 25.780 24.400 ;
        RECT 43.680 21.050 45.780 24.400 ;
        RECT 63.680 21.050 65.780 24.400 ;
        RECT 83.680 21.050 85.780 24.400 ;
        RECT 103.680 21.165 104.730 24.400 ;
        RECT 105.140 21.165 107.140 36.035 ;
        RECT 103.680 21.050 107.140 21.165 ;
        RECT 2.315 18.950 9.130 21.050 ;
        RECT 20.330 18.950 29.130 21.050 ;
        RECT 40.330 18.950 49.130 21.050 ;
        RECT 60.330 18.950 69.130 21.050 ;
        RECT 80.330 18.950 89.130 21.050 ;
        RECT 100.330 18.950 107.140 21.050 ;
        RECT 2.315 18.800 5.780 18.950 ;
        RECT 2.315 3.650 4.315 18.800 ;
        RECT 4.730 15.600 5.780 18.800 ;
        RECT 23.680 15.600 25.780 18.950 ;
        RECT 43.680 15.600 45.780 18.950 ;
        RECT 63.680 15.600 65.780 18.950 ;
        RECT 83.680 15.600 85.780 18.950 ;
        RECT 103.680 18.830 107.140 18.950 ;
        RECT 103.680 15.600 104.730 18.830 ;
        RECT 105.140 17.310 107.140 18.830 ;
        RECT 105.135 16.035 107.140 17.310 ;
        RECT 2.315 2.375 4.325 3.650 ;
        RECT 2.315 1.195 4.315 2.375 ;
        RECT 4.730 1.195 5.780 4.400 ;
        RECT 2.315 1.050 5.780 1.195 ;
        RECT 23.680 1.050 25.780 4.400 ;
        RECT 43.680 1.050 45.780 4.400 ;
        RECT 63.680 1.050 65.780 4.400 ;
        RECT 83.680 1.050 85.780 4.400 ;
        RECT 103.680 1.165 104.730 4.400 ;
        RECT 105.140 1.165 107.140 16.035 ;
        RECT 103.680 1.050 107.140 1.165 ;
        RECT 2.315 0.000 9.130 1.050 ;
        RECT 20.330 0.000 29.130 1.050 ;
        RECT 40.330 0.000 49.130 1.050 ;
        RECT 60.330 0.000 69.130 1.050 ;
        RECT 80.330 0.000 89.130 1.050 ;
        RECT 100.330 0.000 107.140 1.050 ;
    END
  END VSS
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 6.695 191.085 7.615 191.345 ;
        RECT 8.530 191.090 8.865 191.340 ;
        RECT 7.365 188.700 7.695 188.940 ;
      LAYER mcon ;
        RECT 7.395 191.125 7.575 191.300 ;
        RECT 8.575 191.120 8.745 191.290 ;
        RECT 7.405 188.740 7.575 188.910 ;
      LAYER met1 ;
        RECT 7.325 191.340 7.645 191.345 ;
        RECT 7.325 191.090 8.865 191.340 ;
        RECT 7.325 191.085 7.645 191.090 ;
        RECT 7.285 188.690 7.695 188.950 ;
      LAYER via ;
        RECT 7.355 191.085 7.615 191.345 ;
        RECT 7.315 188.690 7.575 188.950 ;
      LAYER met2 ;
        RECT 7.355 191.055 7.615 191.375 ;
        RECT 7.355 188.985 7.520 191.055 ;
        RECT 7.315 188.660 7.575 188.985 ;
    END
  END clk
  PIN vcm
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 20992.000000 ;
    ANTENNADIFFAREA 1.160000 ;
    PORT
      LAYER li1 ;
        RECT 5.930 377.600 9.930 377.800 ;
        RECT 5.930 377.000 6.330 377.600 ;
        RECT 5.930 376.800 9.930 377.000 ;
        RECT 5.930 376.200 6.330 376.800 ;
        RECT 5.930 376.000 9.930 376.200 ;
        RECT 5.930 375.400 6.330 376.000 ;
        RECT 5.930 375.200 9.930 375.400 ;
        RECT 5.930 374.600 6.330 375.200 ;
        RECT 5.930 374.400 9.930 374.600 ;
        RECT 5.930 373.800 6.330 374.400 ;
        RECT 5.930 373.600 9.930 373.800 ;
        RECT 5.930 373.000 6.330 373.600 ;
        RECT 5.930 372.800 9.930 373.000 ;
        RECT 5.930 372.200 6.330 372.800 ;
        RECT 5.930 372.000 9.930 372.200 ;
        RECT 5.930 371.400 6.330 372.000 ;
        RECT 5.930 371.200 9.930 371.400 ;
        RECT 5.930 370.600 6.330 371.200 ;
        RECT 5.930 370.400 9.930 370.600 ;
        RECT 5.930 370.200 6.330 370.400 ;
        RECT 10.680 370.200 10.880 377.800 ;
        RECT 11.480 370.200 11.680 377.800 ;
        RECT 12.280 370.200 12.480 377.800 ;
        RECT 13.080 370.200 13.280 377.800 ;
        RECT 13.880 370.200 14.080 377.800 ;
        RECT 5.930 369.800 14.080 370.200 ;
        RECT 5.930 369.600 6.330 369.800 ;
        RECT 5.930 369.400 9.930 369.600 ;
        RECT 5.930 368.800 6.330 369.400 ;
        RECT 5.930 368.600 9.930 368.800 ;
        RECT 5.930 368.000 6.330 368.600 ;
        RECT 5.930 367.800 9.930 368.000 ;
        RECT 5.930 367.200 6.330 367.800 ;
        RECT 5.930 367.000 9.930 367.200 ;
        RECT 5.930 366.400 6.330 367.000 ;
        RECT 5.930 366.200 9.930 366.400 ;
        RECT 5.930 365.600 6.330 366.200 ;
        RECT 5.930 365.400 9.930 365.600 ;
        RECT 5.930 364.800 6.330 365.400 ;
        RECT 5.930 364.600 9.930 364.800 ;
        RECT 5.930 364.000 6.330 364.600 ;
        RECT 5.930 363.800 9.930 364.000 ;
        RECT 5.930 363.200 6.330 363.800 ;
        RECT 5.930 363.000 9.930 363.200 ;
        RECT 5.930 362.400 6.330 363.000 ;
        RECT 5.930 362.200 9.930 362.400 ;
        RECT 10.680 362.200 10.880 369.800 ;
        RECT 11.480 362.200 11.680 369.800 ;
        RECT 12.280 362.200 12.480 369.800 ;
        RECT 13.080 362.200 13.280 369.800 ;
        RECT 13.880 362.200 14.080 369.800 ;
        RECT 15.380 370.200 15.580 377.800 ;
        RECT 16.180 370.200 16.380 377.800 ;
        RECT 16.980 370.200 17.180 377.800 ;
        RECT 17.780 370.200 17.980 377.800 ;
        RECT 18.580 370.200 18.780 377.800 ;
        RECT 19.530 377.600 23.530 377.800 ;
        RECT 23.130 377.000 23.530 377.600 ;
        RECT 19.530 376.800 23.530 377.000 ;
        RECT 23.130 376.200 23.530 376.800 ;
        RECT 19.530 376.000 23.530 376.200 ;
        RECT 23.130 375.400 23.530 376.000 ;
        RECT 19.530 375.200 23.530 375.400 ;
        RECT 23.130 374.600 23.530 375.200 ;
        RECT 19.530 374.400 23.530 374.600 ;
        RECT 23.130 373.800 23.530 374.400 ;
        RECT 19.530 373.600 23.530 373.800 ;
        RECT 23.130 373.000 23.530 373.600 ;
        RECT 19.530 372.800 23.530 373.000 ;
        RECT 23.130 372.200 23.530 372.800 ;
        RECT 19.530 372.000 23.530 372.200 ;
        RECT 23.130 371.400 23.530 372.000 ;
        RECT 19.530 371.200 23.530 371.400 ;
        RECT 23.130 370.600 23.530 371.200 ;
        RECT 19.530 370.400 23.530 370.600 ;
        RECT 23.130 370.200 23.530 370.400 ;
        RECT 15.380 369.800 23.530 370.200 ;
        RECT 15.380 362.200 15.580 369.800 ;
        RECT 16.180 362.200 16.380 369.800 ;
        RECT 16.980 362.200 17.180 369.800 ;
        RECT 17.780 362.200 17.980 369.800 ;
        RECT 18.580 362.200 18.780 369.800 ;
        RECT 23.130 369.600 23.530 369.800 ;
        RECT 19.530 369.400 23.530 369.600 ;
        RECT 23.130 368.800 23.530 369.400 ;
        RECT 19.530 368.600 23.530 368.800 ;
        RECT 23.130 368.000 23.530 368.600 ;
        RECT 19.530 367.800 23.530 368.000 ;
        RECT 23.130 367.200 23.530 367.800 ;
        RECT 19.530 367.000 23.530 367.200 ;
        RECT 23.130 366.400 23.530 367.000 ;
        RECT 19.530 366.200 23.530 366.400 ;
        RECT 23.130 365.600 23.530 366.200 ;
        RECT 19.530 365.400 23.530 365.600 ;
        RECT 23.130 364.800 23.530 365.400 ;
        RECT 19.530 364.600 23.530 364.800 ;
        RECT 23.130 364.000 23.530 364.600 ;
        RECT 19.530 363.800 23.530 364.000 ;
        RECT 23.130 363.200 23.530 363.800 ;
        RECT 19.530 363.000 23.530 363.200 ;
        RECT 23.130 362.400 23.530 363.000 ;
        RECT 19.530 362.200 23.530 362.400 ;
        RECT 25.930 377.600 29.930 377.800 ;
        RECT 25.930 377.000 26.330 377.600 ;
        RECT 25.930 376.800 29.930 377.000 ;
        RECT 25.930 376.200 26.330 376.800 ;
        RECT 25.930 376.000 29.930 376.200 ;
        RECT 25.930 375.400 26.330 376.000 ;
        RECT 25.930 375.200 29.930 375.400 ;
        RECT 25.930 374.600 26.330 375.200 ;
        RECT 25.930 374.400 29.930 374.600 ;
        RECT 25.930 373.800 26.330 374.400 ;
        RECT 25.930 373.600 29.930 373.800 ;
        RECT 25.930 373.000 26.330 373.600 ;
        RECT 25.930 372.800 29.930 373.000 ;
        RECT 25.930 372.200 26.330 372.800 ;
        RECT 25.930 372.000 29.930 372.200 ;
        RECT 25.930 371.400 26.330 372.000 ;
        RECT 25.930 371.200 29.930 371.400 ;
        RECT 25.930 370.600 26.330 371.200 ;
        RECT 25.930 370.400 29.930 370.600 ;
        RECT 25.930 370.200 26.330 370.400 ;
        RECT 30.680 370.200 30.880 377.800 ;
        RECT 31.480 370.200 31.680 377.800 ;
        RECT 32.280 370.200 32.480 377.800 ;
        RECT 33.080 370.200 33.280 377.800 ;
        RECT 33.880 370.200 34.080 377.800 ;
        RECT 25.930 369.800 34.080 370.200 ;
        RECT 25.930 369.600 26.330 369.800 ;
        RECT 25.930 369.400 29.930 369.600 ;
        RECT 25.930 368.800 26.330 369.400 ;
        RECT 25.930 368.600 29.930 368.800 ;
        RECT 25.930 368.000 26.330 368.600 ;
        RECT 25.930 367.800 29.930 368.000 ;
        RECT 25.930 367.200 26.330 367.800 ;
        RECT 25.930 367.000 29.930 367.200 ;
        RECT 25.930 366.400 26.330 367.000 ;
        RECT 25.930 366.200 29.930 366.400 ;
        RECT 25.930 365.600 26.330 366.200 ;
        RECT 25.930 365.400 29.930 365.600 ;
        RECT 25.930 364.800 26.330 365.400 ;
        RECT 25.930 364.600 29.930 364.800 ;
        RECT 25.930 364.000 26.330 364.600 ;
        RECT 25.930 363.800 29.930 364.000 ;
        RECT 25.930 363.200 26.330 363.800 ;
        RECT 25.930 363.000 29.930 363.200 ;
        RECT 25.930 362.400 26.330 363.000 ;
        RECT 25.930 362.200 29.930 362.400 ;
        RECT 30.680 362.200 30.880 369.800 ;
        RECT 31.480 362.200 31.680 369.800 ;
        RECT 32.280 362.200 32.480 369.800 ;
        RECT 33.080 362.200 33.280 369.800 ;
        RECT 33.880 362.200 34.080 369.800 ;
        RECT 35.380 370.200 35.580 377.800 ;
        RECT 36.180 370.200 36.380 377.800 ;
        RECT 36.980 370.200 37.180 377.800 ;
        RECT 37.780 370.200 37.980 377.800 ;
        RECT 38.580 370.200 38.780 377.800 ;
        RECT 39.530 377.600 43.530 377.800 ;
        RECT 43.130 377.000 43.530 377.600 ;
        RECT 39.530 376.800 43.530 377.000 ;
        RECT 43.130 376.200 43.530 376.800 ;
        RECT 39.530 376.000 43.530 376.200 ;
        RECT 43.130 375.400 43.530 376.000 ;
        RECT 39.530 375.200 43.530 375.400 ;
        RECT 43.130 374.600 43.530 375.200 ;
        RECT 39.530 374.400 43.530 374.600 ;
        RECT 43.130 373.800 43.530 374.400 ;
        RECT 39.530 373.600 43.530 373.800 ;
        RECT 43.130 373.000 43.530 373.600 ;
        RECT 39.530 372.800 43.530 373.000 ;
        RECT 43.130 372.200 43.530 372.800 ;
        RECT 39.530 372.000 43.530 372.200 ;
        RECT 43.130 371.400 43.530 372.000 ;
        RECT 39.530 371.200 43.530 371.400 ;
        RECT 43.130 370.600 43.530 371.200 ;
        RECT 39.530 370.400 43.530 370.600 ;
        RECT 43.130 370.200 43.530 370.400 ;
        RECT 35.380 369.800 43.530 370.200 ;
        RECT 35.380 362.200 35.580 369.800 ;
        RECT 36.180 362.200 36.380 369.800 ;
        RECT 36.980 362.200 37.180 369.800 ;
        RECT 37.780 362.200 37.980 369.800 ;
        RECT 38.580 362.200 38.780 369.800 ;
        RECT 43.130 369.600 43.530 369.800 ;
        RECT 39.530 369.400 43.530 369.600 ;
        RECT 43.130 368.800 43.530 369.400 ;
        RECT 39.530 368.600 43.530 368.800 ;
        RECT 43.130 368.000 43.530 368.600 ;
        RECT 39.530 367.800 43.530 368.000 ;
        RECT 43.130 367.200 43.530 367.800 ;
        RECT 39.530 367.000 43.530 367.200 ;
        RECT 43.130 366.400 43.530 367.000 ;
        RECT 39.530 366.200 43.530 366.400 ;
        RECT 43.130 365.600 43.530 366.200 ;
        RECT 39.530 365.400 43.530 365.600 ;
        RECT 43.130 364.800 43.530 365.400 ;
        RECT 39.530 364.600 43.530 364.800 ;
        RECT 43.130 364.000 43.530 364.600 ;
        RECT 39.530 363.800 43.530 364.000 ;
        RECT 43.130 363.200 43.530 363.800 ;
        RECT 39.530 363.000 43.530 363.200 ;
        RECT 43.130 362.400 43.530 363.000 ;
        RECT 39.530 362.200 43.530 362.400 ;
        RECT 45.930 377.600 49.930 377.800 ;
        RECT 45.930 377.000 46.330 377.600 ;
        RECT 45.930 376.800 49.930 377.000 ;
        RECT 45.930 376.200 46.330 376.800 ;
        RECT 45.930 376.000 49.930 376.200 ;
        RECT 45.930 375.400 46.330 376.000 ;
        RECT 45.930 375.200 49.930 375.400 ;
        RECT 45.930 374.600 46.330 375.200 ;
        RECT 45.930 374.400 49.930 374.600 ;
        RECT 45.930 373.800 46.330 374.400 ;
        RECT 45.930 373.600 49.930 373.800 ;
        RECT 45.930 373.000 46.330 373.600 ;
        RECT 45.930 372.800 49.930 373.000 ;
        RECT 45.930 372.200 46.330 372.800 ;
        RECT 45.930 372.000 49.930 372.200 ;
        RECT 45.930 371.400 46.330 372.000 ;
        RECT 45.930 371.200 49.930 371.400 ;
        RECT 45.930 370.600 46.330 371.200 ;
        RECT 45.930 370.400 49.930 370.600 ;
        RECT 45.930 370.200 46.330 370.400 ;
        RECT 50.680 370.200 50.880 377.800 ;
        RECT 51.480 370.200 51.680 377.800 ;
        RECT 52.280 370.200 52.480 377.800 ;
        RECT 53.080 370.200 53.280 377.800 ;
        RECT 53.880 370.200 54.080 377.800 ;
        RECT 45.930 369.800 54.080 370.200 ;
        RECT 45.930 369.600 46.330 369.800 ;
        RECT 45.930 369.400 49.930 369.600 ;
        RECT 45.930 368.800 46.330 369.400 ;
        RECT 45.930 368.600 49.930 368.800 ;
        RECT 45.930 368.000 46.330 368.600 ;
        RECT 45.930 367.800 49.930 368.000 ;
        RECT 45.930 367.200 46.330 367.800 ;
        RECT 45.930 367.000 49.930 367.200 ;
        RECT 45.930 366.400 46.330 367.000 ;
        RECT 45.930 366.200 49.930 366.400 ;
        RECT 45.930 365.600 46.330 366.200 ;
        RECT 45.930 365.400 49.930 365.600 ;
        RECT 45.930 364.800 46.330 365.400 ;
        RECT 45.930 364.600 49.930 364.800 ;
        RECT 45.930 364.000 46.330 364.600 ;
        RECT 45.930 363.800 49.930 364.000 ;
        RECT 45.930 363.200 46.330 363.800 ;
        RECT 45.930 363.000 49.930 363.200 ;
        RECT 45.930 362.400 46.330 363.000 ;
        RECT 45.930 362.200 49.930 362.400 ;
        RECT 50.680 362.200 50.880 369.800 ;
        RECT 51.480 362.200 51.680 369.800 ;
        RECT 52.280 362.200 52.480 369.800 ;
        RECT 53.080 362.200 53.280 369.800 ;
        RECT 53.880 362.200 54.080 369.800 ;
        RECT 55.380 370.200 55.580 377.800 ;
        RECT 56.180 370.200 56.380 377.800 ;
        RECT 56.980 370.200 57.180 377.800 ;
        RECT 57.780 370.200 57.980 377.800 ;
        RECT 58.580 370.200 58.780 377.800 ;
        RECT 59.530 377.600 63.530 377.800 ;
        RECT 63.130 377.000 63.530 377.600 ;
        RECT 59.530 376.800 63.530 377.000 ;
        RECT 63.130 376.200 63.530 376.800 ;
        RECT 59.530 376.000 63.530 376.200 ;
        RECT 63.130 375.400 63.530 376.000 ;
        RECT 59.530 375.200 63.530 375.400 ;
        RECT 63.130 374.600 63.530 375.200 ;
        RECT 59.530 374.400 63.530 374.600 ;
        RECT 63.130 373.800 63.530 374.400 ;
        RECT 59.530 373.600 63.530 373.800 ;
        RECT 63.130 373.000 63.530 373.600 ;
        RECT 59.530 372.800 63.530 373.000 ;
        RECT 63.130 372.200 63.530 372.800 ;
        RECT 59.530 372.000 63.530 372.200 ;
        RECT 63.130 371.400 63.530 372.000 ;
        RECT 59.530 371.200 63.530 371.400 ;
        RECT 63.130 370.600 63.530 371.200 ;
        RECT 59.530 370.400 63.530 370.600 ;
        RECT 63.130 370.200 63.530 370.400 ;
        RECT 55.380 369.800 63.530 370.200 ;
        RECT 55.380 362.200 55.580 369.800 ;
        RECT 56.180 362.200 56.380 369.800 ;
        RECT 56.980 362.200 57.180 369.800 ;
        RECT 57.780 362.200 57.980 369.800 ;
        RECT 58.580 362.200 58.780 369.800 ;
        RECT 63.130 369.600 63.530 369.800 ;
        RECT 59.530 369.400 63.530 369.600 ;
        RECT 63.130 368.800 63.530 369.400 ;
        RECT 59.530 368.600 63.530 368.800 ;
        RECT 63.130 368.000 63.530 368.600 ;
        RECT 59.530 367.800 63.530 368.000 ;
        RECT 63.130 367.200 63.530 367.800 ;
        RECT 59.530 367.000 63.530 367.200 ;
        RECT 63.130 366.400 63.530 367.000 ;
        RECT 59.530 366.200 63.530 366.400 ;
        RECT 63.130 365.600 63.530 366.200 ;
        RECT 59.530 365.400 63.530 365.600 ;
        RECT 63.130 364.800 63.530 365.400 ;
        RECT 59.530 364.600 63.530 364.800 ;
        RECT 63.130 364.000 63.530 364.600 ;
        RECT 59.530 363.800 63.530 364.000 ;
        RECT 63.130 363.200 63.530 363.800 ;
        RECT 59.530 363.000 63.530 363.200 ;
        RECT 63.130 362.400 63.530 363.000 ;
        RECT 59.530 362.200 63.530 362.400 ;
        RECT 65.930 377.600 69.930 377.800 ;
        RECT 65.930 377.000 66.330 377.600 ;
        RECT 65.930 376.800 69.930 377.000 ;
        RECT 65.930 376.200 66.330 376.800 ;
        RECT 65.930 376.000 69.930 376.200 ;
        RECT 65.930 375.400 66.330 376.000 ;
        RECT 65.930 375.200 69.930 375.400 ;
        RECT 65.930 374.600 66.330 375.200 ;
        RECT 65.930 374.400 69.930 374.600 ;
        RECT 65.930 373.800 66.330 374.400 ;
        RECT 65.930 373.600 69.930 373.800 ;
        RECT 65.930 373.000 66.330 373.600 ;
        RECT 65.930 372.800 69.930 373.000 ;
        RECT 65.930 372.200 66.330 372.800 ;
        RECT 65.930 372.000 69.930 372.200 ;
        RECT 65.930 371.400 66.330 372.000 ;
        RECT 65.930 371.200 69.930 371.400 ;
        RECT 65.930 370.600 66.330 371.200 ;
        RECT 65.930 370.400 69.930 370.600 ;
        RECT 65.930 370.200 66.330 370.400 ;
        RECT 70.680 370.200 70.880 377.800 ;
        RECT 71.480 370.200 71.680 377.800 ;
        RECT 72.280 370.200 72.480 377.800 ;
        RECT 73.080 370.200 73.280 377.800 ;
        RECT 73.880 370.200 74.080 377.800 ;
        RECT 65.930 369.800 74.080 370.200 ;
        RECT 65.930 369.600 66.330 369.800 ;
        RECT 65.930 369.400 69.930 369.600 ;
        RECT 65.930 368.800 66.330 369.400 ;
        RECT 65.930 368.600 69.930 368.800 ;
        RECT 65.930 368.000 66.330 368.600 ;
        RECT 65.930 367.800 69.930 368.000 ;
        RECT 65.930 367.200 66.330 367.800 ;
        RECT 65.930 367.000 69.930 367.200 ;
        RECT 65.930 366.400 66.330 367.000 ;
        RECT 65.930 366.200 69.930 366.400 ;
        RECT 65.930 365.600 66.330 366.200 ;
        RECT 65.930 365.400 69.930 365.600 ;
        RECT 65.930 364.800 66.330 365.400 ;
        RECT 65.930 364.600 69.930 364.800 ;
        RECT 65.930 364.000 66.330 364.600 ;
        RECT 65.930 363.800 69.930 364.000 ;
        RECT 65.930 363.200 66.330 363.800 ;
        RECT 65.930 363.000 69.930 363.200 ;
        RECT 65.930 362.400 66.330 363.000 ;
        RECT 65.930 362.200 69.930 362.400 ;
        RECT 70.680 362.200 70.880 369.800 ;
        RECT 71.480 362.200 71.680 369.800 ;
        RECT 72.280 362.200 72.480 369.800 ;
        RECT 73.080 362.200 73.280 369.800 ;
        RECT 73.880 362.200 74.080 369.800 ;
        RECT 75.380 370.200 75.580 377.800 ;
        RECT 76.180 370.200 76.380 377.800 ;
        RECT 76.980 370.200 77.180 377.800 ;
        RECT 77.780 370.200 77.980 377.800 ;
        RECT 78.580 370.200 78.780 377.800 ;
        RECT 79.530 377.600 83.530 377.800 ;
        RECT 83.130 377.000 83.530 377.600 ;
        RECT 79.530 376.800 83.530 377.000 ;
        RECT 83.130 376.200 83.530 376.800 ;
        RECT 79.530 376.000 83.530 376.200 ;
        RECT 83.130 375.400 83.530 376.000 ;
        RECT 79.530 375.200 83.530 375.400 ;
        RECT 83.130 374.600 83.530 375.200 ;
        RECT 79.530 374.400 83.530 374.600 ;
        RECT 83.130 373.800 83.530 374.400 ;
        RECT 79.530 373.600 83.530 373.800 ;
        RECT 83.130 373.000 83.530 373.600 ;
        RECT 79.530 372.800 83.530 373.000 ;
        RECT 83.130 372.200 83.530 372.800 ;
        RECT 79.530 372.000 83.530 372.200 ;
        RECT 83.130 371.400 83.530 372.000 ;
        RECT 79.530 371.200 83.530 371.400 ;
        RECT 83.130 370.600 83.530 371.200 ;
        RECT 79.530 370.400 83.530 370.600 ;
        RECT 83.130 370.200 83.530 370.400 ;
        RECT 75.380 369.800 83.530 370.200 ;
        RECT 75.380 362.200 75.580 369.800 ;
        RECT 76.180 362.200 76.380 369.800 ;
        RECT 76.980 362.200 77.180 369.800 ;
        RECT 77.780 362.200 77.980 369.800 ;
        RECT 78.580 362.200 78.780 369.800 ;
        RECT 83.130 369.600 83.530 369.800 ;
        RECT 79.530 369.400 83.530 369.600 ;
        RECT 83.130 368.800 83.530 369.400 ;
        RECT 79.530 368.600 83.530 368.800 ;
        RECT 83.130 368.000 83.530 368.600 ;
        RECT 79.530 367.800 83.530 368.000 ;
        RECT 83.130 367.200 83.530 367.800 ;
        RECT 79.530 367.000 83.530 367.200 ;
        RECT 83.130 366.400 83.530 367.000 ;
        RECT 79.530 366.200 83.530 366.400 ;
        RECT 83.130 365.600 83.530 366.200 ;
        RECT 79.530 365.400 83.530 365.600 ;
        RECT 83.130 364.800 83.530 365.400 ;
        RECT 79.530 364.600 83.530 364.800 ;
        RECT 83.130 364.000 83.530 364.600 ;
        RECT 79.530 363.800 83.530 364.000 ;
        RECT 83.130 363.200 83.530 363.800 ;
        RECT 79.530 363.000 83.530 363.200 ;
        RECT 83.130 362.400 83.530 363.000 ;
        RECT 79.530 362.200 83.530 362.400 ;
        RECT 85.930 377.600 89.930 377.800 ;
        RECT 85.930 377.000 86.330 377.600 ;
        RECT 85.930 376.800 89.930 377.000 ;
        RECT 85.930 376.200 86.330 376.800 ;
        RECT 85.930 376.000 89.930 376.200 ;
        RECT 85.930 375.400 86.330 376.000 ;
        RECT 85.930 375.200 89.930 375.400 ;
        RECT 85.930 374.600 86.330 375.200 ;
        RECT 85.930 374.400 89.930 374.600 ;
        RECT 85.930 373.800 86.330 374.400 ;
        RECT 85.930 373.600 89.930 373.800 ;
        RECT 85.930 373.000 86.330 373.600 ;
        RECT 85.930 372.800 89.930 373.000 ;
        RECT 85.930 372.200 86.330 372.800 ;
        RECT 85.930 372.000 89.930 372.200 ;
        RECT 85.930 371.400 86.330 372.000 ;
        RECT 85.930 371.200 89.930 371.400 ;
        RECT 85.930 370.600 86.330 371.200 ;
        RECT 85.930 370.400 89.930 370.600 ;
        RECT 85.930 370.200 86.330 370.400 ;
        RECT 90.680 370.200 90.880 377.800 ;
        RECT 91.480 370.200 91.680 377.800 ;
        RECT 92.280 370.200 92.480 377.800 ;
        RECT 93.080 370.200 93.280 377.800 ;
        RECT 93.880 370.200 94.080 377.800 ;
        RECT 85.930 369.800 94.080 370.200 ;
        RECT 85.930 369.600 86.330 369.800 ;
        RECT 85.930 369.400 89.930 369.600 ;
        RECT 85.930 368.800 86.330 369.400 ;
        RECT 85.930 368.600 89.930 368.800 ;
        RECT 85.930 368.000 86.330 368.600 ;
        RECT 85.930 367.800 89.930 368.000 ;
        RECT 85.930 367.200 86.330 367.800 ;
        RECT 85.930 367.000 89.930 367.200 ;
        RECT 85.930 366.400 86.330 367.000 ;
        RECT 85.930 366.200 89.930 366.400 ;
        RECT 85.930 365.600 86.330 366.200 ;
        RECT 85.930 365.400 89.930 365.600 ;
        RECT 85.930 364.800 86.330 365.400 ;
        RECT 85.930 364.600 89.930 364.800 ;
        RECT 85.930 364.000 86.330 364.600 ;
        RECT 85.930 363.800 89.930 364.000 ;
        RECT 85.930 363.200 86.330 363.800 ;
        RECT 85.930 363.000 89.930 363.200 ;
        RECT 85.930 362.400 86.330 363.000 ;
        RECT 85.930 362.200 89.930 362.400 ;
        RECT 90.680 362.200 90.880 369.800 ;
        RECT 91.480 362.200 91.680 369.800 ;
        RECT 92.280 362.200 92.480 369.800 ;
        RECT 93.080 362.200 93.280 369.800 ;
        RECT 93.880 362.200 94.080 369.800 ;
        RECT 95.380 370.200 95.580 377.800 ;
        RECT 96.180 370.200 96.380 377.800 ;
        RECT 96.980 370.200 97.180 377.800 ;
        RECT 97.780 370.200 97.980 377.800 ;
        RECT 98.580 370.200 98.780 377.800 ;
        RECT 99.530 377.600 103.530 377.800 ;
        RECT 103.130 377.000 103.530 377.600 ;
        RECT 99.530 376.800 103.530 377.000 ;
        RECT 103.130 376.200 103.530 376.800 ;
        RECT 99.530 376.000 103.530 376.200 ;
        RECT 103.130 375.400 103.530 376.000 ;
        RECT 99.530 375.200 103.530 375.400 ;
        RECT 103.130 374.600 103.530 375.200 ;
        RECT 99.530 374.400 103.530 374.600 ;
        RECT 103.130 373.800 103.530 374.400 ;
        RECT 99.530 373.600 103.530 373.800 ;
        RECT 103.130 373.000 103.530 373.600 ;
        RECT 99.530 372.800 103.530 373.000 ;
        RECT 103.130 372.200 103.530 372.800 ;
        RECT 99.530 372.000 103.530 372.200 ;
        RECT 103.130 371.400 103.530 372.000 ;
        RECT 99.530 371.200 103.530 371.400 ;
        RECT 103.130 370.600 103.530 371.200 ;
        RECT 99.530 370.400 103.530 370.600 ;
        RECT 103.130 370.200 103.530 370.400 ;
        RECT 95.380 369.800 103.530 370.200 ;
        RECT 110.050 369.975 110.410 370.355 ;
        RECT 110.680 369.975 111.040 370.355 ;
        RECT 111.280 369.975 111.640 370.355 ;
        RECT 95.380 362.200 95.580 369.800 ;
        RECT 96.180 362.200 96.380 369.800 ;
        RECT 96.980 362.200 97.180 369.800 ;
        RECT 97.780 362.200 97.980 369.800 ;
        RECT 98.580 362.200 98.780 369.800 ;
        RECT 103.130 369.600 103.530 369.800 ;
        RECT 99.530 369.400 103.530 369.600 ;
        RECT 103.130 368.800 103.530 369.400 ;
        RECT 110.050 369.385 110.410 369.765 ;
        RECT 110.680 369.385 111.040 369.765 ;
        RECT 111.280 369.385 111.640 369.765 ;
        RECT 99.530 368.600 103.530 368.800 ;
        RECT 103.130 368.000 103.530 368.600 ;
        RECT 99.530 367.800 103.530 368.000 ;
        RECT 103.130 367.200 103.530 367.800 ;
        RECT 99.530 367.000 103.530 367.200 ;
        RECT 103.130 366.400 103.530 367.000 ;
        RECT 99.530 366.200 103.530 366.400 ;
        RECT 103.130 365.600 103.530 366.200 ;
        RECT 99.530 365.400 103.530 365.600 ;
        RECT 103.130 364.800 103.530 365.400 ;
        RECT 99.530 364.600 103.530 364.800 ;
        RECT 103.130 364.000 103.530 364.600 ;
        RECT 99.530 363.800 103.530 364.000 ;
        RECT 103.130 363.200 103.530 363.800 ;
        RECT 99.530 363.000 103.530 363.200 ;
        RECT 103.130 362.400 103.530 363.000 ;
        RECT 99.530 362.200 103.530 362.400 ;
        RECT 5.930 357.600 9.930 357.800 ;
        RECT 5.930 357.000 6.330 357.600 ;
        RECT 5.930 356.800 9.930 357.000 ;
        RECT 5.930 356.200 6.330 356.800 ;
        RECT 5.930 356.000 9.930 356.200 ;
        RECT 5.930 355.400 6.330 356.000 ;
        RECT 5.930 355.200 9.930 355.400 ;
        RECT 5.930 354.600 6.330 355.200 ;
        RECT 5.930 354.400 9.930 354.600 ;
        RECT 5.930 353.800 6.330 354.400 ;
        RECT 5.930 353.600 9.930 353.800 ;
        RECT 5.930 353.000 6.330 353.600 ;
        RECT 5.930 352.800 9.930 353.000 ;
        RECT 5.930 352.200 6.330 352.800 ;
        RECT 5.930 352.000 9.930 352.200 ;
        RECT 5.930 351.400 6.330 352.000 ;
        RECT 5.930 351.200 9.930 351.400 ;
        RECT 5.930 350.600 6.330 351.200 ;
        RECT 5.930 350.400 9.930 350.600 ;
        RECT 5.930 350.200 6.330 350.400 ;
        RECT 10.680 350.200 10.880 357.800 ;
        RECT 11.480 350.200 11.680 357.800 ;
        RECT 12.280 350.200 12.480 357.800 ;
        RECT 13.080 350.200 13.280 357.800 ;
        RECT 13.880 350.200 14.080 357.800 ;
        RECT 5.930 349.800 14.080 350.200 ;
        RECT 5.930 349.600 6.330 349.800 ;
        RECT 5.930 349.400 9.930 349.600 ;
        RECT 5.930 348.800 6.330 349.400 ;
        RECT 5.930 348.600 9.930 348.800 ;
        RECT 5.930 348.000 6.330 348.600 ;
        RECT 5.930 347.800 9.930 348.000 ;
        RECT 5.930 347.200 6.330 347.800 ;
        RECT 5.930 347.000 9.930 347.200 ;
        RECT 5.930 346.400 6.330 347.000 ;
        RECT 5.930 346.200 9.930 346.400 ;
        RECT 5.930 345.600 6.330 346.200 ;
        RECT 5.930 345.400 9.930 345.600 ;
        RECT 5.930 344.800 6.330 345.400 ;
        RECT 5.930 344.600 9.930 344.800 ;
        RECT 5.930 344.000 6.330 344.600 ;
        RECT 5.930 343.800 9.930 344.000 ;
        RECT 5.930 343.200 6.330 343.800 ;
        RECT 5.930 343.000 9.930 343.200 ;
        RECT 5.930 342.400 6.330 343.000 ;
        RECT 5.930 342.200 9.930 342.400 ;
        RECT 10.680 342.200 10.880 349.800 ;
        RECT 11.480 342.200 11.680 349.800 ;
        RECT 12.280 342.200 12.480 349.800 ;
        RECT 13.080 342.200 13.280 349.800 ;
        RECT 13.880 342.200 14.080 349.800 ;
        RECT 15.380 350.200 15.580 357.800 ;
        RECT 16.180 350.200 16.380 357.800 ;
        RECT 16.980 350.200 17.180 357.800 ;
        RECT 17.780 350.200 17.980 357.800 ;
        RECT 18.580 350.200 18.780 357.800 ;
        RECT 19.530 357.600 23.530 357.800 ;
        RECT 23.130 357.000 23.530 357.600 ;
        RECT 19.530 356.800 23.530 357.000 ;
        RECT 23.130 356.200 23.530 356.800 ;
        RECT 19.530 356.000 23.530 356.200 ;
        RECT 23.130 355.400 23.530 356.000 ;
        RECT 19.530 355.200 23.530 355.400 ;
        RECT 23.130 354.600 23.530 355.200 ;
        RECT 19.530 354.400 23.530 354.600 ;
        RECT 23.130 353.800 23.530 354.400 ;
        RECT 19.530 353.600 23.530 353.800 ;
        RECT 23.130 353.000 23.530 353.600 ;
        RECT 19.530 352.800 23.530 353.000 ;
        RECT 23.130 352.200 23.530 352.800 ;
        RECT 19.530 352.000 23.530 352.200 ;
        RECT 23.130 351.400 23.530 352.000 ;
        RECT 19.530 351.200 23.530 351.400 ;
        RECT 23.130 350.600 23.530 351.200 ;
        RECT 19.530 350.400 23.530 350.600 ;
        RECT 23.130 350.200 23.530 350.400 ;
        RECT 15.380 349.800 23.530 350.200 ;
        RECT 15.380 342.200 15.580 349.800 ;
        RECT 16.180 342.200 16.380 349.800 ;
        RECT 16.980 342.200 17.180 349.800 ;
        RECT 17.780 342.200 17.980 349.800 ;
        RECT 18.580 342.200 18.780 349.800 ;
        RECT 23.130 349.600 23.530 349.800 ;
        RECT 19.530 349.400 23.530 349.600 ;
        RECT 23.130 348.800 23.530 349.400 ;
        RECT 19.530 348.600 23.530 348.800 ;
        RECT 23.130 348.000 23.530 348.600 ;
        RECT 19.530 347.800 23.530 348.000 ;
        RECT 23.130 347.200 23.530 347.800 ;
        RECT 19.530 347.000 23.530 347.200 ;
        RECT 23.130 346.400 23.530 347.000 ;
        RECT 19.530 346.200 23.530 346.400 ;
        RECT 23.130 345.600 23.530 346.200 ;
        RECT 19.530 345.400 23.530 345.600 ;
        RECT 23.130 344.800 23.530 345.400 ;
        RECT 19.530 344.600 23.530 344.800 ;
        RECT 23.130 344.000 23.530 344.600 ;
        RECT 19.530 343.800 23.530 344.000 ;
        RECT 23.130 343.200 23.530 343.800 ;
        RECT 19.530 343.000 23.530 343.200 ;
        RECT 23.130 342.400 23.530 343.000 ;
        RECT 19.530 342.200 23.530 342.400 ;
        RECT 25.930 357.600 29.930 357.800 ;
        RECT 25.930 357.000 26.330 357.600 ;
        RECT 25.930 356.800 29.930 357.000 ;
        RECT 25.930 356.200 26.330 356.800 ;
        RECT 25.930 356.000 29.930 356.200 ;
        RECT 25.930 355.400 26.330 356.000 ;
        RECT 25.930 355.200 29.930 355.400 ;
        RECT 25.930 354.600 26.330 355.200 ;
        RECT 25.930 354.400 29.930 354.600 ;
        RECT 25.930 353.800 26.330 354.400 ;
        RECT 25.930 353.600 29.930 353.800 ;
        RECT 25.930 353.000 26.330 353.600 ;
        RECT 25.930 352.800 29.930 353.000 ;
        RECT 25.930 352.200 26.330 352.800 ;
        RECT 25.930 352.000 29.930 352.200 ;
        RECT 25.930 351.400 26.330 352.000 ;
        RECT 25.930 351.200 29.930 351.400 ;
        RECT 25.930 350.600 26.330 351.200 ;
        RECT 25.930 350.400 29.930 350.600 ;
        RECT 25.930 350.200 26.330 350.400 ;
        RECT 30.680 350.200 30.880 357.800 ;
        RECT 31.480 350.200 31.680 357.800 ;
        RECT 32.280 350.200 32.480 357.800 ;
        RECT 33.080 350.200 33.280 357.800 ;
        RECT 33.880 350.200 34.080 357.800 ;
        RECT 25.930 349.800 34.080 350.200 ;
        RECT 25.930 349.600 26.330 349.800 ;
        RECT 25.930 349.400 29.930 349.600 ;
        RECT 25.930 348.800 26.330 349.400 ;
        RECT 25.930 348.600 29.930 348.800 ;
        RECT 25.930 348.000 26.330 348.600 ;
        RECT 25.930 347.800 29.930 348.000 ;
        RECT 25.930 347.200 26.330 347.800 ;
        RECT 25.930 347.000 29.930 347.200 ;
        RECT 25.930 346.400 26.330 347.000 ;
        RECT 25.930 346.200 29.930 346.400 ;
        RECT 25.930 345.600 26.330 346.200 ;
        RECT 25.930 345.400 29.930 345.600 ;
        RECT 25.930 344.800 26.330 345.400 ;
        RECT 25.930 344.600 29.930 344.800 ;
        RECT 25.930 344.000 26.330 344.600 ;
        RECT 25.930 343.800 29.930 344.000 ;
        RECT 25.930 343.200 26.330 343.800 ;
        RECT 25.930 343.000 29.930 343.200 ;
        RECT 25.930 342.400 26.330 343.000 ;
        RECT 25.930 342.200 29.930 342.400 ;
        RECT 30.680 342.200 30.880 349.800 ;
        RECT 31.480 342.200 31.680 349.800 ;
        RECT 32.280 342.200 32.480 349.800 ;
        RECT 33.080 342.200 33.280 349.800 ;
        RECT 33.880 342.200 34.080 349.800 ;
        RECT 35.380 350.200 35.580 357.800 ;
        RECT 36.180 350.200 36.380 357.800 ;
        RECT 36.980 350.200 37.180 357.800 ;
        RECT 37.780 350.200 37.980 357.800 ;
        RECT 38.580 350.200 38.780 357.800 ;
        RECT 39.530 357.600 43.530 357.800 ;
        RECT 43.130 357.000 43.530 357.600 ;
        RECT 39.530 356.800 43.530 357.000 ;
        RECT 43.130 356.200 43.530 356.800 ;
        RECT 39.530 356.000 43.530 356.200 ;
        RECT 43.130 355.400 43.530 356.000 ;
        RECT 39.530 355.200 43.530 355.400 ;
        RECT 43.130 354.600 43.530 355.200 ;
        RECT 39.530 354.400 43.530 354.600 ;
        RECT 43.130 353.800 43.530 354.400 ;
        RECT 39.530 353.600 43.530 353.800 ;
        RECT 43.130 353.000 43.530 353.600 ;
        RECT 39.530 352.800 43.530 353.000 ;
        RECT 43.130 352.200 43.530 352.800 ;
        RECT 39.530 352.000 43.530 352.200 ;
        RECT 43.130 351.400 43.530 352.000 ;
        RECT 39.530 351.200 43.530 351.400 ;
        RECT 43.130 350.600 43.530 351.200 ;
        RECT 39.530 350.400 43.530 350.600 ;
        RECT 43.130 350.200 43.530 350.400 ;
        RECT 35.380 349.800 43.530 350.200 ;
        RECT 35.380 342.200 35.580 349.800 ;
        RECT 36.180 342.200 36.380 349.800 ;
        RECT 36.980 342.200 37.180 349.800 ;
        RECT 37.780 342.200 37.980 349.800 ;
        RECT 38.580 342.200 38.780 349.800 ;
        RECT 43.130 349.600 43.530 349.800 ;
        RECT 39.530 349.400 43.530 349.600 ;
        RECT 43.130 348.800 43.530 349.400 ;
        RECT 39.530 348.600 43.530 348.800 ;
        RECT 43.130 348.000 43.530 348.600 ;
        RECT 39.530 347.800 43.530 348.000 ;
        RECT 43.130 347.200 43.530 347.800 ;
        RECT 39.530 347.000 43.530 347.200 ;
        RECT 43.130 346.400 43.530 347.000 ;
        RECT 39.530 346.200 43.530 346.400 ;
        RECT 43.130 345.600 43.530 346.200 ;
        RECT 39.530 345.400 43.530 345.600 ;
        RECT 43.130 344.800 43.530 345.400 ;
        RECT 39.530 344.600 43.530 344.800 ;
        RECT 43.130 344.000 43.530 344.600 ;
        RECT 39.530 343.800 43.530 344.000 ;
        RECT 43.130 343.200 43.530 343.800 ;
        RECT 39.530 343.000 43.530 343.200 ;
        RECT 43.130 342.400 43.530 343.000 ;
        RECT 39.530 342.200 43.530 342.400 ;
        RECT 45.930 357.600 49.930 357.800 ;
        RECT 45.930 357.000 46.330 357.600 ;
        RECT 45.930 356.800 49.930 357.000 ;
        RECT 45.930 356.200 46.330 356.800 ;
        RECT 45.930 356.000 49.930 356.200 ;
        RECT 45.930 355.400 46.330 356.000 ;
        RECT 45.930 355.200 49.930 355.400 ;
        RECT 45.930 354.600 46.330 355.200 ;
        RECT 45.930 354.400 49.930 354.600 ;
        RECT 45.930 353.800 46.330 354.400 ;
        RECT 45.930 353.600 49.930 353.800 ;
        RECT 45.930 353.000 46.330 353.600 ;
        RECT 45.930 352.800 49.930 353.000 ;
        RECT 45.930 352.200 46.330 352.800 ;
        RECT 45.930 352.000 49.930 352.200 ;
        RECT 45.930 351.400 46.330 352.000 ;
        RECT 45.930 351.200 49.930 351.400 ;
        RECT 45.930 350.600 46.330 351.200 ;
        RECT 45.930 350.400 49.930 350.600 ;
        RECT 45.930 350.200 46.330 350.400 ;
        RECT 50.680 350.200 50.880 357.800 ;
        RECT 51.480 350.200 51.680 357.800 ;
        RECT 52.280 350.200 52.480 357.800 ;
        RECT 53.080 350.200 53.280 357.800 ;
        RECT 53.880 350.200 54.080 357.800 ;
        RECT 45.930 349.800 54.080 350.200 ;
        RECT 45.930 349.600 46.330 349.800 ;
        RECT 45.930 349.400 49.930 349.600 ;
        RECT 45.930 348.800 46.330 349.400 ;
        RECT 45.930 348.600 49.930 348.800 ;
        RECT 45.930 348.000 46.330 348.600 ;
        RECT 45.930 347.800 49.930 348.000 ;
        RECT 45.930 347.200 46.330 347.800 ;
        RECT 45.930 347.000 49.930 347.200 ;
        RECT 45.930 346.400 46.330 347.000 ;
        RECT 45.930 346.200 49.930 346.400 ;
        RECT 45.930 345.600 46.330 346.200 ;
        RECT 45.930 345.400 49.930 345.600 ;
        RECT 45.930 344.800 46.330 345.400 ;
        RECT 45.930 344.600 49.930 344.800 ;
        RECT 45.930 344.000 46.330 344.600 ;
        RECT 45.930 343.800 49.930 344.000 ;
        RECT 45.930 343.200 46.330 343.800 ;
        RECT 45.930 343.000 49.930 343.200 ;
        RECT 45.930 342.400 46.330 343.000 ;
        RECT 45.930 342.200 49.930 342.400 ;
        RECT 50.680 342.200 50.880 349.800 ;
        RECT 51.480 342.200 51.680 349.800 ;
        RECT 52.280 342.200 52.480 349.800 ;
        RECT 53.080 342.200 53.280 349.800 ;
        RECT 53.880 342.200 54.080 349.800 ;
        RECT 55.380 350.200 55.580 357.800 ;
        RECT 56.180 350.200 56.380 357.800 ;
        RECT 56.980 350.200 57.180 357.800 ;
        RECT 57.780 350.200 57.980 357.800 ;
        RECT 58.580 350.200 58.780 357.800 ;
        RECT 59.530 357.600 63.530 357.800 ;
        RECT 63.130 357.000 63.530 357.600 ;
        RECT 59.530 356.800 63.530 357.000 ;
        RECT 63.130 356.200 63.530 356.800 ;
        RECT 59.530 356.000 63.530 356.200 ;
        RECT 63.130 355.400 63.530 356.000 ;
        RECT 59.530 355.200 63.530 355.400 ;
        RECT 63.130 354.600 63.530 355.200 ;
        RECT 59.530 354.400 63.530 354.600 ;
        RECT 63.130 353.800 63.530 354.400 ;
        RECT 59.530 353.600 63.530 353.800 ;
        RECT 63.130 353.000 63.530 353.600 ;
        RECT 59.530 352.800 63.530 353.000 ;
        RECT 63.130 352.200 63.530 352.800 ;
        RECT 59.530 352.000 63.530 352.200 ;
        RECT 63.130 351.400 63.530 352.000 ;
        RECT 59.530 351.200 63.530 351.400 ;
        RECT 63.130 350.600 63.530 351.200 ;
        RECT 59.530 350.400 63.530 350.600 ;
        RECT 63.130 350.200 63.530 350.400 ;
        RECT 55.380 349.800 63.530 350.200 ;
        RECT 55.380 342.200 55.580 349.800 ;
        RECT 56.180 342.200 56.380 349.800 ;
        RECT 56.980 342.200 57.180 349.800 ;
        RECT 57.780 342.200 57.980 349.800 ;
        RECT 58.580 342.200 58.780 349.800 ;
        RECT 63.130 349.600 63.530 349.800 ;
        RECT 59.530 349.400 63.530 349.600 ;
        RECT 63.130 348.800 63.530 349.400 ;
        RECT 59.530 348.600 63.530 348.800 ;
        RECT 63.130 348.000 63.530 348.600 ;
        RECT 59.530 347.800 63.530 348.000 ;
        RECT 63.130 347.200 63.530 347.800 ;
        RECT 59.530 347.000 63.530 347.200 ;
        RECT 63.130 346.400 63.530 347.000 ;
        RECT 59.530 346.200 63.530 346.400 ;
        RECT 63.130 345.600 63.530 346.200 ;
        RECT 59.530 345.400 63.530 345.600 ;
        RECT 63.130 344.800 63.530 345.400 ;
        RECT 59.530 344.600 63.530 344.800 ;
        RECT 63.130 344.000 63.530 344.600 ;
        RECT 59.530 343.800 63.530 344.000 ;
        RECT 63.130 343.200 63.530 343.800 ;
        RECT 59.530 343.000 63.530 343.200 ;
        RECT 63.130 342.400 63.530 343.000 ;
        RECT 59.530 342.200 63.530 342.400 ;
        RECT 65.930 357.600 69.930 357.800 ;
        RECT 65.930 357.000 66.330 357.600 ;
        RECT 65.930 356.800 69.930 357.000 ;
        RECT 65.930 356.200 66.330 356.800 ;
        RECT 65.930 356.000 69.930 356.200 ;
        RECT 65.930 355.400 66.330 356.000 ;
        RECT 65.930 355.200 69.930 355.400 ;
        RECT 65.930 354.600 66.330 355.200 ;
        RECT 65.930 354.400 69.930 354.600 ;
        RECT 65.930 353.800 66.330 354.400 ;
        RECT 65.930 353.600 69.930 353.800 ;
        RECT 65.930 353.000 66.330 353.600 ;
        RECT 65.930 352.800 69.930 353.000 ;
        RECT 65.930 352.200 66.330 352.800 ;
        RECT 65.930 352.000 69.930 352.200 ;
        RECT 65.930 351.400 66.330 352.000 ;
        RECT 65.930 351.200 69.930 351.400 ;
        RECT 65.930 350.600 66.330 351.200 ;
        RECT 65.930 350.400 69.930 350.600 ;
        RECT 65.930 350.200 66.330 350.400 ;
        RECT 70.680 350.200 70.880 357.800 ;
        RECT 71.480 350.200 71.680 357.800 ;
        RECT 72.280 350.200 72.480 357.800 ;
        RECT 73.080 350.200 73.280 357.800 ;
        RECT 73.880 350.200 74.080 357.800 ;
        RECT 65.930 349.800 74.080 350.200 ;
        RECT 65.930 349.600 66.330 349.800 ;
        RECT 65.930 349.400 69.930 349.600 ;
        RECT 65.930 348.800 66.330 349.400 ;
        RECT 65.930 348.600 69.930 348.800 ;
        RECT 65.930 348.000 66.330 348.600 ;
        RECT 65.930 347.800 69.930 348.000 ;
        RECT 65.930 347.200 66.330 347.800 ;
        RECT 65.930 347.000 69.930 347.200 ;
        RECT 65.930 346.400 66.330 347.000 ;
        RECT 65.930 346.200 69.930 346.400 ;
        RECT 65.930 345.600 66.330 346.200 ;
        RECT 65.930 345.400 69.930 345.600 ;
        RECT 65.930 344.800 66.330 345.400 ;
        RECT 65.930 344.600 69.930 344.800 ;
        RECT 65.930 344.000 66.330 344.600 ;
        RECT 65.930 343.800 69.930 344.000 ;
        RECT 65.930 343.200 66.330 343.800 ;
        RECT 65.930 343.000 69.930 343.200 ;
        RECT 65.930 342.400 66.330 343.000 ;
        RECT 65.930 342.200 69.930 342.400 ;
        RECT 70.680 342.200 70.880 349.800 ;
        RECT 71.480 342.200 71.680 349.800 ;
        RECT 72.280 342.200 72.480 349.800 ;
        RECT 73.080 342.200 73.280 349.800 ;
        RECT 73.880 342.200 74.080 349.800 ;
        RECT 75.380 350.200 75.580 357.800 ;
        RECT 76.180 350.200 76.380 357.800 ;
        RECT 76.980 350.200 77.180 357.800 ;
        RECT 77.780 350.200 77.980 357.800 ;
        RECT 78.580 350.200 78.780 357.800 ;
        RECT 79.530 357.600 83.530 357.800 ;
        RECT 83.130 357.000 83.530 357.600 ;
        RECT 79.530 356.800 83.530 357.000 ;
        RECT 83.130 356.200 83.530 356.800 ;
        RECT 79.530 356.000 83.530 356.200 ;
        RECT 83.130 355.400 83.530 356.000 ;
        RECT 79.530 355.200 83.530 355.400 ;
        RECT 83.130 354.600 83.530 355.200 ;
        RECT 79.530 354.400 83.530 354.600 ;
        RECT 83.130 353.800 83.530 354.400 ;
        RECT 79.530 353.600 83.530 353.800 ;
        RECT 83.130 353.000 83.530 353.600 ;
        RECT 79.530 352.800 83.530 353.000 ;
        RECT 83.130 352.200 83.530 352.800 ;
        RECT 79.530 352.000 83.530 352.200 ;
        RECT 83.130 351.400 83.530 352.000 ;
        RECT 79.530 351.200 83.530 351.400 ;
        RECT 83.130 350.600 83.530 351.200 ;
        RECT 79.530 350.400 83.530 350.600 ;
        RECT 83.130 350.200 83.530 350.400 ;
        RECT 75.380 349.800 83.530 350.200 ;
        RECT 75.380 342.200 75.580 349.800 ;
        RECT 76.180 342.200 76.380 349.800 ;
        RECT 76.980 342.200 77.180 349.800 ;
        RECT 77.780 342.200 77.980 349.800 ;
        RECT 78.580 342.200 78.780 349.800 ;
        RECT 83.130 349.600 83.530 349.800 ;
        RECT 79.530 349.400 83.530 349.600 ;
        RECT 83.130 348.800 83.530 349.400 ;
        RECT 79.530 348.600 83.530 348.800 ;
        RECT 83.130 348.000 83.530 348.600 ;
        RECT 79.530 347.800 83.530 348.000 ;
        RECT 83.130 347.200 83.530 347.800 ;
        RECT 79.530 347.000 83.530 347.200 ;
        RECT 83.130 346.400 83.530 347.000 ;
        RECT 79.530 346.200 83.530 346.400 ;
        RECT 83.130 345.600 83.530 346.200 ;
        RECT 79.530 345.400 83.530 345.600 ;
        RECT 83.130 344.800 83.530 345.400 ;
        RECT 79.530 344.600 83.530 344.800 ;
        RECT 83.130 344.000 83.530 344.600 ;
        RECT 79.530 343.800 83.530 344.000 ;
        RECT 83.130 343.200 83.530 343.800 ;
        RECT 79.530 343.000 83.530 343.200 ;
        RECT 83.130 342.400 83.530 343.000 ;
        RECT 79.530 342.200 83.530 342.400 ;
        RECT 85.930 357.600 89.930 357.800 ;
        RECT 85.930 357.000 86.330 357.600 ;
        RECT 85.930 356.800 89.930 357.000 ;
        RECT 85.930 356.200 86.330 356.800 ;
        RECT 85.930 356.000 89.930 356.200 ;
        RECT 85.930 355.400 86.330 356.000 ;
        RECT 85.930 355.200 89.930 355.400 ;
        RECT 85.930 354.600 86.330 355.200 ;
        RECT 85.930 354.400 89.930 354.600 ;
        RECT 85.930 353.800 86.330 354.400 ;
        RECT 85.930 353.600 89.930 353.800 ;
        RECT 85.930 353.000 86.330 353.600 ;
        RECT 85.930 352.800 89.930 353.000 ;
        RECT 85.930 352.200 86.330 352.800 ;
        RECT 85.930 352.000 89.930 352.200 ;
        RECT 85.930 351.400 86.330 352.000 ;
        RECT 85.930 351.200 89.930 351.400 ;
        RECT 85.930 350.600 86.330 351.200 ;
        RECT 85.930 350.400 89.930 350.600 ;
        RECT 85.930 350.200 86.330 350.400 ;
        RECT 90.680 350.200 90.880 357.800 ;
        RECT 91.480 350.200 91.680 357.800 ;
        RECT 92.280 350.200 92.480 357.800 ;
        RECT 93.080 350.200 93.280 357.800 ;
        RECT 93.880 350.200 94.080 357.800 ;
        RECT 85.930 349.800 94.080 350.200 ;
        RECT 85.930 349.600 86.330 349.800 ;
        RECT 85.930 349.400 89.930 349.600 ;
        RECT 85.930 348.800 86.330 349.400 ;
        RECT 85.930 348.600 89.930 348.800 ;
        RECT 85.930 348.000 86.330 348.600 ;
        RECT 85.930 347.800 89.930 348.000 ;
        RECT 85.930 347.200 86.330 347.800 ;
        RECT 85.930 347.000 89.930 347.200 ;
        RECT 85.930 346.400 86.330 347.000 ;
        RECT 85.930 346.200 89.930 346.400 ;
        RECT 85.930 345.600 86.330 346.200 ;
        RECT 85.930 345.400 89.930 345.600 ;
        RECT 85.930 344.800 86.330 345.400 ;
        RECT 85.930 344.600 89.930 344.800 ;
        RECT 85.930 344.000 86.330 344.600 ;
        RECT 85.930 343.800 89.930 344.000 ;
        RECT 85.930 343.200 86.330 343.800 ;
        RECT 85.930 343.000 89.930 343.200 ;
        RECT 85.930 342.400 86.330 343.000 ;
        RECT 85.930 342.200 89.930 342.400 ;
        RECT 90.680 342.200 90.880 349.800 ;
        RECT 91.480 342.200 91.680 349.800 ;
        RECT 92.280 342.200 92.480 349.800 ;
        RECT 93.080 342.200 93.280 349.800 ;
        RECT 93.880 342.200 94.080 349.800 ;
        RECT 95.380 350.200 95.580 357.800 ;
        RECT 96.180 350.200 96.380 357.800 ;
        RECT 96.980 350.200 97.180 357.800 ;
        RECT 97.780 350.200 97.980 357.800 ;
        RECT 98.580 350.200 98.780 357.800 ;
        RECT 99.530 357.600 103.530 357.800 ;
        RECT 103.130 357.000 103.530 357.600 ;
        RECT 99.530 356.800 103.530 357.000 ;
        RECT 103.130 356.200 103.530 356.800 ;
        RECT 99.530 356.000 103.530 356.200 ;
        RECT 103.130 355.400 103.530 356.000 ;
        RECT 99.530 355.200 103.530 355.400 ;
        RECT 103.130 354.600 103.530 355.200 ;
        RECT 99.530 354.400 103.530 354.600 ;
        RECT 103.130 353.800 103.530 354.400 ;
        RECT 99.530 353.600 103.530 353.800 ;
        RECT 103.130 353.000 103.530 353.600 ;
        RECT 99.530 352.800 103.530 353.000 ;
        RECT 103.130 352.200 103.530 352.800 ;
        RECT 99.530 352.000 103.530 352.200 ;
        RECT 103.130 351.400 103.530 352.000 ;
        RECT 99.530 351.200 103.530 351.400 ;
        RECT 103.130 350.600 103.530 351.200 ;
        RECT 99.530 350.400 103.530 350.600 ;
        RECT 103.130 350.200 103.530 350.400 ;
        RECT 95.380 349.800 103.530 350.200 ;
        RECT 110.050 349.975 110.410 350.355 ;
        RECT 110.680 349.975 111.040 350.355 ;
        RECT 111.280 349.975 111.640 350.355 ;
        RECT 95.380 342.200 95.580 349.800 ;
        RECT 96.180 342.200 96.380 349.800 ;
        RECT 96.980 342.200 97.180 349.800 ;
        RECT 97.780 342.200 97.980 349.800 ;
        RECT 98.580 342.200 98.780 349.800 ;
        RECT 103.130 349.600 103.530 349.800 ;
        RECT 99.530 349.400 103.530 349.600 ;
        RECT 103.130 348.800 103.530 349.400 ;
        RECT 110.050 349.385 110.410 349.765 ;
        RECT 110.680 349.385 111.040 349.765 ;
        RECT 111.280 349.385 111.640 349.765 ;
        RECT 99.530 348.600 103.530 348.800 ;
        RECT 103.130 348.000 103.530 348.600 ;
        RECT 99.530 347.800 103.530 348.000 ;
        RECT 103.130 347.200 103.530 347.800 ;
        RECT 99.530 347.000 103.530 347.200 ;
        RECT 103.130 346.400 103.530 347.000 ;
        RECT 99.530 346.200 103.530 346.400 ;
        RECT 103.130 345.600 103.530 346.200 ;
        RECT 99.530 345.400 103.530 345.600 ;
        RECT 103.130 344.800 103.530 345.400 ;
        RECT 99.530 344.600 103.530 344.800 ;
        RECT 103.130 344.000 103.530 344.600 ;
        RECT 99.530 343.800 103.530 344.000 ;
        RECT 103.130 343.200 103.530 343.800 ;
        RECT 99.530 343.000 103.530 343.200 ;
        RECT 103.130 342.400 103.530 343.000 ;
        RECT 99.530 342.200 103.530 342.400 ;
        RECT 5.930 337.600 9.930 337.800 ;
        RECT 5.930 337.000 6.330 337.600 ;
        RECT 5.930 336.800 9.930 337.000 ;
        RECT 5.930 336.200 6.330 336.800 ;
        RECT 5.930 336.000 9.930 336.200 ;
        RECT 5.930 335.400 6.330 336.000 ;
        RECT 5.930 335.200 9.930 335.400 ;
        RECT 5.930 334.600 6.330 335.200 ;
        RECT 5.930 334.400 9.930 334.600 ;
        RECT 5.930 333.800 6.330 334.400 ;
        RECT 5.930 333.600 9.930 333.800 ;
        RECT 5.930 333.000 6.330 333.600 ;
        RECT 5.930 332.800 9.930 333.000 ;
        RECT 5.930 332.200 6.330 332.800 ;
        RECT 5.930 332.000 9.930 332.200 ;
        RECT 5.930 331.400 6.330 332.000 ;
        RECT 5.930 331.200 9.930 331.400 ;
        RECT 5.930 330.600 6.330 331.200 ;
        RECT 5.930 330.400 9.930 330.600 ;
        RECT 5.930 330.200 6.330 330.400 ;
        RECT 10.680 330.200 10.880 337.800 ;
        RECT 11.480 330.200 11.680 337.800 ;
        RECT 12.280 330.200 12.480 337.800 ;
        RECT 13.080 330.200 13.280 337.800 ;
        RECT 13.880 330.200 14.080 337.800 ;
        RECT 5.930 329.800 14.080 330.200 ;
        RECT 5.930 329.600 6.330 329.800 ;
        RECT 5.930 329.400 9.930 329.600 ;
        RECT 5.930 328.800 6.330 329.400 ;
        RECT 5.930 328.600 9.930 328.800 ;
        RECT 5.930 328.000 6.330 328.600 ;
        RECT 5.930 327.800 9.930 328.000 ;
        RECT 5.930 327.200 6.330 327.800 ;
        RECT 5.930 327.000 9.930 327.200 ;
        RECT 5.930 326.400 6.330 327.000 ;
        RECT 5.930 326.200 9.930 326.400 ;
        RECT 5.930 325.600 6.330 326.200 ;
        RECT 5.930 325.400 9.930 325.600 ;
        RECT 5.930 324.800 6.330 325.400 ;
        RECT 5.930 324.600 9.930 324.800 ;
        RECT 5.930 324.000 6.330 324.600 ;
        RECT 5.930 323.800 9.930 324.000 ;
        RECT 5.930 323.200 6.330 323.800 ;
        RECT 5.930 323.000 9.930 323.200 ;
        RECT 5.930 322.400 6.330 323.000 ;
        RECT 5.930 322.200 9.930 322.400 ;
        RECT 10.680 322.200 10.880 329.800 ;
        RECT 11.480 322.200 11.680 329.800 ;
        RECT 12.280 322.200 12.480 329.800 ;
        RECT 13.080 322.200 13.280 329.800 ;
        RECT 13.880 322.200 14.080 329.800 ;
        RECT 15.380 330.200 15.580 337.800 ;
        RECT 16.180 330.200 16.380 337.800 ;
        RECT 16.980 330.200 17.180 337.800 ;
        RECT 17.780 330.200 17.980 337.800 ;
        RECT 18.580 330.200 18.780 337.800 ;
        RECT 19.530 337.600 23.530 337.800 ;
        RECT 23.130 337.000 23.530 337.600 ;
        RECT 19.530 336.800 23.530 337.000 ;
        RECT 23.130 336.200 23.530 336.800 ;
        RECT 19.530 336.000 23.530 336.200 ;
        RECT 23.130 335.400 23.530 336.000 ;
        RECT 19.530 335.200 23.530 335.400 ;
        RECT 23.130 334.600 23.530 335.200 ;
        RECT 19.530 334.400 23.530 334.600 ;
        RECT 23.130 333.800 23.530 334.400 ;
        RECT 19.530 333.600 23.530 333.800 ;
        RECT 23.130 333.000 23.530 333.600 ;
        RECT 19.530 332.800 23.530 333.000 ;
        RECT 23.130 332.200 23.530 332.800 ;
        RECT 19.530 332.000 23.530 332.200 ;
        RECT 23.130 331.400 23.530 332.000 ;
        RECT 19.530 331.200 23.530 331.400 ;
        RECT 23.130 330.600 23.530 331.200 ;
        RECT 19.530 330.400 23.530 330.600 ;
        RECT 23.130 330.200 23.530 330.400 ;
        RECT 15.380 329.800 23.530 330.200 ;
        RECT 15.380 322.200 15.580 329.800 ;
        RECT 16.180 322.200 16.380 329.800 ;
        RECT 16.980 322.200 17.180 329.800 ;
        RECT 17.780 322.200 17.980 329.800 ;
        RECT 18.580 322.200 18.780 329.800 ;
        RECT 23.130 329.600 23.530 329.800 ;
        RECT 19.530 329.400 23.530 329.600 ;
        RECT 23.130 328.800 23.530 329.400 ;
        RECT 19.530 328.600 23.530 328.800 ;
        RECT 23.130 328.000 23.530 328.600 ;
        RECT 19.530 327.800 23.530 328.000 ;
        RECT 23.130 327.200 23.530 327.800 ;
        RECT 19.530 327.000 23.530 327.200 ;
        RECT 23.130 326.400 23.530 327.000 ;
        RECT 19.530 326.200 23.530 326.400 ;
        RECT 23.130 325.600 23.530 326.200 ;
        RECT 19.530 325.400 23.530 325.600 ;
        RECT 23.130 324.800 23.530 325.400 ;
        RECT 19.530 324.600 23.530 324.800 ;
        RECT 23.130 324.000 23.530 324.600 ;
        RECT 19.530 323.800 23.530 324.000 ;
        RECT 23.130 323.200 23.530 323.800 ;
        RECT 19.530 323.000 23.530 323.200 ;
        RECT 23.130 322.400 23.530 323.000 ;
        RECT 19.530 322.200 23.530 322.400 ;
        RECT 25.930 337.600 29.930 337.800 ;
        RECT 25.930 337.000 26.330 337.600 ;
        RECT 25.930 336.800 29.930 337.000 ;
        RECT 25.930 336.200 26.330 336.800 ;
        RECT 25.930 336.000 29.930 336.200 ;
        RECT 25.930 335.400 26.330 336.000 ;
        RECT 25.930 335.200 29.930 335.400 ;
        RECT 25.930 334.600 26.330 335.200 ;
        RECT 25.930 334.400 29.930 334.600 ;
        RECT 25.930 333.800 26.330 334.400 ;
        RECT 25.930 333.600 29.930 333.800 ;
        RECT 25.930 333.000 26.330 333.600 ;
        RECT 25.930 332.800 29.930 333.000 ;
        RECT 25.930 332.200 26.330 332.800 ;
        RECT 25.930 332.000 29.930 332.200 ;
        RECT 25.930 331.400 26.330 332.000 ;
        RECT 25.930 331.200 29.930 331.400 ;
        RECT 25.930 330.600 26.330 331.200 ;
        RECT 25.930 330.400 29.930 330.600 ;
        RECT 25.930 330.200 26.330 330.400 ;
        RECT 30.680 330.200 30.880 337.800 ;
        RECT 31.480 330.200 31.680 337.800 ;
        RECT 32.280 330.200 32.480 337.800 ;
        RECT 33.080 330.200 33.280 337.800 ;
        RECT 33.880 330.200 34.080 337.800 ;
        RECT 25.930 329.800 34.080 330.200 ;
        RECT 25.930 329.600 26.330 329.800 ;
        RECT 25.930 329.400 29.930 329.600 ;
        RECT 25.930 328.800 26.330 329.400 ;
        RECT 25.930 328.600 29.930 328.800 ;
        RECT 25.930 328.000 26.330 328.600 ;
        RECT 25.930 327.800 29.930 328.000 ;
        RECT 25.930 327.200 26.330 327.800 ;
        RECT 25.930 327.000 29.930 327.200 ;
        RECT 25.930 326.400 26.330 327.000 ;
        RECT 25.930 326.200 29.930 326.400 ;
        RECT 25.930 325.600 26.330 326.200 ;
        RECT 25.930 325.400 29.930 325.600 ;
        RECT 25.930 324.800 26.330 325.400 ;
        RECT 25.930 324.600 29.930 324.800 ;
        RECT 25.930 324.000 26.330 324.600 ;
        RECT 25.930 323.800 29.930 324.000 ;
        RECT 25.930 323.200 26.330 323.800 ;
        RECT 25.930 323.000 29.930 323.200 ;
        RECT 25.930 322.400 26.330 323.000 ;
        RECT 25.930 322.200 29.930 322.400 ;
        RECT 30.680 322.200 30.880 329.800 ;
        RECT 31.480 322.200 31.680 329.800 ;
        RECT 32.280 322.200 32.480 329.800 ;
        RECT 33.080 322.200 33.280 329.800 ;
        RECT 33.880 322.200 34.080 329.800 ;
        RECT 35.380 330.200 35.580 337.800 ;
        RECT 36.180 330.200 36.380 337.800 ;
        RECT 36.980 330.200 37.180 337.800 ;
        RECT 37.780 330.200 37.980 337.800 ;
        RECT 38.580 330.200 38.780 337.800 ;
        RECT 39.530 337.600 43.530 337.800 ;
        RECT 43.130 337.000 43.530 337.600 ;
        RECT 39.530 336.800 43.530 337.000 ;
        RECT 43.130 336.200 43.530 336.800 ;
        RECT 39.530 336.000 43.530 336.200 ;
        RECT 43.130 335.400 43.530 336.000 ;
        RECT 39.530 335.200 43.530 335.400 ;
        RECT 43.130 334.600 43.530 335.200 ;
        RECT 39.530 334.400 43.530 334.600 ;
        RECT 43.130 333.800 43.530 334.400 ;
        RECT 39.530 333.600 43.530 333.800 ;
        RECT 43.130 333.000 43.530 333.600 ;
        RECT 39.530 332.800 43.530 333.000 ;
        RECT 43.130 332.200 43.530 332.800 ;
        RECT 39.530 332.000 43.530 332.200 ;
        RECT 43.130 331.400 43.530 332.000 ;
        RECT 39.530 331.200 43.530 331.400 ;
        RECT 43.130 330.600 43.530 331.200 ;
        RECT 39.530 330.400 43.530 330.600 ;
        RECT 43.130 330.200 43.530 330.400 ;
        RECT 35.380 329.800 43.530 330.200 ;
        RECT 35.380 322.200 35.580 329.800 ;
        RECT 36.180 322.200 36.380 329.800 ;
        RECT 36.980 322.200 37.180 329.800 ;
        RECT 37.780 322.200 37.980 329.800 ;
        RECT 38.580 322.200 38.780 329.800 ;
        RECT 43.130 329.600 43.530 329.800 ;
        RECT 39.530 329.400 43.530 329.600 ;
        RECT 43.130 328.800 43.530 329.400 ;
        RECT 39.530 328.600 43.530 328.800 ;
        RECT 43.130 328.000 43.530 328.600 ;
        RECT 39.530 327.800 43.530 328.000 ;
        RECT 43.130 327.200 43.530 327.800 ;
        RECT 39.530 327.000 43.530 327.200 ;
        RECT 43.130 326.400 43.530 327.000 ;
        RECT 39.530 326.200 43.530 326.400 ;
        RECT 43.130 325.600 43.530 326.200 ;
        RECT 39.530 325.400 43.530 325.600 ;
        RECT 43.130 324.800 43.530 325.400 ;
        RECT 39.530 324.600 43.530 324.800 ;
        RECT 43.130 324.000 43.530 324.600 ;
        RECT 39.530 323.800 43.530 324.000 ;
        RECT 43.130 323.200 43.530 323.800 ;
        RECT 39.530 323.000 43.530 323.200 ;
        RECT 43.130 322.400 43.530 323.000 ;
        RECT 39.530 322.200 43.530 322.400 ;
        RECT 45.930 337.600 49.930 337.800 ;
        RECT 45.930 337.000 46.330 337.600 ;
        RECT 45.930 336.800 49.930 337.000 ;
        RECT 45.930 336.200 46.330 336.800 ;
        RECT 45.930 336.000 49.930 336.200 ;
        RECT 45.930 335.400 46.330 336.000 ;
        RECT 45.930 335.200 49.930 335.400 ;
        RECT 45.930 334.600 46.330 335.200 ;
        RECT 45.930 334.400 49.930 334.600 ;
        RECT 45.930 333.800 46.330 334.400 ;
        RECT 45.930 333.600 49.930 333.800 ;
        RECT 45.930 333.000 46.330 333.600 ;
        RECT 45.930 332.800 49.930 333.000 ;
        RECT 45.930 332.200 46.330 332.800 ;
        RECT 45.930 332.000 49.930 332.200 ;
        RECT 45.930 331.400 46.330 332.000 ;
        RECT 45.930 331.200 49.930 331.400 ;
        RECT 45.930 330.600 46.330 331.200 ;
        RECT 45.930 330.400 49.930 330.600 ;
        RECT 45.930 330.200 46.330 330.400 ;
        RECT 50.680 330.200 50.880 337.800 ;
        RECT 51.480 330.200 51.680 337.800 ;
        RECT 52.280 330.200 52.480 337.800 ;
        RECT 53.080 330.200 53.280 337.800 ;
        RECT 53.880 330.200 54.080 337.800 ;
        RECT 45.930 329.800 54.080 330.200 ;
        RECT 45.930 329.600 46.330 329.800 ;
        RECT 45.930 329.400 49.930 329.600 ;
        RECT 45.930 328.800 46.330 329.400 ;
        RECT 45.930 328.600 49.930 328.800 ;
        RECT 45.930 328.000 46.330 328.600 ;
        RECT 45.930 327.800 49.930 328.000 ;
        RECT 45.930 327.200 46.330 327.800 ;
        RECT 45.930 327.000 49.930 327.200 ;
        RECT 45.930 326.400 46.330 327.000 ;
        RECT 45.930 326.200 49.930 326.400 ;
        RECT 45.930 325.600 46.330 326.200 ;
        RECT 45.930 325.400 49.930 325.600 ;
        RECT 45.930 324.800 46.330 325.400 ;
        RECT 45.930 324.600 49.930 324.800 ;
        RECT 45.930 324.000 46.330 324.600 ;
        RECT 45.930 323.800 49.930 324.000 ;
        RECT 45.930 323.200 46.330 323.800 ;
        RECT 45.930 323.000 49.930 323.200 ;
        RECT 45.930 322.400 46.330 323.000 ;
        RECT 45.930 322.200 49.930 322.400 ;
        RECT 50.680 322.200 50.880 329.800 ;
        RECT 51.480 322.200 51.680 329.800 ;
        RECT 52.280 322.200 52.480 329.800 ;
        RECT 53.080 322.200 53.280 329.800 ;
        RECT 53.880 322.200 54.080 329.800 ;
        RECT 55.380 330.200 55.580 337.800 ;
        RECT 56.180 330.200 56.380 337.800 ;
        RECT 56.980 330.200 57.180 337.800 ;
        RECT 57.780 330.200 57.980 337.800 ;
        RECT 58.580 330.200 58.780 337.800 ;
        RECT 59.530 337.600 63.530 337.800 ;
        RECT 63.130 337.000 63.530 337.600 ;
        RECT 59.530 336.800 63.530 337.000 ;
        RECT 63.130 336.200 63.530 336.800 ;
        RECT 59.530 336.000 63.530 336.200 ;
        RECT 63.130 335.400 63.530 336.000 ;
        RECT 59.530 335.200 63.530 335.400 ;
        RECT 63.130 334.600 63.530 335.200 ;
        RECT 59.530 334.400 63.530 334.600 ;
        RECT 63.130 333.800 63.530 334.400 ;
        RECT 59.530 333.600 63.530 333.800 ;
        RECT 63.130 333.000 63.530 333.600 ;
        RECT 59.530 332.800 63.530 333.000 ;
        RECT 63.130 332.200 63.530 332.800 ;
        RECT 59.530 332.000 63.530 332.200 ;
        RECT 63.130 331.400 63.530 332.000 ;
        RECT 59.530 331.200 63.530 331.400 ;
        RECT 63.130 330.600 63.530 331.200 ;
        RECT 59.530 330.400 63.530 330.600 ;
        RECT 63.130 330.200 63.530 330.400 ;
        RECT 55.380 329.800 63.530 330.200 ;
        RECT 55.380 322.200 55.580 329.800 ;
        RECT 56.180 322.200 56.380 329.800 ;
        RECT 56.980 322.200 57.180 329.800 ;
        RECT 57.780 322.200 57.980 329.800 ;
        RECT 58.580 322.200 58.780 329.800 ;
        RECT 63.130 329.600 63.530 329.800 ;
        RECT 59.530 329.400 63.530 329.600 ;
        RECT 63.130 328.800 63.530 329.400 ;
        RECT 59.530 328.600 63.530 328.800 ;
        RECT 63.130 328.000 63.530 328.600 ;
        RECT 59.530 327.800 63.530 328.000 ;
        RECT 63.130 327.200 63.530 327.800 ;
        RECT 59.530 327.000 63.530 327.200 ;
        RECT 63.130 326.400 63.530 327.000 ;
        RECT 59.530 326.200 63.530 326.400 ;
        RECT 63.130 325.600 63.530 326.200 ;
        RECT 59.530 325.400 63.530 325.600 ;
        RECT 63.130 324.800 63.530 325.400 ;
        RECT 59.530 324.600 63.530 324.800 ;
        RECT 63.130 324.000 63.530 324.600 ;
        RECT 59.530 323.800 63.530 324.000 ;
        RECT 63.130 323.200 63.530 323.800 ;
        RECT 59.530 323.000 63.530 323.200 ;
        RECT 63.130 322.400 63.530 323.000 ;
        RECT 59.530 322.200 63.530 322.400 ;
        RECT 65.930 337.600 69.930 337.800 ;
        RECT 65.930 337.000 66.330 337.600 ;
        RECT 65.930 336.800 69.930 337.000 ;
        RECT 65.930 336.200 66.330 336.800 ;
        RECT 65.930 336.000 69.930 336.200 ;
        RECT 65.930 335.400 66.330 336.000 ;
        RECT 65.930 335.200 69.930 335.400 ;
        RECT 65.930 334.600 66.330 335.200 ;
        RECT 65.930 334.400 69.930 334.600 ;
        RECT 65.930 333.800 66.330 334.400 ;
        RECT 65.930 333.600 69.930 333.800 ;
        RECT 65.930 333.000 66.330 333.600 ;
        RECT 65.930 332.800 69.930 333.000 ;
        RECT 65.930 332.200 66.330 332.800 ;
        RECT 65.930 332.000 69.930 332.200 ;
        RECT 65.930 331.400 66.330 332.000 ;
        RECT 65.930 331.200 69.930 331.400 ;
        RECT 65.930 330.600 66.330 331.200 ;
        RECT 65.930 330.400 69.930 330.600 ;
        RECT 65.930 330.200 66.330 330.400 ;
        RECT 70.680 330.200 70.880 337.800 ;
        RECT 71.480 330.200 71.680 337.800 ;
        RECT 72.280 330.200 72.480 337.800 ;
        RECT 73.080 330.200 73.280 337.800 ;
        RECT 73.880 330.200 74.080 337.800 ;
        RECT 65.930 329.800 74.080 330.200 ;
        RECT 65.930 329.600 66.330 329.800 ;
        RECT 65.930 329.400 69.930 329.600 ;
        RECT 65.930 328.800 66.330 329.400 ;
        RECT 65.930 328.600 69.930 328.800 ;
        RECT 65.930 328.000 66.330 328.600 ;
        RECT 65.930 327.800 69.930 328.000 ;
        RECT 65.930 327.200 66.330 327.800 ;
        RECT 65.930 327.000 69.930 327.200 ;
        RECT 65.930 326.400 66.330 327.000 ;
        RECT 65.930 326.200 69.930 326.400 ;
        RECT 65.930 325.600 66.330 326.200 ;
        RECT 65.930 325.400 69.930 325.600 ;
        RECT 65.930 324.800 66.330 325.400 ;
        RECT 65.930 324.600 69.930 324.800 ;
        RECT 65.930 324.000 66.330 324.600 ;
        RECT 65.930 323.800 69.930 324.000 ;
        RECT 65.930 323.200 66.330 323.800 ;
        RECT 65.930 323.000 69.930 323.200 ;
        RECT 65.930 322.400 66.330 323.000 ;
        RECT 65.930 322.200 69.930 322.400 ;
        RECT 70.680 322.200 70.880 329.800 ;
        RECT 71.480 322.200 71.680 329.800 ;
        RECT 72.280 322.200 72.480 329.800 ;
        RECT 73.080 322.200 73.280 329.800 ;
        RECT 73.880 322.200 74.080 329.800 ;
        RECT 75.380 330.200 75.580 337.800 ;
        RECT 76.180 330.200 76.380 337.800 ;
        RECT 76.980 330.200 77.180 337.800 ;
        RECT 77.780 330.200 77.980 337.800 ;
        RECT 78.580 330.200 78.780 337.800 ;
        RECT 79.530 337.600 83.530 337.800 ;
        RECT 83.130 337.000 83.530 337.600 ;
        RECT 79.530 336.800 83.530 337.000 ;
        RECT 83.130 336.200 83.530 336.800 ;
        RECT 79.530 336.000 83.530 336.200 ;
        RECT 83.130 335.400 83.530 336.000 ;
        RECT 79.530 335.200 83.530 335.400 ;
        RECT 83.130 334.600 83.530 335.200 ;
        RECT 79.530 334.400 83.530 334.600 ;
        RECT 83.130 333.800 83.530 334.400 ;
        RECT 79.530 333.600 83.530 333.800 ;
        RECT 83.130 333.000 83.530 333.600 ;
        RECT 79.530 332.800 83.530 333.000 ;
        RECT 83.130 332.200 83.530 332.800 ;
        RECT 79.530 332.000 83.530 332.200 ;
        RECT 83.130 331.400 83.530 332.000 ;
        RECT 79.530 331.200 83.530 331.400 ;
        RECT 83.130 330.600 83.530 331.200 ;
        RECT 79.530 330.400 83.530 330.600 ;
        RECT 83.130 330.200 83.530 330.400 ;
        RECT 75.380 329.800 83.530 330.200 ;
        RECT 75.380 322.200 75.580 329.800 ;
        RECT 76.180 322.200 76.380 329.800 ;
        RECT 76.980 322.200 77.180 329.800 ;
        RECT 77.780 322.200 77.980 329.800 ;
        RECT 78.580 322.200 78.780 329.800 ;
        RECT 83.130 329.600 83.530 329.800 ;
        RECT 79.530 329.400 83.530 329.600 ;
        RECT 83.130 328.800 83.530 329.400 ;
        RECT 79.530 328.600 83.530 328.800 ;
        RECT 83.130 328.000 83.530 328.600 ;
        RECT 79.530 327.800 83.530 328.000 ;
        RECT 83.130 327.200 83.530 327.800 ;
        RECT 79.530 327.000 83.530 327.200 ;
        RECT 83.130 326.400 83.530 327.000 ;
        RECT 79.530 326.200 83.530 326.400 ;
        RECT 83.130 325.600 83.530 326.200 ;
        RECT 79.530 325.400 83.530 325.600 ;
        RECT 83.130 324.800 83.530 325.400 ;
        RECT 79.530 324.600 83.530 324.800 ;
        RECT 83.130 324.000 83.530 324.600 ;
        RECT 79.530 323.800 83.530 324.000 ;
        RECT 83.130 323.200 83.530 323.800 ;
        RECT 79.530 323.000 83.530 323.200 ;
        RECT 83.130 322.400 83.530 323.000 ;
        RECT 79.530 322.200 83.530 322.400 ;
        RECT 85.930 337.600 89.930 337.800 ;
        RECT 85.930 337.000 86.330 337.600 ;
        RECT 85.930 336.800 89.930 337.000 ;
        RECT 85.930 336.200 86.330 336.800 ;
        RECT 85.930 336.000 89.930 336.200 ;
        RECT 85.930 335.400 86.330 336.000 ;
        RECT 85.930 335.200 89.930 335.400 ;
        RECT 85.930 334.600 86.330 335.200 ;
        RECT 85.930 334.400 89.930 334.600 ;
        RECT 85.930 333.800 86.330 334.400 ;
        RECT 85.930 333.600 89.930 333.800 ;
        RECT 85.930 333.000 86.330 333.600 ;
        RECT 85.930 332.800 89.930 333.000 ;
        RECT 85.930 332.200 86.330 332.800 ;
        RECT 85.930 332.000 89.930 332.200 ;
        RECT 85.930 331.400 86.330 332.000 ;
        RECT 85.930 331.200 89.930 331.400 ;
        RECT 85.930 330.600 86.330 331.200 ;
        RECT 85.930 330.400 89.930 330.600 ;
        RECT 85.930 330.200 86.330 330.400 ;
        RECT 90.680 330.200 90.880 337.800 ;
        RECT 91.480 330.200 91.680 337.800 ;
        RECT 92.280 330.200 92.480 337.800 ;
        RECT 93.080 330.200 93.280 337.800 ;
        RECT 93.880 330.200 94.080 337.800 ;
        RECT 85.930 329.800 94.080 330.200 ;
        RECT 85.930 329.600 86.330 329.800 ;
        RECT 85.930 329.400 89.930 329.600 ;
        RECT 85.930 328.800 86.330 329.400 ;
        RECT 85.930 328.600 89.930 328.800 ;
        RECT 85.930 328.000 86.330 328.600 ;
        RECT 85.930 327.800 89.930 328.000 ;
        RECT 85.930 327.200 86.330 327.800 ;
        RECT 85.930 327.000 89.930 327.200 ;
        RECT 85.930 326.400 86.330 327.000 ;
        RECT 85.930 326.200 89.930 326.400 ;
        RECT 85.930 325.600 86.330 326.200 ;
        RECT 85.930 325.400 89.930 325.600 ;
        RECT 85.930 324.800 86.330 325.400 ;
        RECT 85.930 324.600 89.930 324.800 ;
        RECT 85.930 324.000 86.330 324.600 ;
        RECT 85.930 323.800 89.930 324.000 ;
        RECT 85.930 323.200 86.330 323.800 ;
        RECT 85.930 323.000 89.930 323.200 ;
        RECT 85.930 322.400 86.330 323.000 ;
        RECT 85.930 322.200 89.930 322.400 ;
        RECT 90.680 322.200 90.880 329.800 ;
        RECT 91.480 322.200 91.680 329.800 ;
        RECT 92.280 322.200 92.480 329.800 ;
        RECT 93.080 322.200 93.280 329.800 ;
        RECT 93.880 322.200 94.080 329.800 ;
        RECT 95.380 330.200 95.580 337.800 ;
        RECT 96.180 330.200 96.380 337.800 ;
        RECT 96.980 330.200 97.180 337.800 ;
        RECT 97.780 330.200 97.980 337.800 ;
        RECT 98.580 330.200 98.780 337.800 ;
        RECT 99.530 337.600 103.530 337.800 ;
        RECT 103.130 337.000 103.530 337.600 ;
        RECT 99.530 336.800 103.530 337.000 ;
        RECT 103.130 336.200 103.530 336.800 ;
        RECT 99.530 336.000 103.530 336.200 ;
        RECT 103.130 335.400 103.530 336.000 ;
        RECT 99.530 335.200 103.530 335.400 ;
        RECT 103.130 334.600 103.530 335.200 ;
        RECT 99.530 334.400 103.530 334.600 ;
        RECT 103.130 333.800 103.530 334.400 ;
        RECT 99.530 333.600 103.530 333.800 ;
        RECT 103.130 333.000 103.530 333.600 ;
        RECT 99.530 332.800 103.530 333.000 ;
        RECT 103.130 332.200 103.530 332.800 ;
        RECT 99.530 332.000 103.530 332.200 ;
        RECT 103.130 331.400 103.530 332.000 ;
        RECT 99.530 331.200 103.530 331.400 ;
        RECT 103.130 330.600 103.530 331.200 ;
        RECT 99.530 330.400 103.530 330.600 ;
        RECT 103.130 330.200 103.530 330.400 ;
        RECT 95.380 329.800 103.530 330.200 ;
        RECT 110.050 329.910 110.410 330.290 ;
        RECT 110.680 329.910 111.040 330.290 ;
        RECT 111.280 329.910 111.640 330.290 ;
        RECT 95.380 322.200 95.580 329.800 ;
        RECT 96.180 322.200 96.380 329.800 ;
        RECT 96.980 322.200 97.180 329.800 ;
        RECT 97.780 322.200 97.980 329.800 ;
        RECT 98.580 322.200 98.780 329.800 ;
        RECT 103.130 329.600 103.530 329.800 ;
        RECT 99.530 329.400 103.530 329.600 ;
        RECT 103.130 328.800 103.530 329.400 ;
        RECT 110.050 329.320 110.410 329.700 ;
        RECT 110.680 329.320 111.040 329.700 ;
        RECT 111.280 329.320 111.640 329.700 ;
        RECT 99.530 328.600 103.530 328.800 ;
        RECT 103.130 328.000 103.530 328.600 ;
        RECT 99.530 327.800 103.530 328.000 ;
        RECT 103.130 327.200 103.530 327.800 ;
        RECT 99.530 327.000 103.530 327.200 ;
        RECT 103.130 326.400 103.530 327.000 ;
        RECT 99.530 326.200 103.530 326.400 ;
        RECT 103.130 325.600 103.530 326.200 ;
        RECT 99.530 325.400 103.530 325.600 ;
        RECT 103.130 324.800 103.530 325.400 ;
        RECT 99.530 324.600 103.530 324.800 ;
        RECT 103.130 324.000 103.530 324.600 ;
        RECT 99.530 323.800 103.530 324.000 ;
        RECT 103.130 323.200 103.530 323.800 ;
        RECT 99.530 323.000 103.530 323.200 ;
        RECT 103.130 322.400 103.530 323.000 ;
        RECT 99.530 322.200 103.530 322.400 ;
        RECT 5.930 317.600 9.930 317.800 ;
        RECT 5.930 317.000 6.330 317.600 ;
        RECT 5.930 316.800 9.930 317.000 ;
        RECT 5.930 316.200 6.330 316.800 ;
        RECT 5.930 316.000 9.930 316.200 ;
        RECT 5.930 315.400 6.330 316.000 ;
        RECT 5.930 315.200 9.930 315.400 ;
        RECT 5.930 314.600 6.330 315.200 ;
        RECT 5.930 314.400 9.930 314.600 ;
        RECT 5.930 313.800 6.330 314.400 ;
        RECT 5.930 313.600 9.930 313.800 ;
        RECT 5.930 313.000 6.330 313.600 ;
        RECT 5.930 312.800 9.930 313.000 ;
        RECT 5.930 312.200 6.330 312.800 ;
        RECT 5.930 312.000 9.930 312.200 ;
        RECT 5.930 311.400 6.330 312.000 ;
        RECT 5.930 311.200 9.930 311.400 ;
        RECT 5.930 310.600 6.330 311.200 ;
        RECT 5.930 310.400 9.930 310.600 ;
        RECT 5.930 310.200 6.330 310.400 ;
        RECT 10.680 310.200 10.880 317.800 ;
        RECT 11.480 310.200 11.680 317.800 ;
        RECT 12.280 310.200 12.480 317.800 ;
        RECT 13.080 310.200 13.280 317.800 ;
        RECT 13.880 310.200 14.080 317.800 ;
        RECT 5.930 309.800 14.080 310.200 ;
        RECT 5.930 309.600 6.330 309.800 ;
        RECT 5.930 309.400 9.930 309.600 ;
        RECT 5.930 308.800 6.330 309.400 ;
        RECT 5.930 308.600 9.930 308.800 ;
        RECT 5.930 308.000 6.330 308.600 ;
        RECT 5.930 307.800 9.930 308.000 ;
        RECT 5.930 307.200 6.330 307.800 ;
        RECT 5.930 307.000 9.930 307.200 ;
        RECT 5.930 306.400 6.330 307.000 ;
        RECT 5.930 306.200 9.930 306.400 ;
        RECT 5.930 305.600 6.330 306.200 ;
        RECT 5.930 305.400 9.930 305.600 ;
        RECT 5.930 304.800 6.330 305.400 ;
        RECT 5.930 304.600 9.930 304.800 ;
        RECT 5.930 304.000 6.330 304.600 ;
        RECT 5.930 303.800 9.930 304.000 ;
        RECT 5.930 303.200 6.330 303.800 ;
        RECT 5.930 303.000 9.930 303.200 ;
        RECT 5.930 302.400 6.330 303.000 ;
        RECT 5.930 302.200 9.930 302.400 ;
        RECT 10.680 302.200 10.880 309.800 ;
        RECT 11.480 302.200 11.680 309.800 ;
        RECT 12.280 302.200 12.480 309.800 ;
        RECT 13.080 302.200 13.280 309.800 ;
        RECT 13.880 302.200 14.080 309.800 ;
        RECT 15.380 310.200 15.580 317.800 ;
        RECT 16.180 310.200 16.380 317.800 ;
        RECT 16.980 310.200 17.180 317.800 ;
        RECT 17.780 310.200 17.980 317.800 ;
        RECT 18.580 310.200 18.780 317.800 ;
        RECT 19.530 317.600 23.530 317.800 ;
        RECT 23.130 317.000 23.530 317.600 ;
        RECT 19.530 316.800 23.530 317.000 ;
        RECT 23.130 316.200 23.530 316.800 ;
        RECT 19.530 316.000 23.530 316.200 ;
        RECT 23.130 315.400 23.530 316.000 ;
        RECT 19.530 315.200 23.530 315.400 ;
        RECT 23.130 314.600 23.530 315.200 ;
        RECT 19.530 314.400 23.530 314.600 ;
        RECT 23.130 313.800 23.530 314.400 ;
        RECT 19.530 313.600 23.530 313.800 ;
        RECT 23.130 313.000 23.530 313.600 ;
        RECT 19.530 312.800 23.530 313.000 ;
        RECT 23.130 312.200 23.530 312.800 ;
        RECT 19.530 312.000 23.530 312.200 ;
        RECT 23.130 311.400 23.530 312.000 ;
        RECT 19.530 311.200 23.530 311.400 ;
        RECT 23.130 310.600 23.530 311.200 ;
        RECT 19.530 310.400 23.530 310.600 ;
        RECT 23.130 310.200 23.530 310.400 ;
        RECT 15.380 309.800 23.530 310.200 ;
        RECT 15.380 302.200 15.580 309.800 ;
        RECT 16.180 302.200 16.380 309.800 ;
        RECT 16.980 302.200 17.180 309.800 ;
        RECT 17.780 302.200 17.980 309.800 ;
        RECT 18.580 302.200 18.780 309.800 ;
        RECT 23.130 309.600 23.530 309.800 ;
        RECT 19.530 309.400 23.530 309.600 ;
        RECT 23.130 308.800 23.530 309.400 ;
        RECT 19.530 308.600 23.530 308.800 ;
        RECT 23.130 308.000 23.530 308.600 ;
        RECT 19.530 307.800 23.530 308.000 ;
        RECT 23.130 307.200 23.530 307.800 ;
        RECT 19.530 307.000 23.530 307.200 ;
        RECT 23.130 306.400 23.530 307.000 ;
        RECT 19.530 306.200 23.530 306.400 ;
        RECT 23.130 305.600 23.530 306.200 ;
        RECT 19.530 305.400 23.530 305.600 ;
        RECT 23.130 304.800 23.530 305.400 ;
        RECT 19.530 304.600 23.530 304.800 ;
        RECT 23.130 304.000 23.530 304.600 ;
        RECT 19.530 303.800 23.530 304.000 ;
        RECT 23.130 303.200 23.530 303.800 ;
        RECT 19.530 303.000 23.530 303.200 ;
        RECT 23.130 302.400 23.530 303.000 ;
        RECT 19.530 302.200 23.530 302.400 ;
        RECT 25.930 317.600 29.930 317.800 ;
        RECT 25.930 317.000 26.330 317.600 ;
        RECT 25.930 316.800 29.930 317.000 ;
        RECT 25.930 316.200 26.330 316.800 ;
        RECT 25.930 316.000 29.930 316.200 ;
        RECT 25.930 315.400 26.330 316.000 ;
        RECT 25.930 315.200 29.930 315.400 ;
        RECT 25.930 314.600 26.330 315.200 ;
        RECT 25.930 314.400 29.930 314.600 ;
        RECT 25.930 313.800 26.330 314.400 ;
        RECT 25.930 313.600 29.930 313.800 ;
        RECT 25.930 313.000 26.330 313.600 ;
        RECT 25.930 312.800 29.930 313.000 ;
        RECT 25.930 312.200 26.330 312.800 ;
        RECT 25.930 312.000 29.930 312.200 ;
        RECT 25.930 311.400 26.330 312.000 ;
        RECT 25.930 311.200 29.930 311.400 ;
        RECT 25.930 310.600 26.330 311.200 ;
        RECT 25.930 310.400 29.930 310.600 ;
        RECT 25.930 310.200 26.330 310.400 ;
        RECT 30.680 310.200 30.880 317.800 ;
        RECT 31.480 310.200 31.680 317.800 ;
        RECT 32.280 310.200 32.480 317.800 ;
        RECT 33.080 310.200 33.280 317.800 ;
        RECT 33.880 310.200 34.080 317.800 ;
        RECT 25.930 309.800 34.080 310.200 ;
        RECT 25.930 309.600 26.330 309.800 ;
        RECT 25.930 309.400 29.930 309.600 ;
        RECT 25.930 308.800 26.330 309.400 ;
        RECT 25.930 308.600 29.930 308.800 ;
        RECT 25.930 308.000 26.330 308.600 ;
        RECT 25.930 307.800 29.930 308.000 ;
        RECT 25.930 307.200 26.330 307.800 ;
        RECT 25.930 307.000 29.930 307.200 ;
        RECT 25.930 306.400 26.330 307.000 ;
        RECT 25.930 306.200 29.930 306.400 ;
        RECT 25.930 305.600 26.330 306.200 ;
        RECT 25.930 305.400 29.930 305.600 ;
        RECT 25.930 304.800 26.330 305.400 ;
        RECT 25.930 304.600 29.930 304.800 ;
        RECT 25.930 304.000 26.330 304.600 ;
        RECT 25.930 303.800 29.930 304.000 ;
        RECT 25.930 303.200 26.330 303.800 ;
        RECT 25.930 303.000 29.930 303.200 ;
        RECT 25.930 302.400 26.330 303.000 ;
        RECT 25.930 302.200 29.930 302.400 ;
        RECT 30.680 302.200 30.880 309.800 ;
        RECT 31.480 302.200 31.680 309.800 ;
        RECT 32.280 302.200 32.480 309.800 ;
        RECT 33.080 302.200 33.280 309.800 ;
        RECT 33.880 302.200 34.080 309.800 ;
        RECT 35.380 310.200 35.580 317.800 ;
        RECT 36.180 310.200 36.380 317.800 ;
        RECT 36.980 310.200 37.180 317.800 ;
        RECT 37.780 310.200 37.980 317.800 ;
        RECT 38.580 310.200 38.780 317.800 ;
        RECT 39.530 317.600 43.530 317.800 ;
        RECT 43.130 317.000 43.530 317.600 ;
        RECT 39.530 316.800 43.530 317.000 ;
        RECT 43.130 316.200 43.530 316.800 ;
        RECT 39.530 316.000 43.530 316.200 ;
        RECT 43.130 315.400 43.530 316.000 ;
        RECT 39.530 315.200 43.530 315.400 ;
        RECT 43.130 314.600 43.530 315.200 ;
        RECT 39.530 314.400 43.530 314.600 ;
        RECT 43.130 313.800 43.530 314.400 ;
        RECT 39.530 313.600 43.530 313.800 ;
        RECT 43.130 313.000 43.530 313.600 ;
        RECT 39.530 312.800 43.530 313.000 ;
        RECT 43.130 312.200 43.530 312.800 ;
        RECT 39.530 312.000 43.530 312.200 ;
        RECT 43.130 311.400 43.530 312.000 ;
        RECT 39.530 311.200 43.530 311.400 ;
        RECT 43.130 310.600 43.530 311.200 ;
        RECT 39.530 310.400 43.530 310.600 ;
        RECT 43.130 310.200 43.530 310.400 ;
        RECT 35.380 309.800 43.530 310.200 ;
        RECT 35.380 302.200 35.580 309.800 ;
        RECT 36.180 302.200 36.380 309.800 ;
        RECT 36.980 302.200 37.180 309.800 ;
        RECT 37.780 302.200 37.980 309.800 ;
        RECT 38.580 302.200 38.780 309.800 ;
        RECT 43.130 309.600 43.530 309.800 ;
        RECT 39.530 309.400 43.530 309.600 ;
        RECT 43.130 308.800 43.530 309.400 ;
        RECT 39.530 308.600 43.530 308.800 ;
        RECT 43.130 308.000 43.530 308.600 ;
        RECT 39.530 307.800 43.530 308.000 ;
        RECT 43.130 307.200 43.530 307.800 ;
        RECT 39.530 307.000 43.530 307.200 ;
        RECT 43.130 306.400 43.530 307.000 ;
        RECT 39.530 306.200 43.530 306.400 ;
        RECT 43.130 305.600 43.530 306.200 ;
        RECT 39.530 305.400 43.530 305.600 ;
        RECT 43.130 304.800 43.530 305.400 ;
        RECT 39.530 304.600 43.530 304.800 ;
        RECT 43.130 304.000 43.530 304.600 ;
        RECT 39.530 303.800 43.530 304.000 ;
        RECT 43.130 303.200 43.530 303.800 ;
        RECT 39.530 303.000 43.530 303.200 ;
        RECT 43.130 302.400 43.530 303.000 ;
        RECT 39.530 302.200 43.530 302.400 ;
        RECT 45.930 317.600 49.930 317.800 ;
        RECT 45.930 317.000 46.330 317.600 ;
        RECT 45.930 316.800 49.930 317.000 ;
        RECT 45.930 316.200 46.330 316.800 ;
        RECT 45.930 316.000 49.930 316.200 ;
        RECT 45.930 315.400 46.330 316.000 ;
        RECT 45.930 315.200 49.930 315.400 ;
        RECT 45.930 314.600 46.330 315.200 ;
        RECT 45.930 314.400 49.930 314.600 ;
        RECT 45.930 313.800 46.330 314.400 ;
        RECT 45.930 313.600 49.930 313.800 ;
        RECT 45.930 313.000 46.330 313.600 ;
        RECT 45.930 312.800 49.930 313.000 ;
        RECT 45.930 312.200 46.330 312.800 ;
        RECT 45.930 312.000 49.930 312.200 ;
        RECT 45.930 311.400 46.330 312.000 ;
        RECT 45.930 311.200 49.930 311.400 ;
        RECT 45.930 310.600 46.330 311.200 ;
        RECT 45.930 310.400 49.930 310.600 ;
        RECT 45.930 310.200 46.330 310.400 ;
        RECT 50.680 310.200 50.880 317.800 ;
        RECT 51.480 310.200 51.680 317.800 ;
        RECT 52.280 310.200 52.480 317.800 ;
        RECT 53.080 310.200 53.280 317.800 ;
        RECT 53.880 310.200 54.080 317.800 ;
        RECT 45.930 309.800 54.080 310.200 ;
        RECT 45.930 309.600 46.330 309.800 ;
        RECT 45.930 309.400 49.930 309.600 ;
        RECT 45.930 308.800 46.330 309.400 ;
        RECT 45.930 308.600 49.930 308.800 ;
        RECT 45.930 308.000 46.330 308.600 ;
        RECT 45.930 307.800 49.930 308.000 ;
        RECT 45.930 307.200 46.330 307.800 ;
        RECT 45.930 307.000 49.930 307.200 ;
        RECT 45.930 306.400 46.330 307.000 ;
        RECT 45.930 306.200 49.930 306.400 ;
        RECT 45.930 305.600 46.330 306.200 ;
        RECT 45.930 305.400 49.930 305.600 ;
        RECT 45.930 304.800 46.330 305.400 ;
        RECT 45.930 304.600 49.930 304.800 ;
        RECT 45.930 304.000 46.330 304.600 ;
        RECT 45.930 303.800 49.930 304.000 ;
        RECT 45.930 303.200 46.330 303.800 ;
        RECT 45.930 303.000 49.930 303.200 ;
        RECT 45.930 302.400 46.330 303.000 ;
        RECT 45.930 302.200 49.930 302.400 ;
        RECT 50.680 302.200 50.880 309.800 ;
        RECT 51.480 302.200 51.680 309.800 ;
        RECT 52.280 302.200 52.480 309.800 ;
        RECT 53.080 302.200 53.280 309.800 ;
        RECT 53.880 302.200 54.080 309.800 ;
        RECT 55.380 310.200 55.580 317.800 ;
        RECT 56.180 310.200 56.380 317.800 ;
        RECT 56.980 310.200 57.180 317.800 ;
        RECT 57.780 310.200 57.980 317.800 ;
        RECT 58.580 310.200 58.780 317.800 ;
        RECT 59.530 317.600 63.530 317.800 ;
        RECT 63.130 317.000 63.530 317.600 ;
        RECT 59.530 316.800 63.530 317.000 ;
        RECT 63.130 316.200 63.530 316.800 ;
        RECT 59.530 316.000 63.530 316.200 ;
        RECT 63.130 315.400 63.530 316.000 ;
        RECT 59.530 315.200 63.530 315.400 ;
        RECT 63.130 314.600 63.530 315.200 ;
        RECT 59.530 314.400 63.530 314.600 ;
        RECT 63.130 313.800 63.530 314.400 ;
        RECT 59.530 313.600 63.530 313.800 ;
        RECT 63.130 313.000 63.530 313.600 ;
        RECT 59.530 312.800 63.530 313.000 ;
        RECT 63.130 312.200 63.530 312.800 ;
        RECT 59.530 312.000 63.530 312.200 ;
        RECT 63.130 311.400 63.530 312.000 ;
        RECT 59.530 311.200 63.530 311.400 ;
        RECT 63.130 310.600 63.530 311.200 ;
        RECT 59.530 310.400 63.530 310.600 ;
        RECT 63.130 310.200 63.530 310.400 ;
        RECT 55.380 309.800 63.530 310.200 ;
        RECT 55.380 302.200 55.580 309.800 ;
        RECT 56.180 302.200 56.380 309.800 ;
        RECT 56.980 302.200 57.180 309.800 ;
        RECT 57.780 302.200 57.980 309.800 ;
        RECT 58.580 302.200 58.780 309.800 ;
        RECT 63.130 309.600 63.530 309.800 ;
        RECT 59.530 309.400 63.530 309.600 ;
        RECT 63.130 308.800 63.530 309.400 ;
        RECT 59.530 308.600 63.530 308.800 ;
        RECT 63.130 308.000 63.530 308.600 ;
        RECT 59.530 307.800 63.530 308.000 ;
        RECT 63.130 307.200 63.530 307.800 ;
        RECT 59.530 307.000 63.530 307.200 ;
        RECT 63.130 306.400 63.530 307.000 ;
        RECT 59.530 306.200 63.530 306.400 ;
        RECT 63.130 305.600 63.530 306.200 ;
        RECT 59.530 305.400 63.530 305.600 ;
        RECT 63.130 304.800 63.530 305.400 ;
        RECT 59.530 304.600 63.530 304.800 ;
        RECT 63.130 304.000 63.530 304.600 ;
        RECT 59.530 303.800 63.530 304.000 ;
        RECT 63.130 303.200 63.530 303.800 ;
        RECT 59.530 303.000 63.530 303.200 ;
        RECT 63.130 302.400 63.530 303.000 ;
        RECT 59.530 302.200 63.530 302.400 ;
        RECT 65.930 317.600 69.930 317.800 ;
        RECT 65.930 317.000 66.330 317.600 ;
        RECT 65.930 316.800 69.930 317.000 ;
        RECT 65.930 316.200 66.330 316.800 ;
        RECT 65.930 316.000 69.930 316.200 ;
        RECT 65.930 315.400 66.330 316.000 ;
        RECT 65.930 315.200 69.930 315.400 ;
        RECT 65.930 314.600 66.330 315.200 ;
        RECT 65.930 314.400 69.930 314.600 ;
        RECT 65.930 313.800 66.330 314.400 ;
        RECT 65.930 313.600 69.930 313.800 ;
        RECT 65.930 313.000 66.330 313.600 ;
        RECT 65.930 312.800 69.930 313.000 ;
        RECT 65.930 312.200 66.330 312.800 ;
        RECT 65.930 312.000 69.930 312.200 ;
        RECT 65.930 311.400 66.330 312.000 ;
        RECT 65.930 311.200 69.930 311.400 ;
        RECT 65.930 310.600 66.330 311.200 ;
        RECT 65.930 310.400 69.930 310.600 ;
        RECT 65.930 310.200 66.330 310.400 ;
        RECT 70.680 310.200 70.880 317.800 ;
        RECT 71.480 310.200 71.680 317.800 ;
        RECT 72.280 310.200 72.480 317.800 ;
        RECT 73.080 310.200 73.280 317.800 ;
        RECT 73.880 310.200 74.080 317.800 ;
        RECT 65.930 309.800 74.080 310.200 ;
        RECT 65.930 309.600 66.330 309.800 ;
        RECT 65.930 309.400 69.930 309.600 ;
        RECT 65.930 308.800 66.330 309.400 ;
        RECT 65.930 308.600 69.930 308.800 ;
        RECT 65.930 308.000 66.330 308.600 ;
        RECT 65.930 307.800 69.930 308.000 ;
        RECT 65.930 307.200 66.330 307.800 ;
        RECT 65.930 307.000 69.930 307.200 ;
        RECT 65.930 306.400 66.330 307.000 ;
        RECT 65.930 306.200 69.930 306.400 ;
        RECT 65.930 305.600 66.330 306.200 ;
        RECT 65.930 305.400 69.930 305.600 ;
        RECT 65.930 304.800 66.330 305.400 ;
        RECT 65.930 304.600 69.930 304.800 ;
        RECT 65.930 304.000 66.330 304.600 ;
        RECT 65.930 303.800 69.930 304.000 ;
        RECT 65.930 303.200 66.330 303.800 ;
        RECT 65.930 303.000 69.930 303.200 ;
        RECT 65.930 302.400 66.330 303.000 ;
        RECT 65.930 302.200 69.930 302.400 ;
        RECT 70.680 302.200 70.880 309.800 ;
        RECT 71.480 302.200 71.680 309.800 ;
        RECT 72.280 302.200 72.480 309.800 ;
        RECT 73.080 302.200 73.280 309.800 ;
        RECT 73.880 302.200 74.080 309.800 ;
        RECT 75.380 310.200 75.580 317.800 ;
        RECT 76.180 310.200 76.380 317.800 ;
        RECT 76.980 310.200 77.180 317.800 ;
        RECT 77.780 310.200 77.980 317.800 ;
        RECT 78.580 310.200 78.780 317.800 ;
        RECT 79.530 317.600 83.530 317.800 ;
        RECT 83.130 317.000 83.530 317.600 ;
        RECT 79.530 316.800 83.530 317.000 ;
        RECT 83.130 316.200 83.530 316.800 ;
        RECT 79.530 316.000 83.530 316.200 ;
        RECT 83.130 315.400 83.530 316.000 ;
        RECT 79.530 315.200 83.530 315.400 ;
        RECT 83.130 314.600 83.530 315.200 ;
        RECT 79.530 314.400 83.530 314.600 ;
        RECT 83.130 313.800 83.530 314.400 ;
        RECT 79.530 313.600 83.530 313.800 ;
        RECT 83.130 313.000 83.530 313.600 ;
        RECT 79.530 312.800 83.530 313.000 ;
        RECT 83.130 312.200 83.530 312.800 ;
        RECT 79.530 312.000 83.530 312.200 ;
        RECT 83.130 311.400 83.530 312.000 ;
        RECT 79.530 311.200 83.530 311.400 ;
        RECT 83.130 310.600 83.530 311.200 ;
        RECT 79.530 310.400 83.530 310.600 ;
        RECT 83.130 310.200 83.530 310.400 ;
        RECT 75.380 309.800 83.530 310.200 ;
        RECT 75.380 302.200 75.580 309.800 ;
        RECT 76.180 302.200 76.380 309.800 ;
        RECT 76.980 302.200 77.180 309.800 ;
        RECT 77.780 302.200 77.980 309.800 ;
        RECT 78.580 302.200 78.780 309.800 ;
        RECT 83.130 309.600 83.530 309.800 ;
        RECT 79.530 309.400 83.530 309.600 ;
        RECT 83.130 308.800 83.530 309.400 ;
        RECT 79.530 308.600 83.530 308.800 ;
        RECT 83.130 308.000 83.530 308.600 ;
        RECT 79.530 307.800 83.530 308.000 ;
        RECT 83.130 307.200 83.530 307.800 ;
        RECT 79.530 307.000 83.530 307.200 ;
        RECT 83.130 306.400 83.530 307.000 ;
        RECT 79.530 306.200 83.530 306.400 ;
        RECT 83.130 305.600 83.530 306.200 ;
        RECT 79.530 305.400 83.530 305.600 ;
        RECT 83.130 304.800 83.530 305.400 ;
        RECT 79.530 304.600 83.530 304.800 ;
        RECT 83.130 304.000 83.530 304.600 ;
        RECT 79.530 303.800 83.530 304.000 ;
        RECT 83.130 303.200 83.530 303.800 ;
        RECT 79.530 303.000 83.530 303.200 ;
        RECT 83.130 302.400 83.530 303.000 ;
        RECT 79.530 302.200 83.530 302.400 ;
        RECT 85.930 317.600 89.930 317.800 ;
        RECT 85.930 317.000 86.330 317.600 ;
        RECT 85.930 316.800 89.930 317.000 ;
        RECT 85.930 316.200 86.330 316.800 ;
        RECT 85.930 316.000 89.930 316.200 ;
        RECT 85.930 315.400 86.330 316.000 ;
        RECT 85.930 315.200 89.930 315.400 ;
        RECT 85.930 314.600 86.330 315.200 ;
        RECT 85.930 314.400 89.930 314.600 ;
        RECT 85.930 313.800 86.330 314.400 ;
        RECT 85.930 313.600 89.930 313.800 ;
        RECT 85.930 313.000 86.330 313.600 ;
        RECT 85.930 312.800 89.930 313.000 ;
        RECT 85.930 312.200 86.330 312.800 ;
        RECT 85.930 312.000 89.930 312.200 ;
        RECT 85.930 311.400 86.330 312.000 ;
        RECT 85.930 311.200 89.930 311.400 ;
        RECT 85.930 310.600 86.330 311.200 ;
        RECT 85.930 310.400 89.930 310.600 ;
        RECT 85.930 310.200 86.330 310.400 ;
        RECT 90.680 310.200 90.880 317.800 ;
        RECT 91.480 310.200 91.680 317.800 ;
        RECT 92.280 310.200 92.480 317.800 ;
        RECT 93.080 310.200 93.280 317.800 ;
        RECT 93.880 310.200 94.080 317.800 ;
        RECT 85.930 309.800 94.080 310.200 ;
        RECT 85.930 309.600 86.330 309.800 ;
        RECT 85.930 309.400 89.930 309.600 ;
        RECT 85.930 308.800 86.330 309.400 ;
        RECT 85.930 308.600 89.930 308.800 ;
        RECT 85.930 308.000 86.330 308.600 ;
        RECT 85.930 307.800 89.930 308.000 ;
        RECT 85.930 307.200 86.330 307.800 ;
        RECT 85.930 307.000 89.930 307.200 ;
        RECT 85.930 306.400 86.330 307.000 ;
        RECT 85.930 306.200 89.930 306.400 ;
        RECT 85.930 305.600 86.330 306.200 ;
        RECT 85.930 305.400 89.930 305.600 ;
        RECT 85.930 304.800 86.330 305.400 ;
        RECT 85.930 304.600 89.930 304.800 ;
        RECT 85.930 304.000 86.330 304.600 ;
        RECT 85.930 303.800 89.930 304.000 ;
        RECT 85.930 303.200 86.330 303.800 ;
        RECT 85.930 303.000 89.930 303.200 ;
        RECT 85.930 302.400 86.330 303.000 ;
        RECT 85.930 302.200 89.930 302.400 ;
        RECT 90.680 302.200 90.880 309.800 ;
        RECT 91.480 302.200 91.680 309.800 ;
        RECT 92.280 302.200 92.480 309.800 ;
        RECT 93.080 302.200 93.280 309.800 ;
        RECT 93.880 302.200 94.080 309.800 ;
        RECT 95.380 310.200 95.580 317.800 ;
        RECT 96.180 310.200 96.380 317.800 ;
        RECT 96.980 310.200 97.180 317.800 ;
        RECT 97.780 310.200 97.980 317.800 ;
        RECT 98.580 310.200 98.780 317.800 ;
        RECT 99.530 317.600 103.530 317.800 ;
        RECT 103.130 317.000 103.530 317.600 ;
        RECT 99.530 316.800 103.530 317.000 ;
        RECT 103.130 316.200 103.530 316.800 ;
        RECT 99.530 316.000 103.530 316.200 ;
        RECT 103.130 315.400 103.530 316.000 ;
        RECT 99.530 315.200 103.530 315.400 ;
        RECT 103.130 314.600 103.530 315.200 ;
        RECT 99.530 314.400 103.530 314.600 ;
        RECT 103.130 313.800 103.530 314.400 ;
        RECT 99.530 313.600 103.530 313.800 ;
        RECT 103.130 313.000 103.530 313.600 ;
        RECT 99.530 312.800 103.530 313.000 ;
        RECT 103.130 312.200 103.530 312.800 ;
        RECT 99.530 312.000 103.530 312.200 ;
        RECT 103.130 311.400 103.530 312.000 ;
        RECT 99.530 311.200 103.530 311.400 ;
        RECT 103.130 310.600 103.530 311.200 ;
        RECT 99.530 310.400 103.530 310.600 ;
        RECT 103.130 310.200 103.530 310.400 ;
        RECT 95.380 309.800 103.530 310.200 ;
        RECT 110.050 309.905 110.410 310.285 ;
        RECT 110.680 309.905 111.040 310.285 ;
        RECT 111.280 309.905 111.640 310.285 ;
        RECT 95.380 302.200 95.580 309.800 ;
        RECT 96.180 302.200 96.380 309.800 ;
        RECT 96.980 302.200 97.180 309.800 ;
        RECT 97.780 302.200 97.980 309.800 ;
        RECT 98.580 302.200 98.780 309.800 ;
        RECT 103.130 309.600 103.530 309.800 ;
        RECT 99.530 309.400 103.530 309.600 ;
        RECT 103.130 308.800 103.530 309.400 ;
        RECT 110.050 309.315 110.410 309.695 ;
        RECT 110.680 309.315 111.040 309.695 ;
        RECT 111.280 309.315 111.640 309.695 ;
        RECT 99.530 308.600 103.530 308.800 ;
        RECT 103.130 308.000 103.530 308.600 ;
        RECT 99.530 307.800 103.530 308.000 ;
        RECT 103.130 307.200 103.530 307.800 ;
        RECT 99.530 307.000 103.530 307.200 ;
        RECT 103.130 306.400 103.530 307.000 ;
        RECT 99.530 306.200 103.530 306.400 ;
        RECT 103.130 305.600 103.530 306.200 ;
        RECT 99.530 305.400 103.530 305.600 ;
        RECT 103.130 304.800 103.530 305.400 ;
        RECT 99.530 304.600 103.530 304.800 ;
        RECT 103.130 304.000 103.530 304.600 ;
        RECT 99.530 303.800 103.530 304.000 ;
        RECT 103.130 303.200 103.530 303.800 ;
        RECT 99.530 303.000 103.530 303.200 ;
        RECT 103.130 302.400 103.530 303.000 ;
        RECT 99.530 302.200 103.530 302.400 ;
        RECT 5.930 297.600 9.930 297.800 ;
        RECT 5.930 297.000 6.330 297.600 ;
        RECT 5.930 296.800 9.930 297.000 ;
        RECT 5.930 296.200 6.330 296.800 ;
        RECT 5.930 296.000 9.930 296.200 ;
        RECT 5.930 295.400 6.330 296.000 ;
        RECT 5.930 295.200 9.930 295.400 ;
        RECT 5.930 294.600 6.330 295.200 ;
        RECT 5.930 294.400 9.930 294.600 ;
        RECT 5.930 293.800 6.330 294.400 ;
        RECT 5.930 293.600 9.930 293.800 ;
        RECT 5.930 293.000 6.330 293.600 ;
        RECT 5.930 292.800 9.930 293.000 ;
        RECT 5.930 292.200 6.330 292.800 ;
        RECT 5.930 292.000 9.930 292.200 ;
        RECT 5.930 291.400 6.330 292.000 ;
        RECT 5.930 291.200 9.930 291.400 ;
        RECT 5.930 290.600 6.330 291.200 ;
        RECT 5.930 290.400 9.930 290.600 ;
        RECT 5.930 290.200 6.330 290.400 ;
        RECT 10.680 290.200 10.880 297.800 ;
        RECT 11.480 290.200 11.680 297.800 ;
        RECT 12.280 290.200 12.480 297.800 ;
        RECT 13.080 290.200 13.280 297.800 ;
        RECT 13.880 290.200 14.080 297.800 ;
        RECT 5.930 289.800 14.080 290.200 ;
        RECT 5.930 289.600 6.330 289.800 ;
        RECT 5.930 289.400 9.930 289.600 ;
        RECT 5.930 288.800 6.330 289.400 ;
        RECT 5.930 288.600 9.930 288.800 ;
        RECT 5.930 288.000 6.330 288.600 ;
        RECT 5.930 287.800 9.930 288.000 ;
        RECT 5.930 287.200 6.330 287.800 ;
        RECT 5.930 287.000 9.930 287.200 ;
        RECT 5.930 286.400 6.330 287.000 ;
        RECT 5.930 286.200 9.930 286.400 ;
        RECT 5.930 285.600 6.330 286.200 ;
        RECT 5.930 285.400 9.930 285.600 ;
        RECT 5.930 284.800 6.330 285.400 ;
        RECT 5.930 284.600 9.930 284.800 ;
        RECT 5.930 284.000 6.330 284.600 ;
        RECT 5.930 283.800 9.930 284.000 ;
        RECT 5.930 283.200 6.330 283.800 ;
        RECT 5.930 283.000 9.930 283.200 ;
        RECT 5.930 282.400 6.330 283.000 ;
        RECT 5.930 282.200 9.930 282.400 ;
        RECT 10.680 282.200 10.880 289.800 ;
        RECT 11.480 282.200 11.680 289.800 ;
        RECT 12.280 282.200 12.480 289.800 ;
        RECT 13.080 282.200 13.280 289.800 ;
        RECT 13.880 282.200 14.080 289.800 ;
        RECT 15.380 290.200 15.580 297.800 ;
        RECT 16.180 290.200 16.380 297.800 ;
        RECT 16.980 290.200 17.180 297.800 ;
        RECT 17.780 290.200 17.980 297.800 ;
        RECT 18.580 290.200 18.780 297.800 ;
        RECT 19.530 297.600 23.530 297.800 ;
        RECT 23.130 297.000 23.530 297.600 ;
        RECT 19.530 296.800 23.530 297.000 ;
        RECT 23.130 296.200 23.530 296.800 ;
        RECT 19.530 296.000 23.530 296.200 ;
        RECT 23.130 295.400 23.530 296.000 ;
        RECT 19.530 295.200 23.530 295.400 ;
        RECT 23.130 294.600 23.530 295.200 ;
        RECT 19.530 294.400 23.530 294.600 ;
        RECT 23.130 293.800 23.530 294.400 ;
        RECT 19.530 293.600 23.530 293.800 ;
        RECT 23.130 293.000 23.530 293.600 ;
        RECT 19.530 292.800 23.530 293.000 ;
        RECT 23.130 292.200 23.530 292.800 ;
        RECT 19.530 292.000 23.530 292.200 ;
        RECT 23.130 291.400 23.530 292.000 ;
        RECT 19.530 291.200 23.530 291.400 ;
        RECT 23.130 290.600 23.530 291.200 ;
        RECT 19.530 290.400 23.530 290.600 ;
        RECT 23.130 290.200 23.530 290.400 ;
        RECT 15.380 289.800 23.530 290.200 ;
        RECT 15.380 282.200 15.580 289.800 ;
        RECT 16.180 282.200 16.380 289.800 ;
        RECT 16.980 282.200 17.180 289.800 ;
        RECT 17.780 282.200 17.980 289.800 ;
        RECT 18.580 282.200 18.780 289.800 ;
        RECT 23.130 289.600 23.530 289.800 ;
        RECT 19.530 289.400 23.530 289.600 ;
        RECT 23.130 288.800 23.530 289.400 ;
        RECT 19.530 288.600 23.530 288.800 ;
        RECT 23.130 288.000 23.530 288.600 ;
        RECT 19.530 287.800 23.530 288.000 ;
        RECT 23.130 287.200 23.530 287.800 ;
        RECT 19.530 287.000 23.530 287.200 ;
        RECT 23.130 286.400 23.530 287.000 ;
        RECT 19.530 286.200 23.530 286.400 ;
        RECT 23.130 285.600 23.530 286.200 ;
        RECT 19.530 285.400 23.530 285.600 ;
        RECT 23.130 284.800 23.530 285.400 ;
        RECT 19.530 284.600 23.530 284.800 ;
        RECT 23.130 284.000 23.530 284.600 ;
        RECT 19.530 283.800 23.530 284.000 ;
        RECT 23.130 283.200 23.530 283.800 ;
        RECT 19.530 283.000 23.530 283.200 ;
        RECT 23.130 282.400 23.530 283.000 ;
        RECT 19.530 282.200 23.530 282.400 ;
        RECT 25.930 297.600 29.930 297.800 ;
        RECT 25.930 297.000 26.330 297.600 ;
        RECT 25.930 296.800 29.930 297.000 ;
        RECT 25.930 296.200 26.330 296.800 ;
        RECT 25.930 296.000 29.930 296.200 ;
        RECT 25.930 295.400 26.330 296.000 ;
        RECT 25.930 295.200 29.930 295.400 ;
        RECT 25.930 294.600 26.330 295.200 ;
        RECT 25.930 294.400 29.930 294.600 ;
        RECT 25.930 293.800 26.330 294.400 ;
        RECT 25.930 293.600 29.930 293.800 ;
        RECT 25.930 293.000 26.330 293.600 ;
        RECT 25.930 292.800 29.930 293.000 ;
        RECT 25.930 292.200 26.330 292.800 ;
        RECT 25.930 292.000 29.930 292.200 ;
        RECT 25.930 291.400 26.330 292.000 ;
        RECT 25.930 291.200 29.930 291.400 ;
        RECT 25.930 290.600 26.330 291.200 ;
        RECT 25.930 290.400 29.930 290.600 ;
        RECT 25.930 290.200 26.330 290.400 ;
        RECT 30.680 290.200 30.880 297.800 ;
        RECT 31.480 290.200 31.680 297.800 ;
        RECT 32.280 290.200 32.480 297.800 ;
        RECT 33.080 290.200 33.280 297.800 ;
        RECT 33.880 290.200 34.080 297.800 ;
        RECT 25.930 289.800 34.080 290.200 ;
        RECT 25.930 289.600 26.330 289.800 ;
        RECT 25.930 289.400 29.930 289.600 ;
        RECT 25.930 288.800 26.330 289.400 ;
        RECT 25.930 288.600 29.930 288.800 ;
        RECT 25.930 288.000 26.330 288.600 ;
        RECT 25.930 287.800 29.930 288.000 ;
        RECT 25.930 287.200 26.330 287.800 ;
        RECT 25.930 287.000 29.930 287.200 ;
        RECT 25.930 286.400 26.330 287.000 ;
        RECT 25.930 286.200 29.930 286.400 ;
        RECT 25.930 285.600 26.330 286.200 ;
        RECT 25.930 285.400 29.930 285.600 ;
        RECT 25.930 284.800 26.330 285.400 ;
        RECT 25.930 284.600 29.930 284.800 ;
        RECT 25.930 284.000 26.330 284.600 ;
        RECT 25.930 283.800 29.930 284.000 ;
        RECT 25.930 283.200 26.330 283.800 ;
        RECT 25.930 283.000 29.930 283.200 ;
        RECT 25.930 282.400 26.330 283.000 ;
        RECT 25.930 282.200 29.930 282.400 ;
        RECT 30.680 282.200 30.880 289.800 ;
        RECT 31.480 282.200 31.680 289.800 ;
        RECT 32.280 282.200 32.480 289.800 ;
        RECT 33.080 282.200 33.280 289.800 ;
        RECT 33.880 282.200 34.080 289.800 ;
        RECT 35.380 290.200 35.580 297.800 ;
        RECT 36.180 290.200 36.380 297.800 ;
        RECT 36.980 290.200 37.180 297.800 ;
        RECT 37.780 290.200 37.980 297.800 ;
        RECT 38.580 290.200 38.780 297.800 ;
        RECT 39.530 297.600 43.530 297.800 ;
        RECT 43.130 297.000 43.530 297.600 ;
        RECT 39.530 296.800 43.530 297.000 ;
        RECT 43.130 296.200 43.530 296.800 ;
        RECT 39.530 296.000 43.530 296.200 ;
        RECT 43.130 295.400 43.530 296.000 ;
        RECT 39.530 295.200 43.530 295.400 ;
        RECT 43.130 294.600 43.530 295.200 ;
        RECT 39.530 294.400 43.530 294.600 ;
        RECT 43.130 293.800 43.530 294.400 ;
        RECT 39.530 293.600 43.530 293.800 ;
        RECT 43.130 293.000 43.530 293.600 ;
        RECT 39.530 292.800 43.530 293.000 ;
        RECT 43.130 292.200 43.530 292.800 ;
        RECT 39.530 292.000 43.530 292.200 ;
        RECT 43.130 291.400 43.530 292.000 ;
        RECT 39.530 291.200 43.530 291.400 ;
        RECT 43.130 290.600 43.530 291.200 ;
        RECT 39.530 290.400 43.530 290.600 ;
        RECT 43.130 290.200 43.530 290.400 ;
        RECT 35.380 289.800 43.530 290.200 ;
        RECT 35.380 282.200 35.580 289.800 ;
        RECT 36.180 282.200 36.380 289.800 ;
        RECT 36.980 282.200 37.180 289.800 ;
        RECT 37.780 282.200 37.980 289.800 ;
        RECT 38.580 282.200 38.780 289.800 ;
        RECT 43.130 289.600 43.530 289.800 ;
        RECT 39.530 289.400 43.530 289.600 ;
        RECT 43.130 288.800 43.530 289.400 ;
        RECT 39.530 288.600 43.530 288.800 ;
        RECT 43.130 288.000 43.530 288.600 ;
        RECT 39.530 287.800 43.530 288.000 ;
        RECT 43.130 287.200 43.530 287.800 ;
        RECT 39.530 287.000 43.530 287.200 ;
        RECT 43.130 286.400 43.530 287.000 ;
        RECT 39.530 286.200 43.530 286.400 ;
        RECT 43.130 285.600 43.530 286.200 ;
        RECT 39.530 285.400 43.530 285.600 ;
        RECT 43.130 284.800 43.530 285.400 ;
        RECT 39.530 284.600 43.530 284.800 ;
        RECT 43.130 284.000 43.530 284.600 ;
        RECT 39.530 283.800 43.530 284.000 ;
        RECT 43.130 283.200 43.530 283.800 ;
        RECT 39.530 283.000 43.530 283.200 ;
        RECT 43.130 282.400 43.530 283.000 ;
        RECT 39.530 282.200 43.530 282.400 ;
        RECT 45.930 297.600 49.930 297.800 ;
        RECT 45.930 297.000 46.330 297.600 ;
        RECT 45.930 296.800 49.930 297.000 ;
        RECT 45.930 296.200 46.330 296.800 ;
        RECT 45.930 296.000 49.930 296.200 ;
        RECT 45.930 295.400 46.330 296.000 ;
        RECT 45.930 295.200 49.930 295.400 ;
        RECT 45.930 294.600 46.330 295.200 ;
        RECT 45.930 294.400 49.930 294.600 ;
        RECT 45.930 293.800 46.330 294.400 ;
        RECT 45.930 293.600 49.930 293.800 ;
        RECT 45.930 293.000 46.330 293.600 ;
        RECT 45.930 292.800 49.930 293.000 ;
        RECT 45.930 292.200 46.330 292.800 ;
        RECT 45.930 292.000 49.930 292.200 ;
        RECT 45.930 291.400 46.330 292.000 ;
        RECT 45.930 291.200 49.930 291.400 ;
        RECT 45.930 290.600 46.330 291.200 ;
        RECT 45.930 290.400 49.930 290.600 ;
        RECT 45.930 290.200 46.330 290.400 ;
        RECT 50.680 290.200 50.880 297.800 ;
        RECT 51.480 290.200 51.680 297.800 ;
        RECT 52.280 290.200 52.480 297.800 ;
        RECT 53.080 290.200 53.280 297.800 ;
        RECT 53.880 290.200 54.080 297.800 ;
        RECT 45.930 289.800 54.080 290.200 ;
        RECT 45.930 289.600 46.330 289.800 ;
        RECT 45.930 289.400 49.930 289.600 ;
        RECT 45.930 288.800 46.330 289.400 ;
        RECT 45.930 288.600 49.930 288.800 ;
        RECT 45.930 288.000 46.330 288.600 ;
        RECT 45.930 287.800 49.930 288.000 ;
        RECT 45.930 287.200 46.330 287.800 ;
        RECT 45.930 287.000 49.930 287.200 ;
        RECT 45.930 286.400 46.330 287.000 ;
        RECT 45.930 286.200 49.930 286.400 ;
        RECT 45.930 285.600 46.330 286.200 ;
        RECT 45.930 285.400 49.930 285.600 ;
        RECT 45.930 284.800 46.330 285.400 ;
        RECT 45.930 284.600 49.930 284.800 ;
        RECT 45.930 284.000 46.330 284.600 ;
        RECT 45.930 283.800 49.930 284.000 ;
        RECT 45.930 283.200 46.330 283.800 ;
        RECT 45.930 283.000 49.930 283.200 ;
        RECT 45.930 282.400 46.330 283.000 ;
        RECT 45.930 282.200 49.930 282.400 ;
        RECT 50.680 282.200 50.880 289.800 ;
        RECT 51.480 282.200 51.680 289.800 ;
        RECT 52.280 282.200 52.480 289.800 ;
        RECT 53.080 282.200 53.280 289.800 ;
        RECT 53.880 282.200 54.080 289.800 ;
        RECT 55.380 290.200 55.580 297.800 ;
        RECT 56.180 290.200 56.380 297.800 ;
        RECT 56.980 290.200 57.180 297.800 ;
        RECT 57.780 290.200 57.980 297.800 ;
        RECT 58.580 290.200 58.780 297.800 ;
        RECT 59.530 297.600 63.530 297.800 ;
        RECT 63.130 297.000 63.530 297.600 ;
        RECT 59.530 296.800 63.530 297.000 ;
        RECT 63.130 296.200 63.530 296.800 ;
        RECT 59.530 296.000 63.530 296.200 ;
        RECT 63.130 295.400 63.530 296.000 ;
        RECT 59.530 295.200 63.530 295.400 ;
        RECT 63.130 294.600 63.530 295.200 ;
        RECT 59.530 294.400 63.530 294.600 ;
        RECT 63.130 293.800 63.530 294.400 ;
        RECT 59.530 293.600 63.530 293.800 ;
        RECT 63.130 293.000 63.530 293.600 ;
        RECT 59.530 292.800 63.530 293.000 ;
        RECT 63.130 292.200 63.530 292.800 ;
        RECT 59.530 292.000 63.530 292.200 ;
        RECT 63.130 291.400 63.530 292.000 ;
        RECT 59.530 291.200 63.530 291.400 ;
        RECT 63.130 290.600 63.530 291.200 ;
        RECT 59.530 290.400 63.530 290.600 ;
        RECT 63.130 290.200 63.530 290.400 ;
        RECT 55.380 289.800 63.530 290.200 ;
        RECT 55.380 282.200 55.580 289.800 ;
        RECT 56.180 282.200 56.380 289.800 ;
        RECT 56.980 282.200 57.180 289.800 ;
        RECT 57.780 282.200 57.980 289.800 ;
        RECT 58.580 282.200 58.780 289.800 ;
        RECT 63.130 289.600 63.530 289.800 ;
        RECT 59.530 289.400 63.530 289.600 ;
        RECT 63.130 288.800 63.530 289.400 ;
        RECT 59.530 288.600 63.530 288.800 ;
        RECT 63.130 288.000 63.530 288.600 ;
        RECT 59.530 287.800 63.530 288.000 ;
        RECT 63.130 287.200 63.530 287.800 ;
        RECT 59.530 287.000 63.530 287.200 ;
        RECT 63.130 286.400 63.530 287.000 ;
        RECT 59.530 286.200 63.530 286.400 ;
        RECT 63.130 285.600 63.530 286.200 ;
        RECT 59.530 285.400 63.530 285.600 ;
        RECT 63.130 284.800 63.530 285.400 ;
        RECT 59.530 284.600 63.530 284.800 ;
        RECT 63.130 284.000 63.530 284.600 ;
        RECT 59.530 283.800 63.530 284.000 ;
        RECT 63.130 283.200 63.530 283.800 ;
        RECT 59.530 283.000 63.530 283.200 ;
        RECT 63.130 282.400 63.530 283.000 ;
        RECT 59.530 282.200 63.530 282.400 ;
        RECT 65.930 297.600 69.930 297.800 ;
        RECT 65.930 297.000 66.330 297.600 ;
        RECT 65.930 296.800 69.930 297.000 ;
        RECT 65.930 296.200 66.330 296.800 ;
        RECT 65.930 296.000 69.930 296.200 ;
        RECT 65.930 295.400 66.330 296.000 ;
        RECT 65.930 295.200 69.930 295.400 ;
        RECT 65.930 294.600 66.330 295.200 ;
        RECT 65.930 294.400 69.930 294.600 ;
        RECT 65.930 293.800 66.330 294.400 ;
        RECT 65.930 293.600 69.930 293.800 ;
        RECT 65.930 293.000 66.330 293.600 ;
        RECT 65.930 292.800 69.930 293.000 ;
        RECT 65.930 292.200 66.330 292.800 ;
        RECT 65.930 292.000 69.930 292.200 ;
        RECT 65.930 291.400 66.330 292.000 ;
        RECT 65.930 291.200 69.930 291.400 ;
        RECT 65.930 290.600 66.330 291.200 ;
        RECT 65.930 290.400 69.930 290.600 ;
        RECT 65.930 290.200 66.330 290.400 ;
        RECT 70.680 290.200 70.880 297.800 ;
        RECT 71.480 290.200 71.680 297.800 ;
        RECT 72.280 290.200 72.480 297.800 ;
        RECT 73.080 290.200 73.280 297.800 ;
        RECT 73.880 290.200 74.080 297.800 ;
        RECT 65.930 289.800 74.080 290.200 ;
        RECT 65.930 289.600 66.330 289.800 ;
        RECT 65.930 289.400 69.930 289.600 ;
        RECT 65.930 288.800 66.330 289.400 ;
        RECT 65.930 288.600 69.930 288.800 ;
        RECT 65.930 288.000 66.330 288.600 ;
        RECT 65.930 287.800 69.930 288.000 ;
        RECT 65.930 287.200 66.330 287.800 ;
        RECT 65.930 287.000 69.930 287.200 ;
        RECT 65.930 286.400 66.330 287.000 ;
        RECT 65.930 286.200 69.930 286.400 ;
        RECT 65.930 285.600 66.330 286.200 ;
        RECT 65.930 285.400 69.930 285.600 ;
        RECT 65.930 284.800 66.330 285.400 ;
        RECT 65.930 284.600 69.930 284.800 ;
        RECT 65.930 284.000 66.330 284.600 ;
        RECT 65.930 283.800 69.930 284.000 ;
        RECT 65.930 283.200 66.330 283.800 ;
        RECT 65.930 283.000 69.930 283.200 ;
        RECT 65.930 282.400 66.330 283.000 ;
        RECT 65.930 282.200 69.930 282.400 ;
        RECT 70.680 282.200 70.880 289.800 ;
        RECT 71.480 282.200 71.680 289.800 ;
        RECT 72.280 282.200 72.480 289.800 ;
        RECT 73.080 282.200 73.280 289.800 ;
        RECT 73.880 282.200 74.080 289.800 ;
        RECT 75.380 290.200 75.580 297.800 ;
        RECT 76.180 290.200 76.380 297.800 ;
        RECT 76.980 290.200 77.180 297.800 ;
        RECT 77.780 290.200 77.980 297.800 ;
        RECT 78.580 290.200 78.780 297.800 ;
        RECT 79.530 297.600 83.530 297.800 ;
        RECT 83.130 297.000 83.530 297.600 ;
        RECT 79.530 296.800 83.530 297.000 ;
        RECT 83.130 296.200 83.530 296.800 ;
        RECT 79.530 296.000 83.530 296.200 ;
        RECT 83.130 295.400 83.530 296.000 ;
        RECT 79.530 295.200 83.530 295.400 ;
        RECT 83.130 294.600 83.530 295.200 ;
        RECT 79.530 294.400 83.530 294.600 ;
        RECT 83.130 293.800 83.530 294.400 ;
        RECT 79.530 293.600 83.530 293.800 ;
        RECT 83.130 293.000 83.530 293.600 ;
        RECT 79.530 292.800 83.530 293.000 ;
        RECT 83.130 292.200 83.530 292.800 ;
        RECT 79.530 292.000 83.530 292.200 ;
        RECT 83.130 291.400 83.530 292.000 ;
        RECT 79.530 291.200 83.530 291.400 ;
        RECT 83.130 290.600 83.530 291.200 ;
        RECT 79.530 290.400 83.530 290.600 ;
        RECT 83.130 290.200 83.530 290.400 ;
        RECT 75.380 289.800 83.530 290.200 ;
        RECT 75.380 282.200 75.580 289.800 ;
        RECT 76.180 282.200 76.380 289.800 ;
        RECT 76.980 282.200 77.180 289.800 ;
        RECT 77.780 282.200 77.980 289.800 ;
        RECT 78.580 282.200 78.780 289.800 ;
        RECT 83.130 289.600 83.530 289.800 ;
        RECT 79.530 289.400 83.530 289.600 ;
        RECT 83.130 288.800 83.530 289.400 ;
        RECT 79.530 288.600 83.530 288.800 ;
        RECT 83.130 288.000 83.530 288.600 ;
        RECT 79.530 287.800 83.530 288.000 ;
        RECT 83.130 287.200 83.530 287.800 ;
        RECT 79.530 287.000 83.530 287.200 ;
        RECT 83.130 286.400 83.530 287.000 ;
        RECT 79.530 286.200 83.530 286.400 ;
        RECT 83.130 285.600 83.530 286.200 ;
        RECT 79.530 285.400 83.530 285.600 ;
        RECT 83.130 284.800 83.530 285.400 ;
        RECT 79.530 284.600 83.530 284.800 ;
        RECT 83.130 284.000 83.530 284.600 ;
        RECT 79.530 283.800 83.530 284.000 ;
        RECT 83.130 283.200 83.530 283.800 ;
        RECT 79.530 283.000 83.530 283.200 ;
        RECT 83.130 282.400 83.530 283.000 ;
        RECT 79.530 282.200 83.530 282.400 ;
        RECT 85.930 297.600 89.930 297.800 ;
        RECT 85.930 297.000 86.330 297.600 ;
        RECT 85.930 296.800 89.930 297.000 ;
        RECT 85.930 296.200 86.330 296.800 ;
        RECT 85.930 296.000 89.930 296.200 ;
        RECT 85.930 295.400 86.330 296.000 ;
        RECT 85.930 295.200 89.930 295.400 ;
        RECT 85.930 294.600 86.330 295.200 ;
        RECT 85.930 294.400 89.930 294.600 ;
        RECT 85.930 293.800 86.330 294.400 ;
        RECT 85.930 293.600 89.930 293.800 ;
        RECT 85.930 293.000 86.330 293.600 ;
        RECT 85.930 292.800 89.930 293.000 ;
        RECT 85.930 292.200 86.330 292.800 ;
        RECT 85.930 292.000 89.930 292.200 ;
        RECT 85.930 291.400 86.330 292.000 ;
        RECT 85.930 291.200 89.930 291.400 ;
        RECT 85.930 290.600 86.330 291.200 ;
        RECT 85.930 290.400 89.930 290.600 ;
        RECT 85.930 290.200 86.330 290.400 ;
        RECT 90.680 290.200 90.880 297.800 ;
        RECT 91.480 290.200 91.680 297.800 ;
        RECT 92.280 290.200 92.480 297.800 ;
        RECT 93.080 290.200 93.280 297.800 ;
        RECT 93.880 290.200 94.080 297.800 ;
        RECT 85.930 289.800 94.080 290.200 ;
        RECT 85.930 289.600 86.330 289.800 ;
        RECT 85.930 289.400 89.930 289.600 ;
        RECT 85.930 288.800 86.330 289.400 ;
        RECT 85.930 288.600 89.930 288.800 ;
        RECT 85.930 288.000 86.330 288.600 ;
        RECT 85.930 287.800 89.930 288.000 ;
        RECT 85.930 287.200 86.330 287.800 ;
        RECT 85.930 287.000 89.930 287.200 ;
        RECT 85.930 286.400 86.330 287.000 ;
        RECT 85.930 286.200 89.930 286.400 ;
        RECT 85.930 285.600 86.330 286.200 ;
        RECT 85.930 285.400 89.930 285.600 ;
        RECT 85.930 284.800 86.330 285.400 ;
        RECT 85.930 284.600 89.930 284.800 ;
        RECT 85.930 284.000 86.330 284.600 ;
        RECT 85.930 283.800 89.930 284.000 ;
        RECT 85.930 283.200 86.330 283.800 ;
        RECT 85.930 283.000 89.930 283.200 ;
        RECT 85.930 282.400 86.330 283.000 ;
        RECT 85.930 282.200 89.930 282.400 ;
        RECT 90.680 282.200 90.880 289.800 ;
        RECT 91.480 282.200 91.680 289.800 ;
        RECT 92.280 282.200 92.480 289.800 ;
        RECT 93.080 282.200 93.280 289.800 ;
        RECT 93.880 282.200 94.080 289.800 ;
        RECT 95.380 290.200 95.580 297.800 ;
        RECT 96.180 290.200 96.380 297.800 ;
        RECT 96.980 290.200 97.180 297.800 ;
        RECT 97.780 290.200 97.980 297.800 ;
        RECT 98.580 290.200 98.780 297.800 ;
        RECT 99.530 297.600 103.530 297.800 ;
        RECT 103.130 297.000 103.530 297.600 ;
        RECT 99.530 296.800 103.530 297.000 ;
        RECT 103.130 296.200 103.530 296.800 ;
        RECT 99.530 296.000 103.530 296.200 ;
        RECT 103.130 295.400 103.530 296.000 ;
        RECT 99.530 295.200 103.530 295.400 ;
        RECT 103.130 294.600 103.530 295.200 ;
        RECT 99.530 294.400 103.530 294.600 ;
        RECT 103.130 293.800 103.530 294.400 ;
        RECT 99.530 293.600 103.530 293.800 ;
        RECT 103.130 293.000 103.530 293.600 ;
        RECT 99.530 292.800 103.530 293.000 ;
        RECT 103.130 292.200 103.530 292.800 ;
        RECT 99.530 292.000 103.530 292.200 ;
        RECT 103.130 291.400 103.530 292.000 ;
        RECT 99.530 291.200 103.530 291.400 ;
        RECT 103.130 290.600 103.530 291.200 ;
        RECT 99.530 290.400 103.530 290.600 ;
        RECT 103.130 290.200 103.530 290.400 ;
        RECT 95.380 289.800 103.530 290.200 ;
        RECT 110.050 290.100 110.410 290.480 ;
        RECT 110.680 290.100 111.040 290.480 ;
        RECT 111.280 290.100 111.640 290.480 ;
        RECT 95.380 282.200 95.580 289.800 ;
        RECT 96.180 282.200 96.380 289.800 ;
        RECT 96.980 282.200 97.180 289.800 ;
        RECT 97.780 282.200 97.980 289.800 ;
        RECT 98.580 282.200 98.780 289.800 ;
        RECT 103.130 289.600 103.530 289.800 ;
        RECT 99.530 289.400 103.530 289.600 ;
        RECT 110.050 289.510 110.410 289.890 ;
        RECT 110.680 289.510 111.040 289.890 ;
        RECT 111.280 289.510 111.640 289.890 ;
        RECT 103.130 288.800 103.530 289.400 ;
        RECT 99.530 288.600 103.530 288.800 ;
        RECT 103.130 288.000 103.530 288.600 ;
        RECT 99.530 287.800 103.530 288.000 ;
        RECT 103.130 287.200 103.530 287.800 ;
        RECT 99.530 287.000 103.530 287.200 ;
        RECT 103.130 286.400 103.530 287.000 ;
        RECT 99.530 286.200 103.530 286.400 ;
        RECT 103.130 285.600 103.530 286.200 ;
        RECT 99.530 285.400 103.530 285.600 ;
        RECT 103.130 284.800 103.530 285.400 ;
        RECT 99.530 284.600 103.530 284.800 ;
        RECT 103.130 284.000 103.530 284.600 ;
        RECT 99.530 283.800 103.530 284.000 ;
        RECT 103.130 283.200 103.530 283.800 ;
        RECT 99.530 283.000 103.530 283.200 ;
        RECT 103.130 282.400 103.530 283.000 ;
        RECT 99.530 282.200 103.530 282.400 ;
        RECT 5.930 277.600 9.930 277.800 ;
        RECT 5.930 277.000 6.330 277.600 ;
        RECT 5.930 276.800 9.930 277.000 ;
        RECT 5.930 276.200 6.330 276.800 ;
        RECT 5.930 276.000 9.930 276.200 ;
        RECT 5.930 275.400 6.330 276.000 ;
        RECT 5.930 275.200 9.930 275.400 ;
        RECT 5.930 274.600 6.330 275.200 ;
        RECT 5.930 274.400 9.930 274.600 ;
        RECT 5.930 273.800 6.330 274.400 ;
        RECT 5.930 273.600 9.930 273.800 ;
        RECT 5.930 273.000 6.330 273.600 ;
        RECT 5.930 272.800 9.930 273.000 ;
        RECT 5.930 272.200 6.330 272.800 ;
        RECT 5.930 272.000 9.930 272.200 ;
        RECT 5.930 271.400 6.330 272.000 ;
        RECT 5.930 271.200 9.930 271.400 ;
        RECT 5.930 270.600 6.330 271.200 ;
        RECT 5.930 270.400 9.930 270.600 ;
        RECT 5.930 270.200 6.330 270.400 ;
        RECT 10.680 270.200 10.880 277.800 ;
        RECT 11.480 270.200 11.680 277.800 ;
        RECT 12.280 270.200 12.480 277.800 ;
        RECT 13.080 270.200 13.280 277.800 ;
        RECT 13.880 270.200 14.080 277.800 ;
        RECT 5.930 269.800 14.080 270.200 ;
        RECT 5.930 269.600 6.330 269.800 ;
        RECT 5.930 269.400 9.930 269.600 ;
        RECT 5.930 268.800 6.330 269.400 ;
        RECT 5.930 268.600 9.930 268.800 ;
        RECT 5.930 268.000 6.330 268.600 ;
        RECT 5.930 267.800 9.930 268.000 ;
        RECT 5.930 267.200 6.330 267.800 ;
        RECT 5.930 267.000 9.930 267.200 ;
        RECT 5.930 266.400 6.330 267.000 ;
        RECT 5.930 266.200 9.930 266.400 ;
        RECT 5.930 265.600 6.330 266.200 ;
        RECT 5.930 265.400 9.930 265.600 ;
        RECT 5.930 264.800 6.330 265.400 ;
        RECT 5.930 264.600 9.930 264.800 ;
        RECT 5.930 264.000 6.330 264.600 ;
        RECT 5.930 263.800 9.930 264.000 ;
        RECT 5.930 263.200 6.330 263.800 ;
        RECT 5.930 263.000 9.930 263.200 ;
        RECT 5.930 262.400 6.330 263.000 ;
        RECT 5.930 262.200 9.930 262.400 ;
        RECT 10.680 262.200 10.880 269.800 ;
        RECT 11.480 262.200 11.680 269.800 ;
        RECT 12.280 262.200 12.480 269.800 ;
        RECT 13.080 262.200 13.280 269.800 ;
        RECT 13.880 262.200 14.080 269.800 ;
        RECT 15.380 270.200 15.580 277.800 ;
        RECT 16.180 270.200 16.380 277.800 ;
        RECT 16.980 270.200 17.180 277.800 ;
        RECT 17.780 270.200 17.980 277.800 ;
        RECT 18.580 270.200 18.780 277.800 ;
        RECT 19.530 277.600 23.530 277.800 ;
        RECT 23.130 277.000 23.530 277.600 ;
        RECT 19.530 276.800 23.530 277.000 ;
        RECT 23.130 276.200 23.530 276.800 ;
        RECT 19.530 276.000 23.530 276.200 ;
        RECT 23.130 275.400 23.530 276.000 ;
        RECT 19.530 275.200 23.530 275.400 ;
        RECT 23.130 274.600 23.530 275.200 ;
        RECT 19.530 274.400 23.530 274.600 ;
        RECT 23.130 273.800 23.530 274.400 ;
        RECT 19.530 273.600 23.530 273.800 ;
        RECT 23.130 273.000 23.530 273.600 ;
        RECT 19.530 272.800 23.530 273.000 ;
        RECT 23.130 272.200 23.530 272.800 ;
        RECT 19.530 272.000 23.530 272.200 ;
        RECT 23.130 271.400 23.530 272.000 ;
        RECT 19.530 271.200 23.530 271.400 ;
        RECT 23.130 270.600 23.530 271.200 ;
        RECT 19.530 270.400 23.530 270.600 ;
        RECT 23.130 270.200 23.530 270.400 ;
        RECT 15.380 269.800 23.530 270.200 ;
        RECT 15.380 262.200 15.580 269.800 ;
        RECT 16.180 262.200 16.380 269.800 ;
        RECT 16.980 262.200 17.180 269.800 ;
        RECT 17.780 262.200 17.980 269.800 ;
        RECT 18.580 262.200 18.780 269.800 ;
        RECT 23.130 269.600 23.530 269.800 ;
        RECT 19.530 269.400 23.530 269.600 ;
        RECT 23.130 268.800 23.530 269.400 ;
        RECT 19.530 268.600 23.530 268.800 ;
        RECT 23.130 268.000 23.530 268.600 ;
        RECT 19.530 267.800 23.530 268.000 ;
        RECT 23.130 267.200 23.530 267.800 ;
        RECT 19.530 267.000 23.530 267.200 ;
        RECT 23.130 266.400 23.530 267.000 ;
        RECT 19.530 266.200 23.530 266.400 ;
        RECT 23.130 265.600 23.530 266.200 ;
        RECT 19.530 265.400 23.530 265.600 ;
        RECT 23.130 264.800 23.530 265.400 ;
        RECT 19.530 264.600 23.530 264.800 ;
        RECT 23.130 264.000 23.530 264.600 ;
        RECT 19.530 263.800 23.530 264.000 ;
        RECT 23.130 263.200 23.530 263.800 ;
        RECT 19.530 263.000 23.530 263.200 ;
        RECT 23.130 262.400 23.530 263.000 ;
        RECT 19.530 262.200 23.530 262.400 ;
        RECT 25.930 277.600 29.930 277.800 ;
        RECT 25.930 277.000 26.330 277.600 ;
        RECT 25.930 276.800 29.930 277.000 ;
        RECT 25.930 276.200 26.330 276.800 ;
        RECT 25.930 276.000 29.930 276.200 ;
        RECT 25.930 275.400 26.330 276.000 ;
        RECT 25.930 275.200 29.930 275.400 ;
        RECT 25.930 274.600 26.330 275.200 ;
        RECT 25.930 274.400 29.930 274.600 ;
        RECT 25.930 273.800 26.330 274.400 ;
        RECT 25.930 273.600 29.930 273.800 ;
        RECT 25.930 273.000 26.330 273.600 ;
        RECT 25.930 272.800 29.930 273.000 ;
        RECT 25.930 272.200 26.330 272.800 ;
        RECT 25.930 272.000 29.930 272.200 ;
        RECT 25.930 271.400 26.330 272.000 ;
        RECT 25.930 271.200 29.930 271.400 ;
        RECT 25.930 270.600 26.330 271.200 ;
        RECT 25.930 270.400 29.930 270.600 ;
        RECT 25.930 270.200 26.330 270.400 ;
        RECT 30.680 270.200 30.880 277.800 ;
        RECT 31.480 270.200 31.680 277.800 ;
        RECT 32.280 270.200 32.480 277.800 ;
        RECT 33.080 270.200 33.280 277.800 ;
        RECT 33.880 270.200 34.080 277.800 ;
        RECT 25.930 269.800 34.080 270.200 ;
        RECT 25.930 269.600 26.330 269.800 ;
        RECT 25.930 269.400 29.930 269.600 ;
        RECT 25.930 268.800 26.330 269.400 ;
        RECT 25.930 268.600 29.930 268.800 ;
        RECT 25.930 268.000 26.330 268.600 ;
        RECT 25.930 267.800 29.930 268.000 ;
        RECT 25.930 267.200 26.330 267.800 ;
        RECT 25.930 267.000 29.930 267.200 ;
        RECT 25.930 266.400 26.330 267.000 ;
        RECT 25.930 266.200 29.930 266.400 ;
        RECT 25.930 265.600 26.330 266.200 ;
        RECT 25.930 265.400 29.930 265.600 ;
        RECT 25.930 264.800 26.330 265.400 ;
        RECT 25.930 264.600 29.930 264.800 ;
        RECT 25.930 264.000 26.330 264.600 ;
        RECT 25.930 263.800 29.930 264.000 ;
        RECT 25.930 263.200 26.330 263.800 ;
        RECT 25.930 263.000 29.930 263.200 ;
        RECT 25.930 262.400 26.330 263.000 ;
        RECT 25.930 262.200 29.930 262.400 ;
        RECT 30.680 262.200 30.880 269.800 ;
        RECT 31.480 262.200 31.680 269.800 ;
        RECT 32.280 262.200 32.480 269.800 ;
        RECT 33.080 262.200 33.280 269.800 ;
        RECT 33.880 262.200 34.080 269.800 ;
        RECT 35.380 270.200 35.580 277.800 ;
        RECT 36.180 270.200 36.380 277.800 ;
        RECT 36.980 270.200 37.180 277.800 ;
        RECT 37.780 270.200 37.980 277.800 ;
        RECT 38.580 270.200 38.780 277.800 ;
        RECT 39.530 277.600 43.530 277.800 ;
        RECT 43.130 277.000 43.530 277.600 ;
        RECT 39.530 276.800 43.530 277.000 ;
        RECT 43.130 276.200 43.530 276.800 ;
        RECT 39.530 276.000 43.530 276.200 ;
        RECT 43.130 275.400 43.530 276.000 ;
        RECT 39.530 275.200 43.530 275.400 ;
        RECT 43.130 274.600 43.530 275.200 ;
        RECT 39.530 274.400 43.530 274.600 ;
        RECT 43.130 273.800 43.530 274.400 ;
        RECT 39.530 273.600 43.530 273.800 ;
        RECT 43.130 273.000 43.530 273.600 ;
        RECT 39.530 272.800 43.530 273.000 ;
        RECT 43.130 272.200 43.530 272.800 ;
        RECT 39.530 272.000 43.530 272.200 ;
        RECT 43.130 271.400 43.530 272.000 ;
        RECT 39.530 271.200 43.530 271.400 ;
        RECT 43.130 270.600 43.530 271.200 ;
        RECT 39.530 270.400 43.530 270.600 ;
        RECT 43.130 270.200 43.530 270.400 ;
        RECT 35.380 269.800 43.530 270.200 ;
        RECT 35.380 262.200 35.580 269.800 ;
        RECT 36.180 262.200 36.380 269.800 ;
        RECT 36.980 262.200 37.180 269.800 ;
        RECT 37.780 262.200 37.980 269.800 ;
        RECT 38.580 262.200 38.780 269.800 ;
        RECT 43.130 269.600 43.530 269.800 ;
        RECT 39.530 269.400 43.530 269.600 ;
        RECT 43.130 268.800 43.530 269.400 ;
        RECT 39.530 268.600 43.530 268.800 ;
        RECT 43.130 268.000 43.530 268.600 ;
        RECT 39.530 267.800 43.530 268.000 ;
        RECT 43.130 267.200 43.530 267.800 ;
        RECT 39.530 267.000 43.530 267.200 ;
        RECT 43.130 266.400 43.530 267.000 ;
        RECT 39.530 266.200 43.530 266.400 ;
        RECT 43.130 265.600 43.530 266.200 ;
        RECT 39.530 265.400 43.530 265.600 ;
        RECT 43.130 264.800 43.530 265.400 ;
        RECT 39.530 264.600 43.530 264.800 ;
        RECT 43.130 264.000 43.530 264.600 ;
        RECT 39.530 263.800 43.530 264.000 ;
        RECT 43.130 263.200 43.530 263.800 ;
        RECT 39.530 263.000 43.530 263.200 ;
        RECT 43.130 262.400 43.530 263.000 ;
        RECT 39.530 262.200 43.530 262.400 ;
        RECT 45.930 277.600 49.930 277.800 ;
        RECT 45.930 277.000 46.330 277.600 ;
        RECT 45.930 276.800 49.930 277.000 ;
        RECT 45.930 276.200 46.330 276.800 ;
        RECT 45.930 276.000 49.930 276.200 ;
        RECT 45.930 275.400 46.330 276.000 ;
        RECT 45.930 275.200 49.930 275.400 ;
        RECT 45.930 274.600 46.330 275.200 ;
        RECT 45.930 274.400 49.930 274.600 ;
        RECT 45.930 273.800 46.330 274.400 ;
        RECT 45.930 273.600 49.930 273.800 ;
        RECT 45.930 273.000 46.330 273.600 ;
        RECT 45.930 272.800 49.930 273.000 ;
        RECT 45.930 272.200 46.330 272.800 ;
        RECT 45.930 272.000 49.930 272.200 ;
        RECT 45.930 271.400 46.330 272.000 ;
        RECT 45.930 271.200 49.930 271.400 ;
        RECT 45.930 270.600 46.330 271.200 ;
        RECT 45.930 270.400 49.930 270.600 ;
        RECT 45.930 270.200 46.330 270.400 ;
        RECT 50.680 270.200 50.880 277.800 ;
        RECT 51.480 270.200 51.680 277.800 ;
        RECT 52.280 270.200 52.480 277.800 ;
        RECT 53.080 270.200 53.280 277.800 ;
        RECT 53.880 270.200 54.080 277.800 ;
        RECT 45.930 269.800 54.080 270.200 ;
        RECT 45.930 269.600 46.330 269.800 ;
        RECT 45.930 269.400 49.930 269.600 ;
        RECT 45.930 268.800 46.330 269.400 ;
        RECT 45.930 268.600 49.930 268.800 ;
        RECT 45.930 268.000 46.330 268.600 ;
        RECT 45.930 267.800 49.930 268.000 ;
        RECT 45.930 267.200 46.330 267.800 ;
        RECT 45.930 267.000 49.930 267.200 ;
        RECT 45.930 266.400 46.330 267.000 ;
        RECT 45.930 266.200 49.930 266.400 ;
        RECT 45.930 265.600 46.330 266.200 ;
        RECT 45.930 265.400 49.930 265.600 ;
        RECT 45.930 264.800 46.330 265.400 ;
        RECT 45.930 264.600 49.930 264.800 ;
        RECT 45.930 264.000 46.330 264.600 ;
        RECT 45.930 263.800 49.930 264.000 ;
        RECT 45.930 263.200 46.330 263.800 ;
        RECT 45.930 263.000 49.930 263.200 ;
        RECT 45.930 262.400 46.330 263.000 ;
        RECT 45.930 262.200 49.930 262.400 ;
        RECT 50.680 262.200 50.880 269.800 ;
        RECT 51.480 262.200 51.680 269.800 ;
        RECT 52.280 262.200 52.480 269.800 ;
        RECT 53.080 262.200 53.280 269.800 ;
        RECT 53.880 262.200 54.080 269.800 ;
        RECT 55.380 270.200 55.580 277.800 ;
        RECT 56.180 270.200 56.380 277.800 ;
        RECT 56.980 270.200 57.180 277.800 ;
        RECT 57.780 270.200 57.980 277.800 ;
        RECT 58.580 270.200 58.780 277.800 ;
        RECT 59.530 277.600 63.530 277.800 ;
        RECT 63.130 277.000 63.530 277.600 ;
        RECT 59.530 276.800 63.530 277.000 ;
        RECT 63.130 276.200 63.530 276.800 ;
        RECT 59.530 276.000 63.530 276.200 ;
        RECT 63.130 275.400 63.530 276.000 ;
        RECT 59.530 275.200 63.530 275.400 ;
        RECT 63.130 274.600 63.530 275.200 ;
        RECT 59.530 274.400 63.530 274.600 ;
        RECT 63.130 273.800 63.530 274.400 ;
        RECT 59.530 273.600 63.530 273.800 ;
        RECT 63.130 273.000 63.530 273.600 ;
        RECT 59.530 272.800 63.530 273.000 ;
        RECT 63.130 272.200 63.530 272.800 ;
        RECT 59.530 272.000 63.530 272.200 ;
        RECT 63.130 271.400 63.530 272.000 ;
        RECT 59.530 271.200 63.530 271.400 ;
        RECT 63.130 270.600 63.530 271.200 ;
        RECT 59.530 270.400 63.530 270.600 ;
        RECT 63.130 270.200 63.530 270.400 ;
        RECT 55.380 269.800 63.530 270.200 ;
        RECT 55.380 262.200 55.580 269.800 ;
        RECT 56.180 262.200 56.380 269.800 ;
        RECT 56.980 262.200 57.180 269.800 ;
        RECT 57.780 262.200 57.980 269.800 ;
        RECT 58.580 262.200 58.780 269.800 ;
        RECT 63.130 269.600 63.530 269.800 ;
        RECT 59.530 269.400 63.530 269.600 ;
        RECT 63.130 268.800 63.530 269.400 ;
        RECT 59.530 268.600 63.530 268.800 ;
        RECT 63.130 268.000 63.530 268.600 ;
        RECT 59.530 267.800 63.530 268.000 ;
        RECT 63.130 267.200 63.530 267.800 ;
        RECT 59.530 267.000 63.530 267.200 ;
        RECT 63.130 266.400 63.530 267.000 ;
        RECT 59.530 266.200 63.530 266.400 ;
        RECT 63.130 265.600 63.530 266.200 ;
        RECT 59.530 265.400 63.530 265.600 ;
        RECT 63.130 264.800 63.530 265.400 ;
        RECT 59.530 264.600 63.530 264.800 ;
        RECT 63.130 264.000 63.530 264.600 ;
        RECT 59.530 263.800 63.530 264.000 ;
        RECT 63.130 263.200 63.530 263.800 ;
        RECT 59.530 263.000 63.530 263.200 ;
        RECT 63.130 262.400 63.530 263.000 ;
        RECT 59.530 262.200 63.530 262.400 ;
        RECT 65.930 277.600 69.930 277.800 ;
        RECT 65.930 277.000 66.330 277.600 ;
        RECT 65.930 276.800 69.930 277.000 ;
        RECT 65.930 276.200 66.330 276.800 ;
        RECT 65.930 276.000 69.930 276.200 ;
        RECT 65.930 275.400 66.330 276.000 ;
        RECT 65.930 275.200 69.930 275.400 ;
        RECT 65.930 274.600 66.330 275.200 ;
        RECT 65.930 274.400 69.930 274.600 ;
        RECT 65.930 273.800 66.330 274.400 ;
        RECT 65.930 273.600 69.930 273.800 ;
        RECT 65.930 273.000 66.330 273.600 ;
        RECT 65.930 272.800 69.930 273.000 ;
        RECT 65.930 272.200 66.330 272.800 ;
        RECT 65.930 272.000 69.930 272.200 ;
        RECT 65.930 271.400 66.330 272.000 ;
        RECT 65.930 271.200 69.930 271.400 ;
        RECT 65.930 270.600 66.330 271.200 ;
        RECT 65.930 270.400 69.930 270.600 ;
        RECT 65.930 270.200 66.330 270.400 ;
        RECT 70.680 270.200 70.880 277.800 ;
        RECT 71.480 270.200 71.680 277.800 ;
        RECT 72.280 270.200 72.480 277.800 ;
        RECT 73.080 270.200 73.280 277.800 ;
        RECT 73.880 270.200 74.080 277.800 ;
        RECT 65.930 269.800 74.080 270.200 ;
        RECT 65.930 269.600 66.330 269.800 ;
        RECT 65.930 269.400 69.930 269.600 ;
        RECT 65.930 268.800 66.330 269.400 ;
        RECT 65.930 268.600 69.930 268.800 ;
        RECT 65.930 268.000 66.330 268.600 ;
        RECT 65.930 267.800 69.930 268.000 ;
        RECT 65.930 267.200 66.330 267.800 ;
        RECT 65.930 267.000 69.930 267.200 ;
        RECT 65.930 266.400 66.330 267.000 ;
        RECT 65.930 266.200 69.930 266.400 ;
        RECT 65.930 265.600 66.330 266.200 ;
        RECT 65.930 265.400 69.930 265.600 ;
        RECT 65.930 264.800 66.330 265.400 ;
        RECT 65.930 264.600 69.930 264.800 ;
        RECT 65.930 264.000 66.330 264.600 ;
        RECT 65.930 263.800 69.930 264.000 ;
        RECT 65.930 263.200 66.330 263.800 ;
        RECT 65.930 263.000 69.930 263.200 ;
        RECT 65.930 262.400 66.330 263.000 ;
        RECT 65.930 262.200 69.930 262.400 ;
        RECT 70.680 262.200 70.880 269.800 ;
        RECT 71.480 262.200 71.680 269.800 ;
        RECT 72.280 262.200 72.480 269.800 ;
        RECT 73.080 262.200 73.280 269.800 ;
        RECT 73.880 262.200 74.080 269.800 ;
        RECT 75.380 270.200 75.580 277.800 ;
        RECT 76.180 270.200 76.380 277.800 ;
        RECT 76.980 270.200 77.180 277.800 ;
        RECT 77.780 270.200 77.980 277.800 ;
        RECT 78.580 270.200 78.780 277.800 ;
        RECT 79.530 277.600 83.530 277.800 ;
        RECT 83.130 277.000 83.530 277.600 ;
        RECT 79.530 276.800 83.530 277.000 ;
        RECT 83.130 276.200 83.530 276.800 ;
        RECT 79.530 276.000 83.530 276.200 ;
        RECT 83.130 275.400 83.530 276.000 ;
        RECT 79.530 275.200 83.530 275.400 ;
        RECT 83.130 274.600 83.530 275.200 ;
        RECT 79.530 274.400 83.530 274.600 ;
        RECT 83.130 273.800 83.530 274.400 ;
        RECT 79.530 273.600 83.530 273.800 ;
        RECT 83.130 273.000 83.530 273.600 ;
        RECT 79.530 272.800 83.530 273.000 ;
        RECT 83.130 272.200 83.530 272.800 ;
        RECT 79.530 272.000 83.530 272.200 ;
        RECT 83.130 271.400 83.530 272.000 ;
        RECT 79.530 271.200 83.530 271.400 ;
        RECT 83.130 270.600 83.530 271.200 ;
        RECT 79.530 270.400 83.530 270.600 ;
        RECT 83.130 270.200 83.530 270.400 ;
        RECT 75.380 269.800 83.530 270.200 ;
        RECT 75.380 262.200 75.580 269.800 ;
        RECT 76.180 262.200 76.380 269.800 ;
        RECT 76.980 262.200 77.180 269.800 ;
        RECT 77.780 262.200 77.980 269.800 ;
        RECT 78.580 262.200 78.780 269.800 ;
        RECT 83.130 269.600 83.530 269.800 ;
        RECT 79.530 269.400 83.530 269.600 ;
        RECT 83.130 268.800 83.530 269.400 ;
        RECT 79.530 268.600 83.530 268.800 ;
        RECT 83.130 268.000 83.530 268.600 ;
        RECT 79.530 267.800 83.530 268.000 ;
        RECT 83.130 267.200 83.530 267.800 ;
        RECT 79.530 267.000 83.530 267.200 ;
        RECT 83.130 266.400 83.530 267.000 ;
        RECT 79.530 266.200 83.530 266.400 ;
        RECT 83.130 265.600 83.530 266.200 ;
        RECT 79.530 265.400 83.530 265.600 ;
        RECT 83.130 264.800 83.530 265.400 ;
        RECT 79.530 264.600 83.530 264.800 ;
        RECT 83.130 264.000 83.530 264.600 ;
        RECT 79.530 263.800 83.530 264.000 ;
        RECT 83.130 263.200 83.530 263.800 ;
        RECT 79.530 263.000 83.530 263.200 ;
        RECT 83.130 262.400 83.530 263.000 ;
        RECT 79.530 262.200 83.530 262.400 ;
        RECT 85.930 277.600 89.930 277.800 ;
        RECT 85.930 277.000 86.330 277.600 ;
        RECT 85.930 276.800 89.930 277.000 ;
        RECT 85.930 276.200 86.330 276.800 ;
        RECT 85.930 276.000 89.930 276.200 ;
        RECT 85.930 275.400 86.330 276.000 ;
        RECT 85.930 275.200 89.930 275.400 ;
        RECT 85.930 274.600 86.330 275.200 ;
        RECT 85.930 274.400 89.930 274.600 ;
        RECT 85.930 273.800 86.330 274.400 ;
        RECT 85.930 273.600 89.930 273.800 ;
        RECT 85.930 273.000 86.330 273.600 ;
        RECT 85.930 272.800 89.930 273.000 ;
        RECT 85.930 272.200 86.330 272.800 ;
        RECT 85.930 272.000 89.930 272.200 ;
        RECT 85.930 271.400 86.330 272.000 ;
        RECT 85.930 271.200 89.930 271.400 ;
        RECT 85.930 270.600 86.330 271.200 ;
        RECT 85.930 270.400 89.930 270.600 ;
        RECT 85.930 270.200 86.330 270.400 ;
        RECT 90.680 270.200 90.880 277.800 ;
        RECT 91.480 270.200 91.680 277.800 ;
        RECT 92.280 270.200 92.480 277.800 ;
        RECT 93.080 270.200 93.280 277.800 ;
        RECT 93.880 270.200 94.080 277.800 ;
        RECT 85.930 269.800 94.080 270.200 ;
        RECT 85.930 269.600 86.330 269.800 ;
        RECT 85.930 269.400 89.930 269.600 ;
        RECT 85.930 268.800 86.330 269.400 ;
        RECT 85.930 268.600 89.930 268.800 ;
        RECT 85.930 268.000 86.330 268.600 ;
        RECT 85.930 267.800 89.930 268.000 ;
        RECT 85.930 267.200 86.330 267.800 ;
        RECT 85.930 267.000 89.930 267.200 ;
        RECT 85.930 266.400 86.330 267.000 ;
        RECT 85.930 266.200 89.930 266.400 ;
        RECT 85.930 265.600 86.330 266.200 ;
        RECT 85.930 265.400 89.930 265.600 ;
        RECT 85.930 264.800 86.330 265.400 ;
        RECT 85.930 264.600 89.930 264.800 ;
        RECT 85.930 264.000 86.330 264.600 ;
        RECT 85.930 263.800 89.930 264.000 ;
        RECT 85.930 263.200 86.330 263.800 ;
        RECT 85.930 263.000 89.930 263.200 ;
        RECT 85.930 262.400 86.330 263.000 ;
        RECT 85.930 262.200 89.930 262.400 ;
        RECT 90.680 262.200 90.880 269.800 ;
        RECT 91.480 262.200 91.680 269.800 ;
        RECT 92.280 262.200 92.480 269.800 ;
        RECT 93.080 262.200 93.280 269.800 ;
        RECT 93.880 262.200 94.080 269.800 ;
        RECT 95.380 270.200 95.580 277.800 ;
        RECT 96.180 270.200 96.380 277.800 ;
        RECT 96.980 270.200 97.180 277.800 ;
        RECT 97.780 270.200 97.980 277.800 ;
        RECT 98.580 270.200 98.780 277.800 ;
        RECT 99.530 277.600 103.530 277.800 ;
        RECT 103.130 277.000 103.530 277.600 ;
        RECT 99.530 276.800 103.530 277.000 ;
        RECT 103.130 276.200 103.530 276.800 ;
        RECT 99.530 276.000 103.530 276.200 ;
        RECT 103.130 275.400 103.530 276.000 ;
        RECT 99.530 275.200 103.530 275.400 ;
        RECT 103.130 274.600 103.530 275.200 ;
        RECT 99.530 274.400 103.530 274.600 ;
        RECT 103.130 273.800 103.530 274.400 ;
        RECT 99.530 273.600 103.530 273.800 ;
        RECT 103.130 273.000 103.530 273.600 ;
        RECT 99.530 272.800 103.530 273.000 ;
        RECT 103.130 272.200 103.530 272.800 ;
        RECT 99.530 272.000 103.530 272.200 ;
        RECT 103.130 271.400 103.530 272.000 ;
        RECT 99.530 271.200 103.530 271.400 ;
        RECT 103.130 270.600 103.530 271.200 ;
        RECT 99.530 270.400 103.530 270.600 ;
        RECT 103.130 270.200 103.530 270.400 ;
        RECT 95.380 269.800 103.530 270.200 ;
        RECT 110.050 270.015 110.410 270.395 ;
        RECT 110.680 270.015 111.040 270.395 ;
        RECT 111.280 270.015 111.640 270.395 ;
        RECT 95.380 262.200 95.580 269.800 ;
        RECT 96.180 262.200 96.380 269.800 ;
        RECT 96.980 262.200 97.180 269.800 ;
        RECT 97.780 262.200 97.980 269.800 ;
        RECT 98.580 262.200 98.780 269.800 ;
        RECT 103.130 269.600 103.530 269.800 ;
        RECT 99.530 269.400 103.530 269.600 ;
        RECT 110.050 269.425 110.410 269.805 ;
        RECT 110.680 269.425 111.040 269.805 ;
        RECT 111.280 269.425 111.640 269.805 ;
        RECT 103.130 268.800 103.530 269.400 ;
        RECT 99.530 268.600 103.530 268.800 ;
        RECT 103.130 268.000 103.530 268.600 ;
        RECT 99.530 267.800 103.530 268.000 ;
        RECT 103.130 267.200 103.530 267.800 ;
        RECT 99.530 267.000 103.530 267.200 ;
        RECT 103.130 266.400 103.530 267.000 ;
        RECT 99.530 266.200 103.530 266.400 ;
        RECT 103.130 265.600 103.530 266.200 ;
        RECT 99.530 265.400 103.530 265.600 ;
        RECT 103.130 264.800 103.530 265.400 ;
        RECT 99.530 264.600 103.530 264.800 ;
        RECT 103.130 264.000 103.530 264.600 ;
        RECT 99.530 263.800 103.530 264.000 ;
        RECT 103.130 263.200 103.530 263.800 ;
        RECT 99.530 263.000 103.530 263.200 ;
        RECT 103.130 262.400 103.530 263.000 ;
        RECT 99.530 262.200 103.530 262.400 ;
        RECT 5.930 257.600 9.930 257.800 ;
        RECT 5.930 257.000 6.330 257.600 ;
        RECT 5.930 256.800 9.930 257.000 ;
        RECT 5.930 256.200 6.330 256.800 ;
        RECT 5.930 256.000 9.930 256.200 ;
        RECT 5.930 255.400 6.330 256.000 ;
        RECT 5.930 255.200 9.930 255.400 ;
        RECT 5.930 254.600 6.330 255.200 ;
        RECT 5.930 254.400 9.930 254.600 ;
        RECT 5.930 253.800 6.330 254.400 ;
        RECT 5.930 253.600 9.930 253.800 ;
        RECT 5.930 253.000 6.330 253.600 ;
        RECT 5.930 252.800 9.930 253.000 ;
        RECT 5.930 252.200 6.330 252.800 ;
        RECT 5.930 252.000 9.930 252.200 ;
        RECT 5.930 251.400 6.330 252.000 ;
        RECT 5.930 251.200 9.930 251.400 ;
        RECT 5.930 250.600 6.330 251.200 ;
        RECT 5.930 250.400 9.930 250.600 ;
        RECT 5.930 250.200 6.330 250.400 ;
        RECT 10.680 250.200 10.880 257.800 ;
        RECT 11.480 250.200 11.680 257.800 ;
        RECT 12.280 250.200 12.480 257.800 ;
        RECT 13.080 250.200 13.280 257.800 ;
        RECT 13.880 250.200 14.080 257.800 ;
        RECT 5.930 249.800 14.080 250.200 ;
        RECT 5.930 249.600 6.330 249.800 ;
        RECT 5.930 249.400 9.930 249.600 ;
        RECT 5.930 248.800 6.330 249.400 ;
        RECT 5.930 248.600 9.930 248.800 ;
        RECT 5.930 248.000 6.330 248.600 ;
        RECT 5.930 247.800 9.930 248.000 ;
        RECT 5.930 247.200 6.330 247.800 ;
        RECT 5.930 247.000 9.930 247.200 ;
        RECT 5.930 246.400 6.330 247.000 ;
        RECT 5.930 246.200 9.930 246.400 ;
        RECT 5.930 245.600 6.330 246.200 ;
        RECT 5.930 245.400 9.930 245.600 ;
        RECT 5.930 244.800 6.330 245.400 ;
        RECT 5.930 244.600 9.930 244.800 ;
        RECT 5.930 244.000 6.330 244.600 ;
        RECT 5.930 243.800 9.930 244.000 ;
        RECT 5.930 243.200 6.330 243.800 ;
        RECT 5.930 243.000 9.930 243.200 ;
        RECT 5.930 242.400 6.330 243.000 ;
        RECT 5.930 242.200 9.930 242.400 ;
        RECT 10.680 242.200 10.880 249.800 ;
        RECT 11.480 242.200 11.680 249.800 ;
        RECT 12.280 242.200 12.480 249.800 ;
        RECT 13.080 242.200 13.280 249.800 ;
        RECT 13.880 242.200 14.080 249.800 ;
        RECT 15.380 250.200 15.580 257.800 ;
        RECT 16.180 250.200 16.380 257.800 ;
        RECT 16.980 250.200 17.180 257.800 ;
        RECT 17.780 250.200 17.980 257.800 ;
        RECT 18.580 250.200 18.780 257.800 ;
        RECT 19.530 257.600 23.530 257.800 ;
        RECT 23.130 257.000 23.530 257.600 ;
        RECT 19.530 256.800 23.530 257.000 ;
        RECT 23.130 256.200 23.530 256.800 ;
        RECT 19.530 256.000 23.530 256.200 ;
        RECT 23.130 255.400 23.530 256.000 ;
        RECT 19.530 255.200 23.530 255.400 ;
        RECT 23.130 254.600 23.530 255.200 ;
        RECT 19.530 254.400 23.530 254.600 ;
        RECT 23.130 253.800 23.530 254.400 ;
        RECT 19.530 253.600 23.530 253.800 ;
        RECT 23.130 253.000 23.530 253.600 ;
        RECT 19.530 252.800 23.530 253.000 ;
        RECT 23.130 252.200 23.530 252.800 ;
        RECT 19.530 252.000 23.530 252.200 ;
        RECT 23.130 251.400 23.530 252.000 ;
        RECT 19.530 251.200 23.530 251.400 ;
        RECT 23.130 250.600 23.530 251.200 ;
        RECT 19.530 250.400 23.530 250.600 ;
        RECT 23.130 250.200 23.530 250.400 ;
        RECT 15.380 249.800 23.530 250.200 ;
        RECT 15.380 242.200 15.580 249.800 ;
        RECT 16.180 242.200 16.380 249.800 ;
        RECT 16.980 242.200 17.180 249.800 ;
        RECT 17.780 242.200 17.980 249.800 ;
        RECT 18.580 242.200 18.780 249.800 ;
        RECT 23.130 249.600 23.530 249.800 ;
        RECT 19.530 249.400 23.530 249.600 ;
        RECT 23.130 248.800 23.530 249.400 ;
        RECT 19.530 248.600 23.530 248.800 ;
        RECT 23.130 248.000 23.530 248.600 ;
        RECT 19.530 247.800 23.530 248.000 ;
        RECT 23.130 247.200 23.530 247.800 ;
        RECT 19.530 247.000 23.530 247.200 ;
        RECT 23.130 246.400 23.530 247.000 ;
        RECT 19.530 246.200 23.530 246.400 ;
        RECT 23.130 245.600 23.530 246.200 ;
        RECT 19.530 245.400 23.530 245.600 ;
        RECT 23.130 244.800 23.530 245.400 ;
        RECT 19.530 244.600 23.530 244.800 ;
        RECT 23.130 244.000 23.530 244.600 ;
        RECT 19.530 243.800 23.530 244.000 ;
        RECT 23.130 243.200 23.530 243.800 ;
        RECT 19.530 243.000 23.530 243.200 ;
        RECT 23.130 242.400 23.530 243.000 ;
        RECT 19.530 242.200 23.530 242.400 ;
        RECT 25.930 257.600 29.930 257.800 ;
        RECT 25.930 257.000 26.330 257.600 ;
        RECT 25.930 256.800 29.930 257.000 ;
        RECT 25.930 256.200 26.330 256.800 ;
        RECT 25.930 256.000 29.930 256.200 ;
        RECT 25.930 255.400 26.330 256.000 ;
        RECT 25.930 255.200 29.930 255.400 ;
        RECT 25.930 254.600 26.330 255.200 ;
        RECT 25.930 254.400 29.930 254.600 ;
        RECT 25.930 253.800 26.330 254.400 ;
        RECT 25.930 253.600 29.930 253.800 ;
        RECT 25.930 253.000 26.330 253.600 ;
        RECT 25.930 252.800 29.930 253.000 ;
        RECT 25.930 252.200 26.330 252.800 ;
        RECT 25.930 252.000 29.930 252.200 ;
        RECT 25.930 251.400 26.330 252.000 ;
        RECT 25.930 251.200 29.930 251.400 ;
        RECT 25.930 250.600 26.330 251.200 ;
        RECT 25.930 250.400 29.930 250.600 ;
        RECT 25.930 250.200 26.330 250.400 ;
        RECT 30.680 250.200 30.880 257.800 ;
        RECT 31.480 250.200 31.680 257.800 ;
        RECT 32.280 250.200 32.480 257.800 ;
        RECT 33.080 250.200 33.280 257.800 ;
        RECT 33.880 250.200 34.080 257.800 ;
        RECT 25.930 249.800 34.080 250.200 ;
        RECT 25.930 249.600 26.330 249.800 ;
        RECT 25.930 249.400 29.930 249.600 ;
        RECT 25.930 248.800 26.330 249.400 ;
        RECT 25.930 248.600 29.930 248.800 ;
        RECT 25.930 248.000 26.330 248.600 ;
        RECT 25.930 247.800 29.930 248.000 ;
        RECT 25.930 247.200 26.330 247.800 ;
        RECT 25.930 247.000 29.930 247.200 ;
        RECT 25.930 246.400 26.330 247.000 ;
        RECT 25.930 246.200 29.930 246.400 ;
        RECT 25.930 245.600 26.330 246.200 ;
        RECT 25.930 245.400 29.930 245.600 ;
        RECT 25.930 244.800 26.330 245.400 ;
        RECT 25.930 244.600 29.930 244.800 ;
        RECT 25.930 244.000 26.330 244.600 ;
        RECT 25.930 243.800 29.930 244.000 ;
        RECT 25.930 243.200 26.330 243.800 ;
        RECT 25.930 243.000 29.930 243.200 ;
        RECT 25.930 242.400 26.330 243.000 ;
        RECT 25.930 242.200 29.930 242.400 ;
        RECT 30.680 242.200 30.880 249.800 ;
        RECT 31.480 242.200 31.680 249.800 ;
        RECT 32.280 242.200 32.480 249.800 ;
        RECT 33.080 242.200 33.280 249.800 ;
        RECT 33.880 242.200 34.080 249.800 ;
        RECT 35.380 250.200 35.580 257.800 ;
        RECT 36.180 250.200 36.380 257.800 ;
        RECT 36.980 250.200 37.180 257.800 ;
        RECT 37.780 250.200 37.980 257.800 ;
        RECT 38.580 250.200 38.780 257.800 ;
        RECT 39.530 257.600 43.530 257.800 ;
        RECT 43.130 257.000 43.530 257.600 ;
        RECT 39.530 256.800 43.530 257.000 ;
        RECT 43.130 256.200 43.530 256.800 ;
        RECT 39.530 256.000 43.530 256.200 ;
        RECT 43.130 255.400 43.530 256.000 ;
        RECT 39.530 255.200 43.530 255.400 ;
        RECT 43.130 254.600 43.530 255.200 ;
        RECT 39.530 254.400 43.530 254.600 ;
        RECT 43.130 253.800 43.530 254.400 ;
        RECT 39.530 253.600 43.530 253.800 ;
        RECT 43.130 253.000 43.530 253.600 ;
        RECT 39.530 252.800 43.530 253.000 ;
        RECT 43.130 252.200 43.530 252.800 ;
        RECT 39.530 252.000 43.530 252.200 ;
        RECT 43.130 251.400 43.530 252.000 ;
        RECT 39.530 251.200 43.530 251.400 ;
        RECT 43.130 250.600 43.530 251.200 ;
        RECT 39.530 250.400 43.530 250.600 ;
        RECT 43.130 250.200 43.530 250.400 ;
        RECT 35.380 249.800 43.530 250.200 ;
        RECT 35.380 242.200 35.580 249.800 ;
        RECT 36.180 242.200 36.380 249.800 ;
        RECT 36.980 242.200 37.180 249.800 ;
        RECT 37.780 242.200 37.980 249.800 ;
        RECT 38.580 242.200 38.780 249.800 ;
        RECT 43.130 249.600 43.530 249.800 ;
        RECT 39.530 249.400 43.530 249.600 ;
        RECT 43.130 248.800 43.530 249.400 ;
        RECT 39.530 248.600 43.530 248.800 ;
        RECT 43.130 248.000 43.530 248.600 ;
        RECT 39.530 247.800 43.530 248.000 ;
        RECT 43.130 247.200 43.530 247.800 ;
        RECT 39.530 247.000 43.530 247.200 ;
        RECT 43.130 246.400 43.530 247.000 ;
        RECT 39.530 246.200 43.530 246.400 ;
        RECT 43.130 245.600 43.530 246.200 ;
        RECT 39.530 245.400 43.530 245.600 ;
        RECT 43.130 244.800 43.530 245.400 ;
        RECT 39.530 244.600 43.530 244.800 ;
        RECT 43.130 244.000 43.530 244.600 ;
        RECT 39.530 243.800 43.530 244.000 ;
        RECT 43.130 243.200 43.530 243.800 ;
        RECT 39.530 243.000 43.530 243.200 ;
        RECT 43.130 242.400 43.530 243.000 ;
        RECT 39.530 242.200 43.530 242.400 ;
        RECT 45.930 257.600 49.930 257.800 ;
        RECT 45.930 257.000 46.330 257.600 ;
        RECT 45.930 256.800 49.930 257.000 ;
        RECT 45.930 256.200 46.330 256.800 ;
        RECT 45.930 256.000 49.930 256.200 ;
        RECT 45.930 255.400 46.330 256.000 ;
        RECT 45.930 255.200 49.930 255.400 ;
        RECT 45.930 254.600 46.330 255.200 ;
        RECT 45.930 254.400 49.930 254.600 ;
        RECT 45.930 253.800 46.330 254.400 ;
        RECT 45.930 253.600 49.930 253.800 ;
        RECT 45.930 253.000 46.330 253.600 ;
        RECT 45.930 252.800 49.930 253.000 ;
        RECT 45.930 252.200 46.330 252.800 ;
        RECT 45.930 252.000 49.930 252.200 ;
        RECT 45.930 251.400 46.330 252.000 ;
        RECT 45.930 251.200 49.930 251.400 ;
        RECT 45.930 250.600 46.330 251.200 ;
        RECT 45.930 250.400 49.930 250.600 ;
        RECT 45.930 250.200 46.330 250.400 ;
        RECT 50.680 250.200 50.880 257.800 ;
        RECT 51.480 250.200 51.680 257.800 ;
        RECT 52.280 250.200 52.480 257.800 ;
        RECT 53.080 250.200 53.280 257.800 ;
        RECT 53.880 250.200 54.080 257.800 ;
        RECT 45.930 249.800 54.080 250.200 ;
        RECT 45.930 249.600 46.330 249.800 ;
        RECT 45.930 249.400 49.930 249.600 ;
        RECT 45.930 248.800 46.330 249.400 ;
        RECT 45.930 248.600 49.930 248.800 ;
        RECT 45.930 248.000 46.330 248.600 ;
        RECT 45.930 247.800 49.930 248.000 ;
        RECT 45.930 247.200 46.330 247.800 ;
        RECT 45.930 247.000 49.930 247.200 ;
        RECT 45.930 246.400 46.330 247.000 ;
        RECT 45.930 246.200 49.930 246.400 ;
        RECT 45.930 245.600 46.330 246.200 ;
        RECT 45.930 245.400 49.930 245.600 ;
        RECT 45.930 244.800 46.330 245.400 ;
        RECT 45.930 244.600 49.930 244.800 ;
        RECT 45.930 244.000 46.330 244.600 ;
        RECT 45.930 243.800 49.930 244.000 ;
        RECT 45.930 243.200 46.330 243.800 ;
        RECT 45.930 243.000 49.930 243.200 ;
        RECT 45.930 242.400 46.330 243.000 ;
        RECT 45.930 242.200 49.930 242.400 ;
        RECT 50.680 242.200 50.880 249.800 ;
        RECT 51.480 242.200 51.680 249.800 ;
        RECT 52.280 242.200 52.480 249.800 ;
        RECT 53.080 242.200 53.280 249.800 ;
        RECT 53.880 242.200 54.080 249.800 ;
        RECT 55.380 250.200 55.580 257.800 ;
        RECT 56.180 250.200 56.380 257.800 ;
        RECT 56.980 250.200 57.180 257.800 ;
        RECT 57.780 250.200 57.980 257.800 ;
        RECT 58.580 250.200 58.780 257.800 ;
        RECT 59.530 257.600 63.530 257.800 ;
        RECT 63.130 257.000 63.530 257.600 ;
        RECT 59.530 256.800 63.530 257.000 ;
        RECT 63.130 256.200 63.530 256.800 ;
        RECT 59.530 256.000 63.530 256.200 ;
        RECT 63.130 255.400 63.530 256.000 ;
        RECT 59.530 255.200 63.530 255.400 ;
        RECT 63.130 254.600 63.530 255.200 ;
        RECT 59.530 254.400 63.530 254.600 ;
        RECT 63.130 253.800 63.530 254.400 ;
        RECT 59.530 253.600 63.530 253.800 ;
        RECT 63.130 253.000 63.530 253.600 ;
        RECT 59.530 252.800 63.530 253.000 ;
        RECT 63.130 252.200 63.530 252.800 ;
        RECT 59.530 252.000 63.530 252.200 ;
        RECT 63.130 251.400 63.530 252.000 ;
        RECT 59.530 251.200 63.530 251.400 ;
        RECT 63.130 250.600 63.530 251.200 ;
        RECT 59.530 250.400 63.530 250.600 ;
        RECT 63.130 250.200 63.530 250.400 ;
        RECT 55.380 249.800 63.530 250.200 ;
        RECT 55.380 242.200 55.580 249.800 ;
        RECT 56.180 242.200 56.380 249.800 ;
        RECT 56.980 242.200 57.180 249.800 ;
        RECT 57.780 242.200 57.980 249.800 ;
        RECT 58.580 242.200 58.780 249.800 ;
        RECT 63.130 249.600 63.530 249.800 ;
        RECT 59.530 249.400 63.530 249.600 ;
        RECT 63.130 248.800 63.530 249.400 ;
        RECT 59.530 248.600 63.530 248.800 ;
        RECT 63.130 248.000 63.530 248.600 ;
        RECT 59.530 247.800 63.530 248.000 ;
        RECT 63.130 247.200 63.530 247.800 ;
        RECT 59.530 247.000 63.530 247.200 ;
        RECT 63.130 246.400 63.530 247.000 ;
        RECT 59.530 246.200 63.530 246.400 ;
        RECT 63.130 245.600 63.530 246.200 ;
        RECT 59.530 245.400 63.530 245.600 ;
        RECT 63.130 244.800 63.530 245.400 ;
        RECT 59.530 244.600 63.530 244.800 ;
        RECT 63.130 244.000 63.530 244.600 ;
        RECT 59.530 243.800 63.530 244.000 ;
        RECT 63.130 243.200 63.530 243.800 ;
        RECT 59.530 243.000 63.530 243.200 ;
        RECT 63.130 242.400 63.530 243.000 ;
        RECT 59.530 242.200 63.530 242.400 ;
        RECT 65.930 257.600 69.930 257.800 ;
        RECT 65.930 257.000 66.330 257.600 ;
        RECT 65.930 256.800 69.930 257.000 ;
        RECT 65.930 256.200 66.330 256.800 ;
        RECT 65.930 256.000 69.930 256.200 ;
        RECT 65.930 255.400 66.330 256.000 ;
        RECT 65.930 255.200 69.930 255.400 ;
        RECT 65.930 254.600 66.330 255.200 ;
        RECT 65.930 254.400 69.930 254.600 ;
        RECT 65.930 253.800 66.330 254.400 ;
        RECT 65.930 253.600 69.930 253.800 ;
        RECT 65.930 253.000 66.330 253.600 ;
        RECT 65.930 252.800 69.930 253.000 ;
        RECT 65.930 252.200 66.330 252.800 ;
        RECT 65.930 252.000 69.930 252.200 ;
        RECT 65.930 251.400 66.330 252.000 ;
        RECT 65.930 251.200 69.930 251.400 ;
        RECT 65.930 250.600 66.330 251.200 ;
        RECT 65.930 250.400 69.930 250.600 ;
        RECT 65.930 250.200 66.330 250.400 ;
        RECT 70.680 250.200 70.880 257.800 ;
        RECT 71.480 250.200 71.680 257.800 ;
        RECT 72.280 250.200 72.480 257.800 ;
        RECT 73.080 250.200 73.280 257.800 ;
        RECT 73.880 250.200 74.080 257.800 ;
        RECT 65.930 249.800 74.080 250.200 ;
        RECT 65.930 249.600 66.330 249.800 ;
        RECT 65.930 249.400 69.930 249.600 ;
        RECT 65.930 248.800 66.330 249.400 ;
        RECT 65.930 248.600 69.930 248.800 ;
        RECT 65.930 248.000 66.330 248.600 ;
        RECT 65.930 247.800 69.930 248.000 ;
        RECT 65.930 247.200 66.330 247.800 ;
        RECT 65.930 247.000 69.930 247.200 ;
        RECT 65.930 246.400 66.330 247.000 ;
        RECT 65.930 246.200 69.930 246.400 ;
        RECT 65.930 245.600 66.330 246.200 ;
        RECT 65.930 245.400 69.930 245.600 ;
        RECT 65.930 244.800 66.330 245.400 ;
        RECT 65.930 244.600 69.930 244.800 ;
        RECT 65.930 244.000 66.330 244.600 ;
        RECT 65.930 243.800 69.930 244.000 ;
        RECT 65.930 243.200 66.330 243.800 ;
        RECT 65.930 243.000 69.930 243.200 ;
        RECT 65.930 242.400 66.330 243.000 ;
        RECT 65.930 242.200 69.930 242.400 ;
        RECT 70.680 242.200 70.880 249.800 ;
        RECT 71.480 242.200 71.680 249.800 ;
        RECT 72.280 242.200 72.480 249.800 ;
        RECT 73.080 242.200 73.280 249.800 ;
        RECT 73.880 242.200 74.080 249.800 ;
        RECT 75.380 250.200 75.580 257.800 ;
        RECT 76.180 250.200 76.380 257.800 ;
        RECT 76.980 250.200 77.180 257.800 ;
        RECT 77.780 250.200 77.980 257.800 ;
        RECT 78.580 250.200 78.780 257.800 ;
        RECT 79.530 257.600 83.530 257.800 ;
        RECT 83.130 257.000 83.530 257.600 ;
        RECT 79.530 256.800 83.530 257.000 ;
        RECT 83.130 256.200 83.530 256.800 ;
        RECT 79.530 256.000 83.530 256.200 ;
        RECT 83.130 255.400 83.530 256.000 ;
        RECT 79.530 255.200 83.530 255.400 ;
        RECT 83.130 254.600 83.530 255.200 ;
        RECT 79.530 254.400 83.530 254.600 ;
        RECT 83.130 253.800 83.530 254.400 ;
        RECT 79.530 253.600 83.530 253.800 ;
        RECT 83.130 253.000 83.530 253.600 ;
        RECT 79.530 252.800 83.530 253.000 ;
        RECT 83.130 252.200 83.530 252.800 ;
        RECT 79.530 252.000 83.530 252.200 ;
        RECT 83.130 251.400 83.530 252.000 ;
        RECT 79.530 251.200 83.530 251.400 ;
        RECT 83.130 250.600 83.530 251.200 ;
        RECT 79.530 250.400 83.530 250.600 ;
        RECT 83.130 250.200 83.530 250.400 ;
        RECT 75.380 249.800 83.530 250.200 ;
        RECT 75.380 242.200 75.580 249.800 ;
        RECT 76.180 242.200 76.380 249.800 ;
        RECT 76.980 242.200 77.180 249.800 ;
        RECT 77.780 242.200 77.980 249.800 ;
        RECT 78.580 242.200 78.780 249.800 ;
        RECT 83.130 249.600 83.530 249.800 ;
        RECT 79.530 249.400 83.530 249.600 ;
        RECT 83.130 248.800 83.530 249.400 ;
        RECT 79.530 248.600 83.530 248.800 ;
        RECT 83.130 248.000 83.530 248.600 ;
        RECT 79.530 247.800 83.530 248.000 ;
        RECT 83.130 247.200 83.530 247.800 ;
        RECT 79.530 247.000 83.530 247.200 ;
        RECT 83.130 246.400 83.530 247.000 ;
        RECT 79.530 246.200 83.530 246.400 ;
        RECT 83.130 245.600 83.530 246.200 ;
        RECT 79.530 245.400 83.530 245.600 ;
        RECT 83.130 244.800 83.530 245.400 ;
        RECT 79.530 244.600 83.530 244.800 ;
        RECT 83.130 244.000 83.530 244.600 ;
        RECT 79.530 243.800 83.530 244.000 ;
        RECT 83.130 243.200 83.530 243.800 ;
        RECT 79.530 243.000 83.530 243.200 ;
        RECT 83.130 242.400 83.530 243.000 ;
        RECT 79.530 242.200 83.530 242.400 ;
        RECT 85.930 257.600 89.930 257.800 ;
        RECT 85.930 257.000 86.330 257.600 ;
        RECT 85.930 256.800 89.930 257.000 ;
        RECT 85.930 256.200 86.330 256.800 ;
        RECT 85.930 256.000 89.930 256.200 ;
        RECT 85.930 255.400 86.330 256.000 ;
        RECT 85.930 255.200 89.930 255.400 ;
        RECT 85.930 254.600 86.330 255.200 ;
        RECT 85.930 254.400 89.930 254.600 ;
        RECT 85.930 253.800 86.330 254.400 ;
        RECT 85.930 253.600 89.930 253.800 ;
        RECT 85.930 253.000 86.330 253.600 ;
        RECT 85.930 252.800 89.930 253.000 ;
        RECT 85.930 252.200 86.330 252.800 ;
        RECT 85.930 252.000 89.930 252.200 ;
        RECT 85.930 251.400 86.330 252.000 ;
        RECT 85.930 251.200 89.930 251.400 ;
        RECT 85.930 250.600 86.330 251.200 ;
        RECT 85.930 250.400 89.930 250.600 ;
        RECT 85.930 250.200 86.330 250.400 ;
        RECT 90.680 250.200 90.880 257.800 ;
        RECT 91.480 250.200 91.680 257.800 ;
        RECT 92.280 250.200 92.480 257.800 ;
        RECT 93.080 250.200 93.280 257.800 ;
        RECT 93.880 250.200 94.080 257.800 ;
        RECT 85.930 249.800 94.080 250.200 ;
        RECT 85.930 249.600 86.330 249.800 ;
        RECT 85.930 249.400 89.930 249.600 ;
        RECT 85.930 248.800 86.330 249.400 ;
        RECT 85.930 248.600 89.930 248.800 ;
        RECT 85.930 248.000 86.330 248.600 ;
        RECT 85.930 247.800 89.930 248.000 ;
        RECT 85.930 247.200 86.330 247.800 ;
        RECT 85.930 247.000 89.930 247.200 ;
        RECT 85.930 246.400 86.330 247.000 ;
        RECT 85.930 246.200 89.930 246.400 ;
        RECT 85.930 245.600 86.330 246.200 ;
        RECT 85.930 245.400 89.930 245.600 ;
        RECT 85.930 244.800 86.330 245.400 ;
        RECT 85.930 244.600 89.930 244.800 ;
        RECT 85.930 244.000 86.330 244.600 ;
        RECT 85.930 243.800 89.930 244.000 ;
        RECT 85.930 243.200 86.330 243.800 ;
        RECT 85.930 243.000 89.930 243.200 ;
        RECT 85.930 242.400 86.330 243.000 ;
        RECT 85.930 242.200 89.930 242.400 ;
        RECT 90.680 242.200 90.880 249.800 ;
        RECT 91.480 242.200 91.680 249.800 ;
        RECT 92.280 242.200 92.480 249.800 ;
        RECT 93.080 242.200 93.280 249.800 ;
        RECT 93.880 242.200 94.080 249.800 ;
        RECT 95.380 250.200 95.580 257.800 ;
        RECT 96.180 250.200 96.380 257.800 ;
        RECT 96.980 250.200 97.180 257.800 ;
        RECT 97.780 250.200 97.980 257.800 ;
        RECT 98.580 250.200 98.780 257.800 ;
        RECT 99.530 257.600 103.530 257.800 ;
        RECT 103.130 257.000 103.530 257.600 ;
        RECT 99.530 256.800 103.530 257.000 ;
        RECT 103.130 256.200 103.530 256.800 ;
        RECT 99.530 256.000 103.530 256.200 ;
        RECT 103.130 255.400 103.530 256.000 ;
        RECT 99.530 255.200 103.530 255.400 ;
        RECT 103.130 254.600 103.530 255.200 ;
        RECT 99.530 254.400 103.530 254.600 ;
        RECT 103.130 253.800 103.530 254.400 ;
        RECT 99.530 253.600 103.530 253.800 ;
        RECT 103.130 253.000 103.530 253.600 ;
        RECT 99.530 252.800 103.530 253.000 ;
        RECT 103.130 252.200 103.530 252.800 ;
        RECT 99.530 252.000 103.530 252.200 ;
        RECT 103.130 251.400 103.530 252.000 ;
        RECT 99.530 251.200 103.530 251.400 ;
        RECT 103.130 250.600 103.530 251.200 ;
        RECT 99.530 250.400 103.530 250.600 ;
        RECT 110.050 250.410 110.410 250.790 ;
        RECT 110.680 250.410 111.040 250.790 ;
        RECT 111.280 250.410 111.640 250.790 ;
        RECT 103.130 250.200 103.530 250.400 ;
        RECT 95.380 249.800 103.530 250.200 ;
        RECT 110.050 249.820 110.410 250.200 ;
        RECT 110.680 249.820 111.040 250.200 ;
        RECT 111.280 249.820 111.640 250.200 ;
        RECT 95.380 242.200 95.580 249.800 ;
        RECT 96.180 242.200 96.380 249.800 ;
        RECT 96.980 242.200 97.180 249.800 ;
        RECT 97.780 242.200 97.980 249.800 ;
        RECT 98.580 242.200 98.780 249.800 ;
        RECT 103.130 249.600 103.530 249.800 ;
        RECT 99.530 249.400 103.530 249.600 ;
        RECT 103.130 248.800 103.530 249.400 ;
        RECT 99.530 248.600 103.530 248.800 ;
        RECT 103.130 248.000 103.530 248.600 ;
        RECT 99.530 247.800 103.530 248.000 ;
        RECT 103.130 247.200 103.530 247.800 ;
        RECT 99.530 247.000 103.530 247.200 ;
        RECT 103.130 246.400 103.530 247.000 ;
        RECT 99.530 246.200 103.530 246.400 ;
        RECT 103.130 245.600 103.530 246.200 ;
        RECT 99.530 245.400 103.530 245.600 ;
        RECT 103.130 244.800 103.530 245.400 ;
        RECT 99.530 244.600 103.530 244.800 ;
        RECT 103.130 244.000 103.530 244.600 ;
        RECT 99.530 243.800 103.530 244.000 ;
        RECT 103.130 243.200 103.530 243.800 ;
        RECT 99.530 243.000 103.530 243.200 ;
        RECT 103.130 242.400 103.530 243.000 ;
        RECT 99.530 242.200 103.530 242.400 ;
        RECT 5.930 237.600 9.930 237.800 ;
        RECT 5.930 237.000 6.330 237.600 ;
        RECT 5.930 236.800 9.930 237.000 ;
        RECT 5.930 236.200 6.330 236.800 ;
        RECT 5.930 236.000 9.930 236.200 ;
        RECT 5.930 235.400 6.330 236.000 ;
        RECT 5.930 235.200 9.930 235.400 ;
        RECT 5.930 234.600 6.330 235.200 ;
        RECT 5.930 234.400 9.930 234.600 ;
        RECT 5.930 233.800 6.330 234.400 ;
        RECT 5.930 233.600 9.930 233.800 ;
        RECT 5.930 233.000 6.330 233.600 ;
        RECT 5.930 232.800 9.930 233.000 ;
        RECT 5.930 232.200 6.330 232.800 ;
        RECT 5.930 232.000 9.930 232.200 ;
        RECT 5.930 231.400 6.330 232.000 ;
        RECT 5.930 231.200 9.930 231.400 ;
        RECT 5.930 230.600 6.330 231.200 ;
        RECT 5.930 230.400 9.930 230.600 ;
        RECT 5.930 230.200 6.330 230.400 ;
        RECT 10.680 230.200 10.880 237.800 ;
        RECT 11.480 230.200 11.680 237.800 ;
        RECT 12.280 230.200 12.480 237.800 ;
        RECT 13.080 230.200 13.280 237.800 ;
        RECT 13.880 230.200 14.080 237.800 ;
        RECT 5.930 229.800 14.080 230.200 ;
        RECT 5.930 229.600 6.330 229.800 ;
        RECT 5.930 229.400 9.930 229.600 ;
        RECT 5.930 228.800 6.330 229.400 ;
        RECT 5.930 228.600 9.930 228.800 ;
        RECT 5.930 228.000 6.330 228.600 ;
        RECT 5.930 227.800 9.930 228.000 ;
        RECT 5.930 227.200 6.330 227.800 ;
        RECT 5.930 227.000 9.930 227.200 ;
        RECT 5.930 226.400 6.330 227.000 ;
        RECT 5.930 226.200 9.930 226.400 ;
        RECT 5.930 225.600 6.330 226.200 ;
        RECT 5.930 225.400 9.930 225.600 ;
        RECT 5.930 224.800 6.330 225.400 ;
        RECT 5.930 224.600 9.930 224.800 ;
        RECT 5.930 224.000 6.330 224.600 ;
        RECT 5.930 223.800 9.930 224.000 ;
        RECT 5.930 223.200 6.330 223.800 ;
        RECT 5.930 223.000 9.930 223.200 ;
        RECT 5.930 222.400 6.330 223.000 ;
        RECT 5.930 222.200 9.930 222.400 ;
        RECT 10.680 222.200 10.880 229.800 ;
        RECT 11.480 222.200 11.680 229.800 ;
        RECT 12.280 222.200 12.480 229.800 ;
        RECT 13.080 222.200 13.280 229.800 ;
        RECT 13.880 222.200 14.080 229.800 ;
        RECT 15.380 230.200 15.580 237.800 ;
        RECT 16.180 230.200 16.380 237.800 ;
        RECT 16.980 230.200 17.180 237.800 ;
        RECT 17.780 230.200 17.980 237.800 ;
        RECT 18.580 230.200 18.780 237.800 ;
        RECT 19.530 237.600 23.530 237.800 ;
        RECT 23.130 237.000 23.530 237.600 ;
        RECT 19.530 236.800 23.530 237.000 ;
        RECT 23.130 236.200 23.530 236.800 ;
        RECT 19.530 236.000 23.530 236.200 ;
        RECT 23.130 235.400 23.530 236.000 ;
        RECT 19.530 235.200 23.530 235.400 ;
        RECT 23.130 234.600 23.530 235.200 ;
        RECT 19.530 234.400 23.530 234.600 ;
        RECT 23.130 233.800 23.530 234.400 ;
        RECT 19.530 233.600 23.530 233.800 ;
        RECT 23.130 233.000 23.530 233.600 ;
        RECT 19.530 232.800 23.530 233.000 ;
        RECT 23.130 232.200 23.530 232.800 ;
        RECT 19.530 232.000 23.530 232.200 ;
        RECT 23.130 231.400 23.530 232.000 ;
        RECT 19.530 231.200 23.530 231.400 ;
        RECT 23.130 230.600 23.530 231.200 ;
        RECT 19.530 230.400 23.530 230.600 ;
        RECT 23.130 230.200 23.530 230.400 ;
        RECT 15.380 229.800 23.530 230.200 ;
        RECT 15.380 222.200 15.580 229.800 ;
        RECT 16.180 222.200 16.380 229.800 ;
        RECT 16.980 222.200 17.180 229.800 ;
        RECT 17.780 222.200 17.980 229.800 ;
        RECT 18.580 222.200 18.780 229.800 ;
        RECT 23.130 229.600 23.530 229.800 ;
        RECT 19.530 229.400 23.530 229.600 ;
        RECT 23.130 228.800 23.530 229.400 ;
        RECT 19.530 228.600 23.530 228.800 ;
        RECT 23.130 228.000 23.530 228.600 ;
        RECT 19.530 227.800 23.530 228.000 ;
        RECT 23.130 227.200 23.530 227.800 ;
        RECT 19.530 227.000 23.530 227.200 ;
        RECT 23.130 226.400 23.530 227.000 ;
        RECT 19.530 226.200 23.530 226.400 ;
        RECT 23.130 225.600 23.530 226.200 ;
        RECT 19.530 225.400 23.530 225.600 ;
        RECT 23.130 224.800 23.530 225.400 ;
        RECT 19.530 224.600 23.530 224.800 ;
        RECT 23.130 224.000 23.530 224.600 ;
        RECT 19.530 223.800 23.530 224.000 ;
        RECT 23.130 223.200 23.530 223.800 ;
        RECT 19.530 223.000 23.530 223.200 ;
        RECT 23.130 222.400 23.530 223.000 ;
        RECT 19.530 222.200 23.530 222.400 ;
        RECT 25.930 237.600 29.930 237.800 ;
        RECT 25.930 237.000 26.330 237.600 ;
        RECT 25.930 236.800 29.930 237.000 ;
        RECT 25.930 236.200 26.330 236.800 ;
        RECT 25.930 236.000 29.930 236.200 ;
        RECT 25.930 235.400 26.330 236.000 ;
        RECT 25.930 235.200 29.930 235.400 ;
        RECT 25.930 234.600 26.330 235.200 ;
        RECT 25.930 234.400 29.930 234.600 ;
        RECT 25.930 233.800 26.330 234.400 ;
        RECT 25.930 233.600 29.930 233.800 ;
        RECT 25.930 233.000 26.330 233.600 ;
        RECT 25.930 232.800 29.930 233.000 ;
        RECT 25.930 232.200 26.330 232.800 ;
        RECT 25.930 232.000 29.930 232.200 ;
        RECT 25.930 231.400 26.330 232.000 ;
        RECT 25.930 231.200 29.930 231.400 ;
        RECT 25.930 230.600 26.330 231.200 ;
        RECT 25.930 230.400 29.930 230.600 ;
        RECT 25.930 230.200 26.330 230.400 ;
        RECT 30.680 230.200 30.880 237.800 ;
        RECT 31.480 230.200 31.680 237.800 ;
        RECT 32.280 230.200 32.480 237.800 ;
        RECT 33.080 230.200 33.280 237.800 ;
        RECT 33.880 230.200 34.080 237.800 ;
        RECT 25.930 229.800 34.080 230.200 ;
        RECT 25.930 229.600 26.330 229.800 ;
        RECT 25.930 229.400 29.930 229.600 ;
        RECT 25.930 228.800 26.330 229.400 ;
        RECT 25.930 228.600 29.930 228.800 ;
        RECT 25.930 228.000 26.330 228.600 ;
        RECT 25.930 227.800 29.930 228.000 ;
        RECT 25.930 227.200 26.330 227.800 ;
        RECT 25.930 227.000 29.930 227.200 ;
        RECT 25.930 226.400 26.330 227.000 ;
        RECT 25.930 226.200 29.930 226.400 ;
        RECT 25.930 225.600 26.330 226.200 ;
        RECT 25.930 225.400 29.930 225.600 ;
        RECT 25.930 224.800 26.330 225.400 ;
        RECT 25.930 224.600 29.930 224.800 ;
        RECT 25.930 224.000 26.330 224.600 ;
        RECT 25.930 223.800 29.930 224.000 ;
        RECT 25.930 223.200 26.330 223.800 ;
        RECT 25.930 223.000 29.930 223.200 ;
        RECT 25.930 222.400 26.330 223.000 ;
        RECT 25.930 222.200 29.930 222.400 ;
        RECT 30.680 222.200 30.880 229.800 ;
        RECT 31.480 222.200 31.680 229.800 ;
        RECT 32.280 222.200 32.480 229.800 ;
        RECT 33.080 222.200 33.280 229.800 ;
        RECT 33.880 222.200 34.080 229.800 ;
        RECT 35.380 230.200 35.580 237.800 ;
        RECT 36.180 230.200 36.380 237.800 ;
        RECT 36.980 230.200 37.180 237.800 ;
        RECT 37.780 230.200 37.980 237.800 ;
        RECT 38.580 230.200 38.780 237.800 ;
        RECT 39.530 237.600 43.530 237.800 ;
        RECT 43.130 237.000 43.530 237.600 ;
        RECT 39.530 236.800 43.530 237.000 ;
        RECT 43.130 236.200 43.530 236.800 ;
        RECT 39.530 236.000 43.530 236.200 ;
        RECT 43.130 235.400 43.530 236.000 ;
        RECT 39.530 235.200 43.530 235.400 ;
        RECT 43.130 234.600 43.530 235.200 ;
        RECT 39.530 234.400 43.530 234.600 ;
        RECT 43.130 233.800 43.530 234.400 ;
        RECT 39.530 233.600 43.530 233.800 ;
        RECT 43.130 233.000 43.530 233.600 ;
        RECT 39.530 232.800 43.530 233.000 ;
        RECT 43.130 232.200 43.530 232.800 ;
        RECT 39.530 232.000 43.530 232.200 ;
        RECT 43.130 231.400 43.530 232.000 ;
        RECT 39.530 231.200 43.530 231.400 ;
        RECT 43.130 230.600 43.530 231.200 ;
        RECT 39.530 230.400 43.530 230.600 ;
        RECT 43.130 230.200 43.530 230.400 ;
        RECT 35.380 229.800 43.530 230.200 ;
        RECT 35.380 222.200 35.580 229.800 ;
        RECT 36.180 222.200 36.380 229.800 ;
        RECT 36.980 222.200 37.180 229.800 ;
        RECT 37.780 222.200 37.980 229.800 ;
        RECT 38.580 222.200 38.780 229.800 ;
        RECT 43.130 229.600 43.530 229.800 ;
        RECT 39.530 229.400 43.530 229.600 ;
        RECT 43.130 228.800 43.530 229.400 ;
        RECT 39.530 228.600 43.530 228.800 ;
        RECT 43.130 228.000 43.530 228.600 ;
        RECT 39.530 227.800 43.530 228.000 ;
        RECT 43.130 227.200 43.530 227.800 ;
        RECT 39.530 227.000 43.530 227.200 ;
        RECT 43.130 226.400 43.530 227.000 ;
        RECT 39.530 226.200 43.530 226.400 ;
        RECT 43.130 225.600 43.530 226.200 ;
        RECT 39.530 225.400 43.530 225.600 ;
        RECT 43.130 224.800 43.530 225.400 ;
        RECT 39.530 224.600 43.530 224.800 ;
        RECT 43.130 224.000 43.530 224.600 ;
        RECT 39.530 223.800 43.530 224.000 ;
        RECT 43.130 223.200 43.530 223.800 ;
        RECT 39.530 223.000 43.530 223.200 ;
        RECT 43.130 222.400 43.530 223.000 ;
        RECT 39.530 222.200 43.530 222.400 ;
        RECT 45.930 237.600 49.930 237.800 ;
        RECT 45.930 237.000 46.330 237.600 ;
        RECT 45.930 236.800 49.930 237.000 ;
        RECT 45.930 236.200 46.330 236.800 ;
        RECT 45.930 236.000 49.930 236.200 ;
        RECT 45.930 235.400 46.330 236.000 ;
        RECT 45.930 235.200 49.930 235.400 ;
        RECT 45.930 234.600 46.330 235.200 ;
        RECT 45.930 234.400 49.930 234.600 ;
        RECT 45.930 233.800 46.330 234.400 ;
        RECT 45.930 233.600 49.930 233.800 ;
        RECT 45.930 233.000 46.330 233.600 ;
        RECT 45.930 232.800 49.930 233.000 ;
        RECT 45.930 232.200 46.330 232.800 ;
        RECT 45.930 232.000 49.930 232.200 ;
        RECT 45.930 231.400 46.330 232.000 ;
        RECT 45.930 231.200 49.930 231.400 ;
        RECT 45.930 230.600 46.330 231.200 ;
        RECT 45.930 230.400 49.930 230.600 ;
        RECT 45.930 230.200 46.330 230.400 ;
        RECT 50.680 230.200 50.880 237.800 ;
        RECT 51.480 230.200 51.680 237.800 ;
        RECT 52.280 230.200 52.480 237.800 ;
        RECT 53.080 230.200 53.280 237.800 ;
        RECT 53.880 230.200 54.080 237.800 ;
        RECT 45.930 229.800 54.080 230.200 ;
        RECT 45.930 229.600 46.330 229.800 ;
        RECT 45.930 229.400 49.930 229.600 ;
        RECT 45.930 228.800 46.330 229.400 ;
        RECT 45.930 228.600 49.930 228.800 ;
        RECT 45.930 228.000 46.330 228.600 ;
        RECT 45.930 227.800 49.930 228.000 ;
        RECT 45.930 227.200 46.330 227.800 ;
        RECT 45.930 227.000 49.930 227.200 ;
        RECT 45.930 226.400 46.330 227.000 ;
        RECT 45.930 226.200 49.930 226.400 ;
        RECT 45.930 225.600 46.330 226.200 ;
        RECT 45.930 225.400 49.930 225.600 ;
        RECT 45.930 224.800 46.330 225.400 ;
        RECT 45.930 224.600 49.930 224.800 ;
        RECT 45.930 224.000 46.330 224.600 ;
        RECT 45.930 223.800 49.930 224.000 ;
        RECT 45.930 223.200 46.330 223.800 ;
        RECT 45.930 223.000 49.930 223.200 ;
        RECT 45.930 222.400 46.330 223.000 ;
        RECT 45.930 222.200 49.930 222.400 ;
        RECT 50.680 222.200 50.880 229.800 ;
        RECT 51.480 222.200 51.680 229.800 ;
        RECT 52.280 222.200 52.480 229.800 ;
        RECT 53.080 222.200 53.280 229.800 ;
        RECT 53.880 222.200 54.080 229.800 ;
        RECT 55.380 230.200 55.580 237.800 ;
        RECT 56.180 230.200 56.380 237.800 ;
        RECT 56.980 230.200 57.180 237.800 ;
        RECT 57.780 230.200 57.980 237.800 ;
        RECT 58.580 230.200 58.780 237.800 ;
        RECT 59.530 237.600 63.530 237.800 ;
        RECT 63.130 237.000 63.530 237.600 ;
        RECT 59.530 236.800 63.530 237.000 ;
        RECT 63.130 236.200 63.530 236.800 ;
        RECT 59.530 236.000 63.530 236.200 ;
        RECT 63.130 235.400 63.530 236.000 ;
        RECT 59.530 235.200 63.530 235.400 ;
        RECT 63.130 234.600 63.530 235.200 ;
        RECT 59.530 234.400 63.530 234.600 ;
        RECT 63.130 233.800 63.530 234.400 ;
        RECT 59.530 233.600 63.530 233.800 ;
        RECT 63.130 233.000 63.530 233.600 ;
        RECT 59.530 232.800 63.530 233.000 ;
        RECT 63.130 232.200 63.530 232.800 ;
        RECT 59.530 232.000 63.530 232.200 ;
        RECT 63.130 231.400 63.530 232.000 ;
        RECT 59.530 231.200 63.530 231.400 ;
        RECT 63.130 230.600 63.530 231.200 ;
        RECT 59.530 230.400 63.530 230.600 ;
        RECT 63.130 230.200 63.530 230.400 ;
        RECT 55.380 229.800 63.530 230.200 ;
        RECT 55.380 222.200 55.580 229.800 ;
        RECT 56.180 222.200 56.380 229.800 ;
        RECT 56.980 222.200 57.180 229.800 ;
        RECT 57.780 222.200 57.980 229.800 ;
        RECT 58.580 222.200 58.780 229.800 ;
        RECT 63.130 229.600 63.530 229.800 ;
        RECT 59.530 229.400 63.530 229.600 ;
        RECT 63.130 228.800 63.530 229.400 ;
        RECT 59.530 228.600 63.530 228.800 ;
        RECT 63.130 228.000 63.530 228.600 ;
        RECT 59.530 227.800 63.530 228.000 ;
        RECT 63.130 227.200 63.530 227.800 ;
        RECT 59.530 227.000 63.530 227.200 ;
        RECT 63.130 226.400 63.530 227.000 ;
        RECT 59.530 226.200 63.530 226.400 ;
        RECT 63.130 225.600 63.530 226.200 ;
        RECT 59.530 225.400 63.530 225.600 ;
        RECT 63.130 224.800 63.530 225.400 ;
        RECT 59.530 224.600 63.530 224.800 ;
        RECT 63.130 224.000 63.530 224.600 ;
        RECT 59.530 223.800 63.530 224.000 ;
        RECT 63.130 223.200 63.530 223.800 ;
        RECT 59.530 223.000 63.530 223.200 ;
        RECT 63.130 222.400 63.530 223.000 ;
        RECT 59.530 222.200 63.530 222.400 ;
        RECT 65.930 237.600 69.930 237.800 ;
        RECT 65.930 237.000 66.330 237.600 ;
        RECT 65.930 236.800 69.930 237.000 ;
        RECT 65.930 236.200 66.330 236.800 ;
        RECT 65.930 236.000 69.930 236.200 ;
        RECT 65.930 235.400 66.330 236.000 ;
        RECT 65.930 235.200 69.930 235.400 ;
        RECT 65.930 234.600 66.330 235.200 ;
        RECT 65.930 234.400 69.930 234.600 ;
        RECT 65.930 233.800 66.330 234.400 ;
        RECT 65.930 233.600 69.930 233.800 ;
        RECT 65.930 233.000 66.330 233.600 ;
        RECT 65.930 232.800 69.930 233.000 ;
        RECT 65.930 232.200 66.330 232.800 ;
        RECT 65.930 232.000 69.930 232.200 ;
        RECT 65.930 231.400 66.330 232.000 ;
        RECT 65.930 231.200 69.930 231.400 ;
        RECT 65.930 230.600 66.330 231.200 ;
        RECT 65.930 230.400 69.930 230.600 ;
        RECT 65.930 230.200 66.330 230.400 ;
        RECT 70.680 230.200 70.880 237.800 ;
        RECT 71.480 230.200 71.680 237.800 ;
        RECT 72.280 230.200 72.480 237.800 ;
        RECT 73.080 230.200 73.280 237.800 ;
        RECT 73.880 230.200 74.080 237.800 ;
        RECT 65.930 229.800 74.080 230.200 ;
        RECT 65.930 229.600 66.330 229.800 ;
        RECT 65.930 229.400 69.930 229.600 ;
        RECT 65.930 228.800 66.330 229.400 ;
        RECT 65.930 228.600 69.930 228.800 ;
        RECT 65.930 228.000 66.330 228.600 ;
        RECT 65.930 227.800 69.930 228.000 ;
        RECT 65.930 227.200 66.330 227.800 ;
        RECT 65.930 227.000 69.930 227.200 ;
        RECT 65.930 226.400 66.330 227.000 ;
        RECT 65.930 226.200 69.930 226.400 ;
        RECT 65.930 225.600 66.330 226.200 ;
        RECT 65.930 225.400 69.930 225.600 ;
        RECT 65.930 224.800 66.330 225.400 ;
        RECT 65.930 224.600 69.930 224.800 ;
        RECT 65.930 224.000 66.330 224.600 ;
        RECT 65.930 223.800 69.930 224.000 ;
        RECT 65.930 223.200 66.330 223.800 ;
        RECT 65.930 223.000 69.930 223.200 ;
        RECT 65.930 222.400 66.330 223.000 ;
        RECT 65.930 222.200 69.930 222.400 ;
        RECT 70.680 222.200 70.880 229.800 ;
        RECT 71.480 222.200 71.680 229.800 ;
        RECT 72.280 222.200 72.480 229.800 ;
        RECT 73.080 222.200 73.280 229.800 ;
        RECT 73.880 222.200 74.080 229.800 ;
        RECT 75.380 230.200 75.580 237.800 ;
        RECT 76.180 230.200 76.380 237.800 ;
        RECT 76.980 230.200 77.180 237.800 ;
        RECT 77.780 230.200 77.980 237.800 ;
        RECT 78.580 230.200 78.780 237.800 ;
        RECT 79.530 237.600 83.530 237.800 ;
        RECT 83.130 237.000 83.530 237.600 ;
        RECT 79.530 236.800 83.530 237.000 ;
        RECT 83.130 236.200 83.530 236.800 ;
        RECT 79.530 236.000 83.530 236.200 ;
        RECT 83.130 235.400 83.530 236.000 ;
        RECT 79.530 235.200 83.530 235.400 ;
        RECT 83.130 234.600 83.530 235.200 ;
        RECT 79.530 234.400 83.530 234.600 ;
        RECT 83.130 233.800 83.530 234.400 ;
        RECT 79.530 233.600 83.530 233.800 ;
        RECT 83.130 233.000 83.530 233.600 ;
        RECT 79.530 232.800 83.530 233.000 ;
        RECT 83.130 232.200 83.530 232.800 ;
        RECT 79.530 232.000 83.530 232.200 ;
        RECT 83.130 231.400 83.530 232.000 ;
        RECT 79.530 231.200 83.530 231.400 ;
        RECT 83.130 230.600 83.530 231.200 ;
        RECT 79.530 230.400 83.530 230.600 ;
        RECT 83.130 230.200 83.530 230.400 ;
        RECT 75.380 229.800 83.530 230.200 ;
        RECT 75.380 222.200 75.580 229.800 ;
        RECT 76.180 222.200 76.380 229.800 ;
        RECT 76.980 222.200 77.180 229.800 ;
        RECT 77.780 222.200 77.980 229.800 ;
        RECT 78.580 222.200 78.780 229.800 ;
        RECT 83.130 229.600 83.530 229.800 ;
        RECT 79.530 229.400 83.530 229.600 ;
        RECT 83.130 228.800 83.530 229.400 ;
        RECT 79.530 228.600 83.530 228.800 ;
        RECT 83.130 228.000 83.530 228.600 ;
        RECT 79.530 227.800 83.530 228.000 ;
        RECT 83.130 227.200 83.530 227.800 ;
        RECT 79.530 227.000 83.530 227.200 ;
        RECT 83.130 226.400 83.530 227.000 ;
        RECT 79.530 226.200 83.530 226.400 ;
        RECT 83.130 225.600 83.530 226.200 ;
        RECT 79.530 225.400 83.530 225.600 ;
        RECT 83.130 224.800 83.530 225.400 ;
        RECT 79.530 224.600 83.530 224.800 ;
        RECT 83.130 224.000 83.530 224.600 ;
        RECT 79.530 223.800 83.530 224.000 ;
        RECT 83.130 223.200 83.530 223.800 ;
        RECT 79.530 223.000 83.530 223.200 ;
        RECT 83.130 222.400 83.530 223.000 ;
        RECT 79.530 222.200 83.530 222.400 ;
        RECT 85.930 237.600 89.930 237.800 ;
        RECT 85.930 237.000 86.330 237.600 ;
        RECT 85.930 236.800 89.930 237.000 ;
        RECT 85.930 236.200 86.330 236.800 ;
        RECT 85.930 236.000 89.930 236.200 ;
        RECT 85.930 235.400 86.330 236.000 ;
        RECT 85.930 235.200 89.930 235.400 ;
        RECT 85.930 234.600 86.330 235.200 ;
        RECT 85.930 234.400 89.930 234.600 ;
        RECT 85.930 233.800 86.330 234.400 ;
        RECT 85.930 233.600 89.930 233.800 ;
        RECT 85.930 233.000 86.330 233.600 ;
        RECT 85.930 232.800 89.930 233.000 ;
        RECT 85.930 232.200 86.330 232.800 ;
        RECT 85.930 232.000 89.930 232.200 ;
        RECT 85.930 231.400 86.330 232.000 ;
        RECT 85.930 231.200 89.930 231.400 ;
        RECT 85.930 230.600 86.330 231.200 ;
        RECT 85.930 230.400 89.930 230.600 ;
        RECT 85.930 230.200 86.330 230.400 ;
        RECT 90.680 230.200 90.880 237.800 ;
        RECT 91.480 230.200 91.680 237.800 ;
        RECT 92.280 230.200 92.480 237.800 ;
        RECT 93.080 230.200 93.280 237.800 ;
        RECT 93.880 230.200 94.080 237.800 ;
        RECT 85.930 229.800 94.080 230.200 ;
        RECT 85.930 229.600 86.330 229.800 ;
        RECT 85.930 229.400 89.930 229.600 ;
        RECT 85.930 228.800 86.330 229.400 ;
        RECT 85.930 228.600 89.930 228.800 ;
        RECT 85.930 228.000 86.330 228.600 ;
        RECT 85.930 227.800 89.930 228.000 ;
        RECT 85.930 227.200 86.330 227.800 ;
        RECT 85.930 227.000 89.930 227.200 ;
        RECT 85.930 226.400 86.330 227.000 ;
        RECT 85.930 226.200 89.930 226.400 ;
        RECT 85.930 225.600 86.330 226.200 ;
        RECT 85.930 225.400 89.930 225.600 ;
        RECT 85.930 224.800 86.330 225.400 ;
        RECT 85.930 224.600 89.930 224.800 ;
        RECT 85.930 224.000 86.330 224.600 ;
        RECT 85.930 223.800 89.930 224.000 ;
        RECT 85.930 223.200 86.330 223.800 ;
        RECT 85.930 223.000 89.930 223.200 ;
        RECT 85.930 222.400 86.330 223.000 ;
        RECT 85.930 222.200 89.930 222.400 ;
        RECT 90.680 222.200 90.880 229.800 ;
        RECT 91.480 222.200 91.680 229.800 ;
        RECT 92.280 222.200 92.480 229.800 ;
        RECT 93.080 222.200 93.280 229.800 ;
        RECT 93.880 222.200 94.080 229.800 ;
        RECT 95.380 230.200 95.580 237.800 ;
        RECT 96.180 230.200 96.380 237.800 ;
        RECT 96.980 230.200 97.180 237.800 ;
        RECT 97.780 230.200 97.980 237.800 ;
        RECT 98.580 230.200 98.780 237.800 ;
        RECT 99.530 237.600 103.530 237.800 ;
        RECT 103.130 237.000 103.530 237.600 ;
        RECT 99.530 236.800 103.530 237.000 ;
        RECT 103.130 236.200 103.530 236.800 ;
        RECT 99.530 236.000 103.530 236.200 ;
        RECT 103.130 235.400 103.530 236.000 ;
        RECT 99.530 235.200 103.530 235.400 ;
        RECT 103.130 234.600 103.530 235.200 ;
        RECT 99.530 234.400 103.530 234.600 ;
        RECT 103.130 233.800 103.530 234.400 ;
        RECT 99.530 233.600 103.530 233.800 ;
        RECT 103.130 233.000 103.530 233.600 ;
        RECT 99.530 232.800 103.530 233.000 ;
        RECT 103.130 232.200 103.530 232.800 ;
        RECT 99.530 232.000 103.530 232.200 ;
        RECT 103.130 231.400 103.530 232.000 ;
        RECT 99.530 231.200 103.530 231.400 ;
        RECT 103.130 230.600 103.530 231.200 ;
        RECT 99.530 230.400 103.530 230.600 ;
        RECT 103.130 230.200 103.530 230.400 ;
        RECT 95.380 229.800 103.530 230.200 ;
        RECT 95.380 222.200 95.580 229.800 ;
        RECT 96.180 222.200 96.380 229.800 ;
        RECT 96.980 222.200 97.180 229.800 ;
        RECT 97.780 222.200 97.980 229.800 ;
        RECT 98.580 222.200 98.780 229.800 ;
        RECT 103.130 229.600 103.530 229.800 ;
        RECT 99.530 229.400 103.530 229.600 ;
        RECT 103.130 228.800 103.530 229.400 ;
        RECT 110.050 229.120 110.410 229.500 ;
        RECT 110.680 229.120 111.040 229.500 ;
        RECT 111.280 229.120 111.640 229.500 ;
        RECT 99.530 228.600 103.530 228.800 ;
        RECT 103.130 228.000 103.530 228.600 ;
        RECT 110.050 228.530 110.410 228.910 ;
        RECT 110.680 228.530 111.040 228.910 ;
        RECT 111.280 228.530 111.640 228.910 ;
        RECT 99.530 227.800 103.530 228.000 ;
        RECT 103.130 227.200 103.530 227.800 ;
        RECT 99.530 227.000 103.530 227.200 ;
        RECT 103.130 226.400 103.530 227.000 ;
        RECT 99.530 226.200 103.530 226.400 ;
        RECT 103.130 225.600 103.530 226.200 ;
        RECT 99.530 225.400 103.530 225.600 ;
        RECT 103.130 224.800 103.530 225.400 ;
        RECT 99.530 224.600 103.530 224.800 ;
        RECT 103.130 224.000 103.530 224.600 ;
        RECT 99.530 223.800 103.530 224.000 ;
        RECT 103.130 223.200 103.530 223.800 ;
        RECT 99.530 223.000 103.530 223.200 ;
        RECT 103.130 222.400 103.530 223.000 ;
        RECT 99.530 222.200 103.530 222.400 ;
        RECT 9.340 196.355 12.515 197.050 ;
        RECT 9.340 196.350 10.045 196.355 ;
        RECT 11.755 195.425 12.515 196.355 ;
        RECT 10.175 193.440 10.345 195.425 ;
        RECT 11.755 194.885 12.570 195.425 ;
        RECT 13.965 194.885 14.155 195.425 ;
        RECT 11.755 193.440 11.925 194.885 ;
        RECT 12.395 194.255 12.570 194.885 ;
        RECT 12.400 193.445 12.570 194.255 ;
        RECT 13.980 194.255 14.155 194.885 ;
        RECT 13.980 193.445 14.150 194.255 ;
        RECT 5.930 157.600 9.930 157.800 ;
        RECT 5.930 157.000 6.330 157.600 ;
        RECT 5.930 156.800 9.930 157.000 ;
        RECT 5.930 156.200 6.330 156.800 ;
        RECT 5.930 156.000 9.930 156.200 ;
        RECT 5.930 155.400 6.330 156.000 ;
        RECT 5.930 155.200 9.930 155.400 ;
        RECT 5.930 154.600 6.330 155.200 ;
        RECT 5.930 154.400 9.930 154.600 ;
        RECT 5.930 153.800 6.330 154.400 ;
        RECT 5.930 153.600 9.930 153.800 ;
        RECT 5.930 153.000 6.330 153.600 ;
        RECT 5.930 152.800 9.930 153.000 ;
        RECT 5.930 152.200 6.330 152.800 ;
        RECT 5.930 152.000 9.930 152.200 ;
        RECT 5.930 151.400 6.330 152.000 ;
        RECT 5.930 151.200 9.930 151.400 ;
        RECT 5.930 150.600 6.330 151.200 ;
        RECT 5.930 150.400 9.930 150.600 ;
        RECT 5.930 150.200 6.330 150.400 ;
        RECT 10.680 150.200 10.880 157.800 ;
        RECT 11.480 150.200 11.680 157.800 ;
        RECT 12.280 150.200 12.480 157.800 ;
        RECT 13.080 150.200 13.280 157.800 ;
        RECT 13.880 150.200 14.080 157.800 ;
        RECT 5.930 149.800 14.080 150.200 ;
        RECT 5.930 149.600 6.330 149.800 ;
        RECT 5.930 149.400 9.930 149.600 ;
        RECT 5.930 148.800 6.330 149.400 ;
        RECT 5.930 148.600 9.930 148.800 ;
        RECT 5.930 148.000 6.330 148.600 ;
        RECT 5.930 147.800 9.930 148.000 ;
        RECT 5.930 147.200 6.330 147.800 ;
        RECT 5.930 147.000 9.930 147.200 ;
        RECT 5.930 146.400 6.330 147.000 ;
        RECT 5.930 146.200 9.930 146.400 ;
        RECT 5.930 145.600 6.330 146.200 ;
        RECT 5.930 145.400 9.930 145.600 ;
        RECT 5.930 144.800 6.330 145.400 ;
        RECT 5.930 144.600 9.930 144.800 ;
        RECT 5.930 144.000 6.330 144.600 ;
        RECT 5.930 143.800 9.930 144.000 ;
        RECT 5.930 143.200 6.330 143.800 ;
        RECT 5.930 143.000 9.930 143.200 ;
        RECT 5.930 142.400 6.330 143.000 ;
        RECT 5.930 142.200 9.930 142.400 ;
        RECT 10.680 142.200 10.880 149.800 ;
        RECT 11.480 142.200 11.680 149.800 ;
        RECT 12.280 142.200 12.480 149.800 ;
        RECT 13.080 142.200 13.280 149.800 ;
        RECT 13.880 142.200 14.080 149.800 ;
        RECT 15.380 150.200 15.580 157.800 ;
        RECT 16.180 150.200 16.380 157.800 ;
        RECT 16.980 150.200 17.180 157.800 ;
        RECT 17.780 150.200 17.980 157.800 ;
        RECT 18.580 150.200 18.780 157.800 ;
        RECT 19.530 157.600 23.530 157.800 ;
        RECT 23.130 157.000 23.530 157.600 ;
        RECT 19.530 156.800 23.530 157.000 ;
        RECT 23.130 156.200 23.530 156.800 ;
        RECT 19.530 156.000 23.530 156.200 ;
        RECT 23.130 155.400 23.530 156.000 ;
        RECT 19.530 155.200 23.530 155.400 ;
        RECT 23.130 154.600 23.530 155.200 ;
        RECT 19.530 154.400 23.530 154.600 ;
        RECT 23.130 153.800 23.530 154.400 ;
        RECT 19.530 153.600 23.530 153.800 ;
        RECT 23.130 153.000 23.530 153.600 ;
        RECT 19.530 152.800 23.530 153.000 ;
        RECT 23.130 152.200 23.530 152.800 ;
        RECT 19.530 152.000 23.530 152.200 ;
        RECT 23.130 151.400 23.530 152.000 ;
        RECT 19.530 151.200 23.530 151.400 ;
        RECT 23.130 150.600 23.530 151.200 ;
        RECT 19.530 150.400 23.530 150.600 ;
        RECT 23.130 150.200 23.530 150.400 ;
        RECT 15.380 149.800 23.530 150.200 ;
        RECT 15.380 142.200 15.580 149.800 ;
        RECT 16.180 142.200 16.380 149.800 ;
        RECT 16.980 142.200 17.180 149.800 ;
        RECT 17.780 142.200 17.980 149.800 ;
        RECT 18.580 142.200 18.780 149.800 ;
        RECT 23.130 149.600 23.530 149.800 ;
        RECT 19.530 149.400 23.530 149.600 ;
        RECT 23.130 148.800 23.530 149.400 ;
        RECT 19.530 148.600 23.530 148.800 ;
        RECT 23.130 148.000 23.530 148.600 ;
        RECT 19.530 147.800 23.530 148.000 ;
        RECT 23.130 147.200 23.530 147.800 ;
        RECT 19.530 147.000 23.530 147.200 ;
        RECT 23.130 146.400 23.530 147.000 ;
        RECT 19.530 146.200 23.530 146.400 ;
        RECT 23.130 145.600 23.530 146.200 ;
        RECT 19.530 145.400 23.530 145.600 ;
        RECT 23.130 144.800 23.530 145.400 ;
        RECT 19.530 144.600 23.530 144.800 ;
        RECT 23.130 144.000 23.530 144.600 ;
        RECT 19.530 143.800 23.530 144.000 ;
        RECT 23.130 143.200 23.530 143.800 ;
        RECT 19.530 143.000 23.530 143.200 ;
        RECT 23.130 142.400 23.530 143.000 ;
        RECT 19.530 142.200 23.530 142.400 ;
        RECT 25.930 157.600 29.930 157.800 ;
        RECT 25.930 157.000 26.330 157.600 ;
        RECT 25.930 156.800 29.930 157.000 ;
        RECT 25.930 156.200 26.330 156.800 ;
        RECT 25.930 156.000 29.930 156.200 ;
        RECT 25.930 155.400 26.330 156.000 ;
        RECT 25.930 155.200 29.930 155.400 ;
        RECT 25.930 154.600 26.330 155.200 ;
        RECT 25.930 154.400 29.930 154.600 ;
        RECT 25.930 153.800 26.330 154.400 ;
        RECT 25.930 153.600 29.930 153.800 ;
        RECT 25.930 153.000 26.330 153.600 ;
        RECT 25.930 152.800 29.930 153.000 ;
        RECT 25.930 152.200 26.330 152.800 ;
        RECT 25.930 152.000 29.930 152.200 ;
        RECT 25.930 151.400 26.330 152.000 ;
        RECT 25.930 151.200 29.930 151.400 ;
        RECT 25.930 150.600 26.330 151.200 ;
        RECT 25.930 150.400 29.930 150.600 ;
        RECT 25.930 150.200 26.330 150.400 ;
        RECT 30.680 150.200 30.880 157.800 ;
        RECT 31.480 150.200 31.680 157.800 ;
        RECT 32.280 150.200 32.480 157.800 ;
        RECT 33.080 150.200 33.280 157.800 ;
        RECT 33.880 150.200 34.080 157.800 ;
        RECT 25.930 149.800 34.080 150.200 ;
        RECT 25.930 149.600 26.330 149.800 ;
        RECT 25.930 149.400 29.930 149.600 ;
        RECT 25.930 148.800 26.330 149.400 ;
        RECT 25.930 148.600 29.930 148.800 ;
        RECT 25.930 148.000 26.330 148.600 ;
        RECT 25.930 147.800 29.930 148.000 ;
        RECT 25.930 147.200 26.330 147.800 ;
        RECT 25.930 147.000 29.930 147.200 ;
        RECT 25.930 146.400 26.330 147.000 ;
        RECT 25.930 146.200 29.930 146.400 ;
        RECT 25.930 145.600 26.330 146.200 ;
        RECT 25.930 145.400 29.930 145.600 ;
        RECT 25.930 144.800 26.330 145.400 ;
        RECT 25.930 144.600 29.930 144.800 ;
        RECT 25.930 144.000 26.330 144.600 ;
        RECT 25.930 143.800 29.930 144.000 ;
        RECT 25.930 143.200 26.330 143.800 ;
        RECT 25.930 143.000 29.930 143.200 ;
        RECT 25.930 142.400 26.330 143.000 ;
        RECT 25.930 142.200 29.930 142.400 ;
        RECT 30.680 142.200 30.880 149.800 ;
        RECT 31.480 142.200 31.680 149.800 ;
        RECT 32.280 142.200 32.480 149.800 ;
        RECT 33.080 142.200 33.280 149.800 ;
        RECT 33.880 142.200 34.080 149.800 ;
        RECT 35.380 150.200 35.580 157.800 ;
        RECT 36.180 150.200 36.380 157.800 ;
        RECT 36.980 150.200 37.180 157.800 ;
        RECT 37.780 150.200 37.980 157.800 ;
        RECT 38.580 150.200 38.780 157.800 ;
        RECT 39.530 157.600 43.530 157.800 ;
        RECT 43.130 157.000 43.530 157.600 ;
        RECT 39.530 156.800 43.530 157.000 ;
        RECT 43.130 156.200 43.530 156.800 ;
        RECT 39.530 156.000 43.530 156.200 ;
        RECT 43.130 155.400 43.530 156.000 ;
        RECT 39.530 155.200 43.530 155.400 ;
        RECT 43.130 154.600 43.530 155.200 ;
        RECT 39.530 154.400 43.530 154.600 ;
        RECT 43.130 153.800 43.530 154.400 ;
        RECT 39.530 153.600 43.530 153.800 ;
        RECT 43.130 153.000 43.530 153.600 ;
        RECT 39.530 152.800 43.530 153.000 ;
        RECT 43.130 152.200 43.530 152.800 ;
        RECT 39.530 152.000 43.530 152.200 ;
        RECT 43.130 151.400 43.530 152.000 ;
        RECT 39.530 151.200 43.530 151.400 ;
        RECT 43.130 150.600 43.530 151.200 ;
        RECT 39.530 150.400 43.530 150.600 ;
        RECT 43.130 150.200 43.530 150.400 ;
        RECT 35.380 149.800 43.530 150.200 ;
        RECT 35.380 142.200 35.580 149.800 ;
        RECT 36.180 142.200 36.380 149.800 ;
        RECT 36.980 142.200 37.180 149.800 ;
        RECT 37.780 142.200 37.980 149.800 ;
        RECT 38.580 142.200 38.780 149.800 ;
        RECT 43.130 149.600 43.530 149.800 ;
        RECT 39.530 149.400 43.530 149.600 ;
        RECT 43.130 148.800 43.530 149.400 ;
        RECT 39.530 148.600 43.530 148.800 ;
        RECT 43.130 148.000 43.530 148.600 ;
        RECT 39.530 147.800 43.530 148.000 ;
        RECT 43.130 147.200 43.530 147.800 ;
        RECT 39.530 147.000 43.530 147.200 ;
        RECT 43.130 146.400 43.530 147.000 ;
        RECT 39.530 146.200 43.530 146.400 ;
        RECT 43.130 145.600 43.530 146.200 ;
        RECT 39.530 145.400 43.530 145.600 ;
        RECT 43.130 144.800 43.530 145.400 ;
        RECT 39.530 144.600 43.530 144.800 ;
        RECT 43.130 144.000 43.530 144.600 ;
        RECT 39.530 143.800 43.530 144.000 ;
        RECT 43.130 143.200 43.530 143.800 ;
        RECT 39.530 143.000 43.530 143.200 ;
        RECT 43.130 142.400 43.530 143.000 ;
        RECT 39.530 142.200 43.530 142.400 ;
        RECT 45.930 157.600 49.930 157.800 ;
        RECT 45.930 157.000 46.330 157.600 ;
        RECT 45.930 156.800 49.930 157.000 ;
        RECT 45.930 156.200 46.330 156.800 ;
        RECT 45.930 156.000 49.930 156.200 ;
        RECT 45.930 155.400 46.330 156.000 ;
        RECT 45.930 155.200 49.930 155.400 ;
        RECT 45.930 154.600 46.330 155.200 ;
        RECT 45.930 154.400 49.930 154.600 ;
        RECT 45.930 153.800 46.330 154.400 ;
        RECT 45.930 153.600 49.930 153.800 ;
        RECT 45.930 153.000 46.330 153.600 ;
        RECT 45.930 152.800 49.930 153.000 ;
        RECT 45.930 152.200 46.330 152.800 ;
        RECT 45.930 152.000 49.930 152.200 ;
        RECT 45.930 151.400 46.330 152.000 ;
        RECT 45.930 151.200 49.930 151.400 ;
        RECT 45.930 150.600 46.330 151.200 ;
        RECT 45.930 150.400 49.930 150.600 ;
        RECT 45.930 150.200 46.330 150.400 ;
        RECT 50.680 150.200 50.880 157.800 ;
        RECT 51.480 150.200 51.680 157.800 ;
        RECT 52.280 150.200 52.480 157.800 ;
        RECT 53.080 150.200 53.280 157.800 ;
        RECT 53.880 150.200 54.080 157.800 ;
        RECT 45.930 149.800 54.080 150.200 ;
        RECT 45.930 149.600 46.330 149.800 ;
        RECT 45.930 149.400 49.930 149.600 ;
        RECT 45.930 148.800 46.330 149.400 ;
        RECT 45.930 148.600 49.930 148.800 ;
        RECT 45.930 148.000 46.330 148.600 ;
        RECT 45.930 147.800 49.930 148.000 ;
        RECT 45.930 147.200 46.330 147.800 ;
        RECT 45.930 147.000 49.930 147.200 ;
        RECT 45.930 146.400 46.330 147.000 ;
        RECT 45.930 146.200 49.930 146.400 ;
        RECT 45.930 145.600 46.330 146.200 ;
        RECT 45.930 145.400 49.930 145.600 ;
        RECT 45.930 144.800 46.330 145.400 ;
        RECT 45.930 144.600 49.930 144.800 ;
        RECT 45.930 144.000 46.330 144.600 ;
        RECT 45.930 143.800 49.930 144.000 ;
        RECT 45.930 143.200 46.330 143.800 ;
        RECT 45.930 143.000 49.930 143.200 ;
        RECT 45.930 142.400 46.330 143.000 ;
        RECT 45.930 142.200 49.930 142.400 ;
        RECT 50.680 142.200 50.880 149.800 ;
        RECT 51.480 142.200 51.680 149.800 ;
        RECT 52.280 142.200 52.480 149.800 ;
        RECT 53.080 142.200 53.280 149.800 ;
        RECT 53.880 142.200 54.080 149.800 ;
        RECT 55.380 150.200 55.580 157.800 ;
        RECT 56.180 150.200 56.380 157.800 ;
        RECT 56.980 150.200 57.180 157.800 ;
        RECT 57.780 150.200 57.980 157.800 ;
        RECT 58.580 150.200 58.780 157.800 ;
        RECT 59.530 157.600 63.530 157.800 ;
        RECT 63.130 157.000 63.530 157.600 ;
        RECT 59.530 156.800 63.530 157.000 ;
        RECT 63.130 156.200 63.530 156.800 ;
        RECT 59.530 156.000 63.530 156.200 ;
        RECT 63.130 155.400 63.530 156.000 ;
        RECT 59.530 155.200 63.530 155.400 ;
        RECT 63.130 154.600 63.530 155.200 ;
        RECT 59.530 154.400 63.530 154.600 ;
        RECT 63.130 153.800 63.530 154.400 ;
        RECT 59.530 153.600 63.530 153.800 ;
        RECT 63.130 153.000 63.530 153.600 ;
        RECT 59.530 152.800 63.530 153.000 ;
        RECT 63.130 152.200 63.530 152.800 ;
        RECT 59.530 152.000 63.530 152.200 ;
        RECT 63.130 151.400 63.530 152.000 ;
        RECT 59.530 151.200 63.530 151.400 ;
        RECT 63.130 150.600 63.530 151.200 ;
        RECT 59.530 150.400 63.530 150.600 ;
        RECT 63.130 150.200 63.530 150.400 ;
        RECT 55.380 149.800 63.530 150.200 ;
        RECT 55.380 142.200 55.580 149.800 ;
        RECT 56.180 142.200 56.380 149.800 ;
        RECT 56.980 142.200 57.180 149.800 ;
        RECT 57.780 142.200 57.980 149.800 ;
        RECT 58.580 142.200 58.780 149.800 ;
        RECT 63.130 149.600 63.530 149.800 ;
        RECT 59.530 149.400 63.530 149.600 ;
        RECT 63.130 148.800 63.530 149.400 ;
        RECT 59.530 148.600 63.530 148.800 ;
        RECT 63.130 148.000 63.530 148.600 ;
        RECT 59.530 147.800 63.530 148.000 ;
        RECT 63.130 147.200 63.530 147.800 ;
        RECT 59.530 147.000 63.530 147.200 ;
        RECT 63.130 146.400 63.530 147.000 ;
        RECT 59.530 146.200 63.530 146.400 ;
        RECT 63.130 145.600 63.530 146.200 ;
        RECT 59.530 145.400 63.530 145.600 ;
        RECT 63.130 144.800 63.530 145.400 ;
        RECT 59.530 144.600 63.530 144.800 ;
        RECT 63.130 144.000 63.530 144.600 ;
        RECT 59.530 143.800 63.530 144.000 ;
        RECT 63.130 143.200 63.530 143.800 ;
        RECT 59.530 143.000 63.530 143.200 ;
        RECT 63.130 142.400 63.530 143.000 ;
        RECT 59.530 142.200 63.530 142.400 ;
        RECT 65.930 157.600 69.930 157.800 ;
        RECT 65.930 157.000 66.330 157.600 ;
        RECT 65.930 156.800 69.930 157.000 ;
        RECT 65.930 156.200 66.330 156.800 ;
        RECT 65.930 156.000 69.930 156.200 ;
        RECT 65.930 155.400 66.330 156.000 ;
        RECT 65.930 155.200 69.930 155.400 ;
        RECT 65.930 154.600 66.330 155.200 ;
        RECT 65.930 154.400 69.930 154.600 ;
        RECT 65.930 153.800 66.330 154.400 ;
        RECT 65.930 153.600 69.930 153.800 ;
        RECT 65.930 153.000 66.330 153.600 ;
        RECT 65.930 152.800 69.930 153.000 ;
        RECT 65.930 152.200 66.330 152.800 ;
        RECT 65.930 152.000 69.930 152.200 ;
        RECT 65.930 151.400 66.330 152.000 ;
        RECT 65.930 151.200 69.930 151.400 ;
        RECT 65.930 150.600 66.330 151.200 ;
        RECT 65.930 150.400 69.930 150.600 ;
        RECT 65.930 150.200 66.330 150.400 ;
        RECT 70.680 150.200 70.880 157.800 ;
        RECT 71.480 150.200 71.680 157.800 ;
        RECT 72.280 150.200 72.480 157.800 ;
        RECT 73.080 150.200 73.280 157.800 ;
        RECT 73.880 150.200 74.080 157.800 ;
        RECT 65.930 149.800 74.080 150.200 ;
        RECT 65.930 149.600 66.330 149.800 ;
        RECT 65.930 149.400 69.930 149.600 ;
        RECT 65.930 148.800 66.330 149.400 ;
        RECT 65.930 148.600 69.930 148.800 ;
        RECT 65.930 148.000 66.330 148.600 ;
        RECT 65.930 147.800 69.930 148.000 ;
        RECT 65.930 147.200 66.330 147.800 ;
        RECT 65.930 147.000 69.930 147.200 ;
        RECT 65.930 146.400 66.330 147.000 ;
        RECT 65.930 146.200 69.930 146.400 ;
        RECT 65.930 145.600 66.330 146.200 ;
        RECT 65.930 145.400 69.930 145.600 ;
        RECT 65.930 144.800 66.330 145.400 ;
        RECT 65.930 144.600 69.930 144.800 ;
        RECT 65.930 144.000 66.330 144.600 ;
        RECT 65.930 143.800 69.930 144.000 ;
        RECT 65.930 143.200 66.330 143.800 ;
        RECT 65.930 143.000 69.930 143.200 ;
        RECT 65.930 142.400 66.330 143.000 ;
        RECT 65.930 142.200 69.930 142.400 ;
        RECT 70.680 142.200 70.880 149.800 ;
        RECT 71.480 142.200 71.680 149.800 ;
        RECT 72.280 142.200 72.480 149.800 ;
        RECT 73.080 142.200 73.280 149.800 ;
        RECT 73.880 142.200 74.080 149.800 ;
        RECT 75.380 150.200 75.580 157.800 ;
        RECT 76.180 150.200 76.380 157.800 ;
        RECT 76.980 150.200 77.180 157.800 ;
        RECT 77.780 150.200 77.980 157.800 ;
        RECT 78.580 150.200 78.780 157.800 ;
        RECT 79.530 157.600 83.530 157.800 ;
        RECT 83.130 157.000 83.530 157.600 ;
        RECT 79.530 156.800 83.530 157.000 ;
        RECT 83.130 156.200 83.530 156.800 ;
        RECT 79.530 156.000 83.530 156.200 ;
        RECT 83.130 155.400 83.530 156.000 ;
        RECT 79.530 155.200 83.530 155.400 ;
        RECT 83.130 154.600 83.530 155.200 ;
        RECT 79.530 154.400 83.530 154.600 ;
        RECT 83.130 153.800 83.530 154.400 ;
        RECT 79.530 153.600 83.530 153.800 ;
        RECT 83.130 153.000 83.530 153.600 ;
        RECT 79.530 152.800 83.530 153.000 ;
        RECT 83.130 152.200 83.530 152.800 ;
        RECT 79.530 152.000 83.530 152.200 ;
        RECT 83.130 151.400 83.530 152.000 ;
        RECT 79.530 151.200 83.530 151.400 ;
        RECT 83.130 150.600 83.530 151.200 ;
        RECT 79.530 150.400 83.530 150.600 ;
        RECT 83.130 150.200 83.530 150.400 ;
        RECT 75.380 149.800 83.530 150.200 ;
        RECT 75.380 142.200 75.580 149.800 ;
        RECT 76.180 142.200 76.380 149.800 ;
        RECT 76.980 142.200 77.180 149.800 ;
        RECT 77.780 142.200 77.980 149.800 ;
        RECT 78.580 142.200 78.780 149.800 ;
        RECT 83.130 149.600 83.530 149.800 ;
        RECT 79.530 149.400 83.530 149.600 ;
        RECT 83.130 148.800 83.530 149.400 ;
        RECT 79.530 148.600 83.530 148.800 ;
        RECT 83.130 148.000 83.530 148.600 ;
        RECT 79.530 147.800 83.530 148.000 ;
        RECT 83.130 147.200 83.530 147.800 ;
        RECT 79.530 147.000 83.530 147.200 ;
        RECT 83.130 146.400 83.530 147.000 ;
        RECT 79.530 146.200 83.530 146.400 ;
        RECT 83.130 145.600 83.530 146.200 ;
        RECT 79.530 145.400 83.530 145.600 ;
        RECT 83.130 144.800 83.530 145.400 ;
        RECT 79.530 144.600 83.530 144.800 ;
        RECT 83.130 144.000 83.530 144.600 ;
        RECT 79.530 143.800 83.530 144.000 ;
        RECT 83.130 143.200 83.530 143.800 ;
        RECT 79.530 143.000 83.530 143.200 ;
        RECT 83.130 142.400 83.530 143.000 ;
        RECT 79.530 142.200 83.530 142.400 ;
        RECT 85.930 157.600 89.930 157.800 ;
        RECT 85.930 157.000 86.330 157.600 ;
        RECT 85.930 156.800 89.930 157.000 ;
        RECT 85.930 156.200 86.330 156.800 ;
        RECT 85.930 156.000 89.930 156.200 ;
        RECT 85.930 155.400 86.330 156.000 ;
        RECT 85.930 155.200 89.930 155.400 ;
        RECT 85.930 154.600 86.330 155.200 ;
        RECT 85.930 154.400 89.930 154.600 ;
        RECT 85.930 153.800 86.330 154.400 ;
        RECT 85.930 153.600 89.930 153.800 ;
        RECT 85.930 153.000 86.330 153.600 ;
        RECT 85.930 152.800 89.930 153.000 ;
        RECT 85.930 152.200 86.330 152.800 ;
        RECT 85.930 152.000 89.930 152.200 ;
        RECT 85.930 151.400 86.330 152.000 ;
        RECT 85.930 151.200 89.930 151.400 ;
        RECT 85.930 150.600 86.330 151.200 ;
        RECT 85.930 150.400 89.930 150.600 ;
        RECT 85.930 150.200 86.330 150.400 ;
        RECT 90.680 150.200 90.880 157.800 ;
        RECT 91.480 150.200 91.680 157.800 ;
        RECT 92.280 150.200 92.480 157.800 ;
        RECT 93.080 150.200 93.280 157.800 ;
        RECT 93.880 150.200 94.080 157.800 ;
        RECT 85.930 149.800 94.080 150.200 ;
        RECT 85.930 149.600 86.330 149.800 ;
        RECT 85.930 149.400 89.930 149.600 ;
        RECT 85.930 148.800 86.330 149.400 ;
        RECT 85.930 148.600 89.930 148.800 ;
        RECT 85.930 148.000 86.330 148.600 ;
        RECT 85.930 147.800 89.930 148.000 ;
        RECT 85.930 147.200 86.330 147.800 ;
        RECT 85.930 147.000 89.930 147.200 ;
        RECT 85.930 146.400 86.330 147.000 ;
        RECT 85.930 146.200 89.930 146.400 ;
        RECT 85.930 145.600 86.330 146.200 ;
        RECT 85.930 145.400 89.930 145.600 ;
        RECT 85.930 144.800 86.330 145.400 ;
        RECT 85.930 144.600 89.930 144.800 ;
        RECT 85.930 144.000 86.330 144.600 ;
        RECT 85.930 143.800 89.930 144.000 ;
        RECT 85.930 143.200 86.330 143.800 ;
        RECT 85.930 143.000 89.930 143.200 ;
        RECT 85.930 142.400 86.330 143.000 ;
        RECT 85.930 142.200 89.930 142.400 ;
        RECT 90.680 142.200 90.880 149.800 ;
        RECT 91.480 142.200 91.680 149.800 ;
        RECT 92.280 142.200 92.480 149.800 ;
        RECT 93.080 142.200 93.280 149.800 ;
        RECT 93.880 142.200 94.080 149.800 ;
        RECT 95.380 150.200 95.580 157.800 ;
        RECT 96.180 150.200 96.380 157.800 ;
        RECT 96.980 150.200 97.180 157.800 ;
        RECT 97.780 150.200 97.980 157.800 ;
        RECT 98.580 150.200 98.780 157.800 ;
        RECT 99.530 157.600 103.530 157.800 ;
        RECT 103.130 157.000 103.530 157.600 ;
        RECT 99.530 156.800 103.530 157.000 ;
        RECT 103.130 156.200 103.530 156.800 ;
        RECT 99.530 156.000 103.530 156.200 ;
        RECT 103.130 155.400 103.530 156.000 ;
        RECT 99.530 155.200 103.530 155.400 ;
        RECT 103.130 154.600 103.530 155.200 ;
        RECT 99.530 154.400 103.530 154.600 ;
        RECT 103.130 153.800 103.530 154.400 ;
        RECT 99.530 153.600 103.530 153.800 ;
        RECT 103.130 153.000 103.530 153.600 ;
        RECT 99.530 152.800 103.530 153.000 ;
        RECT 103.130 152.200 103.530 152.800 ;
        RECT 99.530 152.000 103.530 152.200 ;
        RECT 103.130 151.400 103.530 152.000 ;
        RECT 99.530 151.200 103.530 151.400 ;
        RECT 103.130 150.600 103.530 151.200 ;
        RECT 99.530 150.400 103.530 150.600 ;
        RECT 103.130 150.200 103.530 150.400 ;
        RECT 110.050 150.270 110.410 150.650 ;
        RECT 110.680 150.270 111.040 150.650 ;
        RECT 111.280 150.270 111.640 150.650 ;
        RECT 95.380 149.800 103.530 150.200 ;
        RECT 95.380 142.200 95.580 149.800 ;
        RECT 96.180 142.200 96.380 149.800 ;
        RECT 96.980 142.200 97.180 149.800 ;
        RECT 97.780 142.200 97.980 149.800 ;
        RECT 98.580 142.200 98.780 149.800 ;
        RECT 103.130 149.600 103.530 149.800 ;
        RECT 110.050 149.680 110.410 150.060 ;
        RECT 110.680 149.680 111.040 150.060 ;
        RECT 111.280 149.680 111.640 150.060 ;
        RECT 99.530 149.400 103.530 149.600 ;
        RECT 103.130 148.800 103.530 149.400 ;
        RECT 99.530 148.600 103.530 148.800 ;
        RECT 103.130 148.000 103.530 148.600 ;
        RECT 99.530 147.800 103.530 148.000 ;
        RECT 103.130 147.200 103.530 147.800 ;
        RECT 99.530 147.000 103.530 147.200 ;
        RECT 103.130 146.400 103.530 147.000 ;
        RECT 99.530 146.200 103.530 146.400 ;
        RECT 103.130 145.600 103.530 146.200 ;
        RECT 99.530 145.400 103.530 145.600 ;
        RECT 103.130 144.800 103.530 145.400 ;
        RECT 99.530 144.600 103.530 144.800 ;
        RECT 103.130 144.000 103.530 144.600 ;
        RECT 99.530 143.800 103.530 144.000 ;
        RECT 103.130 143.200 103.530 143.800 ;
        RECT 99.530 143.000 103.530 143.200 ;
        RECT 103.130 142.400 103.530 143.000 ;
        RECT 99.530 142.200 103.530 142.400 ;
        RECT 5.930 137.600 9.930 137.800 ;
        RECT 5.930 137.000 6.330 137.600 ;
        RECT 5.930 136.800 9.930 137.000 ;
        RECT 5.930 136.200 6.330 136.800 ;
        RECT 5.930 136.000 9.930 136.200 ;
        RECT 5.930 135.400 6.330 136.000 ;
        RECT 5.930 135.200 9.930 135.400 ;
        RECT 5.930 134.600 6.330 135.200 ;
        RECT 5.930 134.400 9.930 134.600 ;
        RECT 5.930 133.800 6.330 134.400 ;
        RECT 5.930 133.600 9.930 133.800 ;
        RECT 5.930 133.000 6.330 133.600 ;
        RECT 5.930 132.800 9.930 133.000 ;
        RECT 5.930 132.200 6.330 132.800 ;
        RECT 5.930 132.000 9.930 132.200 ;
        RECT 5.930 131.400 6.330 132.000 ;
        RECT 5.930 131.200 9.930 131.400 ;
        RECT 5.930 130.600 6.330 131.200 ;
        RECT 5.930 130.400 9.930 130.600 ;
        RECT 5.930 130.200 6.330 130.400 ;
        RECT 10.680 130.200 10.880 137.800 ;
        RECT 11.480 130.200 11.680 137.800 ;
        RECT 12.280 130.200 12.480 137.800 ;
        RECT 13.080 130.200 13.280 137.800 ;
        RECT 13.880 130.200 14.080 137.800 ;
        RECT 5.930 129.800 14.080 130.200 ;
        RECT 5.930 129.600 6.330 129.800 ;
        RECT 5.930 129.400 9.930 129.600 ;
        RECT 5.930 128.800 6.330 129.400 ;
        RECT 5.930 128.600 9.930 128.800 ;
        RECT 5.930 128.000 6.330 128.600 ;
        RECT 5.930 127.800 9.930 128.000 ;
        RECT 5.930 127.200 6.330 127.800 ;
        RECT 5.930 127.000 9.930 127.200 ;
        RECT 5.930 126.400 6.330 127.000 ;
        RECT 5.930 126.200 9.930 126.400 ;
        RECT 5.930 125.600 6.330 126.200 ;
        RECT 5.930 125.400 9.930 125.600 ;
        RECT 5.930 124.800 6.330 125.400 ;
        RECT 5.930 124.600 9.930 124.800 ;
        RECT 5.930 124.000 6.330 124.600 ;
        RECT 5.930 123.800 9.930 124.000 ;
        RECT 5.930 123.200 6.330 123.800 ;
        RECT 5.930 123.000 9.930 123.200 ;
        RECT 5.930 122.400 6.330 123.000 ;
        RECT 5.930 122.200 9.930 122.400 ;
        RECT 10.680 122.200 10.880 129.800 ;
        RECT 11.480 122.200 11.680 129.800 ;
        RECT 12.280 122.200 12.480 129.800 ;
        RECT 13.080 122.200 13.280 129.800 ;
        RECT 13.880 122.200 14.080 129.800 ;
        RECT 15.380 130.200 15.580 137.800 ;
        RECT 16.180 130.200 16.380 137.800 ;
        RECT 16.980 130.200 17.180 137.800 ;
        RECT 17.780 130.200 17.980 137.800 ;
        RECT 18.580 130.200 18.780 137.800 ;
        RECT 19.530 137.600 23.530 137.800 ;
        RECT 23.130 137.000 23.530 137.600 ;
        RECT 19.530 136.800 23.530 137.000 ;
        RECT 23.130 136.200 23.530 136.800 ;
        RECT 19.530 136.000 23.530 136.200 ;
        RECT 23.130 135.400 23.530 136.000 ;
        RECT 19.530 135.200 23.530 135.400 ;
        RECT 23.130 134.600 23.530 135.200 ;
        RECT 19.530 134.400 23.530 134.600 ;
        RECT 23.130 133.800 23.530 134.400 ;
        RECT 19.530 133.600 23.530 133.800 ;
        RECT 23.130 133.000 23.530 133.600 ;
        RECT 19.530 132.800 23.530 133.000 ;
        RECT 23.130 132.200 23.530 132.800 ;
        RECT 19.530 132.000 23.530 132.200 ;
        RECT 23.130 131.400 23.530 132.000 ;
        RECT 19.530 131.200 23.530 131.400 ;
        RECT 23.130 130.600 23.530 131.200 ;
        RECT 19.530 130.400 23.530 130.600 ;
        RECT 23.130 130.200 23.530 130.400 ;
        RECT 15.380 129.800 23.530 130.200 ;
        RECT 15.380 122.200 15.580 129.800 ;
        RECT 16.180 122.200 16.380 129.800 ;
        RECT 16.980 122.200 17.180 129.800 ;
        RECT 17.780 122.200 17.980 129.800 ;
        RECT 18.580 122.200 18.780 129.800 ;
        RECT 23.130 129.600 23.530 129.800 ;
        RECT 19.530 129.400 23.530 129.600 ;
        RECT 23.130 128.800 23.530 129.400 ;
        RECT 19.530 128.600 23.530 128.800 ;
        RECT 23.130 128.000 23.530 128.600 ;
        RECT 19.530 127.800 23.530 128.000 ;
        RECT 23.130 127.200 23.530 127.800 ;
        RECT 19.530 127.000 23.530 127.200 ;
        RECT 23.130 126.400 23.530 127.000 ;
        RECT 19.530 126.200 23.530 126.400 ;
        RECT 23.130 125.600 23.530 126.200 ;
        RECT 19.530 125.400 23.530 125.600 ;
        RECT 23.130 124.800 23.530 125.400 ;
        RECT 19.530 124.600 23.530 124.800 ;
        RECT 23.130 124.000 23.530 124.600 ;
        RECT 19.530 123.800 23.530 124.000 ;
        RECT 23.130 123.200 23.530 123.800 ;
        RECT 19.530 123.000 23.530 123.200 ;
        RECT 23.130 122.400 23.530 123.000 ;
        RECT 19.530 122.200 23.530 122.400 ;
        RECT 25.930 137.600 29.930 137.800 ;
        RECT 25.930 137.000 26.330 137.600 ;
        RECT 25.930 136.800 29.930 137.000 ;
        RECT 25.930 136.200 26.330 136.800 ;
        RECT 25.930 136.000 29.930 136.200 ;
        RECT 25.930 135.400 26.330 136.000 ;
        RECT 25.930 135.200 29.930 135.400 ;
        RECT 25.930 134.600 26.330 135.200 ;
        RECT 25.930 134.400 29.930 134.600 ;
        RECT 25.930 133.800 26.330 134.400 ;
        RECT 25.930 133.600 29.930 133.800 ;
        RECT 25.930 133.000 26.330 133.600 ;
        RECT 25.930 132.800 29.930 133.000 ;
        RECT 25.930 132.200 26.330 132.800 ;
        RECT 25.930 132.000 29.930 132.200 ;
        RECT 25.930 131.400 26.330 132.000 ;
        RECT 25.930 131.200 29.930 131.400 ;
        RECT 25.930 130.600 26.330 131.200 ;
        RECT 25.930 130.400 29.930 130.600 ;
        RECT 25.930 130.200 26.330 130.400 ;
        RECT 30.680 130.200 30.880 137.800 ;
        RECT 31.480 130.200 31.680 137.800 ;
        RECT 32.280 130.200 32.480 137.800 ;
        RECT 33.080 130.200 33.280 137.800 ;
        RECT 33.880 130.200 34.080 137.800 ;
        RECT 25.930 129.800 34.080 130.200 ;
        RECT 25.930 129.600 26.330 129.800 ;
        RECT 25.930 129.400 29.930 129.600 ;
        RECT 25.930 128.800 26.330 129.400 ;
        RECT 25.930 128.600 29.930 128.800 ;
        RECT 25.930 128.000 26.330 128.600 ;
        RECT 25.930 127.800 29.930 128.000 ;
        RECT 25.930 127.200 26.330 127.800 ;
        RECT 25.930 127.000 29.930 127.200 ;
        RECT 25.930 126.400 26.330 127.000 ;
        RECT 25.930 126.200 29.930 126.400 ;
        RECT 25.930 125.600 26.330 126.200 ;
        RECT 25.930 125.400 29.930 125.600 ;
        RECT 25.930 124.800 26.330 125.400 ;
        RECT 25.930 124.600 29.930 124.800 ;
        RECT 25.930 124.000 26.330 124.600 ;
        RECT 25.930 123.800 29.930 124.000 ;
        RECT 25.930 123.200 26.330 123.800 ;
        RECT 25.930 123.000 29.930 123.200 ;
        RECT 25.930 122.400 26.330 123.000 ;
        RECT 25.930 122.200 29.930 122.400 ;
        RECT 30.680 122.200 30.880 129.800 ;
        RECT 31.480 122.200 31.680 129.800 ;
        RECT 32.280 122.200 32.480 129.800 ;
        RECT 33.080 122.200 33.280 129.800 ;
        RECT 33.880 122.200 34.080 129.800 ;
        RECT 35.380 130.200 35.580 137.800 ;
        RECT 36.180 130.200 36.380 137.800 ;
        RECT 36.980 130.200 37.180 137.800 ;
        RECT 37.780 130.200 37.980 137.800 ;
        RECT 38.580 130.200 38.780 137.800 ;
        RECT 39.530 137.600 43.530 137.800 ;
        RECT 43.130 137.000 43.530 137.600 ;
        RECT 39.530 136.800 43.530 137.000 ;
        RECT 43.130 136.200 43.530 136.800 ;
        RECT 39.530 136.000 43.530 136.200 ;
        RECT 43.130 135.400 43.530 136.000 ;
        RECT 39.530 135.200 43.530 135.400 ;
        RECT 43.130 134.600 43.530 135.200 ;
        RECT 39.530 134.400 43.530 134.600 ;
        RECT 43.130 133.800 43.530 134.400 ;
        RECT 39.530 133.600 43.530 133.800 ;
        RECT 43.130 133.000 43.530 133.600 ;
        RECT 39.530 132.800 43.530 133.000 ;
        RECT 43.130 132.200 43.530 132.800 ;
        RECT 39.530 132.000 43.530 132.200 ;
        RECT 43.130 131.400 43.530 132.000 ;
        RECT 39.530 131.200 43.530 131.400 ;
        RECT 43.130 130.600 43.530 131.200 ;
        RECT 39.530 130.400 43.530 130.600 ;
        RECT 43.130 130.200 43.530 130.400 ;
        RECT 35.380 129.800 43.530 130.200 ;
        RECT 35.380 122.200 35.580 129.800 ;
        RECT 36.180 122.200 36.380 129.800 ;
        RECT 36.980 122.200 37.180 129.800 ;
        RECT 37.780 122.200 37.980 129.800 ;
        RECT 38.580 122.200 38.780 129.800 ;
        RECT 43.130 129.600 43.530 129.800 ;
        RECT 39.530 129.400 43.530 129.600 ;
        RECT 43.130 128.800 43.530 129.400 ;
        RECT 39.530 128.600 43.530 128.800 ;
        RECT 43.130 128.000 43.530 128.600 ;
        RECT 39.530 127.800 43.530 128.000 ;
        RECT 43.130 127.200 43.530 127.800 ;
        RECT 39.530 127.000 43.530 127.200 ;
        RECT 43.130 126.400 43.530 127.000 ;
        RECT 39.530 126.200 43.530 126.400 ;
        RECT 43.130 125.600 43.530 126.200 ;
        RECT 39.530 125.400 43.530 125.600 ;
        RECT 43.130 124.800 43.530 125.400 ;
        RECT 39.530 124.600 43.530 124.800 ;
        RECT 43.130 124.000 43.530 124.600 ;
        RECT 39.530 123.800 43.530 124.000 ;
        RECT 43.130 123.200 43.530 123.800 ;
        RECT 39.530 123.000 43.530 123.200 ;
        RECT 43.130 122.400 43.530 123.000 ;
        RECT 39.530 122.200 43.530 122.400 ;
        RECT 45.930 137.600 49.930 137.800 ;
        RECT 45.930 137.000 46.330 137.600 ;
        RECT 45.930 136.800 49.930 137.000 ;
        RECT 45.930 136.200 46.330 136.800 ;
        RECT 45.930 136.000 49.930 136.200 ;
        RECT 45.930 135.400 46.330 136.000 ;
        RECT 45.930 135.200 49.930 135.400 ;
        RECT 45.930 134.600 46.330 135.200 ;
        RECT 45.930 134.400 49.930 134.600 ;
        RECT 45.930 133.800 46.330 134.400 ;
        RECT 45.930 133.600 49.930 133.800 ;
        RECT 45.930 133.000 46.330 133.600 ;
        RECT 45.930 132.800 49.930 133.000 ;
        RECT 45.930 132.200 46.330 132.800 ;
        RECT 45.930 132.000 49.930 132.200 ;
        RECT 45.930 131.400 46.330 132.000 ;
        RECT 45.930 131.200 49.930 131.400 ;
        RECT 45.930 130.600 46.330 131.200 ;
        RECT 45.930 130.400 49.930 130.600 ;
        RECT 45.930 130.200 46.330 130.400 ;
        RECT 50.680 130.200 50.880 137.800 ;
        RECT 51.480 130.200 51.680 137.800 ;
        RECT 52.280 130.200 52.480 137.800 ;
        RECT 53.080 130.200 53.280 137.800 ;
        RECT 53.880 130.200 54.080 137.800 ;
        RECT 45.930 129.800 54.080 130.200 ;
        RECT 45.930 129.600 46.330 129.800 ;
        RECT 45.930 129.400 49.930 129.600 ;
        RECT 45.930 128.800 46.330 129.400 ;
        RECT 45.930 128.600 49.930 128.800 ;
        RECT 45.930 128.000 46.330 128.600 ;
        RECT 45.930 127.800 49.930 128.000 ;
        RECT 45.930 127.200 46.330 127.800 ;
        RECT 45.930 127.000 49.930 127.200 ;
        RECT 45.930 126.400 46.330 127.000 ;
        RECT 45.930 126.200 49.930 126.400 ;
        RECT 45.930 125.600 46.330 126.200 ;
        RECT 45.930 125.400 49.930 125.600 ;
        RECT 45.930 124.800 46.330 125.400 ;
        RECT 45.930 124.600 49.930 124.800 ;
        RECT 45.930 124.000 46.330 124.600 ;
        RECT 45.930 123.800 49.930 124.000 ;
        RECT 45.930 123.200 46.330 123.800 ;
        RECT 45.930 123.000 49.930 123.200 ;
        RECT 45.930 122.400 46.330 123.000 ;
        RECT 45.930 122.200 49.930 122.400 ;
        RECT 50.680 122.200 50.880 129.800 ;
        RECT 51.480 122.200 51.680 129.800 ;
        RECT 52.280 122.200 52.480 129.800 ;
        RECT 53.080 122.200 53.280 129.800 ;
        RECT 53.880 122.200 54.080 129.800 ;
        RECT 55.380 130.200 55.580 137.800 ;
        RECT 56.180 130.200 56.380 137.800 ;
        RECT 56.980 130.200 57.180 137.800 ;
        RECT 57.780 130.200 57.980 137.800 ;
        RECT 58.580 130.200 58.780 137.800 ;
        RECT 59.530 137.600 63.530 137.800 ;
        RECT 63.130 137.000 63.530 137.600 ;
        RECT 59.530 136.800 63.530 137.000 ;
        RECT 63.130 136.200 63.530 136.800 ;
        RECT 59.530 136.000 63.530 136.200 ;
        RECT 63.130 135.400 63.530 136.000 ;
        RECT 59.530 135.200 63.530 135.400 ;
        RECT 63.130 134.600 63.530 135.200 ;
        RECT 59.530 134.400 63.530 134.600 ;
        RECT 63.130 133.800 63.530 134.400 ;
        RECT 59.530 133.600 63.530 133.800 ;
        RECT 63.130 133.000 63.530 133.600 ;
        RECT 59.530 132.800 63.530 133.000 ;
        RECT 63.130 132.200 63.530 132.800 ;
        RECT 59.530 132.000 63.530 132.200 ;
        RECT 63.130 131.400 63.530 132.000 ;
        RECT 59.530 131.200 63.530 131.400 ;
        RECT 63.130 130.600 63.530 131.200 ;
        RECT 59.530 130.400 63.530 130.600 ;
        RECT 63.130 130.200 63.530 130.400 ;
        RECT 55.380 129.800 63.530 130.200 ;
        RECT 55.380 122.200 55.580 129.800 ;
        RECT 56.180 122.200 56.380 129.800 ;
        RECT 56.980 122.200 57.180 129.800 ;
        RECT 57.780 122.200 57.980 129.800 ;
        RECT 58.580 122.200 58.780 129.800 ;
        RECT 63.130 129.600 63.530 129.800 ;
        RECT 59.530 129.400 63.530 129.600 ;
        RECT 63.130 128.800 63.530 129.400 ;
        RECT 59.530 128.600 63.530 128.800 ;
        RECT 63.130 128.000 63.530 128.600 ;
        RECT 59.530 127.800 63.530 128.000 ;
        RECT 63.130 127.200 63.530 127.800 ;
        RECT 59.530 127.000 63.530 127.200 ;
        RECT 63.130 126.400 63.530 127.000 ;
        RECT 59.530 126.200 63.530 126.400 ;
        RECT 63.130 125.600 63.530 126.200 ;
        RECT 59.530 125.400 63.530 125.600 ;
        RECT 63.130 124.800 63.530 125.400 ;
        RECT 59.530 124.600 63.530 124.800 ;
        RECT 63.130 124.000 63.530 124.600 ;
        RECT 59.530 123.800 63.530 124.000 ;
        RECT 63.130 123.200 63.530 123.800 ;
        RECT 59.530 123.000 63.530 123.200 ;
        RECT 63.130 122.400 63.530 123.000 ;
        RECT 59.530 122.200 63.530 122.400 ;
        RECT 65.930 137.600 69.930 137.800 ;
        RECT 65.930 137.000 66.330 137.600 ;
        RECT 65.930 136.800 69.930 137.000 ;
        RECT 65.930 136.200 66.330 136.800 ;
        RECT 65.930 136.000 69.930 136.200 ;
        RECT 65.930 135.400 66.330 136.000 ;
        RECT 65.930 135.200 69.930 135.400 ;
        RECT 65.930 134.600 66.330 135.200 ;
        RECT 65.930 134.400 69.930 134.600 ;
        RECT 65.930 133.800 66.330 134.400 ;
        RECT 65.930 133.600 69.930 133.800 ;
        RECT 65.930 133.000 66.330 133.600 ;
        RECT 65.930 132.800 69.930 133.000 ;
        RECT 65.930 132.200 66.330 132.800 ;
        RECT 65.930 132.000 69.930 132.200 ;
        RECT 65.930 131.400 66.330 132.000 ;
        RECT 65.930 131.200 69.930 131.400 ;
        RECT 65.930 130.600 66.330 131.200 ;
        RECT 65.930 130.400 69.930 130.600 ;
        RECT 65.930 130.200 66.330 130.400 ;
        RECT 70.680 130.200 70.880 137.800 ;
        RECT 71.480 130.200 71.680 137.800 ;
        RECT 72.280 130.200 72.480 137.800 ;
        RECT 73.080 130.200 73.280 137.800 ;
        RECT 73.880 130.200 74.080 137.800 ;
        RECT 65.930 129.800 74.080 130.200 ;
        RECT 65.930 129.600 66.330 129.800 ;
        RECT 65.930 129.400 69.930 129.600 ;
        RECT 65.930 128.800 66.330 129.400 ;
        RECT 65.930 128.600 69.930 128.800 ;
        RECT 65.930 128.000 66.330 128.600 ;
        RECT 65.930 127.800 69.930 128.000 ;
        RECT 65.930 127.200 66.330 127.800 ;
        RECT 65.930 127.000 69.930 127.200 ;
        RECT 65.930 126.400 66.330 127.000 ;
        RECT 65.930 126.200 69.930 126.400 ;
        RECT 65.930 125.600 66.330 126.200 ;
        RECT 65.930 125.400 69.930 125.600 ;
        RECT 65.930 124.800 66.330 125.400 ;
        RECT 65.930 124.600 69.930 124.800 ;
        RECT 65.930 124.000 66.330 124.600 ;
        RECT 65.930 123.800 69.930 124.000 ;
        RECT 65.930 123.200 66.330 123.800 ;
        RECT 65.930 123.000 69.930 123.200 ;
        RECT 65.930 122.400 66.330 123.000 ;
        RECT 65.930 122.200 69.930 122.400 ;
        RECT 70.680 122.200 70.880 129.800 ;
        RECT 71.480 122.200 71.680 129.800 ;
        RECT 72.280 122.200 72.480 129.800 ;
        RECT 73.080 122.200 73.280 129.800 ;
        RECT 73.880 122.200 74.080 129.800 ;
        RECT 75.380 130.200 75.580 137.800 ;
        RECT 76.180 130.200 76.380 137.800 ;
        RECT 76.980 130.200 77.180 137.800 ;
        RECT 77.780 130.200 77.980 137.800 ;
        RECT 78.580 130.200 78.780 137.800 ;
        RECT 79.530 137.600 83.530 137.800 ;
        RECT 83.130 137.000 83.530 137.600 ;
        RECT 79.530 136.800 83.530 137.000 ;
        RECT 83.130 136.200 83.530 136.800 ;
        RECT 79.530 136.000 83.530 136.200 ;
        RECT 83.130 135.400 83.530 136.000 ;
        RECT 79.530 135.200 83.530 135.400 ;
        RECT 83.130 134.600 83.530 135.200 ;
        RECT 79.530 134.400 83.530 134.600 ;
        RECT 83.130 133.800 83.530 134.400 ;
        RECT 79.530 133.600 83.530 133.800 ;
        RECT 83.130 133.000 83.530 133.600 ;
        RECT 79.530 132.800 83.530 133.000 ;
        RECT 83.130 132.200 83.530 132.800 ;
        RECT 79.530 132.000 83.530 132.200 ;
        RECT 83.130 131.400 83.530 132.000 ;
        RECT 79.530 131.200 83.530 131.400 ;
        RECT 83.130 130.600 83.530 131.200 ;
        RECT 79.530 130.400 83.530 130.600 ;
        RECT 83.130 130.200 83.530 130.400 ;
        RECT 75.380 129.800 83.530 130.200 ;
        RECT 75.380 122.200 75.580 129.800 ;
        RECT 76.180 122.200 76.380 129.800 ;
        RECT 76.980 122.200 77.180 129.800 ;
        RECT 77.780 122.200 77.980 129.800 ;
        RECT 78.580 122.200 78.780 129.800 ;
        RECT 83.130 129.600 83.530 129.800 ;
        RECT 79.530 129.400 83.530 129.600 ;
        RECT 83.130 128.800 83.530 129.400 ;
        RECT 79.530 128.600 83.530 128.800 ;
        RECT 83.130 128.000 83.530 128.600 ;
        RECT 79.530 127.800 83.530 128.000 ;
        RECT 83.130 127.200 83.530 127.800 ;
        RECT 79.530 127.000 83.530 127.200 ;
        RECT 83.130 126.400 83.530 127.000 ;
        RECT 79.530 126.200 83.530 126.400 ;
        RECT 83.130 125.600 83.530 126.200 ;
        RECT 79.530 125.400 83.530 125.600 ;
        RECT 83.130 124.800 83.530 125.400 ;
        RECT 79.530 124.600 83.530 124.800 ;
        RECT 83.130 124.000 83.530 124.600 ;
        RECT 79.530 123.800 83.530 124.000 ;
        RECT 83.130 123.200 83.530 123.800 ;
        RECT 79.530 123.000 83.530 123.200 ;
        RECT 83.130 122.400 83.530 123.000 ;
        RECT 79.530 122.200 83.530 122.400 ;
        RECT 85.930 137.600 89.930 137.800 ;
        RECT 85.930 137.000 86.330 137.600 ;
        RECT 85.930 136.800 89.930 137.000 ;
        RECT 85.930 136.200 86.330 136.800 ;
        RECT 85.930 136.000 89.930 136.200 ;
        RECT 85.930 135.400 86.330 136.000 ;
        RECT 85.930 135.200 89.930 135.400 ;
        RECT 85.930 134.600 86.330 135.200 ;
        RECT 85.930 134.400 89.930 134.600 ;
        RECT 85.930 133.800 86.330 134.400 ;
        RECT 85.930 133.600 89.930 133.800 ;
        RECT 85.930 133.000 86.330 133.600 ;
        RECT 85.930 132.800 89.930 133.000 ;
        RECT 85.930 132.200 86.330 132.800 ;
        RECT 85.930 132.000 89.930 132.200 ;
        RECT 85.930 131.400 86.330 132.000 ;
        RECT 85.930 131.200 89.930 131.400 ;
        RECT 85.930 130.600 86.330 131.200 ;
        RECT 85.930 130.400 89.930 130.600 ;
        RECT 85.930 130.200 86.330 130.400 ;
        RECT 90.680 130.200 90.880 137.800 ;
        RECT 91.480 130.200 91.680 137.800 ;
        RECT 92.280 130.200 92.480 137.800 ;
        RECT 93.080 130.200 93.280 137.800 ;
        RECT 93.880 130.200 94.080 137.800 ;
        RECT 85.930 129.800 94.080 130.200 ;
        RECT 85.930 129.600 86.330 129.800 ;
        RECT 85.930 129.400 89.930 129.600 ;
        RECT 85.930 128.800 86.330 129.400 ;
        RECT 85.930 128.600 89.930 128.800 ;
        RECT 85.930 128.000 86.330 128.600 ;
        RECT 85.930 127.800 89.930 128.000 ;
        RECT 85.930 127.200 86.330 127.800 ;
        RECT 85.930 127.000 89.930 127.200 ;
        RECT 85.930 126.400 86.330 127.000 ;
        RECT 85.930 126.200 89.930 126.400 ;
        RECT 85.930 125.600 86.330 126.200 ;
        RECT 85.930 125.400 89.930 125.600 ;
        RECT 85.930 124.800 86.330 125.400 ;
        RECT 85.930 124.600 89.930 124.800 ;
        RECT 85.930 124.000 86.330 124.600 ;
        RECT 85.930 123.800 89.930 124.000 ;
        RECT 85.930 123.200 86.330 123.800 ;
        RECT 85.930 123.000 89.930 123.200 ;
        RECT 85.930 122.400 86.330 123.000 ;
        RECT 85.930 122.200 89.930 122.400 ;
        RECT 90.680 122.200 90.880 129.800 ;
        RECT 91.480 122.200 91.680 129.800 ;
        RECT 92.280 122.200 92.480 129.800 ;
        RECT 93.080 122.200 93.280 129.800 ;
        RECT 93.880 122.200 94.080 129.800 ;
        RECT 95.380 130.200 95.580 137.800 ;
        RECT 96.180 130.200 96.380 137.800 ;
        RECT 96.980 130.200 97.180 137.800 ;
        RECT 97.780 130.200 97.980 137.800 ;
        RECT 98.580 130.200 98.780 137.800 ;
        RECT 99.530 137.600 103.530 137.800 ;
        RECT 103.130 137.000 103.530 137.600 ;
        RECT 99.530 136.800 103.530 137.000 ;
        RECT 103.130 136.200 103.530 136.800 ;
        RECT 99.530 136.000 103.530 136.200 ;
        RECT 103.130 135.400 103.530 136.000 ;
        RECT 99.530 135.200 103.530 135.400 ;
        RECT 103.130 134.600 103.530 135.200 ;
        RECT 99.530 134.400 103.530 134.600 ;
        RECT 103.130 133.800 103.530 134.400 ;
        RECT 99.530 133.600 103.530 133.800 ;
        RECT 103.130 133.000 103.530 133.600 ;
        RECT 99.530 132.800 103.530 133.000 ;
        RECT 103.130 132.200 103.530 132.800 ;
        RECT 99.530 132.000 103.530 132.200 ;
        RECT 103.130 131.400 103.530 132.000 ;
        RECT 99.530 131.200 103.530 131.400 ;
        RECT 103.130 130.600 103.530 131.200 ;
        RECT 99.530 130.400 103.530 130.600 ;
        RECT 103.130 130.200 103.530 130.400 ;
        RECT 95.380 129.800 103.530 130.200 ;
        RECT 95.380 122.200 95.580 129.800 ;
        RECT 96.180 122.200 96.380 129.800 ;
        RECT 96.980 122.200 97.180 129.800 ;
        RECT 97.780 122.200 97.980 129.800 ;
        RECT 98.580 122.200 98.780 129.800 ;
        RECT 103.130 129.600 103.530 129.800 ;
        RECT 99.530 129.400 103.530 129.600 ;
        RECT 110.050 129.475 110.410 129.855 ;
        RECT 110.680 129.475 111.040 129.855 ;
        RECT 111.280 129.475 111.640 129.855 ;
        RECT 103.130 128.800 103.530 129.400 ;
        RECT 110.050 128.885 110.410 129.265 ;
        RECT 110.680 128.885 111.040 129.265 ;
        RECT 111.280 128.885 111.640 129.265 ;
        RECT 99.530 128.600 103.530 128.800 ;
        RECT 103.130 128.000 103.530 128.600 ;
        RECT 99.530 127.800 103.530 128.000 ;
        RECT 103.130 127.200 103.530 127.800 ;
        RECT 99.530 127.000 103.530 127.200 ;
        RECT 103.130 126.400 103.530 127.000 ;
        RECT 99.530 126.200 103.530 126.400 ;
        RECT 103.130 125.600 103.530 126.200 ;
        RECT 99.530 125.400 103.530 125.600 ;
        RECT 103.130 124.800 103.530 125.400 ;
        RECT 99.530 124.600 103.530 124.800 ;
        RECT 103.130 124.000 103.530 124.600 ;
        RECT 99.530 123.800 103.530 124.000 ;
        RECT 103.130 123.200 103.530 123.800 ;
        RECT 99.530 123.000 103.530 123.200 ;
        RECT 103.130 122.400 103.530 123.000 ;
        RECT 99.530 122.200 103.530 122.400 ;
        RECT 5.930 117.600 9.930 117.800 ;
        RECT 5.930 117.000 6.330 117.600 ;
        RECT 5.930 116.800 9.930 117.000 ;
        RECT 5.930 116.200 6.330 116.800 ;
        RECT 5.930 116.000 9.930 116.200 ;
        RECT 5.930 115.400 6.330 116.000 ;
        RECT 5.930 115.200 9.930 115.400 ;
        RECT 5.930 114.600 6.330 115.200 ;
        RECT 5.930 114.400 9.930 114.600 ;
        RECT 5.930 113.800 6.330 114.400 ;
        RECT 5.930 113.600 9.930 113.800 ;
        RECT 5.930 113.000 6.330 113.600 ;
        RECT 5.930 112.800 9.930 113.000 ;
        RECT 5.930 112.200 6.330 112.800 ;
        RECT 5.930 112.000 9.930 112.200 ;
        RECT 5.930 111.400 6.330 112.000 ;
        RECT 5.930 111.200 9.930 111.400 ;
        RECT 5.930 110.600 6.330 111.200 ;
        RECT 5.930 110.400 9.930 110.600 ;
        RECT 5.930 110.200 6.330 110.400 ;
        RECT 10.680 110.200 10.880 117.800 ;
        RECT 11.480 110.200 11.680 117.800 ;
        RECT 12.280 110.200 12.480 117.800 ;
        RECT 13.080 110.200 13.280 117.800 ;
        RECT 13.880 110.200 14.080 117.800 ;
        RECT 5.930 109.800 14.080 110.200 ;
        RECT 5.930 109.600 6.330 109.800 ;
        RECT 5.930 109.400 9.930 109.600 ;
        RECT 5.930 108.800 6.330 109.400 ;
        RECT 5.930 108.600 9.930 108.800 ;
        RECT 5.930 108.000 6.330 108.600 ;
        RECT 5.930 107.800 9.930 108.000 ;
        RECT 5.930 107.200 6.330 107.800 ;
        RECT 5.930 107.000 9.930 107.200 ;
        RECT 5.930 106.400 6.330 107.000 ;
        RECT 5.930 106.200 9.930 106.400 ;
        RECT 5.930 105.600 6.330 106.200 ;
        RECT 5.930 105.400 9.930 105.600 ;
        RECT 5.930 104.800 6.330 105.400 ;
        RECT 5.930 104.600 9.930 104.800 ;
        RECT 5.930 104.000 6.330 104.600 ;
        RECT 5.930 103.800 9.930 104.000 ;
        RECT 5.930 103.200 6.330 103.800 ;
        RECT 5.930 103.000 9.930 103.200 ;
        RECT 5.930 102.400 6.330 103.000 ;
        RECT 5.930 102.200 9.930 102.400 ;
        RECT 10.680 102.200 10.880 109.800 ;
        RECT 11.480 102.200 11.680 109.800 ;
        RECT 12.280 102.200 12.480 109.800 ;
        RECT 13.080 102.200 13.280 109.800 ;
        RECT 13.880 102.200 14.080 109.800 ;
        RECT 15.380 110.200 15.580 117.800 ;
        RECT 16.180 110.200 16.380 117.800 ;
        RECT 16.980 110.200 17.180 117.800 ;
        RECT 17.780 110.200 17.980 117.800 ;
        RECT 18.580 110.200 18.780 117.800 ;
        RECT 19.530 117.600 23.530 117.800 ;
        RECT 23.130 117.000 23.530 117.600 ;
        RECT 19.530 116.800 23.530 117.000 ;
        RECT 23.130 116.200 23.530 116.800 ;
        RECT 19.530 116.000 23.530 116.200 ;
        RECT 23.130 115.400 23.530 116.000 ;
        RECT 19.530 115.200 23.530 115.400 ;
        RECT 23.130 114.600 23.530 115.200 ;
        RECT 19.530 114.400 23.530 114.600 ;
        RECT 23.130 113.800 23.530 114.400 ;
        RECT 19.530 113.600 23.530 113.800 ;
        RECT 23.130 113.000 23.530 113.600 ;
        RECT 19.530 112.800 23.530 113.000 ;
        RECT 23.130 112.200 23.530 112.800 ;
        RECT 19.530 112.000 23.530 112.200 ;
        RECT 23.130 111.400 23.530 112.000 ;
        RECT 19.530 111.200 23.530 111.400 ;
        RECT 23.130 110.600 23.530 111.200 ;
        RECT 19.530 110.400 23.530 110.600 ;
        RECT 23.130 110.200 23.530 110.400 ;
        RECT 15.380 109.800 23.530 110.200 ;
        RECT 15.380 102.200 15.580 109.800 ;
        RECT 16.180 102.200 16.380 109.800 ;
        RECT 16.980 102.200 17.180 109.800 ;
        RECT 17.780 102.200 17.980 109.800 ;
        RECT 18.580 102.200 18.780 109.800 ;
        RECT 23.130 109.600 23.530 109.800 ;
        RECT 19.530 109.400 23.530 109.600 ;
        RECT 23.130 108.800 23.530 109.400 ;
        RECT 19.530 108.600 23.530 108.800 ;
        RECT 23.130 108.000 23.530 108.600 ;
        RECT 19.530 107.800 23.530 108.000 ;
        RECT 23.130 107.200 23.530 107.800 ;
        RECT 19.530 107.000 23.530 107.200 ;
        RECT 23.130 106.400 23.530 107.000 ;
        RECT 19.530 106.200 23.530 106.400 ;
        RECT 23.130 105.600 23.530 106.200 ;
        RECT 19.530 105.400 23.530 105.600 ;
        RECT 23.130 104.800 23.530 105.400 ;
        RECT 19.530 104.600 23.530 104.800 ;
        RECT 23.130 104.000 23.530 104.600 ;
        RECT 19.530 103.800 23.530 104.000 ;
        RECT 23.130 103.200 23.530 103.800 ;
        RECT 19.530 103.000 23.530 103.200 ;
        RECT 23.130 102.400 23.530 103.000 ;
        RECT 19.530 102.200 23.530 102.400 ;
        RECT 25.930 117.600 29.930 117.800 ;
        RECT 25.930 117.000 26.330 117.600 ;
        RECT 25.930 116.800 29.930 117.000 ;
        RECT 25.930 116.200 26.330 116.800 ;
        RECT 25.930 116.000 29.930 116.200 ;
        RECT 25.930 115.400 26.330 116.000 ;
        RECT 25.930 115.200 29.930 115.400 ;
        RECT 25.930 114.600 26.330 115.200 ;
        RECT 25.930 114.400 29.930 114.600 ;
        RECT 25.930 113.800 26.330 114.400 ;
        RECT 25.930 113.600 29.930 113.800 ;
        RECT 25.930 113.000 26.330 113.600 ;
        RECT 25.930 112.800 29.930 113.000 ;
        RECT 25.930 112.200 26.330 112.800 ;
        RECT 25.930 112.000 29.930 112.200 ;
        RECT 25.930 111.400 26.330 112.000 ;
        RECT 25.930 111.200 29.930 111.400 ;
        RECT 25.930 110.600 26.330 111.200 ;
        RECT 25.930 110.400 29.930 110.600 ;
        RECT 25.930 110.200 26.330 110.400 ;
        RECT 30.680 110.200 30.880 117.800 ;
        RECT 31.480 110.200 31.680 117.800 ;
        RECT 32.280 110.200 32.480 117.800 ;
        RECT 33.080 110.200 33.280 117.800 ;
        RECT 33.880 110.200 34.080 117.800 ;
        RECT 25.930 109.800 34.080 110.200 ;
        RECT 25.930 109.600 26.330 109.800 ;
        RECT 25.930 109.400 29.930 109.600 ;
        RECT 25.930 108.800 26.330 109.400 ;
        RECT 25.930 108.600 29.930 108.800 ;
        RECT 25.930 108.000 26.330 108.600 ;
        RECT 25.930 107.800 29.930 108.000 ;
        RECT 25.930 107.200 26.330 107.800 ;
        RECT 25.930 107.000 29.930 107.200 ;
        RECT 25.930 106.400 26.330 107.000 ;
        RECT 25.930 106.200 29.930 106.400 ;
        RECT 25.930 105.600 26.330 106.200 ;
        RECT 25.930 105.400 29.930 105.600 ;
        RECT 25.930 104.800 26.330 105.400 ;
        RECT 25.930 104.600 29.930 104.800 ;
        RECT 25.930 104.000 26.330 104.600 ;
        RECT 25.930 103.800 29.930 104.000 ;
        RECT 25.930 103.200 26.330 103.800 ;
        RECT 25.930 103.000 29.930 103.200 ;
        RECT 25.930 102.400 26.330 103.000 ;
        RECT 25.930 102.200 29.930 102.400 ;
        RECT 30.680 102.200 30.880 109.800 ;
        RECT 31.480 102.200 31.680 109.800 ;
        RECT 32.280 102.200 32.480 109.800 ;
        RECT 33.080 102.200 33.280 109.800 ;
        RECT 33.880 102.200 34.080 109.800 ;
        RECT 35.380 110.200 35.580 117.800 ;
        RECT 36.180 110.200 36.380 117.800 ;
        RECT 36.980 110.200 37.180 117.800 ;
        RECT 37.780 110.200 37.980 117.800 ;
        RECT 38.580 110.200 38.780 117.800 ;
        RECT 39.530 117.600 43.530 117.800 ;
        RECT 43.130 117.000 43.530 117.600 ;
        RECT 39.530 116.800 43.530 117.000 ;
        RECT 43.130 116.200 43.530 116.800 ;
        RECT 39.530 116.000 43.530 116.200 ;
        RECT 43.130 115.400 43.530 116.000 ;
        RECT 39.530 115.200 43.530 115.400 ;
        RECT 43.130 114.600 43.530 115.200 ;
        RECT 39.530 114.400 43.530 114.600 ;
        RECT 43.130 113.800 43.530 114.400 ;
        RECT 39.530 113.600 43.530 113.800 ;
        RECT 43.130 113.000 43.530 113.600 ;
        RECT 39.530 112.800 43.530 113.000 ;
        RECT 43.130 112.200 43.530 112.800 ;
        RECT 39.530 112.000 43.530 112.200 ;
        RECT 43.130 111.400 43.530 112.000 ;
        RECT 39.530 111.200 43.530 111.400 ;
        RECT 43.130 110.600 43.530 111.200 ;
        RECT 39.530 110.400 43.530 110.600 ;
        RECT 43.130 110.200 43.530 110.400 ;
        RECT 35.380 109.800 43.530 110.200 ;
        RECT 35.380 102.200 35.580 109.800 ;
        RECT 36.180 102.200 36.380 109.800 ;
        RECT 36.980 102.200 37.180 109.800 ;
        RECT 37.780 102.200 37.980 109.800 ;
        RECT 38.580 102.200 38.780 109.800 ;
        RECT 43.130 109.600 43.530 109.800 ;
        RECT 39.530 109.400 43.530 109.600 ;
        RECT 43.130 108.800 43.530 109.400 ;
        RECT 39.530 108.600 43.530 108.800 ;
        RECT 43.130 108.000 43.530 108.600 ;
        RECT 39.530 107.800 43.530 108.000 ;
        RECT 43.130 107.200 43.530 107.800 ;
        RECT 39.530 107.000 43.530 107.200 ;
        RECT 43.130 106.400 43.530 107.000 ;
        RECT 39.530 106.200 43.530 106.400 ;
        RECT 43.130 105.600 43.530 106.200 ;
        RECT 39.530 105.400 43.530 105.600 ;
        RECT 43.130 104.800 43.530 105.400 ;
        RECT 39.530 104.600 43.530 104.800 ;
        RECT 43.130 104.000 43.530 104.600 ;
        RECT 39.530 103.800 43.530 104.000 ;
        RECT 43.130 103.200 43.530 103.800 ;
        RECT 39.530 103.000 43.530 103.200 ;
        RECT 43.130 102.400 43.530 103.000 ;
        RECT 39.530 102.200 43.530 102.400 ;
        RECT 45.930 117.600 49.930 117.800 ;
        RECT 45.930 117.000 46.330 117.600 ;
        RECT 45.930 116.800 49.930 117.000 ;
        RECT 45.930 116.200 46.330 116.800 ;
        RECT 45.930 116.000 49.930 116.200 ;
        RECT 45.930 115.400 46.330 116.000 ;
        RECT 45.930 115.200 49.930 115.400 ;
        RECT 45.930 114.600 46.330 115.200 ;
        RECT 45.930 114.400 49.930 114.600 ;
        RECT 45.930 113.800 46.330 114.400 ;
        RECT 45.930 113.600 49.930 113.800 ;
        RECT 45.930 113.000 46.330 113.600 ;
        RECT 45.930 112.800 49.930 113.000 ;
        RECT 45.930 112.200 46.330 112.800 ;
        RECT 45.930 112.000 49.930 112.200 ;
        RECT 45.930 111.400 46.330 112.000 ;
        RECT 45.930 111.200 49.930 111.400 ;
        RECT 45.930 110.600 46.330 111.200 ;
        RECT 45.930 110.400 49.930 110.600 ;
        RECT 45.930 110.200 46.330 110.400 ;
        RECT 50.680 110.200 50.880 117.800 ;
        RECT 51.480 110.200 51.680 117.800 ;
        RECT 52.280 110.200 52.480 117.800 ;
        RECT 53.080 110.200 53.280 117.800 ;
        RECT 53.880 110.200 54.080 117.800 ;
        RECT 45.930 109.800 54.080 110.200 ;
        RECT 45.930 109.600 46.330 109.800 ;
        RECT 45.930 109.400 49.930 109.600 ;
        RECT 45.930 108.800 46.330 109.400 ;
        RECT 45.930 108.600 49.930 108.800 ;
        RECT 45.930 108.000 46.330 108.600 ;
        RECT 45.930 107.800 49.930 108.000 ;
        RECT 45.930 107.200 46.330 107.800 ;
        RECT 45.930 107.000 49.930 107.200 ;
        RECT 45.930 106.400 46.330 107.000 ;
        RECT 45.930 106.200 49.930 106.400 ;
        RECT 45.930 105.600 46.330 106.200 ;
        RECT 45.930 105.400 49.930 105.600 ;
        RECT 45.930 104.800 46.330 105.400 ;
        RECT 45.930 104.600 49.930 104.800 ;
        RECT 45.930 104.000 46.330 104.600 ;
        RECT 45.930 103.800 49.930 104.000 ;
        RECT 45.930 103.200 46.330 103.800 ;
        RECT 45.930 103.000 49.930 103.200 ;
        RECT 45.930 102.400 46.330 103.000 ;
        RECT 45.930 102.200 49.930 102.400 ;
        RECT 50.680 102.200 50.880 109.800 ;
        RECT 51.480 102.200 51.680 109.800 ;
        RECT 52.280 102.200 52.480 109.800 ;
        RECT 53.080 102.200 53.280 109.800 ;
        RECT 53.880 102.200 54.080 109.800 ;
        RECT 55.380 110.200 55.580 117.800 ;
        RECT 56.180 110.200 56.380 117.800 ;
        RECT 56.980 110.200 57.180 117.800 ;
        RECT 57.780 110.200 57.980 117.800 ;
        RECT 58.580 110.200 58.780 117.800 ;
        RECT 59.530 117.600 63.530 117.800 ;
        RECT 63.130 117.000 63.530 117.600 ;
        RECT 59.530 116.800 63.530 117.000 ;
        RECT 63.130 116.200 63.530 116.800 ;
        RECT 59.530 116.000 63.530 116.200 ;
        RECT 63.130 115.400 63.530 116.000 ;
        RECT 59.530 115.200 63.530 115.400 ;
        RECT 63.130 114.600 63.530 115.200 ;
        RECT 59.530 114.400 63.530 114.600 ;
        RECT 63.130 113.800 63.530 114.400 ;
        RECT 59.530 113.600 63.530 113.800 ;
        RECT 63.130 113.000 63.530 113.600 ;
        RECT 59.530 112.800 63.530 113.000 ;
        RECT 63.130 112.200 63.530 112.800 ;
        RECT 59.530 112.000 63.530 112.200 ;
        RECT 63.130 111.400 63.530 112.000 ;
        RECT 59.530 111.200 63.530 111.400 ;
        RECT 63.130 110.600 63.530 111.200 ;
        RECT 59.530 110.400 63.530 110.600 ;
        RECT 63.130 110.200 63.530 110.400 ;
        RECT 55.380 109.800 63.530 110.200 ;
        RECT 55.380 102.200 55.580 109.800 ;
        RECT 56.180 102.200 56.380 109.800 ;
        RECT 56.980 102.200 57.180 109.800 ;
        RECT 57.780 102.200 57.980 109.800 ;
        RECT 58.580 102.200 58.780 109.800 ;
        RECT 63.130 109.600 63.530 109.800 ;
        RECT 59.530 109.400 63.530 109.600 ;
        RECT 63.130 108.800 63.530 109.400 ;
        RECT 59.530 108.600 63.530 108.800 ;
        RECT 63.130 108.000 63.530 108.600 ;
        RECT 59.530 107.800 63.530 108.000 ;
        RECT 63.130 107.200 63.530 107.800 ;
        RECT 59.530 107.000 63.530 107.200 ;
        RECT 63.130 106.400 63.530 107.000 ;
        RECT 59.530 106.200 63.530 106.400 ;
        RECT 63.130 105.600 63.530 106.200 ;
        RECT 59.530 105.400 63.530 105.600 ;
        RECT 63.130 104.800 63.530 105.400 ;
        RECT 59.530 104.600 63.530 104.800 ;
        RECT 63.130 104.000 63.530 104.600 ;
        RECT 59.530 103.800 63.530 104.000 ;
        RECT 63.130 103.200 63.530 103.800 ;
        RECT 59.530 103.000 63.530 103.200 ;
        RECT 63.130 102.400 63.530 103.000 ;
        RECT 59.530 102.200 63.530 102.400 ;
        RECT 65.930 117.600 69.930 117.800 ;
        RECT 65.930 117.000 66.330 117.600 ;
        RECT 65.930 116.800 69.930 117.000 ;
        RECT 65.930 116.200 66.330 116.800 ;
        RECT 65.930 116.000 69.930 116.200 ;
        RECT 65.930 115.400 66.330 116.000 ;
        RECT 65.930 115.200 69.930 115.400 ;
        RECT 65.930 114.600 66.330 115.200 ;
        RECT 65.930 114.400 69.930 114.600 ;
        RECT 65.930 113.800 66.330 114.400 ;
        RECT 65.930 113.600 69.930 113.800 ;
        RECT 65.930 113.000 66.330 113.600 ;
        RECT 65.930 112.800 69.930 113.000 ;
        RECT 65.930 112.200 66.330 112.800 ;
        RECT 65.930 112.000 69.930 112.200 ;
        RECT 65.930 111.400 66.330 112.000 ;
        RECT 65.930 111.200 69.930 111.400 ;
        RECT 65.930 110.600 66.330 111.200 ;
        RECT 65.930 110.400 69.930 110.600 ;
        RECT 65.930 110.200 66.330 110.400 ;
        RECT 70.680 110.200 70.880 117.800 ;
        RECT 71.480 110.200 71.680 117.800 ;
        RECT 72.280 110.200 72.480 117.800 ;
        RECT 73.080 110.200 73.280 117.800 ;
        RECT 73.880 110.200 74.080 117.800 ;
        RECT 65.930 109.800 74.080 110.200 ;
        RECT 65.930 109.600 66.330 109.800 ;
        RECT 65.930 109.400 69.930 109.600 ;
        RECT 65.930 108.800 66.330 109.400 ;
        RECT 65.930 108.600 69.930 108.800 ;
        RECT 65.930 108.000 66.330 108.600 ;
        RECT 65.930 107.800 69.930 108.000 ;
        RECT 65.930 107.200 66.330 107.800 ;
        RECT 65.930 107.000 69.930 107.200 ;
        RECT 65.930 106.400 66.330 107.000 ;
        RECT 65.930 106.200 69.930 106.400 ;
        RECT 65.930 105.600 66.330 106.200 ;
        RECT 65.930 105.400 69.930 105.600 ;
        RECT 65.930 104.800 66.330 105.400 ;
        RECT 65.930 104.600 69.930 104.800 ;
        RECT 65.930 104.000 66.330 104.600 ;
        RECT 65.930 103.800 69.930 104.000 ;
        RECT 65.930 103.200 66.330 103.800 ;
        RECT 65.930 103.000 69.930 103.200 ;
        RECT 65.930 102.400 66.330 103.000 ;
        RECT 65.930 102.200 69.930 102.400 ;
        RECT 70.680 102.200 70.880 109.800 ;
        RECT 71.480 102.200 71.680 109.800 ;
        RECT 72.280 102.200 72.480 109.800 ;
        RECT 73.080 102.200 73.280 109.800 ;
        RECT 73.880 102.200 74.080 109.800 ;
        RECT 75.380 110.200 75.580 117.800 ;
        RECT 76.180 110.200 76.380 117.800 ;
        RECT 76.980 110.200 77.180 117.800 ;
        RECT 77.780 110.200 77.980 117.800 ;
        RECT 78.580 110.200 78.780 117.800 ;
        RECT 79.530 117.600 83.530 117.800 ;
        RECT 83.130 117.000 83.530 117.600 ;
        RECT 79.530 116.800 83.530 117.000 ;
        RECT 83.130 116.200 83.530 116.800 ;
        RECT 79.530 116.000 83.530 116.200 ;
        RECT 83.130 115.400 83.530 116.000 ;
        RECT 79.530 115.200 83.530 115.400 ;
        RECT 83.130 114.600 83.530 115.200 ;
        RECT 79.530 114.400 83.530 114.600 ;
        RECT 83.130 113.800 83.530 114.400 ;
        RECT 79.530 113.600 83.530 113.800 ;
        RECT 83.130 113.000 83.530 113.600 ;
        RECT 79.530 112.800 83.530 113.000 ;
        RECT 83.130 112.200 83.530 112.800 ;
        RECT 79.530 112.000 83.530 112.200 ;
        RECT 83.130 111.400 83.530 112.000 ;
        RECT 79.530 111.200 83.530 111.400 ;
        RECT 83.130 110.600 83.530 111.200 ;
        RECT 79.530 110.400 83.530 110.600 ;
        RECT 83.130 110.200 83.530 110.400 ;
        RECT 75.380 109.800 83.530 110.200 ;
        RECT 75.380 102.200 75.580 109.800 ;
        RECT 76.180 102.200 76.380 109.800 ;
        RECT 76.980 102.200 77.180 109.800 ;
        RECT 77.780 102.200 77.980 109.800 ;
        RECT 78.580 102.200 78.780 109.800 ;
        RECT 83.130 109.600 83.530 109.800 ;
        RECT 79.530 109.400 83.530 109.600 ;
        RECT 83.130 108.800 83.530 109.400 ;
        RECT 79.530 108.600 83.530 108.800 ;
        RECT 83.130 108.000 83.530 108.600 ;
        RECT 79.530 107.800 83.530 108.000 ;
        RECT 83.130 107.200 83.530 107.800 ;
        RECT 79.530 107.000 83.530 107.200 ;
        RECT 83.130 106.400 83.530 107.000 ;
        RECT 79.530 106.200 83.530 106.400 ;
        RECT 83.130 105.600 83.530 106.200 ;
        RECT 79.530 105.400 83.530 105.600 ;
        RECT 83.130 104.800 83.530 105.400 ;
        RECT 79.530 104.600 83.530 104.800 ;
        RECT 83.130 104.000 83.530 104.600 ;
        RECT 79.530 103.800 83.530 104.000 ;
        RECT 83.130 103.200 83.530 103.800 ;
        RECT 79.530 103.000 83.530 103.200 ;
        RECT 83.130 102.400 83.530 103.000 ;
        RECT 79.530 102.200 83.530 102.400 ;
        RECT 85.930 117.600 89.930 117.800 ;
        RECT 85.930 117.000 86.330 117.600 ;
        RECT 85.930 116.800 89.930 117.000 ;
        RECT 85.930 116.200 86.330 116.800 ;
        RECT 85.930 116.000 89.930 116.200 ;
        RECT 85.930 115.400 86.330 116.000 ;
        RECT 85.930 115.200 89.930 115.400 ;
        RECT 85.930 114.600 86.330 115.200 ;
        RECT 85.930 114.400 89.930 114.600 ;
        RECT 85.930 113.800 86.330 114.400 ;
        RECT 85.930 113.600 89.930 113.800 ;
        RECT 85.930 113.000 86.330 113.600 ;
        RECT 85.930 112.800 89.930 113.000 ;
        RECT 85.930 112.200 86.330 112.800 ;
        RECT 85.930 112.000 89.930 112.200 ;
        RECT 85.930 111.400 86.330 112.000 ;
        RECT 85.930 111.200 89.930 111.400 ;
        RECT 85.930 110.600 86.330 111.200 ;
        RECT 85.930 110.400 89.930 110.600 ;
        RECT 85.930 110.200 86.330 110.400 ;
        RECT 90.680 110.200 90.880 117.800 ;
        RECT 91.480 110.200 91.680 117.800 ;
        RECT 92.280 110.200 92.480 117.800 ;
        RECT 93.080 110.200 93.280 117.800 ;
        RECT 93.880 110.200 94.080 117.800 ;
        RECT 85.930 109.800 94.080 110.200 ;
        RECT 85.930 109.600 86.330 109.800 ;
        RECT 85.930 109.400 89.930 109.600 ;
        RECT 85.930 108.800 86.330 109.400 ;
        RECT 85.930 108.600 89.930 108.800 ;
        RECT 85.930 108.000 86.330 108.600 ;
        RECT 85.930 107.800 89.930 108.000 ;
        RECT 85.930 107.200 86.330 107.800 ;
        RECT 85.930 107.000 89.930 107.200 ;
        RECT 85.930 106.400 86.330 107.000 ;
        RECT 85.930 106.200 89.930 106.400 ;
        RECT 85.930 105.600 86.330 106.200 ;
        RECT 85.930 105.400 89.930 105.600 ;
        RECT 85.930 104.800 86.330 105.400 ;
        RECT 85.930 104.600 89.930 104.800 ;
        RECT 85.930 104.000 86.330 104.600 ;
        RECT 85.930 103.800 89.930 104.000 ;
        RECT 85.930 103.200 86.330 103.800 ;
        RECT 85.930 103.000 89.930 103.200 ;
        RECT 85.930 102.400 86.330 103.000 ;
        RECT 85.930 102.200 89.930 102.400 ;
        RECT 90.680 102.200 90.880 109.800 ;
        RECT 91.480 102.200 91.680 109.800 ;
        RECT 92.280 102.200 92.480 109.800 ;
        RECT 93.080 102.200 93.280 109.800 ;
        RECT 93.880 102.200 94.080 109.800 ;
        RECT 95.380 110.200 95.580 117.800 ;
        RECT 96.180 110.200 96.380 117.800 ;
        RECT 96.980 110.200 97.180 117.800 ;
        RECT 97.780 110.200 97.980 117.800 ;
        RECT 98.580 110.200 98.780 117.800 ;
        RECT 99.530 117.600 103.530 117.800 ;
        RECT 103.130 117.000 103.530 117.600 ;
        RECT 99.530 116.800 103.530 117.000 ;
        RECT 103.130 116.200 103.530 116.800 ;
        RECT 99.530 116.000 103.530 116.200 ;
        RECT 103.130 115.400 103.530 116.000 ;
        RECT 99.530 115.200 103.530 115.400 ;
        RECT 103.130 114.600 103.530 115.200 ;
        RECT 99.530 114.400 103.530 114.600 ;
        RECT 103.130 113.800 103.530 114.400 ;
        RECT 99.530 113.600 103.530 113.800 ;
        RECT 103.130 113.000 103.530 113.600 ;
        RECT 99.530 112.800 103.530 113.000 ;
        RECT 103.130 112.200 103.530 112.800 ;
        RECT 99.530 112.000 103.530 112.200 ;
        RECT 103.130 111.400 103.530 112.000 ;
        RECT 99.530 111.200 103.530 111.400 ;
        RECT 103.130 110.600 103.530 111.200 ;
        RECT 99.530 110.400 103.530 110.600 ;
        RECT 110.050 110.525 110.410 110.905 ;
        RECT 110.680 110.525 111.040 110.905 ;
        RECT 111.280 110.525 111.640 110.905 ;
        RECT 103.130 110.200 103.530 110.400 ;
        RECT 95.380 109.800 103.530 110.200 ;
        RECT 110.050 109.935 110.410 110.315 ;
        RECT 110.680 109.935 111.040 110.315 ;
        RECT 111.280 109.935 111.640 110.315 ;
        RECT 95.380 102.200 95.580 109.800 ;
        RECT 96.180 102.200 96.380 109.800 ;
        RECT 96.980 102.200 97.180 109.800 ;
        RECT 97.780 102.200 97.980 109.800 ;
        RECT 98.580 102.200 98.780 109.800 ;
        RECT 103.130 109.600 103.530 109.800 ;
        RECT 99.530 109.400 103.530 109.600 ;
        RECT 103.130 108.800 103.530 109.400 ;
        RECT 99.530 108.600 103.530 108.800 ;
        RECT 103.130 108.000 103.530 108.600 ;
        RECT 99.530 107.800 103.530 108.000 ;
        RECT 103.130 107.200 103.530 107.800 ;
        RECT 99.530 107.000 103.530 107.200 ;
        RECT 103.130 106.400 103.530 107.000 ;
        RECT 99.530 106.200 103.530 106.400 ;
        RECT 103.130 105.600 103.530 106.200 ;
        RECT 99.530 105.400 103.530 105.600 ;
        RECT 103.130 104.800 103.530 105.400 ;
        RECT 99.530 104.600 103.530 104.800 ;
        RECT 103.130 104.000 103.530 104.600 ;
        RECT 99.530 103.800 103.530 104.000 ;
        RECT 103.130 103.200 103.530 103.800 ;
        RECT 99.530 103.000 103.530 103.200 ;
        RECT 103.130 102.400 103.530 103.000 ;
        RECT 99.530 102.200 103.530 102.400 ;
        RECT 5.930 97.600 9.930 97.800 ;
        RECT 5.930 97.000 6.330 97.600 ;
        RECT 5.930 96.800 9.930 97.000 ;
        RECT 5.930 96.200 6.330 96.800 ;
        RECT 5.930 96.000 9.930 96.200 ;
        RECT 5.930 95.400 6.330 96.000 ;
        RECT 5.930 95.200 9.930 95.400 ;
        RECT 5.930 94.600 6.330 95.200 ;
        RECT 5.930 94.400 9.930 94.600 ;
        RECT 5.930 93.800 6.330 94.400 ;
        RECT 5.930 93.600 9.930 93.800 ;
        RECT 5.930 93.000 6.330 93.600 ;
        RECT 5.930 92.800 9.930 93.000 ;
        RECT 5.930 92.200 6.330 92.800 ;
        RECT 5.930 92.000 9.930 92.200 ;
        RECT 5.930 91.400 6.330 92.000 ;
        RECT 5.930 91.200 9.930 91.400 ;
        RECT 5.930 90.600 6.330 91.200 ;
        RECT 5.930 90.400 9.930 90.600 ;
        RECT 5.930 90.200 6.330 90.400 ;
        RECT 10.680 90.200 10.880 97.800 ;
        RECT 11.480 90.200 11.680 97.800 ;
        RECT 12.280 90.200 12.480 97.800 ;
        RECT 13.080 90.200 13.280 97.800 ;
        RECT 13.880 90.200 14.080 97.800 ;
        RECT 5.930 89.800 14.080 90.200 ;
        RECT 5.930 89.600 6.330 89.800 ;
        RECT 5.930 89.400 9.930 89.600 ;
        RECT 5.930 88.800 6.330 89.400 ;
        RECT 5.930 88.600 9.930 88.800 ;
        RECT 5.930 88.000 6.330 88.600 ;
        RECT 5.930 87.800 9.930 88.000 ;
        RECT 5.930 87.200 6.330 87.800 ;
        RECT 5.930 87.000 9.930 87.200 ;
        RECT 5.930 86.400 6.330 87.000 ;
        RECT 5.930 86.200 9.930 86.400 ;
        RECT 5.930 85.600 6.330 86.200 ;
        RECT 5.930 85.400 9.930 85.600 ;
        RECT 5.930 84.800 6.330 85.400 ;
        RECT 5.930 84.600 9.930 84.800 ;
        RECT 5.930 84.000 6.330 84.600 ;
        RECT 5.930 83.800 9.930 84.000 ;
        RECT 5.930 83.200 6.330 83.800 ;
        RECT 5.930 83.000 9.930 83.200 ;
        RECT 5.930 82.400 6.330 83.000 ;
        RECT 5.930 82.200 9.930 82.400 ;
        RECT 10.680 82.200 10.880 89.800 ;
        RECT 11.480 82.200 11.680 89.800 ;
        RECT 12.280 82.200 12.480 89.800 ;
        RECT 13.080 82.200 13.280 89.800 ;
        RECT 13.880 82.200 14.080 89.800 ;
        RECT 15.380 90.200 15.580 97.800 ;
        RECT 16.180 90.200 16.380 97.800 ;
        RECT 16.980 90.200 17.180 97.800 ;
        RECT 17.780 90.200 17.980 97.800 ;
        RECT 18.580 90.200 18.780 97.800 ;
        RECT 19.530 97.600 23.530 97.800 ;
        RECT 23.130 97.000 23.530 97.600 ;
        RECT 19.530 96.800 23.530 97.000 ;
        RECT 23.130 96.200 23.530 96.800 ;
        RECT 19.530 96.000 23.530 96.200 ;
        RECT 23.130 95.400 23.530 96.000 ;
        RECT 19.530 95.200 23.530 95.400 ;
        RECT 23.130 94.600 23.530 95.200 ;
        RECT 19.530 94.400 23.530 94.600 ;
        RECT 23.130 93.800 23.530 94.400 ;
        RECT 19.530 93.600 23.530 93.800 ;
        RECT 23.130 93.000 23.530 93.600 ;
        RECT 19.530 92.800 23.530 93.000 ;
        RECT 23.130 92.200 23.530 92.800 ;
        RECT 19.530 92.000 23.530 92.200 ;
        RECT 23.130 91.400 23.530 92.000 ;
        RECT 19.530 91.200 23.530 91.400 ;
        RECT 23.130 90.600 23.530 91.200 ;
        RECT 19.530 90.400 23.530 90.600 ;
        RECT 23.130 90.200 23.530 90.400 ;
        RECT 15.380 89.800 23.530 90.200 ;
        RECT 15.380 82.200 15.580 89.800 ;
        RECT 16.180 82.200 16.380 89.800 ;
        RECT 16.980 82.200 17.180 89.800 ;
        RECT 17.780 82.200 17.980 89.800 ;
        RECT 18.580 82.200 18.780 89.800 ;
        RECT 23.130 89.600 23.530 89.800 ;
        RECT 19.530 89.400 23.530 89.600 ;
        RECT 23.130 88.800 23.530 89.400 ;
        RECT 19.530 88.600 23.530 88.800 ;
        RECT 23.130 88.000 23.530 88.600 ;
        RECT 19.530 87.800 23.530 88.000 ;
        RECT 23.130 87.200 23.530 87.800 ;
        RECT 19.530 87.000 23.530 87.200 ;
        RECT 23.130 86.400 23.530 87.000 ;
        RECT 19.530 86.200 23.530 86.400 ;
        RECT 23.130 85.600 23.530 86.200 ;
        RECT 19.530 85.400 23.530 85.600 ;
        RECT 23.130 84.800 23.530 85.400 ;
        RECT 19.530 84.600 23.530 84.800 ;
        RECT 23.130 84.000 23.530 84.600 ;
        RECT 19.530 83.800 23.530 84.000 ;
        RECT 23.130 83.200 23.530 83.800 ;
        RECT 19.530 83.000 23.530 83.200 ;
        RECT 23.130 82.400 23.530 83.000 ;
        RECT 19.530 82.200 23.530 82.400 ;
        RECT 25.930 97.600 29.930 97.800 ;
        RECT 25.930 97.000 26.330 97.600 ;
        RECT 25.930 96.800 29.930 97.000 ;
        RECT 25.930 96.200 26.330 96.800 ;
        RECT 25.930 96.000 29.930 96.200 ;
        RECT 25.930 95.400 26.330 96.000 ;
        RECT 25.930 95.200 29.930 95.400 ;
        RECT 25.930 94.600 26.330 95.200 ;
        RECT 25.930 94.400 29.930 94.600 ;
        RECT 25.930 93.800 26.330 94.400 ;
        RECT 25.930 93.600 29.930 93.800 ;
        RECT 25.930 93.000 26.330 93.600 ;
        RECT 25.930 92.800 29.930 93.000 ;
        RECT 25.930 92.200 26.330 92.800 ;
        RECT 25.930 92.000 29.930 92.200 ;
        RECT 25.930 91.400 26.330 92.000 ;
        RECT 25.930 91.200 29.930 91.400 ;
        RECT 25.930 90.600 26.330 91.200 ;
        RECT 25.930 90.400 29.930 90.600 ;
        RECT 25.930 90.200 26.330 90.400 ;
        RECT 30.680 90.200 30.880 97.800 ;
        RECT 31.480 90.200 31.680 97.800 ;
        RECT 32.280 90.200 32.480 97.800 ;
        RECT 33.080 90.200 33.280 97.800 ;
        RECT 33.880 90.200 34.080 97.800 ;
        RECT 25.930 89.800 34.080 90.200 ;
        RECT 25.930 89.600 26.330 89.800 ;
        RECT 25.930 89.400 29.930 89.600 ;
        RECT 25.930 88.800 26.330 89.400 ;
        RECT 25.930 88.600 29.930 88.800 ;
        RECT 25.930 88.000 26.330 88.600 ;
        RECT 25.930 87.800 29.930 88.000 ;
        RECT 25.930 87.200 26.330 87.800 ;
        RECT 25.930 87.000 29.930 87.200 ;
        RECT 25.930 86.400 26.330 87.000 ;
        RECT 25.930 86.200 29.930 86.400 ;
        RECT 25.930 85.600 26.330 86.200 ;
        RECT 25.930 85.400 29.930 85.600 ;
        RECT 25.930 84.800 26.330 85.400 ;
        RECT 25.930 84.600 29.930 84.800 ;
        RECT 25.930 84.000 26.330 84.600 ;
        RECT 25.930 83.800 29.930 84.000 ;
        RECT 25.930 83.200 26.330 83.800 ;
        RECT 25.930 83.000 29.930 83.200 ;
        RECT 25.930 82.400 26.330 83.000 ;
        RECT 25.930 82.200 29.930 82.400 ;
        RECT 30.680 82.200 30.880 89.800 ;
        RECT 31.480 82.200 31.680 89.800 ;
        RECT 32.280 82.200 32.480 89.800 ;
        RECT 33.080 82.200 33.280 89.800 ;
        RECT 33.880 82.200 34.080 89.800 ;
        RECT 35.380 90.200 35.580 97.800 ;
        RECT 36.180 90.200 36.380 97.800 ;
        RECT 36.980 90.200 37.180 97.800 ;
        RECT 37.780 90.200 37.980 97.800 ;
        RECT 38.580 90.200 38.780 97.800 ;
        RECT 39.530 97.600 43.530 97.800 ;
        RECT 43.130 97.000 43.530 97.600 ;
        RECT 39.530 96.800 43.530 97.000 ;
        RECT 43.130 96.200 43.530 96.800 ;
        RECT 39.530 96.000 43.530 96.200 ;
        RECT 43.130 95.400 43.530 96.000 ;
        RECT 39.530 95.200 43.530 95.400 ;
        RECT 43.130 94.600 43.530 95.200 ;
        RECT 39.530 94.400 43.530 94.600 ;
        RECT 43.130 93.800 43.530 94.400 ;
        RECT 39.530 93.600 43.530 93.800 ;
        RECT 43.130 93.000 43.530 93.600 ;
        RECT 39.530 92.800 43.530 93.000 ;
        RECT 43.130 92.200 43.530 92.800 ;
        RECT 39.530 92.000 43.530 92.200 ;
        RECT 43.130 91.400 43.530 92.000 ;
        RECT 39.530 91.200 43.530 91.400 ;
        RECT 43.130 90.600 43.530 91.200 ;
        RECT 39.530 90.400 43.530 90.600 ;
        RECT 43.130 90.200 43.530 90.400 ;
        RECT 35.380 89.800 43.530 90.200 ;
        RECT 35.380 82.200 35.580 89.800 ;
        RECT 36.180 82.200 36.380 89.800 ;
        RECT 36.980 82.200 37.180 89.800 ;
        RECT 37.780 82.200 37.980 89.800 ;
        RECT 38.580 82.200 38.780 89.800 ;
        RECT 43.130 89.600 43.530 89.800 ;
        RECT 39.530 89.400 43.530 89.600 ;
        RECT 43.130 88.800 43.530 89.400 ;
        RECT 39.530 88.600 43.530 88.800 ;
        RECT 43.130 88.000 43.530 88.600 ;
        RECT 39.530 87.800 43.530 88.000 ;
        RECT 43.130 87.200 43.530 87.800 ;
        RECT 39.530 87.000 43.530 87.200 ;
        RECT 43.130 86.400 43.530 87.000 ;
        RECT 39.530 86.200 43.530 86.400 ;
        RECT 43.130 85.600 43.530 86.200 ;
        RECT 39.530 85.400 43.530 85.600 ;
        RECT 43.130 84.800 43.530 85.400 ;
        RECT 39.530 84.600 43.530 84.800 ;
        RECT 43.130 84.000 43.530 84.600 ;
        RECT 39.530 83.800 43.530 84.000 ;
        RECT 43.130 83.200 43.530 83.800 ;
        RECT 39.530 83.000 43.530 83.200 ;
        RECT 43.130 82.400 43.530 83.000 ;
        RECT 39.530 82.200 43.530 82.400 ;
        RECT 45.930 97.600 49.930 97.800 ;
        RECT 45.930 97.000 46.330 97.600 ;
        RECT 45.930 96.800 49.930 97.000 ;
        RECT 45.930 96.200 46.330 96.800 ;
        RECT 45.930 96.000 49.930 96.200 ;
        RECT 45.930 95.400 46.330 96.000 ;
        RECT 45.930 95.200 49.930 95.400 ;
        RECT 45.930 94.600 46.330 95.200 ;
        RECT 45.930 94.400 49.930 94.600 ;
        RECT 45.930 93.800 46.330 94.400 ;
        RECT 45.930 93.600 49.930 93.800 ;
        RECT 45.930 93.000 46.330 93.600 ;
        RECT 45.930 92.800 49.930 93.000 ;
        RECT 45.930 92.200 46.330 92.800 ;
        RECT 45.930 92.000 49.930 92.200 ;
        RECT 45.930 91.400 46.330 92.000 ;
        RECT 45.930 91.200 49.930 91.400 ;
        RECT 45.930 90.600 46.330 91.200 ;
        RECT 45.930 90.400 49.930 90.600 ;
        RECT 45.930 90.200 46.330 90.400 ;
        RECT 50.680 90.200 50.880 97.800 ;
        RECT 51.480 90.200 51.680 97.800 ;
        RECT 52.280 90.200 52.480 97.800 ;
        RECT 53.080 90.200 53.280 97.800 ;
        RECT 53.880 90.200 54.080 97.800 ;
        RECT 45.930 89.800 54.080 90.200 ;
        RECT 45.930 89.600 46.330 89.800 ;
        RECT 45.930 89.400 49.930 89.600 ;
        RECT 45.930 88.800 46.330 89.400 ;
        RECT 45.930 88.600 49.930 88.800 ;
        RECT 45.930 88.000 46.330 88.600 ;
        RECT 45.930 87.800 49.930 88.000 ;
        RECT 45.930 87.200 46.330 87.800 ;
        RECT 45.930 87.000 49.930 87.200 ;
        RECT 45.930 86.400 46.330 87.000 ;
        RECT 45.930 86.200 49.930 86.400 ;
        RECT 45.930 85.600 46.330 86.200 ;
        RECT 45.930 85.400 49.930 85.600 ;
        RECT 45.930 84.800 46.330 85.400 ;
        RECT 45.930 84.600 49.930 84.800 ;
        RECT 45.930 84.000 46.330 84.600 ;
        RECT 45.930 83.800 49.930 84.000 ;
        RECT 45.930 83.200 46.330 83.800 ;
        RECT 45.930 83.000 49.930 83.200 ;
        RECT 45.930 82.400 46.330 83.000 ;
        RECT 45.930 82.200 49.930 82.400 ;
        RECT 50.680 82.200 50.880 89.800 ;
        RECT 51.480 82.200 51.680 89.800 ;
        RECT 52.280 82.200 52.480 89.800 ;
        RECT 53.080 82.200 53.280 89.800 ;
        RECT 53.880 82.200 54.080 89.800 ;
        RECT 55.380 90.200 55.580 97.800 ;
        RECT 56.180 90.200 56.380 97.800 ;
        RECT 56.980 90.200 57.180 97.800 ;
        RECT 57.780 90.200 57.980 97.800 ;
        RECT 58.580 90.200 58.780 97.800 ;
        RECT 59.530 97.600 63.530 97.800 ;
        RECT 63.130 97.000 63.530 97.600 ;
        RECT 59.530 96.800 63.530 97.000 ;
        RECT 63.130 96.200 63.530 96.800 ;
        RECT 59.530 96.000 63.530 96.200 ;
        RECT 63.130 95.400 63.530 96.000 ;
        RECT 59.530 95.200 63.530 95.400 ;
        RECT 63.130 94.600 63.530 95.200 ;
        RECT 59.530 94.400 63.530 94.600 ;
        RECT 63.130 93.800 63.530 94.400 ;
        RECT 59.530 93.600 63.530 93.800 ;
        RECT 63.130 93.000 63.530 93.600 ;
        RECT 59.530 92.800 63.530 93.000 ;
        RECT 63.130 92.200 63.530 92.800 ;
        RECT 59.530 92.000 63.530 92.200 ;
        RECT 63.130 91.400 63.530 92.000 ;
        RECT 59.530 91.200 63.530 91.400 ;
        RECT 63.130 90.600 63.530 91.200 ;
        RECT 59.530 90.400 63.530 90.600 ;
        RECT 63.130 90.200 63.530 90.400 ;
        RECT 55.380 89.800 63.530 90.200 ;
        RECT 55.380 82.200 55.580 89.800 ;
        RECT 56.180 82.200 56.380 89.800 ;
        RECT 56.980 82.200 57.180 89.800 ;
        RECT 57.780 82.200 57.980 89.800 ;
        RECT 58.580 82.200 58.780 89.800 ;
        RECT 63.130 89.600 63.530 89.800 ;
        RECT 59.530 89.400 63.530 89.600 ;
        RECT 63.130 88.800 63.530 89.400 ;
        RECT 59.530 88.600 63.530 88.800 ;
        RECT 63.130 88.000 63.530 88.600 ;
        RECT 59.530 87.800 63.530 88.000 ;
        RECT 63.130 87.200 63.530 87.800 ;
        RECT 59.530 87.000 63.530 87.200 ;
        RECT 63.130 86.400 63.530 87.000 ;
        RECT 59.530 86.200 63.530 86.400 ;
        RECT 63.130 85.600 63.530 86.200 ;
        RECT 59.530 85.400 63.530 85.600 ;
        RECT 63.130 84.800 63.530 85.400 ;
        RECT 59.530 84.600 63.530 84.800 ;
        RECT 63.130 84.000 63.530 84.600 ;
        RECT 59.530 83.800 63.530 84.000 ;
        RECT 63.130 83.200 63.530 83.800 ;
        RECT 59.530 83.000 63.530 83.200 ;
        RECT 63.130 82.400 63.530 83.000 ;
        RECT 59.530 82.200 63.530 82.400 ;
        RECT 65.930 97.600 69.930 97.800 ;
        RECT 65.930 97.000 66.330 97.600 ;
        RECT 65.930 96.800 69.930 97.000 ;
        RECT 65.930 96.200 66.330 96.800 ;
        RECT 65.930 96.000 69.930 96.200 ;
        RECT 65.930 95.400 66.330 96.000 ;
        RECT 65.930 95.200 69.930 95.400 ;
        RECT 65.930 94.600 66.330 95.200 ;
        RECT 65.930 94.400 69.930 94.600 ;
        RECT 65.930 93.800 66.330 94.400 ;
        RECT 65.930 93.600 69.930 93.800 ;
        RECT 65.930 93.000 66.330 93.600 ;
        RECT 65.930 92.800 69.930 93.000 ;
        RECT 65.930 92.200 66.330 92.800 ;
        RECT 65.930 92.000 69.930 92.200 ;
        RECT 65.930 91.400 66.330 92.000 ;
        RECT 65.930 91.200 69.930 91.400 ;
        RECT 65.930 90.600 66.330 91.200 ;
        RECT 65.930 90.400 69.930 90.600 ;
        RECT 65.930 90.200 66.330 90.400 ;
        RECT 70.680 90.200 70.880 97.800 ;
        RECT 71.480 90.200 71.680 97.800 ;
        RECT 72.280 90.200 72.480 97.800 ;
        RECT 73.080 90.200 73.280 97.800 ;
        RECT 73.880 90.200 74.080 97.800 ;
        RECT 65.930 89.800 74.080 90.200 ;
        RECT 65.930 89.600 66.330 89.800 ;
        RECT 65.930 89.400 69.930 89.600 ;
        RECT 65.930 88.800 66.330 89.400 ;
        RECT 65.930 88.600 69.930 88.800 ;
        RECT 65.930 88.000 66.330 88.600 ;
        RECT 65.930 87.800 69.930 88.000 ;
        RECT 65.930 87.200 66.330 87.800 ;
        RECT 65.930 87.000 69.930 87.200 ;
        RECT 65.930 86.400 66.330 87.000 ;
        RECT 65.930 86.200 69.930 86.400 ;
        RECT 65.930 85.600 66.330 86.200 ;
        RECT 65.930 85.400 69.930 85.600 ;
        RECT 65.930 84.800 66.330 85.400 ;
        RECT 65.930 84.600 69.930 84.800 ;
        RECT 65.930 84.000 66.330 84.600 ;
        RECT 65.930 83.800 69.930 84.000 ;
        RECT 65.930 83.200 66.330 83.800 ;
        RECT 65.930 83.000 69.930 83.200 ;
        RECT 65.930 82.400 66.330 83.000 ;
        RECT 65.930 82.200 69.930 82.400 ;
        RECT 70.680 82.200 70.880 89.800 ;
        RECT 71.480 82.200 71.680 89.800 ;
        RECT 72.280 82.200 72.480 89.800 ;
        RECT 73.080 82.200 73.280 89.800 ;
        RECT 73.880 82.200 74.080 89.800 ;
        RECT 75.380 90.200 75.580 97.800 ;
        RECT 76.180 90.200 76.380 97.800 ;
        RECT 76.980 90.200 77.180 97.800 ;
        RECT 77.780 90.200 77.980 97.800 ;
        RECT 78.580 90.200 78.780 97.800 ;
        RECT 79.530 97.600 83.530 97.800 ;
        RECT 83.130 97.000 83.530 97.600 ;
        RECT 79.530 96.800 83.530 97.000 ;
        RECT 83.130 96.200 83.530 96.800 ;
        RECT 79.530 96.000 83.530 96.200 ;
        RECT 83.130 95.400 83.530 96.000 ;
        RECT 79.530 95.200 83.530 95.400 ;
        RECT 83.130 94.600 83.530 95.200 ;
        RECT 79.530 94.400 83.530 94.600 ;
        RECT 83.130 93.800 83.530 94.400 ;
        RECT 79.530 93.600 83.530 93.800 ;
        RECT 83.130 93.000 83.530 93.600 ;
        RECT 79.530 92.800 83.530 93.000 ;
        RECT 83.130 92.200 83.530 92.800 ;
        RECT 79.530 92.000 83.530 92.200 ;
        RECT 83.130 91.400 83.530 92.000 ;
        RECT 79.530 91.200 83.530 91.400 ;
        RECT 83.130 90.600 83.530 91.200 ;
        RECT 79.530 90.400 83.530 90.600 ;
        RECT 83.130 90.200 83.530 90.400 ;
        RECT 75.380 89.800 83.530 90.200 ;
        RECT 75.380 82.200 75.580 89.800 ;
        RECT 76.180 82.200 76.380 89.800 ;
        RECT 76.980 82.200 77.180 89.800 ;
        RECT 77.780 82.200 77.980 89.800 ;
        RECT 78.580 82.200 78.780 89.800 ;
        RECT 83.130 89.600 83.530 89.800 ;
        RECT 79.530 89.400 83.530 89.600 ;
        RECT 83.130 88.800 83.530 89.400 ;
        RECT 79.530 88.600 83.530 88.800 ;
        RECT 83.130 88.000 83.530 88.600 ;
        RECT 79.530 87.800 83.530 88.000 ;
        RECT 83.130 87.200 83.530 87.800 ;
        RECT 79.530 87.000 83.530 87.200 ;
        RECT 83.130 86.400 83.530 87.000 ;
        RECT 79.530 86.200 83.530 86.400 ;
        RECT 83.130 85.600 83.530 86.200 ;
        RECT 79.530 85.400 83.530 85.600 ;
        RECT 83.130 84.800 83.530 85.400 ;
        RECT 79.530 84.600 83.530 84.800 ;
        RECT 83.130 84.000 83.530 84.600 ;
        RECT 79.530 83.800 83.530 84.000 ;
        RECT 83.130 83.200 83.530 83.800 ;
        RECT 79.530 83.000 83.530 83.200 ;
        RECT 83.130 82.400 83.530 83.000 ;
        RECT 79.530 82.200 83.530 82.400 ;
        RECT 85.930 97.600 89.930 97.800 ;
        RECT 85.930 97.000 86.330 97.600 ;
        RECT 85.930 96.800 89.930 97.000 ;
        RECT 85.930 96.200 86.330 96.800 ;
        RECT 85.930 96.000 89.930 96.200 ;
        RECT 85.930 95.400 86.330 96.000 ;
        RECT 85.930 95.200 89.930 95.400 ;
        RECT 85.930 94.600 86.330 95.200 ;
        RECT 85.930 94.400 89.930 94.600 ;
        RECT 85.930 93.800 86.330 94.400 ;
        RECT 85.930 93.600 89.930 93.800 ;
        RECT 85.930 93.000 86.330 93.600 ;
        RECT 85.930 92.800 89.930 93.000 ;
        RECT 85.930 92.200 86.330 92.800 ;
        RECT 85.930 92.000 89.930 92.200 ;
        RECT 85.930 91.400 86.330 92.000 ;
        RECT 85.930 91.200 89.930 91.400 ;
        RECT 85.930 90.600 86.330 91.200 ;
        RECT 85.930 90.400 89.930 90.600 ;
        RECT 85.930 90.200 86.330 90.400 ;
        RECT 90.680 90.200 90.880 97.800 ;
        RECT 91.480 90.200 91.680 97.800 ;
        RECT 92.280 90.200 92.480 97.800 ;
        RECT 93.080 90.200 93.280 97.800 ;
        RECT 93.880 90.200 94.080 97.800 ;
        RECT 85.930 89.800 94.080 90.200 ;
        RECT 85.930 89.600 86.330 89.800 ;
        RECT 85.930 89.400 89.930 89.600 ;
        RECT 85.930 88.800 86.330 89.400 ;
        RECT 85.930 88.600 89.930 88.800 ;
        RECT 85.930 88.000 86.330 88.600 ;
        RECT 85.930 87.800 89.930 88.000 ;
        RECT 85.930 87.200 86.330 87.800 ;
        RECT 85.930 87.000 89.930 87.200 ;
        RECT 85.930 86.400 86.330 87.000 ;
        RECT 85.930 86.200 89.930 86.400 ;
        RECT 85.930 85.600 86.330 86.200 ;
        RECT 85.930 85.400 89.930 85.600 ;
        RECT 85.930 84.800 86.330 85.400 ;
        RECT 85.930 84.600 89.930 84.800 ;
        RECT 85.930 84.000 86.330 84.600 ;
        RECT 85.930 83.800 89.930 84.000 ;
        RECT 85.930 83.200 86.330 83.800 ;
        RECT 85.930 83.000 89.930 83.200 ;
        RECT 85.930 82.400 86.330 83.000 ;
        RECT 85.930 82.200 89.930 82.400 ;
        RECT 90.680 82.200 90.880 89.800 ;
        RECT 91.480 82.200 91.680 89.800 ;
        RECT 92.280 82.200 92.480 89.800 ;
        RECT 93.080 82.200 93.280 89.800 ;
        RECT 93.880 82.200 94.080 89.800 ;
        RECT 95.380 90.200 95.580 97.800 ;
        RECT 96.180 90.200 96.380 97.800 ;
        RECT 96.980 90.200 97.180 97.800 ;
        RECT 97.780 90.200 97.980 97.800 ;
        RECT 98.580 90.200 98.780 97.800 ;
        RECT 99.530 97.600 103.530 97.800 ;
        RECT 103.130 97.000 103.530 97.600 ;
        RECT 99.530 96.800 103.530 97.000 ;
        RECT 103.130 96.200 103.530 96.800 ;
        RECT 99.530 96.000 103.530 96.200 ;
        RECT 103.130 95.400 103.530 96.000 ;
        RECT 99.530 95.200 103.530 95.400 ;
        RECT 103.130 94.600 103.530 95.200 ;
        RECT 99.530 94.400 103.530 94.600 ;
        RECT 103.130 93.800 103.530 94.400 ;
        RECT 99.530 93.600 103.530 93.800 ;
        RECT 103.130 93.000 103.530 93.600 ;
        RECT 99.530 92.800 103.530 93.000 ;
        RECT 103.130 92.200 103.530 92.800 ;
        RECT 99.530 92.000 103.530 92.200 ;
        RECT 103.130 91.400 103.530 92.000 ;
        RECT 99.530 91.200 103.530 91.400 ;
        RECT 103.130 90.600 103.530 91.200 ;
        RECT 99.530 90.400 103.530 90.600 ;
        RECT 103.130 90.200 103.530 90.400 ;
        RECT 95.380 89.800 103.530 90.200 ;
        RECT 110.050 89.990 110.410 90.370 ;
        RECT 110.680 89.990 111.040 90.370 ;
        RECT 111.280 89.990 111.640 90.370 ;
        RECT 95.380 82.200 95.580 89.800 ;
        RECT 96.180 82.200 96.380 89.800 ;
        RECT 96.980 82.200 97.180 89.800 ;
        RECT 97.780 82.200 97.980 89.800 ;
        RECT 98.580 82.200 98.780 89.800 ;
        RECT 103.130 89.600 103.530 89.800 ;
        RECT 99.530 89.400 103.530 89.600 ;
        RECT 110.050 89.400 110.410 89.780 ;
        RECT 110.680 89.400 111.040 89.780 ;
        RECT 111.280 89.400 111.640 89.780 ;
        RECT 103.130 88.800 103.530 89.400 ;
        RECT 99.530 88.600 103.530 88.800 ;
        RECT 103.130 88.000 103.530 88.600 ;
        RECT 99.530 87.800 103.530 88.000 ;
        RECT 103.130 87.200 103.530 87.800 ;
        RECT 99.530 87.000 103.530 87.200 ;
        RECT 103.130 86.400 103.530 87.000 ;
        RECT 99.530 86.200 103.530 86.400 ;
        RECT 103.130 85.600 103.530 86.200 ;
        RECT 99.530 85.400 103.530 85.600 ;
        RECT 103.130 84.800 103.530 85.400 ;
        RECT 99.530 84.600 103.530 84.800 ;
        RECT 103.130 84.000 103.530 84.600 ;
        RECT 99.530 83.800 103.530 84.000 ;
        RECT 103.130 83.200 103.530 83.800 ;
        RECT 99.530 83.000 103.530 83.200 ;
        RECT 103.130 82.400 103.530 83.000 ;
        RECT 99.530 82.200 103.530 82.400 ;
        RECT 5.930 77.600 9.930 77.800 ;
        RECT 5.930 77.000 6.330 77.600 ;
        RECT 5.930 76.800 9.930 77.000 ;
        RECT 5.930 76.200 6.330 76.800 ;
        RECT 5.930 76.000 9.930 76.200 ;
        RECT 5.930 75.400 6.330 76.000 ;
        RECT 5.930 75.200 9.930 75.400 ;
        RECT 5.930 74.600 6.330 75.200 ;
        RECT 5.930 74.400 9.930 74.600 ;
        RECT 5.930 73.800 6.330 74.400 ;
        RECT 5.930 73.600 9.930 73.800 ;
        RECT 5.930 73.000 6.330 73.600 ;
        RECT 5.930 72.800 9.930 73.000 ;
        RECT 5.930 72.200 6.330 72.800 ;
        RECT 5.930 72.000 9.930 72.200 ;
        RECT 5.930 71.400 6.330 72.000 ;
        RECT 5.930 71.200 9.930 71.400 ;
        RECT 5.930 70.600 6.330 71.200 ;
        RECT 5.930 70.400 9.930 70.600 ;
        RECT 5.930 70.200 6.330 70.400 ;
        RECT 10.680 70.200 10.880 77.800 ;
        RECT 11.480 70.200 11.680 77.800 ;
        RECT 12.280 70.200 12.480 77.800 ;
        RECT 13.080 70.200 13.280 77.800 ;
        RECT 13.880 70.200 14.080 77.800 ;
        RECT 5.930 69.800 14.080 70.200 ;
        RECT 5.930 69.600 6.330 69.800 ;
        RECT 5.930 69.400 9.930 69.600 ;
        RECT 5.930 68.800 6.330 69.400 ;
        RECT 5.930 68.600 9.930 68.800 ;
        RECT 5.930 68.000 6.330 68.600 ;
        RECT 5.930 67.800 9.930 68.000 ;
        RECT 5.930 67.200 6.330 67.800 ;
        RECT 5.930 67.000 9.930 67.200 ;
        RECT 5.930 66.400 6.330 67.000 ;
        RECT 5.930 66.200 9.930 66.400 ;
        RECT 5.930 65.600 6.330 66.200 ;
        RECT 5.930 65.400 9.930 65.600 ;
        RECT 5.930 64.800 6.330 65.400 ;
        RECT 5.930 64.600 9.930 64.800 ;
        RECT 5.930 64.000 6.330 64.600 ;
        RECT 5.930 63.800 9.930 64.000 ;
        RECT 5.930 63.200 6.330 63.800 ;
        RECT 5.930 63.000 9.930 63.200 ;
        RECT 5.930 62.400 6.330 63.000 ;
        RECT 5.930 62.200 9.930 62.400 ;
        RECT 10.680 62.200 10.880 69.800 ;
        RECT 11.480 62.200 11.680 69.800 ;
        RECT 12.280 62.200 12.480 69.800 ;
        RECT 13.080 62.200 13.280 69.800 ;
        RECT 13.880 62.200 14.080 69.800 ;
        RECT 15.380 70.200 15.580 77.800 ;
        RECT 16.180 70.200 16.380 77.800 ;
        RECT 16.980 70.200 17.180 77.800 ;
        RECT 17.780 70.200 17.980 77.800 ;
        RECT 18.580 70.200 18.780 77.800 ;
        RECT 19.530 77.600 23.530 77.800 ;
        RECT 23.130 77.000 23.530 77.600 ;
        RECT 19.530 76.800 23.530 77.000 ;
        RECT 23.130 76.200 23.530 76.800 ;
        RECT 19.530 76.000 23.530 76.200 ;
        RECT 23.130 75.400 23.530 76.000 ;
        RECT 19.530 75.200 23.530 75.400 ;
        RECT 23.130 74.600 23.530 75.200 ;
        RECT 19.530 74.400 23.530 74.600 ;
        RECT 23.130 73.800 23.530 74.400 ;
        RECT 19.530 73.600 23.530 73.800 ;
        RECT 23.130 73.000 23.530 73.600 ;
        RECT 19.530 72.800 23.530 73.000 ;
        RECT 23.130 72.200 23.530 72.800 ;
        RECT 19.530 72.000 23.530 72.200 ;
        RECT 23.130 71.400 23.530 72.000 ;
        RECT 19.530 71.200 23.530 71.400 ;
        RECT 23.130 70.600 23.530 71.200 ;
        RECT 19.530 70.400 23.530 70.600 ;
        RECT 23.130 70.200 23.530 70.400 ;
        RECT 15.380 69.800 23.530 70.200 ;
        RECT 15.380 62.200 15.580 69.800 ;
        RECT 16.180 62.200 16.380 69.800 ;
        RECT 16.980 62.200 17.180 69.800 ;
        RECT 17.780 62.200 17.980 69.800 ;
        RECT 18.580 62.200 18.780 69.800 ;
        RECT 23.130 69.600 23.530 69.800 ;
        RECT 19.530 69.400 23.530 69.600 ;
        RECT 23.130 68.800 23.530 69.400 ;
        RECT 19.530 68.600 23.530 68.800 ;
        RECT 23.130 68.000 23.530 68.600 ;
        RECT 19.530 67.800 23.530 68.000 ;
        RECT 23.130 67.200 23.530 67.800 ;
        RECT 19.530 67.000 23.530 67.200 ;
        RECT 23.130 66.400 23.530 67.000 ;
        RECT 19.530 66.200 23.530 66.400 ;
        RECT 23.130 65.600 23.530 66.200 ;
        RECT 19.530 65.400 23.530 65.600 ;
        RECT 23.130 64.800 23.530 65.400 ;
        RECT 19.530 64.600 23.530 64.800 ;
        RECT 23.130 64.000 23.530 64.600 ;
        RECT 19.530 63.800 23.530 64.000 ;
        RECT 23.130 63.200 23.530 63.800 ;
        RECT 19.530 63.000 23.530 63.200 ;
        RECT 23.130 62.400 23.530 63.000 ;
        RECT 19.530 62.200 23.530 62.400 ;
        RECT 25.930 77.600 29.930 77.800 ;
        RECT 25.930 77.000 26.330 77.600 ;
        RECT 25.930 76.800 29.930 77.000 ;
        RECT 25.930 76.200 26.330 76.800 ;
        RECT 25.930 76.000 29.930 76.200 ;
        RECT 25.930 75.400 26.330 76.000 ;
        RECT 25.930 75.200 29.930 75.400 ;
        RECT 25.930 74.600 26.330 75.200 ;
        RECT 25.930 74.400 29.930 74.600 ;
        RECT 25.930 73.800 26.330 74.400 ;
        RECT 25.930 73.600 29.930 73.800 ;
        RECT 25.930 73.000 26.330 73.600 ;
        RECT 25.930 72.800 29.930 73.000 ;
        RECT 25.930 72.200 26.330 72.800 ;
        RECT 25.930 72.000 29.930 72.200 ;
        RECT 25.930 71.400 26.330 72.000 ;
        RECT 25.930 71.200 29.930 71.400 ;
        RECT 25.930 70.600 26.330 71.200 ;
        RECT 25.930 70.400 29.930 70.600 ;
        RECT 25.930 70.200 26.330 70.400 ;
        RECT 30.680 70.200 30.880 77.800 ;
        RECT 31.480 70.200 31.680 77.800 ;
        RECT 32.280 70.200 32.480 77.800 ;
        RECT 33.080 70.200 33.280 77.800 ;
        RECT 33.880 70.200 34.080 77.800 ;
        RECT 25.930 69.800 34.080 70.200 ;
        RECT 25.930 69.600 26.330 69.800 ;
        RECT 25.930 69.400 29.930 69.600 ;
        RECT 25.930 68.800 26.330 69.400 ;
        RECT 25.930 68.600 29.930 68.800 ;
        RECT 25.930 68.000 26.330 68.600 ;
        RECT 25.930 67.800 29.930 68.000 ;
        RECT 25.930 67.200 26.330 67.800 ;
        RECT 25.930 67.000 29.930 67.200 ;
        RECT 25.930 66.400 26.330 67.000 ;
        RECT 25.930 66.200 29.930 66.400 ;
        RECT 25.930 65.600 26.330 66.200 ;
        RECT 25.930 65.400 29.930 65.600 ;
        RECT 25.930 64.800 26.330 65.400 ;
        RECT 25.930 64.600 29.930 64.800 ;
        RECT 25.930 64.000 26.330 64.600 ;
        RECT 25.930 63.800 29.930 64.000 ;
        RECT 25.930 63.200 26.330 63.800 ;
        RECT 25.930 63.000 29.930 63.200 ;
        RECT 25.930 62.400 26.330 63.000 ;
        RECT 25.930 62.200 29.930 62.400 ;
        RECT 30.680 62.200 30.880 69.800 ;
        RECT 31.480 62.200 31.680 69.800 ;
        RECT 32.280 62.200 32.480 69.800 ;
        RECT 33.080 62.200 33.280 69.800 ;
        RECT 33.880 62.200 34.080 69.800 ;
        RECT 35.380 70.200 35.580 77.800 ;
        RECT 36.180 70.200 36.380 77.800 ;
        RECT 36.980 70.200 37.180 77.800 ;
        RECT 37.780 70.200 37.980 77.800 ;
        RECT 38.580 70.200 38.780 77.800 ;
        RECT 39.530 77.600 43.530 77.800 ;
        RECT 43.130 77.000 43.530 77.600 ;
        RECT 39.530 76.800 43.530 77.000 ;
        RECT 43.130 76.200 43.530 76.800 ;
        RECT 39.530 76.000 43.530 76.200 ;
        RECT 43.130 75.400 43.530 76.000 ;
        RECT 39.530 75.200 43.530 75.400 ;
        RECT 43.130 74.600 43.530 75.200 ;
        RECT 39.530 74.400 43.530 74.600 ;
        RECT 43.130 73.800 43.530 74.400 ;
        RECT 39.530 73.600 43.530 73.800 ;
        RECT 43.130 73.000 43.530 73.600 ;
        RECT 39.530 72.800 43.530 73.000 ;
        RECT 43.130 72.200 43.530 72.800 ;
        RECT 39.530 72.000 43.530 72.200 ;
        RECT 43.130 71.400 43.530 72.000 ;
        RECT 39.530 71.200 43.530 71.400 ;
        RECT 43.130 70.600 43.530 71.200 ;
        RECT 39.530 70.400 43.530 70.600 ;
        RECT 43.130 70.200 43.530 70.400 ;
        RECT 35.380 69.800 43.530 70.200 ;
        RECT 35.380 62.200 35.580 69.800 ;
        RECT 36.180 62.200 36.380 69.800 ;
        RECT 36.980 62.200 37.180 69.800 ;
        RECT 37.780 62.200 37.980 69.800 ;
        RECT 38.580 62.200 38.780 69.800 ;
        RECT 43.130 69.600 43.530 69.800 ;
        RECT 39.530 69.400 43.530 69.600 ;
        RECT 43.130 68.800 43.530 69.400 ;
        RECT 39.530 68.600 43.530 68.800 ;
        RECT 43.130 68.000 43.530 68.600 ;
        RECT 39.530 67.800 43.530 68.000 ;
        RECT 43.130 67.200 43.530 67.800 ;
        RECT 39.530 67.000 43.530 67.200 ;
        RECT 43.130 66.400 43.530 67.000 ;
        RECT 39.530 66.200 43.530 66.400 ;
        RECT 43.130 65.600 43.530 66.200 ;
        RECT 39.530 65.400 43.530 65.600 ;
        RECT 43.130 64.800 43.530 65.400 ;
        RECT 39.530 64.600 43.530 64.800 ;
        RECT 43.130 64.000 43.530 64.600 ;
        RECT 39.530 63.800 43.530 64.000 ;
        RECT 43.130 63.200 43.530 63.800 ;
        RECT 39.530 63.000 43.530 63.200 ;
        RECT 43.130 62.400 43.530 63.000 ;
        RECT 39.530 62.200 43.530 62.400 ;
        RECT 45.930 77.600 49.930 77.800 ;
        RECT 45.930 77.000 46.330 77.600 ;
        RECT 45.930 76.800 49.930 77.000 ;
        RECT 45.930 76.200 46.330 76.800 ;
        RECT 45.930 76.000 49.930 76.200 ;
        RECT 45.930 75.400 46.330 76.000 ;
        RECT 45.930 75.200 49.930 75.400 ;
        RECT 45.930 74.600 46.330 75.200 ;
        RECT 45.930 74.400 49.930 74.600 ;
        RECT 45.930 73.800 46.330 74.400 ;
        RECT 45.930 73.600 49.930 73.800 ;
        RECT 45.930 73.000 46.330 73.600 ;
        RECT 45.930 72.800 49.930 73.000 ;
        RECT 45.930 72.200 46.330 72.800 ;
        RECT 45.930 72.000 49.930 72.200 ;
        RECT 45.930 71.400 46.330 72.000 ;
        RECT 45.930 71.200 49.930 71.400 ;
        RECT 45.930 70.600 46.330 71.200 ;
        RECT 45.930 70.400 49.930 70.600 ;
        RECT 45.930 70.200 46.330 70.400 ;
        RECT 50.680 70.200 50.880 77.800 ;
        RECT 51.480 70.200 51.680 77.800 ;
        RECT 52.280 70.200 52.480 77.800 ;
        RECT 53.080 70.200 53.280 77.800 ;
        RECT 53.880 70.200 54.080 77.800 ;
        RECT 45.930 69.800 54.080 70.200 ;
        RECT 45.930 69.600 46.330 69.800 ;
        RECT 45.930 69.400 49.930 69.600 ;
        RECT 45.930 68.800 46.330 69.400 ;
        RECT 45.930 68.600 49.930 68.800 ;
        RECT 45.930 68.000 46.330 68.600 ;
        RECT 45.930 67.800 49.930 68.000 ;
        RECT 45.930 67.200 46.330 67.800 ;
        RECT 45.930 67.000 49.930 67.200 ;
        RECT 45.930 66.400 46.330 67.000 ;
        RECT 45.930 66.200 49.930 66.400 ;
        RECT 45.930 65.600 46.330 66.200 ;
        RECT 45.930 65.400 49.930 65.600 ;
        RECT 45.930 64.800 46.330 65.400 ;
        RECT 45.930 64.600 49.930 64.800 ;
        RECT 45.930 64.000 46.330 64.600 ;
        RECT 45.930 63.800 49.930 64.000 ;
        RECT 45.930 63.200 46.330 63.800 ;
        RECT 45.930 63.000 49.930 63.200 ;
        RECT 45.930 62.400 46.330 63.000 ;
        RECT 45.930 62.200 49.930 62.400 ;
        RECT 50.680 62.200 50.880 69.800 ;
        RECT 51.480 62.200 51.680 69.800 ;
        RECT 52.280 62.200 52.480 69.800 ;
        RECT 53.080 62.200 53.280 69.800 ;
        RECT 53.880 62.200 54.080 69.800 ;
        RECT 55.380 70.200 55.580 77.800 ;
        RECT 56.180 70.200 56.380 77.800 ;
        RECT 56.980 70.200 57.180 77.800 ;
        RECT 57.780 70.200 57.980 77.800 ;
        RECT 58.580 70.200 58.780 77.800 ;
        RECT 59.530 77.600 63.530 77.800 ;
        RECT 63.130 77.000 63.530 77.600 ;
        RECT 59.530 76.800 63.530 77.000 ;
        RECT 63.130 76.200 63.530 76.800 ;
        RECT 59.530 76.000 63.530 76.200 ;
        RECT 63.130 75.400 63.530 76.000 ;
        RECT 59.530 75.200 63.530 75.400 ;
        RECT 63.130 74.600 63.530 75.200 ;
        RECT 59.530 74.400 63.530 74.600 ;
        RECT 63.130 73.800 63.530 74.400 ;
        RECT 59.530 73.600 63.530 73.800 ;
        RECT 63.130 73.000 63.530 73.600 ;
        RECT 59.530 72.800 63.530 73.000 ;
        RECT 63.130 72.200 63.530 72.800 ;
        RECT 59.530 72.000 63.530 72.200 ;
        RECT 63.130 71.400 63.530 72.000 ;
        RECT 59.530 71.200 63.530 71.400 ;
        RECT 63.130 70.600 63.530 71.200 ;
        RECT 59.530 70.400 63.530 70.600 ;
        RECT 63.130 70.200 63.530 70.400 ;
        RECT 55.380 69.800 63.530 70.200 ;
        RECT 55.380 62.200 55.580 69.800 ;
        RECT 56.180 62.200 56.380 69.800 ;
        RECT 56.980 62.200 57.180 69.800 ;
        RECT 57.780 62.200 57.980 69.800 ;
        RECT 58.580 62.200 58.780 69.800 ;
        RECT 63.130 69.600 63.530 69.800 ;
        RECT 59.530 69.400 63.530 69.600 ;
        RECT 63.130 68.800 63.530 69.400 ;
        RECT 59.530 68.600 63.530 68.800 ;
        RECT 63.130 68.000 63.530 68.600 ;
        RECT 59.530 67.800 63.530 68.000 ;
        RECT 63.130 67.200 63.530 67.800 ;
        RECT 59.530 67.000 63.530 67.200 ;
        RECT 63.130 66.400 63.530 67.000 ;
        RECT 59.530 66.200 63.530 66.400 ;
        RECT 63.130 65.600 63.530 66.200 ;
        RECT 59.530 65.400 63.530 65.600 ;
        RECT 63.130 64.800 63.530 65.400 ;
        RECT 59.530 64.600 63.530 64.800 ;
        RECT 63.130 64.000 63.530 64.600 ;
        RECT 59.530 63.800 63.530 64.000 ;
        RECT 63.130 63.200 63.530 63.800 ;
        RECT 59.530 63.000 63.530 63.200 ;
        RECT 63.130 62.400 63.530 63.000 ;
        RECT 59.530 62.200 63.530 62.400 ;
        RECT 65.930 77.600 69.930 77.800 ;
        RECT 65.930 77.000 66.330 77.600 ;
        RECT 65.930 76.800 69.930 77.000 ;
        RECT 65.930 76.200 66.330 76.800 ;
        RECT 65.930 76.000 69.930 76.200 ;
        RECT 65.930 75.400 66.330 76.000 ;
        RECT 65.930 75.200 69.930 75.400 ;
        RECT 65.930 74.600 66.330 75.200 ;
        RECT 65.930 74.400 69.930 74.600 ;
        RECT 65.930 73.800 66.330 74.400 ;
        RECT 65.930 73.600 69.930 73.800 ;
        RECT 65.930 73.000 66.330 73.600 ;
        RECT 65.930 72.800 69.930 73.000 ;
        RECT 65.930 72.200 66.330 72.800 ;
        RECT 65.930 72.000 69.930 72.200 ;
        RECT 65.930 71.400 66.330 72.000 ;
        RECT 65.930 71.200 69.930 71.400 ;
        RECT 65.930 70.600 66.330 71.200 ;
        RECT 65.930 70.400 69.930 70.600 ;
        RECT 65.930 70.200 66.330 70.400 ;
        RECT 70.680 70.200 70.880 77.800 ;
        RECT 71.480 70.200 71.680 77.800 ;
        RECT 72.280 70.200 72.480 77.800 ;
        RECT 73.080 70.200 73.280 77.800 ;
        RECT 73.880 70.200 74.080 77.800 ;
        RECT 65.930 69.800 74.080 70.200 ;
        RECT 65.930 69.600 66.330 69.800 ;
        RECT 65.930 69.400 69.930 69.600 ;
        RECT 65.930 68.800 66.330 69.400 ;
        RECT 65.930 68.600 69.930 68.800 ;
        RECT 65.930 68.000 66.330 68.600 ;
        RECT 65.930 67.800 69.930 68.000 ;
        RECT 65.930 67.200 66.330 67.800 ;
        RECT 65.930 67.000 69.930 67.200 ;
        RECT 65.930 66.400 66.330 67.000 ;
        RECT 65.930 66.200 69.930 66.400 ;
        RECT 65.930 65.600 66.330 66.200 ;
        RECT 65.930 65.400 69.930 65.600 ;
        RECT 65.930 64.800 66.330 65.400 ;
        RECT 65.930 64.600 69.930 64.800 ;
        RECT 65.930 64.000 66.330 64.600 ;
        RECT 65.930 63.800 69.930 64.000 ;
        RECT 65.930 63.200 66.330 63.800 ;
        RECT 65.930 63.000 69.930 63.200 ;
        RECT 65.930 62.400 66.330 63.000 ;
        RECT 65.930 62.200 69.930 62.400 ;
        RECT 70.680 62.200 70.880 69.800 ;
        RECT 71.480 62.200 71.680 69.800 ;
        RECT 72.280 62.200 72.480 69.800 ;
        RECT 73.080 62.200 73.280 69.800 ;
        RECT 73.880 62.200 74.080 69.800 ;
        RECT 75.380 70.200 75.580 77.800 ;
        RECT 76.180 70.200 76.380 77.800 ;
        RECT 76.980 70.200 77.180 77.800 ;
        RECT 77.780 70.200 77.980 77.800 ;
        RECT 78.580 70.200 78.780 77.800 ;
        RECT 79.530 77.600 83.530 77.800 ;
        RECT 83.130 77.000 83.530 77.600 ;
        RECT 79.530 76.800 83.530 77.000 ;
        RECT 83.130 76.200 83.530 76.800 ;
        RECT 79.530 76.000 83.530 76.200 ;
        RECT 83.130 75.400 83.530 76.000 ;
        RECT 79.530 75.200 83.530 75.400 ;
        RECT 83.130 74.600 83.530 75.200 ;
        RECT 79.530 74.400 83.530 74.600 ;
        RECT 83.130 73.800 83.530 74.400 ;
        RECT 79.530 73.600 83.530 73.800 ;
        RECT 83.130 73.000 83.530 73.600 ;
        RECT 79.530 72.800 83.530 73.000 ;
        RECT 83.130 72.200 83.530 72.800 ;
        RECT 79.530 72.000 83.530 72.200 ;
        RECT 83.130 71.400 83.530 72.000 ;
        RECT 79.530 71.200 83.530 71.400 ;
        RECT 83.130 70.600 83.530 71.200 ;
        RECT 79.530 70.400 83.530 70.600 ;
        RECT 83.130 70.200 83.530 70.400 ;
        RECT 75.380 69.800 83.530 70.200 ;
        RECT 75.380 62.200 75.580 69.800 ;
        RECT 76.180 62.200 76.380 69.800 ;
        RECT 76.980 62.200 77.180 69.800 ;
        RECT 77.780 62.200 77.980 69.800 ;
        RECT 78.580 62.200 78.780 69.800 ;
        RECT 83.130 69.600 83.530 69.800 ;
        RECT 79.530 69.400 83.530 69.600 ;
        RECT 83.130 68.800 83.530 69.400 ;
        RECT 79.530 68.600 83.530 68.800 ;
        RECT 83.130 68.000 83.530 68.600 ;
        RECT 79.530 67.800 83.530 68.000 ;
        RECT 83.130 67.200 83.530 67.800 ;
        RECT 79.530 67.000 83.530 67.200 ;
        RECT 83.130 66.400 83.530 67.000 ;
        RECT 79.530 66.200 83.530 66.400 ;
        RECT 83.130 65.600 83.530 66.200 ;
        RECT 79.530 65.400 83.530 65.600 ;
        RECT 83.130 64.800 83.530 65.400 ;
        RECT 79.530 64.600 83.530 64.800 ;
        RECT 83.130 64.000 83.530 64.600 ;
        RECT 79.530 63.800 83.530 64.000 ;
        RECT 83.130 63.200 83.530 63.800 ;
        RECT 79.530 63.000 83.530 63.200 ;
        RECT 83.130 62.400 83.530 63.000 ;
        RECT 79.530 62.200 83.530 62.400 ;
        RECT 85.930 77.600 89.930 77.800 ;
        RECT 85.930 77.000 86.330 77.600 ;
        RECT 85.930 76.800 89.930 77.000 ;
        RECT 85.930 76.200 86.330 76.800 ;
        RECT 85.930 76.000 89.930 76.200 ;
        RECT 85.930 75.400 86.330 76.000 ;
        RECT 85.930 75.200 89.930 75.400 ;
        RECT 85.930 74.600 86.330 75.200 ;
        RECT 85.930 74.400 89.930 74.600 ;
        RECT 85.930 73.800 86.330 74.400 ;
        RECT 85.930 73.600 89.930 73.800 ;
        RECT 85.930 73.000 86.330 73.600 ;
        RECT 85.930 72.800 89.930 73.000 ;
        RECT 85.930 72.200 86.330 72.800 ;
        RECT 85.930 72.000 89.930 72.200 ;
        RECT 85.930 71.400 86.330 72.000 ;
        RECT 85.930 71.200 89.930 71.400 ;
        RECT 85.930 70.600 86.330 71.200 ;
        RECT 85.930 70.400 89.930 70.600 ;
        RECT 85.930 70.200 86.330 70.400 ;
        RECT 90.680 70.200 90.880 77.800 ;
        RECT 91.480 70.200 91.680 77.800 ;
        RECT 92.280 70.200 92.480 77.800 ;
        RECT 93.080 70.200 93.280 77.800 ;
        RECT 93.880 70.200 94.080 77.800 ;
        RECT 85.930 69.800 94.080 70.200 ;
        RECT 85.930 69.600 86.330 69.800 ;
        RECT 85.930 69.400 89.930 69.600 ;
        RECT 85.930 68.800 86.330 69.400 ;
        RECT 85.930 68.600 89.930 68.800 ;
        RECT 85.930 68.000 86.330 68.600 ;
        RECT 85.930 67.800 89.930 68.000 ;
        RECT 85.930 67.200 86.330 67.800 ;
        RECT 85.930 67.000 89.930 67.200 ;
        RECT 85.930 66.400 86.330 67.000 ;
        RECT 85.930 66.200 89.930 66.400 ;
        RECT 85.930 65.600 86.330 66.200 ;
        RECT 85.930 65.400 89.930 65.600 ;
        RECT 85.930 64.800 86.330 65.400 ;
        RECT 85.930 64.600 89.930 64.800 ;
        RECT 85.930 64.000 86.330 64.600 ;
        RECT 85.930 63.800 89.930 64.000 ;
        RECT 85.930 63.200 86.330 63.800 ;
        RECT 85.930 63.000 89.930 63.200 ;
        RECT 85.930 62.400 86.330 63.000 ;
        RECT 85.930 62.200 89.930 62.400 ;
        RECT 90.680 62.200 90.880 69.800 ;
        RECT 91.480 62.200 91.680 69.800 ;
        RECT 92.280 62.200 92.480 69.800 ;
        RECT 93.080 62.200 93.280 69.800 ;
        RECT 93.880 62.200 94.080 69.800 ;
        RECT 95.380 70.200 95.580 77.800 ;
        RECT 96.180 70.200 96.380 77.800 ;
        RECT 96.980 70.200 97.180 77.800 ;
        RECT 97.780 70.200 97.980 77.800 ;
        RECT 98.580 70.200 98.780 77.800 ;
        RECT 99.530 77.600 103.530 77.800 ;
        RECT 103.130 77.000 103.530 77.600 ;
        RECT 99.530 76.800 103.530 77.000 ;
        RECT 103.130 76.200 103.530 76.800 ;
        RECT 99.530 76.000 103.530 76.200 ;
        RECT 103.130 75.400 103.530 76.000 ;
        RECT 99.530 75.200 103.530 75.400 ;
        RECT 103.130 74.600 103.530 75.200 ;
        RECT 99.530 74.400 103.530 74.600 ;
        RECT 103.130 73.800 103.530 74.400 ;
        RECT 99.530 73.600 103.530 73.800 ;
        RECT 103.130 73.000 103.530 73.600 ;
        RECT 99.530 72.800 103.530 73.000 ;
        RECT 103.130 72.200 103.530 72.800 ;
        RECT 99.530 72.000 103.530 72.200 ;
        RECT 103.130 71.400 103.530 72.000 ;
        RECT 99.530 71.200 103.530 71.400 ;
        RECT 103.130 70.600 103.530 71.200 ;
        RECT 110.050 70.900 110.410 71.280 ;
        RECT 110.680 70.900 111.040 71.280 ;
        RECT 111.280 70.900 111.640 71.280 ;
        RECT 99.530 70.400 103.530 70.600 ;
        RECT 103.130 70.200 103.530 70.400 ;
        RECT 110.050 70.310 110.410 70.690 ;
        RECT 110.680 70.310 111.040 70.690 ;
        RECT 111.280 70.310 111.640 70.690 ;
        RECT 95.380 69.800 103.530 70.200 ;
        RECT 95.380 62.200 95.580 69.800 ;
        RECT 96.180 62.200 96.380 69.800 ;
        RECT 96.980 62.200 97.180 69.800 ;
        RECT 97.780 62.200 97.980 69.800 ;
        RECT 98.580 62.200 98.780 69.800 ;
        RECT 103.130 69.600 103.530 69.800 ;
        RECT 99.530 69.400 103.530 69.600 ;
        RECT 103.130 68.800 103.530 69.400 ;
        RECT 99.530 68.600 103.530 68.800 ;
        RECT 103.130 68.000 103.530 68.600 ;
        RECT 99.530 67.800 103.530 68.000 ;
        RECT 103.130 67.200 103.530 67.800 ;
        RECT 99.530 67.000 103.530 67.200 ;
        RECT 103.130 66.400 103.530 67.000 ;
        RECT 99.530 66.200 103.530 66.400 ;
        RECT 103.130 65.600 103.530 66.200 ;
        RECT 99.530 65.400 103.530 65.600 ;
        RECT 103.130 64.800 103.530 65.400 ;
        RECT 99.530 64.600 103.530 64.800 ;
        RECT 103.130 64.000 103.530 64.600 ;
        RECT 99.530 63.800 103.530 64.000 ;
        RECT 103.130 63.200 103.530 63.800 ;
        RECT 99.530 63.000 103.530 63.200 ;
        RECT 103.130 62.400 103.530 63.000 ;
        RECT 99.530 62.200 103.530 62.400 ;
        RECT 5.930 57.600 9.930 57.800 ;
        RECT 5.930 57.000 6.330 57.600 ;
        RECT 5.930 56.800 9.930 57.000 ;
        RECT 5.930 56.200 6.330 56.800 ;
        RECT 5.930 56.000 9.930 56.200 ;
        RECT 5.930 55.400 6.330 56.000 ;
        RECT 5.930 55.200 9.930 55.400 ;
        RECT 5.930 54.600 6.330 55.200 ;
        RECT 5.930 54.400 9.930 54.600 ;
        RECT 5.930 53.800 6.330 54.400 ;
        RECT 5.930 53.600 9.930 53.800 ;
        RECT 5.930 53.000 6.330 53.600 ;
        RECT 5.930 52.800 9.930 53.000 ;
        RECT 5.930 52.200 6.330 52.800 ;
        RECT 5.930 52.000 9.930 52.200 ;
        RECT 5.930 51.400 6.330 52.000 ;
        RECT 5.930 51.200 9.930 51.400 ;
        RECT 5.930 50.600 6.330 51.200 ;
        RECT 5.930 50.400 9.930 50.600 ;
        RECT 5.930 50.200 6.330 50.400 ;
        RECT 10.680 50.200 10.880 57.800 ;
        RECT 11.480 50.200 11.680 57.800 ;
        RECT 12.280 50.200 12.480 57.800 ;
        RECT 13.080 50.200 13.280 57.800 ;
        RECT 13.880 50.200 14.080 57.800 ;
        RECT 5.930 49.800 14.080 50.200 ;
        RECT 5.930 49.600 6.330 49.800 ;
        RECT 5.930 49.400 9.930 49.600 ;
        RECT 5.930 48.800 6.330 49.400 ;
        RECT 5.930 48.600 9.930 48.800 ;
        RECT 5.930 48.000 6.330 48.600 ;
        RECT 5.930 47.800 9.930 48.000 ;
        RECT 5.930 47.200 6.330 47.800 ;
        RECT 5.930 47.000 9.930 47.200 ;
        RECT 5.930 46.400 6.330 47.000 ;
        RECT 5.930 46.200 9.930 46.400 ;
        RECT 5.930 45.600 6.330 46.200 ;
        RECT 5.930 45.400 9.930 45.600 ;
        RECT 5.930 44.800 6.330 45.400 ;
        RECT 5.930 44.600 9.930 44.800 ;
        RECT 5.930 44.000 6.330 44.600 ;
        RECT 5.930 43.800 9.930 44.000 ;
        RECT 5.930 43.200 6.330 43.800 ;
        RECT 5.930 43.000 9.930 43.200 ;
        RECT 5.930 42.400 6.330 43.000 ;
        RECT 5.930 42.200 9.930 42.400 ;
        RECT 10.680 42.200 10.880 49.800 ;
        RECT 11.480 42.200 11.680 49.800 ;
        RECT 12.280 42.200 12.480 49.800 ;
        RECT 13.080 42.200 13.280 49.800 ;
        RECT 13.880 42.200 14.080 49.800 ;
        RECT 15.380 50.200 15.580 57.800 ;
        RECT 16.180 50.200 16.380 57.800 ;
        RECT 16.980 50.200 17.180 57.800 ;
        RECT 17.780 50.200 17.980 57.800 ;
        RECT 18.580 50.200 18.780 57.800 ;
        RECT 19.530 57.600 23.530 57.800 ;
        RECT 23.130 57.000 23.530 57.600 ;
        RECT 19.530 56.800 23.530 57.000 ;
        RECT 23.130 56.200 23.530 56.800 ;
        RECT 19.530 56.000 23.530 56.200 ;
        RECT 23.130 55.400 23.530 56.000 ;
        RECT 19.530 55.200 23.530 55.400 ;
        RECT 23.130 54.600 23.530 55.200 ;
        RECT 19.530 54.400 23.530 54.600 ;
        RECT 23.130 53.800 23.530 54.400 ;
        RECT 19.530 53.600 23.530 53.800 ;
        RECT 23.130 53.000 23.530 53.600 ;
        RECT 19.530 52.800 23.530 53.000 ;
        RECT 23.130 52.200 23.530 52.800 ;
        RECT 19.530 52.000 23.530 52.200 ;
        RECT 23.130 51.400 23.530 52.000 ;
        RECT 19.530 51.200 23.530 51.400 ;
        RECT 23.130 50.600 23.530 51.200 ;
        RECT 19.530 50.400 23.530 50.600 ;
        RECT 23.130 50.200 23.530 50.400 ;
        RECT 15.380 49.800 23.530 50.200 ;
        RECT 15.380 42.200 15.580 49.800 ;
        RECT 16.180 42.200 16.380 49.800 ;
        RECT 16.980 42.200 17.180 49.800 ;
        RECT 17.780 42.200 17.980 49.800 ;
        RECT 18.580 42.200 18.780 49.800 ;
        RECT 23.130 49.600 23.530 49.800 ;
        RECT 19.530 49.400 23.530 49.600 ;
        RECT 23.130 48.800 23.530 49.400 ;
        RECT 19.530 48.600 23.530 48.800 ;
        RECT 23.130 48.000 23.530 48.600 ;
        RECT 19.530 47.800 23.530 48.000 ;
        RECT 23.130 47.200 23.530 47.800 ;
        RECT 19.530 47.000 23.530 47.200 ;
        RECT 23.130 46.400 23.530 47.000 ;
        RECT 19.530 46.200 23.530 46.400 ;
        RECT 23.130 45.600 23.530 46.200 ;
        RECT 19.530 45.400 23.530 45.600 ;
        RECT 23.130 44.800 23.530 45.400 ;
        RECT 19.530 44.600 23.530 44.800 ;
        RECT 23.130 44.000 23.530 44.600 ;
        RECT 19.530 43.800 23.530 44.000 ;
        RECT 23.130 43.200 23.530 43.800 ;
        RECT 19.530 43.000 23.530 43.200 ;
        RECT 23.130 42.400 23.530 43.000 ;
        RECT 19.530 42.200 23.530 42.400 ;
        RECT 25.930 57.600 29.930 57.800 ;
        RECT 25.930 57.000 26.330 57.600 ;
        RECT 25.930 56.800 29.930 57.000 ;
        RECT 25.930 56.200 26.330 56.800 ;
        RECT 25.930 56.000 29.930 56.200 ;
        RECT 25.930 55.400 26.330 56.000 ;
        RECT 25.930 55.200 29.930 55.400 ;
        RECT 25.930 54.600 26.330 55.200 ;
        RECT 25.930 54.400 29.930 54.600 ;
        RECT 25.930 53.800 26.330 54.400 ;
        RECT 25.930 53.600 29.930 53.800 ;
        RECT 25.930 53.000 26.330 53.600 ;
        RECT 25.930 52.800 29.930 53.000 ;
        RECT 25.930 52.200 26.330 52.800 ;
        RECT 25.930 52.000 29.930 52.200 ;
        RECT 25.930 51.400 26.330 52.000 ;
        RECT 25.930 51.200 29.930 51.400 ;
        RECT 25.930 50.600 26.330 51.200 ;
        RECT 25.930 50.400 29.930 50.600 ;
        RECT 25.930 50.200 26.330 50.400 ;
        RECT 30.680 50.200 30.880 57.800 ;
        RECT 31.480 50.200 31.680 57.800 ;
        RECT 32.280 50.200 32.480 57.800 ;
        RECT 33.080 50.200 33.280 57.800 ;
        RECT 33.880 50.200 34.080 57.800 ;
        RECT 25.930 49.800 34.080 50.200 ;
        RECT 25.930 49.600 26.330 49.800 ;
        RECT 25.930 49.400 29.930 49.600 ;
        RECT 25.930 48.800 26.330 49.400 ;
        RECT 25.930 48.600 29.930 48.800 ;
        RECT 25.930 48.000 26.330 48.600 ;
        RECT 25.930 47.800 29.930 48.000 ;
        RECT 25.930 47.200 26.330 47.800 ;
        RECT 25.930 47.000 29.930 47.200 ;
        RECT 25.930 46.400 26.330 47.000 ;
        RECT 25.930 46.200 29.930 46.400 ;
        RECT 25.930 45.600 26.330 46.200 ;
        RECT 25.930 45.400 29.930 45.600 ;
        RECT 25.930 44.800 26.330 45.400 ;
        RECT 25.930 44.600 29.930 44.800 ;
        RECT 25.930 44.000 26.330 44.600 ;
        RECT 25.930 43.800 29.930 44.000 ;
        RECT 25.930 43.200 26.330 43.800 ;
        RECT 25.930 43.000 29.930 43.200 ;
        RECT 25.930 42.400 26.330 43.000 ;
        RECT 25.930 42.200 29.930 42.400 ;
        RECT 30.680 42.200 30.880 49.800 ;
        RECT 31.480 42.200 31.680 49.800 ;
        RECT 32.280 42.200 32.480 49.800 ;
        RECT 33.080 42.200 33.280 49.800 ;
        RECT 33.880 42.200 34.080 49.800 ;
        RECT 35.380 50.200 35.580 57.800 ;
        RECT 36.180 50.200 36.380 57.800 ;
        RECT 36.980 50.200 37.180 57.800 ;
        RECT 37.780 50.200 37.980 57.800 ;
        RECT 38.580 50.200 38.780 57.800 ;
        RECT 39.530 57.600 43.530 57.800 ;
        RECT 43.130 57.000 43.530 57.600 ;
        RECT 39.530 56.800 43.530 57.000 ;
        RECT 43.130 56.200 43.530 56.800 ;
        RECT 39.530 56.000 43.530 56.200 ;
        RECT 43.130 55.400 43.530 56.000 ;
        RECT 39.530 55.200 43.530 55.400 ;
        RECT 43.130 54.600 43.530 55.200 ;
        RECT 39.530 54.400 43.530 54.600 ;
        RECT 43.130 53.800 43.530 54.400 ;
        RECT 39.530 53.600 43.530 53.800 ;
        RECT 43.130 53.000 43.530 53.600 ;
        RECT 39.530 52.800 43.530 53.000 ;
        RECT 43.130 52.200 43.530 52.800 ;
        RECT 39.530 52.000 43.530 52.200 ;
        RECT 43.130 51.400 43.530 52.000 ;
        RECT 39.530 51.200 43.530 51.400 ;
        RECT 43.130 50.600 43.530 51.200 ;
        RECT 39.530 50.400 43.530 50.600 ;
        RECT 43.130 50.200 43.530 50.400 ;
        RECT 35.380 49.800 43.530 50.200 ;
        RECT 35.380 42.200 35.580 49.800 ;
        RECT 36.180 42.200 36.380 49.800 ;
        RECT 36.980 42.200 37.180 49.800 ;
        RECT 37.780 42.200 37.980 49.800 ;
        RECT 38.580 42.200 38.780 49.800 ;
        RECT 43.130 49.600 43.530 49.800 ;
        RECT 39.530 49.400 43.530 49.600 ;
        RECT 43.130 48.800 43.530 49.400 ;
        RECT 39.530 48.600 43.530 48.800 ;
        RECT 43.130 48.000 43.530 48.600 ;
        RECT 39.530 47.800 43.530 48.000 ;
        RECT 43.130 47.200 43.530 47.800 ;
        RECT 39.530 47.000 43.530 47.200 ;
        RECT 43.130 46.400 43.530 47.000 ;
        RECT 39.530 46.200 43.530 46.400 ;
        RECT 43.130 45.600 43.530 46.200 ;
        RECT 39.530 45.400 43.530 45.600 ;
        RECT 43.130 44.800 43.530 45.400 ;
        RECT 39.530 44.600 43.530 44.800 ;
        RECT 43.130 44.000 43.530 44.600 ;
        RECT 39.530 43.800 43.530 44.000 ;
        RECT 43.130 43.200 43.530 43.800 ;
        RECT 39.530 43.000 43.530 43.200 ;
        RECT 43.130 42.400 43.530 43.000 ;
        RECT 39.530 42.200 43.530 42.400 ;
        RECT 45.930 57.600 49.930 57.800 ;
        RECT 45.930 57.000 46.330 57.600 ;
        RECT 45.930 56.800 49.930 57.000 ;
        RECT 45.930 56.200 46.330 56.800 ;
        RECT 45.930 56.000 49.930 56.200 ;
        RECT 45.930 55.400 46.330 56.000 ;
        RECT 45.930 55.200 49.930 55.400 ;
        RECT 45.930 54.600 46.330 55.200 ;
        RECT 45.930 54.400 49.930 54.600 ;
        RECT 45.930 53.800 46.330 54.400 ;
        RECT 45.930 53.600 49.930 53.800 ;
        RECT 45.930 53.000 46.330 53.600 ;
        RECT 45.930 52.800 49.930 53.000 ;
        RECT 45.930 52.200 46.330 52.800 ;
        RECT 45.930 52.000 49.930 52.200 ;
        RECT 45.930 51.400 46.330 52.000 ;
        RECT 45.930 51.200 49.930 51.400 ;
        RECT 45.930 50.600 46.330 51.200 ;
        RECT 45.930 50.400 49.930 50.600 ;
        RECT 45.930 50.200 46.330 50.400 ;
        RECT 50.680 50.200 50.880 57.800 ;
        RECT 51.480 50.200 51.680 57.800 ;
        RECT 52.280 50.200 52.480 57.800 ;
        RECT 53.080 50.200 53.280 57.800 ;
        RECT 53.880 50.200 54.080 57.800 ;
        RECT 45.930 49.800 54.080 50.200 ;
        RECT 45.930 49.600 46.330 49.800 ;
        RECT 45.930 49.400 49.930 49.600 ;
        RECT 45.930 48.800 46.330 49.400 ;
        RECT 45.930 48.600 49.930 48.800 ;
        RECT 45.930 48.000 46.330 48.600 ;
        RECT 45.930 47.800 49.930 48.000 ;
        RECT 45.930 47.200 46.330 47.800 ;
        RECT 45.930 47.000 49.930 47.200 ;
        RECT 45.930 46.400 46.330 47.000 ;
        RECT 45.930 46.200 49.930 46.400 ;
        RECT 45.930 45.600 46.330 46.200 ;
        RECT 45.930 45.400 49.930 45.600 ;
        RECT 45.930 44.800 46.330 45.400 ;
        RECT 45.930 44.600 49.930 44.800 ;
        RECT 45.930 44.000 46.330 44.600 ;
        RECT 45.930 43.800 49.930 44.000 ;
        RECT 45.930 43.200 46.330 43.800 ;
        RECT 45.930 43.000 49.930 43.200 ;
        RECT 45.930 42.400 46.330 43.000 ;
        RECT 45.930 42.200 49.930 42.400 ;
        RECT 50.680 42.200 50.880 49.800 ;
        RECT 51.480 42.200 51.680 49.800 ;
        RECT 52.280 42.200 52.480 49.800 ;
        RECT 53.080 42.200 53.280 49.800 ;
        RECT 53.880 42.200 54.080 49.800 ;
        RECT 55.380 50.200 55.580 57.800 ;
        RECT 56.180 50.200 56.380 57.800 ;
        RECT 56.980 50.200 57.180 57.800 ;
        RECT 57.780 50.200 57.980 57.800 ;
        RECT 58.580 50.200 58.780 57.800 ;
        RECT 59.530 57.600 63.530 57.800 ;
        RECT 63.130 57.000 63.530 57.600 ;
        RECT 59.530 56.800 63.530 57.000 ;
        RECT 63.130 56.200 63.530 56.800 ;
        RECT 59.530 56.000 63.530 56.200 ;
        RECT 63.130 55.400 63.530 56.000 ;
        RECT 59.530 55.200 63.530 55.400 ;
        RECT 63.130 54.600 63.530 55.200 ;
        RECT 59.530 54.400 63.530 54.600 ;
        RECT 63.130 53.800 63.530 54.400 ;
        RECT 59.530 53.600 63.530 53.800 ;
        RECT 63.130 53.000 63.530 53.600 ;
        RECT 59.530 52.800 63.530 53.000 ;
        RECT 63.130 52.200 63.530 52.800 ;
        RECT 59.530 52.000 63.530 52.200 ;
        RECT 63.130 51.400 63.530 52.000 ;
        RECT 59.530 51.200 63.530 51.400 ;
        RECT 63.130 50.600 63.530 51.200 ;
        RECT 59.530 50.400 63.530 50.600 ;
        RECT 63.130 50.200 63.530 50.400 ;
        RECT 55.380 49.800 63.530 50.200 ;
        RECT 55.380 42.200 55.580 49.800 ;
        RECT 56.180 42.200 56.380 49.800 ;
        RECT 56.980 42.200 57.180 49.800 ;
        RECT 57.780 42.200 57.980 49.800 ;
        RECT 58.580 42.200 58.780 49.800 ;
        RECT 63.130 49.600 63.530 49.800 ;
        RECT 59.530 49.400 63.530 49.600 ;
        RECT 63.130 48.800 63.530 49.400 ;
        RECT 59.530 48.600 63.530 48.800 ;
        RECT 63.130 48.000 63.530 48.600 ;
        RECT 59.530 47.800 63.530 48.000 ;
        RECT 63.130 47.200 63.530 47.800 ;
        RECT 59.530 47.000 63.530 47.200 ;
        RECT 63.130 46.400 63.530 47.000 ;
        RECT 59.530 46.200 63.530 46.400 ;
        RECT 63.130 45.600 63.530 46.200 ;
        RECT 59.530 45.400 63.530 45.600 ;
        RECT 63.130 44.800 63.530 45.400 ;
        RECT 59.530 44.600 63.530 44.800 ;
        RECT 63.130 44.000 63.530 44.600 ;
        RECT 59.530 43.800 63.530 44.000 ;
        RECT 63.130 43.200 63.530 43.800 ;
        RECT 59.530 43.000 63.530 43.200 ;
        RECT 63.130 42.400 63.530 43.000 ;
        RECT 59.530 42.200 63.530 42.400 ;
        RECT 65.930 57.600 69.930 57.800 ;
        RECT 65.930 57.000 66.330 57.600 ;
        RECT 65.930 56.800 69.930 57.000 ;
        RECT 65.930 56.200 66.330 56.800 ;
        RECT 65.930 56.000 69.930 56.200 ;
        RECT 65.930 55.400 66.330 56.000 ;
        RECT 65.930 55.200 69.930 55.400 ;
        RECT 65.930 54.600 66.330 55.200 ;
        RECT 65.930 54.400 69.930 54.600 ;
        RECT 65.930 53.800 66.330 54.400 ;
        RECT 65.930 53.600 69.930 53.800 ;
        RECT 65.930 53.000 66.330 53.600 ;
        RECT 65.930 52.800 69.930 53.000 ;
        RECT 65.930 52.200 66.330 52.800 ;
        RECT 65.930 52.000 69.930 52.200 ;
        RECT 65.930 51.400 66.330 52.000 ;
        RECT 65.930 51.200 69.930 51.400 ;
        RECT 65.930 50.600 66.330 51.200 ;
        RECT 65.930 50.400 69.930 50.600 ;
        RECT 65.930 50.200 66.330 50.400 ;
        RECT 70.680 50.200 70.880 57.800 ;
        RECT 71.480 50.200 71.680 57.800 ;
        RECT 72.280 50.200 72.480 57.800 ;
        RECT 73.080 50.200 73.280 57.800 ;
        RECT 73.880 50.200 74.080 57.800 ;
        RECT 65.930 49.800 74.080 50.200 ;
        RECT 65.930 49.600 66.330 49.800 ;
        RECT 65.930 49.400 69.930 49.600 ;
        RECT 65.930 48.800 66.330 49.400 ;
        RECT 65.930 48.600 69.930 48.800 ;
        RECT 65.930 48.000 66.330 48.600 ;
        RECT 65.930 47.800 69.930 48.000 ;
        RECT 65.930 47.200 66.330 47.800 ;
        RECT 65.930 47.000 69.930 47.200 ;
        RECT 65.930 46.400 66.330 47.000 ;
        RECT 65.930 46.200 69.930 46.400 ;
        RECT 65.930 45.600 66.330 46.200 ;
        RECT 65.930 45.400 69.930 45.600 ;
        RECT 65.930 44.800 66.330 45.400 ;
        RECT 65.930 44.600 69.930 44.800 ;
        RECT 65.930 44.000 66.330 44.600 ;
        RECT 65.930 43.800 69.930 44.000 ;
        RECT 65.930 43.200 66.330 43.800 ;
        RECT 65.930 43.000 69.930 43.200 ;
        RECT 65.930 42.400 66.330 43.000 ;
        RECT 65.930 42.200 69.930 42.400 ;
        RECT 70.680 42.200 70.880 49.800 ;
        RECT 71.480 42.200 71.680 49.800 ;
        RECT 72.280 42.200 72.480 49.800 ;
        RECT 73.080 42.200 73.280 49.800 ;
        RECT 73.880 42.200 74.080 49.800 ;
        RECT 75.380 50.200 75.580 57.800 ;
        RECT 76.180 50.200 76.380 57.800 ;
        RECT 76.980 50.200 77.180 57.800 ;
        RECT 77.780 50.200 77.980 57.800 ;
        RECT 78.580 50.200 78.780 57.800 ;
        RECT 79.530 57.600 83.530 57.800 ;
        RECT 83.130 57.000 83.530 57.600 ;
        RECT 79.530 56.800 83.530 57.000 ;
        RECT 83.130 56.200 83.530 56.800 ;
        RECT 79.530 56.000 83.530 56.200 ;
        RECT 83.130 55.400 83.530 56.000 ;
        RECT 79.530 55.200 83.530 55.400 ;
        RECT 83.130 54.600 83.530 55.200 ;
        RECT 79.530 54.400 83.530 54.600 ;
        RECT 83.130 53.800 83.530 54.400 ;
        RECT 79.530 53.600 83.530 53.800 ;
        RECT 83.130 53.000 83.530 53.600 ;
        RECT 79.530 52.800 83.530 53.000 ;
        RECT 83.130 52.200 83.530 52.800 ;
        RECT 79.530 52.000 83.530 52.200 ;
        RECT 83.130 51.400 83.530 52.000 ;
        RECT 79.530 51.200 83.530 51.400 ;
        RECT 83.130 50.600 83.530 51.200 ;
        RECT 79.530 50.400 83.530 50.600 ;
        RECT 83.130 50.200 83.530 50.400 ;
        RECT 75.380 49.800 83.530 50.200 ;
        RECT 75.380 42.200 75.580 49.800 ;
        RECT 76.180 42.200 76.380 49.800 ;
        RECT 76.980 42.200 77.180 49.800 ;
        RECT 77.780 42.200 77.980 49.800 ;
        RECT 78.580 42.200 78.780 49.800 ;
        RECT 83.130 49.600 83.530 49.800 ;
        RECT 79.530 49.400 83.530 49.600 ;
        RECT 83.130 48.800 83.530 49.400 ;
        RECT 79.530 48.600 83.530 48.800 ;
        RECT 83.130 48.000 83.530 48.600 ;
        RECT 79.530 47.800 83.530 48.000 ;
        RECT 83.130 47.200 83.530 47.800 ;
        RECT 79.530 47.000 83.530 47.200 ;
        RECT 83.130 46.400 83.530 47.000 ;
        RECT 79.530 46.200 83.530 46.400 ;
        RECT 83.130 45.600 83.530 46.200 ;
        RECT 79.530 45.400 83.530 45.600 ;
        RECT 83.130 44.800 83.530 45.400 ;
        RECT 79.530 44.600 83.530 44.800 ;
        RECT 83.130 44.000 83.530 44.600 ;
        RECT 79.530 43.800 83.530 44.000 ;
        RECT 83.130 43.200 83.530 43.800 ;
        RECT 79.530 43.000 83.530 43.200 ;
        RECT 83.130 42.400 83.530 43.000 ;
        RECT 79.530 42.200 83.530 42.400 ;
        RECT 85.930 57.600 89.930 57.800 ;
        RECT 85.930 57.000 86.330 57.600 ;
        RECT 85.930 56.800 89.930 57.000 ;
        RECT 85.930 56.200 86.330 56.800 ;
        RECT 85.930 56.000 89.930 56.200 ;
        RECT 85.930 55.400 86.330 56.000 ;
        RECT 85.930 55.200 89.930 55.400 ;
        RECT 85.930 54.600 86.330 55.200 ;
        RECT 85.930 54.400 89.930 54.600 ;
        RECT 85.930 53.800 86.330 54.400 ;
        RECT 85.930 53.600 89.930 53.800 ;
        RECT 85.930 53.000 86.330 53.600 ;
        RECT 85.930 52.800 89.930 53.000 ;
        RECT 85.930 52.200 86.330 52.800 ;
        RECT 85.930 52.000 89.930 52.200 ;
        RECT 85.930 51.400 86.330 52.000 ;
        RECT 85.930 51.200 89.930 51.400 ;
        RECT 85.930 50.600 86.330 51.200 ;
        RECT 85.930 50.400 89.930 50.600 ;
        RECT 85.930 50.200 86.330 50.400 ;
        RECT 90.680 50.200 90.880 57.800 ;
        RECT 91.480 50.200 91.680 57.800 ;
        RECT 92.280 50.200 92.480 57.800 ;
        RECT 93.080 50.200 93.280 57.800 ;
        RECT 93.880 50.200 94.080 57.800 ;
        RECT 85.930 49.800 94.080 50.200 ;
        RECT 85.930 49.600 86.330 49.800 ;
        RECT 85.930 49.400 89.930 49.600 ;
        RECT 85.930 48.800 86.330 49.400 ;
        RECT 85.930 48.600 89.930 48.800 ;
        RECT 85.930 48.000 86.330 48.600 ;
        RECT 85.930 47.800 89.930 48.000 ;
        RECT 85.930 47.200 86.330 47.800 ;
        RECT 85.930 47.000 89.930 47.200 ;
        RECT 85.930 46.400 86.330 47.000 ;
        RECT 85.930 46.200 89.930 46.400 ;
        RECT 85.930 45.600 86.330 46.200 ;
        RECT 85.930 45.400 89.930 45.600 ;
        RECT 85.930 44.800 86.330 45.400 ;
        RECT 85.930 44.600 89.930 44.800 ;
        RECT 85.930 44.000 86.330 44.600 ;
        RECT 85.930 43.800 89.930 44.000 ;
        RECT 85.930 43.200 86.330 43.800 ;
        RECT 85.930 43.000 89.930 43.200 ;
        RECT 85.930 42.400 86.330 43.000 ;
        RECT 85.930 42.200 89.930 42.400 ;
        RECT 90.680 42.200 90.880 49.800 ;
        RECT 91.480 42.200 91.680 49.800 ;
        RECT 92.280 42.200 92.480 49.800 ;
        RECT 93.080 42.200 93.280 49.800 ;
        RECT 93.880 42.200 94.080 49.800 ;
        RECT 95.380 50.200 95.580 57.800 ;
        RECT 96.180 50.200 96.380 57.800 ;
        RECT 96.980 50.200 97.180 57.800 ;
        RECT 97.780 50.200 97.980 57.800 ;
        RECT 98.580 50.200 98.780 57.800 ;
        RECT 99.530 57.600 103.530 57.800 ;
        RECT 103.130 57.000 103.530 57.600 ;
        RECT 99.530 56.800 103.530 57.000 ;
        RECT 103.130 56.200 103.530 56.800 ;
        RECT 99.530 56.000 103.530 56.200 ;
        RECT 103.130 55.400 103.530 56.000 ;
        RECT 99.530 55.200 103.530 55.400 ;
        RECT 103.130 54.600 103.530 55.200 ;
        RECT 99.530 54.400 103.530 54.600 ;
        RECT 103.130 53.800 103.530 54.400 ;
        RECT 99.530 53.600 103.530 53.800 ;
        RECT 103.130 53.000 103.530 53.600 ;
        RECT 99.530 52.800 103.530 53.000 ;
        RECT 103.130 52.200 103.530 52.800 ;
        RECT 99.530 52.000 103.530 52.200 ;
        RECT 103.130 51.400 103.530 52.000 ;
        RECT 99.530 51.200 103.530 51.400 ;
        RECT 103.130 50.600 103.530 51.200 ;
        RECT 110.050 51.080 110.410 51.460 ;
        RECT 110.680 51.080 111.040 51.460 ;
        RECT 111.280 51.080 111.640 51.460 ;
        RECT 99.530 50.400 103.530 50.600 ;
        RECT 110.050 50.490 110.410 50.870 ;
        RECT 110.680 50.490 111.040 50.870 ;
        RECT 111.280 50.490 111.640 50.870 ;
        RECT 103.130 50.200 103.530 50.400 ;
        RECT 95.380 49.800 103.530 50.200 ;
        RECT 95.380 42.200 95.580 49.800 ;
        RECT 96.180 42.200 96.380 49.800 ;
        RECT 96.980 42.200 97.180 49.800 ;
        RECT 97.780 42.200 97.980 49.800 ;
        RECT 98.580 42.200 98.780 49.800 ;
        RECT 103.130 49.600 103.530 49.800 ;
        RECT 99.530 49.400 103.530 49.600 ;
        RECT 103.130 48.800 103.530 49.400 ;
        RECT 99.530 48.600 103.530 48.800 ;
        RECT 103.130 48.000 103.530 48.600 ;
        RECT 99.530 47.800 103.530 48.000 ;
        RECT 103.130 47.200 103.530 47.800 ;
        RECT 99.530 47.000 103.530 47.200 ;
        RECT 103.130 46.400 103.530 47.000 ;
        RECT 99.530 46.200 103.530 46.400 ;
        RECT 103.130 45.600 103.530 46.200 ;
        RECT 99.530 45.400 103.530 45.600 ;
        RECT 103.130 44.800 103.530 45.400 ;
        RECT 99.530 44.600 103.530 44.800 ;
        RECT 103.130 44.000 103.530 44.600 ;
        RECT 99.530 43.800 103.530 44.000 ;
        RECT 103.130 43.200 103.530 43.800 ;
        RECT 99.530 43.000 103.530 43.200 ;
        RECT 103.130 42.400 103.530 43.000 ;
        RECT 99.530 42.200 103.530 42.400 ;
        RECT 5.930 37.600 9.930 37.800 ;
        RECT 5.930 37.000 6.330 37.600 ;
        RECT 5.930 36.800 9.930 37.000 ;
        RECT 5.930 36.200 6.330 36.800 ;
        RECT 5.930 36.000 9.930 36.200 ;
        RECT 5.930 35.400 6.330 36.000 ;
        RECT 5.930 35.200 9.930 35.400 ;
        RECT 5.930 34.600 6.330 35.200 ;
        RECT 5.930 34.400 9.930 34.600 ;
        RECT 5.930 33.800 6.330 34.400 ;
        RECT 5.930 33.600 9.930 33.800 ;
        RECT 5.930 33.000 6.330 33.600 ;
        RECT 5.930 32.800 9.930 33.000 ;
        RECT 5.930 32.200 6.330 32.800 ;
        RECT 5.930 32.000 9.930 32.200 ;
        RECT 5.930 31.400 6.330 32.000 ;
        RECT 5.930 31.200 9.930 31.400 ;
        RECT 5.930 30.600 6.330 31.200 ;
        RECT 5.930 30.400 9.930 30.600 ;
        RECT 5.930 30.200 6.330 30.400 ;
        RECT 10.680 30.200 10.880 37.800 ;
        RECT 11.480 30.200 11.680 37.800 ;
        RECT 12.280 30.200 12.480 37.800 ;
        RECT 13.080 30.200 13.280 37.800 ;
        RECT 13.880 30.200 14.080 37.800 ;
        RECT 5.930 29.800 14.080 30.200 ;
        RECT 5.930 29.600 6.330 29.800 ;
        RECT 5.930 29.400 9.930 29.600 ;
        RECT 5.930 28.800 6.330 29.400 ;
        RECT 5.930 28.600 9.930 28.800 ;
        RECT 5.930 28.000 6.330 28.600 ;
        RECT 5.930 27.800 9.930 28.000 ;
        RECT 5.930 27.200 6.330 27.800 ;
        RECT 5.930 27.000 9.930 27.200 ;
        RECT 5.930 26.400 6.330 27.000 ;
        RECT 5.930 26.200 9.930 26.400 ;
        RECT 5.930 25.600 6.330 26.200 ;
        RECT 5.930 25.400 9.930 25.600 ;
        RECT 5.930 24.800 6.330 25.400 ;
        RECT 5.930 24.600 9.930 24.800 ;
        RECT 5.930 24.000 6.330 24.600 ;
        RECT 5.930 23.800 9.930 24.000 ;
        RECT 5.930 23.200 6.330 23.800 ;
        RECT 5.930 23.000 9.930 23.200 ;
        RECT 5.930 22.400 6.330 23.000 ;
        RECT 5.930 22.200 9.930 22.400 ;
        RECT 10.680 22.200 10.880 29.800 ;
        RECT 11.480 22.200 11.680 29.800 ;
        RECT 12.280 22.200 12.480 29.800 ;
        RECT 13.080 22.200 13.280 29.800 ;
        RECT 13.880 22.200 14.080 29.800 ;
        RECT 15.380 30.200 15.580 37.800 ;
        RECT 16.180 30.200 16.380 37.800 ;
        RECT 16.980 30.200 17.180 37.800 ;
        RECT 17.780 30.200 17.980 37.800 ;
        RECT 18.580 30.200 18.780 37.800 ;
        RECT 19.530 37.600 23.530 37.800 ;
        RECT 23.130 37.000 23.530 37.600 ;
        RECT 19.530 36.800 23.530 37.000 ;
        RECT 23.130 36.200 23.530 36.800 ;
        RECT 19.530 36.000 23.530 36.200 ;
        RECT 23.130 35.400 23.530 36.000 ;
        RECT 19.530 35.200 23.530 35.400 ;
        RECT 23.130 34.600 23.530 35.200 ;
        RECT 19.530 34.400 23.530 34.600 ;
        RECT 23.130 33.800 23.530 34.400 ;
        RECT 19.530 33.600 23.530 33.800 ;
        RECT 23.130 33.000 23.530 33.600 ;
        RECT 19.530 32.800 23.530 33.000 ;
        RECT 23.130 32.200 23.530 32.800 ;
        RECT 19.530 32.000 23.530 32.200 ;
        RECT 23.130 31.400 23.530 32.000 ;
        RECT 19.530 31.200 23.530 31.400 ;
        RECT 23.130 30.600 23.530 31.200 ;
        RECT 19.530 30.400 23.530 30.600 ;
        RECT 23.130 30.200 23.530 30.400 ;
        RECT 15.380 29.800 23.530 30.200 ;
        RECT 15.380 22.200 15.580 29.800 ;
        RECT 16.180 22.200 16.380 29.800 ;
        RECT 16.980 22.200 17.180 29.800 ;
        RECT 17.780 22.200 17.980 29.800 ;
        RECT 18.580 22.200 18.780 29.800 ;
        RECT 23.130 29.600 23.530 29.800 ;
        RECT 19.530 29.400 23.530 29.600 ;
        RECT 23.130 28.800 23.530 29.400 ;
        RECT 19.530 28.600 23.530 28.800 ;
        RECT 23.130 28.000 23.530 28.600 ;
        RECT 19.530 27.800 23.530 28.000 ;
        RECT 23.130 27.200 23.530 27.800 ;
        RECT 19.530 27.000 23.530 27.200 ;
        RECT 23.130 26.400 23.530 27.000 ;
        RECT 19.530 26.200 23.530 26.400 ;
        RECT 23.130 25.600 23.530 26.200 ;
        RECT 19.530 25.400 23.530 25.600 ;
        RECT 23.130 24.800 23.530 25.400 ;
        RECT 19.530 24.600 23.530 24.800 ;
        RECT 23.130 24.000 23.530 24.600 ;
        RECT 19.530 23.800 23.530 24.000 ;
        RECT 23.130 23.200 23.530 23.800 ;
        RECT 19.530 23.000 23.530 23.200 ;
        RECT 23.130 22.400 23.530 23.000 ;
        RECT 19.530 22.200 23.530 22.400 ;
        RECT 25.930 37.600 29.930 37.800 ;
        RECT 25.930 37.000 26.330 37.600 ;
        RECT 25.930 36.800 29.930 37.000 ;
        RECT 25.930 36.200 26.330 36.800 ;
        RECT 25.930 36.000 29.930 36.200 ;
        RECT 25.930 35.400 26.330 36.000 ;
        RECT 25.930 35.200 29.930 35.400 ;
        RECT 25.930 34.600 26.330 35.200 ;
        RECT 25.930 34.400 29.930 34.600 ;
        RECT 25.930 33.800 26.330 34.400 ;
        RECT 25.930 33.600 29.930 33.800 ;
        RECT 25.930 33.000 26.330 33.600 ;
        RECT 25.930 32.800 29.930 33.000 ;
        RECT 25.930 32.200 26.330 32.800 ;
        RECT 25.930 32.000 29.930 32.200 ;
        RECT 25.930 31.400 26.330 32.000 ;
        RECT 25.930 31.200 29.930 31.400 ;
        RECT 25.930 30.600 26.330 31.200 ;
        RECT 25.930 30.400 29.930 30.600 ;
        RECT 25.930 30.200 26.330 30.400 ;
        RECT 30.680 30.200 30.880 37.800 ;
        RECT 31.480 30.200 31.680 37.800 ;
        RECT 32.280 30.200 32.480 37.800 ;
        RECT 33.080 30.200 33.280 37.800 ;
        RECT 33.880 30.200 34.080 37.800 ;
        RECT 25.930 29.800 34.080 30.200 ;
        RECT 25.930 29.600 26.330 29.800 ;
        RECT 25.930 29.400 29.930 29.600 ;
        RECT 25.930 28.800 26.330 29.400 ;
        RECT 25.930 28.600 29.930 28.800 ;
        RECT 25.930 28.000 26.330 28.600 ;
        RECT 25.930 27.800 29.930 28.000 ;
        RECT 25.930 27.200 26.330 27.800 ;
        RECT 25.930 27.000 29.930 27.200 ;
        RECT 25.930 26.400 26.330 27.000 ;
        RECT 25.930 26.200 29.930 26.400 ;
        RECT 25.930 25.600 26.330 26.200 ;
        RECT 25.930 25.400 29.930 25.600 ;
        RECT 25.930 24.800 26.330 25.400 ;
        RECT 25.930 24.600 29.930 24.800 ;
        RECT 25.930 24.000 26.330 24.600 ;
        RECT 25.930 23.800 29.930 24.000 ;
        RECT 25.930 23.200 26.330 23.800 ;
        RECT 25.930 23.000 29.930 23.200 ;
        RECT 25.930 22.400 26.330 23.000 ;
        RECT 25.930 22.200 29.930 22.400 ;
        RECT 30.680 22.200 30.880 29.800 ;
        RECT 31.480 22.200 31.680 29.800 ;
        RECT 32.280 22.200 32.480 29.800 ;
        RECT 33.080 22.200 33.280 29.800 ;
        RECT 33.880 22.200 34.080 29.800 ;
        RECT 35.380 30.200 35.580 37.800 ;
        RECT 36.180 30.200 36.380 37.800 ;
        RECT 36.980 30.200 37.180 37.800 ;
        RECT 37.780 30.200 37.980 37.800 ;
        RECT 38.580 30.200 38.780 37.800 ;
        RECT 39.530 37.600 43.530 37.800 ;
        RECT 43.130 37.000 43.530 37.600 ;
        RECT 39.530 36.800 43.530 37.000 ;
        RECT 43.130 36.200 43.530 36.800 ;
        RECT 39.530 36.000 43.530 36.200 ;
        RECT 43.130 35.400 43.530 36.000 ;
        RECT 39.530 35.200 43.530 35.400 ;
        RECT 43.130 34.600 43.530 35.200 ;
        RECT 39.530 34.400 43.530 34.600 ;
        RECT 43.130 33.800 43.530 34.400 ;
        RECT 39.530 33.600 43.530 33.800 ;
        RECT 43.130 33.000 43.530 33.600 ;
        RECT 39.530 32.800 43.530 33.000 ;
        RECT 43.130 32.200 43.530 32.800 ;
        RECT 39.530 32.000 43.530 32.200 ;
        RECT 43.130 31.400 43.530 32.000 ;
        RECT 39.530 31.200 43.530 31.400 ;
        RECT 43.130 30.600 43.530 31.200 ;
        RECT 39.530 30.400 43.530 30.600 ;
        RECT 43.130 30.200 43.530 30.400 ;
        RECT 35.380 29.800 43.530 30.200 ;
        RECT 35.380 22.200 35.580 29.800 ;
        RECT 36.180 22.200 36.380 29.800 ;
        RECT 36.980 22.200 37.180 29.800 ;
        RECT 37.780 22.200 37.980 29.800 ;
        RECT 38.580 22.200 38.780 29.800 ;
        RECT 43.130 29.600 43.530 29.800 ;
        RECT 39.530 29.400 43.530 29.600 ;
        RECT 43.130 28.800 43.530 29.400 ;
        RECT 39.530 28.600 43.530 28.800 ;
        RECT 43.130 28.000 43.530 28.600 ;
        RECT 39.530 27.800 43.530 28.000 ;
        RECT 43.130 27.200 43.530 27.800 ;
        RECT 39.530 27.000 43.530 27.200 ;
        RECT 43.130 26.400 43.530 27.000 ;
        RECT 39.530 26.200 43.530 26.400 ;
        RECT 43.130 25.600 43.530 26.200 ;
        RECT 39.530 25.400 43.530 25.600 ;
        RECT 43.130 24.800 43.530 25.400 ;
        RECT 39.530 24.600 43.530 24.800 ;
        RECT 43.130 24.000 43.530 24.600 ;
        RECT 39.530 23.800 43.530 24.000 ;
        RECT 43.130 23.200 43.530 23.800 ;
        RECT 39.530 23.000 43.530 23.200 ;
        RECT 43.130 22.400 43.530 23.000 ;
        RECT 39.530 22.200 43.530 22.400 ;
        RECT 45.930 37.600 49.930 37.800 ;
        RECT 45.930 37.000 46.330 37.600 ;
        RECT 45.930 36.800 49.930 37.000 ;
        RECT 45.930 36.200 46.330 36.800 ;
        RECT 45.930 36.000 49.930 36.200 ;
        RECT 45.930 35.400 46.330 36.000 ;
        RECT 45.930 35.200 49.930 35.400 ;
        RECT 45.930 34.600 46.330 35.200 ;
        RECT 45.930 34.400 49.930 34.600 ;
        RECT 45.930 33.800 46.330 34.400 ;
        RECT 45.930 33.600 49.930 33.800 ;
        RECT 45.930 33.000 46.330 33.600 ;
        RECT 45.930 32.800 49.930 33.000 ;
        RECT 45.930 32.200 46.330 32.800 ;
        RECT 45.930 32.000 49.930 32.200 ;
        RECT 45.930 31.400 46.330 32.000 ;
        RECT 45.930 31.200 49.930 31.400 ;
        RECT 45.930 30.600 46.330 31.200 ;
        RECT 45.930 30.400 49.930 30.600 ;
        RECT 45.930 30.200 46.330 30.400 ;
        RECT 50.680 30.200 50.880 37.800 ;
        RECT 51.480 30.200 51.680 37.800 ;
        RECT 52.280 30.200 52.480 37.800 ;
        RECT 53.080 30.200 53.280 37.800 ;
        RECT 53.880 30.200 54.080 37.800 ;
        RECT 45.930 29.800 54.080 30.200 ;
        RECT 45.930 29.600 46.330 29.800 ;
        RECT 45.930 29.400 49.930 29.600 ;
        RECT 45.930 28.800 46.330 29.400 ;
        RECT 45.930 28.600 49.930 28.800 ;
        RECT 45.930 28.000 46.330 28.600 ;
        RECT 45.930 27.800 49.930 28.000 ;
        RECT 45.930 27.200 46.330 27.800 ;
        RECT 45.930 27.000 49.930 27.200 ;
        RECT 45.930 26.400 46.330 27.000 ;
        RECT 45.930 26.200 49.930 26.400 ;
        RECT 45.930 25.600 46.330 26.200 ;
        RECT 45.930 25.400 49.930 25.600 ;
        RECT 45.930 24.800 46.330 25.400 ;
        RECT 45.930 24.600 49.930 24.800 ;
        RECT 45.930 24.000 46.330 24.600 ;
        RECT 45.930 23.800 49.930 24.000 ;
        RECT 45.930 23.200 46.330 23.800 ;
        RECT 45.930 23.000 49.930 23.200 ;
        RECT 45.930 22.400 46.330 23.000 ;
        RECT 45.930 22.200 49.930 22.400 ;
        RECT 50.680 22.200 50.880 29.800 ;
        RECT 51.480 22.200 51.680 29.800 ;
        RECT 52.280 22.200 52.480 29.800 ;
        RECT 53.080 22.200 53.280 29.800 ;
        RECT 53.880 22.200 54.080 29.800 ;
        RECT 55.380 30.200 55.580 37.800 ;
        RECT 56.180 30.200 56.380 37.800 ;
        RECT 56.980 30.200 57.180 37.800 ;
        RECT 57.780 30.200 57.980 37.800 ;
        RECT 58.580 30.200 58.780 37.800 ;
        RECT 59.530 37.600 63.530 37.800 ;
        RECT 63.130 37.000 63.530 37.600 ;
        RECT 59.530 36.800 63.530 37.000 ;
        RECT 63.130 36.200 63.530 36.800 ;
        RECT 59.530 36.000 63.530 36.200 ;
        RECT 63.130 35.400 63.530 36.000 ;
        RECT 59.530 35.200 63.530 35.400 ;
        RECT 63.130 34.600 63.530 35.200 ;
        RECT 59.530 34.400 63.530 34.600 ;
        RECT 63.130 33.800 63.530 34.400 ;
        RECT 59.530 33.600 63.530 33.800 ;
        RECT 63.130 33.000 63.530 33.600 ;
        RECT 59.530 32.800 63.530 33.000 ;
        RECT 63.130 32.200 63.530 32.800 ;
        RECT 59.530 32.000 63.530 32.200 ;
        RECT 63.130 31.400 63.530 32.000 ;
        RECT 59.530 31.200 63.530 31.400 ;
        RECT 63.130 30.600 63.530 31.200 ;
        RECT 59.530 30.400 63.530 30.600 ;
        RECT 63.130 30.200 63.530 30.400 ;
        RECT 55.380 29.800 63.530 30.200 ;
        RECT 55.380 22.200 55.580 29.800 ;
        RECT 56.180 22.200 56.380 29.800 ;
        RECT 56.980 22.200 57.180 29.800 ;
        RECT 57.780 22.200 57.980 29.800 ;
        RECT 58.580 22.200 58.780 29.800 ;
        RECT 63.130 29.600 63.530 29.800 ;
        RECT 59.530 29.400 63.530 29.600 ;
        RECT 63.130 28.800 63.530 29.400 ;
        RECT 59.530 28.600 63.530 28.800 ;
        RECT 63.130 28.000 63.530 28.600 ;
        RECT 59.530 27.800 63.530 28.000 ;
        RECT 63.130 27.200 63.530 27.800 ;
        RECT 59.530 27.000 63.530 27.200 ;
        RECT 63.130 26.400 63.530 27.000 ;
        RECT 59.530 26.200 63.530 26.400 ;
        RECT 63.130 25.600 63.530 26.200 ;
        RECT 59.530 25.400 63.530 25.600 ;
        RECT 63.130 24.800 63.530 25.400 ;
        RECT 59.530 24.600 63.530 24.800 ;
        RECT 63.130 24.000 63.530 24.600 ;
        RECT 59.530 23.800 63.530 24.000 ;
        RECT 63.130 23.200 63.530 23.800 ;
        RECT 59.530 23.000 63.530 23.200 ;
        RECT 63.130 22.400 63.530 23.000 ;
        RECT 59.530 22.200 63.530 22.400 ;
        RECT 65.930 37.600 69.930 37.800 ;
        RECT 65.930 37.000 66.330 37.600 ;
        RECT 65.930 36.800 69.930 37.000 ;
        RECT 65.930 36.200 66.330 36.800 ;
        RECT 65.930 36.000 69.930 36.200 ;
        RECT 65.930 35.400 66.330 36.000 ;
        RECT 65.930 35.200 69.930 35.400 ;
        RECT 65.930 34.600 66.330 35.200 ;
        RECT 65.930 34.400 69.930 34.600 ;
        RECT 65.930 33.800 66.330 34.400 ;
        RECT 65.930 33.600 69.930 33.800 ;
        RECT 65.930 33.000 66.330 33.600 ;
        RECT 65.930 32.800 69.930 33.000 ;
        RECT 65.930 32.200 66.330 32.800 ;
        RECT 65.930 32.000 69.930 32.200 ;
        RECT 65.930 31.400 66.330 32.000 ;
        RECT 65.930 31.200 69.930 31.400 ;
        RECT 65.930 30.600 66.330 31.200 ;
        RECT 65.930 30.400 69.930 30.600 ;
        RECT 65.930 30.200 66.330 30.400 ;
        RECT 70.680 30.200 70.880 37.800 ;
        RECT 71.480 30.200 71.680 37.800 ;
        RECT 72.280 30.200 72.480 37.800 ;
        RECT 73.080 30.200 73.280 37.800 ;
        RECT 73.880 30.200 74.080 37.800 ;
        RECT 65.930 29.800 74.080 30.200 ;
        RECT 65.930 29.600 66.330 29.800 ;
        RECT 65.930 29.400 69.930 29.600 ;
        RECT 65.930 28.800 66.330 29.400 ;
        RECT 65.930 28.600 69.930 28.800 ;
        RECT 65.930 28.000 66.330 28.600 ;
        RECT 65.930 27.800 69.930 28.000 ;
        RECT 65.930 27.200 66.330 27.800 ;
        RECT 65.930 27.000 69.930 27.200 ;
        RECT 65.930 26.400 66.330 27.000 ;
        RECT 65.930 26.200 69.930 26.400 ;
        RECT 65.930 25.600 66.330 26.200 ;
        RECT 65.930 25.400 69.930 25.600 ;
        RECT 65.930 24.800 66.330 25.400 ;
        RECT 65.930 24.600 69.930 24.800 ;
        RECT 65.930 24.000 66.330 24.600 ;
        RECT 65.930 23.800 69.930 24.000 ;
        RECT 65.930 23.200 66.330 23.800 ;
        RECT 65.930 23.000 69.930 23.200 ;
        RECT 65.930 22.400 66.330 23.000 ;
        RECT 65.930 22.200 69.930 22.400 ;
        RECT 70.680 22.200 70.880 29.800 ;
        RECT 71.480 22.200 71.680 29.800 ;
        RECT 72.280 22.200 72.480 29.800 ;
        RECT 73.080 22.200 73.280 29.800 ;
        RECT 73.880 22.200 74.080 29.800 ;
        RECT 75.380 30.200 75.580 37.800 ;
        RECT 76.180 30.200 76.380 37.800 ;
        RECT 76.980 30.200 77.180 37.800 ;
        RECT 77.780 30.200 77.980 37.800 ;
        RECT 78.580 30.200 78.780 37.800 ;
        RECT 79.530 37.600 83.530 37.800 ;
        RECT 83.130 37.000 83.530 37.600 ;
        RECT 79.530 36.800 83.530 37.000 ;
        RECT 83.130 36.200 83.530 36.800 ;
        RECT 79.530 36.000 83.530 36.200 ;
        RECT 83.130 35.400 83.530 36.000 ;
        RECT 79.530 35.200 83.530 35.400 ;
        RECT 83.130 34.600 83.530 35.200 ;
        RECT 79.530 34.400 83.530 34.600 ;
        RECT 83.130 33.800 83.530 34.400 ;
        RECT 79.530 33.600 83.530 33.800 ;
        RECT 83.130 33.000 83.530 33.600 ;
        RECT 79.530 32.800 83.530 33.000 ;
        RECT 83.130 32.200 83.530 32.800 ;
        RECT 79.530 32.000 83.530 32.200 ;
        RECT 83.130 31.400 83.530 32.000 ;
        RECT 79.530 31.200 83.530 31.400 ;
        RECT 83.130 30.600 83.530 31.200 ;
        RECT 79.530 30.400 83.530 30.600 ;
        RECT 83.130 30.200 83.530 30.400 ;
        RECT 75.380 29.800 83.530 30.200 ;
        RECT 75.380 22.200 75.580 29.800 ;
        RECT 76.180 22.200 76.380 29.800 ;
        RECT 76.980 22.200 77.180 29.800 ;
        RECT 77.780 22.200 77.980 29.800 ;
        RECT 78.580 22.200 78.780 29.800 ;
        RECT 83.130 29.600 83.530 29.800 ;
        RECT 79.530 29.400 83.530 29.600 ;
        RECT 83.130 28.800 83.530 29.400 ;
        RECT 79.530 28.600 83.530 28.800 ;
        RECT 83.130 28.000 83.530 28.600 ;
        RECT 79.530 27.800 83.530 28.000 ;
        RECT 83.130 27.200 83.530 27.800 ;
        RECT 79.530 27.000 83.530 27.200 ;
        RECT 83.130 26.400 83.530 27.000 ;
        RECT 79.530 26.200 83.530 26.400 ;
        RECT 83.130 25.600 83.530 26.200 ;
        RECT 79.530 25.400 83.530 25.600 ;
        RECT 83.130 24.800 83.530 25.400 ;
        RECT 79.530 24.600 83.530 24.800 ;
        RECT 83.130 24.000 83.530 24.600 ;
        RECT 79.530 23.800 83.530 24.000 ;
        RECT 83.130 23.200 83.530 23.800 ;
        RECT 79.530 23.000 83.530 23.200 ;
        RECT 83.130 22.400 83.530 23.000 ;
        RECT 79.530 22.200 83.530 22.400 ;
        RECT 85.930 37.600 89.930 37.800 ;
        RECT 85.930 37.000 86.330 37.600 ;
        RECT 85.930 36.800 89.930 37.000 ;
        RECT 85.930 36.200 86.330 36.800 ;
        RECT 85.930 36.000 89.930 36.200 ;
        RECT 85.930 35.400 86.330 36.000 ;
        RECT 85.930 35.200 89.930 35.400 ;
        RECT 85.930 34.600 86.330 35.200 ;
        RECT 85.930 34.400 89.930 34.600 ;
        RECT 85.930 33.800 86.330 34.400 ;
        RECT 85.930 33.600 89.930 33.800 ;
        RECT 85.930 33.000 86.330 33.600 ;
        RECT 85.930 32.800 89.930 33.000 ;
        RECT 85.930 32.200 86.330 32.800 ;
        RECT 85.930 32.000 89.930 32.200 ;
        RECT 85.930 31.400 86.330 32.000 ;
        RECT 85.930 31.200 89.930 31.400 ;
        RECT 85.930 30.600 86.330 31.200 ;
        RECT 85.930 30.400 89.930 30.600 ;
        RECT 85.930 30.200 86.330 30.400 ;
        RECT 90.680 30.200 90.880 37.800 ;
        RECT 91.480 30.200 91.680 37.800 ;
        RECT 92.280 30.200 92.480 37.800 ;
        RECT 93.080 30.200 93.280 37.800 ;
        RECT 93.880 30.200 94.080 37.800 ;
        RECT 85.930 29.800 94.080 30.200 ;
        RECT 85.930 29.600 86.330 29.800 ;
        RECT 85.930 29.400 89.930 29.600 ;
        RECT 85.930 28.800 86.330 29.400 ;
        RECT 85.930 28.600 89.930 28.800 ;
        RECT 85.930 28.000 86.330 28.600 ;
        RECT 85.930 27.800 89.930 28.000 ;
        RECT 85.930 27.200 86.330 27.800 ;
        RECT 85.930 27.000 89.930 27.200 ;
        RECT 85.930 26.400 86.330 27.000 ;
        RECT 85.930 26.200 89.930 26.400 ;
        RECT 85.930 25.600 86.330 26.200 ;
        RECT 85.930 25.400 89.930 25.600 ;
        RECT 85.930 24.800 86.330 25.400 ;
        RECT 85.930 24.600 89.930 24.800 ;
        RECT 85.930 24.000 86.330 24.600 ;
        RECT 85.930 23.800 89.930 24.000 ;
        RECT 85.930 23.200 86.330 23.800 ;
        RECT 85.930 23.000 89.930 23.200 ;
        RECT 85.930 22.400 86.330 23.000 ;
        RECT 85.930 22.200 89.930 22.400 ;
        RECT 90.680 22.200 90.880 29.800 ;
        RECT 91.480 22.200 91.680 29.800 ;
        RECT 92.280 22.200 92.480 29.800 ;
        RECT 93.080 22.200 93.280 29.800 ;
        RECT 93.880 22.200 94.080 29.800 ;
        RECT 95.380 30.200 95.580 37.800 ;
        RECT 96.180 30.200 96.380 37.800 ;
        RECT 96.980 30.200 97.180 37.800 ;
        RECT 97.780 30.200 97.980 37.800 ;
        RECT 98.580 30.200 98.780 37.800 ;
        RECT 99.530 37.600 103.530 37.800 ;
        RECT 103.130 37.000 103.530 37.600 ;
        RECT 99.530 36.800 103.530 37.000 ;
        RECT 103.130 36.200 103.530 36.800 ;
        RECT 99.530 36.000 103.530 36.200 ;
        RECT 103.130 35.400 103.530 36.000 ;
        RECT 99.530 35.200 103.530 35.400 ;
        RECT 103.130 34.600 103.530 35.200 ;
        RECT 99.530 34.400 103.530 34.600 ;
        RECT 103.130 33.800 103.530 34.400 ;
        RECT 99.530 33.600 103.530 33.800 ;
        RECT 103.130 33.000 103.530 33.600 ;
        RECT 99.530 32.800 103.530 33.000 ;
        RECT 103.130 32.200 103.530 32.800 ;
        RECT 99.530 32.000 103.530 32.200 ;
        RECT 103.130 31.400 103.530 32.000 ;
        RECT 99.530 31.200 103.530 31.400 ;
        RECT 103.130 30.600 103.530 31.200 ;
        RECT 110.050 31.020 110.410 31.400 ;
        RECT 110.680 31.020 111.040 31.400 ;
        RECT 111.280 31.020 111.640 31.400 ;
        RECT 99.530 30.400 103.530 30.600 ;
        RECT 110.050 30.430 110.410 30.810 ;
        RECT 110.680 30.430 111.040 30.810 ;
        RECT 111.280 30.430 111.640 30.810 ;
        RECT 103.130 30.200 103.530 30.400 ;
        RECT 95.380 29.800 103.530 30.200 ;
        RECT 95.380 22.200 95.580 29.800 ;
        RECT 96.180 22.200 96.380 29.800 ;
        RECT 96.980 22.200 97.180 29.800 ;
        RECT 97.780 22.200 97.980 29.800 ;
        RECT 98.580 22.200 98.780 29.800 ;
        RECT 103.130 29.600 103.530 29.800 ;
        RECT 99.530 29.400 103.530 29.600 ;
        RECT 103.130 28.800 103.530 29.400 ;
        RECT 99.530 28.600 103.530 28.800 ;
        RECT 103.130 28.000 103.530 28.600 ;
        RECT 99.530 27.800 103.530 28.000 ;
        RECT 103.130 27.200 103.530 27.800 ;
        RECT 99.530 27.000 103.530 27.200 ;
        RECT 103.130 26.400 103.530 27.000 ;
        RECT 99.530 26.200 103.530 26.400 ;
        RECT 103.130 25.600 103.530 26.200 ;
        RECT 99.530 25.400 103.530 25.600 ;
        RECT 103.130 24.800 103.530 25.400 ;
        RECT 99.530 24.600 103.530 24.800 ;
        RECT 103.130 24.000 103.530 24.600 ;
        RECT 99.530 23.800 103.530 24.000 ;
        RECT 103.130 23.200 103.530 23.800 ;
        RECT 99.530 23.000 103.530 23.200 ;
        RECT 103.130 22.400 103.530 23.000 ;
        RECT 99.530 22.200 103.530 22.400 ;
        RECT 5.930 17.600 9.930 17.800 ;
        RECT 5.930 17.000 6.330 17.600 ;
        RECT 5.930 16.800 9.930 17.000 ;
        RECT 5.930 16.200 6.330 16.800 ;
        RECT 5.930 16.000 9.930 16.200 ;
        RECT 5.930 15.400 6.330 16.000 ;
        RECT 5.930 15.200 9.930 15.400 ;
        RECT 5.930 14.600 6.330 15.200 ;
        RECT 5.930 14.400 9.930 14.600 ;
        RECT 5.930 13.800 6.330 14.400 ;
        RECT 5.930 13.600 9.930 13.800 ;
        RECT 5.930 13.000 6.330 13.600 ;
        RECT 5.930 12.800 9.930 13.000 ;
        RECT 5.930 12.200 6.330 12.800 ;
        RECT 5.930 12.000 9.930 12.200 ;
        RECT 5.930 11.400 6.330 12.000 ;
        RECT 5.930 11.200 9.930 11.400 ;
        RECT 5.930 10.600 6.330 11.200 ;
        RECT 5.930 10.400 9.930 10.600 ;
        RECT 5.930 10.200 6.330 10.400 ;
        RECT 10.680 10.200 10.880 17.800 ;
        RECT 11.480 10.200 11.680 17.800 ;
        RECT 12.280 10.200 12.480 17.800 ;
        RECT 13.080 10.200 13.280 17.800 ;
        RECT 13.880 10.200 14.080 17.800 ;
        RECT 5.930 9.800 14.080 10.200 ;
        RECT 5.930 9.600 6.330 9.800 ;
        RECT 5.930 9.400 9.930 9.600 ;
        RECT 5.930 8.800 6.330 9.400 ;
        RECT 5.930 8.600 9.930 8.800 ;
        RECT 5.930 8.000 6.330 8.600 ;
        RECT 5.930 7.800 9.930 8.000 ;
        RECT 5.930 7.200 6.330 7.800 ;
        RECT 5.930 7.000 9.930 7.200 ;
        RECT 5.930 6.400 6.330 7.000 ;
        RECT 5.930 6.200 9.930 6.400 ;
        RECT 5.930 5.600 6.330 6.200 ;
        RECT 5.930 5.400 9.930 5.600 ;
        RECT 5.930 4.800 6.330 5.400 ;
        RECT 5.930 4.600 9.930 4.800 ;
        RECT 5.930 4.000 6.330 4.600 ;
        RECT 5.930 3.800 9.930 4.000 ;
        RECT 5.930 3.200 6.330 3.800 ;
        RECT 5.930 3.000 9.930 3.200 ;
        RECT 5.930 2.400 6.330 3.000 ;
        RECT 5.930 2.200 9.930 2.400 ;
        RECT 10.680 2.200 10.880 9.800 ;
        RECT 11.480 2.200 11.680 9.800 ;
        RECT 12.280 2.200 12.480 9.800 ;
        RECT 13.080 2.200 13.280 9.800 ;
        RECT 13.880 2.200 14.080 9.800 ;
        RECT 15.380 10.200 15.580 17.800 ;
        RECT 16.180 10.200 16.380 17.800 ;
        RECT 16.980 10.200 17.180 17.800 ;
        RECT 17.780 10.200 17.980 17.800 ;
        RECT 18.580 10.200 18.780 17.800 ;
        RECT 19.530 17.600 23.530 17.800 ;
        RECT 23.130 17.000 23.530 17.600 ;
        RECT 19.530 16.800 23.530 17.000 ;
        RECT 23.130 16.200 23.530 16.800 ;
        RECT 19.530 16.000 23.530 16.200 ;
        RECT 23.130 15.400 23.530 16.000 ;
        RECT 19.530 15.200 23.530 15.400 ;
        RECT 23.130 14.600 23.530 15.200 ;
        RECT 19.530 14.400 23.530 14.600 ;
        RECT 23.130 13.800 23.530 14.400 ;
        RECT 19.530 13.600 23.530 13.800 ;
        RECT 23.130 13.000 23.530 13.600 ;
        RECT 19.530 12.800 23.530 13.000 ;
        RECT 23.130 12.200 23.530 12.800 ;
        RECT 19.530 12.000 23.530 12.200 ;
        RECT 23.130 11.400 23.530 12.000 ;
        RECT 19.530 11.200 23.530 11.400 ;
        RECT 23.130 10.600 23.530 11.200 ;
        RECT 19.530 10.400 23.530 10.600 ;
        RECT 23.130 10.200 23.530 10.400 ;
        RECT 15.380 9.800 23.530 10.200 ;
        RECT 15.380 2.200 15.580 9.800 ;
        RECT 16.180 2.200 16.380 9.800 ;
        RECT 16.980 2.200 17.180 9.800 ;
        RECT 17.780 2.200 17.980 9.800 ;
        RECT 18.580 2.200 18.780 9.800 ;
        RECT 23.130 9.600 23.530 9.800 ;
        RECT 19.530 9.400 23.530 9.600 ;
        RECT 23.130 8.800 23.530 9.400 ;
        RECT 19.530 8.600 23.530 8.800 ;
        RECT 23.130 8.000 23.530 8.600 ;
        RECT 19.530 7.800 23.530 8.000 ;
        RECT 23.130 7.200 23.530 7.800 ;
        RECT 19.530 7.000 23.530 7.200 ;
        RECT 23.130 6.400 23.530 7.000 ;
        RECT 19.530 6.200 23.530 6.400 ;
        RECT 23.130 5.600 23.530 6.200 ;
        RECT 19.530 5.400 23.530 5.600 ;
        RECT 23.130 4.800 23.530 5.400 ;
        RECT 19.530 4.600 23.530 4.800 ;
        RECT 23.130 4.000 23.530 4.600 ;
        RECT 19.530 3.800 23.530 4.000 ;
        RECT 23.130 3.200 23.530 3.800 ;
        RECT 19.530 3.000 23.530 3.200 ;
        RECT 23.130 2.400 23.530 3.000 ;
        RECT 19.530 2.200 23.530 2.400 ;
        RECT 25.930 17.600 29.930 17.800 ;
        RECT 25.930 17.000 26.330 17.600 ;
        RECT 25.930 16.800 29.930 17.000 ;
        RECT 25.930 16.200 26.330 16.800 ;
        RECT 25.930 16.000 29.930 16.200 ;
        RECT 25.930 15.400 26.330 16.000 ;
        RECT 25.930 15.200 29.930 15.400 ;
        RECT 25.930 14.600 26.330 15.200 ;
        RECT 25.930 14.400 29.930 14.600 ;
        RECT 25.930 13.800 26.330 14.400 ;
        RECT 25.930 13.600 29.930 13.800 ;
        RECT 25.930 13.000 26.330 13.600 ;
        RECT 25.930 12.800 29.930 13.000 ;
        RECT 25.930 12.200 26.330 12.800 ;
        RECT 25.930 12.000 29.930 12.200 ;
        RECT 25.930 11.400 26.330 12.000 ;
        RECT 25.930 11.200 29.930 11.400 ;
        RECT 25.930 10.600 26.330 11.200 ;
        RECT 25.930 10.400 29.930 10.600 ;
        RECT 25.930 10.200 26.330 10.400 ;
        RECT 30.680 10.200 30.880 17.800 ;
        RECT 31.480 10.200 31.680 17.800 ;
        RECT 32.280 10.200 32.480 17.800 ;
        RECT 33.080 10.200 33.280 17.800 ;
        RECT 33.880 10.200 34.080 17.800 ;
        RECT 25.930 9.800 34.080 10.200 ;
        RECT 25.930 9.600 26.330 9.800 ;
        RECT 25.930 9.400 29.930 9.600 ;
        RECT 25.930 8.800 26.330 9.400 ;
        RECT 25.930 8.600 29.930 8.800 ;
        RECT 25.930 8.000 26.330 8.600 ;
        RECT 25.930 7.800 29.930 8.000 ;
        RECT 25.930 7.200 26.330 7.800 ;
        RECT 25.930 7.000 29.930 7.200 ;
        RECT 25.930 6.400 26.330 7.000 ;
        RECT 25.930 6.200 29.930 6.400 ;
        RECT 25.930 5.600 26.330 6.200 ;
        RECT 25.930 5.400 29.930 5.600 ;
        RECT 25.930 4.800 26.330 5.400 ;
        RECT 25.930 4.600 29.930 4.800 ;
        RECT 25.930 4.000 26.330 4.600 ;
        RECT 25.930 3.800 29.930 4.000 ;
        RECT 25.930 3.200 26.330 3.800 ;
        RECT 25.930 3.000 29.930 3.200 ;
        RECT 25.930 2.400 26.330 3.000 ;
        RECT 25.930 2.200 29.930 2.400 ;
        RECT 30.680 2.200 30.880 9.800 ;
        RECT 31.480 2.200 31.680 9.800 ;
        RECT 32.280 2.200 32.480 9.800 ;
        RECT 33.080 2.200 33.280 9.800 ;
        RECT 33.880 2.200 34.080 9.800 ;
        RECT 35.380 10.200 35.580 17.800 ;
        RECT 36.180 10.200 36.380 17.800 ;
        RECT 36.980 10.200 37.180 17.800 ;
        RECT 37.780 10.200 37.980 17.800 ;
        RECT 38.580 10.200 38.780 17.800 ;
        RECT 39.530 17.600 43.530 17.800 ;
        RECT 43.130 17.000 43.530 17.600 ;
        RECT 39.530 16.800 43.530 17.000 ;
        RECT 43.130 16.200 43.530 16.800 ;
        RECT 39.530 16.000 43.530 16.200 ;
        RECT 43.130 15.400 43.530 16.000 ;
        RECT 39.530 15.200 43.530 15.400 ;
        RECT 43.130 14.600 43.530 15.200 ;
        RECT 39.530 14.400 43.530 14.600 ;
        RECT 43.130 13.800 43.530 14.400 ;
        RECT 39.530 13.600 43.530 13.800 ;
        RECT 43.130 13.000 43.530 13.600 ;
        RECT 39.530 12.800 43.530 13.000 ;
        RECT 43.130 12.200 43.530 12.800 ;
        RECT 39.530 12.000 43.530 12.200 ;
        RECT 43.130 11.400 43.530 12.000 ;
        RECT 39.530 11.200 43.530 11.400 ;
        RECT 43.130 10.600 43.530 11.200 ;
        RECT 39.530 10.400 43.530 10.600 ;
        RECT 43.130 10.200 43.530 10.400 ;
        RECT 35.380 9.800 43.530 10.200 ;
        RECT 35.380 2.200 35.580 9.800 ;
        RECT 36.180 2.200 36.380 9.800 ;
        RECT 36.980 2.200 37.180 9.800 ;
        RECT 37.780 2.200 37.980 9.800 ;
        RECT 38.580 2.200 38.780 9.800 ;
        RECT 43.130 9.600 43.530 9.800 ;
        RECT 39.530 9.400 43.530 9.600 ;
        RECT 43.130 8.800 43.530 9.400 ;
        RECT 39.530 8.600 43.530 8.800 ;
        RECT 43.130 8.000 43.530 8.600 ;
        RECT 39.530 7.800 43.530 8.000 ;
        RECT 43.130 7.200 43.530 7.800 ;
        RECT 39.530 7.000 43.530 7.200 ;
        RECT 43.130 6.400 43.530 7.000 ;
        RECT 39.530 6.200 43.530 6.400 ;
        RECT 43.130 5.600 43.530 6.200 ;
        RECT 39.530 5.400 43.530 5.600 ;
        RECT 43.130 4.800 43.530 5.400 ;
        RECT 39.530 4.600 43.530 4.800 ;
        RECT 43.130 4.000 43.530 4.600 ;
        RECT 39.530 3.800 43.530 4.000 ;
        RECT 43.130 3.200 43.530 3.800 ;
        RECT 39.530 3.000 43.530 3.200 ;
        RECT 43.130 2.400 43.530 3.000 ;
        RECT 39.530 2.200 43.530 2.400 ;
        RECT 45.930 17.600 49.930 17.800 ;
        RECT 45.930 17.000 46.330 17.600 ;
        RECT 45.930 16.800 49.930 17.000 ;
        RECT 45.930 16.200 46.330 16.800 ;
        RECT 45.930 16.000 49.930 16.200 ;
        RECT 45.930 15.400 46.330 16.000 ;
        RECT 45.930 15.200 49.930 15.400 ;
        RECT 45.930 14.600 46.330 15.200 ;
        RECT 45.930 14.400 49.930 14.600 ;
        RECT 45.930 13.800 46.330 14.400 ;
        RECT 45.930 13.600 49.930 13.800 ;
        RECT 45.930 13.000 46.330 13.600 ;
        RECT 45.930 12.800 49.930 13.000 ;
        RECT 45.930 12.200 46.330 12.800 ;
        RECT 45.930 12.000 49.930 12.200 ;
        RECT 45.930 11.400 46.330 12.000 ;
        RECT 45.930 11.200 49.930 11.400 ;
        RECT 45.930 10.600 46.330 11.200 ;
        RECT 45.930 10.400 49.930 10.600 ;
        RECT 45.930 10.200 46.330 10.400 ;
        RECT 50.680 10.200 50.880 17.800 ;
        RECT 51.480 10.200 51.680 17.800 ;
        RECT 52.280 10.200 52.480 17.800 ;
        RECT 53.080 10.200 53.280 17.800 ;
        RECT 53.880 10.200 54.080 17.800 ;
        RECT 45.930 9.800 54.080 10.200 ;
        RECT 45.930 9.600 46.330 9.800 ;
        RECT 45.930 9.400 49.930 9.600 ;
        RECT 45.930 8.800 46.330 9.400 ;
        RECT 45.930 8.600 49.930 8.800 ;
        RECT 45.930 8.000 46.330 8.600 ;
        RECT 45.930 7.800 49.930 8.000 ;
        RECT 45.930 7.200 46.330 7.800 ;
        RECT 45.930 7.000 49.930 7.200 ;
        RECT 45.930 6.400 46.330 7.000 ;
        RECT 45.930 6.200 49.930 6.400 ;
        RECT 45.930 5.600 46.330 6.200 ;
        RECT 45.930 5.400 49.930 5.600 ;
        RECT 45.930 4.800 46.330 5.400 ;
        RECT 45.930 4.600 49.930 4.800 ;
        RECT 45.930 4.000 46.330 4.600 ;
        RECT 45.930 3.800 49.930 4.000 ;
        RECT 45.930 3.200 46.330 3.800 ;
        RECT 45.930 3.000 49.930 3.200 ;
        RECT 45.930 2.400 46.330 3.000 ;
        RECT 45.930 2.200 49.930 2.400 ;
        RECT 50.680 2.200 50.880 9.800 ;
        RECT 51.480 2.200 51.680 9.800 ;
        RECT 52.280 2.200 52.480 9.800 ;
        RECT 53.080 2.200 53.280 9.800 ;
        RECT 53.880 2.200 54.080 9.800 ;
        RECT 55.380 10.200 55.580 17.800 ;
        RECT 56.180 10.200 56.380 17.800 ;
        RECT 56.980 10.200 57.180 17.800 ;
        RECT 57.780 10.200 57.980 17.800 ;
        RECT 58.580 10.200 58.780 17.800 ;
        RECT 59.530 17.600 63.530 17.800 ;
        RECT 63.130 17.000 63.530 17.600 ;
        RECT 59.530 16.800 63.530 17.000 ;
        RECT 63.130 16.200 63.530 16.800 ;
        RECT 59.530 16.000 63.530 16.200 ;
        RECT 63.130 15.400 63.530 16.000 ;
        RECT 59.530 15.200 63.530 15.400 ;
        RECT 63.130 14.600 63.530 15.200 ;
        RECT 59.530 14.400 63.530 14.600 ;
        RECT 63.130 13.800 63.530 14.400 ;
        RECT 59.530 13.600 63.530 13.800 ;
        RECT 63.130 13.000 63.530 13.600 ;
        RECT 59.530 12.800 63.530 13.000 ;
        RECT 63.130 12.200 63.530 12.800 ;
        RECT 59.530 12.000 63.530 12.200 ;
        RECT 63.130 11.400 63.530 12.000 ;
        RECT 59.530 11.200 63.530 11.400 ;
        RECT 63.130 10.600 63.530 11.200 ;
        RECT 59.530 10.400 63.530 10.600 ;
        RECT 63.130 10.200 63.530 10.400 ;
        RECT 55.380 9.800 63.530 10.200 ;
        RECT 55.380 2.200 55.580 9.800 ;
        RECT 56.180 2.200 56.380 9.800 ;
        RECT 56.980 2.200 57.180 9.800 ;
        RECT 57.780 2.200 57.980 9.800 ;
        RECT 58.580 2.200 58.780 9.800 ;
        RECT 63.130 9.600 63.530 9.800 ;
        RECT 59.530 9.400 63.530 9.600 ;
        RECT 63.130 8.800 63.530 9.400 ;
        RECT 59.530 8.600 63.530 8.800 ;
        RECT 63.130 8.000 63.530 8.600 ;
        RECT 59.530 7.800 63.530 8.000 ;
        RECT 63.130 7.200 63.530 7.800 ;
        RECT 59.530 7.000 63.530 7.200 ;
        RECT 63.130 6.400 63.530 7.000 ;
        RECT 59.530 6.200 63.530 6.400 ;
        RECT 63.130 5.600 63.530 6.200 ;
        RECT 59.530 5.400 63.530 5.600 ;
        RECT 63.130 4.800 63.530 5.400 ;
        RECT 59.530 4.600 63.530 4.800 ;
        RECT 63.130 4.000 63.530 4.600 ;
        RECT 59.530 3.800 63.530 4.000 ;
        RECT 63.130 3.200 63.530 3.800 ;
        RECT 59.530 3.000 63.530 3.200 ;
        RECT 63.130 2.400 63.530 3.000 ;
        RECT 59.530 2.200 63.530 2.400 ;
        RECT 65.930 17.600 69.930 17.800 ;
        RECT 65.930 17.000 66.330 17.600 ;
        RECT 65.930 16.800 69.930 17.000 ;
        RECT 65.930 16.200 66.330 16.800 ;
        RECT 65.930 16.000 69.930 16.200 ;
        RECT 65.930 15.400 66.330 16.000 ;
        RECT 65.930 15.200 69.930 15.400 ;
        RECT 65.930 14.600 66.330 15.200 ;
        RECT 65.930 14.400 69.930 14.600 ;
        RECT 65.930 13.800 66.330 14.400 ;
        RECT 65.930 13.600 69.930 13.800 ;
        RECT 65.930 13.000 66.330 13.600 ;
        RECT 65.930 12.800 69.930 13.000 ;
        RECT 65.930 12.200 66.330 12.800 ;
        RECT 65.930 12.000 69.930 12.200 ;
        RECT 65.930 11.400 66.330 12.000 ;
        RECT 65.930 11.200 69.930 11.400 ;
        RECT 65.930 10.600 66.330 11.200 ;
        RECT 65.930 10.400 69.930 10.600 ;
        RECT 65.930 10.200 66.330 10.400 ;
        RECT 70.680 10.200 70.880 17.800 ;
        RECT 71.480 10.200 71.680 17.800 ;
        RECT 72.280 10.200 72.480 17.800 ;
        RECT 73.080 10.200 73.280 17.800 ;
        RECT 73.880 10.200 74.080 17.800 ;
        RECT 65.930 9.800 74.080 10.200 ;
        RECT 65.930 9.600 66.330 9.800 ;
        RECT 65.930 9.400 69.930 9.600 ;
        RECT 65.930 8.800 66.330 9.400 ;
        RECT 65.930 8.600 69.930 8.800 ;
        RECT 65.930 8.000 66.330 8.600 ;
        RECT 65.930 7.800 69.930 8.000 ;
        RECT 65.930 7.200 66.330 7.800 ;
        RECT 65.930 7.000 69.930 7.200 ;
        RECT 65.930 6.400 66.330 7.000 ;
        RECT 65.930 6.200 69.930 6.400 ;
        RECT 65.930 5.600 66.330 6.200 ;
        RECT 65.930 5.400 69.930 5.600 ;
        RECT 65.930 4.800 66.330 5.400 ;
        RECT 65.930 4.600 69.930 4.800 ;
        RECT 65.930 4.000 66.330 4.600 ;
        RECT 65.930 3.800 69.930 4.000 ;
        RECT 65.930 3.200 66.330 3.800 ;
        RECT 65.930 3.000 69.930 3.200 ;
        RECT 65.930 2.400 66.330 3.000 ;
        RECT 65.930 2.200 69.930 2.400 ;
        RECT 70.680 2.200 70.880 9.800 ;
        RECT 71.480 2.200 71.680 9.800 ;
        RECT 72.280 2.200 72.480 9.800 ;
        RECT 73.080 2.200 73.280 9.800 ;
        RECT 73.880 2.200 74.080 9.800 ;
        RECT 75.380 10.200 75.580 17.800 ;
        RECT 76.180 10.200 76.380 17.800 ;
        RECT 76.980 10.200 77.180 17.800 ;
        RECT 77.780 10.200 77.980 17.800 ;
        RECT 78.580 10.200 78.780 17.800 ;
        RECT 79.530 17.600 83.530 17.800 ;
        RECT 83.130 17.000 83.530 17.600 ;
        RECT 79.530 16.800 83.530 17.000 ;
        RECT 83.130 16.200 83.530 16.800 ;
        RECT 79.530 16.000 83.530 16.200 ;
        RECT 83.130 15.400 83.530 16.000 ;
        RECT 79.530 15.200 83.530 15.400 ;
        RECT 83.130 14.600 83.530 15.200 ;
        RECT 79.530 14.400 83.530 14.600 ;
        RECT 83.130 13.800 83.530 14.400 ;
        RECT 79.530 13.600 83.530 13.800 ;
        RECT 83.130 13.000 83.530 13.600 ;
        RECT 79.530 12.800 83.530 13.000 ;
        RECT 83.130 12.200 83.530 12.800 ;
        RECT 79.530 12.000 83.530 12.200 ;
        RECT 83.130 11.400 83.530 12.000 ;
        RECT 79.530 11.200 83.530 11.400 ;
        RECT 83.130 10.600 83.530 11.200 ;
        RECT 79.530 10.400 83.530 10.600 ;
        RECT 83.130 10.200 83.530 10.400 ;
        RECT 75.380 9.800 83.530 10.200 ;
        RECT 75.380 2.200 75.580 9.800 ;
        RECT 76.180 2.200 76.380 9.800 ;
        RECT 76.980 2.200 77.180 9.800 ;
        RECT 77.780 2.200 77.980 9.800 ;
        RECT 78.580 2.200 78.780 9.800 ;
        RECT 83.130 9.600 83.530 9.800 ;
        RECT 79.530 9.400 83.530 9.600 ;
        RECT 83.130 8.800 83.530 9.400 ;
        RECT 79.530 8.600 83.530 8.800 ;
        RECT 83.130 8.000 83.530 8.600 ;
        RECT 79.530 7.800 83.530 8.000 ;
        RECT 83.130 7.200 83.530 7.800 ;
        RECT 79.530 7.000 83.530 7.200 ;
        RECT 83.130 6.400 83.530 7.000 ;
        RECT 79.530 6.200 83.530 6.400 ;
        RECT 83.130 5.600 83.530 6.200 ;
        RECT 79.530 5.400 83.530 5.600 ;
        RECT 83.130 4.800 83.530 5.400 ;
        RECT 79.530 4.600 83.530 4.800 ;
        RECT 83.130 4.000 83.530 4.600 ;
        RECT 79.530 3.800 83.530 4.000 ;
        RECT 83.130 3.200 83.530 3.800 ;
        RECT 79.530 3.000 83.530 3.200 ;
        RECT 83.130 2.400 83.530 3.000 ;
        RECT 79.530 2.200 83.530 2.400 ;
        RECT 85.930 17.600 89.930 17.800 ;
        RECT 85.930 17.000 86.330 17.600 ;
        RECT 85.930 16.800 89.930 17.000 ;
        RECT 85.930 16.200 86.330 16.800 ;
        RECT 85.930 16.000 89.930 16.200 ;
        RECT 85.930 15.400 86.330 16.000 ;
        RECT 85.930 15.200 89.930 15.400 ;
        RECT 85.930 14.600 86.330 15.200 ;
        RECT 85.930 14.400 89.930 14.600 ;
        RECT 85.930 13.800 86.330 14.400 ;
        RECT 85.930 13.600 89.930 13.800 ;
        RECT 85.930 13.000 86.330 13.600 ;
        RECT 85.930 12.800 89.930 13.000 ;
        RECT 85.930 12.200 86.330 12.800 ;
        RECT 85.930 12.000 89.930 12.200 ;
        RECT 85.930 11.400 86.330 12.000 ;
        RECT 85.930 11.200 89.930 11.400 ;
        RECT 85.930 10.600 86.330 11.200 ;
        RECT 85.930 10.400 89.930 10.600 ;
        RECT 85.930 10.200 86.330 10.400 ;
        RECT 90.680 10.200 90.880 17.800 ;
        RECT 91.480 10.200 91.680 17.800 ;
        RECT 92.280 10.200 92.480 17.800 ;
        RECT 93.080 10.200 93.280 17.800 ;
        RECT 93.880 10.200 94.080 17.800 ;
        RECT 85.930 9.800 94.080 10.200 ;
        RECT 85.930 9.600 86.330 9.800 ;
        RECT 85.930 9.400 89.930 9.600 ;
        RECT 85.930 8.800 86.330 9.400 ;
        RECT 85.930 8.600 89.930 8.800 ;
        RECT 85.930 8.000 86.330 8.600 ;
        RECT 85.930 7.800 89.930 8.000 ;
        RECT 85.930 7.200 86.330 7.800 ;
        RECT 85.930 7.000 89.930 7.200 ;
        RECT 85.930 6.400 86.330 7.000 ;
        RECT 85.930 6.200 89.930 6.400 ;
        RECT 85.930 5.600 86.330 6.200 ;
        RECT 85.930 5.400 89.930 5.600 ;
        RECT 85.930 4.800 86.330 5.400 ;
        RECT 85.930 4.600 89.930 4.800 ;
        RECT 85.930 4.000 86.330 4.600 ;
        RECT 85.930 3.800 89.930 4.000 ;
        RECT 85.930 3.200 86.330 3.800 ;
        RECT 85.930 3.000 89.930 3.200 ;
        RECT 85.930 2.400 86.330 3.000 ;
        RECT 85.930 2.200 89.930 2.400 ;
        RECT 90.680 2.200 90.880 9.800 ;
        RECT 91.480 2.200 91.680 9.800 ;
        RECT 92.280 2.200 92.480 9.800 ;
        RECT 93.080 2.200 93.280 9.800 ;
        RECT 93.880 2.200 94.080 9.800 ;
        RECT 95.380 10.200 95.580 17.800 ;
        RECT 96.180 10.200 96.380 17.800 ;
        RECT 96.980 10.200 97.180 17.800 ;
        RECT 97.780 10.200 97.980 17.800 ;
        RECT 98.580 10.200 98.780 17.800 ;
        RECT 99.530 17.600 103.530 17.800 ;
        RECT 103.130 17.000 103.530 17.600 ;
        RECT 99.530 16.800 103.530 17.000 ;
        RECT 103.130 16.200 103.530 16.800 ;
        RECT 99.530 16.000 103.530 16.200 ;
        RECT 103.130 15.400 103.530 16.000 ;
        RECT 99.530 15.200 103.530 15.400 ;
        RECT 103.130 14.600 103.530 15.200 ;
        RECT 99.530 14.400 103.530 14.600 ;
        RECT 103.130 13.800 103.530 14.400 ;
        RECT 99.530 13.600 103.530 13.800 ;
        RECT 103.130 13.000 103.530 13.600 ;
        RECT 99.530 12.800 103.530 13.000 ;
        RECT 103.130 12.200 103.530 12.800 ;
        RECT 99.530 12.000 103.530 12.200 ;
        RECT 103.130 11.400 103.530 12.000 ;
        RECT 99.530 11.200 103.530 11.400 ;
        RECT 103.130 10.600 103.530 11.200 ;
        RECT 110.050 11.020 110.410 11.400 ;
        RECT 110.680 11.020 111.040 11.400 ;
        RECT 111.280 11.020 111.640 11.400 ;
        RECT 99.530 10.400 103.530 10.600 ;
        RECT 110.050 10.430 110.410 10.810 ;
        RECT 110.680 10.430 111.040 10.810 ;
        RECT 111.280 10.430 111.640 10.810 ;
        RECT 103.130 10.200 103.530 10.400 ;
        RECT 95.380 9.800 103.530 10.200 ;
        RECT 95.380 2.200 95.580 9.800 ;
        RECT 96.180 2.200 96.380 9.800 ;
        RECT 96.980 2.200 97.180 9.800 ;
        RECT 97.780 2.200 97.980 9.800 ;
        RECT 98.580 2.200 98.780 9.800 ;
        RECT 103.130 9.600 103.530 9.800 ;
        RECT 99.530 9.400 103.530 9.600 ;
        RECT 103.130 8.800 103.530 9.400 ;
        RECT 99.530 8.600 103.530 8.800 ;
        RECT 103.130 8.000 103.530 8.600 ;
        RECT 99.530 7.800 103.530 8.000 ;
        RECT 103.130 7.200 103.530 7.800 ;
        RECT 99.530 7.000 103.530 7.200 ;
        RECT 103.130 6.400 103.530 7.000 ;
        RECT 99.530 6.200 103.530 6.400 ;
        RECT 103.130 5.600 103.530 6.200 ;
        RECT 99.530 5.400 103.530 5.600 ;
        RECT 103.130 4.800 103.530 5.400 ;
        RECT 99.530 4.600 103.530 4.800 ;
        RECT 103.130 4.000 103.530 4.600 ;
        RECT 99.530 3.800 103.530 4.000 ;
        RECT 103.130 3.200 103.530 3.800 ;
        RECT 99.530 3.000 103.530 3.200 ;
        RECT 103.130 2.400 103.530 3.000 ;
        RECT 99.530 2.200 103.530 2.400 ;
      LAYER mcon ;
        RECT 5.980 374.300 6.280 374.750 ;
        RECT 5.980 373.550 6.280 374.000 ;
        RECT 5.980 372.800 6.280 373.250 ;
        RECT 5.980 372.050 6.280 372.500 ;
        RECT 5.980 371.300 6.280 371.750 ;
        RECT 5.980 370.550 6.280 371.000 ;
        RECT 5.980 369.800 6.280 370.250 ;
        RECT 5.980 369.050 6.280 369.500 ;
        RECT 5.980 368.300 6.280 368.750 ;
        RECT 5.980 367.550 6.280 368.000 ;
        RECT 5.980 366.800 6.280 367.250 ;
        RECT 5.980 366.050 6.280 366.500 ;
        RECT 5.980 365.300 6.280 365.750 ;
        RECT 23.180 374.300 23.480 374.750 ;
        RECT 23.180 373.550 23.480 374.000 ;
        RECT 23.180 372.800 23.480 373.250 ;
        RECT 23.180 372.050 23.480 372.500 ;
        RECT 23.180 371.300 23.480 371.750 ;
        RECT 23.180 370.550 23.480 371.000 ;
        RECT 23.180 369.800 23.480 370.250 ;
        RECT 23.180 369.050 23.480 369.500 ;
        RECT 23.180 368.300 23.480 368.750 ;
        RECT 23.180 367.550 23.480 368.000 ;
        RECT 23.180 366.800 23.480 367.250 ;
        RECT 23.180 366.050 23.480 366.500 ;
        RECT 23.180 365.300 23.480 365.750 ;
        RECT 25.980 374.300 26.280 374.750 ;
        RECT 25.980 373.550 26.280 374.000 ;
        RECT 25.980 372.800 26.280 373.250 ;
        RECT 25.980 372.050 26.280 372.500 ;
        RECT 25.980 371.300 26.280 371.750 ;
        RECT 25.980 370.550 26.280 371.000 ;
        RECT 25.980 369.800 26.280 370.250 ;
        RECT 25.980 369.050 26.280 369.500 ;
        RECT 25.980 368.300 26.280 368.750 ;
        RECT 25.980 367.550 26.280 368.000 ;
        RECT 25.980 366.800 26.280 367.250 ;
        RECT 25.980 366.050 26.280 366.500 ;
        RECT 25.980 365.300 26.280 365.750 ;
        RECT 43.180 374.300 43.480 374.750 ;
        RECT 43.180 373.550 43.480 374.000 ;
        RECT 43.180 372.800 43.480 373.250 ;
        RECT 43.180 372.050 43.480 372.500 ;
        RECT 43.180 371.300 43.480 371.750 ;
        RECT 43.180 370.550 43.480 371.000 ;
        RECT 43.180 369.800 43.480 370.250 ;
        RECT 43.180 369.050 43.480 369.500 ;
        RECT 43.180 368.300 43.480 368.750 ;
        RECT 43.180 367.550 43.480 368.000 ;
        RECT 43.180 366.800 43.480 367.250 ;
        RECT 43.180 366.050 43.480 366.500 ;
        RECT 43.180 365.300 43.480 365.750 ;
        RECT 45.980 374.300 46.280 374.750 ;
        RECT 45.980 373.550 46.280 374.000 ;
        RECT 45.980 372.800 46.280 373.250 ;
        RECT 45.980 372.050 46.280 372.500 ;
        RECT 45.980 371.300 46.280 371.750 ;
        RECT 45.980 370.550 46.280 371.000 ;
        RECT 45.980 369.800 46.280 370.250 ;
        RECT 45.980 369.050 46.280 369.500 ;
        RECT 45.980 368.300 46.280 368.750 ;
        RECT 45.980 367.550 46.280 368.000 ;
        RECT 45.980 366.800 46.280 367.250 ;
        RECT 45.980 366.050 46.280 366.500 ;
        RECT 45.980 365.300 46.280 365.750 ;
        RECT 63.180 374.300 63.480 374.750 ;
        RECT 63.180 373.550 63.480 374.000 ;
        RECT 63.180 372.800 63.480 373.250 ;
        RECT 63.180 372.050 63.480 372.500 ;
        RECT 63.180 371.300 63.480 371.750 ;
        RECT 63.180 370.550 63.480 371.000 ;
        RECT 63.180 369.800 63.480 370.250 ;
        RECT 63.180 369.050 63.480 369.500 ;
        RECT 63.180 368.300 63.480 368.750 ;
        RECT 63.180 367.550 63.480 368.000 ;
        RECT 63.180 366.800 63.480 367.250 ;
        RECT 63.180 366.050 63.480 366.500 ;
        RECT 63.180 365.300 63.480 365.750 ;
        RECT 65.980 374.300 66.280 374.750 ;
        RECT 65.980 373.550 66.280 374.000 ;
        RECT 65.980 372.800 66.280 373.250 ;
        RECT 65.980 372.050 66.280 372.500 ;
        RECT 65.980 371.300 66.280 371.750 ;
        RECT 65.980 370.550 66.280 371.000 ;
        RECT 65.980 369.800 66.280 370.250 ;
        RECT 65.980 369.050 66.280 369.500 ;
        RECT 65.980 368.300 66.280 368.750 ;
        RECT 65.980 367.550 66.280 368.000 ;
        RECT 65.980 366.800 66.280 367.250 ;
        RECT 65.980 366.050 66.280 366.500 ;
        RECT 65.980 365.300 66.280 365.750 ;
        RECT 83.180 374.300 83.480 374.750 ;
        RECT 83.180 373.550 83.480 374.000 ;
        RECT 83.180 372.800 83.480 373.250 ;
        RECT 83.180 372.050 83.480 372.500 ;
        RECT 83.180 371.300 83.480 371.750 ;
        RECT 83.180 370.550 83.480 371.000 ;
        RECT 83.180 369.800 83.480 370.250 ;
        RECT 83.180 369.050 83.480 369.500 ;
        RECT 83.180 368.300 83.480 368.750 ;
        RECT 83.180 367.550 83.480 368.000 ;
        RECT 83.180 366.800 83.480 367.250 ;
        RECT 83.180 366.050 83.480 366.500 ;
        RECT 83.180 365.300 83.480 365.750 ;
        RECT 85.980 374.300 86.280 374.750 ;
        RECT 85.980 373.550 86.280 374.000 ;
        RECT 85.980 372.800 86.280 373.250 ;
        RECT 85.980 372.050 86.280 372.500 ;
        RECT 85.980 371.300 86.280 371.750 ;
        RECT 85.980 370.550 86.280 371.000 ;
        RECT 85.980 369.800 86.280 370.250 ;
        RECT 85.980 369.050 86.280 369.500 ;
        RECT 85.980 368.300 86.280 368.750 ;
        RECT 85.980 367.550 86.280 368.000 ;
        RECT 85.980 366.800 86.280 367.250 ;
        RECT 85.980 366.050 86.280 366.500 ;
        RECT 85.980 365.300 86.280 365.750 ;
        RECT 103.180 374.300 103.480 374.750 ;
        RECT 103.180 373.550 103.480 374.000 ;
        RECT 103.180 372.800 103.480 373.250 ;
        RECT 103.180 372.050 103.480 372.500 ;
        RECT 103.180 371.300 103.480 371.750 ;
        RECT 103.180 370.550 103.480 371.000 ;
        RECT 103.180 369.800 103.480 370.250 ;
        RECT 103.180 369.050 103.480 369.500 ;
        RECT 103.180 368.300 103.480 368.750 ;
        RECT 103.180 367.550 103.480 368.000 ;
        RECT 103.180 366.800 103.480 367.250 ;
        RECT 103.180 366.050 103.480 366.500 ;
        RECT 103.180 365.300 103.480 365.750 ;
        RECT 5.980 354.300 6.280 354.750 ;
        RECT 5.980 353.550 6.280 354.000 ;
        RECT 5.980 352.800 6.280 353.250 ;
        RECT 5.980 352.050 6.280 352.500 ;
        RECT 5.980 351.300 6.280 351.750 ;
        RECT 5.980 350.550 6.280 351.000 ;
        RECT 5.980 349.800 6.280 350.250 ;
        RECT 5.980 349.050 6.280 349.500 ;
        RECT 5.980 348.300 6.280 348.750 ;
        RECT 5.980 347.550 6.280 348.000 ;
        RECT 5.980 346.800 6.280 347.250 ;
        RECT 5.980 346.050 6.280 346.500 ;
        RECT 5.980 345.300 6.280 345.750 ;
        RECT 23.180 354.300 23.480 354.750 ;
        RECT 23.180 353.550 23.480 354.000 ;
        RECT 23.180 352.800 23.480 353.250 ;
        RECT 23.180 352.050 23.480 352.500 ;
        RECT 23.180 351.300 23.480 351.750 ;
        RECT 23.180 350.550 23.480 351.000 ;
        RECT 23.180 349.800 23.480 350.250 ;
        RECT 23.180 349.050 23.480 349.500 ;
        RECT 23.180 348.300 23.480 348.750 ;
        RECT 23.180 347.550 23.480 348.000 ;
        RECT 23.180 346.800 23.480 347.250 ;
        RECT 23.180 346.050 23.480 346.500 ;
        RECT 23.180 345.300 23.480 345.750 ;
        RECT 25.980 354.300 26.280 354.750 ;
        RECT 25.980 353.550 26.280 354.000 ;
        RECT 25.980 352.800 26.280 353.250 ;
        RECT 25.980 352.050 26.280 352.500 ;
        RECT 25.980 351.300 26.280 351.750 ;
        RECT 25.980 350.550 26.280 351.000 ;
        RECT 25.980 349.800 26.280 350.250 ;
        RECT 25.980 349.050 26.280 349.500 ;
        RECT 25.980 348.300 26.280 348.750 ;
        RECT 25.980 347.550 26.280 348.000 ;
        RECT 25.980 346.800 26.280 347.250 ;
        RECT 25.980 346.050 26.280 346.500 ;
        RECT 25.980 345.300 26.280 345.750 ;
        RECT 43.180 354.300 43.480 354.750 ;
        RECT 43.180 353.550 43.480 354.000 ;
        RECT 43.180 352.800 43.480 353.250 ;
        RECT 43.180 352.050 43.480 352.500 ;
        RECT 43.180 351.300 43.480 351.750 ;
        RECT 43.180 350.550 43.480 351.000 ;
        RECT 43.180 349.800 43.480 350.250 ;
        RECT 43.180 349.050 43.480 349.500 ;
        RECT 43.180 348.300 43.480 348.750 ;
        RECT 43.180 347.550 43.480 348.000 ;
        RECT 43.180 346.800 43.480 347.250 ;
        RECT 43.180 346.050 43.480 346.500 ;
        RECT 43.180 345.300 43.480 345.750 ;
        RECT 45.980 354.300 46.280 354.750 ;
        RECT 45.980 353.550 46.280 354.000 ;
        RECT 45.980 352.800 46.280 353.250 ;
        RECT 45.980 352.050 46.280 352.500 ;
        RECT 45.980 351.300 46.280 351.750 ;
        RECT 45.980 350.550 46.280 351.000 ;
        RECT 45.980 349.800 46.280 350.250 ;
        RECT 45.980 349.050 46.280 349.500 ;
        RECT 45.980 348.300 46.280 348.750 ;
        RECT 45.980 347.550 46.280 348.000 ;
        RECT 45.980 346.800 46.280 347.250 ;
        RECT 45.980 346.050 46.280 346.500 ;
        RECT 45.980 345.300 46.280 345.750 ;
        RECT 63.180 354.300 63.480 354.750 ;
        RECT 63.180 353.550 63.480 354.000 ;
        RECT 63.180 352.800 63.480 353.250 ;
        RECT 63.180 352.050 63.480 352.500 ;
        RECT 63.180 351.300 63.480 351.750 ;
        RECT 63.180 350.550 63.480 351.000 ;
        RECT 63.180 349.800 63.480 350.250 ;
        RECT 63.180 349.050 63.480 349.500 ;
        RECT 63.180 348.300 63.480 348.750 ;
        RECT 63.180 347.550 63.480 348.000 ;
        RECT 63.180 346.800 63.480 347.250 ;
        RECT 63.180 346.050 63.480 346.500 ;
        RECT 63.180 345.300 63.480 345.750 ;
        RECT 65.980 354.300 66.280 354.750 ;
        RECT 65.980 353.550 66.280 354.000 ;
        RECT 65.980 352.800 66.280 353.250 ;
        RECT 65.980 352.050 66.280 352.500 ;
        RECT 65.980 351.300 66.280 351.750 ;
        RECT 65.980 350.550 66.280 351.000 ;
        RECT 65.980 349.800 66.280 350.250 ;
        RECT 65.980 349.050 66.280 349.500 ;
        RECT 65.980 348.300 66.280 348.750 ;
        RECT 65.980 347.550 66.280 348.000 ;
        RECT 65.980 346.800 66.280 347.250 ;
        RECT 65.980 346.050 66.280 346.500 ;
        RECT 65.980 345.300 66.280 345.750 ;
        RECT 83.180 354.300 83.480 354.750 ;
        RECT 83.180 353.550 83.480 354.000 ;
        RECT 83.180 352.800 83.480 353.250 ;
        RECT 83.180 352.050 83.480 352.500 ;
        RECT 83.180 351.300 83.480 351.750 ;
        RECT 83.180 350.550 83.480 351.000 ;
        RECT 83.180 349.800 83.480 350.250 ;
        RECT 83.180 349.050 83.480 349.500 ;
        RECT 83.180 348.300 83.480 348.750 ;
        RECT 83.180 347.550 83.480 348.000 ;
        RECT 83.180 346.800 83.480 347.250 ;
        RECT 83.180 346.050 83.480 346.500 ;
        RECT 83.180 345.300 83.480 345.750 ;
        RECT 85.980 354.300 86.280 354.750 ;
        RECT 85.980 353.550 86.280 354.000 ;
        RECT 85.980 352.800 86.280 353.250 ;
        RECT 85.980 352.050 86.280 352.500 ;
        RECT 85.980 351.300 86.280 351.750 ;
        RECT 85.980 350.550 86.280 351.000 ;
        RECT 85.980 349.800 86.280 350.250 ;
        RECT 85.980 349.050 86.280 349.500 ;
        RECT 85.980 348.300 86.280 348.750 ;
        RECT 85.980 347.550 86.280 348.000 ;
        RECT 85.980 346.800 86.280 347.250 ;
        RECT 85.980 346.050 86.280 346.500 ;
        RECT 85.980 345.300 86.280 345.750 ;
        RECT 103.180 354.300 103.480 354.750 ;
        RECT 103.180 353.550 103.480 354.000 ;
        RECT 103.180 352.800 103.480 353.250 ;
        RECT 103.180 352.050 103.480 352.500 ;
        RECT 103.180 351.300 103.480 351.750 ;
        RECT 103.180 350.550 103.480 351.000 ;
        RECT 103.180 349.800 103.480 350.250 ;
        RECT 103.180 349.050 103.480 349.500 ;
        RECT 103.180 348.300 103.480 348.750 ;
        RECT 103.180 347.550 103.480 348.000 ;
        RECT 103.180 346.800 103.480 347.250 ;
        RECT 103.180 346.050 103.480 346.500 ;
        RECT 103.180 345.300 103.480 345.750 ;
        RECT 5.980 334.300 6.280 334.750 ;
        RECT 5.980 333.550 6.280 334.000 ;
        RECT 5.980 332.800 6.280 333.250 ;
        RECT 5.980 332.050 6.280 332.500 ;
        RECT 5.980 331.300 6.280 331.750 ;
        RECT 5.980 330.550 6.280 331.000 ;
        RECT 5.980 329.800 6.280 330.250 ;
        RECT 5.980 329.050 6.280 329.500 ;
        RECT 5.980 328.300 6.280 328.750 ;
        RECT 5.980 327.550 6.280 328.000 ;
        RECT 5.980 326.800 6.280 327.250 ;
        RECT 5.980 326.050 6.280 326.500 ;
        RECT 5.980 325.300 6.280 325.750 ;
        RECT 23.180 334.300 23.480 334.750 ;
        RECT 23.180 333.550 23.480 334.000 ;
        RECT 23.180 332.800 23.480 333.250 ;
        RECT 23.180 332.050 23.480 332.500 ;
        RECT 23.180 331.300 23.480 331.750 ;
        RECT 23.180 330.550 23.480 331.000 ;
        RECT 23.180 329.800 23.480 330.250 ;
        RECT 23.180 329.050 23.480 329.500 ;
        RECT 23.180 328.300 23.480 328.750 ;
        RECT 23.180 327.550 23.480 328.000 ;
        RECT 23.180 326.800 23.480 327.250 ;
        RECT 23.180 326.050 23.480 326.500 ;
        RECT 23.180 325.300 23.480 325.750 ;
        RECT 25.980 334.300 26.280 334.750 ;
        RECT 25.980 333.550 26.280 334.000 ;
        RECT 25.980 332.800 26.280 333.250 ;
        RECT 25.980 332.050 26.280 332.500 ;
        RECT 25.980 331.300 26.280 331.750 ;
        RECT 25.980 330.550 26.280 331.000 ;
        RECT 25.980 329.800 26.280 330.250 ;
        RECT 25.980 329.050 26.280 329.500 ;
        RECT 25.980 328.300 26.280 328.750 ;
        RECT 25.980 327.550 26.280 328.000 ;
        RECT 25.980 326.800 26.280 327.250 ;
        RECT 25.980 326.050 26.280 326.500 ;
        RECT 25.980 325.300 26.280 325.750 ;
        RECT 43.180 334.300 43.480 334.750 ;
        RECT 43.180 333.550 43.480 334.000 ;
        RECT 43.180 332.800 43.480 333.250 ;
        RECT 43.180 332.050 43.480 332.500 ;
        RECT 43.180 331.300 43.480 331.750 ;
        RECT 43.180 330.550 43.480 331.000 ;
        RECT 43.180 329.800 43.480 330.250 ;
        RECT 43.180 329.050 43.480 329.500 ;
        RECT 43.180 328.300 43.480 328.750 ;
        RECT 43.180 327.550 43.480 328.000 ;
        RECT 43.180 326.800 43.480 327.250 ;
        RECT 43.180 326.050 43.480 326.500 ;
        RECT 43.180 325.300 43.480 325.750 ;
        RECT 45.980 334.300 46.280 334.750 ;
        RECT 45.980 333.550 46.280 334.000 ;
        RECT 45.980 332.800 46.280 333.250 ;
        RECT 45.980 332.050 46.280 332.500 ;
        RECT 45.980 331.300 46.280 331.750 ;
        RECT 45.980 330.550 46.280 331.000 ;
        RECT 45.980 329.800 46.280 330.250 ;
        RECT 45.980 329.050 46.280 329.500 ;
        RECT 45.980 328.300 46.280 328.750 ;
        RECT 45.980 327.550 46.280 328.000 ;
        RECT 45.980 326.800 46.280 327.250 ;
        RECT 45.980 326.050 46.280 326.500 ;
        RECT 45.980 325.300 46.280 325.750 ;
        RECT 63.180 334.300 63.480 334.750 ;
        RECT 63.180 333.550 63.480 334.000 ;
        RECT 63.180 332.800 63.480 333.250 ;
        RECT 63.180 332.050 63.480 332.500 ;
        RECT 63.180 331.300 63.480 331.750 ;
        RECT 63.180 330.550 63.480 331.000 ;
        RECT 63.180 329.800 63.480 330.250 ;
        RECT 63.180 329.050 63.480 329.500 ;
        RECT 63.180 328.300 63.480 328.750 ;
        RECT 63.180 327.550 63.480 328.000 ;
        RECT 63.180 326.800 63.480 327.250 ;
        RECT 63.180 326.050 63.480 326.500 ;
        RECT 63.180 325.300 63.480 325.750 ;
        RECT 65.980 334.300 66.280 334.750 ;
        RECT 65.980 333.550 66.280 334.000 ;
        RECT 65.980 332.800 66.280 333.250 ;
        RECT 65.980 332.050 66.280 332.500 ;
        RECT 65.980 331.300 66.280 331.750 ;
        RECT 65.980 330.550 66.280 331.000 ;
        RECT 65.980 329.800 66.280 330.250 ;
        RECT 65.980 329.050 66.280 329.500 ;
        RECT 65.980 328.300 66.280 328.750 ;
        RECT 65.980 327.550 66.280 328.000 ;
        RECT 65.980 326.800 66.280 327.250 ;
        RECT 65.980 326.050 66.280 326.500 ;
        RECT 65.980 325.300 66.280 325.750 ;
        RECT 83.180 334.300 83.480 334.750 ;
        RECT 83.180 333.550 83.480 334.000 ;
        RECT 83.180 332.800 83.480 333.250 ;
        RECT 83.180 332.050 83.480 332.500 ;
        RECT 83.180 331.300 83.480 331.750 ;
        RECT 83.180 330.550 83.480 331.000 ;
        RECT 83.180 329.800 83.480 330.250 ;
        RECT 83.180 329.050 83.480 329.500 ;
        RECT 83.180 328.300 83.480 328.750 ;
        RECT 83.180 327.550 83.480 328.000 ;
        RECT 83.180 326.800 83.480 327.250 ;
        RECT 83.180 326.050 83.480 326.500 ;
        RECT 83.180 325.300 83.480 325.750 ;
        RECT 85.980 334.300 86.280 334.750 ;
        RECT 85.980 333.550 86.280 334.000 ;
        RECT 85.980 332.800 86.280 333.250 ;
        RECT 85.980 332.050 86.280 332.500 ;
        RECT 85.980 331.300 86.280 331.750 ;
        RECT 85.980 330.550 86.280 331.000 ;
        RECT 85.980 329.800 86.280 330.250 ;
        RECT 85.980 329.050 86.280 329.500 ;
        RECT 85.980 328.300 86.280 328.750 ;
        RECT 85.980 327.550 86.280 328.000 ;
        RECT 85.980 326.800 86.280 327.250 ;
        RECT 85.980 326.050 86.280 326.500 ;
        RECT 85.980 325.300 86.280 325.750 ;
        RECT 103.180 334.300 103.480 334.750 ;
        RECT 103.180 333.550 103.480 334.000 ;
        RECT 103.180 332.800 103.480 333.250 ;
        RECT 103.180 332.050 103.480 332.500 ;
        RECT 103.180 331.300 103.480 331.750 ;
        RECT 103.180 330.550 103.480 331.000 ;
        RECT 103.180 329.800 103.480 330.250 ;
        RECT 103.180 329.050 103.480 329.500 ;
        RECT 103.180 328.300 103.480 328.750 ;
        RECT 103.180 327.550 103.480 328.000 ;
        RECT 103.180 326.800 103.480 327.250 ;
        RECT 103.180 326.050 103.480 326.500 ;
        RECT 103.180 325.300 103.480 325.750 ;
        RECT 5.980 314.300 6.280 314.750 ;
        RECT 5.980 313.550 6.280 314.000 ;
        RECT 5.980 312.800 6.280 313.250 ;
        RECT 5.980 312.050 6.280 312.500 ;
        RECT 5.980 311.300 6.280 311.750 ;
        RECT 5.980 310.550 6.280 311.000 ;
        RECT 5.980 309.800 6.280 310.250 ;
        RECT 5.980 309.050 6.280 309.500 ;
        RECT 5.980 308.300 6.280 308.750 ;
        RECT 5.980 307.550 6.280 308.000 ;
        RECT 5.980 306.800 6.280 307.250 ;
        RECT 5.980 306.050 6.280 306.500 ;
        RECT 5.980 305.300 6.280 305.750 ;
        RECT 23.180 314.300 23.480 314.750 ;
        RECT 23.180 313.550 23.480 314.000 ;
        RECT 23.180 312.800 23.480 313.250 ;
        RECT 23.180 312.050 23.480 312.500 ;
        RECT 23.180 311.300 23.480 311.750 ;
        RECT 23.180 310.550 23.480 311.000 ;
        RECT 23.180 309.800 23.480 310.250 ;
        RECT 23.180 309.050 23.480 309.500 ;
        RECT 23.180 308.300 23.480 308.750 ;
        RECT 23.180 307.550 23.480 308.000 ;
        RECT 23.180 306.800 23.480 307.250 ;
        RECT 23.180 306.050 23.480 306.500 ;
        RECT 23.180 305.300 23.480 305.750 ;
        RECT 25.980 314.300 26.280 314.750 ;
        RECT 25.980 313.550 26.280 314.000 ;
        RECT 25.980 312.800 26.280 313.250 ;
        RECT 25.980 312.050 26.280 312.500 ;
        RECT 25.980 311.300 26.280 311.750 ;
        RECT 25.980 310.550 26.280 311.000 ;
        RECT 25.980 309.800 26.280 310.250 ;
        RECT 25.980 309.050 26.280 309.500 ;
        RECT 25.980 308.300 26.280 308.750 ;
        RECT 25.980 307.550 26.280 308.000 ;
        RECT 25.980 306.800 26.280 307.250 ;
        RECT 25.980 306.050 26.280 306.500 ;
        RECT 25.980 305.300 26.280 305.750 ;
        RECT 43.180 314.300 43.480 314.750 ;
        RECT 43.180 313.550 43.480 314.000 ;
        RECT 43.180 312.800 43.480 313.250 ;
        RECT 43.180 312.050 43.480 312.500 ;
        RECT 43.180 311.300 43.480 311.750 ;
        RECT 43.180 310.550 43.480 311.000 ;
        RECT 43.180 309.800 43.480 310.250 ;
        RECT 43.180 309.050 43.480 309.500 ;
        RECT 43.180 308.300 43.480 308.750 ;
        RECT 43.180 307.550 43.480 308.000 ;
        RECT 43.180 306.800 43.480 307.250 ;
        RECT 43.180 306.050 43.480 306.500 ;
        RECT 43.180 305.300 43.480 305.750 ;
        RECT 45.980 314.300 46.280 314.750 ;
        RECT 45.980 313.550 46.280 314.000 ;
        RECT 45.980 312.800 46.280 313.250 ;
        RECT 45.980 312.050 46.280 312.500 ;
        RECT 45.980 311.300 46.280 311.750 ;
        RECT 45.980 310.550 46.280 311.000 ;
        RECT 45.980 309.800 46.280 310.250 ;
        RECT 45.980 309.050 46.280 309.500 ;
        RECT 45.980 308.300 46.280 308.750 ;
        RECT 45.980 307.550 46.280 308.000 ;
        RECT 45.980 306.800 46.280 307.250 ;
        RECT 45.980 306.050 46.280 306.500 ;
        RECT 45.980 305.300 46.280 305.750 ;
        RECT 63.180 314.300 63.480 314.750 ;
        RECT 63.180 313.550 63.480 314.000 ;
        RECT 63.180 312.800 63.480 313.250 ;
        RECT 63.180 312.050 63.480 312.500 ;
        RECT 63.180 311.300 63.480 311.750 ;
        RECT 63.180 310.550 63.480 311.000 ;
        RECT 63.180 309.800 63.480 310.250 ;
        RECT 63.180 309.050 63.480 309.500 ;
        RECT 63.180 308.300 63.480 308.750 ;
        RECT 63.180 307.550 63.480 308.000 ;
        RECT 63.180 306.800 63.480 307.250 ;
        RECT 63.180 306.050 63.480 306.500 ;
        RECT 63.180 305.300 63.480 305.750 ;
        RECT 65.980 314.300 66.280 314.750 ;
        RECT 65.980 313.550 66.280 314.000 ;
        RECT 65.980 312.800 66.280 313.250 ;
        RECT 65.980 312.050 66.280 312.500 ;
        RECT 65.980 311.300 66.280 311.750 ;
        RECT 65.980 310.550 66.280 311.000 ;
        RECT 65.980 309.800 66.280 310.250 ;
        RECT 65.980 309.050 66.280 309.500 ;
        RECT 65.980 308.300 66.280 308.750 ;
        RECT 65.980 307.550 66.280 308.000 ;
        RECT 65.980 306.800 66.280 307.250 ;
        RECT 65.980 306.050 66.280 306.500 ;
        RECT 65.980 305.300 66.280 305.750 ;
        RECT 83.180 314.300 83.480 314.750 ;
        RECT 83.180 313.550 83.480 314.000 ;
        RECT 83.180 312.800 83.480 313.250 ;
        RECT 83.180 312.050 83.480 312.500 ;
        RECT 83.180 311.300 83.480 311.750 ;
        RECT 83.180 310.550 83.480 311.000 ;
        RECT 83.180 309.800 83.480 310.250 ;
        RECT 83.180 309.050 83.480 309.500 ;
        RECT 83.180 308.300 83.480 308.750 ;
        RECT 83.180 307.550 83.480 308.000 ;
        RECT 83.180 306.800 83.480 307.250 ;
        RECT 83.180 306.050 83.480 306.500 ;
        RECT 83.180 305.300 83.480 305.750 ;
        RECT 85.980 314.300 86.280 314.750 ;
        RECT 85.980 313.550 86.280 314.000 ;
        RECT 85.980 312.800 86.280 313.250 ;
        RECT 85.980 312.050 86.280 312.500 ;
        RECT 85.980 311.300 86.280 311.750 ;
        RECT 85.980 310.550 86.280 311.000 ;
        RECT 85.980 309.800 86.280 310.250 ;
        RECT 85.980 309.050 86.280 309.500 ;
        RECT 85.980 308.300 86.280 308.750 ;
        RECT 85.980 307.550 86.280 308.000 ;
        RECT 85.980 306.800 86.280 307.250 ;
        RECT 85.980 306.050 86.280 306.500 ;
        RECT 85.980 305.300 86.280 305.750 ;
        RECT 103.180 314.300 103.480 314.750 ;
        RECT 103.180 313.550 103.480 314.000 ;
        RECT 103.180 312.800 103.480 313.250 ;
        RECT 103.180 312.050 103.480 312.500 ;
        RECT 103.180 311.300 103.480 311.750 ;
        RECT 103.180 310.550 103.480 311.000 ;
        RECT 103.180 309.800 103.480 310.250 ;
        RECT 103.180 309.050 103.480 309.500 ;
        RECT 103.180 308.300 103.480 308.750 ;
        RECT 103.180 307.550 103.480 308.000 ;
        RECT 103.180 306.800 103.480 307.250 ;
        RECT 103.180 306.050 103.480 306.500 ;
        RECT 103.180 305.300 103.480 305.750 ;
        RECT 5.980 294.300 6.280 294.750 ;
        RECT 5.980 293.550 6.280 294.000 ;
        RECT 5.980 292.800 6.280 293.250 ;
        RECT 5.980 292.050 6.280 292.500 ;
        RECT 5.980 291.300 6.280 291.750 ;
        RECT 5.980 290.550 6.280 291.000 ;
        RECT 5.980 289.800 6.280 290.250 ;
        RECT 5.980 289.050 6.280 289.500 ;
        RECT 5.980 288.300 6.280 288.750 ;
        RECT 5.980 287.550 6.280 288.000 ;
        RECT 5.980 286.800 6.280 287.250 ;
        RECT 5.980 286.050 6.280 286.500 ;
        RECT 5.980 285.300 6.280 285.750 ;
        RECT 23.180 294.300 23.480 294.750 ;
        RECT 23.180 293.550 23.480 294.000 ;
        RECT 23.180 292.800 23.480 293.250 ;
        RECT 23.180 292.050 23.480 292.500 ;
        RECT 23.180 291.300 23.480 291.750 ;
        RECT 23.180 290.550 23.480 291.000 ;
        RECT 23.180 289.800 23.480 290.250 ;
        RECT 23.180 289.050 23.480 289.500 ;
        RECT 23.180 288.300 23.480 288.750 ;
        RECT 23.180 287.550 23.480 288.000 ;
        RECT 23.180 286.800 23.480 287.250 ;
        RECT 23.180 286.050 23.480 286.500 ;
        RECT 23.180 285.300 23.480 285.750 ;
        RECT 25.980 294.300 26.280 294.750 ;
        RECT 25.980 293.550 26.280 294.000 ;
        RECT 25.980 292.800 26.280 293.250 ;
        RECT 25.980 292.050 26.280 292.500 ;
        RECT 25.980 291.300 26.280 291.750 ;
        RECT 25.980 290.550 26.280 291.000 ;
        RECT 25.980 289.800 26.280 290.250 ;
        RECT 25.980 289.050 26.280 289.500 ;
        RECT 25.980 288.300 26.280 288.750 ;
        RECT 25.980 287.550 26.280 288.000 ;
        RECT 25.980 286.800 26.280 287.250 ;
        RECT 25.980 286.050 26.280 286.500 ;
        RECT 25.980 285.300 26.280 285.750 ;
        RECT 43.180 294.300 43.480 294.750 ;
        RECT 43.180 293.550 43.480 294.000 ;
        RECT 43.180 292.800 43.480 293.250 ;
        RECT 43.180 292.050 43.480 292.500 ;
        RECT 43.180 291.300 43.480 291.750 ;
        RECT 43.180 290.550 43.480 291.000 ;
        RECT 43.180 289.800 43.480 290.250 ;
        RECT 43.180 289.050 43.480 289.500 ;
        RECT 43.180 288.300 43.480 288.750 ;
        RECT 43.180 287.550 43.480 288.000 ;
        RECT 43.180 286.800 43.480 287.250 ;
        RECT 43.180 286.050 43.480 286.500 ;
        RECT 43.180 285.300 43.480 285.750 ;
        RECT 45.980 294.300 46.280 294.750 ;
        RECT 45.980 293.550 46.280 294.000 ;
        RECT 45.980 292.800 46.280 293.250 ;
        RECT 45.980 292.050 46.280 292.500 ;
        RECT 45.980 291.300 46.280 291.750 ;
        RECT 45.980 290.550 46.280 291.000 ;
        RECT 45.980 289.800 46.280 290.250 ;
        RECT 45.980 289.050 46.280 289.500 ;
        RECT 45.980 288.300 46.280 288.750 ;
        RECT 45.980 287.550 46.280 288.000 ;
        RECT 45.980 286.800 46.280 287.250 ;
        RECT 45.980 286.050 46.280 286.500 ;
        RECT 45.980 285.300 46.280 285.750 ;
        RECT 63.180 294.300 63.480 294.750 ;
        RECT 63.180 293.550 63.480 294.000 ;
        RECT 63.180 292.800 63.480 293.250 ;
        RECT 63.180 292.050 63.480 292.500 ;
        RECT 63.180 291.300 63.480 291.750 ;
        RECT 63.180 290.550 63.480 291.000 ;
        RECT 63.180 289.800 63.480 290.250 ;
        RECT 63.180 289.050 63.480 289.500 ;
        RECT 63.180 288.300 63.480 288.750 ;
        RECT 63.180 287.550 63.480 288.000 ;
        RECT 63.180 286.800 63.480 287.250 ;
        RECT 63.180 286.050 63.480 286.500 ;
        RECT 63.180 285.300 63.480 285.750 ;
        RECT 65.980 294.300 66.280 294.750 ;
        RECT 65.980 293.550 66.280 294.000 ;
        RECT 65.980 292.800 66.280 293.250 ;
        RECT 65.980 292.050 66.280 292.500 ;
        RECT 65.980 291.300 66.280 291.750 ;
        RECT 65.980 290.550 66.280 291.000 ;
        RECT 65.980 289.800 66.280 290.250 ;
        RECT 65.980 289.050 66.280 289.500 ;
        RECT 65.980 288.300 66.280 288.750 ;
        RECT 65.980 287.550 66.280 288.000 ;
        RECT 65.980 286.800 66.280 287.250 ;
        RECT 65.980 286.050 66.280 286.500 ;
        RECT 65.980 285.300 66.280 285.750 ;
        RECT 83.180 294.300 83.480 294.750 ;
        RECT 83.180 293.550 83.480 294.000 ;
        RECT 83.180 292.800 83.480 293.250 ;
        RECT 83.180 292.050 83.480 292.500 ;
        RECT 83.180 291.300 83.480 291.750 ;
        RECT 83.180 290.550 83.480 291.000 ;
        RECT 83.180 289.800 83.480 290.250 ;
        RECT 83.180 289.050 83.480 289.500 ;
        RECT 83.180 288.300 83.480 288.750 ;
        RECT 83.180 287.550 83.480 288.000 ;
        RECT 83.180 286.800 83.480 287.250 ;
        RECT 83.180 286.050 83.480 286.500 ;
        RECT 83.180 285.300 83.480 285.750 ;
        RECT 85.980 294.300 86.280 294.750 ;
        RECT 85.980 293.550 86.280 294.000 ;
        RECT 85.980 292.800 86.280 293.250 ;
        RECT 85.980 292.050 86.280 292.500 ;
        RECT 85.980 291.300 86.280 291.750 ;
        RECT 85.980 290.550 86.280 291.000 ;
        RECT 85.980 289.800 86.280 290.250 ;
        RECT 85.980 289.050 86.280 289.500 ;
        RECT 85.980 288.300 86.280 288.750 ;
        RECT 85.980 287.550 86.280 288.000 ;
        RECT 85.980 286.800 86.280 287.250 ;
        RECT 85.980 286.050 86.280 286.500 ;
        RECT 85.980 285.300 86.280 285.750 ;
        RECT 103.180 294.300 103.480 294.750 ;
        RECT 103.180 293.550 103.480 294.000 ;
        RECT 103.180 292.800 103.480 293.250 ;
        RECT 103.180 292.050 103.480 292.500 ;
        RECT 103.180 291.300 103.480 291.750 ;
        RECT 103.180 290.550 103.480 291.000 ;
        RECT 103.180 289.800 103.480 290.250 ;
        RECT 103.180 289.050 103.480 289.500 ;
        RECT 103.180 288.300 103.480 288.750 ;
        RECT 103.180 287.550 103.480 288.000 ;
        RECT 103.180 286.800 103.480 287.250 ;
        RECT 103.180 286.050 103.480 286.500 ;
        RECT 103.180 285.300 103.480 285.750 ;
        RECT 5.980 274.300 6.280 274.750 ;
        RECT 5.980 273.550 6.280 274.000 ;
        RECT 5.980 272.800 6.280 273.250 ;
        RECT 5.980 272.050 6.280 272.500 ;
        RECT 5.980 271.300 6.280 271.750 ;
        RECT 5.980 270.550 6.280 271.000 ;
        RECT 5.980 269.800 6.280 270.250 ;
        RECT 5.980 269.050 6.280 269.500 ;
        RECT 5.980 268.300 6.280 268.750 ;
        RECT 5.980 267.550 6.280 268.000 ;
        RECT 5.980 266.800 6.280 267.250 ;
        RECT 5.980 266.050 6.280 266.500 ;
        RECT 5.980 265.300 6.280 265.750 ;
        RECT 23.180 274.300 23.480 274.750 ;
        RECT 23.180 273.550 23.480 274.000 ;
        RECT 23.180 272.800 23.480 273.250 ;
        RECT 23.180 272.050 23.480 272.500 ;
        RECT 23.180 271.300 23.480 271.750 ;
        RECT 23.180 270.550 23.480 271.000 ;
        RECT 23.180 269.800 23.480 270.250 ;
        RECT 23.180 269.050 23.480 269.500 ;
        RECT 23.180 268.300 23.480 268.750 ;
        RECT 23.180 267.550 23.480 268.000 ;
        RECT 23.180 266.800 23.480 267.250 ;
        RECT 23.180 266.050 23.480 266.500 ;
        RECT 23.180 265.300 23.480 265.750 ;
        RECT 25.980 274.300 26.280 274.750 ;
        RECT 25.980 273.550 26.280 274.000 ;
        RECT 25.980 272.800 26.280 273.250 ;
        RECT 25.980 272.050 26.280 272.500 ;
        RECT 25.980 271.300 26.280 271.750 ;
        RECT 25.980 270.550 26.280 271.000 ;
        RECT 25.980 269.800 26.280 270.250 ;
        RECT 25.980 269.050 26.280 269.500 ;
        RECT 25.980 268.300 26.280 268.750 ;
        RECT 25.980 267.550 26.280 268.000 ;
        RECT 25.980 266.800 26.280 267.250 ;
        RECT 25.980 266.050 26.280 266.500 ;
        RECT 25.980 265.300 26.280 265.750 ;
        RECT 43.180 274.300 43.480 274.750 ;
        RECT 43.180 273.550 43.480 274.000 ;
        RECT 43.180 272.800 43.480 273.250 ;
        RECT 43.180 272.050 43.480 272.500 ;
        RECT 43.180 271.300 43.480 271.750 ;
        RECT 43.180 270.550 43.480 271.000 ;
        RECT 43.180 269.800 43.480 270.250 ;
        RECT 43.180 269.050 43.480 269.500 ;
        RECT 43.180 268.300 43.480 268.750 ;
        RECT 43.180 267.550 43.480 268.000 ;
        RECT 43.180 266.800 43.480 267.250 ;
        RECT 43.180 266.050 43.480 266.500 ;
        RECT 43.180 265.300 43.480 265.750 ;
        RECT 45.980 274.300 46.280 274.750 ;
        RECT 45.980 273.550 46.280 274.000 ;
        RECT 45.980 272.800 46.280 273.250 ;
        RECT 45.980 272.050 46.280 272.500 ;
        RECT 45.980 271.300 46.280 271.750 ;
        RECT 45.980 270.550 46.280 271.000 ;
        RECT 45.980 269.800 46.280 270.250 ;
        RECT 45.980 269.050 46.280 269.500 ;
        RECT 45.980 268.300 46.280 268.750 ;
        RECT 45.980 267.550 46.280 268.000 ;
        RECT 45.980 266.800 46.280 267.250 ;
        RECT 45.980 266.050 46.280 266.500 ;
        RECT 45.980 265.300 46.280 265.750 ;
        RECT 63.180 274.300 63.480 274.750 ;
        RECT 63.180 273.550 63.480 274.000 ;
        RECT 63.180 272.800 63.480 273.250 ;
        RECT 63.180 272.050 63.480 272.500 ;
        RECT 63.180 271.300 63.480 271.750 ;
        RECT 63.180 270.550 63.480 271.000 ;
        RECT 63.180 269.800 63.480 270.250 ;
        RECT 63.180 269.050 63.480 269.500 ;
        RECT 63.180 268.300 63.480 268.750 ;
        RECT 63.180 267.550 63.480 268.000 ;
        RECT 63.180 266.800 63.480 267.250 ;
        RECT 63.180 266.050 63.480 266.500 ;
        RECT 63.180 265.300 63.480 265.750 ;
        RECT 65.980 274.300 66.280 274.750 ;
        RECT 65.980 273.550 66.280 274.000 ;
        RECT 65.980 272.800 66.280 273.250 ;
        RECT 65.980 272.050 66.280 272.500 ;
        RECT 65.980 271.300 66.280 271.750 ;
        RECT 65.980 270.550 66.280 271.000 ;
        RECT 65.980 269.800 66.280 270.250 ;
        RECT 65.980 269.050 66.280 269.500 ;
        RECT 65.980 268.300 66.280 268.750 ;
        RECT 65.980 267.550 66.280 268.000 ;
        RECT 65.980 266.800 66.280 267.250 ;
        RECT 65.980 266.050 66.280 266.500 ;
        RECT 65.980 265.300 66.280 265.750 ;
        RECT 83.180 274.300 83.480 274.750 ;
        RECT 83.180 273.550 83.480 274.000 ;
        RECT 83.180 272.800 83.480 273.250 ;
        RECT 83.180 272.050 83.480 272.500 ;
        RECT 83.180 271.300 83.480 271.750 ;
        RECT 83.180 270.550 83.480 271.000 ;
        RECT 83.180 269.800 83.480 270.250 ;
        RECT 83.180 269.050 83.480 269.500 ;
        RECT 83.180 268.300 83.480 268.750 ;
        RECT 83.180 267.550 83.480 268.000 ;
        RECT 83.180 266.800 83.480 267.250 ;
        RECT 83.180 266.050 83.480 266.500 ;
        RECT 83.180 265.300 83.480 265.750 ;
        RECT 85.980 274.300 86.280 274.750 ;
        RECT 85.980 273.550 86.280 274.000 ;
        RECT 85.980 272.800 86.280 273.250 ;
        RECT 85.980 272.050 86.280 272.500 ;
        RECT 85.980 271.300 86.280 271.750 ;
        RECT 85.980 270.550 86.280 271.000 ;
        RECT 85.980 269.800 86.280 270.250 ;
        RECT 85.980 269.050 86.280 269.500 ;
        RECT 85.980 268.300 86.280 268.750 ;
        RECT 85.980 267.550 86.280 268.000 ;
        RECT 85.980 266.800 86.280 267.250 ;
        RECT 85.980 266.050 86.280 266.500 ;
        RECT 85.980 265.300 86.280 265.750 ;
        RECT 103.180 274.300 103.480 274.750 ;
        RECT 103.180 273.550 103.480 274.000 ;
        RECT 103.180 272.800 103.480 273.250 ;
        RECT 103.180 272.050 103.480 272.500 ;
        RECT 103.180 271.300 103.480 271.750 ;
        RECT 103.180 270.550 103.480 271.000 ;
        RECT 103.180 269.800 103.480 270.250 ;
        RECT 103.180 269.050 103.480 269.500 ;
        RECT 103.180 268.300 103.480 268.750 ;
        RECT 103.180 267.550 103.480 268.000 ;
        RECT 103.180 266.800 103.480 267.250 ;
        RECT 103.180 266.050 103.480 266.500 ;
        RECT 103.180 265.300 103.480 265.750 ;
        RECT 5.980 254.300 6.280 254.750 ;
        RECT 5.980 253.550 6.280 254.000 ;
        RECT 5.980 252.800 6.280 253.250 ;
        RECT 5.980 252.050 6.280 252.500 ;
        RECT 5.980 251.300 6.280 251.750 ;
        RECT 5.980 250.550 6.280 251.000 ;
        RECT 5.980 249.800 6.280 250.250 ;
        RECT 5.980 249.050 6.280 249.500 ;
        RECT 5.980 248.300 6.280 248.750 ;
        RECT 5.980 247.550 6.280 248.000 ;
        RECT 5.980 246.800 6.280 247.250 ;
        RECT 5.980 246.050 6.280 246.500 ;
        RECT 5.980 245.300 6.280 245.750 ;
        RECT 23.180 254.300 23.480 254.750 ;
        RECT 23.180 253.550 23.480 254.000 ;
        RECT 23.180 252.800 23.480 253.250 ;
        RECT 23.180 252.050 23.480 252.500 ;
        RECT 23.180 251.300 23.480 251.750 ;
        RECT 23.180 250.550 23.480 251.000 ;
        RECT 23.180 249.800 23.480 250.250 ;
        RECT 23.180 249.050 23.480 249.500 ;
        RECT 23.180 248.300 23.480 248.750 ;
        RECT 23.180 247.550 23.480 248.000 ;
        RECT 23.180 246.800 23.480 247.250 ;
        RECT 23.180 246.050 23.480 246.500 ;
        RECT 23.180 245.300 23.480 245.750 ;
        RECT 25.980 254.300 26.280 254.750 ;
        RECT 25.980 253.550 26.280 254.000 ;
        RECT 25.980 252.800 26.280 253.250 ;
        RECT 25.980 252.050 26.280 252.500 ;
        RECT 25.980 251.300 26.280 251.750 ;
        RECT 25.980 250.550 26.280 251.000 ;
        RECT 25.980 249.800 26.280 250.250 ;
        RECT 25.980 249.050 26.280 249.500 ;
        RECT 25.980 248.300 26.280 248.750 ;
        RECT 25.980 247.550 26.280 248.000 ;
        RECT 25.980 246.800 26.280 247.250 ;
        RECT 25.980 246.050 26.280 246.500 ;
        RECT 25.980 245.300 26.280 245.750 ;
        RECT 43.180 254.300 43.480 254.750 ;
        RECT 43.180 253.550 43.480 254.000 ;
        RECT 43.180 252.800 43.480 253.250 ;
        RECT 43.180 252.050 43.480 252.500 ;
        RECT 43.180 251.300 43.480 251.750 ;
        RECT 43.180 250.550 43.480 251.000 ;
        RECT 43.180 249.800 43.480 250.250 ;
        RECT 43.180 249.050 43.480 249.500 ;
        RECT 43.180 248.300 43.480 248.750 ;
        RECT 43.180 247.550 43.480 248.000 ;
        RECT 43.180 246.800 43.480 247.250 ;
        RECT 43.180 246.050 43.480 246.500 ;
        RECT 43.180 245.300 43.480 245.750 ;
        RECT 45.980 254.300 46.280 254.750 ;
        RECT 45.980 253.550 46.280 254.000 ;
        RECT 45.980 252.800 46.280 253.250 ;
        RECT 45.980 252.050 46.280 252.500 ;
        RECT 45.980 251.300 46.280 251.750 ;
        RECT 45.980 250.550 46.280 251.000 ;
        RECT 45.980 249.800 46.280 250.250 ;
        RECT 45.980 249.050 46.280 249.500 ;
        RECT 45.980 248.300 46.280 248.750 ;
        RECT 45.980 247.550 46.280 248.000 ;
        RECT 45.980 246.800 46.280 247.250 ;
        RECT 45.980 246.050 46.280 246.500 ;
        RECT 45.980 245.300 46.280 245.750 ;
        RECT 63.180 254.300 63.480 254.750 ;
        RECT 63.180 253.550 63.480 254.000 ;
        RECT 63.180 252.800 63.480 253.250 ;
        RECT 63.180 252.050 63.480 252.500 ;
        RECT 63.180 251.300 63.480 251.750 ;
        RECT 63.180 250.550 63.480 251.000 ;
        RECT 63.180 249.800 63.480 250.250 ;
        RECT 63.180 249.050 63.480 249.500 ;
        RECT 63.180 248.300 63.480 248.750 ;
        RECT 63.180 247.550 63.480 248.000 ;
        RECT 63.180 246.800 63.480 247.250 ;
        RECT 63.180 246.050 63.480 246.500 ;
        RECT 63.180 245.300 63.480 245.750 ;
        RECT 65.980 254.300 66.280 254.750 ;
        RECT 65.980 253.550 66.280 254.000 ;
        RECT 65.980 252.800 66.280 253.250 ;
        RECT 65.980 252.050 66.280 252.500 ;
        RECT 65.980 251.300 66.280 251.750 ;
        RECT 65.980 250.550 66.280 251.000 ;
        RECT 65.980 249.800 66.280 250.250 ;
        RECT 65.980 249.050 66.280 249.500 ;
        RECT 65.980 248.300 66.280 248.750 ;
        RECT 65.980 247.550 66.280 248.000 ;
        RECT 65.980 246.800 66.280 247.250 ;
        RECT 65.980 246.050 66.280 246.500 ;
        RECT 65.980 245.300 66.280 245.750 ;
        RECT 83.180 254.300 83.480 254.750 ;
        RECT 83.180 253.550 83.480 254.000 ;
        RECT 83.180 252.800 83.480 253.250 ;
        RECT 83.180 252.050 83.480 252.500 ;
        RECT 83.180 251.300 83.480 251.750 ;
        RECT 83.180 250.550 83.480 251.000 ;
        RECT 83.180 249.800 83.480 250.250 ;
        RECT 83.180 249.050 83.480 249.500 ;
        RECT 83.180 248.300 83.480 248.750 ;
        RECT 83.180 247.550 83.480 248.000 ;
        RECT 83.180 246.800 83.480 247.250 ;
        RECT 83.180 246.050 83.480 246.500 ;
        RECT 83.180 245.300 83.480 245.750 ;
        RECT 85.980 254.300 86.280 254.750 ;
        RECT 85.980 253.550 86.280 254.000 ;
        RECT 85.980 252.800 86.280 253.250 ;
        RECT 85.980 252.050 86.280 252.500 ;
        RECT 85.980 251.300 86.280 251.750 ;
        RECT 85.980 250.550 86.280 251.000 ;
        RECT 85.980 249.800 86.280 250.250 ;
        RECT 85.980 249.050 86.280 249.500 ;
        RECT 85.980 248.300 86.280 248.750 ;
        RECT 85.980 247.550 86.280 248.000 ;
        RECT 85.980 246.800 86.280 247.250 ;
        RECT 85.980 246.050 86.280 246.500 ;
        RECT 85.980 245.300 86.280 245.750 ;
        RECT 103.180 254.300 103.480 254.750 ;
        RECT 103.180 253.550 103.480 254.000 ;
        RECT 103.180 252.800 103.480 253.250 ;
        RECT 103.180 252.050 103.480 252.500 ;
        RECT 103.180 251.300 103.480 251.750 ;
        RECT 103.180 250.550 103.480 251.000 ;
        RECT 103.180 249.800 103.480 250.250 ;
        RECT 103.180 249.050 103.480 249.500 ;
        RECT 103.180 248.300 103.480 248.750 ;
        RECT 103.180 247.550 103.480 248.000 ;
        RECT 103.180 246.800 103.480 247.250 ;
        RECT 103.180 246.050 103.480 246.500 ;
        RECT 103.180 245.300 103.480 245.750 ;
        RECT 5.980 234.300 6.280 234.750 ;
        RECT 5.980 233.550 6.280 234.000 ;
        RECT 5.980 232.800 6.280 233.250 ;
        RECT 5.980 232.050 6.280 232.500 ;
        RECT 5.980 231.300 6.280 231.750 ;
        RECT 5.980 230.550 6.280 231.000 ;
        RECT 5.980 229.800 6.280 230.250 ;
        RECT 5.980 229.050 6.280 229.500 ;
        RECT 5.980 228.300 6.280 228.750 ;
        RECT 5.980 227.550 6.280 228.000 ;
        RECT 5.980 226.800 6.280 227.250 ;
        RECT 5.980 226.050 6.280 226.500 ;
        RECT 5.980 225.300 6.280 225.750 ;
        RECT 23.180 234.300 23.480 234.750 ;
        RECT 23.180 233.550 23.480 234.000 ;
        RECT 23.180 232.800 23.480 233.250 ;
        RECT 23.180 232.050 23.480 232.500 ;
        RECT 23.180 231.300 23.480 231.750 ;
        RECT 23.180 230.550 23.480 231.000 ;
        RECT 23.180 229.800 23.480 230.250 ;
        RECT 23.180 229.050 23.480 229.500 ;
        RECT 23.180 228.300 23.480 228.750 ;
        RECT 23.180 227.550 23.480 228.000 ;
        RECT 23.180 226.800 23.480 227.250 ;
        RECT 23.180 226.050 23.480 226.500 ;
        RECT 23.180 225.300 23.480 225.750 ;
        RECT 25.980 234.300 26.280 234.750 ;
        RECT 25.980 233.550 26.280 234.000 ;
        RECT 25.980 232.800 26.280 233.250 ;
        RECT 25.980 232.050 26.280 232.500 ;
        RECT 25.980 231.300 26.280 231.750 ;
        RECT 25.980 230.550 26.280 231.000 ;
        RECT 25.980 229.800 26.280 230.250 ;
        RECT 25.980 229.050 26.280 229.500 ;
        RECT 25.980 228.300 26.280 228.750 ;
        RECT 25.980 227.550 26.280 228.000 ;
        RECT 25.980 226.800 26.280 227.250 ;
        RECT 25.980 226.050 26.280 226.500 ;
        RECT 25.980 225.300 26.280 225.750 ;
        RECT 43.180 234.300 43.480 234.750 ;
        RECT 43.180 233.550 43.480 234.000 ;
        RECT 43.180 232.800 43.480 233.250 ;
        RECT 43.180 232.050 43.480 232.500 ;
        RECT 43.180 231.300 43.480 231.750 ;
        RECT 43.180 230.550 43.480 231.000 ;
        RECT 43.180 229.800 43.480 230.250 ;
        RECT 43.180 229.050 43.480 229.500 ;
        RECT 43.180 228.300 43.480 228.750 ;
        RECT 43.180 227.550 43.480 228.000 ;
        RECT 43.180 226.800 43.480 227.250 ;
        RECT 43.180 226.050 43.480 226.500 ;
        RECT 43.180 225.300 43.480 225.750 ;
        RECT 45.980 234.300 46.280 234.750 ;
        RECT 45.980 233.550 46.280 234.000 ;
        RECT 45.980 232.800 46.280 233.250 ;
        RECT 45.980 232.050 46.280 232.500 ;
        RECT 45.980 231.300 46.280 231.750 ;
        RECT 45.980 230.550 46.280 231.000 ;
        RECT 45.980 229.800 46.280 230.250 ;
        RECT 45.980 229.050 46.280 229.500 ;
        RECT 45.980 228.300 46.280 228.750 ;
        RECT 45.980 227.550 46.280 228.000 ;
        RECT 45.980 226.800 46.280 227.250 ;
        RECT 45.980 226.050 46.280 226.500 ;
        RECT 45.980 225.300 46.280 225.750 ;
        RECT 63.180 234.300 63.480 234.750 ;
        RECT 63.180 233.550 63.480 234.000 ;
        RECT 63.180 232.800 63.480 233.250 ;
        RECT 63.180 232.050 63.480 232.500 ;
        RECT 63.180 231.300 63.480 231.750 ;
        RECT 63.180 230.550 63.480 231.000 ;
        RECT 63.180 229.800 63.480 230.250 ;
        RECT 63.180 229.050 63.480 229.500 ;
        RECT 63.180 228.300 63.480 228.750 ;
        RECT 63.180 227.550 63.480 228.000 ;
        RECT 63.180 226.800 63.480 227.250 ;
        RECT 63.180 226.050 63.480 226.500 ;
        RECT 63.180 225.300 63.480 225.750 ;
        RECT 65.980 234.300 66.280 234.750 ;
        RECT 65.980 233.550 66.280 234.000 ;
        RECT 65.980 232.800 66.280 233.250 ;
        RECT 65.980 232.050 66.280 232.500 ;
        RECT 65.980 231.300 66.280 231.750 ;
        RECT 65.980 230.550 66.280 231.000 ;
        RECT 65.980 229.800 66.280 230.250 ;
        RECT 65.980 229.050 66.280 229.500 ;
        RECT 65.980 228.300 66.280 228.750 ;
        RECT 65.980 227.550 66.280 228.000 ;
        RECT 65.980 226.800 66.280 227.250 ;
        RECT 65.980 226.050 66.280 226.500 ;
        RECT 65.980 225.300 66.280 225.750 ;
        RECT 83.180 234.300 83.480 234.750 ;
        RECT 83.180 233.550 83.480 234.000 ;
        RECT 83.180 232.800 83.480 233.250 ;
        RECT 83.180 232.050 83.480 232.500 ;
        RECT 83.180 231.300 83.480 231.750 ;
        RECT 83.180 230.550 83.480 231.000 ;
        RECT 83.180 229.800 83.480 230.250 ;
        RECT 83.180 229.050 83.480 229.500 ;
        RECT 83.180 228.300 83.480 228.750 ;
        RECT 83.180 227.550 83.480 228.000 ;
        RECT 83.180 226.800 83.480 227.250 ;
        RECT 83.180 226.050 83.480 226.500 ;
        RECT 83.180 225.300 83.480 225.750 ;
        RECT 85.980 234.300 86.280 234.750 ;
        RECT 85.980 233.550 86.280 234.000 ;
        RECT 85.980 232.800 86.280 233.250 ;
        RECT 85.980 232.050 86.280 232.500 ;
        RECT 85.980 231.300 86.280 231.750 ;
        RECT 85.980 230.550 86.280 231.000 ;
        RECT 85.980 229.800 86.280 230.250 ;
        RECT 85.980 229.050 86.280 229.500 ;
        RECT 85.980 228.300 86.280 228.750 ;
        RECT 85.980 227.550 86.280 228.000 ;
        RECT 85.980 226.800 86.280 227.250 ;
        RECT 85.980 226.050 86.280 226.500 ;
        RECT 85.980 225.300 86.280 225.750 ;
        RECT 103.180 234.300 103.480 234.750 ;
        RECT 103.180 233.550 103.480 234.000 ;
        RECT 103.180 232.800 103.480 233.250 ;
        RECT 103.180 232.050 103.480 232.500 ;
        RECT 103.180 231.300 103.480 231.750 ;
        RECT 103.180 230.550 103.480 231.000 ;
        RECT 103.180 229.800 103.480 230.250 ;
        RECT 103.180 229.050 103.480 229.500 ;
        RECT 103.180 228.300 103.480 228.750 ;
        RECT 103.180 227.550 103.480 228.000 ;
        RECT 103.180 226.800 103.480 227.250 ;
        RECT 103.180 226.050 103.480 226.500 ;
        RECT 103.180 225.300 103.480 225.750 ;
        RECT 9.425 196.405 10.015 196.975 ;
        RECT 10.205 196.405 10.795 196.975 ;
        RECT 10.985 196.405 11.575 196.975 ;
        RECT 10.175 194.445 10.345 194.720 ;
        RECT 11.755 194.445 11.925 194.720 ;
        RECT 12.395 194.445 12.570 194.745 ;
        RECT 13.985 194.450 14.155 194.745 ;
        RECT 5.980 154.300 6.280 154.750 ;
        RECT 5.980 153.550 6.280 154.000 ;
        RECT 5.980 152.800 6.280 153.250 ;
        RECT 5.980 152.050 6.280 152.500 ;
        RECT 5.980 151.300 6.280 151.750 ;
        RECT 5.980 150.550 6.280 151.000 ;
        RECT 5.980 149.800 6.280 150.250 ;
        RECT 5.980 149.050 6.280 149.500 ;
        RECT 5.980 148.300 6.280 148.750 ;
        RECT 5.980 147.550 6.280 148.000 ;
        RECT 5.980 146.800 6.280 147.250 ;
        RECT 5.980 146.050 6.280 146.500 ;
        RECT 5.980 145.300 6.280 145.750 ;
        RECT 23.180 154.300 23.480 154.750 ;
        RECT 23.180 153.550 23.480 154.000 ;
        RECT 23.180 152.800 23.480 153.250 ;
        RECT 23.180 152.050 23.480 152.500 ;
        RECT 23.180 151.300 23.480 151.750 ;
        RECT 23.180 150.550 23.480 151.000 ;
        RECT 23.180 149.800 23.480 150.250 ;
        RECT 23.180 149.050 23.480 149.500 ;
        RECT 23.180 148.300 23.480 148.750 ;
        RECT 23.180 147.550 23.480 148.000 ;
        RECT 23.180 146.800 23.480 147.250 ;
        RECT 23.180 146.050 23.480 146.500 ;
        RECT 23.180 145.300 23.480 145.750 ;
        RECT 25.980 154.300 26.280 154.750 ;
        RECT 25.980 153.550 26.280 154.000 ;
        RECT 25.980 152.800 26.280 153.250 ;
        RECT 25.980 152.050 26.280 152.500 ;
        RECT 25.980 151.300 26.280 151.750 ;
        RECT 25.980 150.550 26.280 151.000 ;
        RECT 25.980 149.800 26.280 150.250 ;
        RECT 25.980 149.050 26.280 149.500 ;
        RECT 25.980 148.300 26.280 148.750 ;
        RECT 25.980 147.550 26.280 148.000 ;
        RECT 25.980 146.800 26.280 147.250 ;
        RECT 25.980 146.050 26.280 146.500 ;
        RECT 25.980 145.300 26.280 145.750 ;
        RECT 43.180 154.300 43.480 154.750 ;
        RECT 43.180 153.550 43.480 154.000 ;
        RECT 43.180 152.800 43.480 153.250 ;
        RECT 43.180 152.050 43.480 152.500 ;
        RECT 43.180 151.300 43.480 151.750 ;
        RECT 43.180 150.550 43.480 151.000 ;
        RECT 43.180 149.800 43.480 150.250 ;
        RECT 43.180 149.050 43.480 149.500 ;
        RECT 43.180 148.300 43.480 148.750 ;
        RECT 43.180 147.550 43.480 148.000 ;
        RECT 43.180 146.800 43.480 147.250 ;
        RECT 43.180 146.050 43.480 146.500 ;
        RECT 43.180 145.300 43.480 145.750 ;
        RECT 45.980 154.300 46.280 154.750 ;
        RECT 45.980 153.550 46.280 154.000 ;
        RECT 45.980 152.800 46.280 153.250 ;
        RECT 45.980 152.050 46.280 152.500 ;
        RECT 45.980 151.300 46.280 151.750 ;
        RECT 45.980 150.550 46.280 151.000 ;
        RECT 45.980 149.800 46.280 150.250 ;
        RECT 45.980 149.050 46.280 149.500 ;
        RECT 45.980 148.300 46.280 148.750 ;
        RECT 45.980 147.550 46.280 148.000 ;
        RECT 45.980 146.800 46.280 147.250 ;
        RECT 45.980 146.050 46.280 146.500 ;
        RECT 45.980 145.300 46.280 145.750 ;
        RECT 63.180 154.300 63.480 154.750 ;
        RECT 63.180 153.550 63.480 154.000 ;
        RECT 63.180 152.800 63.480 153.250 ;
        RECT 63.180 152.050 63.480 152.500 ;
        RECT 63.180 151.300 63.480 151.750 ;
        RECT 63.180 150.550 63.480 151.000 ;
        RECT 63.180 149.800 63.480 150.250 ;
        RECT 63.180 149.050 63.480 149.500 ;
        RECT 63.180 148.300 63.480 148.750 ;
        RECT 63.180 147.550 63.480 148.000 ;
        RECT 63.180 146.800 63.480 147.250 ;
        RECT 63.180 146.050 63.480 146.500 ;
        RECT 63.180 145.300 63.480 145.750 ;
        RECT 65.980 154.300 66.280 154.750 ;
        RECT 65.980 153.550 66.280 154.000 ;
        RECT 65.980 152.800 66.280 153.250 ;
        RECT 65.980 152.050 66.280 152.500 ;
        RECT 65.980 151.300 66.280 151.750 ;
        RECT 65.980 150.550 66.280 151.000 ;
        RECT 65.980 149.800 66.280 150.250 ;
        RECT 65.980 149.050 66.280 149.500 ;
        RECT 65.980 148.300 66.280 148.750 ;
        RECT 65.980 147.550 66.280 148.000 ;
        RECT 65.980 146.800 66.280 147.250 ;
        RECT 65.980 146.050 66.280 146.500 ;
        RECT 65.980 145.300 66.280 145.750 ;
        RECT 83.180 154.300 83.480 154.750 ;
        RECT 83.180 153.550 83.480 154.000 ;
        RECT 83.180 152.800 83.480 153.250 ;
        RECT 83.180 152.050 83.480 152.500 ;
        RECT 83.180 151.300 83.480 151.750 ;
        RECT 83.180 150.550 83.480 151.000 ;
        RECT 83.180 149.800 83.480 150.250 ;
        RECT 83.180 149.050 83.480 149.500 ;
        RECT 83.180 148.300 83.480 148.750 ;
        RECT 83.180 147.550 83.480 148.000 ;
        RECT 83.180 146.800 83.480 147.250 ;
        RECT 83.180 146.050 83.480 146.500 ;
        RECT 83.180 145.300 83.480 145.750 ;
        RECT 85.980 154.300 86.280 154.750 ;
        RECT 85.980 153.550 86.280 154.000 ;
        RECT 85.980 152.800 86.280 153.250 ;
        RECT 85.980 152.050 86.280 152.500 ;
        RECT 85.980 151.300 86.280 151.750 ;
        RECT 85.980 150.550 86.280 151.000 ;
        RECT 85.980 149.800 86.280 150.250 ;
        RECT 85.980 149.050 86.280 149.500 ;
        RECT 85.980 148.300 86.280 148.750 ;
        RECT 85.980 147.550 86.280 148.000 ;
        RECT 85.980 146.800 86.280 147.250 ;
        RECT 85.980 146.050 86.280 146.500 ;
        RECT 85.980 145.300 86.280 145.750 ;
        RECT 103.180 154.300 103.480 154.750 ;
        RECT 103.180 153.550 103.480 154.000 ;
        RECT 103.180 152.800 103.480 153.250 ;
        RECT 103.180 152.050 103.480 152.500 ;
        RECT 103.180 151.300 103.480 151.750 ;
        RECT 103.180 150.550 103.480 151.000 ;
        RECT 103.180 149.800 103.480 150.250 ;
        RECT 103.180 149.050 103.480 149.500 ;
        RECT 103.180 148.300 103.480 148.750 ;
        RECT 103.180 147.550 103.480 148.000 ;
        RECT 103.180 146.800 103.480 147.250 ;
        RECT 103.180 146.050 103.480 146.500 ;
        RECT 103.180 145.300 103.480 145.750 ;
        RECT 5.980 134.300 6.280 134.750 ;
        RECT 5.980 133.550 6.280 134.000 ;
        RECT 5.980 132.800 6.280 133.250 ;
        RECT 5.980 132.050 6.280 132.500 ;
        RECT 5.980 131.300 6.280 131.750 ;
        RECT 5.980 130.550 6.280 131.000 ;
        RECT 5.980 129.800 6.280 130.250 ;
        RECT 5.980 129.050 6.280 129.500 ;
        RECT 5.980 128.300 6.280 128.750 ;
        RECT 5.980 127.550 6.280 128.000 ;
        RECT 5.980 126.800 6.280 127.250 ;
        RECT 5.980 126.050 6.280 126.500 ;
        RECT 5.980 125.300 6.280 125.750 ;
        RECT 23.180 134.300 23.480 134.750 ;
        RECT 23.180 133.550 23.480 134.000 ;
        RECT 23.180 132.800 23.480 133.250 ;
        RECT 23.180 132.050 23.480 132.500 ;
        RECT 23.180 131.300 23.480 131.750 ;
        RECT 23.180 130.550 23.480 131.000 ;
        RECT 23.180 129.800 23.480 130.250 ;
        RECT 23.180 129.050 23.480 129.500 ;
        RECT 23.180 128.300 23.480 128.750 ;
        RECT 23.180 127.550 23.480 128.000 ;
        RECT 23.180 126.800 23.480 127.250 ;
        RECT 23.180 126.050 23.480 126.500 ;
        RECT 23.180 125.300 23.480 125.750 ;
        RECT 25.980 134.300 26.280 134.750 ;
        RECT 25.980 133.550 26.280 134.000 ;
        RECT 25.980 132.800 26.280 133.250 ;
        RECT 25.980 132.050 26.280 132.500 ;
        RECT 25.980 131.300 26.280 131.750 ;
        RECT 25.980 130.550 26.280 131.000 ;
        RECT 25.980 129.800 26.280 130.250 ;
        RECT 25.980 129.050 26.280 129.500 ;
        RECT 25.980 128.300 26.280 128.750 ;
        RECT 25.980 127.550 26.280 128.000 ;
        RECT 25.980 126.800 26.280 127.250 ;
        RECT 25.980 126.050 26.280 126.500 ;
        RECT 25.980 125.300 26.280 125.750 ;
        RECT 43.180 134.300 43.480 134.750 ;
        RECT 43.180 133.550 43.480 134.000 ;
        RECT 43.180 132.800 43.480 133.250 ;
        RECT 43.180 132.050 43.480 132.500 ;
        RECT 43.180 131.300 43.480 131.750 ;
        RECT 43.180 130.550 43.480 131.000 ;
        RECT 43.180 129.800 43.480 130.250 ;
        RECT 43.180 129.050 43.480 129.500 ;
        RECT 43.180 128.300 43.480 128.750 ;
        RECT 43.180 127.550 43.480 128.000 ;
        RECT 43.180 126.800 43.480 127.250 ;
        RECT 43.180 126.050 43.480 126.500 ;
        RECT 43.180 125.300 43.480 125.750 ;
        RECT 45.980 134.300 46.280 134.750 ;
        RECT 45.980 133.550 46.280 134.000 ;
        RECT 45.980 132.800 46.280 133.250 ;
        RECT 45.980 132.050 46.280 132.500 ;
        RECT 45.980 131.300 46.280 131.750 ;
        RECT 45.980 130.550 46.280 131.000 ;
        RECT 45.980 129.800 46.280 130.250 ;
        RECT 45.980 129.050 46.280 129.500 ;
        RECT 45.980 128.300 46.280 128.750 ;
        RECT 45.980 127.550 46.280 128.000 ;
        RECT 45.980 126.800 46.280 127.250 ;
        RECT 45.980 126.050 46.280 126.500 ;
        RECT 45.980 125.300 46.280 125.750 ;
        RECT 63.180 134.300 63.480 134.750 ;
        RECT 63.180 133.550 63.480 134.000 ;
        RECT 63.180 132.800 63.480 133.250 ;
        RECT 63.180 132.050 63.480 132.500 ;
        RECT 63.180 131.300 63.480 131.750 ;
        RECT 63.180 130.550 63.480 131.000 ;
        RECT 63.180 129.800 63.480 130.250 ;
        RECT 63.180 129.050 63.480 129.500 ;
        RECT 63.180 128.300 63.480 128.750 ;
        RECT 63.180 127.550 63.480 128.000 ;
        RECT 63.180 126.800 63.480 127.250 ;
        RECT 63.180 126.050 63.480 126.500 ;
        RECT 63.180 125.300 63.480 125.750 ;
        RECT 65.980 134.300 66.280 134.750 ;
        RECT 65.980 133.550 66.280 134.000 ;
        RECT 65.980 132.800 66.280 133.250 ;
        RECT 65.980 132.050 66.280 132.500 ;
        RECT 65.980 131.300 66.280 131.750 ;
        RECT 65.980 130.550 66.280 131.000 ;
        RECT 65.980 129.800 66.280 130.250 ;
        RECT 65.980 129.050 66.280 129.500 ;
        RECT 65.980 128.300 66.280 128.750 ;
        RECT 65.980 127.550 66.280 128.000 ;
        RECT 65.980 126.800 66.280 127.250 ;
        RECT 65.980 126.050 66.280 126.500 ;
        RECT 65.980 125.300 66.280 125.750 ;
        RECT 83.180 134.300 83.480 134.750 ;
        RECT 83.180 133.550 83.480 134.000 ;
        RECT 83.180 132.800 83.480 133.250 ;
        RECT 83.180 132.050 83.480 132.500 ;
        RECT 83.180 131.300 83.480 131.750 ;
        RECT 83.180 130.550 83.480 131.000 ;
        RECT 83.180 129.800 83.480 130.250 ;
        RECT 83.180 129.050 83.480 129.500 ;
        RECT 83.180 128.300 83.480 128.750 ;
        RECT 83.180 127.550 83.480 128.000 ;
        RECT 83.180 126.800 83.480 127.250 ;
        RECT 83.180 126.050 83.480 126.500 ;
        RECT 83.180 125.300 83.480 125.750 ;
        RECT 85.980 134.300 86.280 134.750 ;
        RECT 85.980 133.550 86.280 134.000 ;
        RECT 85.980 132.800 86.280 133.250 ;
        RECT 85.980 132.050 86.280 132.500 ;
        RECT 85.980 131.300 86.280 131.750 ;
        RECT 85.980 130.550 86.280 131.000 ;
        RECT 85.980 129.800 86.280 130.250 ;
        RECT 85.980 129.050 86.280 129.500 ;
        RECT 85.980 128.300 86.280 128.750 ;
        RECT 85.980 127.550 86.280 128.000 ;
        RECT 85.980 126.800 86.280 127.250 ;
        RECT 85.980 126.050 86.280 126.500 ;
        RECT 85.980 125.300 86.280 125.750 ;
        RECT 103.180 134.300 103.480 134.750 ;
        RECT 103.180 133.550 103.480 134.000 ;
        RECT 103.180 132.800 103.480 133.250 ;
        RECT 103.180 132.050 103.480 132.500 ;
        RECT 103.180 131.300 103.480 131.750 ;
        RECT 103.180 130.550 103.480 131.000 ;
        RECT 103.180 129.800 103.480 130.250 ;
        RECT 103.180 129.050 103.480 129.500 ;
        RECT 103.180 128.300 103.480 128.750 ;
        RECT 103.180 127.550 103.480 128.000 ;
        RECT 103.180 126.800 103.480 127.250 ;
        RECT 103.180 126.050 103.480 126.500 ;
        RECT 103.180 125.300 103.480 125.750 ;
        RECT 5.980 114.300 6.280 114.750 ;
        RECT 5.980 113.550 6.280 114.000 ;
        RECT 5.980 112.800 6.280 113.250 ;
        RECT 5.980 112.050 6.280 112.500 ;
        RECT 5.980 111.300 6.280 111.750 ;
        RECT 5.980 110.550 6.280 111.000 ;
        RECT 5.980 109.800 6.280 110.250 ;
        RECT 5.980 109.050 6.280 109.500 ;
        RECT 5.980 108.300 6.280 108.750 ;
        RECT 5.980 107.550 6.280 108.000 ;
        RECT 5.980 106.800 6.280 107.250 ;
        RECT 5.980 106.050 6.280 106.500 ;
        RECT 5.980 105.300 6.280 105.750 ;
        RECT 23.180 114.300 23.480 114.750 ;
        RECT 23.180 113.550 23.480 114.000 ;
        RECT 23.180 112.800 23.480 113.250 ;
        RECT 23.180 112.050 23.480 112.500 ;
        RECT 23.180 111.300 23.480 111.750 ;
        RECT 23.180 110.550 23.480 111.000 ;
        RECT 23.180 109.800 23.480 110.250 ;
        RECT 23.180 109.050 23.480 109.500 ;
        RECT 23.180 108.300 23.480 108.750 ;
        RECT 23.180 107.550 23.480 108.000 ;
        RECT 23.180 106.800 23.480 107.250 ;
        RECT 23.180 106.050 23.480 106.500 ;
        RECT 23.180 105.300 23.480 105.750 ;
        RECT 25.980 114.300 26.280 114.750 ;
        RECT 25.980 113.550 26.280 114.000 ;
        RECT 25.980 112.800 26.280 113.250 ;
        RECT 25.980 112.050 26.280 112.500 ;
        RECT 25.980 111.300 26.280 111.750 ;
        RECT 25.980 110.550 26.280 111.000 ;
        RECT 25.980 109.800 26.280 110.250 ;
        RECT 25.980 109.050 26.280 109.500 ;
        RECT 25.980 108.300 26.280 108.750 ;
        RECT 25.980 107.550 26.280 108.000 ;
        RECT 25.980 106.800 26.280 107.250 ;
        RECT 25.980 106.050 26.280 106.500 ;
        RECT 25.980 105.300 26.280 105.750 ;
        RECT 43.180 114.300 43.480 114.750 ;
        RECT 43.180 113.550 43.480 114.000 ;
        RECT 43.180 112.800 43.480 113.250 ;
        RECT 43.180 112.050 43.480 112.500 ;
        RECT 43.180 111.300 43.480 111.750 ;
        RECT 43.180 110.550 43.480 111.000 ;
        RECT 43.180 109.800 43.480 110.250 ;
        RECT 43.180 109.050 43.480 109.500 ;
        RECT 43.180 108.300 43.480 108.750 ;
        RECT 43.180 107.550 43.480 108.000 ;
        RECT 43.180 106.800 43.480 107.250 ;
        RECT 43.180 106.050 43.480 106.500 ;
        RECT 43.180 105.300 43.480 105.750 ;
        RECT 45.980 114.300 46.280 114.750 ;
        RECT 45.980 113.550 46.280 114.000 ;
        RECT 45.980 112.800 46.280 113.250 ;
        RECT 45.980 112.050 46.280 112.500 ;
        RECT 45.980 111.300 46.280 111.750 ;
        RECT 45.980 110.550 46.280 111.000 ;
        RECT 45.980 109.800 46.280 110.250 ;
        RECT 45.980 109.050 46.280 109.500 ;
        RECT 45.980 108.300 46.280 108.750 ;
        RECT 45.980 107.550 46.280 108.000 ;
        RECT 45.980 106.800 46.280 107.250 ;
        RECT 45.980 106.050 46.280 106.500 ;
        RECT 45.980 105.300 46.280 105.750 ;
        RECT 63.180 114.300 63.480 114.750 ;
        RECT 63.180 113.550 63.480 114.000 ;
        RECT 63.180 112.800 63.480 113.250 ;
        RECT 63.180 112.050 63.480 112.500 ;
        RECT 63.180 111.300 63.480 111.750 ;
        RECT 63.180 110.550 63.480 111.000 ;
        RECT 63.180 109.800 63.480 110.250 ;
        RECT 63.180 109.050 63.480 109.500 ;
        RECT 63.180 108.300 63.480 108.750 ;
        RECT 63.180 107.550 63.480 108.000 ;
        RECT 63.180 106.800 63.480 107.250 ;
        RECT 63.180 106.050 63.480 106.500 ;
        RECT 63.180 105.300 63.480 105.750 ;
        RECT 65.980 114.300 66.280 114.750 ;
        RECT 65.980 113.550 66.280 114.000 ;
        RECT 65.980 112.800 66.280 113.250 ;
        RECT 65.980 112.050 66.280 112.500 ;
        RECT 65.980 111.300 66.280 111.750 ;
        RECT 65.980 110.550 66.280 111.000 ;
        RECT 65.980 109.800 66.280 110.250 ;
        RECT 65.980 109.050 66.280 109.500 ;
        RECT 65.980 108.300 66.280 108.750 ;
        RECT 65.980 107.550 66.280 108.000 ;
        RECT 65.980 106.800 66.280 107.250 ;
        RECT 65.980 106.050 66.280 106.500 ;
        RECT 65.980 105.300 66.280 105.750 ;
        RECT 83.180 114.300 83.480 114.750 ;
        RECT 83.180 113.550 83.480 114.000 ;
        RECT 83.180 112.800 83.480 113.250 ;
        RECT 83.180 112.050 83.480 112.500 ;
        RECT 83.180 111.300 83.480 111.750 ;
        RECT 83.180 110.550 83.480 111.000 ;
        RECT 83.180 109.800 83.480 110.250 ;
        RECT 83.180 109.050 83.480 109.500 ;
        RECT 83.180 108.300 83.480 108.750 ;
        RECT 83.180 107.550 83.480 108.000 ;
        RECT 83.180 106.800 83.480 107.250 ;
        RECT 83.180 106.050 83.480 106.500 ;
        RECT 83.180 105.300 83.480 105.750 ;
        RECT 85.980 114.300 86.280 114.750 ;
        RECT 85.980 113.550 86.280 114.000 ;
        RECT 85.980 112.800 86.280 113.250 ;
        RECT 85.980 112.050 86.280 112.500 ;
        RECT 85.980 111.300 86.280 111.750 ;
        RECT 85.980 110.550 86.280 111.000 ;
        RECT 85.980 109.800 86.280 110.250 ;
        RECT 85.980 109.050 86.280 109.500 ;
        RECT 85.980 108.300 86.280 108.750 ;
        RECT 85.980 107.550 86.280 108.000 ;
        RECT 85.980 106.800 86.280 107.250 ;
        RECT 85.980 106.050 86.280 106.500 ;
        RECT 85.980 105.300 86.280 105.750 ;
        RECT 103.180 114.300 103.480 114.750 ;
        RECT 103.180 113.550 103.480 114.000 ;
        RECT 103.180 112.800 103.480 113.250 ;
        RECT 103.180 112.050 103.480 112.500 ;
        RECT 103.180 111.300 103.480 111.750 ;
        RECT 103.180 110.550 103.480 111.000 ;
        RECT 103.180 109.800 103.480 110.250 ;
        RECT 103.180 109.050 103.480 109.500 ;
        RECT 103.180 108.300 103.480 108.750 ;
        RECT 103.180 107.550 103.480 108.000 ;
        RECT 103.180 106.800 103.480 107.250 ;
        RECT 103.180 106.050 103.480 106.500 ;
        RECT 103.180 105.300 103.480 105.750 ;
        RECT 5.980 94.300 6.280 94.750 ;
        RECT 5.980 93.550 6.280 94.000 ;
        RECT 5.980 92.800 6.280 93.250 ;
        RECT 5.980 92.050 6.280 92.500 ;
        RECT 5.980 91.300 6.280 91.750 ;
        RECT 5.980 90.550 6.280 91.000 ;
        RECT 5.980 89.800 6.280 90.250 ;
        RECT 5.980 89.050 6.280 89.500 ;
        RECT 5.980 88.300 6.280 88.750 ;
        RECT 5.980 87.550 6.280 88.000 ;
        RECT 5.980 86.800 6.280 87.250 ;
        RECT 5.980 86.050 6.280 86.500 ;
        RECT 5.980 85.300 6.280 85.750 ;
        RECT 23.180 94.300 23.480 94.750 ;
        RECT 23.180 93.550 23.480 94.000 ;
        RECT 23.180 92.800 23.480 93.250 ;
        RECT 23.180 92.050 23.480 92.500 ;
        RECT 23.180 91.300 23.480 91.750 ;
        RECT 23.180 90.550 23.480 91.000 ;
        RECT 23.180 89.800 23.480 90.250 ;
        RECT 23.180 89.050 23.480 89.500 ;
        RECT 23.180 88.300 23.480 88.750 ;
        RECT 23.180 87.550 23.480 88.000 ;
        RECT 23.180 86.800 23.480 87.250 ;
        RECT 23.180 86.050 23.480 86.500 ;
        RECT 23.180 85.300 23.480 85.750 ;
        RECT 25.980 94.300 26.280 94.750 ;
        RECT 25.980 93.550 26.280 94.000 ;
        RECT 25.980 92.800 26.280 93.250 ;
        RECT 25.980 92.050 26.280 92.500 ;
        RECT 25.980 91.300 26.280 91.750 ;
        RECT 25.980 90.550 26.280 91.000 ;
        RECT 25.980 89.800 26.280 90.250 ;
        RECT 25.980 89.050 26.280 89.500 ;
        RECT 25.980 88.300 26.280 88.750 ;
        RECT 25.980 87.550 26.280 88.000 ;
        RECT 25.980 86.800 26.280 87.250 ;
        RECT 25.980 86.050 26.280 86.500 ;
        RECT 25.980 85.300 26.280 85.750 ;
        RECT 43.180 94.300 43.480 94.750 ;
        RECT 43.180 93.550 43.480 94.000 ;
        RECT 43.180 92.800 43.480 93.250 ;
        RECT 43.180 92.050 43.480 92.500 ;
        RECT 43.180 91.300 43.480 91.750 ;
        RECT 43.180 90.550 43.480 91.000 ;
        RECT 43.180 89.800 43.480 90.250 ;
        RECT 43.180 89.050 43.480 89.500 ;
        RECT 43.180 88.300 43.480 88.750 ;
        RECT 43.180 87.550 43.480 88.000 ;
        RECT 43.180 86.800 43.480 87.250 ;
        RECT 43.180 86.050 43.480 86.500 ;
        RECT 43.180 85.300 43.480 85.750 ;
        RECT 45.980 94.300 46.280 94.750 ;
        RECT 45.980 93.550 46.280 94.000 ;
        RECT 45.980 92.800 46.280 93.250 ;
        RECT 45.980 92.050 46.280 92.500 ;
        RECT 45.980 91.300 46.280 91.750 ;
        RECT 45.980 90.550 46.280 91.000 ;
        RECT 45.980 89.800 46.280 90.250 ;
        RECT 45.980 89.050 46.280 89.500 ;
        RECT 45.980 88.300 46.280 88.750 ;
        RECT 45.980 87.550 46.280 88.000 ;
        RECT 45.980 86.800 46.280 87.250 ;
        RECT 45.980 86.050 46.280 86.500 ;
        RECT 45.980 85.300 46.280 85.750 ;
        RECT 63.180 94.300 63.480 94.750 ;
        RECT 63.180 93.550 63.480 94.000 ;
        RECT 63.180 92.800 63.480 93.250 ;
        RECT 63.180 92.050 63.480 92.500 ;
        RECT 63.180 91.300 63.480 91.750 ;
        RECT 63.180 90.550 63.480 91.000 ;
        RECT 63.180 89.800 63.480 90.250 ;
        RECT 63.180 89.050 63.480 89.500 ;
        RECT 63.180 88.300 63.480 88.750 ;
        RECT 63.180 87.550 63.480 88.000 ;
        RECT 63.180 86.800 63.480 87.250 ;
        RECT 63.180 86.050 63.480 86.500 ;
        RECT 63.180 85.300 63.480 85.750 ;
        RECT 65.980 94.300 66.280 94.750 ;
        RECT 65.980 93.550 66.280 94.000 ;
        RECT 65.980 92.800 66.280 93.250 ;
        RECT 65.980 92.050 66.280 92.500 ;
        RECT 65.980 91.300 66.280 91.750 ;
        RECT 65.980 90.550 66.280 91.000 ;
        RECT 65.980 89.800 66.280 90.250 ;
        RECT 65.980 89.050 66.280 89.500 ;
        RECT 65.980 88.300 66.280 88.750 ;
        RECT 65.980 87.550 66.280 88.000 ;
        RECT 65.980 86.800 66.280 87.250 ;
        RECT 65.980 86.050 66.280 86.500 ;
        RECT 65.980 85.300 66.280 85.750 ;
        RECT 83.180 94.300 83.480 94.750 ;
        RECT 83.180 93.550 83.480 94.000 ;
        RECT 83.180 92.800 83.480 93.250 ;
        RECT 83.180 92.050 83.480 92.500 ;
        RECT 83.180 91.300 83.480 91.750 ;
        RECT 83.180 90.550 83.480 91.000 ;
        RECT 83.180 89.800 83.480 90.250 ;
        RECT 83.180 89.050 83.480 89.500 ;
        RECT 83.180 88.300 83.480 88.750 ;
        RECT 83.180 87.550 83.480 88.000 ;
        RECT 83.180 86.800 83.480 87.250 ;
        RECT 83.180 86.050 83.480 86.500 ;
        RECT 83.180 85.300 83.480 85.750 ;
        RECT 85.980 94.300 86.280 94.750 ;
        RECT 85.980 93.550 86.280 94.000 ;
        RECT 85.980 92.800 86.280 93.250 ;
        RECT 85.980 92.050 86.280 92.500 ;
        RECT 85.980 91.300 86.280 91.750 ;
        RECT 85.980 90.550 86.280 91.000 ;
        RECT 85.980 89.800 86.280 90.250 ;
        RECT 85.980 89.050 86.280 89.500 ;
        RECT 85.980 88.300 86.280 88.750 ;
        RECT 85.980 87.550 86.280 88.000 ;
        RECT 85.980 86.800 86.280 87.250 ;
        RECT 85.980 86.050 86.280 86.500 ;
        RECT 85.980 85.300 86.280 85.750 ;
        RECT 103.180 94.300 103.480 94.750 ;
        RECT 103.180 93.550 103.480 94.000 ;
        RECT 103.180 92.800 103.480 93.250 ;
        RECT 103.180 92.050 103.480 92.500 ;
        RECT 103.180 91.300 103.480 91.750 ;
        RECT 103.180 90.550 103.480 91.000 ;
        RECT 103.180 89.800 103.480 90.250 ;
        RECT 103.180 89.050 103.480 89.500 ;
        RECT 103.180 88.300 103.480 88.750 ;
        RECT 103.180 87.550 103.480 88.000 ;
        RECT 103.180 86.800 103.480 87.250 ;
        RECT 103.180 86.050 103.480 86.500 ;
        RECT 103.180 85.300 103.480 85.750 ;
        RECT 5.980 74.300 6.280 74.750 ;
        RECT 5.980 73.550 6.280 74.000 ;
        RECT 5.980 72.800 6.280 73.250 ;
        RECT 5.980 72.050 6.280 72.500 ;
        RECT 5.980 71.300 6.280 71.750 ;
        RECT 5.980 70.550 6.280 71.000 ;
        RECT 5.980 69.800 6.280 70.250 ;
        RECT 5.980 69.050 6.280 69.500 ;
        RECT 5.980 68.300 6.280 68.750 ;
        RECT 5.980 67.550 6.280 68.000 ;
        RECT 5.980 66.800 6.280 67.250 ;
        RECT 5.980 66.050 6.280 66.500 ;
        RECT 5.980 65.300 6.280 65.750 ;
        RECT 23.180 74.300 23.480 74.750 ;
        RECT 23.180 73.550 23.480 74.000 ;
        RECT 23.180 72.800 23.480 73.250 ;
        RECT 23.180 72.050 23.480 72.500 ;
        RECT 23.180 71.300 23.480 71.750 ;
        RECT 23.180 70.550 23.480 71.000 ;
        RECT 23.180 69.800 23.480 70.250 ;
        RECT 23.180 69.050 23.480 69.500 ;
        RECT 23.180 68.300 23.480 68.750 ;
        RECT 23.180 67.550 23.480 68.000 ;
        RECT 23.180 66.800 23.480 67.250 ;
        RECT 23.180 66.050 23.480 66.500 ;
        RECT 23.180 65.300 23.480 65.750 ;
        RECT 25.980 74.300 26.280 74.750 ;
        RECT 25.980 73.550 26.280 74.000 ;
        RECT 25.980 72.800 26.280 73.250 ;
        RECT 25.980 72.050 26.280 72.500 ;
        RECT 25.980 71.300 26.280 71.750 ;
        RECT 25.980 70.550 26.280 71.000 ;
        RECT 25.980 69.800 26.280 70.250 ;
        RECT 25.980 69.050 26.280 69.500 ;
        RECT 25.980 68.300 26.280 68.750 ;
        RECT 25.980 67.550 26.280 68.000 ;
        RECT 25.980 66.800 26.280 67.250 ;
        RECT 25.980 66.050 26.280 66.500 ;
        RECT 25.980 65.300 26.280 65.750 ;
        RECT 43.180 74.300 43.480 74.750 ;
        RECT 43.180 73.550 43.480 74.000 ;
        RECT 43.180 72.800 43.480 73.250 ;
        RECT 43.180 72.050 43.480 72.500 ;
        RECT 43.180 71.300 43.480 71.750 ;
        RECT 43.180 70.550 43.480 71.000 ;
        RECT 43.180 69.800 43.480 70.250 ;
        RECT 43.180 69.050 43.480 69.500 ;
        RECT 43.180 68.300 43.480 68.750 ;
        RECT 43.180 67.550 43.480 68.000 ;
        RECT 43.180 66.800 43.480 67.250 ;
        RECT 43.180 66.050 43.480 66.500 ;
        RECT 43.180 65.300 43.480 65.750 ;
        RECT 45.980 74.300 46.280 74.750 ;
        RECT 45.980 73.550 46.280 74.000 ;
        RECT 45.980 72.800 46.280 73.250 ;
        RECT 45.980 72.050 46.280 72.500 ;
        RECT 45.980 71.300 46.280 71.750 ;
        RECT 45.980 70.550 46.280 71.000 ;
        RECT 45.980 69.800 46.280 70.250 ;
        RECT 45.980 69.050 46.280 69.500 ;
        RECT 45.980 68.300 46.280 68.750 ;
        RECT 45.980 67.550 46.280 68.000 ;
        RECT 45.980 66.800 46.280 67.250 ;
        RECT 45.980 66.050 46.280 66.500 ;
        RECT 45.980 65.300 46.280 65.750 ;
        RECT 63.180 74.300 63.480 74.750 ;
        RECT 63.180 73.550 63.480 74.000 ;
        RECT 63.180 72.800 63.480 73.250 ;
        RECT 63.180 72.050 63.480 72.500 ;
        RECT 63.180 71.300 63.480 71.750 ;
        RECT 63.180 70.550 63.480 71.000 ;
        RECT 63.180 69.800 63.480 70.250 ;
        RECT 63.180 69.050 63.480 69.500 ;
        RECT 63.180 68.300 63.480 68.750 ;
        RECT 63.180 67.550 63.480 68.000 ;
        RECT 63.180 66.800 63.480 67.250 ;
        RECT 63.180 66.050 63.480 66.500 ;
        RECT 63.180 65.300 63.480 65.750 ;
        RECT 65.980 74.300 66.280 74.750 ;
        RECT 65.980 73.550 66.280 74.000 ;
        RECT 65.980 72.800 66.280 73.250 ;
        RECT 65.980 72.050 66.280 72.500 ;
        RECT 65.980 71.300 66.280 71.750 ;
        RECT 65.980 70.550 66.280 71.000 ;
        RECT 65.980 69.800 66.280 70.250 ;
        RECT 65.980 69.050 66.280 69.500 ;
        RECT 65.980 68.300 66.280 68.750 ;
        RECT 65.980 67.550 66.280 68.000 ;
        RECT 65.980 66.800 66.280 67.250 ;
        RECT 65.980 66.050 66.280 66.500 ;
        RECT 65.980 65.300 66.280 65.750 ;
        RECT 83.180 74.300 83.480 74.750 ;
        RECT 83.180 73.550 83.480 74.000 ;
        RECT 83.180 72.800 83.480 73.250 ;
        RECT 83.180 72.050 83.480 72.500 ;
        RECT 83.180 71.300 83.480 71.750 ;
        RECT 83.180 70.550 83.480 71.000 ;
        RECT 83.180 69.800 83.480 70.250 ;
        RECT 83.180 69.050 83.480 69.500 ;
        RECT 83.180 68.300 83.480 68.750 ;
        RECT 83.180 67.550 83.480 68.000 ;
        RECT 83.180 66.800 83.480 67.250 ;
        RECT 83.180 66.050 83.480 66.500 ;
        RECT 83.180 65.300 83.480 65.750 ;
        RECT 85.980 74.300 86.280 74.750 ;
        RECT 85.980 73.550 86.280 74.000 ;
        RECT 85.980 72.800 86.280 73.250 ;
        RECT 85.980 72.050 86.280 72.500 ;
        RECT 85.980 71.300 86.280 71.750 ;
        RECT 85.980 70.550 86.280 71.000 ;
        RECT 85.980 69.800 86.280 70.250 ;
        RECT 85.980 69.050 86.280 69.500 ;
        RECT 85.980 68.300 86.280 68.750 ;
        RECT 85.980 67.550 86.280 68.000 ;
        RECT 85.980 66.800 86.280 67.250 ;
        RECT 85.980 66.050 86.280 66.500 ;
        RECT 85.980 65.300 86.280 65.750 ;
        RECT 103.180 74.300 103.480 74.750 ;
        RECT 103.180 73.550 103.480 74.000 ;
        RECT 103.180 72.800 103.480 73.250 ;
        RECT 103.180 72.050 103.480 72.500 ;
        RECT 103.180 71.300 103.480 71.750 ;
        RECT 103.180 70.550 103.480 71.000 ;
        RECT 103.180 69.800 103.480 70.250 ;
        RECT 103.180 69.050 103.480 69.500 ;
        RECT 103.180 68.300 103.480 68.750 ;
        RECT 103.180 67.550 103.480 68.000 ;
        RECT 103.180 66.800 103.480 67.250 ;
        RECT 103.180 66.050 103.480 66.500 ;
        RECT 103.180 65.300 103.480 65.750 ;
        RECT 5.980 54.300 6.280 54.750 ;
        RECT 5.980 53.550 6.280 54.000 ;
        RECT 5.980 52.800 6.280 53.250 ;
        RECT 5.980 52.050 6.280 52.500 ;
        RECT 5.980 51.300 6.280 51.750 ;
        RECT 5.980 50.550 6.280 51.000 ;
        RECT 5.980 49.800 6.280 50.250 ;
        RECT 5.980 49.050 6.280 49.500 ;
        RECT 5.980 48.300 6.280 48.750 ;
        RECT 5.980 47.550 6.280 48.000 ;
        RECT 5.980 46.800 6.280 47.250 ;
        RECT 5.980 46.050 6.280 46.500 ;
        RECT 5.980 45.300 6.280 45.750 ;
        RECT 23.180 54.300 23.480 54.750 ;
        RECT 23.180 53.550 23.480 54.000 ;
        RECT 23.180 52.800 23.480 53.250 ;
        RECT 23.180 52.050 23.480 52.500 ;
        RECT 23.180 51.300 23.480 51.750 ;
        RECT 23.180 50.550 23.480 51.000 ;
        RECT 23.180 49.800 23.480 50.250 ;
        RECT 23.180 49.050 23.480 49.500 ;
        RECT 23.180 48.300 23.480 48.750 ;
        RECT 23.180 47.550 23.480 48.000 ;
        RECT 23.180 46.800 23.480 47.250 ;
        RECT 23.180 46.050 23.480 46.500 ;
        RECT 23.180 45.300 23.480 45.750 ;
        RECT 25.980 54.300 26.280 54.750 ;
        RECT 25.980 53.550 26.280 54.000 ;
        RECT 25.980 52.800 26.280 53.250 ;
        RECT 25.980 52.050 26.280 52.500 ;
        RECT 25.980 51.300 26.280 51.750 ;
        RECT 25.980 50.550 26.280 51.000 ;
        RECT 25.980 49.800 26.280 50.250 ;
        RECT 25.980 49.050 26.280 49.500 ;
        RECT 25.980 48.300 26.280 48.750 ;
        RECT 25.980 47.550 26.280 48.000 ;
        RECT 25.980 46.800 26.280 47.250 ;
        RECT 25.980 46.050 26.280 46.500 ;
        RECT 25.980 45.300 26.280 45.750 ;
        RECT 43.180 54.300 43.480 54.750 ;
        RECT 43.180 53.550 43.480 54.000 ;
        RECT 43.180 52.800 43.480 53.250 ;
        RECT 43.180 52.050 43.480 52.500 ;
        RECT 43.180 51.300 43.480 51.750 ;
        RECT 43.180 50.550 43.480 51.000 ;
        RECT 43.180 49.800 43.480 50.250 ;
        RECT 43.180 49.050 43.480 49.500 ;
        RECT 43.180 48.300 43.480 48.750 ;
        RECT 43.180 47.550 43.480 48.000 ;
        RECT 43.180 46.800 43.480 47.250 ;
        RECT 43.180 46.050 43.480 46.500 ;
        RECT 43.180 45.300 43.480 45.750 ;
        RECT 45.980 54.300 46.280 54.750 ;
        RECT 45.980 53.550 46.280 54.000 ;
        RECT 45.980 52.800 46.280 53.250 ;
        RECT 45.980 52.050 46.280 52.500 ;
        RECT 45.980 51.300 46.280 51.750 ;
        RECT 45.980 50.550 46.280 51.000 ;
        RECT 45.980 49.800 46.280 50.250 ;
        RECT 45.980 49.050 46.280 49.500 ;
        RECT 45.980 48.300 46.280 48.750 ;
        RECT 45.980 47.550 46.280 48.000 ;
        RECT 45.980 46.800 46.280 47.250 ;
        RECT 45.980 46.050 46.280 46.500 ;
        RECT 45.980 45.300 46.280 45.750 ;
        RECT 63.180 54.300 63.480 54.750 ;
        RECT 63.180 53.550 63.480 54.000 ;
        RECT 63.180 52.800 63.480 53.250 ;
        RECT 63.180 52.050 63.480 52.500 ;
        RECT 63.180 51.300 63.480 51.750 ;
        RECT 63.180 50.550 63.480 51.000 ;
        RECT 63.180 49.800 63.480 50.250 ;
        RECT 63.180 49.050 63.480 49.500 ;
        RECT 63.180 48.300 63.480 48.750 ;
        RECT 63.180 47.550 63.480 48.000 ;
        RECT 63.180 46.800 63.480 47.250 ;
        RECT 63.180 46.050 63.480 46.500 ;
        RECT 63.180 45.300 63.480 45.750 ;
        RECT 65.980 54.300 66.280 54.750 ;
        RECT 65.980 53.550 66.280 54.000 ;
        RECT 65.980 52.800 66.280 53.250 ;
        RECT 65.980 52.050 66.280 52.500 ;
        RECT 65.980 51.300 66.280 51.750 ;
        RECT 65.980 50.550 66.280 51.000 ;
        RECT 65.980 49.800 66.280 50.250 ;
        RECT 65.980 49.050 66.280 49.500 ;
        RECT 65.980 48.300 66.280 48.750 ;
        RECT 65.980 47.550 66.280 48.000 ;
        RECT 65.980 46.800 66.280 47.250 ;
        RECT 65.980 46.050 66.280 46.500 ;
        RECT 65.980 45.300 66.280 45.750 ;
        RECT 83.180 54.300 83.480 54.750 ;
        RECT 83.180 53.550 83.480 54.000 ;
        RECT 83.180 52.800 83.480 53.250 ;
        RECT 83.180 52.050 83.480 52.500 ;
        RECT 83.180 51.300 83.480 51.750 ;
        RECT 83.180 50.550 83.480 51.000 ;
        RECT 83.180 49.800 83.480 50.250 ;
        RECT 83.180 49.050 83.480 49.500 ;
        RECT 83.180 48.300 83.480 48.750 ;
        RECT 83.180 47.550 83.480 48.000 ;
        RECT 83.180 46.800 83.480 47.250 ;
        RECT 83.180 46.050 83.480 46.500 ;
        RECT 83.180 45.300 83.480 45.750 ;
        RECT 85.980 54.300 86.280 54.750 ;
        RECT 85.980 53.550 86.280 54.000 ;
        RECT 85.980 52.800 86.280 53.250 ;
        RECT 85.980 52.050 86.280 52.500 ;
        RECT 85.980 51.300 86.280 51.750 ;
        RECT 85.980 50.550 86.280 51.000 ;
        RECT 85.980 49.800 86.280 50.250 ;
        RECT 85.980 49.050 86.280 49.500 ;
        RECT 85.980 48.300 86.280 48.750 ;
        RECT 85.980 47.550 86.280 48.000 ;
        RECT 85.980 46.800 86.280 47.250 ;
        RECT 85.980 46.050 86.280 46.500 ;
        RECT 85.980 45.300 86.280 45.750 ;
        RECT 103.180 54.300 103.480 54.750 ;
        RECT 103.180 53.550 103.480 54.000 ;
        RECT 103.180 52.800 103.480 53.250 ;
        RECT 103.180 52.050 103.480 52.500 ;
        RECT 103.180 51.300 103.480 51.750 ;
        RECT 103.180 50.550 103.480 51.000 ;
        RECT 103.180 49.800 103.480 50.250 ;
        RECT 103.180 49.050 103.480 49.500 ;
        RECT 103.180 48.300 103.480 48.750 ;
        RECT 103.180 47.550 103.480 48.000 ;
        RECT 103.180 46.800 103.480 47.250 ;
        RECT 103.180 46.050 103.480 46.500 ;
        RECT 103.180 45.300 103.480 45.750 ;
        RECT 5.980 34.300 6.280 34.750 ;
        RECT 5.980 33.550 6.280 34.000 ;
        RECT 5.980 32.800 6.280 33.250 ;
        RECT 5.980 32.050 6.280 32.500 ;
        RECT 5.980 31.300 6.280 31.750 ;
        RECT 5.980 30.550 6.280 31.000 ;
        RECT 5.980 29.800 6.280 30.250 ;
        RECT 5.980 29.050 6.280 29.500 ;
        RECT 5.980 28.300 6.280 28.750 ;
        RECT 5.980 27.550 6.280 28.000 ;
        RECT 5.980 26.800 6.280 27.250 ;
        RECT 5.980 26.050 6.280 26.500 ;
        RECT 5.980 25.300 6.280 25.750 ;
        RECT 23.180 34.300 23.480 34.750 ;
        RECT 23.180 33.550 23.480 34.000 ;
        RECT 23.180 32.800 23.480 33.250 ;
        RECT 23.180 32.050 23.480 32.500 ;
        RECT 23.180 31.300 23.480 31.750 ;
        RECT 23.180 30.550 23.480 31.000 ;
        RECT 23.180 29.800 23.480 30.250 ;
        RECT 23.180 29.050 23.480 29.500 ;
        RECT 23.180 28.300 23.480 28.750 ;
        RECT 23.180 27.550 23.480 28.000 ;
        RECT 23.180 26.800 23.480 27.250 ;
        RECT 23.180 26.050 23.480 26.500 ;
        RECT 23.180 25.300 23.480 25.750 ;
        RECT 25.980 34.300 26.280 34.750 ;
        RECT 25.980 33.550 26.280 34.000 ;
        RECT 25.980 32.800 26.280 33.250 ;
        RECT 25.980 32.050 26.280 32.500 ;
        RECT 25.980 31.300 26.280 31.750 ;
        RECT 25.980 30.550 26.280 31.000 ;
        RECT 25.980 29.800 26.280 30.250 ;
        RECT 25.980 29.050 26.280 29.500 ;
        RECT 25.980 28.300 26.280 28.750 ;
        RECT 25.980 27.550 26.280 28.000 ;
        RECT 25.980 26.800 26.280 27.250 ;
        RECT 25.980 26.050 26.280 26.500 ;
        RECT 25.980 25.300 26.280 25.750 ;
        RECT 43.180 34.300 43.480 34.750 ;
        RECT 43.180 33.550 43.480 34.000 ;
        RECT 43.180 32.800 43.480 33.250 ;
        RECT 43.180 32.050 43.480 32.500 ;
        RECT 43.180 31.300 43.480 31.750 ;
        RECT 43.180 30.550 43.480 31.000 ;
        RECT 43.180 29.800 43.480 30.250 ;
        RECT 43.180 29.050 43.480 29.500 ;
        RECT 43.180 28.300 43.480 28.750 ;
        RECT 43.180 27.550 43.480 28.000 ;
        RECT 43.180 26.800 43.480 27.250 ;
        RECT 43.180 26.050 43.480 26.500 ;
        RECT 43.180 25.300 43.480 25.750 ;
        RECT 45.980 34.300 46.280 34.750 ;
        RECT 45.980 33.550 46.280 34.000 ;
        RECT 45.980 32.800 46.280 33.250 ;
        RECT 45.980 32.050 46.280 32.500 ;
        RECT 45.980 31.300 46.280 31.750 ;
        RECT 45.980 30.550 46.280 31.000 ;
        RECT 45.980 29.800 46.280 30.250 ;
        RECT 45.980 29.050 46.280 29.500 ;
        RECT 45.980 28.300 46.280 28.750 ;
        RECT 45.980 27.550 46.280 28.000 ;
        RECT 45.980 26.800 46.280 27.250 ;
        RECT 45.980 26.050 46.280 26.500 ;
        RECT 45.980 25.300 46.280 25.750 ;
        RECT 63.180 34.300 63.480 34.750 ;
        RECT 63.180 33.550 63.480 34.000 ;
        RECT 63.180 32.800 63.480 33.250 ;
        RECT 63.180 32.050 63.480 32.500 ;
        RECT 63.180 31.300 63.480 31.750 ;
        RECT 63.180 30.550 63.480 31.000 ;
        RECT 63.180 29.800 63.480 30.250 ;
        RECT 63.180 29.050 63.480 29.500 ;
        RECT 63.180 28.300 63.480 28.750 ;
        RECT 63.180 27.550 63.480 28.000 ;
        RECT 63.180 26.800 63.480 27.250 ;
        RECT 63.180 26.050 63.480 26.500 ;
        RECT 63.180 25.300 63.480 25.750 ;
        RECT 65.980 34.300 66.280 34.750 ;
        RECT 65.980 33.550 66.280 34.000 ;
        RECT 65.980 32.800 66.280 33.250 ;
        RECT 65.980 32.050 66.280 32.500 ;
        RECT 65.980 31.300 66.280 31.750 ;
        RECT 65.980 30.550 66.280 31.000 ;
        RECT 65.980 29.800 66.280 30.250 ;
        RECT 65.980 29.050 66.280 29.500 ;
        RECT 65.980 28.300 66.280 28.750 ;
        RECT 65.980 27.550 66.280 28.000 ;
        RECT 65.980 26.800 66.280 27.250 ;
        RECT 65.980 26.050 66.280 26.500 ;
        RECT 65.980 25.300 66.280 25.750 ;
        RECT 83.180 34.300 83.480 34.750 ;
        RECT 83.180 33.550 83.480 34.000 ;
        RECT 83.180 32.800 83.480 33.250 ;
        RECT 83.180 32.050 83.480 32.500 ;
        RECT 83.180 31.300 83.480 31.750 ;
        RECT 83.180 30.550 83.480 31.000 ;
        RECT 83.180 29.800 83.480 30.250 ;
        RECT 83.180 29.050 83.480 29.500 ;
        RECT 83.180 28.300 83.480 28.750 ;
        RECT 83.180 27.550 83.480 28.000 ;
        RECT 83.180 26.800 83.480 27.250 ;
        RECT 83.180 26.050 83.480 26.500 ;
        RECT 83.180 25.300 83.480 25.750 ;
        RECT 85.980 34.300 86.280 34.750 ;
        RECT 85.980 33.550 86.280 34.000 ;
        RECT 85.980 32.800 86.280 33.250 ;
        RECT 85.980 32.050 86.280 32.500 ;
        RECT 85.980 31.300 86.280 31.750 ;
        RECT 85.980 30.550 86.280 31.000 ;
        RECT 85.980 29.800 86.280 30.250 ;
        RECT 85.980 29.050 86.280 29.500 ;
        RECT 85.980 28.300 86.280 28.750 ;
        RECT 85.980 27.550 86.280 28.000 ;
        RECT 85.980 26.800 86.280 27.250 ;
        RECT 85.980 26.050 86.280 26.500 ;
        RECT 85.980 25.300 86.280 25.750 ;
        RECT 103.180 34.300 103.480 34.750 ;
        RECT 103.180 33.550 103.480 34.000 ;
        RECT 103.180 32.800 103.480 33.250 ;
        RECT 103.180 32.050 103.480 32.500 ;
        RECT 103.180 31.300 103.480 31.750 ;
        RECT 103.180 30.550 103.480 31.000 ;
        RECT 103.180 29.800 103.480 30.250 ;
        RECT 103.180 29.050 103.480 29.500 ;
        RECT 103.180 28.300 103.480 28.750 ;
        RECT 103.180 27.550 103.480 28.000 ;
        RECT 103.180 26.800 103.480 27.250 ;
        RECT 103.180 26.050 103.480 26.500 ;
        RECT 103.180 25.300 103.480 25.750 ;
        RECT 5.980 14.300 6.280 14.750 ;
        RECT 5.980 13.550 6.280 14.000 ;
        RECT 5.980 12.800 6.280 13.250 ;
        RECT 5.980 12.050 6.280 12.500 ;
        RECT 5.980 11.300 6.280 11.750 ;
        RECT 5.980 10.550 6.280 11.000 ;
        RECT 5.980 9.800 6.280 10.250 ;
        RECT 5.980 9.050 6.280 9.500 ;
        RECT 5.980 8.300 6.280 8.750 ;
        RECT 5.980 7.550 6.280 8.000 ;
        RECT 5.980 6.800 6.280 7.250 ;
        RECT 5.980 6.050 6.280 6.500 ;
        RECT 5.980 5.300 6.280 5.750 ;
        RECT 23.180 14.300 23.480 14.750 ;
        RECT 23.180 13.550 23.480 14.000 ;
        RECT 23.180 12.800 23.480 13.250 ;
        RECT 23.180 12.050 23.480 12.500 ;
        RECT 23.180 11.300 23.480 11.750 ;
        RECT 23.180 10.550 23.480 11.000 ;
        RECT 23.180 9.800 23.480 10.250 ;
        RECT 23.180 9.050 23.480 9.500 ;
        RECT 23.180 8.300 23.480 8.750 ;
        RECT 23.180 7.550 23.480 8.000 ;
        RECT 23.180 6.800 23.480 7.250 ;
        RECT 23.180 6.050 23.480 6.500 ;
        RECT 23.180 5.300 23.480 5.750 ;
        RECT 25.980 14.300 26.280 14.750 ;
        RECT 25.980 13.550 26.280 14.000 ;
        RECT 25.980 12.800 26.280 13.250 ;
        RECT 25.980 12.050 26.280 12.500 ;
        RECT 25.980 11.300 26.280 11.750 ;
        RECT 25.980 10.550 26.280 11.000 ;
        RECT 25.980 9.800 26.280 10.250 ;
        RECT 25.980 9.050 26.280 9.500 ;
        RECT 25.980 8.300 26.280 8.750 ;
        RECT 25.980 7.550 26.280 8.000 ;
        RECT 25.980 6.800 26.280 7.250 ;
        RECT 25.980 6.050 26.280 6.500 ;
        RECT 25.980 5.300 26.280 5.750 ;
        RECT 43.180 14.300 43.480 14.750 ;
        RECT 43.180 13.550 43.480 14.000 ;
        RECT 43.180 12.800 43.480 13.250 ;
        RECT 43.180 12.050 43.480 12.500 ;
        RECT 43.180 11.300 43.480 11.750 ;
        RECT 43.180 10.550 43.480 11.000 ;
        RECT 43.180 9.800 43.480 10.250 ;
        RECT 43.180 9.050 43.480 9.500 ;
        RECT 43.180 8.300 43.480 8.750 ;
        RECT 43.180 7.550 43.480 8.000 ;
        RECT 43.180 6.800 43.480 7.250 ;
        RECT 43.180 6.050 43.480 6.500 ;
        RECT 43.180 5.300 43.480 5.750 ;
        RECT 45.980 14.300 46.280 14.750 ;
        RECT 45.980 13.550 46.280 14.000 ;
        RECT 45.980 12.800 46.280 13.250 ;
        RECT 45.980 12.050 46.280 12.500 ;
        RECT 45.980 11.300 46.280 11.750 ;
        RECT 45.980 10.550 46.280 11.000 ;
        RECT 45.980 9.800 46.280 10.250 ;
        RECT 45.980 9.050 46.280 9.500 ;
        RECT 45.980 8.300 46.280 8.750 ;
        RECT 45.980 7.550 46.280 8.000 ;
        RECT 45.980 6.800 46.280 7.250 ;
        RECT 45.980 6.050 46.280 6.500 ;
        RECT 45.980 5.300 46.280 5.750 ;
        RECT 63.180 14.300 63.480 14.750 ;
        RECT 63.180 13.550 63.480 14.000 ;
        RECT 63.180 12.800 63.480 13.250 ;
        RECT 63.180 12.050 63.480 12.500 ;
        RECT 63.180 11.300 63.480 11.750 ;
        RECT 63.180 10.550 63.480 11.000 ;
        RECT 63.180 9.800 63.480 10.250 ;
        RECT 63.180 9.050 63.480 9.500 ;
        RECT 63.180 8.300 63.480 8.750 ;
        RECT 63.180 7.550 63.480 8.000 ;
        RECT 63.180 6.800 63.480 7.250 ;
        RECT 63.180 6.050 63.480 6.500 ;
        RECT 63.180 5.300 63.480 5.750 ;
        RECT 65.980 14.300 66.280 14.750 ;
        RECT 65.980 13.550 66.280 14.000 ;
        RECT 65.980 12.800 66.280 13.250 ;
        RECT 65.980 12.050 66.280 12.500 ;
        RECT 65.980 11.300 66.280 11.750 ;
        RECT 65.980 10.550 66.280 11.000 ;
        RECT 65.980 9.800 66.280 10.250 ;
        RECT 65.980 9.050 66.280 9.500 ;
        RECT 65.980 8.300 66.280 8.750 ;
        RECT 65.980 7.550 66.280 8.000 ;
        RECT 65.980 6.800 66.280 7.250 ;
        RECT 65.980 6.050 66.280 6.500 ;
        RECT 65.980 5.300 66.280 5.750 ;
        RECT 83.180 14.300 83.480 14.750 ;
        RECT 83.180 13.550 83.480 14.000 ;
        RECT 83.180 12.800 83.480 13.250 ;
        RECT 83.180 12.050 83.480 12.500 ;
        RECT 83.180 11.300 83.480 11.750 ;
        RECT 83.180 10.550 83.480 11.000 ;
        RECT 83.180 9.800 83.480 10.250 ;
        RECT 83.180 9.050 83.480 9.500 ;
        RECT 83.180 8.300 83.480 8.750 ;
        RECT 83.180 7.550 83.480 8.000 ;
        RECT 83.180 6.800 83.480 7.250 ;
        RECT 83.180 6.050 83.480 6.500 ;
        RECT 83.180 5.300 83.480 5.750 ;
        RECT 85.980 14.300 86.280 14.750 ;
        RECT 85.980 13.550 86.280 14.000 ;
        RECT 85.980 12.800 86.280 13.250 ;
        RECT 85.980 12.050 86.280 12.500 ;
        RECT 85.980 11.300 86.280 11.750 ;
        RECT 85.980 10.550 86.280 11.000 ;
        RECT 85.980 9.800 86.280 10.250 ;
        RECT 85.980 9.050 86.280 9.500 ;
        RECT 85.980 8.300 86.280 8.750 ;
        RECT 85.980 7.550 86.280 8.000 ;
        RECT 85.980 6.800 86.280 7.250 ;
        RECT 85.980 6.050 86.280 6.500 ;
        RECT 85.980 5.300 86.280 5.750 ;
        RECT 103.180 14.300 103.480 14.750 ;
        RECT 103.180 13.550 103.480 14.000 ;
        RECT 103.180 12.800 103.480 13.250 ;
        RECT 103.180 12.050 103.480 12.500 ;
        RECT 103.180 11.300 103.480 11.750 ;
        RECT 103.180 10.550 103.480 11.000 ;
        RECT 103.180 9.800 103.480 10.250 ;
        RECT 103.180 9.050 103.480 9.500 ;
        RECT 103.180 8.300 103.480 8.750 ;
        RECT 103.180 7.550 103.480 8.000 ;
        RECT 103.180 6.800 103.480 7.250 ;
        RECT 103.180 6.050 103.480 6.500 ;
        RECT 103.180 5.300 103.480 5.750 ;
      LAYER met1 ;
        RECT 11.530 378.800 17.930 380.000 ;
        RECT 31.530 378.800 37.930 380.000 ;
        RECT 51.530 378.800 57.930 380.000 ;
        RECT 71.530 378.800 77.930 380.000 ;
        RECT 91.530 378.800 97.930 380.000 ;
        RECT 14.230 378.150 15.230 378.800 ;
        RECT 34.230 378.150 35.230 378.800 ;
        RECT 54.230 378.150 55.230 378.800 ;
        RECT 74.230 378.150 75.230 378.800 ;
        RECT 94.230 378.150 95.230 378.800 ;
        RECT 10.880 378.000 18.580 378.150 ;
        RECT 30.880 378.000 38.580 378.150 ;
        RECT 50.880 378.000 58.580 378.150 ;
        RECT 70.880 378.000 78.580 378.150 ;
        RECT 90.880 378.000 98.580 378.150 ;
        RECT 5.930 373.200 6.680 375.000 ;
        RECT 4.730 370.450 6.680 373.200 ;
        RECT 4.730 369.550 4.880 370.450 ;
        RECT 5.530 370.300 6.680 370.450 ;
        RECT 6.830 370.300 6.980 377.850 ;
        RECT 7.430 370.300 7.580 377.850 ;
        RECT 8.030 370.300 8.180 377.850 ;
        RECT 8.630 370.300 8.780 377.850 ;
        RECT 9.230 370.300 9.380 377.850 ;
        RECT 9.830 370.300 9.980 377.850 ;
        RECT 14.230 377.550 15.230 378.000 ;
        RECT 10.880 377.400 18.580 377.550 ;
        RECT 14.230 376.950 15.230 377.400 ;
        RECT 10.880 376.800 18.580 376.950 ;
        RECT 14.230 376.350 15.230 376.800 ;
        RECT 10.880 376.200 18.580 376.350 ;
        RECT 14.230 375.750 15.230 376.200 ;
        RECT 10.880 375.600 18.580 375.750 ;
        RECT 14.230 375.150 15.230 375.600 ;
        RECT 10.880 375.000 18.580 375.150 ;
        RECT 14.230 374.550 15.230 375.000 ;
        RECT 10.880 374.400 18.580 374.550 ;
        RECT 14.230 373.950 15.230 374.400 ;
        RECT 10.880 373.800 18.580 373.950 ;
        RECT 14.230 373.350 15.230 373.800 ;
        RECT 10.880 373.200 18.580 373.350 ;
        RECT 14.230 372.750 15.230 373.200 ;
        RECT 10.880 372.600 18.580 372.750 ;
        RECT 14.230 372.150 15.230 372.600 ;
        RECT 10.880 372.000 18.580 372.150 ;
        RECT 14.230 371.550 15.230 372.000 ;
        RECT 10.880 371.400 18.580 371.550 ;
        RECT 14.230 370.950 15.230 371.400 ;
        RECT 10.880 370.800 18.580 370.950 ;
        RECT 14.230 370.300 15.230 370.800 ;
        RECT 19.480 370.300 19.630 377.850 ;
        RECT 20.080 370.300 20.230 377.850 ;
        RECT 20.680 370.300 20.830 377.850 ;
        RECT 21.280 370.300 21.430 377.850 ;
        RECT 21.880 370.300 22.030 377.850 ;
        RECT 22.480 370.300 22.630 377.850 ;
        RECT 22.780 373.200 23.530 375.000 ;
        RECT 25.930 373.200 26.680 375.000 ;
        RECT 22.780 370.450 26.680 373.200 ;
        RECT 22.780 370.300 23.930 370.450 ;
        RECT 5.530 369.700 23.930 370.300 ;
        RECT 5.530 369.550 6.680 369.700 ;
        RECT 4.730 366.800 6.680 369.550 ;
        RECT 5.930 365.050 6.680 366.800 ;
        RECT 6.830 362.150 6.980 369.700 ;
        RECT 7.430 362.150 7.580 369.700 ;
        RECT 8.030 362.150 8.180 369.700 ;
        RECT 8.630 362.150 8.780 369.700 ;
        RECT 9.230 362.150 9.380 369.700 ;
        RECT 9.830 362.150 9.980 369.700 ;
        RECT 14.230 369.200 15.230 369.700 ;
        RECT 10.880 369.050 18.580 369.200 ;
        RECT 14.230 368.600 15.230 369.050 ;
        RECT 10.880 368.450 18.580 368.600 ;
        RECT 14.230 368.000 15.230 368.450 ;
        RECT 10.880 367.850 18.580 368.000 ;
        RECT 14.230 367.400 15.230 367.850 ;
        RECT 10.880 367.250 18.580 367.400 ;
        RECT 14.230 366.800 15.230 367.250 ;
        RECT 10.880 366.650 18.580 366.800 ;
        RECT 14.230 366.200 15.230 366.650 ;
        RECT 10.880 366.050 18.580 366.200 ;
        RECT 14.230 365.600 15.230 366.050 ;
        RECT 10.880 365.450 18.580 365.600 ;
        RECT 14.230 365.000 15.230 365.450 ;
        RECT 10.880 364.850 18.580 365.000 ;
        RECT 14.230 364.400 15.230 364.850 ;
        RECT 10.880 364.250 18.580 364.400 ;
        RECT 14.230 363.800 15.230 364.250 ;
        RECT 10.880 363.650 18.580 363.800 ;
        RECT 14.230 363.200 15.230 363.650 ;
        RECT 10.880 363.050 18.580 363.200 ;
        RECT 14.230 362.600 15.230 363.050 ;
        RECT 10.880 362.450 18.580 362.600 ;
        RECT 14.230 362.000 15.230 362.450 ;
        RECT 19.480 362.150 19.630 369.700 ;
        RECT 20.080 362.150 20.230 369.700 ;
        RECT 20.680 362.150 20.830 369.700 ;
        RECT 21.280 362.150 21.430 369.700 ;
        RECT 21.880 362.150 22.030 369.700 ;
        RECT 22.480 362.150 22.630 369.700 ;
        RECT 22.780 369.550 23.930 369.700 ;
        RECT 24.580 369.550 24.880 370.450 ;
        RECT 25.530 370.300 26.680 370.450 ;
        RECT 26.830 370.300 26.980 377.850 ;
        RECT 27.430 370.300 27.580 377.850 ;
        RECT 28.030 370.300 28.180 377.850 ;
        RECT 28.630 370.300 28.780 377.850 ;
        RECT 29.230 370.300 29.380 377.850 ;
        RECT 29.830 370.300 29.980 377.850 ;
        RECT 34.230 377.550 35.230 378.000 ;
        RECT 30.880 377.400 38.580 377.550 ;
        RECT 34.230 376.950 35.230 377.400 ;
        RECT 30.880 376.800 38.580 376.950 ;
        RECT 34.230 376.350 35.230 376.800 ;
        RECT 30.880 376.200 38.580 376.350 ;
        RECT 34.230 375.750 35.230 376.200 ;
        RECT 30.880 375.600 38.580 375.750 ;
        RECT 34.230 375.150 35.230 375.600 ;
        RECT 30.880 375.000 38.580 375.150 ;
        RECT 34.230 374.550 35.230 375.000 ;
        RECT 30.880 374.400 38.580 374.550 ;
        RECT 34.230 373.950 35.230 374.400 ;
        RECT 30.880 373.800 38.580 373.950 ;
        RECT 34.230 373.350 35.230 373.800 ;
        RECT 30.880 373.200 38.580 373.350 ;
        RECT 34.230 372.750 35.230 373.200 ;
        RECT 30.880 372.600 38.580 372.750 ;
        RECT 34.230 372.150 35.230 372.600 ;
        RECT 30.880 372.000 38.580 372.150 ;
        RECT 34.230 371.550 35.230 372.000 ;
        RECT 30.880 371.400 38.580 371.550 ;
        RECT 34.230 370.950 35.230 371.400 ;
        RECT 30.880 370.800 38.580 370.950 ;
        RECT 34.230 370.300 35.230 370.800 ;
        RECT 39.480 370.300 39.630 377.850 ;
        RECT 40.080 370.300 40.230 377.850 ;
        RECT 40.680 370.300 40.830 377.850 ;
        RECT 41.280 370.300 41.430 377.850 ;
        RECT 41.880 370.300 42.030 377.850 ;
        RECT 42.480 370.300 42.630 377.850 ;
        RECT 42.780 373.200 43.530 375.000 ;
        RECT 45.930 373.200 46.680 375.000 ;
        RECT 42.780 370.450 46.680 373.200 ;
        RECT 42.780 370.300 43.930 370.450 ;
        RECT 25.530 369.700 43.930 370.300 ;
        RECT 25.530 369.550 26.680 369.700 ;
        RECT 22.780 366.800 26.680 369.550 ;
        RECT 22.780 365.050 23.530 366.800 ;
        RECT 25.930 365.050 26.680 366.800 ;
        RECT 26.830 362.150 26.980 369.700 ;
        RECT 27.430 362.150 27.580 369.700 ;
        RECT 28.030 362.150 28.180 369.700 ;
        RECT 28.630 362.150 28.780 369.700 ;
        RECT 29.230 362.150 29.380 369.700 ;
        RECT 29.830 362.150 29.980 369.700 ;
        RECT 34.230 369.200 35.230 369.700 ;
        RECT 30.880 369.050 38.580 369.200 ;
        RECT 34.230 368.600 35.230 369.050 ;
        RECT 30.880 368.450 38.580 368.600 ;
        RECT 34.230 368.000 35.230 368.450 ;
        RECT 30.880 367.850 38.580 368.000 ;
        RECT 34.230 367.400 35.230 367.850 ;
        RECT 30.880 367.250 38.580 367.400 ;
        RECT 34.230 366.800 35.230 367.250 ;
        RECT 30.880 366.650 38.580 366.800 ;
        RECT 34.230 366.200 35.230 366.650 ;
        RECT 30.880 366.050 38.580 366.200 ;
        RECT 34.230 365.600 35.230 366.050 ;
        RECT 30.880 365.450 38.580 365.600 ;
        RECT 34.230 365.000 35.230 365.450 ;
        RECT 30.880 364.850 38.580 365.000 ;
        RECT 34.230 364.400 35.230 364.850 ;
        RECT 30.880 364.250 38.580 364.400 ;
        RECT 34.230 363.800 35.230 364.250 ;
        RECT 30.880 363.650 38.580 363.800 ;
        RECT 34.230 363.200 35.230 363.650 ;
        RECT 30.880 363.050 38.580 363.200 ;
        RECT 34.230 362.600 35.230 363.050 ;
        RECT 30.880 362.450 38.580 362.600 ;
        RECT 34.230 362.000 35.230 362.450 ;
        RECT 39.480 362.150 39.630 369.700 ;
        RECT 40.080 362.150 40.230 369.700 ;
        RECT 40.680 362.150 40.830 369.700 ;
        RECT 41.280 362.150 41.430 369.700 ;
        RECT 41.880 362.150 42.030 369.700 ;
        RECT 42.480 362.150 42.630 369.700 ;
        RECT 42.780 369.550 43.930 369.700 ;
        RECT 44.580 369.550 44.880 370.450 ;
        RECT 45.530 370.300 46.680 370.450 ;
        RECT 46.830 370.300 46.980 377.850 ;
        RECT 47.430 370.300 47.580 377.850 ;
        RECT 48.030 370.300 48.180 377.850 ;
        RECT 48.630 370.300 48.780 377.850 ;
        RECT 49.230 370.300 49.380 377.850 ;
        RECT 49.830 370.300 49.980 377.850 ;
        RECT 54.230 377.550 55.230 378.000 ;
        RECT 50.880 377.400 58.580 377.550 ;
        RECT 54.230 376.950 55.230 377.400 ;
        RECT 50.880 376.800 58.580 376.950 ;
        RECT 54.230 376.350 55.230 376.800 ;
        RECT 50.880 376.200 58.580 376.350 ;
        RECT 54.230 375.750 55.230 376.200 ;
        RECT 50.880 375.600 58.580 375.750 ;
        RECT 54.230 375.150 55.230 375.600 ;
        RECT 50.880 375.000 58.580 375.150 ;
        RECT 54.230 374.550 55.230 375.000 ;
        RECT 50.880 374.400 58.580 374.550 ;
        RECT 54.230 373.950 55.230 374.400 ;
        RECT 50.880 373.800 58.580 373.950 ;
        RECT 54.230 373.350 55.230 373.800 ;
        RECT 50.880 373.200 58.580 373.350 ;
        RECT 54.230 372.750 55.230 373.200 ;
        RECT 50.880 372.600 58.580 372.750 ;
        RECT 54.230 372.150 55.230 372.600 ;
        RECT 50.880 372.000 58.580 372.150 ;
        RECT 54.230 371.550 55.230 372.000 ;
        RECT 50.880 371.400 58.580 371.550 ;
        RECT 54.230 370.950 55.230 371.400 ;
        RECT 50.880 370.800 58.580 370.950 ;
        RECT 54.230 370.300 55.230 370.800 ;
        RECT 59.480 370.300 59.630 377.850 ;
        RECT 60.080 370.300 60.230 377.850 ;
        RECT 60.680 370.300 60.830 377.850 ;
        RECT 61.280 370.300 61.430 377.850 ;
        RECT 61.880 370.300 62.030 377.850 ;
        RECT 62.480 370.300 62.630 377.850 ;
        RECT 62.780 373.200 63.530 375.000 ;
        RECT 65.930 373.200 66.680 375.000 ;
        RECT 62.780 370.450 66.680 373.200 ;
        RECT 62.780 370.300 63.930 370.450 ;
        RECT 45.530 369.700 63.930 370.300 ;
        RECT 45.530 369.550 46.680 369.700 ;
        RECT 42.780 366.800 46.680 369.550 ;
        RECT 42.780 365.050 43.530 366.800 ;
        RECT 45.930 365.050 46.680 366.800 ;
        RECT 46.830 362.150 46.980 369.700 ;
        RECT 47.430 362.150 47.580 369.700 ;
        RECT 48.030 362.150 48.180 369.700 ;
        RECT 48.630 362.150 48.780 369.700 ;
        RECT 49.230 362.150 49.380 369.700 ;
        RECT 49.830 362.150 49.980 369.700 ;
        RECT 54.230 369.200 55.230 369.700 ;
        RECT 50.880 369.050 58.580 369.200 ;
        RECT 54.230 368.600 55.230 369.050 ;
        RECT 50.880 368.450 58.580 368.600 ;
        RECT 54.230 368.000 55.230 368.450 ;
        RECT 50.880 367.850 58.580 368.000 ;
        RECT 54.230 367.400 55.230 367.850 ;
        RECT 50.880 367.250 58.580 367.400 ;
        RECT 54.230 366.800 55.230 367.250 ;
        RECT 50.880 366.650 58.580 366.800 ;
        RECT 54.230 366.200 55.230 366.650 ;
        RECT 50.880 366.050 58.580 366.200 ;
        RECT 54.230 365.600 55.230 366.050 ;
        RECT 50.880 365.450 58.580 365.600 ;
        RECT 54.230 365.000 55.230 365.450 ;
        RECT 50.880 364.850 58.580 365.000 ;
        RECT 54.230 364.400 55.230 364.850 ;
        RECT 50.880 364.250 58.580 364.400 ;
        RECT 54.230 363.800 55.230 364.250 ;
        RECT 50.880 363.650 58.580 363.800 ;
        RECT 54.230 363.200 55.230 363.650 ;
        RECT 50.880 363.050 58.580 363.200 ;
        RECT 54.230 362.600 55.230 363.050 ;
        RECT 50.880 362.450 58.580 362.600 ;
        RECT 54.230 362.000 55.230 362.450 ;
        RECT 59.480 362.150 59.630 369.700 ;
        RECT 60.080 362.150 60.230 369.700 ;
        RECT 60.680 362.150 60.830 369.700 ;
        RECT 61.280 362.150 61.430 369.700 ;
        RECT 61.880 362.150 62.030 369.700 ;
        RECT 62.480 362.150 62.630 369.700 ;
        RECT 62.780 369.550 63.930 369.700 ;
        RECT 64.580 369.550 64.880 370.450 ;
        RECT 65.530 370.300 66.680 370.450 ;
        RECT 66.830 370.300 66.980 377.850 ;
        RECT 67.430 370.300 67.580 377.850 ;
        RECT 68.030 370.300 68.180 377.850 ;
        RECT 68.630 370.300 68.780 377.850 ;
        RECT 69.230 370.300 69.380 377.850 ;
        RECT 69.830 370.300 69.980 377.850 ;
        RECT 74.230 377.550 75.230 378.000 ;
        RECT 70.880 377.400 78.580 377.550 ;
        RECT 74.230 376.950 75.230 377.400 ;
        RECT 70.880 376.800 78.580 376.950 ;
        RECT 74.230 376.350 75.230 376.800 ;
        RECT 70.880 376.200 78.580 376.350 ;
        RECT 74.230 375.750 75.230 376.200 ;
        RECT 70.880 375.600 78.580 375.750 ;
        RECT 74.230 375.150 75.230 375.600 ;
        RECT 70.880 375.000 78.580 375.150 ;
        RECT 74.230 374.550 75.230 375.000 ;
        RECT 70.880 374.400 78.580 374.550 ;
        RECT 74.230 373.950 75.230 374.400 ;
        RECT 70.880 373.800 78.580 373.950 ;
        RECT 74.230 373.350 75.230 373.800 ;
        RECT 70.880 373.200 78.580 373.350 ;
        RECT 74.230 372.750 75.230 373.200 ;
        RECT 70.880 372.600 78.580 372.750 ;
        RECT 74.230 372.150 75.230 372.600 ;
        RECT 70.880 372.000 78.580 372.150 ;
        RECT 74.230 371.550 75.230 372.000 ;
        RECT 70.880 371.400 78.580 371.550 ;
        RECT 74.230 370.950 75.230 371.400 ;
        RECT 70.880 370.800 78.580 370.950 ;
        RECT 74.230 370.300 75.230 370.800 ;
        RECT 79.480 370.300 79.630 377.850 ;
        RECT 80.080 370.300 80.230 377.850 ;
        RECT 80.680 370.300 80.830 377.850 ;
        RECT 81.280 370.300 81.430 377.850 ;
        RECT 81.880 370.300 82.030 377.850 ;
        RECT 82.480 370.300 82.630 377.850 ;
        RECT 82.780 373.200 83.530 375.000 ;
        RECT 85.930 373.200 86.680 375.000 ;
        RECT 82.780 370.450 86.680 373.200 ;
        RECT 82.780 370.300 83.930 370.450 ;
        RECT 65.530 369.700 83.930 370.300 ;
        RECT 65.530 369.550 66.680 369.700 ;
        RECT 62.780 366.800 66.680 369.550 ;
        RECT 62.780 365.050 63.530 366.800 ;
        RECT 65.930 365.050 66.680 366.800 ;
        RECT 66.830 362.150 66.980 369.700 ;
        RECT 67.430 362.150 67.580 369.700 ;
        RECT 68.030 362.150 68.180 369.700 ;
        RECT 68.630 362.150 68.780 369.700 ;
        RECT 69.230 362.150 69.380 369.700 ;
        RECT 69.830 362.150 69.980 369.700 ;
        RECT 74.230 369.200 75.230 369.700 ;
        RECT 70.880 369.050 78.580 369.200 ;
        RECT 74.230 368.600 75.230 369.050 ;
        RECT 70.880 368.450 78.580 368.600 ;
        RECT 74.230 368.000 75.230 368.450 ;
        RECT 70.880 367.850 78.580 368.000 ;
        RECT 74.230 367.400 75.230 367.850 ;
        RECT 70.880 367.250 78.580 367.400 ;
        RECT 74.230 366.800 75.230 367.250 ;
        RECT 70.880 366.650 78.580 366.800 ;
        RECT 74.230 366.200 75.230 366.650 ;
        RECT 70.880 366.050 78.580 366.200 ;
        RECT 74.230 365.600 75.230 366.050 ;
        RECT 70.880 365.450 78.580 365.600 ;
        RECT 74.230 365.000 75.230 365.450 ;
        RECT 70.880 364.850 78.580 365.000 ;
        RECT 74.230 364.400 75.230 364.850 ;
        RECT 70.880 364.250 78.580 364.400 ;
        RECT 74.230 363.800 75.230 364.250 ;
        RECT 70.880 363.650 78.580 363.800 ;
        RECT 74.230 363.200 75.230 363.650 ;
        RECT 70.880 363.050 78.580 363.200 ;
        RECT 74.230 362.600 75.230 363.050 ;
        RECT 70.880 362.450 78.580 362.600 ;
        RECT 74.230 362.000 75.230 362.450 ;
        RECT 79.480 362.150 79.630 369.700 ;
        RECT 80.080 362.150 80.230 369.700 ;
        RECT 80.680 362.150 80.830 369.700 ;
        RECT 81.280 362.150 81.430 369.700 ;
        RECT 81.880 362.150 82.030 369.700 ;
        RECT 82.480 362.150 82.630 369.700 ;
        RECT 82.780 369.550 83.930 369.700 ;
        RECT 84.580 369.550 84.880 370.450 ;
        RECT 85.530 370.300 86.680 370.450 ;
        RECT 86.830 370.300 86.980 377.850 ;
        RECT 87.430 370.300 87.580 377.850 ;
        RECT 88.030 370.300 88.180 377.850 ;
        RECT 88.630 370.300 88.780 377.850 ;
        RECT 89.230 370.300 89.380 377.850 ;
        RECT 89.830 370.300 89.980 377.850 ;
        RECT 94.230 377.550 95.230 378.000 ;
        RECT 90.880 377.400 98.580 377.550 ;
        RECT 94.230 376.950 95.230 377.400 ;
        RECT 90.880 376.800 98.580 376.950 ;
        RECT 94.230 376.350 95.230 376.800 ;
        RECT 90.880 376.200 98.580 376.350 ;
        RECT 94.230 375.750 95.230 376.200 ;
        RECT 90.880 375.600 98.580 375.750 ;
        RECT 94.230 375.150 95.230 375.600 ;
        RECT 90.880 375.000 98.580 375.150 ;
        RECT 94.230 374.550 95.230 375.000 ;
        RECT 90.880 374.400 98.580 374.550 ;
        RECT 94.230 373.950 95.230 374.400 ;
        RECT 90.880 373.800 98.580 373.950 ;
        RECT 94.230 373.350 95.230 373.800 ;
        RECT 90.880 373.200 98.580 373.350 ;
        RECT 94.230 372.750 95.230 373.200 ;
        RECT 90.880 372.600 98.580 372.750 ;
        RECT 94.230 372.150 95.230 372.600 ;
        RECT 90.880 372.000 98.580 372.150 ;
        RECT 94.230 371.550 95.230 372.000 ;
        RECT 90.880 371.400 98.580 371.550 ;
        RECT 94.230 370.950 95.230 371.400 ;
        RECT 90.880 370.800 98.580 370.950 ;
        RECT 94.230 370.300 95.230 370.800 ;
        RECT 99.480 370.300 99.630 377.850 ;
        RECT 100.080 370.300 100.230 377.850 ;
        RECT 100.680 370.300 100.830 377.850 ;
        RECT 101.280 370.300 101.430 377.850 ;
        RECT 101.880 370.300 102.030 377.850 ;
        RECT 102.480 370.300 102.630 377.850 ;
        RECT 102.780 373.200 103.530 375.000 ;
        RECT 102.780 370.480 104.730 373.200 ;
        RECT 102.780 370.450 111.850 370.480 ;
        RECT 102.780 370.300 103.930 370.450 ;
        RECT 85.530 369.700 103.930 370.300 ;
        RECT 85.530 369.550 86.680 369.700 ;
        RECT 82.780 366.800 86.680 369.550 ;
        RECT 82.780 365.050 83.530 366.800 ;
        RECT 85.930 365.050 86.680 366.800 ;
        RECT 86.830 362.150 86.980 369.700 ;
        RECT 87.430 362.150 87.580 369.700 ;
        RECT 88.030 362.150 88.180 369.700 ;
        RECT 88.630 362.150 88.780 369.700 ;
        RECT 89.230 362.150 89.380 369.700 ;
        RECT 89.830 362.150 89.980 369.700 ;
        RECT 94.230 369.200 95.230 369.700 ;
        RECT 90.880 369.050 98.580 369.200 ;
        RECT 94.230 368.600 95.230 369.050 ;
        RECT 90.880 368.450 98.580 368.600 ;
        RECT 94.230 368.000 95.230 368.450 ;
        RECT 90.880 367.850 98.580 368.000 ;
        RECT 94.230 367.400 95.230 367.850 ;
        RECT 90.880 367.250 98.580 367.400 ;
        RECT 94.230 366.800 95.230 367.250 ;
        RECT 90.880 366.650 98.580 366.800 ;
        RECT 94.230 366.200 95.230 366.650 ;
        RECT 90.880 366.050 98.580 366.200 ;
        RECT 94.230 365.600 95.230 366.050 ;
        RECT 90.880 365.450 98.580 365.600 ;
        RECT 94.230 365.000 95.230 365.450 ;
        RECT 90.880 364.850 98.580 365.000 ;
        RECT 94.230 364.400 95.230 364.850 ;
        RECT 90.880 364.250 98.580 364.400 ;
        RECT 94.230 363.800 95.230 364.250 ;
        RECT 90.880 363.650 98.580 363.800 ;
        RECT 94.230 363.200 95.230 363.650 ;
        RECT 90.880 363.050 98.580 363.200 ;
        RECT 94.230 362.600 95.230 363.050 ;
        RECT 90.880 362.450 98.580 362.600 ;
        RECT 94.230 362.000 95.230 362.450 ;
        RECT 99.480 362.150 99.630 369.700 ;
        RECT 100.080 362.150 100.230 369.700 ;
        RECT 100.680 362.150 100.830 369.700 ;
        RECT 101.280 362.150 101.430 369.700 ;
        RECT 101.880 362.150 102.030 369.700 ;
        RECT 102.480 362.150 102.630 369.700 ;
        RECT 102.780 369.550 103.930 369.700 ;
        RECT 104.580 369.550 111.850 370.450 ;
        RECT 102.780 369.205 111.850 369.550 ;
        RECT 102.780 366.800 104.730 369.205 ;
        RECT 102.780 365.050 103.530 366.800 ;
        RECT 10.880 361.850 18.580 362.000 ;
        RECT 30.880 361.850 38.580 362.000 ;
        RECT 50.880 361.850 58.580 362.000 ;
        RECT 70.880 361.850 78.580 362.000 ;
        RECT 90.880 361.850 98.580 362.000 ;
        RECT 14.230 361.200 15.230 361.850 ;
        RECT 34.230 361.200 35.230 361.850 ;
        RECT 54.230 361.200 55.230 361.850 ;
        RECT 74.230 361.200 75.230 361.850 ;
        RECT 94.230 361.200 95.230 361.850 ;
        RECT 11.530 358.800 17.930 361.200 ;
        RECT 31.530 358.800 37.930 361.200 ;
        RECT 51.530 358.800 57.930 361.200 ;
        RECT 71.530 358.800 77.930 361.200 ;
        RECT 91.530 358.800 97.930 361.200 ;
        RECT 14.230 358.150 15.230 358.800 ;
        RECT 34.230 358.150 35.230 358.800 ;
        RECT 54.230 358.150 55.230 358.800 ;
        RECT 74.230 358.150 75.230 358.800 ;
        RECT 94.230 358.150 95.230 358.800 ;
        RECT 10.880 358.000 18.580 358.150 ;
        RECT 30.880 358.000 38.580 358.150 ;
        RECT 50.880 358.000 58.580 358.150 ;
        RECT 70.880 358.000 78.580 358.150 ;
        RECT 90.880 358.000 98.580 358.150 ;
        RECT 5.930 353.200 6.680 355.000 ;
        RECT 4.730 350.450 6.680 353.200 ;
        RECT 4.730 349.550 4.880 350.450 ;
        RECT 5.530 350.300 6.680 350.450 ;
        RECT 6.830 350.300 6.980 357.850 ;
        RECT 7.430 350.300 7.580 357.850 ;
        RECT 8.030 350.300 8.180 357.850 ;
        RECT 8.630 350.300 8.780 357.850 ;
        RECT 9.230 350.300 9.380 357.850 ;
        RECT 9.830 350.300 9.980 357.850 ;
        RECT 14.230 357.550 15.230 358.000 ;
        RECT 10.880 357.400 18.580 357.550 ;
        RECT 14.230 356.950 15.230 357.400 ;
        RECT 10.880 356.800 18.580 356.950 ;
        RECT 14.230 356.350 15.230 356.800 ;
        RECT 10.880 356.200 18.580 356.350 ;
        RECT 14.230 355.750 15.230 356.200 ;
        RECT 10.880 355.600 18.580 355.750 ;
        RECT 14.230 355.150 15.230 355.600 ;
        RECT 10.880 355.000 18.580 355.150 ;
        RECT 14.230 354.550 15.230 355.000 ;
        RECT 10.880 354.400 18.580 354.550 ;
        RECT 14.230 353.950 15.230 354.400 ;
        RECT 10.880 353.800 18.580 353.950 ;
        RECT 14.230 353.350 15.230 353.800 ;
        RECT 10.880 353.200 18.580 353.350 ;
        RECT 14.230 352.750 15.230 353.200 ;
        RECT 10.880 352.600 18.580 352.750 ;
        RECT 14.230 352.150 15.230 352.600 ;
        RECT 10.880 352.000 18.580 352.150 ;
        RECT 14.230 351.550 15.230 352.000 ;
        RECT 10.880 351.400 18.580 351.550 ;
        RECT 14.230 350.950 15.230 351.400 ;
        RECT 10.880 350.800 18.580 350.950 ;
        RECT 14.230 350.300 15.230 350.800 ;
        RECT 19.480 350.300 19.630 357.850 ;
        RECT 20.080 350.300 20.230 357.850 ;
        RECT 20.680 350.300 20.830 357.850 ;
        RECT 21.280 350.300 21.430 357.850 ;
        RECT 21.880 350.300 22.030 357.850 ;
        RECT 22.480 350.300 22.630 357.850 ;
        RECT 22.780 353.200 23.530 355.000 ;
        RECT 25.930 353.200 26.680 355.000 ;
        RECT 22.780 350.450 26.680 353.200 ;
        RECT 22.780 350.300 23.930 350.450 ;
        RECT 5.530 349.700 23.930 350.300 ;
        RECT 5.530 349.550 6.680 349.700 ;
        RECT 4.730 346.800 6.680 349.550 ;
        RECT 5.930 345.050 6.680 346.800 ;
        RECT 6.830 342.150 6.980 349.700 ;
        RECT 7.430 342.150 7.580 349.700 ;
        RECT 8.030 342.150 8.180 349.700 ;
        RECT 8.630 342.150 8.780 349.700 ;
        RECT 9.230 342.150 9.380 349.700 ;
        RECT 9.830 342.150 9.980 349.700 ;
        RECT 14.230 349.200 15.230 349.700 ;
        RECT 10.880 349.050 18.580 349.200 ;
        RECT 14.230 348.600 15.230 349.050 ;
        RECT 10.880 348.450 18.580 348.600 ;
        RECT 14.230 348.000 15.230 348.450 ;
        RECT 10.880 347.850 18.580 348.000 ;
        RECT 14.230 347.400 15.230 347.850 ;
        RECT 10.880 347.250 18.580 347.400 ;
        RECT 14.230 346.800 15.230 347.250 ;
        RECT 10.880 346.650 18.580 346.800 ;
        RECT 14.230 346.200 15.230 346.650 ;
        RECT 10.880 346.050 18.580 346.200 ;
        RECT 14.230 345.600 15.230 346.050 ;
        RECT 10.880 345.450 18.580 345.600 ;
        RECT 14.230 345.000 15.230 345.450 ;
        RECT 10.880 344.850 18.580 345.000 ;
        RECT 14.230 344.400 15.230 344.850 ;
        RECT 10.880 344.250 18.580 344.400 ;
        RECT 14.230 343.800 15.230 344.250 ;
        RECT 10.880 343.650 18.580 343.800 ;
        RECT 14.230 343.200 15.230 343.650 ;
        RECT 10.880 343.050 18.580 343.200 ;
        RECT 14.230 342.600 15.230 343.050 ;
        RECT 10.880 342.450 18.580 342.600 ;
        RECT 14.230 342.000 15.230 342.450 ;
        RECT 19.480 342.150 19.630 349.700 ;
        RECT 20.080 342.150 20.230 349.700 ;
        RECT 20.680 342.150 20.830 349.700 ;
        RECT 21.280 342.150 21.430 349.700 ;
        RECT 21.880 342.150 22.030 349.700 ;
        RECT 22.480 342.150 22.630 349.700 ;
        RECT 22.780 349.550 23.930 349.700 ;
        RECT 24.580 349.550 24.880 350.450 ;
        RECT 25.530 350.300 26.680 350.450 ;
        RECT 26.830 350.300 26.980 357.850 ;
        RECT 27.430 350.300 27.580 357.850 ;
        RECT 28.030 350.300 28.180 357.850 ;
        RECT 28.630 350.300 28.780 357.850 ;
        RECT 29.230 350.300 29.380 357.850 ;
        RECT 29.830 350.300 29.980 357.850 ;
        RECT 34.230 357.550 35.230 358.000 ;
        RECT 30.880 357.400 38.580 357.550 ;
        RECT 34.230 356.950 35.230 357.400 ;
        RECT 30.880 356.800 38.580 356.950 ;
        RECT 34.230 356.350 35.230 356.800 ;
        RECT 30.880 356.200 38.580 356.350 ;
        RECT 34.230 355.750 35.230 356.200 ;
        RECT 30.880 355.600 38.580 355.750 ;
        RECT 34.230 355.150 35.230 355.600 ;
        RECT 30.880 355.000 38.580 355.150 ;
        RECT 34.230 354.550 35.230 355.000 ;
        RECT 30.880 354.400 38.580 354.550 ;
        RECT 34.230 353.950 35.230 354.400 ;
        RECT 30.880 353.800 38.580 353.950 ;
        RECT 34.230 353.350 35.230 353.800 ;
        RECT 30.880 353.200 38.580 353.350 ;
        RECT 34.230 352.750 35.230 353.200 ;
        RECT 30.880 352.600 38.580 352.750 ;
        RECT 34.230 352.150 35.230 352.600 ;
        RECT 30.880 352.000 38.580 352.150 ;
        RECT 34.230 351.550 35.230 352.000 ;
        RECT 30.880 351.400 38.580 351.550 ;
        RECT 34.230 350.950 35.230 351.400 ;
        RECT 30.880 350.800 38.580 350.950 ;
        RECT 34.230 350.300 35.230 350.800 ;
        RECT 39.480 350.300 39.630 357.850 ;
        RECT 40.080 350.300 40.230 357.850 ;
        RECT 40.680 350.300 40.830 357.850 ;
        RECT 41.280 350.300 41.430 357.850 ;
        RECT 41.880 350.300 42.030 357.850 ;
        RECT 42.480 350.300 42.630 357.850 ;
        RECT 42.780 353.200 43.530 355.000 ;
        RECT 45.930 353.200 46.680 355.000 ;
        RECT 42.780 350.450 46.680 353.200 ;
        RECT 42.780 350.300 43.930 350.450 ;
        RECT 25.530 349.700 43.930 350.300 ;
        RECT 25.530 349.550 26.680 349.700 ;
        RECT 22.780 346.800 26.680 349.550 ;
        RECT 22.780 345.050 23.530 346.800 ;
        RECT 25.930 345.050 26.680 346.800 ;
        RECT 26.830 342.150 26.980 349.700 ;
        RECT 27.430 342.150 27.580 349.700 ;
        RECT 28.030 342.150 28.180 349.700 ;
        RECT 28.630 342.150 28.780 349.700 ;
        RECT 29.230 342.150 29.380 349.700 ;
        RECT 29.830 342.150 29.980 349.700 ;
        RECT 34.230 349.200 35.230 349.700 ;
        RECT 30.880 349.050 38.580 349.200 ;
        RECT 34.230 348.600 35.230 349.050 ;
        RECT 30.880 348.450 38.580 348.600 ;
        RECT 34.230 348.000 35.230 348.450 ;
        RECT 30.880 347.850 38.580 348.000 ;
        RECT 34.230 347.400 35.230 347.850 ;
        RECT 30.880 347.250 38.580 347.400 ;
        RECT 34.230 346.800 35.230 347.250 ;
        RECT 30.880 346.650 38.580 346.800 ;
        RECT 34.230 346.200 35.230 346.650 ;
        RECT 30.880 346.050 38.580 346.200 ;
        RECT 34.230 345.600 35.230 346.050 ;
        RECT 30.880 345.450 38.580 345.600 ;
        RECT 34.230 345.000 35.230 345.450 ;
        RECT 30.880 344.850 38.580 345.000 ;
        RECT 34.230 344.400 35.230 344.850 ;
        RECT 30.880 344.250 38.580 344.400 ;
        RECT 34.230 343.800 35.230 344.250 ;
        RECT 30.880 343.650 38.580 343.800 ;
        RECT 34.230 343.200 35.230 343.650 ;
        RECT 30.880 343.050 38.580 343.200 ;
        RECT 34.230 342.600 35.230 343.050 ;
        RECT 30.880 342.450 38.580 342.600 ;
        RECT 34.230 342.000 35.230 342.450 ;
        RECT 39.480 342.150 39.630 349.700 ;
        RECT 40.080 342.150 40.230 349.700 ;
        RECT 40.680 342.150 40.830 349.700 ;
        RECT 41.280 342.150 41.430 349.700 ;
        RECT 41.880 342.150 42.030 349.700 ;
        RECT 42.480 342.150 42.630 349.700 ;
        RECT 42.780 349.550 43.930 349.700 ;
        RECT 44.580 349.550 44.880 350.450 ;
        RECT 45.530 350.300 46.680 350.450 ;
        RECT 46.830 350.300 46.980 357.850 ;
        RECT 47.430 350.300 47.580 357.850 ;
        RECT 48.030 350.300 48.180 357.850 ;
        RECT 48.630 350.300 48.780 357.850 ;
        RECT 49.230 350.300 49.380 357.850 ;
        RECT 49.830 350.300 49.980 357.850 ;
        RECT 54.230 357.550 55.230 358.000 ;
        RECT 50.880 357.400 58.580 357.550 ;
        RECT 54.230 356.950 55.230 357.400 ;
        RECT 50.880 356.800 58.580 356.950 ;
        RECT 54.230 356.350 55.230 356.800 ;
        RECT 50.880 356.200 58.580 356.350 ;
        RECT 54.230 355.750 55.230 356.200 ;
        RECT 50.880 355.600 58.580 355.750 ;
        RECT 54.230 355.150 55.230 355.600 ;
        RECT 50.880 355.000 58.580 355.150 ;
        RECT 54.230 354.550 55.230 355.000 ;
        RECT 50.880 354.400 58.580 354.550 ;
        RECT 54.230 353.950 55.230 354.400 ;
        RECT 50.880 353.800 58.580 353.950 ;
        RECT 54.230 353.350 55.230 353.800 ;
        RECT 50.880 353.200 58.580 353.350 ;
        RECT 54.230 352.750 55.230 353.200 ;
        RECT 50.880 352.600 58.580 352.750 ;
        RECT 54.230 352.150 55.230 352.600 ;
        RECT 50.880 352.000 58.580 352.150 ;
        RECT 54.230 351.550 55.230 352.000 ;
        RECT 50.880 351.400 58.580 351.550 ;
        RECT 54.230 350.950 55.230 351.400 ;
        RECT 50.880 350.800 58.580 350.950 ;
        RECT 54.230 350.300 55.230 350.800 ;
        RECT 59.480 350.300 59.630 357.850 ;
        RECT 60.080 350.300 60.230 357.850 ;
        RECT 60.680 350.300 60.830 357.850 ;
        RECT 61.280 350.300 61.430 357.850 ;
        RECT 61.880 350.300 62.030 357.850 ;
        RECT 62.480 350.300 62.630 357.850 ;
        RECT 62.780 353.200 63.530 355.000 ;
        RECT 65.930 353.200 66.680 355.000 ;
        RECT 62.780 350.450 66.680 353.200 ;
        RECT 62.780 350.300 63.930 350.450 ;
        RECT 45.530 349.700 63.930 350.300 ;
        RECT 45.530 349.550 46.680 349.700 ;
        RECT 42.780 346.800 46.680 349.550 ;
        RECT 42.780 345.050 43.530 346.800 ;
        RECT 45.930 345.050 46.680 346.800 ;
        RECT 46.830 342.150 46.980 349.700 ;
        RECT 47.430 342.150 47.580 349.700 ;
        RECT 48.030 342.150 48.180 349.700 ;
        RECT 48.630 342.150 48.780 349.700 ;
        RECT 49.230 342.150 49.380 349.700 ;
        RECT 49.830 342.150 49.980 349.700 ;
        RECT 54.230 349.200 55.230 349.700 ;
        RECT 50.880 349.050 58.580 349.200 ;
        RECT 54.230 348.600 55.230 349.050 ;
        RECT 50.880 348.450 58.580 348.600 ;
        RECT 54.230 348.000 55.230 348.450 ;
        RECT 50.880 347.850 58.580 348.000 ;
        RECT 54.230 347.400 55.230 347.850 ;
        RECT 50.880 347.250 58.580 347.400 ;
        RECT 54.230 346.800 55.230 347.250 ;
        RECT 50.880 346.650 58.580 346.800 ;
        RECT 54.230 346.200 55.230 346.650 ;
        RECT 50.880 346.050 58.580 346.200 ;
        RECT 54.230 345.600 55.230 346.050 ;
        RECT 50.880 345.450 58.580 345.600 ;
        RECT 54.230 345.000 55.230 345.450 ;
        RECT 50.880 344.850 58.580 345.000 ;
        RECT 54.230 344.400 55.230 344.850 ;
        RECT 50.880 344.250 58.580 344.400 ;
        RECT 54.230 343.800 55.230 344.250 ;
        RECT 50.880 343.650 58.580 343.800 ;
        RECT 54.230 343.200 55.230 343.650 ;
        RECT 50.880 343.050 58.580 343.200 ;
        RECT 54.230 342.600 55.230 343.050 ;
        RECT 50.880 342.450 58.580 342.600 ;
        RECT 54.230 342.000 55.230 342.450 ;
        RECT 59.480 342.150 59.630 349.700 ;
        RECT 60.080 342.150 60.230 349.700 ;
        RECT 60.680 342.150 60.830 349.700 ;
        RECT 61.280 342.150 61.430 349.700 ;
        RECT 61.880 342.150 62.030 349.700 ;
        RECT 62.480 342.150 62.630 349.700 ;
        RECT 62.780 349.550 63.930 349.700 ;
        RECT 64.580 349.550 64.880 350.450 ;
        RECT 65.530 350.300 66.680 350.450 ;
        RECT 66.830 350.300 66.980 357.850 ;
        RECT 67.430 350.300 67.580 357.850 ;
        RECT 68.030 350.300 68.180 357.850 ;
        RECT 68.630 350.300 68.780 357.850 ;
        RECT 69.230 350.300 69.380 357.850 ;
        RECT 69.830 350.300 69.980 357.850 ;
        RECT 74.230 357.550 75.230 358.000 ;
        RECT 70.880 357.400 78.580 357.550 ;
        RECT 74.230 356.950 75.230 357.400 ;
        RECT 70.880 356.800 78.580 356.950 ;
        RECT 74.230 356.350 75.230 356.800 ;
        RECT 70.880 356.200 78.580 356.350 ;
        RECT 74.230 355.750 75.230 356.200 ;
        RECT 70.880 355.600 78.580 355.750 ;
        RECT 74.230 355.150 75.230 355.600 ;
        RECT 70.880 355.000 78.580 355.150 ;
        RECT 74.230 354.550 75.230 355.000 ;
        RECT 70.880 354.400 78.580 354.550 ;
        RECT 74.230 353.950 75.230 354.400 ;
        RECT 70.880 353.800 78.580 353.950 ;
        RECT 74.230 353.350 75.230 353.800 ;
        RECT 70.880 353.200 78.580 353.350 ;
        RECT 74.230 352.750 75.230 353.200 ;
        RECT 70.880 352.600 78.580 352.750 ;
        RECT 74.230 352.150 75.230 352.600 ;
        RECT 70.880 352.000 78.580 352.150 ;
        RECT 74.230 351.550 75.230 352.000 ;
        RECT 70.880 351.400 78.580 351.550 ;
        RECT 74.230 350.950 75.230 351.400 ;
        RECT 70.880 350.800 78.580 350.950 ;
        RECT 74.230 350.300 75.230 350.800 ;
        RECT 79.480 350.300 79.630 357.850 ;
        RECT 80.080 350.300 80.230 357.850 ;
        RECT 80.680 350.300 80.830 357.850 ;
        RECT 81.280 350.300 81.430 357.850 ;
        RECT 81.880 350.300 82.030 357.850 ;
        RECT 82.480 350.300 82.630 357.850 ;
        RECT 82.780 353.200 83.530 355.000 ;
        RECT 85.930 353.200 86.680 355.000 ;
        RECT 82.780 350.450 86.680 353.200 ;
        RECT 82.780 350.300 83.930 350.450 ;
        RECT 65.530 349.700 83.930 350.300 ;
        RECT 65.530 349.550 66.680 349.700 ;
        RECT 62.780 346.800 66.680 349.550 ;
        RECT 62.780 345.050 63.530 346.800 ;
        RECT 65.930 345.050 66.680 346.800 ;
        RECT 66.830 342.150 66.980 349.700 ;
        RECT 67.430 342.150 67.580 349.700 ;
        RECT 68.030 342.150 68.180 349.700 ;
        RECT 68.630 342.150 68.780 349.700 ;
        RECT 69.230 342.150 69.380 349.700 ;
        RECT 69.830 342.150 69.980 349.700 ;
        RECT 74.230 349.200 75.230 349.700 ;
        RECT 70.880 349.050 78.580 349.200 ;
        RECT 74.230 348.600 75.230 349.050 ;
        RECT 70.880 348.450 78.580 348.600 ;
        RECT 74.230 348.000 75.230 348.450 ;
        RECT 70.880 347.850 78.580 348.000 ;
        RECT 74.230 347.400 75.230 347.850 ;
        RECT 70.880 347.250 78.580 347.400 ;
        RECT 74.230 346.800 75.230 347.250 ;
        RECT 70.880 346.650 78.580 346.800 ;
        RECT 74.230 346.200 75.230 346.650 ;
        RECT 70.880 346.050 78.580 346.200 ;
        RECT 74.230 345.600 75.230 346.050 ;
        RECT 70.880 345.450 78.580 345.600 ;
        RECT 74.230 345.000 75.230 345.450 ;
        RECT 70.880 344.850 78.580 345.000 ;
        RECT 74.230 344.400 75.230 344.850 ;
        RECT 70.880 344.250 78.580 344.400 ;
        RECT 74.230 343.800 75.230 344.250 ;
        RECT 70.880 343.650 78.580 343.800 ;
        RECT 74.230 343.200 75.230 343.650 ;
        RECT 70.880 343.050 78.580 343.200 ;
        RECT 74.230 342.600 75.230 343.050 ;
        RECT 70.880 342.450 78.580 342.600 ;
        RECT 74.230 342.000 75.230 342.450 ;
        RECT 79.480 342.150 79.630 349.700 ;
        RECT 80.080 342.150 80.230 349.700 ;
        RECT 80.680 342.150 80.830 349.700 ;
        RECT 81.280 342.150 81.430 349.700 ;
        RECT 81.880 342.150 82.030 349.700 ;
        RECT 82.480 342.150 82.630 349.700 ;
        RECT 82.780 349.550 83.930 349.700 ;
        RECT 84.580 349.550 84.880 350.450 ;
        RECT 85.530 350.300 86.680 350.450 ;
        RECT 86.830 350.300 86.980 357.850 ;
        RECT 87.430 350.300 87.580 357.850 ;
        RECT 88.030 350.300 88.180 357.850 ;
        RECT 88.630 350.300 88.780 357.850 ;
        RECT 89.230 350.300 89.380 357.850 ;
        RECT 89.830 350.300 89.980 357.850 ;
        RECT 94.230 357.550 95.230 358.000 ;
        RECT 90.880 357.400 98.580 357.550 ;
        RECT 94.230 356.950 95.230 357.400 ;
        RECT 90.880 356.800 98.580 356.950 ;
        RECT 94.230 356.350 95.230 356.800 ;
        RECT 90.880 356.200 98.580 356.350 ;
        RECT 94.230 355.750 95.230 356.200 ;
        RECT 90.880 355.600 98.580 355.750 ;
        RECT 94.230 355.150 95.230 355.600 ;
        RECT 90.880 355.000 98.580 355.150 ;
        RECT 94.230 354.550 95.230 355.000 ;
        RECT 90.880 354.400 98.580 354.550 ;
        RECT 94.230 353.950 95.230 354.400 ;
        RECT 90.880 353.800 98.580 353.950 ;
        RECT 94.230 353.350 95.230 353.800 ;
        RECT 90.880 353.200 98.580 353.350 ;
        RECT 94.230 352.750 95.230 353.200 ;
        RECT 90.880 352.600 98.580 352.750 ;
        RECT 94.230 352.150 95.230 352.600 ;
        RECT 90.880 352.000 98.580 352.150 ;
        RECT 94.230 351.550 95.230 352.000 ;
        RECT 90.880 351.400 98.580 351.550 ;
        RECT 94.230 350.950 95.230 351.400 ;
        RECT 90.880 350.800 98.580 350.950 ;
        RECT 94.230 350.300 95.230 350.800 ;
        RECT 99.480 350.300 99.630 357.850 ;
        RECT 100.080 350.300 100.230 357.850 ;
        RECT 100.680 350.300 100.830 357.850 ;
        RECT 101.280 350.300 101.430 357.850 ;
        RECT 101.880 350.300 102.030 357.850 ;
        RECT 102.480 350.300 102.630 357.850 ;
        RECT 102.780 353.200 103.530 355.000 ;
        RECT 102.780 350.480 104.730 353.200 ;
        RECT 102.780 350.450 111.850 350.480 ;
        RECT 102.780 350.300 103.930 350.450 ;
        RECT 85.530 349.700 103.930 350.300 ;
        RECT 85.530 349.550 86.680 349.700 ;
        RECT 82.780 346.800 86.680 349.550 ;
        RECT 82.780 345.050 83.530 346.800 ;
        RECT 85.930 345.050 86.680 346.800 ;
        RECT 86.830 342.150 86.980 349.700 ;
        RECT 87.430 342.150 87.580 349.700 ;
        RECT 88.030 342.150 88.180 349.700 ;
        RECT 88.630 342.150 88.780 349.700 ;
        RECT 89.230 342.150 89.380 349.700 ;
        RECT 89.830 342.150 89.980 349.700 ;
        RECT 94.230 349.200 95.230 349.700 ;
        RECT 90.880 349.050 98.580 349.200 ;
        RECT 94.230 348.600 95.230 349.050 ;
        RECT 90.880 348.450 98.580 348.600 ;
        RECT 94.230 348.000 95.230 348.450 ;
        RECT 90.880 347.850 98.580 348.000 ;
        RECT 94.230 347.400 95.230 347.850 ;
        RECT 90.880 347.250 98.580 347.400 ;
        RECT 94.230 346.800 95.230 347.250 ;
        RECT 90.880 346.650 98.580 346.800 ;
        RECT 94.230 346.200 95.230 346.650 ;
        RECT 90.880 346.050 98.580 346.200 ;
        RECT 94.230 345.600 95.230 346.050 ;
        RECT 90.880 345.450 98.580 345.600 ;
        RECT 94.230 345.000 95.230 345.450 ;
        RECT 90.880 344.850 98.580 345.000 ;
        RECT 94.230 344.400 95.230 344.850 ;
        RECT 90.880 344.250 98.580 344.400 ;
        RECT 94.230 343.800 95.230 344.250 ;
        RECT 90.880 343.650 98.580 343.800 ;
        RECT 94.230 343.200 95.230 343.650 ;
        RECT 90.880 343.050 98.580 343.200 ;
        RECT 94.230 342.600 95.230 343.050 ;
        RECT 90.880 342.450 98.580 342.600 ;
        RECT 94.230 342.000 95.230 342.450 ;
        RECT 99.480 342.150 99.630 349.700 ;
        RECT 100.080 342.150 100.230 349.700 ;
        RECT 100.680 342.150 100.830 349.700 ;
        RECT 101.280 342.150 101.430 349.700 ;
        RECT 101.880 342.150 102.030 349.700 ;
        RECT 102.480 342.150 102.630 349.700 ;
        RECT 102.780 349.550 103.930 349.700 ;
        RECT 104.580 349.550 111.850 350.450 ;
        RECT 102.780 349.205 111.850 349.550 ;
        RECT 102.780 346.800 104.730 349.205 ;
        RECT 102.780 345.050 103.530 346.800 ;
        RECT 10.880 341.850 18.580 342.000 ;
        RECT 30.880 341.850 38.580 342.000 ;
        RECT 50.880 341.850 58.580 342.000 ;
        RECT 70.880 341.850 78.580 342.000 ;
        RECT 90.880 341.850 98.580 342.000 ;
        RECT 14.230 341.200 15.230 341.850 ;
        RECT 34.230 341.200 35.230 341.850 ;
        RECT 54.230 341.200 55.230 341.850 ;
        RECT 74.230 341.200 75.230 341.850 ;
        RECT 94.230 341.200 95.230 341.850 ;
        RECT 11.530 338.800 17.930 341.200 ;
        RECT 31.530 338.800 37.930 341.200 ;
        RECT 51.530 338.800 57.930 341.200 ;
        RECT 71.530 338.800 77.930 341.200 ;
        RECT 91.530 338.800 97.930 341.200 ;
        RECT 14.230 338.150 15.230 338.800 ;
        RECT 34.230 338.150 35.230 338.800 ;
        RECT 54.230 338.150 55.230 338.800 ;
        RECT 74.230 338.150 75.230 338.800 ;
        RECT 94.230 338.150 95.230 338.800 ;
        RECT 10.880 338.000 18.580 338.150 ;
        RECT 30.880 338.000 38.580 338.150 ;
        RECT 50.880 338.000 58.580 338.150 ;
        RECT 70.880 338.000 78.580 338.150 ;
        RECT 90.880 338.000 98.580 338.150 ;
        RECT 5.930 333.200 6.680 335.000 ;
        RECT 4.730 330.450 6.680 333.200 ;
        RECT 4.730 329.550 4.880 330.450 ;
        RECT 5.530 330.300 6.680 330.450 ;
        RECT 6.830 330.300 6.980 337.850 ;
        RECT 7.430 330.300 7.580 337.850 ;
        RECT 8.030 330.300 8.180 337.850 ;
        RECT 8.630 330.300 8.780 337.850 ;
        RECT 9.230 330.300 9.380 337.850 ;
        RECT 9.830 330.300 9.980 337.850 ;
        RECT 14.230 337.550 15.230 338.000 ;
        RECT 10.880 337.400 18.580 337.550 ;
        RECT 14.230 336.950 15.230 337.400 ;
        RECT 10.880 336.800 18.580 336.950 ;
        RECT 14.230 336.350 15.230 336.800 ;
        RECT 10.880 336.200 18.580 336.350 ;
        RECT 14.230 335.750 15.230 336.200 ;
        RECT 10.880 335.600 18.580 335.750 ;
        RECT 14.230 335.150 15.230 335.600 ;
        RECT 10.880 335.000 18.580 335.150 ;
        RECT 14.230 334.550 15.230 335.000 ;
        RECT 10.880 334.400 18.580 334.550 ;
        RECT 14.230 333.950 15.230 334.400 ;
        RECT 10.880 333.800 18.580 333.950 ;
        RECT 14.230 333.350 15.230 333.800 ;
        RECT 10.880 333.200 18.580 333.350 ;
        RECT 14.230 332.750 15.230 333.200 ;
        RECT 10.880 332.600 18.580 332.750 ;
        RECT 14.230 332.150 15.230 332.600 ;
        RECT 10.880 332.000 18.580 332.150 ;
        RECT 14.230 331.550 15.230 332.000 ;
        RECT 10.880 331.400 18.580 331.550 ;
        RECT 14.230 330.950 15.230 331.400 ;
        RECT 10.880 330.800 18.580 330.950 ;
        RECT 14.230 330.300 15.230 330.800 ;
        RECT 19.480 330.300 19.630 337.850 ;
        RECT 20.080 330.300 20.230 337.850 ;
        RECT 20.680 330.300 20.830 337.850 ;
        RECT 21.280 330.300 21.430 337.850 ;
        RECT 21.880 330.300 22.030 337.850 ;
        RECT 22.480 330.300 22.630 337.850 ;
        RECT 22.780 333.200 23.530 335.000 ;
        RECT 25.930 333.200 26.680 335.000 ;
        RECT 22.780 330.450 26.680 333.200 ;
        RECT 22.780 330.300 23.930 330.450 ;
        RECT 5.530 329.700 23.930 330.300 ;
        RECT 5.530 329.550 6.680 329.700 ;
        RECT 4.730 326.800 6.680 329.550 ;
        RECT 5.930 325.050 6.680 326.800 ;
        RECT 6.830 322.150 6.980 329.700 ;
        RECT 7.430 322.150 7.580 329.700 ;
        RECT 8.030 322.150 8.180 329.700 ;
        RECT 8.630 322.150 8.780 329.700 ;
        RECT 9.230 322.150 9.380 329.700 ;
        RECT 9.830 322.150 9.980 329.700 ;
        RECT 14.230 329.200 15.230 329.700 ;
        RECT 10.880 329.050 18.580 329.200 ;
        RECT 14.230 328.600 15.230 329.050 ;
        RECT 10.880 328.450 18.580 328.600 ;
        RECT 14.230 328.000 15.230 328.450 ;
        RECT 10.880 327.850 18.580 328.000 ;
        RECT 14.230 327.400 15.230 327.850 ;
        RECT 10.880 327.250 18.580 327.400 ;
        RECT 14.230 326.800 15.230 327.250 ;
        RECT 10.880 326.650 18.580 326.800 ;
        RECT 14.230 326.200 15.230 326.650 ;
        RECT 10.880 326.050 18.580 326.200 ;
        RECT 14.230 325.600 15.230 326.050 ;
        RECT 10.880 325.450 18.580 325.600 ;
        RECT 14.230 325.000 15.230 325.450 ;
        RECT 10.880 324.850 18.580 325.000 ;
        RECT 14.230 324.400 15.230 324.850 ;
        RECT 10.880 324.250 18.580 324.400 ;
        RECT 14.230 323.800 15.230 324.250 ;
        RECT 10.880 323.650 18.580 323.800 ;
        RECT 14.230 323.200 15.230 323.650 ;
        RECT 10.880 323.050 18.580 323.200 ;
        RECT 14.230 322.600 15.230 323.050 ;
        RECT 10.880 322.450 18.580 322.600 ;
        RECT 14.230 322.000 15.230 322.450 ;
        RECT 19.480 322.150 19.630 329.700 ;
        RECT 20.080 322.150 20.230 329.700 ;
        RECT 20.680 322.150 20.830 329.700 ;
        RECT 21.280 322.150 21.430 329.700 ;
        RECT 21.880 322.150 22.030 329.700 ;
        RECT 22.480 322.150 22.630 329.700 ;
        RECT 22.780 329.550 23.930 329.700 ;
        RECT 24.580 329.550 24.880 330.450 ;
        RECT 25.530 330.300 26.680 330.450 ;
        RECT 26.830 330.300 26.980 337.850 ;
        RECT 27.430 330.300 27.580 337.850 ;
        RECT 28.030 330.300 28.180 337.850 ;
        RECT 28.630 330.300 28.780 337.850 ;
        RECT 29.230 330.300 29.380 337.850 ;
        RECT 29.830 330.300 29.980 337.850 ;
        RECT 34.230 337.550 35.230 338.000 ;
        RECT 30.880 337.400 38.580 337.550 ;
        RECT 34.230 336.950 35.230 337.400 ;
        RECT 30.880 336.800 38.580 336.950 ;
        RECT 34.230 336.350 35.230 336.800 ;
        RECT 30.880 336.200 38.580 336.350 ;
        RECT 34.230 335.750 35.230 336.200 ;
        RECT 30.880 335.600 38.580 335.750 ;
        RECT 34.230 335.150 35.230 335.600 ;
        RECT 30.880 335.000 38.580 335.150 ;
        RECT 34.230 334.550 35.230 335.000 ;
        RECT 30.880 334.400 38.580 334.550 ;
        RECT 34.230 333.950 35.230 334.400 ;
        RECT 30.880 333.800 38.580 333.950 ;
        RECT 34.230 333.350 35.230 333.800 ;
        RECT 30.880 333.200 38.580 333.350 ;
        RECT 34.230 332.750 35.230 333.200 ;
        RECT 30.880 332.600 38.580 332.750 ;
        RECT 34.230 332.150 35.230 332.600 ;
        RECT 30.880 332.000 38.580 332.150 ;
        RECT 34.230 331.550 35.230 332.000 ;
        RECT 30.880 331.400 38.580 331.550 ;
        RECT 34.230 330.950 35.230 331.400 ;
        RECT 30.880 330.800 38.580 330.950 ;
        RECT 34.230 330.300 35.230 330.800 ;
        RECT 39.480 330.300 39.630 337.850 ;
        RECT 40.080 330.300 40.230 337.850 ;
        RECT 40.680 330.300 40.830 337.850 ;
        RECT 41.280 330.300 41.430 337.850 ;
        RECT 41.880 330.300 42.030 337.850 ;
        RECT 42.480 330.300 42.630 337.850 ;
        RECT 42.780 333.200 43.530 335.000 ;
        RECT 45.930 333.200 46.680 335.000 ;
        RECT 42.780 330.450 46.680 333.200 ;
        RECT 42.780 330.300 43.930 330.450 ;
        RECT 25.530 329.700 43.930 330.300 ;
        RECT 25.530 329.550 26.680 329.700 ;
        RECT 22.780 326.800 26.680 329.550 ;
        RECT 22.780 325.050 23.530 326.800 ;
        RECT 25.930 325.050 26.680 326.800 ;
        RECT 26.830 322.150 26.980 329.700 ;
        RECT 27.430 322.150 27.580 329.700 ;
        RECT 28.030 322.150 28.180 329.700 ;
        RECT 28.630 322.150 28.780 329.700 ;
        RECT 29.230 322.150 29.380 329.700 ;
        RECT 29.830 322.150 29.980 329.700 ;
        RECT 34.230 329.200 35.230 329.700 ;
        RECT 30.880 329.050 38.580 329.200 ;
        RECT 34.230 328.600 35.230 329.050 ;
        RECT 30.880 328.450 38.580 328.600 ;
        RECT 34.230 328.000 35.230 328.450 ;
        RECT 30.880 327.850 38.580 328.000 ;
        RECT 34.230 327.400 35.230 327.850 ;
        RECT 30.880 327.250 38.580 327.400 ;
        RECT 34.230 326.800 35.230 327.250 ;
        RECT 30.880 326.650 38.580 326.800 ;
        RECT 34.230 326.200 35.230 326.650 ;
        RECT 30.880 326.050 38.580 326.200 ;
        RECT 34.230 325.600 35.230 326.050 ;
        RECT 30.880 325.450 38.580 325.600 ;
        RECT 34.230 325.000 35.230 325.450 ;
        RECT 30.880 324.850 38.580 325.000 ;
        RECT 34.230 324.400 35.230 324.850 ;
        RECT 30.880 324.250 38.580 324.400 ;
        RECT 34.230 323.800 35.230 324.250 ;
        RECT 30.880 323.650 38.580 323.800 ;
        RECT 34.230 323.200 35.230 323.650 ;
        RECT 30.880 323.050 38.580 323.200 ;
        RECT 34.230 322.600 35.230 323.050 ;
        RECT 30.880 322.450 38.580 322.600 ;
        RECT 34.230 322.000 35.230 322.450 ;
        RECT 39.480 322.150 39.630 329.700 ;
        RECT 40.080 322.150 40.230 329.700 ;
        RECT 40.680 322.150 40.830 329.700 ;
        RECT 41.280 322.150 41.430 329.700 ;
        RECT 41.880 322.150 42.030 329.700 ;
        RECT 42.480 322.150 42.630 329.700 ;
        RECT 42.780 329.550 43.930 329.700 ;
        RECT 44.580 329.550 44.880 330.450 ;
        RECT 45.530 330.300 46.680 330.450 ;
        RECT 46.830 330.300 46.980 337.850 ;
        RECT 47.430 330.300 47.580 337.850 ;
        RECT 48.030 330.300 48.180 337.850 ;
        RECT 48.630 330.300 48.780 337.850 ;
        RECT 49.230 330.300 49.380 337.850 ;
        RECT 49.830 330.300 49.980 337.850 ;
        RECT 54.230 337.550 55.230 338.000 ;
        RECT 50.880 337.400 58.580 337.550 ;
        RECT 54.230 336.950 55.230 337.400 ;
        RECT 50.880 336.800 58.580 336.950 ;
        RECT 54.230 336.350 55.230 336.800 ;
        RECT 50.880 336.200 58.580 336.350 ;
        RECT 54.230 335.750 55.230 336.200 ;
        RECT 50.880 335.600 58.580 335.750 ;
        RECT 54.230 335.150 55.230 335.600 ;
        RECT 50.880 335.000 58.580 335.150 ;
        RECT 54.230 334.550 55.230 335.000 ;
        RECT 50.880 334.400 58.580 334.550 ;
        RECT 54.230 333.950 55.230 334.400 ;
        RECT 50.880 333.800 58.580 333.950 ;
        RECT 54.230 333.350 55.230 333.800 ;
        RECT 50.880 333.200 58.580 333.350 ;
        RECT 54.230 332.750 55.230 333.200 ;
        RECT 50.880 332.600 58.580 332.750 ;
        RECT 54.230 332.150 55.230 332.600 ;
        RECT 50.880 332.000 58.580 332.150 ;
        RECT 54.230 331.550 55.230 332.000 ;
        RECT 50.880 331.400 58.580 331.550 ;
        RECT 54.230 330.950 55.230 331.400 ;
        RECT 50.880 330.800 58.580 330.950 ;
        RECT 54.230 330.300 55.230 330.800 ;
        RECT 59.480 330.300 59.630 337.850 ;
        RECT 60.080 330.300 60.230 337.850 ;
        RECT 60.680 330.300 60.830 337.850 ;
        RECT 61.280 330.300 61.430 337.850 ;
        RECT 61.880 330.300 62.030 337.850 ;
        RECT 62.480 330.300 62.630 337.850 ;
        RECT 62.780 333.200 63.530 335.000 ;
        RECT 65.930 333.200 66.680 335.000 ;
        RECT 62.780 330.450 66.680 333.200 ;
        RECT 62.780 330.300 63.930 330.450 ;
        RECT 45.530 329.700 63.930 330.300 ;
        RECT 45.530 329.550 46.680 329.700 ;
        RECT 42.780 326.800 46.680 329.550 ;
        RECT 42.780 325.050 43.530 326.800 ;
        RECT 45.930 325.050 46.680 326.800 ;
        RECT 46.830 322.150 46.980 329.700 ;
        RECT 47.430 322.150 47.580 329.700 ;
        RECT 48.030 322.150 48.180 329.700 ;
        RECT 48.630 322.150 48.780 329.700 ;
        RECT 49.230 322.150 49.380 329.700 ;
        RECT 49.830 322.150 49.980 329.700 ;
        RECT 54.230 329.200 55.230 329.700 ;
        RECT 50.880 329.050 58.580 329.200 ;
        RECT 54.230 328.600 55.230 329.050 ;
        RECT 50.880 328.450 58.580 328.600 ;
        RECT 54.230 328.000 55.230 328.450 ;
        RECT 50.880 327.850 58.580 328.000 ;
        RECT 54.230 327.400 55.230 327.850 ;
        RECT 50.880 327.250 58.580 327.400 ;
        RECT 54.230 326.800 55.230 327.250 ;
        RECT 50.880 326.650 58.580 326.800 ;
        RECT 54.230 326.200 55.230 326.650 ;
        RECT 50.880 326.050 58.580 326.200 ;
        RECT 54.230 325.600 55.230 326.050 ;
        RECT 50.880 325.450 58.580 325.600 ;
        RECT 54.230 325.000 55.230 325.450 ;
        RECT 50.880 324.850 58.580 325.000 ;
        RECT 54.230 324.400 55.230 324.850 ;
        RECT 50.880 324.250 58.580 324.400 ;
        RECT 54.230 323.800 55.230 324.250 ;
        RECT 50.880 323.650 58.580 323.800 ;
        RECT 54.230 323.200 55.230 323.650 ;
        RECT 50.880 323.050 58.580 323.200 ;
        RECT 54.230 322.600 55.230 323.050 ;
        RECT 50.880 322.450 58.580 322.600 ;
        RECT 54.230 322.000 55.230 322.450 ;
        RECT 59.480 322.150 59.630 329.700 ;
        RECT 60.080 322.150 60.230 329.700 ;
        RECT 60.680 322.150 60.830 329.700 ;
        RECT 61.280 322.150 61.430 329.700 ;
        RECT 61.880 322.150 62.030 329.700 ;
        RECT 62.480 322.150 62.630 329.700 ;
        RECT 62.780 329.550 63.930 329.700 ;
        RECT 64.580 329.550 64.880 330.450 ;
        RECT 65.530 330.300 66.680 330.450 ;
        RECT 66.830 330.300 66.980 337.850 ;
        RECT 67.430 330.300 67.580 337.850 ;
        RECT 68.030 330.300 68.180 337.850 ;
        RECT 68.630 330.300 68.780 337.850 ;
        RECT 69.230 330.300 69.380 337.850 ;
        RECT 69.830 330.300 69.980 337.850 ;
        RECT 74.230 337.550 75.230 338.000 ;
        RECT 70.880 337.400 78.580 337.550 ;
        RECT 74.230 336.950 75.230 337.400 ;
        RECT 70.880 336.800 78.580 336.950 ;
        RECT 74.230 336.350 75.230 336.800 ;
        RECT 70.880 336.200 78.580 336.350 ;
        RECT 74.230 335.750 75.230 336.200 ;
        RECT 70.880 335.600 78.580 335.750 ;
        RECT 74.230 335.150 75.230 335.600 ;
        RECT 70.880 335.000 78.580 335.150 ;
        RECT 74.230 334.550 75.230 335.000 ;
        RECT 70.880 334.400 78.580 334.550 ;
        RECT 74.230 333.950 75.230 334.400 ;
        RECT 70.880 333.800 78.580 333.950 ;
        RECT 74.230 333.350 75.230 333.800 ;
        RECT 70.880 333.200 78.580 333.350 ;
        RECT 74.230 332.750 75.230 333.200 ;
        RECT 70.880 332.600 78.580 332.750 ;
        RECT 74.230 332.150 75.230 332.600 ;
        RECT 70.880 332.000 78.580 332.150 ;
        RECT 74.230 331.550 75.230 332.000 ;
        RECT 70.880 331.400 78.580 331.550 ;
        RECT 74.230 330.950 75.230 331.400 ;
        RECT 70.880 330.800 78.580 330.950 ;
        RECT 74.230 330.300 75.230 330.800 ;
        RECT 79.480 330.300 79.630 337.850 ;
        RECT 80.080 330.300 80.230 337.850 ;
        RECT 80.680 330.300 80.830 337.850 ;
        RECT 81.280 330.300 81.430 337.850 ;
        RECT 81.880 330.300 82.030 337.850 ;
        RECT 82.480 330.300 82.630 337.850 ;
        RECT 82.780 333.200 83.530 335.000 ;
        RECT 85.930 333.200 86.680 335.000 ;
        RECT 82.780 330.450 86.680 333.200 ;
        RECT 82.780 330.300 83.930 330.450 ;
        RECT 65.530 329.700 83.930 330.300 ;
        RECT 65.530 329.550 66.680 329.700 ;
        RECT 62.780 326.800 66.680 329.550 ;
        RECT 62.780 325.050 63.530 326.800 ;
        RECT 65.930 325.050 66.680 326.800 ;
        RECT 66.830 322.150 66.980 329.700 ;
        RECT 67.430 322.150 67.580 329.700 ;
        RECT 68.030 322.150 68.180 329.700 ;
        RECT 68.630 322.150 68.780 329.700 ;
        RECT 69.230 322.150 69.380 329.700 ;
        RECT 69.830 322.150 69.980 329.700 ;
        RECT 74.230 329.200 75.230 329.700 ;
        RECT 70.880 329.050 78.580 329.200 ;
        RECT 74.230 328.600 75.230 329.050 ;
        RECT 70.880 328.450 78.580 328.600 ;
        RECT 74.230 328.000 75.230 328.450 ;
        RECT 70.880 327.850 78.580 328.000 ;
        RECT 74.230 327.400 75.230 327.850 ;
        RECT 70.880 327.250 78.580 327.400 ;
        RECT 74.230 326.800 75.230 327.250 ;
        RECT 70.880 326.650 78.580 326.800 ;
        RECT 74.230 326.200 75.230 326.650 ;
        RECT 70.880 326.050 78.580 326.200 ;
        RECT 74.230 325.600 75.230 326.050 ;
        RECT 70.880 325.450 78.580 325.600 ;
        RECT 74.230 325.000 75.230 325.450 ;
        RECT 70.880 324.850 78.580 325.000 ;
        RECT 74.230 324.400 75.230 324.850 ;
        RECT 70.880 324.250 78.580 324.400 ;
        RECT 74.230 323.800 75.230 324.250 ;
        RECT 70.880 323.650 78.580 323.800 ;
        RECT 74.230 323.200 75.230 323.650 ;
        RECT 70.880 323.050 78.580 323.200 ;
        RECT 74.230 322.600 75.230 323.050 ;
        RECT 70.880 322.450 78.580 322.600 ;
        RECT 74.230 322.000 75.230 322.450 ;
        RECT 79.480 322.150 79.630 329.700 ;
        RECT 80.080 322.150 80.230 329.700 ;
        RECT 80.680 322.150 80.830 329.700 ;
        RECT 81.280 322.150 81.430 329.700 ;
        RECT 81.880 322.150 82.030 329.700 ;
        RECT 82.480 322.150 82.630 329.700 ;
        RECT 82.780 329.550 83.930 329.700 ;
        RECT 84.580 329.550 84.880 330.450 ;
        RECT 85.530 330.300 86.680 330.450 ;
        RECT 86.830 330.300 86.980 337.850 ;
        RECT 87.430 330.300 87.580 337.850 ;
        RECT 88.030 330.300 88.180 337.850 ;
        RECT 88.630 330.300 88.780 337.850 ;
        RECT 89.230 330.300 89.380 337.850 ;
        RECT 89.830 330.300 89.980 337.850 ;
        RECT 94.230 337.550 95.230 338.000 ;
        RECT 90.880 337.400 98.580 337.550 ;
        RECT 94.230 336.950 95.230 337.400 ;
        RECT 90.880 336.800 98.580 336.950 ;
        RECT 94.230 336.350 95.230 336.800 ;
        RECT 90.880 336.200 98.580 336.350 ;
        RECT 94.230 335.750 95.230 336.200 ;
        RECT 90.880 335.600 98.580 335.750 ;
        RECT 94.230 335.150 95.230 335.600 ;
        RECT 90.880 335.000 98.580 335.150 ;
        RECT 94.230 334.550 95.230 335.000 ;
        RECT 90.880 334.400 98.580 334.550 ;
        RECT 94.230 333.950 95.230 334.400 ;
        RECT 90.880 333.800 98.580 333.950 ;
        RECT 94.230 333.350 95.230 333.800 ;
        RECT 90.880 333.200 98.580 333.350 ;
        RECT 94.230 332.750 95.230 333.200 ;
        RECT 90.880 332.600 98.580 332.750 ;
        RECT 94.230 332.150 95.230 332.600 ;
        RECT 90.880 332.000 98.580 332.150 ;
        RECT 94.230 331.550 95.230 332.000 ;
        RECT 90.880 331.400 98.580 331.550 ;
        RECT 94.230 330.950 95.230 331.400 ;
        RECT 90.880 330.800 98.580 330.950 ;
        RECT 94.230 330.300 95.230 330.800 ;
        RECT 99.480 330.300 99.630 337.850 ;
        RECT 100.080 330.300 100.230 337.850 ;
        RECT 100.680 330.300 100.830 337.850 ;
        RECT 101.280 330.300 101.430 337.850 ;
        RECT 101.880 330.300 102.030 337.850 ;
        RECT 102.480 330.300 102.630 337.850 ;
        RECT 102.780 333.200 103.530 335.000 ;
        RECT 102.780 330.450 104.730 333.200 ;
        RECT 102.780 330.300 103.930 330.450 ;
        RECT 85.530 329.700 103.930 330.300 ;
        RECT 85.530 329.550 86.680 329.700 ;
        RECT 82.780 326.800 86.680 329.550 ;
        RECT 82.780 325.050 83.530 326.800 ;
        RECT 85.930 325.050 86.680 326.800 ;
        RECT 86.830 322.150 86.980 329.700 ;
        RECT 87.430 322.150 87.580 329.700 ;
        RECT 88.030 322.150 88.180 329.700 ;
        RECT 88.630 322.150 88.780 329.700 ;
        RECT 89.230 322.150 89.380 329.700 ;
        RECT 89.830 322.150 89.980 329.700 ;
        RECT 94.230 329.200 95.230 329.700 ;
        RECT 90.880 329.050 98.580 329.200 ;
        RECT 94.230 328.600 95.230 329.050 ;
        RECT 90.880 328.450 98.580 328.600 ;
        RECT 94.230 328.000 95.230 328.450 ;
        RECT 90.880 327.850 98.580 328.000 ;
        RECT 94.230 327.400 95.230 327.850 ;
        RECT 90.880 327.250 98.580 327.400 ;
        RECT 94.230 326.800 95.230 327.250 ;
        RECT 90.880 326.650 98.580 326.800 ;
        RECT 94.230 326.200 95.230 326.650 ;
        RECT 90.880 326.050 98.580 326.200 ;
        RECT 94.230 325.600 95.230 326.050 ;
        RECT 90.880 325.450 98.580 325.600 ;
        RECT 94.230 325.000 95.230 325.450 ;
        RECT 90.880 324.850 98.580 325.000 ;
        RECT 94.230 324.400 95.230 324.850 ;
        RECT 90.880 324.250 98.580 324.400 ;
        RECT 94.230 323.800 95.230 324.250 ;
        RECT 90.880 323.650 98.580 323.800 ;
        RECT 94.230 323.200 95.230 323.650 ;
        RECT 90.880 323.050 98.580 323.200 ;
        RECT 94.230 322.600 95.230 323.050 ;
        RECT 90.880 322.450 98.580 322.600 ;
        RECT 94.230 322.000 95.230 322.450 ;
        RECT 99.480 322.150 99.630 329.700 ;
        RECT 100.080 322.150 100.230 329.700 ;
        RECT 100.680 322.150 100.830 329.700 ;
        RECT 101.280 322.150 101.430 329.700 ;
        RECT 101.880 322.150 102.030 329.700 ;
        RECT 102.480 322.150 102.630 329.700 ;
        RECT 102.780 329.550 103.930 329.700 ;
        RECT 104.580 330.415 104.730 330.450 ;
        RECT 104.580 329.550 111.850 330.415 ;
        RECT 102.780 329.140 111.850 329.550 ;
        RECT 102.780 326.800 104.730 329.140 ;
        RECT 102.780 325.050 103.530 326.800 ;
        RECT 10.880 321.850 18.580 322.000 ;
        RECT 30.880 321.850 38.580 322.000 ;
        RECT 50.880 321.850 58.580 322.000 ;
        RECT 70.880 321.850 78.580 322.000 ;
        RECT 90.880 321.850 98.580 322.000 ;
        RECT 14.230 321.200 15.230 321.850 ;
        RECT 34.230 321.200 35.230 321.850 ;
        RECT 54.230 321.200 55.230 321.850 ;
        RECT 74.230 321.200 75.230 321.850 ;
        RECT 94.230 321.200 95.230 321.850 ;
        RECT 11.530 318.800 17.930 321.200 ;
        RECT 31.530 318.800 37.930 321.200 ;
        RECT 51.530 318.800 57.930 321.200 ;
        RECT 71.530 318.800 77.930 321.200 ;
        RECT 91.530 318.800 97.930 321.200 ;
        RECT 14.230 318.150 15.230 318.800 ;
        RECT 34.230 318.150 35.230 318.800 ;
        RECT 54.230 318.150 55.230 318.800 ;
        RECT 74.230 318.150 75.230 318.800 ;
        RECT 94.230 318.150 95.230 318.800 ;
        RECT 10.880 318.000 18.580 318.150 ;
        RECT 30.880 318.000 38.580 318.150 ;
        RECT 50.880 318.000 58.580 318.150 ;
        RECT 70.880 318.000 78.580 318.150 ;
        RECT 90.880 318.000 98.580 318.150 ;
        RECT 5.930 313.200 6.680 315.000 ;
        RECT 4.730 310.450 6.680 313.200 ;
        RECT 4.730 309.550 4.880 310.450 ;
        RECT 5.530 310.300 6.680 310.450 ;
        RECT 6.830 310.300 6.980 317.850 ;
        RECT 7.430 310.300 7.580 317.850 ;
        RECT 8.030 310.300 8.180 317.850 ;
        RECT 8.630 310.300 8.780 317.850 ;
        RECT 9.230 310.300 9.380 317.850 ;
        RECT 9.830 310.300 9.980 317.850 ;
        RECT 14.230 317.550 15.230 318.000 ;
        RECT 10.880 317.400 18.580 317.550 ;
        RECT 14.230 316.950 15.230 317.400 ;
        RECT 10.880 316.800 18.580 316.950 ;
        RECT 14.230 316.350 15.230 316.800 ;
        RECT 10.880 316.200 18.580 316.350 ;
        RECT 14.230 315.750 15.230 316.200 ;
        RECT 10.880 315.600 18.580 315.750 ;
        RECT 14.230 315.150 15.230 315.600 ;
        RECT 10.880 315.000 18.580 315.150 ;
        RECT 14.230 314.550 15.230 315.000 ;
        RECT 10.880 314.400 18.580 314.550 ;
        RECT 14.230 313.950 15.230 314.400 ;
        RECT 10.880 313.800 18.580 313.950 ;
        RECT 14.230 313.350 15.230 313.800 ;
        RECT 10.880 313.200 18.580 313.350 ;
        RECT 14.230 312.750 15.230 313.200 ;
        RECT 10.880 312.600 18.580 312.750 ;
        RECT 14.230 312.150 15.230 312.600 ;
        RECT 10.880 312.000 18.580 312.150 ;
        RECT 14.230 311.550 15.230 312.000 ;
        RECT 10.880 311.400 18.580 311.550 ;
        RECT 14.230 310.950 15.230 311.400 ;
        RECT 10.880 310.800 18.580 310.950 ;
        RECT 14.230 310.300 15.230 310.800 ;
        RECT 19.480 310.300 19.630 317.850 ;
        RECT 20.080 310.300 20.230 317.850 ;
        RECT 20.680 310.300 20.830 317.850 ;
        RECT 21.280 310.300 21.430 317.850 ;
        RECT 21.880 310.300 22.030 317.850 ;
        RECT 22.480 310.300 22.630 317.850 ;
        RECT 22.780 313.200 23.530 315.000 ;
        RECT 25.930 313.200 26.680 315.000 ;
        RECT 22.780 310.450 26.680 313.200 ;
        RECT 22.780 310.300 23.930 310.450 ;
        RECT 5.530 309.700 23.930 310.300 ;
        RECT 5.530 309.550 6.680 309.700 ;
        RECT 4.730 306.800 6.680 309.550 ;
        RECT 5.930 305.050 6.680 306.800 ;
        RECT 6.830 302.150 6.980 309.700 ;
        RECT 7.430 302.150 7.580 309.700 ;
        RECT 8.030 302.150 8.180 309.700 ;
        RECT 8.630 302.150 8.780 309.700 ;
        RECT 9.230 302.150 9.380 309.700 ;
        RECT 9.830 302.150 9.980 309.700 ;
        RECT 14.230 309.200 15.230 309.700 ;
        RECT 10.880 309.050 18.580 309.200 ;
        RECT 14.230 308.600 15.230 309.050 ;
        RECT 10.880 308.450 18.580 308.600 ;
        RECT 14.230 308.000 15.230 308.450 ;
        RECT 10.880 307.850 18.580 308.000 ;
        RECT 14.230 307.400 15.230 307.850 ;
        RECT 10.880 307.250 18.580 307.400 ;
        RECT 14.230 306.800 15.230 307.250 ;
        RECT 10.880 306.650 18.580 306.800 ;
        RECT 14.230 306.200 15.230 306.650 ;
        RECT 10.880 306.050 18.580 306.200 ;
        RECT 14.230 305.600 15.230 306.050 ;
        RECT 10.880 305.450 18.580 305.600 ;
        RECT 14.230 305.000 15.230 305.450 ;
        RECT 10.880 304.850 18.580 305.000 ;
        RECT 14.230 304.400 15.230 304.850 ;
        RECT 10.880 304.250 18.580 304.400 ;
        RECT 14.230 303.800 15.230 304.250 ;
        RECT 10.880 303.650 18.580 303.800 ;
        RECT 14.230 303.200 15.230 303.650 ;
        RECT 10.880 303.050 18.580 303.200 ;
        RECT 14.230 302.600 15.230 303.050 ;
        RECT 10.880 302.450 18.580 302.600 ;
        RECT 14.230 302.000 15.230 302.450 ;
        RECT 19.480 302.150 19.630 309.700 ;
        RECT 20.080 302.150 20.230 309.700 ;
        RECT 20.680 302.150 20.830 309.700 ;
        RECT 21.280 302.150 21.430 309.700 ;
        RECT 21.880 302.150 22.030 309.700 ;
        RECT 22.480 302.150 22.630 309.700 ;
        RECT 22.780 309.550 23.930 309.700 ;
        RECT 24.580 309.550 24.880 310.450 ;
        RECT 25.530 310.300 26.680 310.450 ;
        RECT 26.830 310.300 26.980 317.850 ;
        RECT 27.430 310.300 27.580 317.850 ;
        RECT 28.030 310.300 28.180 317.850 ;
        RECT 28.630 310.300 28.780 317.850 ;
        RECT 29.230 310.300 29.380 317.850 ;
        RECT 29.830 310.300 29.980 317.850 ;
        RECT 34.230 317.550 35.230 318.000 ;
        RECT 30.880 317.400 38.580 317.550 ;
        RECT 34.230 316.950 35.230 317.400 ;
        RECT 30.880 316.800 38.580 316.950 ;
        RECT 34.230 316.350 35.230 316.800 ;
        RECT 30.880 316.200 38.580 316.350 ;
        RECT 34.230 315.750 35.230 316.200 ;
        RECT 30.880 315.600 38.580 315.750 ;
        RECT 34.230 315.150 35.230 315.600 ;
        RECT 30.880 315.000 38.580 315.150 ;
        RECT 34.230 314.550 35.230 315.000 ;
        RECT 30.880 314.400 38.580 314.550 ;
        RECT 34.230 313.950 35.230 314.400 ;
        RECT 30.880 313.800 38.580 313.950 ;
        RECT 34.230 313.350 35.230 313.800 ;
        RECT 30.880 313.200 38.580 313.350 ;
        RECT 34.230 312.750 35.230 313.200 ;
        RECT 30.880 312.600 38.580 312.750 ;
        RECT 34.230 312.150 35.230 312.600 ;
        RECT 30.880 312.000 38.580 312.150 ;
        RECT 34.230 311.550 35.230 312.000 ;
        RECT 30.880 311.400 38.580 311.550 ;
        RECT 34.230 310.950 35.230 311.400 ;
        RECT 30.880 310.800 38.580 310.950 ;
        RECT 34.230 310.300 35.230 310.800 ;
        RECT 39.480 310.300 39.630 317.850 ;
        RECT 40.080 310.300 40.230 317.850 ;
        RECT 40.680 310.300 40.830 317.850 ;
        RECT 41.280 310.300 41.430 317.850 ;
        RECT 41.880 310.300 42.030 317.850 ;
        RECT 42.480 310.300 42.630 317.850 ;
        RECT 42.780 313.200 43.530 315.000 ;
        RECT 45.930 313.200 46.680 315.000 ;
        RECT 42.780 310.450 46.680 313.200 ;
        RECT 42.780 310.300 43.930 310.450 ;
        RECT 25.530 309.700 43.930 310.300 ;
        RECT 25.530 309.550 26.680 309.700 ;
        RECT 22.780 306.800 26.680 309.550 ;
        RECT 22.780 305.050 23.530 306.800 ;
        RECT 25.930 305.050 26.680 306.800 ;
        RECT 26.830 302.150 26.980 309.700 ;
        RECT 27.430 302.150 27.580 309.700 ;
        RECT 28.030 302.150 28.180 309.700 ;
        RECT 28.630 302.150 28.780 309.700 ;
        RECT 29.230 302.150 29.380 309.700 ;
        RECT 29.830 302.150 29.980 309.700 ;
        RECT 34.230 309.200 35.230 309.700 ;
        RECT 30.880 309.050 38.580 309.200 ;
        RECT 34.230 308.600 35.230 309.050 ;
        RECT 30.880 308.450 38.580 308.600 ;
        RECT 34.230 308.000 35.230 308.450 ;
        RECT 30.880 307.850 38.580 308.000 ;
        RECT 34.230 307.400 35.230 307.850 ;
        RECT 30.880 307.250 38.580 307.400 ;
        RECT 34.230 306.800 35.230 307.250 ;
        RECT 30.880 306.650 38.580 306.800 ;
        RECT 34.230 306.200 35.230 306.650 ;
        RECT 30.880 306.050 38.580 306.200 ;
        RECT 34.230 305.600 35.230 306.050 ;
        RECT 30.880 305.450 38.580 305.600 ;
        RECT 34.230 305.000 35.230 305.450 ;
        RECT 30.880 304.850 38.580 305.000 ;
        RECT 34.230 304.400 35.230 304.850 ;
        RECT 30.880 304.250 38.580 304.400 ;
        RECT 34.230 303.800 35.230 304.250 ;
        RECT 30.880 303.650 38.580 303.800 ;
        RECT 34.230 303.200 35.230 303.650 ;
        RECT 30.880 303.050 38.580 303.200 ;
        RECT 34.230 302.600 35.230 303.050 ;
        RECT 30.880 302.450 38.580 302.600 ;
        RECT 34.230 302.000 35.230 302.450 ;
        RECT 39.480 302.150 39.630 309.700 ;
        RECT 40.080 302.150 40.230 309.700 ;
        RECT 40.680 302.150 40.830 309.700 ;
        RECT 41.280 302.150 41.430 309.700 ;
        RECT 41.880 302.150 42.030 309.700 ;
        RECT 42.480 302.150 42.630 309.700 ;
        RECT 42.780 309.550 43.930 309.700 ;
        RECT 44.580 309.550 44.880 310.450 ;
        RECT 45.530 310.300 46.680 310.450 ;
        RECT 46.830 310.300 46.980 317.850 ;
        RECT 47.430 310.300 47.580 317.850 ;
        RECT 48.030 310.300 48.180 317.850 ;
        RECT 48.630 310.300 48.780 317.850 ;
        RECT 49.230 310.300 49.380 317.850 ;
        RECT 49.830 310.300 49.980 317.850 ;
        RECT 54.230 317.550 55.230 318.000 ;
        RECT 50.880 317.400 58.580 317.550 ;
        RECT 54.230 316.950 55.230 317.400 ;
        RECT 50.880 316.800 58.580 316.950 ;
        RECT 54.230 316.350 55.230 316.800 ;
        RECT 50.880 316.200 58.580 316.350 ;
        RECT 54.230 315.750 55.230 316.200 ;
        RECT 50.880 315.600 58.580 315.750 ;
        RECT 54.230 315.150 55.230 315.600 ;
        RECT 50.880 315.000 58.580 315.150 ;
        RECT 54.230 314.550 55.230 315.000 ;
        RECT 50.880 314.400 58.580 314.550 ;
        RECT 54.230 313.950 55.230 314.400 ;
        RECT 50.880 313.800 58.580 313.950 ;
        RECT 54.230 313.350 55.230 313.800 ;
        RECT 50.880 313.200 58.580 313.350 ;
        RECT 54.230 312.750 55.230 313.200 ;
        RECT 50.880 312.600 58.580 312.750 ;
        RECT 54.230 312.150 55.230 312.600 ;
        RECT 50.880 312.000 58.580 312.150 ;
        RECT 54.230 311.550 55.230 312.000 ;
        RECT 50.880 311.400 58.580 311.550 ;
        RECT 54.230 310.950 55.230 311.400 ;
        RECT 50.880 310.800 58.580 310.950 ;
        RECT 54.230 310.300 55.230 310.800 ;
        RECT 59.480 310.300 59.630 317.850 ;
        RECT 60.080 310.300 60.230 317.850 ;
        RECT 60.680 310.300 60.830 317.850 ;
        RECT 61.280 310.300 61.430 317.850 ;
        RECT 61.880 310.300 62.030 317.850 ;
        RECT 62.480 310.300 62.630 317.850 ;
        RECT 62.780 313.200 63.530 315.000 ;
        RECT 65.930 313.200 66.680 315.000 ;
        RECT 62.780 310.450 66.680 313.200 ;
        RECT 62.780 310.300 63.930 310.450 ;
        RECT 45.530 309.700 63.930 310.300 ;
        RECT 45.530 309.550 46.680 309.700 ;
        RECT 42.780 306.800 46.680 309.550 ;
        RECT 42.780 305.050 43.530 306.800 ;
        RECT 45.930 305.050 46.680 306.800 ;
        RECT 46.830 302.150 46.980 309.700 ;
        RECT 47.430 302.150 47.580 309.700 ;
        RECT 48.030 302.150 48.180 309.700 ;
        RECT 48.630 302.150 48.780 309.700 ;
        RECT 49.230 302.150 49.380 309.700 ;
        RECT 49.830 302.150 49.980 309.700 ;
        RECT 54.230 309.200 55.230 309.700 ;
        RECT 50.880 309.050 58.580 309.200 ;
        RECT 54.230 308.600 55.230 309.050 ;
        RECT 50.880 308.450 58.580 308.600 ;
        RECT 54.230 308.000 55.230 308.450 ;
        RECT 50.880 307.850 58.580 308.000 ;
        RECT 54.230 307.400 55.230 307.850 ;
        RECT 50.880 307.250 58.580 307.400 ;
        RECT 54.230 306.800 55.230 307.250 ;
        RECT 50.880 306.650 58.580 306.800 ;
        RECT 54.230 306.200 55.230 306.650 ;
        RECT 50.880 306.050 58.580 306.200 ;
        RECT 54.230 305.600 55.230 306.050 ;
        RECT 50.880 305.450 58.580 305.600 ;
        RECT 54.230 305.000 55.230 305.450 ;
        RECT 50.880 304.850 58.580 305.000 ;
        RECT 54.230 304.400 55.230 304.850 ;
        RECT 50.880 304.250 58.580 304.400 ;
        RECT 54.230 303.800 55.230 304.250 ;
        RECT 50.880 303.650 58.580 303.800 ;
        RECT 54.230 303.200 55.230 303.650 ;
        RECT 50.880 303.050 58.580 303.200 ;
        RECT 54.230 302.600 55.230 303.050 ;
        RECT 50.880 302.450 58.580 302.600 ;
        RECT 54.230 302.000 55.230 302.450 ;
        RECT 59.480 302.150 59.630 309.700 ;
        RECT 60.080 302.150 60.230 309.700 ;
        RECT 60.680 302.150 60.830 309.700 ;
        RECT 61.280 302.150 61.430 309.700 ;
        RECT 61.880 302.150 62.030 309.700 ;
        RECT 62.480 302.150 62.630 309.700 ;
        RECT 62.780 309.550 63.930 309.700 ;
        RECT 64.580 309.550 64.880 310.450 ;
        RECT 65.530 310.300 66.680 310.450 ;
        RECT 66.830 310.300 66.980 317.850 ;
        RECT 67.430 310.300 67.580 317.850 ;
        RECT 68.030 310.300 68.180 317.850 ;
        RECT 68.630 310.300 68.780 317.850 ;
        RECT 69.230 310.300 69.380 317.850 ;
        RECT 69.830 310.300 69.980 317.850 ;
        RECT 74.230 317.550 75.230 318.000 ;
        RECT 70.880 317.400 78.580 317.550 ;
        RECT 74.230 316.950 75.230 317.400 ;
        RECT 70.880 316.800 78.580 316.950 ;
        RECT 74.230 316.350 75.230 316.800 ;
        RECT 70.880 316.200 78.580 316.350 ;
        RECT 74.230 315.750 75.230 316.200 ;
        RECT 70.880 315.600 78.580 315.750 ;
        RECT 74.230 315.150 75.230 315.600 ;
        RECT 70.880 315.000 78.580 315.150 ;
        RECT 74.230 314.550 75.230 315.000 ;
        RECT 70.880 314.400 78.580 314.550 ;
        RECT 74.230 313.950 75.230 314.400 ;
        RECT 70.880 313.800 78.580 313.950 ;
        RECT 74.230 313.350 75.230 313.800 ;
        RECT 70.880 313.200 78.580 313.350 ;
        RECT 74.230 312.750 75.230 313.200 ;
        RECT 70.880 312.600 78.580 312.750 ;
        RECT 74.230 312.150 75.230 312.600 ;
        RECT 70.880 312.000 78.580 312.150 ;
        RECT 74.230 311.550 75.230 312.000 ;
        RECT 70.880 311.400 78.580 311.550 ;
        RECT 74.230 310.950 75.230 311.400 ;
        RECT 70.880 310.800 78.580 310.950 ;
        RECT 74.230 310.300 75.230 310.800 ;
        RECT 79.480 310.300 79.630 317.850 ;
        RECT 80.080 310.300 80.230 317.850 ;
        RECT 80.680 310.300 80.830 317.850 ;
        RECT 81.280 310.300 81.430 317.850 ;
        RECT 81.880 310.300 82.030 317.850 ;
        RECT 82.480 310.300 82.630 317.850 ;
        RECT 82.780 313.200 83.530 315.000 ;
        RECT 85.930 313.200 86.680 315.000 ;
        RECT 82.780 310.450 86.680 313.200 ;
        RECT 82.780 310.300 83.930 310.450 ;
        RECT 65.530 309.700 83.930 310.300 ;
        RECT 65.530 309.550 66.680 309.700 ;
        RECT 62.780 306.800 66.680 309.550 ;
        RECT 62.780 305.050 63.530 306.800 ;
        RECT 65.930 305.050 66.680 306.800 ;
        RECT 66.830 302.150 66.980 309.700 ;
        RECT 67.430 302.150 67.580 309.700 ;
        RECT 68.030 302.150 68.180 309.700 ;
        RECT 68.630 302.150 68.780 309.700 ;
        RECT 69.230 302.150 69.380 309.700 ;
        RECT 69.830 302.150 69.980 309.700 ;
        RECT 74.230 309.200 75.230 309.700 ;
        RECT 70.880 309.050 78.580 309.200 ;
        RECT 74.230 308.600 75.230 309.050 ;
        RECT 70.880 308.450 78.580 308.600 ;
        RECT 74.230 308.000 75.230 308.450 ;
        RECT 70.880 307.850 78.580 308.000 ;
        RECT 74.230 307.400 75.230 307.850 ;
        RECT 70.880 307.250 78.580 307.400 ;
        RECT 74.230 306.800 75.230 307.250 ;
        RECT 70.880 306.650 78.580 306.800 ;
        RECT 74.230 306.200 75.230 306.650 ;
        RECT 70.880 306.050 78.580 306.200 ;
        RECT 74.230 305.600 75.230 306.050 ;
        RECT 70.880 305.450 78.580 305.600 ;
        RECT 74.230 305.000 75.230 305.450 ;
        RECT 70.880 304.850 78.580 305.000 ;
        RECT 74.230 304.400 75.230 304.850 ;
        RECT 70.880 304.250 78.580 304.400 ;
        RECT 74.230 303.800 75.230 304.250 ;
        RECT 70.880 303.650 78.580 303.800 ;
        RECT 74.230 303.200 75.230 303.650 ;
        RECT 70.880 303.050 78.580 303.200 ;
        RECT 74.230 302.600 75.230 303.050 ;
        RECT 70.880 302.450 78.580 302.600 ;
        RECT 74.230 302.000 75.230 302.450 ;
        RECT 79.480 302.150 79.630 309.700 ;
        RECT 80.080 302.150 80.230 309.700 ;
        RECT 80.680 302.150 80.830 309.700 ;
        RECT 81.280 302.150 81.430 309.700 ;
        RECT 81.880 302.150 82.030 309.700 ;
        RECT 82.480 302.150 82.630 309.700 ;
        RECT 82.780 309.550 83.930 309.700 ;
        RECT 84.580 309.550 84.880 310.450 ;
        RECT 85.530 310.300 86.680 310.450 ;
        RECT 86.830 310.300 86.980 317.850 ;
        RECT 87.430 310.300 87.580 317.850 ;
        RECT 88.030 310.300 88.180 317.850 ;
        RECT 88.630 310.300 88.780 317.850 ;
        RECT 89.230 310.300 89.380 317.850 ;
        RECT 89.830 310.300 89.980 317.850 ;
        RECT 94.230 317.550 95.230 318.000 ;
        RECT 90.880 317.400 98.580 317.550 ;
        RECT 94.230 316.950 95.230 317.400 ;
        RECT 90.880 316.800 98.580 316.950 ;
        RECT 94.230 316.350 95.230 316.800 ;
        RECT 90.880 316.200 98.580 316.350 ;
        RECT 94.230 315.750 95.230 316.200 ;
        RECT 90.880 315.600 98.580 315.750 ;
        RECT 94.230 315.150 95.230 315.600 ;
        RECT 90.880 315.000 98.580 315.150 ;
        RECT 94.230 314.550 95.230 315.000 ;
        RECT 90.880 314.400 98.580 314.550 ;
        RECT 94.230 313.950 95.230 314.400 ;
        RECT 90.880 313.800 98.580 313.950 ;
        RECT 94.230 313.350 95.230 313.800 ;
        RECT 90.880 313.200 98.580 313.350 ;
        RECT 94.230 312.750 95.230 313.200 ;
        RECT 90.880 312.600 98.580 312.750 ;
        RECT 94.230 312.150 95.230 312.600 ;
        RECT 90.880 312.000 98.580 312.150 ;
        RECT 94.230 311.550 95.230 312.000 ;
        RECT 90.880 311.400 98.580 311.550 ;
        RECT 94.230 310.950 95.230 311.400 ;
        RECT 90.880 310.800 98.580 310.950 ;
        RECT 94.230 310.300 95.230 310.800 ;
        RECT 99.480 310.300 99.630 317.850 ;
        RECT 100.080 310.300 100.230 317.850 ;
        RECT 100.680 310.300 100.830 317.850 ;
        RECT 101.280 310.300 101.430 317.850 ;
        RECT 101.880 310.300 102.030 317.850 ;
        RECT 102.480 310.300 102.630 317.850 ;
        RECT 102.780 313.200 103.530 315.000 ;
        RECT 102.780 310.450 104.730 313.200 ;
        RECT 102.780 310.300 103.930 310.450 ;
        RECT 85.530 309.700 103.930 310.300 ;
        RECT 85.530 309.550 86.680 309.700 ;
        RECT 82.780 306.800 86.680 309.550 ;
        RECT 82.780 305.050 83.530 306.800 ;
        RECT 85.930 305.050 86.680 306.800 ;
        RECT 86.830 302.150 86.980 309.700 ;
        RECT 87.430 302.150 87.580 309.700 ;
        RECT 88.030 302.150 88.180 309.700 ;
        RECT 88.630 302.150 88.780 309.700 ;
        RECT 89.230 302.150 89.380 309.700 ;
        RECT 89.830 302.150 89.980 309.700 ;
        RECT 94.230 309.200 95.230 309.700 ;
        RECT 90.880 309.050 98.580 309.200 ;
        RECT 94.230 308.600 95.230 309.050 ;
        RECT 90.880 308.450 98.580 308.600 ;
        RECT 94.230 308.000 95.230 308.450 ;
        RECT 90.880 307.850 98.580 308.000 ;
        RECT 94.230 307.400 95.230 307.850 ;
        RECT 90.880 307.250 98.580 307.400 ;
        RECT 94.230 306.800 95.230 307.250 ;
        RECT 90.880 306.650 98.580 306.800 ;
        RECT 94.230 306.200 95.230 306.650 ;
        RECT 90.880 306.050 98.580 306.200 ;
        RECT 94.230 305.600 95.230 306.050 ;
        RECT 90.880 305.450 98.580 305.600 ;
        RECT 94.230 305.000 95.230 305.450 ;
        RECT 90.880 304.850 98.580 305.000 ;
        RECT 94.230 304.400 95.230 304.850 ;
        RECT 90.880 304.250 98.580 304.400 ;
        RECT 94.230 303.800 95.230 304.250 ;
        RECT 90.880 303.650 98.580 303.800 ;
        RECT 94.230 303.200 95.230 303.650 ;
        RECT 90.880 303.050 98.580 303.200 ;
        RECT 94.230 302.600 95.230 303.050 ;
        RECT 90.880 302.450 98.580 302.600 ;
        RECT 94.230 302.000 95.230 302.450 ;
        RECT 99.480 302.150 99.630 309.700 ;
        RECT 100.080 302.150 100.230 309.700 ;
        RECT 100.680 302.150 100.830 309.700 ;
        RECT 101.280 302.150 101.430 309.700 ;
        RECT 101.880 302.150 102.030 309.700 ;
        RECT 102.480 302.150 102.630 309.700 ;
        RECT 102.780 309.550 103.930 309.700 ;
        RECT 104.580 310.410 104.730 310.450 ;
        RECT 104.580 309.550 111.850 310.410 ;
        RECT 102.780 309.135 111.850 309.550 ;
        RECT 102.780 306.800 104.730 309.135 ;
        RECT 102.780 305.050 103.530 306.800 ;
        RECT 10.880 301.850 18.580 302.000 ;
        RECT 30.880 301.850 38.580 302.000 ;
        RECT 50.880 301.850 58.580 302.000 ;
        RECT 70.880 301.850 78.580 302.000 ;
        RECT 90.880 301.850 98.580 302.000 ;
        RECT 14.230 301.200 15.230 301.850 ;
        RECT 34.230 301.200 35.230 301.850 ;
        RECT 54.230 301.200 55.230 301.850 ;
        RECT 74.230 301.200 75.230 301.850 ;
        RECT 94.230 301.200 95.230 301.850 ;
        RECT 11.530 298.800 17.930 301.200 ;
        RECT 31.530 298.800 37.930 301.200 ;
        RECT 51.530 298.800 57.930 301.200 ;
        RECT 71.530 298.800 77.930 301.200 ;
        RECT 91.530 298.800 97.930 301.200 ;
        RECT 14.230 298.150 15.230 298.800 ;
        RECT 34.230 298.150 35.230 298.800 ;
        RECT 54.230 298.150 55.230 298.800 ;
        RECT 74.230 298.150 75.230 298.800 ;
        RECT 94.230 298.150 95.230 298.800 ;
        RECT 10.880 298.000 18.580 298.150 ;
        RECT 30.880 298.000 38.580 298.150 ;
        RECT 50.880 298.000 58.580 298.150 ;
        RECT 70.880 298.000 78.580 298.150 ;
        RECT 90.880 298.000 98.580 298.150 ;
        RECT 5.930 293.200 6.680 295.000 ;
        RECT 4.730 290.450 6.680 293.200 ;
        RECT 4.730 289.550 4.880 290.450 ;
        RECT 5.530 290.300 6.680 290.450 ;
        RECT 6.830 290.300 6.980 297.850 ;
        RECT 7.430 290.300 7.580 297.850 ;
        RECT 8.030 290.300 8.180 297.850 ;
        RECT 8.630 290.300 8.780 297.850 ;
        RECT 9.230 290.300 9.380 297.850 ;
        RECT 9.830 290.300 9.980 297.850 ;
        RECT 14.230 297.550 15.230 298.000 ;
        RECT 10.880 297.400 18.580 297.550 ;
        RECT 14.230 296.950 15.230 297.400 ;
        RECT 10.880 296.800 18.580 296.950 ;
        RECT 14.230 296.350 15.230 296.800 ;
        RECT 10.880 296.200 18.580 296.350 ;
        RECT 14.230 295.750 15.230 296.200 ;
        RECT 10.880 295.600 18.580 295.750 ;
        RECT 14.230 295.150 15.230 295.600 ;
        RECT 10.880 295.000 18.580 295.150 ;
        RECT 14.230 294.550 15.230 295.000 ;
        RECT 10.880 294.400 18.580 294.550 ;
        RECT 14.230 293.950 15.230 294.400 ;
        RECT 10.880 293.800 18.580 293.950 ;
        RECT 14.230 293.350 15.230 293.800 ;
        RECT 10.880 293.200 18.580 293.350 ;
        RECT 14.230 292.750 15.230 293.200 ;
        RECT 10.880 292.600 18.580 292.750 ;
        RECT 14.230 292.150 15.230 292.600 ;
        RECT 10.880 292.000 18.580 292.150 ;
        RECT 14.230 291.550 15.230 292.000 ;
        RECT 10.880 291.400 18.580 291.550 ;
        RECT 14.230 290.950 15.230 291.400 ;
        RECT 10.880 290.800 18.580 290.950 ;
        RECT 14.230 290.300 15.230 290.800 ;
        RECT 19.480 290.300 19.630 297.850 ;
        RECT 20.080 290.300 20.230 297.850 ;
        RECT 20.680 290.300 20.830 297.850 ;
        RECT 21.280 290.300 21.430 297.850 ;
        RECT 21.880 290.300 22.030 297.850 ;
        RECT 22.480 290.300 22.630 297.850 ;
        RECT 22.780 293.200 23.530 295.000 ;
        RECT 25.930 293.200 26.680 295.000 ;
        RECT 22.780 290.450 26.680 293.200 ;
        RECT 22.780 290.300 23.930 290.450 ;
        RECT 5.530 289.700 23.930 290.300 ;
        RECT 5.530 289.550 6.680 289.700 ;
        RECT 4.730 286.800 6.680 289.550 ;
        RECT 5.930 285.050 6.680 286.800 ;
        RECT 6.830 282.150 6.980 289.700 ;
        RECT 7.430 282.150 7.580 289.700 ;
        RECT 8.030 282.150 8.180 289.700 ;
        RECT 8.630 282.150 8.780 289.700 ;
        RECT 9.230 282.150 9.380 289.700 ;
        RECT 9.830 282.150 9.980 289.700 ;
        RECT 14.230 289.200 15.230 289.700 ;
        RECT 10.880 289.050 18.580 289.200 ;
        RECT 14.230 288.600 15.230 289.050 ;
        RECT 10.880 288.450 18.580 288.600 ;
        RECT 14.230 288.000 15.230 288.450 ;
        RECT 10.880 287.850 18.580 288.000 ;
        RECT 14.230 287.400 15.230 287.850 ;
        RECT 10.880 287.250 18.580 287.400 ;
        RECT 14.230 286.800 15.230 287.250 ;
        RECT 10.880 286.650 18.580 286.800 ;
        RECT 14.230 286.200 15.230 286.650 ;
        RECT 10.880 286.050 18.580 286.200 ;
        RECT 14.230 285.600 15.230 286.050 ;
        RECT 10.880 285.450 18.580 285.600 ;
        RECT 14.230 285.000 15.230 285.450 ;
        RECT 10.880 284.850 18.580 285.000 ;
        RECT 14.230 284.400 15.230 284.850 ;
        RECT 10.880 284.250 18.580 284.400 ;
        RECT 14.230 283.800 15.230 284.250 ;
        RECT 10.880 283.650 18.580 283.800 ;
        RECT 14.230 283.200 15.230 283.650 ;
        RECT 10.880 283.050 18.580 283.200 ;
        RECT 14.230 282.600 15.230 283.050 ;
        RECT 10.880 282.450 18.580 282.600 ;
        RECT 14.230 282.000 15.230 282.450 ;
        RECT 19.480 282.150 19.630 289.700 ;
        RECT 20.080 282.150 20.230 289.700 ;
        RECT 20.680 282.150 20.830 289.700 ;
        RECT 21.280 282.150 21.430 289.700 ;
        RECT 21.880 282.150 22.030 289.700 ;
        RECT 22.480 282.150 22.630 289.700 ;
        RECT 22.780 289.550 23.930 289.700 ;
        RECT 24.580 289.550 24.880 290.450 ;
        RECT 25.530 290.300 26.680 290.450 ;
        RECT 26.830 290.300 26.980 297.850 ;
        RECT 27.430 290.300 27.580 297.850 ;
        RECT 28.030 290.300 28.180 297.850 ;
        RECT 28.630 290.300 28.780 297.850 ;
        RECT 29.230 290.300 29.380 297.850 ;
        RECT 29.830 290.300 29.980 297.850 ;
        RECT 34.230 297.550 35.230 298.000 ;
        RECT 30.880 297.400 38.580 297.550 ;
        RECT 34.230 296.950 35.230 297.400 ;
        RECT 30.880 296.800 38.580 296.950 ;
        RECT 34.230 296.350 35.230 296.800 ;
        RECT 30.880 296.200 38.580 296.350 ;
        RECT 34.230 295.750 35.230 296.200 ;
        RECT 30.880 295.600 38.580 295.750 ;
        RECT 34.230 295.150 35.230 295.600 ;
        RECT 30.880 295.000 38.580 295.150 ;
        RECT 34.230 294.550 35.230 295.000 ;
        RECT 30.880 294.400 38.580 294.550 ;
        RECT 34.230 293.950 35.230 294.400 ;
        RECT 30.880 293.800 38.580 293.950 ;
        RECT 34.230 293.350 35.230 293.800 ;
        RECT 30.880 293.200 38.580 293.350 ;
        RECT 34.230 292.750 35.230 293.200 ;
        RECT 30.880 292.600 38.580 292.750 ;
        RECT 34.230 292.150 35.230 292.600 ;
        RECT 30.880 292.000 38.580 292.150 ;
        RECT 34.230 291.550 35.230 292.000 ;
        RECT 30.880 291.400 38.580 291.550 ;
        RECT 34.230 290.950 35.230 291.400 ;
        RECT 30.880 290.800 38.580 290.950 ;
        RECT 34.230 290.300 35.230 290.800 ;
        RECT 39.480 290.300 39.630 297.850 ;
        RECT 40.080 290.300 40.230 297.850 ;
        RECT 40.680 290.300 40.830 297.850 ;
        RECT 41.280 290.300 41.430 297.850 ;
        RECT 41.880 290.300 42.030 297.850 ;
        RECT 42.480 290.300 42.630 297.850 ;
        RECT 42.780 293.200 43.530 295.000 ;
        RECT 45.930 293.200 46.680 295.000 ;
        RECT 42.780 290.450 46.680 293.200 ;
        RECT 42.780 290.300 43.930 290.450 ;
        RECT 25.530 289.700 43.930 290.300 ;
        RECT 25.530 289.550 26.680 289.700 ;
        RECT 22.780 286.800 26.680 289.550 ;
        RECT 22.780 285.050 23.530 286.800 ;
        RECT 25.930 285.050 26.680 286.800 ;
        RECT 26.830 282.150 26.980 289.700 ;
        RECT 27.430 282.150 27.580 289.700 ;
        RECT 28.030 282.150 28.180 289.700 ;
        RECT 28.630 282.150 28.780 289.700 ;
        RECT 29.230 282.150 29.380 289.700 ;
        RECT 29.830 282.150 29.980 289.700 ;
        RECT 34.230 289.200 35.230 289.700 ;
        RECT 30.880 289.050 38.580 289.200 ;
        RECT 34.230 288.600 35.230 289.050 ;
        RECT 30.880 288.450 38.580 288.600 ;
        RECT 34.230 288.000 35.230 288.450 ;
        RECT 30.880 287.850 38.580 288.000 ;
        RECT 34.230 287.400 35.230 287.850 ;
        RECT 30.880 287.250 38.580 287.400 ;
        RECT 34.230 286.800 35.230 287.250 ;
        RECT 30.880 286.650 38.580 286.800 ;
        RECT 34.230 286.200 35.230 286.650 ;
        RECT 30.880 286.050 38.580 286.200 ;
        RECT 34.230 285.600 35.230 286.050 ;
        RECT 30.880 285.450 38.580 285.600 ;
        RECT 34.230 285.000 35.230 285.450 ;
        RECT 30.880 284.850 38.580 285.000 ;
        RECT 34.230 284.400 35.230 284.850 ;
        RECT 30.880 284.250 38.580 284.400 ;
        RECT 34.230 283.800 35.230 284.250 ;
        RECT 30.880 283.650 38.580 283.800 ;
        RECT 34.230 283.200 35.230 283.650 ;
        RECT 30.880 283.050 38.580 283.200 ;
        RECT 34.230 282.600 35.230 283.050 ;
        RECT 30.880 282.450 38.580 282.600 ;
        RECT 34.230 282.000 35.230 282.450 ;
        RECT 39.480 282.150 39.630 289.700 ;
        RECT 40.080 282.150 40.230 289.700 ;
        RECT 40.680 282.150 40.830 289.700 ;
        RECT 41.280 282.150 41.430 289.700 ;
        RECT 41.880 282.150 42.030 289.700 ;
        RECT 42.480 282.150 42.630 289.700 ;
        RECT 42.780 289.550 43.930 289.700 ;
        RECT 44.580 289.550 44.880 290.450 ;
        RECT 45.530 290.300 46.680 290.450 ;
        RECT 46.830 290.300 46.980 297.850 ;
        RECT 47.430 290.300 47.580 297.850 ;
        RECT 48.030 290.300 48.180 297.850 ;
        RECT 48.630 290.300 48.780 297.850 ;
        RECT 49.230 290.300 49.380 297.850 ;
        RECT 49.830 290.300 49.980 297.850 ;
        RECT 54.230 297.550 55.230 298.000 ;
        RECT 50.880 297.400 58.580 297.550 ;
        RECT 54.230 296.950 55.230 297.400 ;
        RECT 50.880 296.800 58.580 296.950 ;
        RECT 54.230 296.350 55.230 296.800 ;
        RECT 50.880 296.200 58.580 296.350 ;
        RECT 54.230 295.750 55.230 296.200 ;
        RECT 50.880 295.600 58.580 295.750 ;
        RECT 54.230 295.150 55.230 295.600 ;
        RECT 50.880 295.000 58.580 295.150 ;
        RECT 54.230 294.550 55.230 295.000 ;
        RECT 50.880 294.400 58.580 294.550 ;
        RECT 54.230 293.950 55.230 294.400 ;
        RECT 50.880 293.800 58.580 293.950 ;
        RECT 54.230 293.350 55.230 293.800 ;
        RECT 50.880 293.200 58.580 293.350 ;
        RECT 54.230 292.750 55.230 293.200 ;
        RECT 50.880 292.600 58.580 292.750 ;
        RECT 54.230 292.150 55.230 292.600 ;
        RECT 50.880 292.000 58.580 292.150 ;
        RECT 54.230 291.550 55.230 292.000 ;
        RECT 50.880 291.400 58.580 291.550 ;
        RECT 54.230 290.950 55.230 291.400 ;
        RECT 50.880 290.800 58.580 290.950 ;
        RECT 54.230 290.300 55.230 290.800 ;
        RECT 59.480 290.300 59.630 297.850 ;
        RECT 60.080 290.300 60.230 297.850 ;
        RECT 60.680 290.300 60.830 297.850 ;
        RECT 61.280 290.300 61.430 297.850 ;
        RECT 61.880 290.300 62.030 297.850 ;
        RECT 62.480 290.300 62.630 297.850 ;
        RECT 62.780 293.200 63.530 295.000 ;
        RECT 65.930 293.200 66.680 295.000 ;
        RECT 62.780 290.450 66.680 293.200 ;
        RECT 62.780 290.300 63.930 290.450 ;
        RECT 45.530 289.700 63.930 290.300 ;
        RECT 45.530 289.550 46.680 289.700 ;
        RECT 42.780 286.800 46.680 289.550 ;
        RECT 42.780 285.050 43.530 286.800 ;
        RECT 45.930 285.050 46.680 286.800 ;
        RECT 46.830 282.150 46.980 289.700 ;
        RECT 47.430 282.150 47.580 289.700 ;
        RECT 48.030 282.150 48.180 289.700 ;
        RECT 48.630 282.150 48.780 289.700 ;
        RECT 49.230 282.150 49.380 289.700 ;
        RECT 49.830 282.150 49.980 289.700 ;
        RECT 54.230 289.200 55.230 289.700 ;
        RECT 50.880 289.050 58.580 289.200 ;
        RECT 54.230 288.600 55.230 289.050 ;
        RECT 50.880 288.450 58.580 288.600 ;
        RECT 54.230 288.000 55.230 288.450 ;
        RECT 50.880 287.850 58.580 288.000 ;
        RECT 54.230 287.400 55.230 287.850 ;
        RECT 50.880 287.250 58.580 287.400 ;
        RECT 54.230 286.800 55.230 287.250 ;
        RECT 50.880 286.650 58.580 286.800 ;
        RECT 54.230 286.200 55.230 286.650 ;
        RECT 50.880 286.050 58.580 286.200 ;
        RECT 54.230 285.600 55.230 286.050 ;
        RECT 50.880 285.450 58.580 285.600 ;
        RECT 54.230 285.000 55.230 285.450 ;
        RECT 50.880 284.850 58.580 285.000 ;
        RECT 54.230 284.400 55.230 284.850 ;
        RECT 50.880 284.250 58.580 284.400 ;
        RECT 54.230 283.800 55.230 284.250 ;
        RECT 50.880 283.650 58.580 283.800 ;
        RECT 54.230 283.200 55.230 283.650 ;
        RECT 50.880 283.050 58.580 283.200 ;
        RECT 54.230 282.600 55.230 283.050 ;
        RECT 50.880 282.450 58.580 282.600 ;
        RECT 54.230 282.000 55.230 282.450 ;
        RECT 59.480 282.150 59.630 289.700 ;
        RECT 60.080 282.150 60.230 289.700 ;
        RECT 60.680 282.150 60.830 289.700 ;
        RECT 61.280 282.150 61.430 289.700 ;
        RECT 61.880 282.150 62.030 289.700 ;
        RECT 62.480 282.150 62.630 289.700 ;
        RECT 62.780 289.550 63.930 289.700 ;
        RECT 64.580 289.550 64.880 290.450 ;
        RECT 65.530 290.300 66.680 290.450 ;
        RECT 66.830 290.300 66.980 297.850 ;
        RECT 67.430 290.300 67.580 297.850 ;
        RECT 68.030 290.300 68.180 297.850 ;
        RECT 68.630 290.300 68.780 297.850 ;
        RECT 69.230 290.300 69.380 297.850 ;
        RECT 69.830 290.300 69.980 297.850 ;
        RECT 74.230 297.550 75.230 298.000 ;
        RECT 70.880 297.400 78.580 297.550 ;
        RECT 74.230 296.950 75.230 297.400 ;
        RECT 70.880 296.800 78.580 296.950 ;
        RECT 74.230 296.350 75.230 296.800 ;
        RECT 70.880 296.200 78.580 296.350 ;
        RECT 74.230 295.750 75.230 296.200 ;
        RECT 70.880 295.600 78.580 295.750 ;
        RECT 74.230 295.150 75.230 295.600 ;
        RECT 70.880 295.000 78.580 295.150 ;
        RECT 74.230 294.550 75.230 295.000 ;
        RECT 70.880 294.400 78.580 294.550 ;
        RECT 74.230 293.950 75.230 294.400 ;
        RECT 70.880 293.800 78.580 293.950 ;
        RECT 74.230 293.350 75.230 293.800 ;
        RECT 70.880 293.200 78.580 293.350 ;
        RECT 74.230 292.750 75.230 293.200 ;
        RECT 70.880 292.600 78.580 292.750 ;
        RECT 74.230 292.150 75.230 292.600 ;
        RECT 70.880 292.000 78.580 292.150 ;
        RECT 74.230 291.550 75.230 292.000 ;
        RECT 70.880 291.400 78.580 291.550 ;
        RECT 74.230 290.950 75.230 291.400 ;
        RECT 70.880 290.800 78.580 290.950 ;
        RECT 74.230 290.300 75.230 290.800 ;
        RECT 79.480 290.300 79.630 297.850 ;
        RECT 80.080 290.300 80.230 297.850 ;
        RECT 80.680 290.300 80.830 297.850 ;
        RECT 81.280 290.300 81.430 297.850 ;
        RECT 81.880 290.300 82.030 297.850 ;
        RECT 82.480 290.300 82.630 297.850 ;
        RECT 82.780 293.200 83.530 295.000 ;
        RECT 85.930 293.200 86.680 295.000 ;
        RECT 82.780 290.450 86.680 293.200 ;
        RECT 82.780 290.300 83.930 290.450 ;
        RECT 65.530 289.700 83.930 290.300 ;
        RECT 65.530 289.550 66.680 289.700 ;
        RECT 62.780 286.800 66.680 289.550 ;
        RECT 62.780 285.050 63.530 286.800 ;
        RECT 65.930 285.050 66.680 286.800 ;
        RECT 66.830 282.150 66.980 289.700 ;
        RECT 67.430 282.150 67.580 289.700 ;
        RECT 68.030 282.150 68.180 289.700 ;
        RECT 68.630 282.150 68.780 289.700 ;
        RECT 69.230 282.150 69.380 289.700 ;
        RECT 69.830 282.150 69.980 289.700 ;
        RECT 74.230 289.200 75.230 289.700 ;
        RECT 70.880 289.050 78.580 289.200 ;
        RECT 74.230 288.600 75.230 289.050 ;
        RECT 70.880 288.450 78.580 288.600 ;
        RECT 74.230 288.000 75.230 288.450 ;
        RECT 70.880 287.850 78.580 288.000 ;
        RECT 74.230 287.400 75.230 287.850 ;
        RECT 70.880 287.250 78.580 287.400 ;
        RECT 74.230 286.800 75.230 287.250 ;
        RECT 70.880 286.650 78.580 286.800 ;
        RECT 74.230 286.200 75.230 286.650 ;
        RECT 70.880 286.050 78.580 286.200 ;
        RECT 74.230 285.600 75.230 286.050 ;
        RECT 70.880 285.450 78.580 285.600 ;
        RECT 74.230 285.000 75.230 285.450 ;
        RECT 70.880 284.850 78.580 285.000 ;
        RECT 74.230 284.400 75.230 284.850 ;
        RECT 70.880 284.250 78.580 284.400 ;
        RECT 74.230 283.800 75.230 284.250 ;
        RECT 70.880 283.650 78.580 283.800 ;
        RECT 74.230 283.200 75.230 283.650 ;
        RECT 70.880 283.050 78.580 283.200 ;
        RECT 74.230 282.600 75.230 283.050 ;
        RECT 70.880 282.450 78.580 282.600 ;
        RECT 74.230 282.000 75.230 282.450 ;
        RECT 79.480 282.150 79.630 289.700 ;
        RECT 80.080 282.150 80.230 289.700 ;
        RECT 80.680 282.150 80.830 289.700 ;
        RECT 81.280 282.150 81.430 289.700 ;
        RECT 81.880 282.150 82.030 289.700 ;
        RECT 82.480 282.150 82.630 289.700 ;
        RECT 82.780 289.550 83.930 289.700 ;
        RECT 84.580 289.550 84.880 290.450 ;
        RECT 85.530 290.300 86.680 290.450 ;
        RECT 86.830 290.300 86.980 297.850 ;
        RECT 87.430 290.300 87.580 297.850 ;
        RECT 88.030 290.300 88.180 297.850 ;
        RECT 88.630 290.300 88.780 297.850 ;
        RECT 89.230 290.300 89.380 297.850 ;
        RECT 89.830 290.300 89.980 297.850 ;
        RECT 94.230 297.550 95.230 298.000 ;
        RECT 90.880 297.400 98.580 297.550 ;
        RECT 94.230 296.950 95.230 297.400 ;
        RECT 90.880 296.800 98.580 296.950 ;
        RECT 94.230 296.350 95.230 296.800 ;
        RECT 90.880 296.200 98.580 296.350 ;
        RECT 94.230 295.750 95.230 296.200 ;
        RECT 90.880 295.600 98.580 295.750 ;
        RECT 94.230 295.150 95.230 295.600 ;
        RECT 90.880 295.000 98.580 295.150 ;
        RECT 94.230 294.550 95.230 295.000 ;
        RECT 90.880 294.400 98.580 294.550 ;
        RECT 94.230 293.950 95.230 294.400 ;
        RECT 90.880 293.800 98.580 293.950 ;
        RECT 94.230 293.350 95.230 293.800 ;
        RECT 90.880 293.200 98.580 293.350 ;
        RECT 94.230 292.750 95.230 293.200 ;
        RECT 90.880 292.600 98.580 292.750 ;
        RECT 94.230 292.150 95.230 292.600 ;
        RECT 90.880 292.000 98.580 292.150 ;
        RECT 94.230 291.550 95.230 292.000 ;
        RECT 90.880 291.400 98.580 291.550 ;
        RECT 94.230 290.950 95.230 291.400 ;
        RECT 90.880 290.800 98.580 290.950 ;
        RECT 94.230 290.300 95.230 290.800 ;
        RECT 99.480 290.300 99.630 297.850 ;
        RECT 100.080 290.300 100.230 297.850 ;
        RECT 100.680 290.300 100.830 297.850 ;
        RECT 101.280 290.300 101.430 297.850 ;
        RECT 101.880 290.300 102.030 297.850 ;
        RECT 102.480 290.300 102.630 297.850 ;
        RECT 102.780 293.200 103.530 295.000 ;
        RECT 102.780 290.605 104.730 293.200 ;
        RECT 102.780 290.450 111.850 290.605 ;
        RECT 102.780 290.300 103.930 290.450 ;
        RECT 85.530 289.700 103.930 290.300 ;
        RECT 85.530 289.550 86.680 289.700 ;
        RECT 82.780 286.800 86.680 289.550 ;
        RECT 82.780 285.050 83.530 286.800 ;
        RECT 85.930 285.050 86.680 286.800 ;
        RECT 86.830 282.150 86.980 289.700 ;
        RECT 87.430 282.150 87.580 289.700 ;
        RECT 88.030 282.150 88.180 289.700 ;
        RECT 88.630 282.150 88.780 289.700 ;
        RECT 89.230 282.150 89.380 289.700 ;
        RECT 89.830 282.150 89.980 289.700 ;
        RECT 94.230 289.200 95.230 289.700 ;
        RECT 90.880 289.050 98.580 289.200 ;
        RECT 94.230 288.600 95.230 289.050 ;
        RECT 90.880 288.450 98.580 288.600 ;
        RECT 94.230 288.000 95.230 288.450 ;
        RECT 90.880 287.850 98.580 288.000 ;
        RECT 94.230 287.400 95.230 287.850 ;
        RECT 90.880 287.250 98.580 287.400 ;
        RECT 94.230 286.800 95.230 287.250 ;
        RECT 90.880 286.650 98.580 286.800 ;
        RECT 94.230 286.200 95.230 286.650 ;
        RECT 90.880 286.050 98.580 286.200 ;
        RECT 94.230 285.600 95.230 286.050 ;
        RECT 90.880 285.450 98.580 285.600 ;
        RECT 94.230 285.000 95.230 285.450 ;
        RECT 90.880 284.850 98.580 285.000 ;
        RECT 94.230 284.400 95.230 284.850 ;
        RECT 90.880 284.250 98.580 284.400 ;
        RECT 94.230 283.800 95.230 284.250 ;
        RECT 90.880 283.650 98.580 283.800 ;
        RECT 94.230 283.200 95.230 283.650 ;
        RECT 90.880 283.050 98.580 283.200 ;
        RECT 94.230 282.600 95.230 283.050 ;
        RECT 90.880 282.450 98.580 282.600 ;
        RECT 94.230 282.000 95.230 282.450 ;
        RECT 99.480 282.150 99.630 289.700 ;
        RECT 100.080 282.150 100.230 289.700 ;
        RECT 100.680 282.150 100.830 289.700 ;
        RECT 101.280 282.150 101.430 289.700 ;
        RECT 101.880 282.150 102.030 289.700 ;
        RECT 102.480 282.150 102.630 289.700 ;
        RECT 102.780 289.550 103.930 289.700 ;
        RECT 104.580 289.550 111.850 290.450 ;
        RECT 102.780 289.330 111.850 289.550 ;
        RECT 102.780 286.800 104.730 289.330 ;
        RECT 102.780 285.050 103.530 286.800 ;
        RECT 10.880 281.850 18.580 282.000 ;
        RECT 30.880 281.850 38.580 282.000 ;
        RECT 50.880 281.850 58.580 282.000 ;
        RECT 70.880 281.850 78.580 282.000 ;
        RECT 90.880 281.850 98.580 282.000 ;
        RECT 14.230 281.200 15.230 281.850 ;
        RECT 34.230 281.200 35.230 281.850 ;
        RECT 54.230 281.200 55.230 281.850 ;
        RECT 74.230 281.200 75.230 281.850 ;
        RECT 94.230 281.200 95.230 281.850 ;
        RECT 11.530 278.800 17.930 281.200 ;
        RECT 31.530 278.800 37.930 281.200 ;
        RECT 51.530 278.800 57.930 281.200 ;
        RECT 71.530 278.800 77.930 281.200 ;
        RECT 91.530 278.800 97.930 281.200 ;
        RECT 14.230 278.150 15.230 278.800 ;
        RECT 34.230 278.150 35.230 278.800 ;
        RECT 54.230 278.150 55.230 278.800 ;
        RECT 74.230 278.150 75.230 278.800 ;
        RECT 94.230 278.150 95.230 278.800 ;
        RECT 10.880 278.000 18.580 278.150 ;
        RECT 30.880 278.000 38.580 278.150 ;
        RECT 50.880 278.000 58.580 278.150 ;
        RECT 70.880 278.000 78.580 278.150 ;
        RECT 90.880 278.000 98.580 278.150 ;
        RECT 5.930 273.200 6.680 275.000 ;
        RECT 4.730 270.450 6.680 273.200 ;
        RECT 4.730 269.550 4.880 270.450 ;
        RECT 5.530 270.300 6.680 270.450 ;
        RECT 6.830 270.300 6.980 277.850 ;
        RECT 7.430 270.300 7.580 277.850 ;
        RECT 8.030 270.300 8.180 277.850 ;
        RECT 8.630 270.300 8.780 277.850 ;
        RECT 9.230 270.300 9.380 277.850 ;
        RECT 9.830 270.300 9.980 277.850 ;
        RECT 14.230 277.550 15.230 278.000 ;
        RECT 10.880 277.400 18.580 277.550 ;
        RECT 14.230 276.950 15.230 277.400 ;
        RECT 10.880 276.800 18.580 276.950 ;
        RECT 14.230 276.350 15.230 276.800 ;
        RECT 10.880 276.200 18.580 276.350 ;
        RECT 14.230 275.750 15.230 276.200 ;
        RECT 10.880 275.600 18.580 275.750 ;
        RECT 14.230 275.150 15.230 275.600 ;
        RECT 10.880 275.000 18.580 275.150 ;
        RECT 14.230 274.550 15.230 275.000 ;
        RECT 10.880 274.400 18.580 274.550 ;
        RECT 14.230 273.950 15.230 274.400 ;
        RECT 10.880 273.800 18.580 273.950 ;
        RECT 14.230 273.350 15.230 273.800 ;
        RECT 10.880 273.200 18.580 273.350 ;
        RECT 14.230 272.750 15.230 273.200 ;
        RECT 10.880 272.600 18.580 272.750 ;
        RECT 14.230 272.150 15.230 272.600 ;
        RECT 10.880 272.000 18.580 272.150 ;
        RECT 14.230 271.550 15.230 272.000 ;
        RECT 10.880 271.400 18.580 271.550 ;
        RECT 14.230 270.950 15.230 271.400 ;
        RECT 10.880 270.800 18.580 270.950 ;
        RECT 14.230 270.300 15.230 270.800 ;
        RECT 19.480 270.300 19.630 277.850 ;
        RECT 20.080 270.300 20.230 277.850 ;
        RECT 20.680 270.300 20.830 277.850 ;
        RECT 21.280 270.300 21.430 277.850 ;
        RECT 21.880 270.300 22.030 277.850 ;
        RECT 22.480 270.300 22.630 277.850 ;
        RECT 22.780 273.200 23.530 275.000 ;
        RECT 25.930 273.200 26.680 275.000 ;
        RECT 22.780 270.450 26.680 273.200 ;
        RECT 22.780 270.300 23.930 270.450 ;
        RECT 5.530 269.700 23.930 270.300 ;
        RECT 5.530 269.550 6.680 269.700 ;
        RECT 4.730 266.800 6.680 269.550 ;
        RECT 5.930 265.050 6.680 266.800 ;
        RECT 6.830 262.150 6.980 269.700 ;
        RECT 7.430 262.150 7.580 269.700 ;
        RECT 8.030 262.150 8.180 269.700 ;
        RECT 8.630 262.150 8.780 269.700 ;
        RECT 9.230 262.150 9.380 269.700 ;
        RECT 9.830 262.150 9.980 269.700 ;
        RECT 14.230 269.200 15.230 269.700 ;
        RECT 10.880 269.050 18.580 269.200 ;
        RECT 14.230 268.600 15.230 269.050 ;
        RECT 10.880 268.450 18.580 268.600 ;
        RECT 14.230 268.000 15.230 268.450 ;
        RECT 10.880 267.850 18.580 268.000 ;
        RECT 14.230 267.400 15.230 267.850 ;
        RECT 10.880 267.250 18.580 267.400 ;
        RECT 14.230 266.800 15.230 267.250 ;
        RECT 10.880 266.650 18.580 266.800 ;
        RECT 14.230 266.200 15.230 266.650 ;
        RECT 10.880 266.050 18.580 266.200 ;
        RECT 14.230 265.600 15.230 266.050 ;
        RECT 10.880 265.450 18.580 265.600 ;
        RECT 14.230 265.000 15.230 265.450 ;
        RECT 10.880 264.850 18.580 265.000 ;
        RECT 14.230 264.400 15.230 264.850 ;
        RECT 10.880 264.250 18.580 264.400 ;
        RECT 14.230 263.800 15.230 264.250 ;
        RECT 10.880 263.650 18.580 263.800 ;
        RECT 14.230 263.200 15.230 263.650 ;
        RECT 10.880 263.050 18.580 263.200 ;
        RECT 14.230 262.600 15.230 263.050 ;
        RECT 10.880 262.450 18.580 262.600 ;
        RECT 14.230 262.000 15.230 262.450 ;
        RECT 19.480 262.150 19.630 269.700 ;
        RECT 20.080 262.150 20.230 269.700 ;
        RECT 20.680 262.150 20.830 269.700 ;
        RECT 21.280 262.150 21.430 269.700 ;
        RECT 21.880 262.150 22.030 269.700 ;
        RECT 22.480 262.150 22.630 269.700 ;
        RECT 22.780 269.550 23.930 269.700 ;
        RECT 24.580 269.550 24.880 270.450 ;
        RECT 25.530 270.300 26.680 270.450 ;
        RECT 26.830 270.300 26.980 277.850 ;
        RECT 27.430 270.300 27.580 277.850 ;
        RECT 28.030 270.300 28.180 277.850 ;
        RECT 28.630 270.300 28.780 277.850 ;
        RECT 29.230 270.300 29.380 277.850 ;
        RECT 29.830 270.300 29.980 277.850 ;
        RECT 34.230 277.550 35.230 278.000 ;
        RECT 30.880 277.400 38.580 277.550 ;
        RECT 34.230 276.950 35.230 277.400 ;
        RECT 30.880 276.800 38.580 276.950 ;
        RECT 34.230 276.350 35.230 276.800 ;
        RECT 30.880 276.200 38.580 276.350 ;
        RECT 34.230 275.750 35.230 276.200 ;
        RECT 30.880 275.600 38.580 275.750 ;
        RECT 34.230 275.150 35.230 275.600 ;
        RECT 30.880 275.000 38.580 275.150 ;
        RECT 34.230 274.550 35.230 275.000 ;
        RECT 30.880 274.400 38.580 274.550 ;
        RECT 34.230 273.950 35.230 274.400 ;
        RECT 30.880 273.800 38.580 273.950 ;
        RECT 34.230 273.350 35.230 273.800 ;
        RECT 30.880 273.200 38.580 273.350 ;
        RECT 34.230 272.750 35.230 273.200 ;
        RECT 30.880 272.600 38.580 272.750 ;
        RECT 34.230 272.150 35.230 272.600 ;
        RECT 30.880 272.000 38.580 272.150 ;
        RECT 34.230 271.550 35.230 272.000 ;
        RECT 30.880 271.400 38.580 271.550 ;
        RECT 34.230 270.950 35.230 271.400 ;
        RECT 30.880 270.800 38.580 270.950 ;
        RECT 34.230 270.300 35.230 270.800 ;
        RECT 39.480 270.300 39.630 277.850 ;
        RECT 40.080 270.300 40.230 277.850 ;
        RECT 40.680 270.300 40.830 277.850 ;
        RECT 41.280 270.300 41.430 277.850 ;
        RECT 41.880 270.300 42.030 277.850 ;
        RECT 42.480 270.300 42.630 277.850 ;
        RECT 42.780 273.200 43.530 275.000 ;
        RECT 45.930 273.200 46.680 275.000 ;
        RECT 42.780 270.450 46.680 273.200 ;
        RECT 42.780 270.300 43.930 270.450 ;
        RECT 25.530 269.700 43.930 270.300 ;
        RECT 25.530 269.550 26.680 269.700 ;
        RECT 22.780 266.800 26.680 269.550 ;
        RECT 22.780 265.050 23.530 266.800 ;
        RECT 25.930 265.050 26.680 266.800 ;
        RECT 26.830 262.150 26.980 269.700 ;
        RECT 27.430 262.150 27.580 269.700 ;
        RECT 28.030 262.150 28.180 269.700 ;
        RECT 28.630 262.150 28.780 269.700 ;
        RECT 29.230 262.150 29.380 269.700 ;
        RECT 29.830 262.150 29.980 269.700 ;
        RECT 34.230 269.200 35.230 269.700 ;
        RECT 30.880 269.050 38.580 269.200 ;
        RECT 34.230 268.600 35.230 269.050 ;
        RECT 30.880 268.450 38.580 268.600 ;
        RECT 34.230 268.000 35.230 268.450 ;
        RECT 30.880 267.850 38.580 268.000 ;
        RECT 34.230 267.400 35.230 267.850 ;
        RECT 30.880 267.250 38.580 267.400 ;
        RECT 34.230 266.800 35.230 267.250 ;
        RECT 30.880 266.650 38.580 266.800 ;
        RECT 34.230 266.200 35.230 266.650 ;
        RECT 30.880 266.050 38.580 266.200 ;
        RECT 34.230 265.600 35.230 266.050 ;
        RECT 30.880 265.450 38.580 265.600 ;
        RECT 34.230 265.000 35.230 265.450 ;
        RECT 30.880 264.850 38.580 265.000 ;
        RECT 34.230 264.400 35.230 264.850 ;
        RECT 30.880 264.250 38.580 264.400 ;
        RECT 34.230 263.800 35.230 264.250 ;
        RECT 30.880 263.650 38.580 263.800 ;
        RECT 34.230 263.200 35.230 263.650 ;
        RECT 30.880 263.050 38.580 263.200 ;
        RECT 34.230 262.600 35.230 263.050 ;
        RECT 30.880 262.450 38.580 262.600 ;
        RECT 34.230 262.000 35.230 262.450 ;
        RECT 39.480 262.150 39.630 269.700 ;
        RECT 40.080 262.150 40.230 269.700 ;
        RECT 40.680 262.150 40.830 269.700 ;
        RECT 41.280 262.150 41.430 269.700 ;
        RECT 41.880 262.150 42.030 269.700 ;
        RECT 42.480 262.150 42.630 269.700 ;
        RECT 42.780 269.550 43.930 269.700 ;
        RECT 44.580 269.550 44.880 270.450 ;
        RECT 45.530 270.300 46.680 270.450 ;
        RECT 46.830 270.300 46.980 277.850 ;
        RECT 47.430 270.300 47.580 277.850 ;
        RECT 48.030 270.300 48.180 277.850 ;
        RECT 48.630 270.300 48.780 277.850 ;
        RECT 49.230 270.300 49.380 277.850 ;
        RECT 49.830 270.300 49.980 277.850 ;
        RECT 54.230 277.550 55.230 278.000 ;
        RECT 50.880 277.400 58.580 277.550 ;
        RECT 54.230 276.950 55.230 277.400 ;
        RECT 50.880 276.800 58.580 276.950 ;
        RECT 54.230 276.350 55.230 276.800 ;
        RECT 50.880 276.200 58.580 276.350 ;
        RECT 54.230 275.750 55.230 276.200 ;
        RECT 50.880 275.600 58.580 275.750 ;
        RECT 54.230 275.150 55.230 275.600 ;
        RECT 50.880 275.000 58.580 275.150 ;
        RECT 54.230 274.550 55.230 275.000 ;
        RECT 50.880 274.400 58.580 274.550 ;
        RECT 54.230 273.950 55.230 274.400 ;
        RECT 50.880 273.800 58.580 273.950 ;
        RECT 54.230 273.350 55.230 273.800 ;
        RECT 50.880 273.200 58.580 273.350 ;
        RECT 54.230 272.750 55.230 273.200 ;
        RECT 50.880 272.600 58.580 272.750 ;
        RECT 54.230 272.150 55.230 272.600 ;
        RECT 50.880 272.000 58.580 272.150 ;
        RECT 54.230 271.550 55.230 272.000 ;
        RECT 50.880 271.400 58.580 271.550 ;
        RECT 54.230 270.950 55.230 271.400 ;
        RECT 50.880 270.800 58.580 270.950 ;
        RECT 54.230 270.300 55.230 270.800 ;
        RECT 59.480 270.300 59.630 277.850 ;
        RECT 60.080 270.300 60.230 277.850 ;
        RECT 60.680 270.300 60.830 277.850 ;
        RECT 61.280 270.300 61.430 277.850 ;
        RECT 61.880 270.300 62.030 277.850 ;
        RECT 62.480 270.300 62.630 277.850 ;
        RECT 62.780 273.200 63.530 275.000 ;
        RECT 65.930 273.200 66.680 275.000 ;
        RECT 62.780 270.450 66.680 273.200 ;
        RECT 62.780 270.300 63.930 270.450 ;
        RECT 45.530 269.700 63.930 270.300 ;
        RECT 45.530 269.550 46.680 269.700 ;
        RECT 42.780 266.800 46.680 269.550 ;
        RECT 42.780 265.050 43.530 266.800 ;
        RECT 45.930 265.050 46.680 266.800 ;
        RECT 46.830 262.150 46.980 269.700 ;
        RECT 47.430 262.150 47.580 269.700 ;
        RECT 48.030 262.150 48.180 269.700 ;
        RECT 48.630 262.150 48.780 269.700 ;
        RECT 49.230 262.150 49.380 269.700 ;
        RECT 49.830 262.150 49.980 269.700 ;
        RECT 54.230 269.200 55.230 269.700 ;
        RECT 50.880 269.050 58.580 269.200 ;
        RECT 54.230 268.600 55.230 269.050 ;
        RECT 50.880 268.450 58.580 268.600 ;
        RECT 54.230 268.000 55.230 268.450 ;
        RECT 50.880 267.850 58.580 268.000 ;
        RECT 54.230 267.400 55.230 267.850 ;
        RECT 50.880 267.250 58.580 267.400 ;
        RECT 54.230 266.800 55.230 267.250 ;
        RECT 50.880 266.650 58.580 266.800 ;
        RECT 54.230 266.200 55.230 266.650 ;
        RECT 50.880 266.050 58.580 266.200 ;
        RECT 54.230 265.600 55.230 266.050 ;
        RECT 50.880 265.450 58.580 265.600 ;
        RECT 54.230 265.000 55.230 265.450 ;
        RECT 50.880 264.850 58.580 265.000 ;
        RECT 54.230 264.400 55.230 264.850 ;
        RECT 50.880 264.250 58.580 264.400 ;
        RECT 54.230 263.800 55.230 264.250 ;
        RECT 50.880 263.650 58.580 263.800 ;
        RECT 54.230 263.200 55.230 263.650 ;
        RECT 50.880 263.050 58.580 263.200 ;
        RECT 54.230 262.600 55.230 263.050 ;
        RECT 50.880 262.450 58.580 262.600 ;
        RECT 54.230 262.000 55.230 262.450 ;
        RECT 59.480 262.150 59.630 269.700 ;
        RECT 60.080 262.150 60.230 269.700 ;
        RECT 60.680 262.150 60.830 269.700 ;
        RECT 61.280 262.150 61.430 269.700 ;
        RECT 61.880 262.150 62.030 269.700 ;
        RECT 62.480 262.150 62.630 269.700 ;
        RECT 62.780 269.550 63.930 269.700 ;
        RECT 64.580 269.550 64.880 270.450 ;
        RECT 65.530 270.300 66.680 270.450 ;
        RECT 66.830 270.300 66.980 277.850 ;
        RECT 67.430 270.300 67.580 277.850 ;
        RECT 68.030 270.300 68.180 277.850 ;
        RECT 68.630 270.300 68.780 277.850 ;
        RECT 69.230 270.300 69.380 277.850 ;
        RECT 69.830 270.300 69.980 277.850 ;
        RECT 74.230 277.550 75.230 278.000 ;
        RECT 70.880 277.400 78.580 277.550 ;
        RECT 74.230 276.950 75.230 277.400 ;
        RECT 70.880 276.800 78.580 276.950 ;
        RECT 74.230 276.350 75.230 276.800 ;
        RECT 70.880 276.200 78.580 276.350 ;
        RECT 74.230 275.750 75.230 276.200 ;
        RECT 70.880 275.600 78.580 275.750 ;
        RECT 74.230 275.150 75.230 275.600 ;
        RECT 70.880 275.000 78.580 275.150 ;
        RECT 74.230 274.550 75.230 275.000 ;
        RECT 70.880 274.400 78.580 274.550 ;
        RECT 74.230 273.950 75.230 274.400 ;
        RECT 70.880 273.800 78.580 273.950 ;
        RECT 74.230 273.350 75.230 273.800 ;
        RECT 70.880 273.200 78.580 273.350 ;
        RECT 74.230 272.750 75.230 273.200 ;
        RECT 70.880 272.600 78.580 272.750 ;
        RECT 74.230 272.150 75.230 272.600 ;
        RECT 70.880 272.000 78.580 272.150 ;
        RECT 74.230 271.550 75.230 272.000 ;
        RECT 70.880 271.400 78.580 271.550 ;
        RECT 74.230 270.950 75.230 271.400 ;
        RECT 70.880 270.800 78.580 270.950 ;
        RECT 74.230 270.300 75.230 270.800 ;
        RECT 79.480 270.300 79.630 277.850 ;
        RECT 80.080 270.300 80.230 277.850 ;
        RECT 80.680 270.300 80.830 277.850 ;
        RECT 81.280 270.300 81.430 277.850 ;
        RECT 81.880 270.300 82.030 277.850 ;
        RECT 82.480 270.300 82.630 277.850 ;
        RECT 82.780 273.200 83.530 275.000 ;
        RECT 85.930 273.200 86.680 275.000 ;
        RECT 82.780 270.450 86.680 273.200 ;
        RECT 82.780 270.300 83.930 270.450 ;
        RECT 65.530 269.700 83.930 270.300 ;
        RECT 65.530 269.550 66.680 269.700 ;
        RECT 62.780 266.800 66.680 269.550 ;
        RECT 62.780 265.050 63.530 266.800 ;
        RECT 65.930 265.050 66.680 266.800 ;
        RECT 66.830 262.150 66.980 269.700 ;
        RECT 67.430 262.150 67.580 269.700 ;
        RECT 68.030 262.150 68.180 269.700 ;
        RECT 68.630 262.150 68.780 269.700 ;
        RECT 69.230 262.150 69.380 269.700 ;
        RECT 69.830 262.150 69.980 269.700 ;
        RECT 74.230 269.200 75.230 269.700 ;
        RECT 70.880 269.050 78.580 269.200 ;
        RECT 74.230 268.600 75.230 269.050 ;
        RECT 70.880 268.450 78.580 268.600 ;
        RECT 74.230 268.000 75.230 268.450 ;
        RECT 70.880 267.850 78.580 268.000 ;
        RECT 74.230 267.400 75.230 267.850 ;
        RECT 70.880 267.250 78.580 267.400 ;
        RECT 74.230 266.800 75.230 267.250 ;
        RECT 70.880 266.650 78.580 266.800 ;
        RECT 74.230 266.200 75.230 266.650 ;
        RECT 70.880 266.050 78.580 266.200 ;
        RECT 74.230 265.600 75.230 266.050 ;
        RECT 70.880 265.450 78.580 265.600 ;
        RECT 74.230 265.000 75.230 265.450 ;
        RECT 70.880 264.850 78.580 265.000 ;
        RECT 74.230 264.400 75.230 264.850 ;
        RECT 70.880 264.250 78.580 264.400 ;
        RECT 74.230 263.800 75.230 264.250 ;
        RECT 70.880 263.650 78.580 263.800 ;
        RECT 74.230 263.200 75.230 263.650 ;
        RECT 70.880 263.050 78.580 263.200 ;
        RECT 74.230 262.600 75.230 263.050 ;
        RECT 70.880 262.450 78.580 262.600 ;
        RECT 74.230 262.000 75.230 262.450 ;
        RECT 79.480 262.150 79.630 269.700 ;
        RECT 80.080 262.150 80.230 269.700 ;
        RECT 80.680 262.150 80.830 269.700 ;
        RECT 81.280 262.150 81.430 269.700 ;
        RECT 81.880 262.150 82.030 269.700 ;
        RECT 82.480 262.150 82.630 269.700 ;
        RECT 82.780 269.550 83.930 269.700 ;
        RECT 84.580 269.550 84.880 270.450 ;
        RECT 85.530 270.300 86.680 270.450 ;
        RECT 86.830 270.300 86.980 277.850 ;
        RECT 87.430 270.300 87.580 277.850 ;
        RECT 88.030 270.300 88.180 277.850 ;
        RECT 88.630 270.300 88.780 277.850 ;
        RECT 89.230 270.300 89.380 277.850 ;
        RECT 89.830 270.300 89.980 277.850 ;
        RECT 94.230 277.550 95.230 278.000 ;
        RECT 90.880 277.400 98.580 277.550 ;
        RECT 94.230 276.950 95.230 277.400 ;
        RECT 90.880 276.800 98.580 276.950 ;
        RECT 94.230 276.350 95.230 276.800 ;
        RECT 90.880 276.200 98.580 276.350 ;
        RECT 94.230 275.750 95.230 276.200 ;
        RECT 90.880 275.600 98.580 275.750 ;
        RECT 94.230 275.150 95.230 275.600 ;
        RECT 90.880 275.000 98.580 275.150 ;
        RECT 94.230 274.550 95.230 275.000 ;
        RECT 90.880 274.400 98.580 274.550 ;
        RECT 94.230 273.950 95.230 274.400 ;
        RECT 90.880 273.800 98.580 273.950 ;
        RECT 94.230 273.350 95.230 273.800 ;
        RECT 90.880 273.200 98.580 273.350 ;
        RECT 94.230 272.750 95.230 273.200 ;
        RECT 90.880 272.600 98.580 272.750 ;
        RECT 94.230 272.150 95.230 272.600 ;
        RECT 90.880 272.000 98.580 272.150 ;
        RECT 94.230 271.550 95.230 272.000 ;
        RECT 90.880 271.400 98.580 271.550 ;
        RECT 94.230 270.950 95.230 271.400 ;
        RECT 90.880 270.800 98.580 270.950 ;
        RECT 94.230 270.300 95.230 270.800 ;
        RECT 99.480 270.300 99.630 277.850 ;
        RECT 100.080 270.300 100.230 277.850 ;
        RECT 100.680 270.300 100.830 277.850 ;
        RECT 101.280 270.300 101.430 277.850 ;
        RECT 101.880 270.300 102.030 277.850 ;
        RECT 102.480 270.300 102.630 277.850 ;
        RECT 102.780 273.200 103.530 275.000 ;
        RECT 102.780 270.520 104.730 273.200 ;
        RECT 102.780 270.450 111.850 270.520 ;
        RECT 102.780 270.300 103.930 270.450 ;
        RECT 85.530 269.700 103.930 270.300 ;
        RECT 85.530 269.550 86.680 269.700 ;
        RECT 82.780 266.800 86.680 269.550 ;
        RECT 82.780 265.050 83.530 266.800 ;
        RECT 85.930 265.050 86.680 266.800 ;
        RECT 86.830 262.150 86.980 269.700 ;
        RECT 87.430 262.150 87.580 269.700 ;
        RECT 88.030 262.150 88.180 269.700 ;
        RECT 88.630 262.150 88.780 269.700 ;
        RECT 89.230 262.150 89.380 269.700 ;
        RECT 89.830 262.150 89.980 269.700 ;
        RECT 94.230 269.200 95.230 269.700 ;
        RECT 90.880 269.050 98.580 269.200 ;
        RECT 94.230 268.600 95.230 269.050 ;
        RECT 90.880 268.450 98.580 268.600 ;
        RECT 94.230 268.000 95.230 268.450 ;
        RECT 90.880 267.850 98.580 268.000 ;
        RECT 94.230 267.400 95.230 267.850 ;
        RECT 90.880 267.250 98.580 267.400 ;
        RECT 94.230 266.800 95.230 267.250 ;
        RECT 90.880 266.650 98.580 266.800 ;
        RECT 94.230 266.200 95.230 266.650 ;
        RECT 90.880 266.050 98.580 266.200 ;
        RECT 94.230 265.600 95.230 266.050 ;
        RECT 90.880 265.450 98.580 265.600 ;
        RECT 94.230 265.000 95.230 265.450 ;
        RECT 90.880 264.850 98.580 265.000 ;
        RECT 94.230 264.400 95.230 264.850 ;
        RECT 90.880 264.250 98.580 264.400 ;
        RECT 94.230 263.800 95.230 264.250 ;
        RECT 90.880 263.650 98.580 263.800 ;
        RECT 94.230 263.200 95.230 263.650 ;
        RECT 90.880 263.050 98.580 263.200 ;
        RECT 94.230 262.600 95.230 263.050 ;
        RECT 90.880 262.450 98.580 262.600 ;
        RECT 94.230 262.000 95.230 262.450 ;
        RECT 99.480 262.150 99.630 269.700 ;
        RECT 100.080 262.150 100.230 269.700 ;
        RECT 100.680 262.150 100.830 269.700 ;
        RECT 101.280 262.150 101.430 269.700 ;
        RECT 101.880 262.150 102.030 269.700 ;
        RECT 102.480 262.150 102.630 269.700 ;
        RECT 102.780 269.550 103.930 269.700 ;
        RECT 104.580 269.550 111.850 270.450 ;
        RECT 102.780 269.245 111.850 269.550 ;
        RECT 102.780 266.800 104.730 269.245 ;
        RECT 102.780 265.050 103.530 266.800 ;
        RECT 10.880 261.850 18.580 262.000 ;
        RECT 30.880 261.850 38.580 262.000 ;
        RECT 50.880 261.850 58.580 262.000 ;
        RECT 70.880 261.850 78.580 262.000 ;
        RECT 90.880 261.850 98.580 262.000 ;
        RECT 14.230 261.200 15.230 261.850 ;
        RECT 34.230 261.200 35.230 261.850 ;
        RECT 54.230 261.200 55.230 261.850 ;
        RECT 74.230 261.200 75.230 261.850 ;
        RECT 94.230 261.200 95.230 261.850 ;
        RECT 11.530 258.800 17.930 261.200 ;
        RECT 31.530 258.800 37.930 261.200 ;
        RECT 51.530 258.800 57.930 261.200 ;
        RECT 71.530 258.800 77.930 261.200 ;
        RECT 91.530 258.800 97.930 261.200 ;
        RECT 14.230 258.150 15.230 258.800 ;
        RECT 34.230 258.150 35.230 258.800 ;
        RECT 54.230 258.150 55.230 258.800 ;
        RECT 74.230 258.150 75.230 258.800 ;
        RECT 94.230 258.150 95.230 258.800 ;
        RECT 10.880 258.000 18.580 258.150 ;
        RECT 30.880 258.000 38.580 258.150 ;
        RECT 50.880 258.000 58.580 258.150 ;
        RECT 70.880 258.000 78.580 258.150 ;
        RECT 90.880 258.000 98.580 258.150 ;
        RECT 5.930 253.200 6.680 255.000 ;
        RECT 4.730 250.450 6.680 253.200 ;
        RECT 4.730 249.550 4.880 250.450 ;
        RECT 5.530 250.300 6.680 250.450 ;
        RECT 6.830 250.300 6.980 257.850 ;
        RECT 7.430 250.300 7.580 257.850 ;
        RECT 8.030 250.300 8.180 257.850 ;
        RECT 8.630 250.300 8.780 257.850 ;
        RECT 9.230 250.300 9.380 257.850 ;
        RECT 9.830 250.300 9.980 257.850 ;
        RECT 14.230 257.550 15.230 258.000 ;
        RECT 10.880 257.400 18.580 257.550 ;
        RECT 14.230 256.950 15.230 257.400 ;
        RECT 10.880 256.800 18.580 256.950 ;
        RECT 14.230 256.350 15.230 256.800 ;
        RECT 10.880 256.200 18.580 256.350 ;
        RECT 14.230 255.750 15.230 256.200 ;
        RECT 10.880 255.600 18.580 255.750 ;
        RECT 14.230 255.150 15.230 255.600 ;
        RECT 10.880 255.000 18.580 255.150 ;
        RECT 14.230 254.550 15.230 255.000 ;
        RECT 10.880 254.400 18.580 254.550 ;
        RECT 14.230 253.950 15.230 254.400 ;
        RECT 10.880 253.800 18.580 253.950 ;
        RECT 14.230 253.350 15.230 253.800 ;
        RECT 10.880 253.200 18.580 253.350 ;
        RECT 14.230 252.750 15.230 253.200 ;
        RECT 10.880 252.600 18.580 252.750 ;
        RECT 14.230 252.150 15.230 252.600 ;
        RECT 10.880 252.000 18.580 252.150 ;
        RECT 14.230 251.550 15.230 252.000 ;
        RECT 10.880 251.400 18.580 251.550 ;
        RECT 14.230 250.950 15.230 251.400 ;
        RECT 10.880 250.800 18.580 250.950 ;
        RECT 14.230 250.300 15.230 250.800 ;
        RECT 19.480 250.300 19.630 257.850 ;
        RECT 20.080 250.300 20.230 257.850 ;
        RECT 20.680 250.300 20.830 257.850 ;
        RECT 21.280 250.300 21.430 257.850 ;
        RECT 21.880 250.300 22.030 257.850 ;
        RECT 22.480 250.300 22.630 257.850 ;
        RECT 22.780 253.200 23.530 255.000 ;
        RECT 25.930 253.200 26.680 255.000 ;
        RECT 22.780 250.450 26.680 253.200 ;
        RECT 22.780 250.300 23.930 250.450 ;
        RECT 5.530 249.700 23.930 250.300 ;
        RECT 5.530 249.550 6.680 249.700 ;
        RECT 4.730 246.800 6.680 249.550 ;
        RECT 5.930 245.050 6.680 246.800 ;
        RECT 6.830 242.150 6.980 249.700 ;
        RECT 7.430 242.150 7.580 249.700 ;
        RECT 8.030 242.150 8.180 249.700 ;
        RECT 8.630 242.150 8.780 249.700 ;
        RECT 9.230 242.150 9.380 249.700 ;
        RECT 9.830 242.150 9.980 249.700 ;
        RECT 14.230 249.200 15.230 249.700 ;
        RECT 10.880 249.050 18.580 249.200 ;
        RECT 14.230 248.600 15.230 249.050 ;
        RECT 10.880 248.450 18.580 248.600 ;
        RECT 14.230 248.000 15.230 248.450 ;
        RECT 10.880 247.850 18.580 248.000 ;
        RECT 14.230 247.400 15.230 247.850 ;
        RECT 10.880 247.250 18.580 247.400 ;
        RECT 14.230 246.800 15.230 247.250 ;
        RECT 10.880 246.650 18.580 246.800 ;
        RECT 14.230 246.200 15.230 246.650 ;
        RECT 10.880 246.050 18.580 246.200 ;
        RECT 14.230 245.600 15.230 246.050 ;
        RECT 10.880 245.450 18.580 245.600 ;
        RECT 14.230 245.000 15.230 245.450 ;
        RECT 10.880 244.850 18.580 245.000 ;
        RECT 14.230 244.400 15.230 244.850 ;
        RECT 10.880 244.250 18.580 244.400 ;
        RECT 14.230 243.800 15.230 244.250 ;
        RECT 10.880 243.650 18.580 243.800 ;
        RECT 14.230 243.200 15.230 243.650 ;
        RECT 10.880 243.050 18.580 243.200 ;
        RECT 14.230 242.600 15.230 243.050 ;
        RECT 10.880 242.450 18.580 242.600 ;
        RECT 14.230 242.000 15.230 242.450 ;
        RECT 19.480 242.150 19.630 249.700 ;
        RECT 20.080 242.150 20.230 249.700 ;
        RECT 20.680 242.150 20.830 249.700 ;
        RECT 21.280 242.150 21.430 249.700 ;
        RECT 21.880 242.150 22.030 249.700 ;
        RECT 22.480 242.150 22.630 249.700 ;
        RECT 22.780 249.550 23.930 249.700 ;
        RECT 24.580 249.550 24.880 250.450 ;
        RECT 25.530 250.300 26.680 250.450 ;
        RECT 26.830 250.300 26.980 257.850 ;
        RECT 27.430 250.300 27.580 257.850 ;
        RECT 28.030 250.300 28.180 257.850 ;
        RECT 28.630 250.300 28.780 257.850 ;
        RECT 29.230 250.300 29.380 257.850 ;
        RECT 29.830 250.300 29.980 257.850 ;
        RECT 34.230 257.550 35.230 258.000 ;
        RECT 30.880 257.400 38.580 257.550 ;
        RECT 34.230 256.950 35.230 257.400 ;
        RECT 30.880 256.800 38.580 256.950 ;
        RECT 34.230 256.350 35.230 256.800 ;
        RECT 30.880 256.200 38.580 256.350 ;
        RECT 34.230 255.750 35.230 256.200 ;
        RECT 30.880 255.600 38.580 255.750 ;
        RECT 34.230 255.150 35.230 255.600 ;
        RECT 30.880 255.000 38.580 255.150 ;
        RECT 34.230 254.550 35.230 255.000 ;
        RECT 30.880 254.400 38.580 254.550 ;
        RECT 34.230 253.950 35.230 254.400 ;
        RECT 30.880 253.800 38.580 253.950 ;
        RECT 34.230 253.350 35.230 253.800 ;
        RECT 30.880 253.200 38.580 253.350 ;
        RECT 34.230 252.750 35.230 253.200 ;
        RECT 30.880 252.600 38.580 252.750 ;
        RECT 34.230 252.150 35.230 252.600 ;
        RECT 30.880 252.000 38.580 252.150 ;
        RECT 34.230 251.550 35.230 252.000 ;
        RECT 30.880 251.400 38.580 251.550 ;
        RECT 34.230 250.950 35.230 251.400 ;
        RECT 30.880 250.800 38.580 250.950 ;
        RECT 34.230 250.300 35.230 250.800 ;
        RECT 39.480 250.300 39.630 257.850 ;
        RECT 40.080 250.300 40.230 257.850 ;
        RECT 40.680 250.300 40.830 257.850 ;
        RECT 41.280 250.300 41.430 257.850 ;
        RECT 41.880 250.300 42.030 257.850 ;
        RECT 42.480 250.300 42.630 257.850 ;
        RECT 42.780 253.200 43.530 255.000 ;
        RECT 45.930 253.200 46.680 255.000 ;
        RECT 42.780 250.450 46.680 253.200 ;
        RECT 42.780 250.300 43.930 250.450 ;
        RECT 25.530 249.700 43.930 250.300 ;
        RECT 25.530 249.550 26.680 249.700 ;
        RECT 22.780 246.800 26.680 249.550 ;
        RECT 22.780 245.050 23.530 246.800 ;
        RECT 25.930 245.050 26.680 246.800 ;
        RECT 26.830 242.150 26.980 249.700 ;
        RECT 27.430 242.150 27.580 249.700 ;
        RECT 28.030 242.150 28.180 249.700 ;
        RECT 28.630 242.150 28.780 249.700 ;
        RECT 29.230 242.150 29.380 249.700 ;
        RECT 29.830 242.150 29.980 249.700 ;
        RECT 34.230 249.200 35.230 249.700 ;
        RECT 30.880 249.050 38.580 249.200 ;
        RECT 34.230 248.600 35.230 249.050 ;
        RECT 30.880 248.450 38.580 248.600 ;
        RECT 34.230 248.000 35.230 248.450 ;
        RECT 30.880 247.850 38.580 248.000 ;
        RECT 34.230 247.400 35.230 247.850 ;
        RECT 30.880 247.250 38.580 247.400 ;
        RECT 34.230 246.800 35.230 247.250 ;
        RECT 30.880 246.650 38.580 246.800 ;
        RECT 34.230 246.200 35.230 246.650 ;
        RECT 30.880 246.050 38.580 246.200 ;
        RECT 34.230 245.600 35.230 246.050 ;
        RECT 30.880 245.450 38.580 245.600 ;
        RECT 34.230 245.000 35.230 245.450 ;
        RECT 30.880 244.850 38.580 245.000 ;
        RECT 34.230 244.400 35.230 244.850 ;
        RECT 30.880 244.250 38.580 244.400 ;
        RECT 34.230 243.800 35.230 244.250 ;
        RECT 30.880 243.650 38.580 243.800 ;
        RECT 34.230 243.200 35.230 243.650 ;
        RECT 30.880 243.050 38.580 243.200 ;
        RECT 34.230 242.600 35.230 243.050 ;
        RECT 30.880 242.450 38.580 242.600 ;
        RECT 34.230 242.000 35.230 242.450 ;
        RECT 39.480 242.150 39.630 249.700 ;
        RECT 40.080 242.150 40.230 249.700 ;
        RECT 40.680 242.150 40.830 249.700 ;
        RECT 41.280 242.150 41.430 249.700 ;
        RECT 41.880 242.150 42.030 249.700 ;
        RECT 42.480 242.150 42.630 249.700 ;
        RECT 42.780 249.550 43.930 249.700 ;
        RECT 44.580 249.550 44.880 250.450 ;
        RECT 45.530 250.300 46.680 250.450 ;
        RECT 46.830 250.300 46.980 257.850 ;
        RECT 47.430 250.300 47.580 257.850 ;
        RECT 48.030 250.300 48.180 257.850 ;
        RECT 48.630 250.300 48.780 257.850 ;
        RECT 49.230 250.300 49.380 257.850 ;
        RECT 49.830 250.300 49.980 257.850 ;
        RECT 54.230 257.550 55.230 258.000 ;
        RECT 50.880 257.400 58.580 257.550 ;
        RECT 54.230 256.950 55.230 257.400 ;
        RECT 50.880 256.800 58.580 256.950 ;
        RECT 54.230 256.350 55.230 256.800 ;
        RECT 50.880 256.200 58.580 256.350 ;
        RECT 54.230 255.750 55.230 256.200 ;
        RECT 50.880 255.600 58.580 255.750 ;
        RECT 54.230 255.150 55.230 255.600 ;
        RECT 50.880 255.000 58.580 255.150 ;
        RECT 54.230 254.550 55.230 255.000 ;
        RECT 50.880 254.400 58.580 254.550 ;
        RECT 54.230 253.950 55.230 254.400 ;
        RECT 50.880 253.800 58.580 253.950 ;
        RECT 54.230 253.350 55.230 253.800 ;
        RECT 50.880 253.200 58.580 253.350 ;
        RECT 54.230 252.750 55.230 253.200 ;
        RECT 50.880 252.600 58.580 252.750 ;
        RECT 54.230 252.150 55.230 252.600 ;
        RECT 50.880 252.000 58.580 252.150 ;
        RECT 54.230 251.550 55.230 252.000 ;
        RECT 50.880 251.400 58.580 251.550 ;
        RECT 54.230 250.950 55.230 251.400 ;
        RECT 50.880 250.800 58.580 250.950 ;
        RECT 54.230 250.300 55.230 250.800 ;
        RECT 59.480 250.300 59.630 257.850 ;
        RECT 60.080 250.300 60.230 257.850 ;
        RECT 60.680 250.300 60.830 257.850 ;
        RECT 61.280 250.300 61.430 257.850 ;
        RECT 61.880 250.300 62.030 257.850 ;
        RECT 62.480 250.300 62.630 257.850 ;
        RECT 62.780 253.200 63.530 255.000 ;
        RECT 65.930 253.200 66.680 255.000 ;
        RECT 62.780 250.450 66.680 253.200 ;
        RECT 62.780 250.300 63.930 250.450 ;
        RECT 45.530 249.700 63.930 250.300 ;
        RECT 45.530 249.550 46.680 249.700 ;
        RECT 42.780 246.800 46.680 249.550 ;
        RECT 42.780 245.050 43.530 246.800 ;
        RECT 45.930 245.050 46.680 246.800 ;
        RECT 46.830 242.150 46.980 249.700 ;
        RECT 47.430 242.150 47.580 249.700 ;
        RECT 48.030 242.150 48.180 249.700 ;
        RECT 48.630 242.150 48.780 249.700 ;
        RECT 49.230 242.150 49.380 249.700 ;
        RECT 49.830 242.150 49.980 249.700 ;
        RECT 54.230 249.200 55.230 249.700 ;
        RECT 50.880 249.050 58.580 249.200 ;
        RECT 54.230 248.600 55.230 249.050 ;
        RECT 50.880 248.450 58.580 248.600 ;
        RECT 54.230 248.000 55.230 248.450 ;
        RECT 50.880 247.850 58.580 248.000 ;
        RECT 54.230 247.400 55.230 247.850 ;
        RECT 50.880 247.250 58.580 247.400 ;
        RECT 54.230 246.800 55.230 247.250 ;
        RECT 50.880 246.650 58.580 246.800 ;
        RECT 54.230 246.200 55.230 246.650 ;
        RECT 50.880 246.050 58.580 246.200 ;
        RECT 54.230 245.600 55.230 246.050 ;
        RECT 50.880 245.450 58.580 245.600 ;
        RECT 54.230 245.000 55.230 245.450 ;
        RECT 50.880 244.850 58.580 245.000 ;
        RECT 54.230 244.400 55.230 244.850 ;
        RECT 50.880 244.250 58.580 244.400 ;
        RECT 54.230 243.800 55.230 244.250 ;
        RECT 50.880 243.650 58.580 243.800 ;
        RECT 54.230 243.200 55.230 243.650 ;
        RECT 50.880 243.050 58.580 243.200 ;
        RECT 54.230 242.600 55.230 243.050 ;
        RECT 50.880 242.450 58.580 242.600 ;
        RECT 54.230 242.000 55.230 242.450 ;
        RECT 59.480 242.150 59.630 249.700 ;
        RECT 60.080 242.150 60.230 249.700 ;
        RECT 60.680 242.150 60.830 249.700 ;
        RECT 61.280 242.150 61.430 249.700 ;
        RECT 61.880 242.150 62.030 249.700 ;
        RECT 62.480 242.150 62.630 249.700 ;
        RECT 62.780 249.550 63.930 249.700 ;
        RECT 64.580 249.550 64.880 250.450 ;
        RECT 65.530 250.300 66.680 250.450 ;
        RECT 66.830 250.300 66.980 257.850 ;
        RECT 67.430 250.300 67.580 257.850 ;
        RECT 68.030 250.300 68.180 257.850 ;
        RECT 68.630 250.300 68.780 257.850 ;
        RECT 69.230 250.300 69.380 257.850 ;
        RECT 69.830 250.300 69.980 257.850 ;
        RECT 74.230 257.550 75.230 258.000 ;
        RECT 70.880 257.400 78.580 257.550 ;
        RECT 74.230 256.950 75.230 257.400 ;
        RECT 70.880 256.800 78.580 256.950 ;
        RECT 74.230 256.350 75.230 256.800 ;
        RECT 70.880 256.200 78.580 256.350 ;
        RECT 74.230 255.750 75.230 256.200 ;
        RECT 70.880 255.600 78.580 255.750 ;
        RECT 74.230 255.150 75.230 255.600 ;
        RECT 70.880 255.000 78.580 255.150 ;
        RECT 74.230 254.550 75.230 255.000 ;
        RECT 70.880 254.400 78.580 254.550 ;
        RECT 74.230 253.950 75.230 254.400 ;
        RECT 70.880 253.800 78.580 253.950 ;
        RECT 74.230 253.350 75.230 253.800 ;
        RECT 70.880 253.200 78.580 253.350 ;
        RECT 74.230 252.750 75.230 253.200 ;
        RECT 70.880 252.600 78.580 252.750 ;
        RECT 74.230 252.150 75.230 252.600 ;
        RECT 70.880 252.000 78.580 252.150 ;
        RECT 74.230 251.550 75.230 252.000 ;
        RECT 70.880 251.400 78.580 251.550 ;
        RECT 74.230 250.950 75.230 251.400 ;
        RECT 70.880 250.800 78.580 250.950 ;
        RECT 74.230 250.300 75.230 250.800 ;
        RECT 79.480 250.300 79.630 257.850 ;
        RECT 80.080 250.300 80.230 257.850 ;
        RECT 80.680 250.300 80.830 257.850 ;
        RECT 81.280 250.300 81.430 257.850 ;
        RECT 81.880 250.300 82.030 257.850 ;
        RECT 82.480 250.300 82.630 257.850 ;
        RECT 82.780 253.200 83.530 255.000 ;
        RECT 85.930 253.200 86.680 255.000 ;
        RECT 82.780 250.450 86.680 253.200 ;
        RECT 82.780 250.300 83.930 250.450 ;
        RECT 65.530 249.700 83.930 250.300 ;
        RECT 65.530 249.550 66.680 249.700 ;
        RECT 62.780 246.800 66.680 249.550 ;
        RECT 62.780 245.050 63.530 246.800 ;
        RECT 65.930 245.050 66.680 246.800 ;
        RECT 66.830 242.150 66.980 249.700 ;
        RECT 67.430 242.150 67.580 249.700 ;
        RECT 68.030 242.150 68.180 249.700 ;
        RECT 68.630 242.150 68.780 249.700 ;
        RECT 69.230 242.150 69.380 249.700 ;
        RECT 69.830 242.150 69.980 249.700 ;
        RECT 74.230 249.200 75.230 249.700 ;
        RECT 70.880 249.050 78.580 249.200 ;
        RECT 74.230 248.600 75.230 249.050 ;
        RECT 70.880 248.450 78.580 248.600 ;
        RECT 74.230 248.000 75.230 248.450 ;
        RECT 70.880 247.850 78.580 248.000 ;
        RECT 74.230 247.400 75.230 247.850 ;
        RECT 70.880 247.250 78.580 247.400 ;
        RECT 74.230 246.800 75.230 247.250 ;
        RECT 70.880 246.650 78.580 246.800 ;
        RECT 74.230 246.200 75.230 246.650 ;
        RECT 70.880 246.050 78.580 246.200 ;
        RECT 74.230 245.600 75.230 246.050 ;
        RECT 70.880 245.450 78.580 245.600 ;
        RECT 74.230 245.000 75.230 245.450 ;
        RECT 70.880 244.850 78.580 245.000 ;
        RECT 74.230 244.400 75.230 244.850 ;
        RECT 70.880 244.250 78.580 244.400 ;
        RECT 74.230 243.800 75.230 244.250 ;
        RECT 70.880 243.650 78.580 243.800 ;
        RECT 74.230 243.200 75.230 243.650 ;
        RECT 70.880 243.050 78.580 243.200 ;
        RECT 74.230 242.600 75.230 243.050 ;
        RECT 70.880 242.450 78.580 242.600 ;
        RECT 74.230 242.000 75.230 242.450 ;
        RECT 79.480 242.150 79.630 249.700 ;
        RECT 80.080 242.150 80.230 249.700 ;
        RECT 80.680 242.150 80.830 249.700 ;
        RECT 81.280 242.150 81.430 249.700 ;
        RECT 81.880 242.150 82.030 249.700 ;
        RECT 82.480 242.150 82.630 249.700 ;
        RECT 82.780 249.550 83.930 249.700 ;
        RECT 84.580 249.550 84.880 250.450 ;
        RECT 85.530 250.300 86.680 250.450 ;
        RECT 86.830 250.300 86.980 257.850 ;
        RECT 87.430 250.300 87.580 257.850 ;
        RECT 88.030 250.300 88.180 257.850 ;
        RECT 88.630 250.300 88.780 257.850 ;
        RECT 89.230 250.300 89.380 257.850 ;
        RECT 89.830 250.300 89.980 257.850 ;
        RECT 94.230 257.550 95.230 258.000 ;
        RECT 90.880 257.400 98.580 257.550 ;
        RECT 94.230 256.950 95.230 257.400 ;
        RECT 90.880 256.800 98.580 256.950 ;
        RECT 94.230 256.350 95.230 256.800 ;
        RECT 90.880 256.200 98.580 256.350 ;
        RECT 94.230 255.750 95.230 256.200 ;
        RECT 90.880 255.600 98.580 255.750 ;
        RECT 94.230 255.150 95.230 255.600 ;
        RECT 90.880 255.000 98.580 255.150 ;
        RECT 94.230 254.550 95.230 255.000 ;
        RECT 90.880 254.400 98.580 254.550 ;
        RECT 94.230 253.950 95.230 254.400 ;
        RECT 90.880 253.800 98.580 253.950 ;
        RECT 94.230 253.350 95.230 253.800 ;
        RECT 90.880 253.200 98.580 253.350 ;
        RECT 94.230 252.750 95.230 253.200 ;
        RECT 90.880 252.600 98.580 252.750 ;
        RECT 94.230 252.150 95.230 252.600 ;
        RECT 90.880 252.000 98.580 252.150 ;
        RECT 94.230 251.550 95.230 252.000 ;
        RECT 90.880 251.400 98.580 251.550 ;
        RECT 94.230 250.950 95.230 251.400 ;
        RECT 90.880 250.800 98.580 250.950 ;
        RECT 94.230 250.300 95.230 250.800 ;
        RECT 99.480 250.300 99.630 257.850 ;
        RECT 100.080 250.300 100.230 257.850 ;
        RECT 100.680 250.300 100.830 257.850 ;
        RECT 101.280 250.300 101.430 257.850 ;
        RECT 101.880 250.300 102.030 257.850 ;
        RECT 102.480 250.300 102.630 257.850 ;
        RECT 102.780 253.200 103.530 255.000 ;
        RECT 102.780 250.915 104.730 253.200 ;
        RECT 102.780 250.450 111.850 250.915 ;
        RECT 102.780 250.300 103.930 250.450 ;
        RECT 85.530 249.700 103.930 250.300 ;
        RECT 85.530 249.550 86.680 249.700 ;
        RECT 82.780 246.800 86.680 249.550 ;
        RECT 82.780 245.050 83.530 246.800 ;
        RECT 85.930 245.050 86.680 246.800 ;
        RECT 86.830 242.150 86.980 249.700 ;
        RECT 87.430 242.150 87.580 249.700 ;
        RECT 88.030 242.150 88.180 249.700 ;
        RECT 88.630 242.150 88.780 249.700 ;
        RECT 89.230 242.150 89.380 249.700 ;
        RECT 89.830 242.150 89.980 249.700 ;
        RECT 94.230 249.200 95.230 249.700 ;
        RECT 90.880 249.050 98.580 249.200 ;
        RECT 94.230 248.600 95.230 249.050 ;
        RECT 90.880 248.450 98.580 248.600 ;
        RECT 94.230 248.000 95.230 248.450 ;
        RECT 90.880 247.850 98.580 248.000 ;
        RECT 94.230 247.400 95.230 247.850 ;
        RECT 90.880 247.250 98.580 247.400 ;
        RECT 94.230 246.800 95.230 247.250 ;
        RECT 90.880 246.650 98.580 246.800 ;
        RECT 94.230 246.200 95.230 246.650 ;
        RECT 90.880 246.050 98.580 246.200 ;
        RECT 94.230 245.600 95.230 246.050 ;
        RECT 90.880 245.450 98.580 245.600 ;
        RECT 94.230 245.000 95.230 245.450 ;
        RECT 90.880 244.850 98.580 245.000 ;
        RECT 94.230 244.400 95.230 244.850 ;
        RECT 90.880 244.250 98.580 244.400 ;
        RECT 94.230 243.800 95.230 244.250 ;
        RECT 90.880 243.650 98.580 243.800 ;
        RECT 94.230 243.200 95.230 243.650 ;
        RECT 90.880 243.050 98.580 243.200 ;
        RECT 94.230 242.600 95.230 243.050 ;
        RECT 90.880 242.450 98.580 242.600 ;
        RECT 94.230 242.000 95.230 242.450 ;
        RECT 99.480 242.150 99.630 249.700 ;
        RECT 100.080 242.150 100.230 249.700 ;
        RECT 100.680 242.150 100.830 249.700 ;
        RECT 101.280 242.150 101.430 249.700 ;
        RECT 101.880 242.150 102.030 249.700 ;
        RECT 102.480 242.150 102.630 249.700 ;
        RECT 102.780 249.550 103.930 249.700 ;
        RECT 104.580 249.640 111.850 250.450 ;
        RECT 104.580 249.550 104.730 249.640 ;
        RECT 102.780 246.800 104.730 249.550 ;
        RECT 102.780 245.050 103.530 246.800 ;
        RECT 10.880 241.850 18.580 242.000 ;
        RECT 30.880 241.850 38.580 242.000 ;
        RECT 50.880 241.850 58.580 242.000 ;
        RECT 70.880 241.850 78.580 242.000 ;
        RECT 90.880 241.850 98.580 242.000 ;
        RECT 14.230 241.200 15.230 241.850 ;
        RECT 34.230 241.200 35.230 241.850 ;
        RECT 54.230 241.200 55.230 241.850 ;
        RECT 74.230 241.200 75.230 241.850 ;
        RECT 94.230 241.200 95.230 241.850 ;
        RECT 11.530 238.800 17.930 241.200 ;
        RECT 31.530 238.800 37.930 241.200 ;
        RECT 51.530 238.800 57.930 241.200 ;
        RECT 71.530 238.800 77.930 241.200 ;
        RECT 91.530 238.800 97.930 241.200 ;
        RECT 14.230 238.150 15.230 238.800 ;
        RECT 34.230 238.150 35.230 238.800 ;
        RECT 54.230 238.150 55.230 238.800 ;
        RECT 74.230 238.150 75.230 238.800 ;
        RECT 94.230 238.150 95.230 238.800 ;
        RECT 10.880 238.000 18.580 238.150 ;
        RECT 30.880 238.000 38.580 238.150 ;
        RECT 50.880 238.000 58.580 238.150 ;
        RECT 70.880 238.000 78.580 238.150 ;
        RECT 90.880 238.000 98.580 238.150 ;
        RECT 5.930 233.200 6.680 235.000 ;
        RECT 4.730 230.450 6.680 233.200 ;
        RECT 4.730 229.550 4.880 230.450 ;
        RECT 5.530 230.300 6.680 230.450 ;
        RECT 6.830 230.300 6.980 237.850 ;
        RECT 7.430 230.300 7.580 237.850 ;
        RECT 8.030 230.300 8.180 237.850 ;
        RECT 8.630 230.300 8.780 237.850 ;
        RECT 9.230 230.300 9.380 237.850 ;
        RECT 9.830 230.300 9.980 237.850 ;
        RECT 14.230 237.550 15.230 238.000 ;
        RECT 10.880 237.400 18.580 237.550 ;
        RECT 14.230 236.950 15.230 237.400 ;
        RECT 10.880 236.800 18.580 236.950 ;
        RECT 14.230 236.350 15.230 236.800 ;
        RECT 10.880 236.200 18.580 236.350 ;
        RECT 14.230 235.750 15.230 236.200 ;
        RECT 10.880 235.600 18.580 235.750 ;
        RECT 14.230 235.150 15.230 235.600 ;
        RECT 10.880 235.000 18.580 235.150 ;
        RECT 14.230 234.550 15.230 235.000 ;
        RECT 10.880 234.400 18.580 234.550 ;
        RECT 14.230 233.950 15.230 234.400 ;
        RECT 10.880 233.800 18.580 233.950 ;
        RECT 14.230 233.350 15.230 233.800 ;
        RECT 10.880 233.200 18.580 233.350 ;
        RECT 14.230 232.750 15.230 233.200 ;
        RECT 10.880 232.600 18.580 232.750 ;
        RECT 14.230 232.150 15.230 232.600 ;
        RECT 10.880 232.000 18.580 232.150 ;
        RECT 14.230 231.550 15.230 232.000 ;
        RECT 10.880 231.400 18.580 231.550 ;
        RECT 14.230 230.950 15.230 231.400 ;
        RECT 10.880 230.800 18.580 230.950 ;
        RECT 14.230 230.300 15.230 230.800 ;
        RECT 19.480 230.300 19.630 237.850 ;
        RECT 20.080 230.300 20.230 237.850 ;
        RECT 20.680 230.300 20.830 237.850 ;
        RECT 21.280 230.300 21.430 237.850 ;
        RECT 21.880 230.300 22.030 237.850 ;
        RECT 22.480 230.300 22.630 237.850 ;
        RECT 22.780 233.200 23.530 235.000 ;
        RECT 25.930 233.200 26.680 235.000 ;
        RECT 22.780 230.450 26.680 233.200 ;
        RECT 22.780 230.300 23.930 230.450 ;
        RECT 5.530 229.700 23.930 230.300 ;
        RECT 5.530 229.550 6.680 229.700 ;
        RECT 4.730 226.800 6.680 229.550 ;
        RECT 5.930 225.050 6.680 226.800 ;
        RECT 6.830 222.150 6.980 229.700 ;
        RECT 7.430 222.150 7.580 229.700 ;
        RECT 8.030 222.150 8.180 229.700 ;
        RECT 8.630 222.150 8.780 229.700 ;
        RECT 9.230 222.150 9.380 229.700 ;
        RECT 9.830 222.150 9.980 229.700 ;
        RECT 14.230 229.200 15.230 229.700 ;
        RECT 10.880 229.050 18.580 229.200 ;
        RECT 14.230 228.600 15.230 229.050 ;
        RECT 10.880 228.450 18.580 228.600 ;
        RECT 14.230 228.000 15.230 228.450 ;
        RECT 10.880 227.850 18.580 228.000 ;
        RECT 14.230 227.400 15.230 227.850 ;
        RECT 10.880 227.250 18.580 227.400 ;
        RECT 14.230 226.800 15.230 227.250 ;
        RECT 10.880 226.650 18.580 226.800 ;
        RECT 14.230 226.200 15.230 226.650 ;
        RECT 10.880 226.050 18.580 226.200 ;
        RECT 14.230 225.600 15.230 226.050 ;
        RECT 10.880 225.450 18.580 225.600 ;
        RECT 14.230 225.000 15.230 225.450 ;
        RECT 10.880 224.850 18.580 225.000 ;
        RECT 14.230 224.400 15.230 224.850 ;
        RECT 10.880 224.250 18.580 224.400 ;
        RECT 14.230 223.800 15.230 224.250 ;
        RECT 10.880 223.650 18.580 223.800 ;
        RECT 14.230 223.200 15.230 223.650 ;
        RECT 10.880 223.050 18.580 223.200 ;
        RECT 14.230 222.600 15.230 223.050 ;
        RECT 10.880 222.450 18.580 222.600 ;
        RECT 14.230 222.000 15.230 222.450 ;
        RECT 19.480 222.150 19.630 229.700 ;
        RECT 20.080 222.150 20.230 229.700 ;
        RECT 20.680 222.150 20.830 229.700 ;
        RECT 21.280 222.150 21.430 229.700 ;
        RECT 21.880 222.150 22.030 229.700 ;
        RECT 22.480 222.150 22.630 229.700 ;
        RECT 22.780 229.550 23.930 229.700 ;
        RECT 24.580 229.550 24.880 230.450 ;
        RECT 25.530 230.300 26.680 230.450 ;
        RECT 26.830 230.300 26.980 237.850 ;
        RECT 27.430 230.300 27.580 237.850 ;
        RECT 28.030 230.300 28.180 237.850 ;
        RECT 28.630 230.300 28.780 237.850 ;
        RECT 29.230 230.300 29.380 237.850 ;
        RECT 29.830 230.300 29.980 237.850 ;
        RECT 34.230 237.550 35.230 238.000 ;
        RECT 30.880 237.400 38.580 237.550 ;
        RECT 34.230 236.950 35.230 237.400 ;
        RECT 30.880 236.800 38.580 236.950 ;
        RECT 34.230 236.350 35.230 236.800 ;
        RECT 30.880 236.200 38.580 236.350 ;
        RECT 34.230 235.750 35.230 236.200 ;
        RECT 30.880 235.600 38.580 235.750 ;
        RECT 34.230 235.150 35.230 235.600 ;
        RECT 30.880 235.000 38.580 235.150 ;
        RECT 34.230 234.550 35.230 235.000 ;
        RECT 30.880 234.400 38.580 234.550 ;
        RECT 34.230 233.950 35.230 234.400 ;
        RECT 30.880 233.800 38.580 233.950 ;
        RECT 34.230 233.350 35.230 233.800 ;
        RECT 30.880 233.200 38.580 233.350 ;
        RECT 34.230 232.750 35.230 233.200 ;
        RECT 30.880 232.600 38.580 232.750 ;
        RECT 34.230 232.150 35.230 232.600 ;
        RECT 30.880 232.000 38.580 232.150 ;
        RECT 34.230 231.550 35.230 232.000 ;
        RECT 30.880 231.400 38.580 231.550 ;
        RECT 34.230 230.950 35.230 231.400 ;
        RECT 30.880 230.800 38.580 230.950 ;
        RECT 34.230 230.300 35.230 230.800 ;
        RECT 39.480 230.300 39.630 237.850 ;
        RECT 40.080 230.300 40.230 237.850 ;
        RECT 40.680 230.300 40.830 237.850 ;
        RECT 41.280 230.300 41.430 237.850 ;
        RECT 41.880 230.300 42.030 237.850 ;
        RECT 42.480 230.300 42.630 237.850 ;
        RECT 42.780 233.200 43.530 235.000 ;
        RECT 45.930 233.200 46.680 235.000 ;
        RECT 42.780 230.450 46.680 233.200 ;
        RECT 42.780 230.300 43.930 230.450 ;
        RECT 25.530 229.700 43.930 230.300 ;
        RECT 25.530 229.550 26.680 229.700 ;
        RECT 22.780 226.800 26.680 229.550 ;
        RECT 22.780 225.050 23.530 226.800 ;
        RECT 25.930 225.050 26.680 226.800 ;
        RECT 26.830 222.150 26.980 229.700 ;
        RECT 27.430 222.150 27.580 229.700 ;
        RECT 28.030 222.150 28.180 229.700 ;
        RECT 28.630 222.150 28.780 229.700 ;
        RECT 29.230 222.150 29.380 229.700 ;
        RECT 29.830 222.150 29.980 229.700 ;
        RECT 34.230 229.200 35.230 229.700 ;
        RECT 30.880 229.050 38.580 229.200 ;
        RECT 34.230 228.600 35.230 229.050 ;
        RECT 30.880 228.450 38.580 228.600 ;
        RECT 34.230 228.000 35.230 228.450 ;
        RECT 30.880 227.850 38.580 228.000 ;
        RECT 34.230 227.400 35.230 227.850 ;
        RECT 30.880 227.250 38.580 227.400 ;
        RECT 34.230 226.800 35.230 227.250 ;
        RECT 30.880 226.650 38.580 226.800 ;
        RECT 34.230 226.200 35.230 226.650 ;
        RECT 30.880 226.050 38.580 226.200 ;
        RECT 34.230 225.600 35.230 226.050 ;
        RECT 30.880 225.450 38.580 225.600 ;
        RECT 34.230 225.000 35.230 225.450 ;
        RECT 30.880 224.850 38.580 225.000 ;
        RECT 34.230 224.400 35.230 224.850 ;
        RECT 30.880 224.250 38.580 224.400 ;
        RECT 34.230 223.800 35.230 224.250 ;
        RECT 30.880 223.650 38.580 223.800 ;
        RECT 34.230 223.200 35.230 223.650 ;
        RECT 30.880 223.050 38.580 223.200 ;
        RECT 34.230 222.600 35.230 223.050 ;
        RECT 30.880 222.450 38.580 222.600 ;
        RECT 34.230 222.000 35.230 222.450 ;
        RECT 39.480 222.150 39.630 229.700 ;
        RECT 40.080 222.150 40.230 229.700 ;
        RECT 40.680 222.150 40.830 229.700 ;
        RECT 41.280 222.150 41.430 229.700 ;
        RECT 41.880 222.150 42.030 229.700 ;
        RECT 42.480 222.150 42.630 229.700 ;
        RECT 42.780 229.550 43.930 229.700 ;
        RECT 44.580 229.550 44.880 230.450 ;
        RECT 45.530 230.300 46.680 230.450 ;
        RECT 46.830 230.300 46.980 237.850 ;
        RECT 47.430 230.300 47.580 237.850 ;
        RECT 48.030 230.300 48.180 237.850 ;
        RECT 48.630 230.300 48.780 237.850 ;
        RECT 49.230 230.300 49.380 237.850 ;
        RECT 49.830 230.300 49.980 237.850 ;
        RECT 54.230 237.550 55.230 238.000 ;
        RECT 50.880 237.400 58.580 237.550 ;
        RECT 54.230 236.950 55.230 237.400 ;
        RECT 50.880 236.800 58.580 236.950 ;
        RECT 54.230 236.350 55.230 236.800 ;
        RECT 50.880 236.200 58.580 236.350 ;
        RECT 54.230 235.750 55.230 236.200 ;
        RECT 50.880 235.600 58.580 235.750 ;
        RECT 54.230 235.150 55.230 235.600 ;
        RECT 50.880 235.000 58.580 235.150 ;
        RECT 54.230 234.550 55.230 235.000 ;
        RECT 50.880 234.400 58.580 234.550 ;
        RECT 54.230 233.950 55.230 234.400 ;
        RECT 50.880 233.800 58.580 233.950 ;
        RECT 54.230 233.350 55.230 233.800 ;
        RECT 50.880 233.200 58.580 233.350 ;
        RECT 54.230 232.750 55.230 233.200 ;
        RECT 50.880 232.600 58.580 232.750 ;
        RECT 54.230 232.150 55.230 232.600 ;
        RECT 50.880 232.000 58.580 232.150 ;
        RECT 54.230 231.550 55.230 232.000 ;
        RECT 50.880 231.400 58.580 231.550 ;
        RECT 54.230 230.950 55.230 231.400 ;
        RECT 50.880 230.800 58.580 230.950 ;
        RECT 54.230 230.300 55.230 230.800 ;
        RECT 59.480 230.300 59.630 237.850 ;
        RECT 60.080 230.300 60.230 237.850 ;
        RECT 60.680 230.300 60.830 237.850 ;
        RECT 61.280 230.300 61.430 237.850 ;
        RECT 61.880 230.300 62.030 237.850 ;
        RECT 62.480 230.300 62.630 237.850 ;
        RECT 62.780 233.200 63.530 235.000 ;
        RECT 65.930 233.200 66.680 235.000 ;
        RECT 62.780 230.450 66.680 233.200 ;
        RECT 62.780 230.300 63.930 230.450 ;
        RECT 45.530 229.700 63.930 230.300 ;
        RECT 45.530 229.550 46.680 229.700 ;
        RECT 42.780 226.800 46.680 229.550 ;
        RECT 42.780 225.050 43.530 226.800 ;
        RECT 45.930 225.050 46.680 226.800 ;
        RECT 46.830 222.150 46.980 229.700 ;
        RECT 47.430 222.150 47.580 229.700 ;
        RECT 48.030 222.150 48.180 229.700 ;
        RECT 48.630 222.150 48.780 229.700 ;
        RECT 49.230 222.150 49.380 229.700 ;
        RECT 49.830 222.150 49.980 229.700 ;
        RECT 54.230 229.200 55.230 229.700 ;
        RECT 50.880 229.050 58.580 229.200 ;
        RECT 54.230 228.600 55.230 229.050 ;
        RECT 50.880 228.450 58.580 228.600 ;
        RECT 54.230 228.000 55.230 228.450 ;
        RECT 50.880 227.850 58.580 228.000 ;
        RECT 54.230 227.400 55.230 227.850 ;
        RECT 50.880 227.250 58.580 227.400 ;
        RECT 54.230 226.800 55.230 227.250 ;
        RECT 50.880 226.650 58.580 226.800 ;
        RECT 54.230 226.200 55.230 226.650 ;
        RECT 50.880 226.050 58.580 226.200 ;
        RECT 54.230 225.600 55.230 226.050 ;
        RECT 50.880 225.450 58.580 225.600 ;
        RECT 54.230 225.000 55.230 225.450 ;
        RECT 50.880 224.850 58.580 225.000 ;
        RECT 54.230 224.400 55.230 224.850 ;
        RECT 50.880 224.250 58.580 224.400 ;
        RECT 54.230 223.800 55.230 224.250 ;
        RECT 50.880 223.650 58.580 223.800 ;
        RECT 54.230 223.200 55.230 223.650 ;
        RECT 50.880 223.050 58.580 223.200 ;
        RECT 54.230 222.600 55.230 223.050 ;
        RECT 50.880 222.450 58.580 222.600 ;
        RECT 54.230 222.000 55.230 222.450 ;
        RECT 59.480 222.150 59.630 229.700 ;
        RECT 60.080 222.150 60.230 229.700 ;
        RECT 60.680 222.150 60.830 229.700 ;
        RECT 61.280 222.150 61.430 229.700 ;
        RECT 61.880 222.150 62.030 229.700 ;
        RECT 62.480 222.150 62.630 229.700 ;
        RECT 62.780 229.550 63.930 229.700 ;
        RECT 64.580 229.550 64.880 230.450 ;
        RECT 65.530 230.300 66.680 230.450 ;
        RECT 66.830 230.300 66.980 237.850 ;
        RECT 67.430 230.300 67.580 237.850 ;
        RECT 68.030 230.300 68.180 237.850 ;
        RECT 68.630 230.300 68.780 237.850 ;
        RECT 69.230 230.300 69.380 237.850 ;
        RECT 69.830 230.300 69.980 237.850 ;
        RECT 74.230 237.550 75.230 238.000 ;
        RECT 70.880 237.400 78.580 237.550 ;
        RECT 74.230 236.950 75.230 237.400 ;
        RECT 70.880 236.800 78.580 236.950 ;
        RECT 74.230 236.350 75.230 236.800 ;
        RECT 70.880 236.200 78.580 236.350 ;
        RECT 74.230 235.750 75.230 236.200 ;
        RECT 70.880 235.600 78.580 235.750 ;
        RECT 74.230 235.150 75.230 235.600 ;
        RECT 70.880 235.000 78.580 235.150 ;
        RECT 74.230 234.550 75.230 235.000 ;
        RECT 70.880 234.400 78.580 234.550 ;
        RECT 74.230 233.950 75.230 234.400 ;
        RECT 70.880 233.800 78.580 233.950 ;
        RECT 74.230 233.350 75.230 233.800 ;
        RECT 70.880 233.200 78.580 233.350 ;
        RECT 74.230 232.750 75.230 233.200 ;
        RECT 70.880 232.600 78.580 232.750 ;
        RECT 74.230 232.150 75.230 232.600 ;
        RECT 70.880 232.000 78.580 232.150 ;
        RECT 74.230 231.550 75.230 232.000 ;
        RECT 70.880 231.400 78.580 231.550 ;
        RECT 74.230 230.950 75.230 231.400 ;
        RECT 70.880 230.800 78.580 230.950 ;
        RECT 74.230 230.300 75.230 230.800 ;
        RECT 79.480 230.300 79.630 237.850 ;
        RECT 80.080 230.300 80.230 237.850 ;
        RECT 80.680 230.300 80.830 237.850 ;
        RECT 81.280 230.300 81.430 237.850 ;
        RECT 81.880 230.300 82.030 237.850 ;
        RECT 82.480 230.300 82.630 237.850 ;
        RECT 82.780 233.200 83.530 235.000 ;
        RECT 85.930 233.200 86.680 235.000 ;
        RECT 82.780 230.450 86.680 233.200 ;
        RECT 82.780 230.300 83.930 230.450 ;
        RECT 65.530 229.700 83.930 230.300 ;
        RECT 65.530 229.550 66.680 229.700 ;
        RECT 62.780 226.800 66.680 229.550 ;
        RECT 62.780 225.050 63.530 226.800 ;
        RECT 65.930 225.050 66.680 226.800 ;
        RECT 66.830 222.150 66.980 229.700 ;
        RECT 67.430 222.150 67.580 229.700 ;
        RECT 68.030 222.150 68.180 229.700 ;
        RECT 68.630 222.150 68.780 229.700 ;
        RECT 69.230 222.150 69.380 229.700 ;
        RECT 69.830 222.150 69.980 229.700 ;
        RECT 74.230 229.200 75.230 229.700 ;
        RECT 70.880 229.050 78.580 229.200 ;
        RECT 74.230 228.600 75.230 229.050 ;
        RECT 70.880 228.450 78.580 228.600 ;
        RECT 74.230 228.000 75.230 228.450 ;
        RECT 70.880 227.850 78.580 228.000 ;
        RECT 74.230 227.400 75.230 227.850 ;
        RECT 70.880 227.250 78.580 227.400 ;
        RECT 74.230 226.800 75.230 227.250 ;
        RECT 70.880 226.650 78.580 226.800 ;
        RECT 74.230 226.200 75.230 226.650 ;
        RECT 70.880 226.050 78.580 226.200 ;
        RECT 74.230 225.600 75.230 226.050 ;
        RECT 70.880 225.450 78.580 225.600 ;
        RECT 74.230 225.000 75.230 225.450 ;
        RECT 70.880 224.850 78.580 225.000 ;
        RECT 74.230 224.400 75.230 224.850 ;
        RECT 70.880 224.250 78.580 224.400 ;
        RECT 74.230 223.800 75.230 224.250 ;
        RECT 70.880 223.650 78.580 223.800 ;
        RECT 74.230 223.200 75.230 223.650 ;
        RECT 70.880 223.050 78.580 223.200 ;
        RECT 74.230 222.600 75.230 223.050 ;
        RECT 70.880 222.450 78.580 222.600 ;
        RECT 74.230 222.000 75.230 222.450 ;
        RECT 79.480 222.150 79.630 229.700 ;
        RECT 80.080 222.150 80.230 229.700 ;
        RECT 80.680 222.150 80.830 229.700 ;
        RECT 81.280 222.150 81.430 229.700 ;
        RECT 81.880 222.150 82.030 229.700 ;
        RECT 82.480 222.150 82.630 229.700 ;
        RECT 82.780 229.550 83.930 229.700 ;
        RECT 84.580 229.550 84.880 230.450 ;
        RECT 85.530 230.300 86.680 230.450 ;
        RECT 86.830 230.300 86.980 237.850 ;
        RECT 87.430 230.300 87.580 237.850 ;
        RECT 88.030 230.300 88.180 237.850 ;
        RECT 88.630 230.300 88.780 237.850 ;
        RECT 89.230 230.300 89.380 237.850 ;
        RECT 89.830 230.300 89.980 237.850 ;
        RECT 94.230 237.550 95.230 238.000 ;
        RECT 90.880 237.400 98.580 237.550 ;
        RECT 94.230 236.950 95.230 237.400 ;
        RECT 90.880 236.800 98.580 236.950 ;
        RECT 94.230 236.350 95.230 236.800 ;
        RECT 90.880 236.200 98.580 236.350 ;
        RECT 94.230 235.750 95.230 236.200 ;
        RECT 90.880 235.600 98.580 235.750 ;
        RECT 94.230 235.150 95.230 235.600 ;
        RECT 90.880 235.000 98.580 235.150 ;
        RECT 94.230 234.550 95.230 235.000 ;
        RECT 90.880 234.400 98.580 234.550 ;
        RECT 94.230 233.950 95.230 234.400 ;
        RECT 90.880 233.800 98.580 233.950 ;
        RECT 94.230 233.350 95.230 233.800 ;
        RECT 90.880 233.200 98.580 233.350 ;
        RECT 94.230 232.750 95.230 233.200 ;
        RECT 90.880 232.600 98.580 232.750 ;
        RECT 94.230 232.150 95.230 232.600 ;
        RECT 90.880 232.000 98.580 232.150 ;
        RECT 94.230 231.550 95.230 232.000 ;
        RECT 90.880 231.400 98.580 231.550 ;
        RECT 94.230 230.950 95.230 231.400 ;
        RECT 90.880 230.800 98.580 230.950 ;
        RECT 94.230 230.300 95.230 230.800 ;
        RECT 99.480 230.300 99.630 237.850 ;
        RECT 100.080 230.300 100.230 237.850 ;
        RECT 100.680 230.300 100.830 237.850 ;
        RECT 101.280 230.300 101.430 237.850 ;
        RECT 101.880 230.300 102.030 237.850 ;
        RECT 102.480 230.300 102.630 237.850 ;
        RECT 102.780 233.200 103.530 235.000 ;
        RECT 102.780 230.450 104.730 233.200 ;
        RECT 102.780 230.300 103.930 230.450 ;
        RECT 85.530 229.700 103.930 230.300 ;
        RECT 85.530 229.550 86.680 229.700 ;
        RECT 82.780 226.800 86.680 229.550 ;
        RECT 82.780 225.050 83.530 226.800 ;
        RECT 85.930 225.050 86.680 226.800 ;
        RECT 86.830 222.150 86.980 229.700 ;
        RECT 87.430 222.150 87.580 229.700 ;
        RECT 88.030 222.150 88.180 229.700 ;
        RECT 88.630 222.150 88.780 229.700 ;
        RECT 89.230 222.150 89.380 229.700 ;
        RECT 89.830 222.150 89.980 229.700 ;
        RECT 94.230 229.200 95.230 229.700 ;
        RECT 90.880 229.050 98.580 229.200 ;
        RECT 94.230 228.600 95.230 229.050 ;
        RECT 90.880 228.450 98.580 228.600 ;
        RECT 94.230 228.000 95.230 228.450 ;
        RECT 90.880 227.850 98.580 228.000 ;
        RECT 94.230 227.400 95.230 227.850 ;
        RECT 90.880 227.250 98.580 227.400 ;
        RECT 94.230 226.800 95.230 227.250 ;
        RECT 90.880 226.650 98.580 226.800 ;
        RECT 94.230 226.200 95.230 226.650 ;
        RECT 90.880 226.050 98.580 226.200 ;
        RECT 94.230 225.600 95.230 226.050 ;
        RECT 90.880 225.450 98.580 225.600 ;
        RECT 94.230 225.000 95.230 225.450 ;
        RECT 90.880 224.850 98.580 225.000 ;
        RECT 94.230 224.400 95.230 224.850 ;
        RECT 90.880 224.250 98.580 224.400 ;
        RECT 94.230 223.800 95.230 224.250 ;
        RECT 90.880 223.650 98.580 223.800 ;
        RECT 94.230 223.200 95.230 223.650 ;
        RECT 90.880 223.050 98.580 223.200 ;
        RECT 94.230 222.600 95.230 223.050 ;
        RECT 90.880 222.450 98.580 222.600 ;
        RECT 94.230 222.000 95.230 222.450 ;
        RECT 99.480 222.150 99.630 229.700 ;
        RECT 100.080 222.150 100.230 229.700 ;
        RECT 100.680 222.150 100.830 229.700 ;
        RECT 101.280 222.150 101.430 229.700 ;
        RECT 101.880 222.150 102.030 229.700 ;
        RECT 102.480 222.150 102.630 229.700 ;
        RECT 102.780 229.550 103.930 229.700 ;
        RECT 104.580 229.625 104.730 230.450 ;
        RECT 104.580 229.550 111.850 229.625 ;
        RECT 102.780 228.350 111.850 229.550 ;
        RECT 102.780 226.800 104.730 228.350 ;
        RECT 102.780 225.050 103.530 226.800 ;
        RECT 10.880 221.850 18.580 222.000 ;
        RECT 30.880 221.850 38.580 222.000 ;
        RECT 50.880 221.850 58.580 222.000 ;
        RECT 70.880 221.850 78.580 222.000 ;
        RECT 90.880 221.850 98.580 222.000 ;
        RECT 14.230 221.200 15.230 221.850 ;
        RECT 34.230 221.200 35.230 221.850 ;
        RECT 54.230 221.200 55.230 221.850 ;
        RECT 74.230 221.200 75.230 221.850 ;
        RECT 94.230 221.200 95.230 221.850 ;
        RECT 11.530 220.000 17.930 221.200 ;
        RECT 31.530 220.000 37.930 221.200 ;
        RECT 51.530 220.000 57.930 221.200 ;
        RECT 71.530 220.000 77.930 221.200 ;
        RECT 91.530 220.000 97.930 221.200 ;
        RECT 9.340 196.350 11.675 197.050 ;
        RECT 10.110 194.410 11.985 194.770 ;
        RECT 12.335 194.415 14.215 194.775 ;
        RECT 11.530 158.800 17.930 160.000 ;
        RECT 31.530 158.800 37.930 160.000 ;
        RECT 51.530 158.800 57.930 160.000 ;
        RECT 71.530 158.800 77.930 160.000 ;
        RECT 91.530 158.800 97.930 160.000 ;
        RECT 14.230 158.150 15.230 158.800 ;
        RECT 34.230 158.150 35.230 158.800 ;
        RECT 54.230 158.150 55.230 158.800 ;
        RECT 74.230 158.150 75.230 158.800 ;
        RECT 94.230 158.150 95.230 158.800 ;
        RECT 10.880 158.000 18.580 158.150 ;
        RECT 30.880 158.000 38.580 158.150 ;
        RECT 50.880 158.000 58.580 158.150 ;
        RECT 70.880 158.000 78.580 158.150 ;
        RECT 90.880 158.000 98.580 158.150 ;
        RECT 5.930 153.200 6.680 155.000 ;
        RECT 4.730 150.450 6.680 153.200 ;
        RECT 4.730 149.550 4.880 150.450 ;
        RECT 5.530 150.300 6.680 150.450 ;
        RECT 6.830 150.300 6.980 157.850 ;
        RECT 7.430 150.300 7.580 157.850 ;
        RECT 8.030 150.300 8.180 157.850 ;
        RECT 8.630 150.300 8.780 157.850 ;
        RECT 9.230 150.300 9.380 157.850 ;
        RECT 9.830 150.300 9.980 157.850 ;
        RECT 14.230 157.550 15.230 158.000 ;
        RECT 10.880 157.400 18.580 157.550 ;
        RECT 14.230 156.950 15.230 157.400 ;
        RECT 10.880 156.800 18.580 156.950 ;
        RECT 14.230 156.350 15.230 156.800 ;
        RECT 10.880 156.200 18.580 156.350 ;
        RECT 14.230 155.750 15.230 156.200 ;
        RECT 10.880 155.600 18.580 155.750 ;
        RECT 14.230 155.150 15.230 155.600 ;
        RECT 10.880 155.000 18.580 155.150 ;
        RECT 14.230 154.550 15.230 155.000 ;
        RECT 10.880 154.400 18.580 154.550 ;
        RECT 14.230 153.950 15.230 154.400 ;
        RECT 10.880 153.800 18.580 153.950 ;
        RECT 14.230 153.350 15.230 153.800 ;
        RECT 10.880 153.200 18.580 153.350 ;
        RECT 14.230 152.750 15.230 153.200 ;
        RECT 10.880 152.600 18.580 152.750 ;
        RECT 14.230 152.150 15.230 152.600 ;
        RECT 10.880 152.000 18.580 152.150 ;
        RECT 14.230 151.550 15.230 152.000 ;
        RECT 10.880 151.400 18.580 151.550 ;
        RECT 14.230 150.950 15.230 151.400 ;
        RECT 10.880 150.800 18.580 150.950 ;
        RECT 14.230 150.300 15.230 150.800 ;
        RECT 19.480 150.300 19.630 157.850 ;
        RECT 20.080 150.300 20.230 157.850 ;
        RECT 20.680 150.300 20.830 157.850 ;
        RECT 21.280 150.300 21.430 157.850 ;
        RECT 21.880 150.300 22.030 157.850 ;
        RECT 22.480 150.300 22.630 157.850 ;
        RECT 22.780 153.200 23.530 155.000 ;
        RECT 25.930 153.200 26.680 155.000 ;
        RECT 22.780 150.450 26.680 153.200 ;
        RECT 22.780 150.300 23.930 150.450 ;
        RECT 5.530 149.700 23.930 150.300 ;
        RECT 5.530 149.550 6.680 149.700 ;
        RECT 4.730 146.800 6.680 149.550 ;
        RECT 5.930 145.050 6.680 146.800 ;
        RECT 6.830 142.150 6.980 149.700 ;
        RECT 7.430 142.150 7.580 149.700 ;
        RECT 8.030 142.150 8.180 149.700 ;
        RECT 8.630 142.150 8.780 149.700 ;
        RECT 9.230 142.150 9.380 149.700 ;
        RECT 9.830 142.150 9.980 149.700 ;
        RECT 14.230 149.200 15.230 149.700 ;
        RECT 10.880 149.050 18.580 149.200 ;
        RECT 14.230 148.600 15.230 149.050 ;
        RECT 10.880 148.450 18.580 148.600 ;
        RECT 14.230 148.000 15.230 148.450 ;
        RECT 10.880 147.850 18.580 148.000 ;
        RECT 14.230 147.400 15.230 147.850 ;
        RECT 10.880 147.250 18.580 147.400 ;
        RECT 14.230 146.800 15.230 147.250 ;
        RECT 10.880 146.650 18.580 146.800 ;
        RECT 14.230 146.200 15.230 146.650 ;
        RECT 10.880 146.050 18.580 146.200 ;
        RECT 14.230 145.600 15.230 146.050 ;
        RECT 10.880 145.450 18.580 145.600 ;
        RECT 14.230 145.000 15.230 145.450 ;
        RECT 10.880 144.850 18.580 145.000 ;
        RECT 14.230 144.400 15.230 144.850 ;
        RECT 10.880 144.250 18.580 144.400 ;
        RECT 14.230 143.800 15.230 144.250 ;
        RECT 10.880 143.650 18.580 143.800 ;
        RECT 14.230 143.200 15.230 143.650 ;
        RECT 10.880 143.050 18.580 143.200 ;
        RECT 14.230 142.600 15.230 143.050 ;
        RECT 10.880 142.450 18.580 142.600 ;
        RECT 14.230 142.000 15.230 142.450 ;
        RECT 19.480 142.150 19.630 149.700 ;
        RECT 20.080 142.150 20.230 149.700 ;
        RECT 20.680 142.150 20.830 149.700 ;
        RECT 21.280 142.150 21.430 149.700 ;
        RECT 21.880 142.150 22.030 149.700 ;
        RECT 22.480 142.150 22.630 149.700 ;
        RECT 22.780 149.550 23.930 149.700 ;
        RECT 24.580 149.550 24.880 150.450 ;
        RECT 25.530 150.300 26.680 150.450 ;
        RECT 26.830 150.300 26.980 157.850 ;
        RECT 27.430 150.300 27.580 157.850 ;
        RECT 28.030 150.300 28.180 157.850 ;
        RECT 28.630 150.300 28.780 157.850 ;
        RECT 29.230 150.300 29.380 157.850 ;
        RECT 29.830 150.300 29.980 157.850 ;
        RECT 34.230 157.550 35.230 158.000 ;
        RECT 30.880 157.400 38.580 157.550 ;
        RECT 34.230 156.950 35.230 157.400 ;
        RECT 30.880 156.800 38.580 156.950 ;
        RECT 34.230 156.350 35.230 156.800 ;
        RECT 30.880 156.200 38.580 156.350 ;
        RECT 34.230 155.750 35.230 156.200 ;
        RECT 30.880 155.600 38.580 155.750 ;
        RECT 34.230 155.150 35.230 155.600 ;
        RECT 30.880 155.000 38.580 155.150 ;
        RECT 34.230 154.550 35.230 155.000 ;
        RECT 30.880 154.400 38.580 154.550 ;
        RECT 34.230 153.950 35.230 154.400 ;
        RECT 30.880 153.800 38.580 153.950 ;
        RECT 34.230 153.350 35.230 153.800 ;
        RECT 30.880 153.200 38.580 153.350 ;
        RECT 34.230 152.750 35.230 153.200 ;
        RECT 30.880 152.600 38.580 152.750 ;
        RECT 34.230 152.150 35.230 152.600 ;
        RECT 30.880 152.000 38.580 152.150 ;
        RECT 34.230 151.550 35.230 152.000 ;
        RECT 30.880 151.400 38.580 151.550 ;
        RECT 34.230 150.950 35.230 151.400 ;
        RECT 30.880 150.800 38.580 150.950 ;
        RECT 34.230 150.300 35.230 150.800 ;
        RECT 39.480 150.300 39.630 157.850 ;
        RECT 40.080 150.300 40.230 157.850 ;
        RECT 40.680 150.300 40.830 157.850 ;
        RECT 41.280 150.300 41.430 157.850 ;
        RECT 41.880 150.300 42.030 157.850 ;
        RECT 42.480 150.300 42.630 157.850 ;
        RECT 42.780 153.200 43.530 155.000 ;
        RECT 45.930 153.200 46.680 155.000 ;
        RECT 42.780 150.450 46.680 153.200 ;
        RECT 42.780 150.300 43.930 150.450 ;
        RECT 25.530 149.700 43.930 150.300 ;
        RECT 25.530 149.550 26.680 149.700 ;
        RECT 22.780 146.800 26.680 149.550 ;
        RECT 22.780 145.050 23.530 146.800 ;
        RECT 25.930 145.050 26.680 146.800 ;
        RECT 26.830 142.150 26.980 149.700 ;
        RECT 27.430 142.150 27.580 149.700 ;
        RECT 28.030 142.150 28.180 149.700 ;
        RECT 28.630 142.150 28.780 149.700 ;
        RECT 29.230 142.150 29.380 149.700 ;
        RECT 29.830 142.150 29.980 149.700 ;
        RECT 34.230 149.200 35.230 149.700 ;
        RECT 30.880 149.050 38.580 149.200 ;
        RECT 34.230 148.600 35.230 149.050 ;
        RECT 30.880 148.450 38.580 148.600 ;
        RECT 34.230 148.000 35.230 148.450 ;
        RECT 30.880 147.850 38.580 148.000 ;
        RECT 34.230 147.400 35.230 147.850 ;
        RECT 30.880 147.250 38.580 147.400 ;
        RECT 34.230 146.800 35.230 147.250 ;
        RECT 30.880 146.650 38.580 146.800 ;
        RECT 34.230 146.200 35.230 146.650 ;
        RECT 30.880 146.050 38.580 146.200 ;
        RECT 34.230 145.600 35.230 146.050 ;
        RECT 30.880 145.450 38.580 145.600 ;
        RECT 34.230 145.000 35.230 145.450 ;
        RECT 30.880 144.850 38.580 145.000 ;
        RECT 34.230 144.400 35.230 144.850 ;
        RECT 30.880 144.250 38.580 144.400 ;
        RECT 34.230 143.800 35.230 144.250 ;
        RECT 30.880 143.650 38.580 143.800 ;
        RECT 34.230 143.200 35.230 143.650 ;
        RECT 30.880 143.050 38.580 143.200 ;
        RECT 34.230 142.600 35.230 143.050 ;
        RECT 30.880 142.450 38.580 142.600 ;
        RECT 34.230 142.000 35.230 142.450 ;
        RECT 39.480 142.150 39.630 149.700 ;
        RECT 40.080 142.150 40.230 149.700 ;
        RECT 40.680 142.150 40.830 149.700 ;
        RECT 41.280 142.150 41.430 149.700 ;
        RECT 41.880 142.150 42.030 149.700 ;
        RECT 42.480 142.150 42.630 149.700 ;
        RECT 42.780 149.550 43.930 149.700 ;
        RECT 44.580 149.550 44.880 150.450 ;
        RECT 45.530 150.300 46.680 150.450 ;
        RECT 46.830 150.300 46.980 157.850 ;
        RECT 47.430 150.300 47.580 157.850 ;
        RECT 48.030 150.300 48.180 157.850 ;
        RECT 48.630 150.300 48.780 157.850 ;
        RECT 49.230 150.300 49.380 157.850 ;
        RECT 49.830 150.300 49.980 157.850 ;
        RECT 54.230 157.550 55.230 158.000 ;
        RECT 50.880 157.400 58.580 157.550 ;
        RECT 54.230 156.950 55.230 157.400 ;
        RECT 50.880 156.800 58.580 156.950 ;
        RECT 54.230 156.350 55.230 156.800 ;
        RECT 50.880 156.200 58.580 156.350 ;
        RECT 54.230 155.750 55.230 156.200 ;
        RECT 50.880 155.600 58.580 155.750 ;
        RECT 54.230 155.150 55.230 155.600 ;
        RECT 50.880 155.000 58.580 155.150 ;
        RECT 54.230 154.550 55.230 155.000 ;
        RECT 50.880 154.400 58.580 154.550 ;
        RECT 54.230 153.950 55.230 154.400 ;
        RECT 50.880 153.800 58.580 153.950 ;
        RECT 54.230 153.350 55.230 153.800 ;
        RECT 50.880 153.200 58.580 153.350 ;
        RECT 54.230 152.750 55.230 153.200 ;
        RECT 50.880 152.600 58.580 152.750 ;
        RECT 54.230 152.150 55.230 152.600 ;
        RECT 50.880 152.000 58.580 152.150 ;
        RECT 54.230 151.550 55.230 152.000 ;
        RECT 50.880 151.400 58.580 151.550 ;
        RECT 54.230 150.950 55.230 151.400 ;
        RECT 50.880 150.800 58.580 150.950 ;
        RECT 54.230 150.300 55.230 150.800 ;
        RECT 59.480 150.300 59.630 157.850 ;
        RECT 60.080 150.300 60.230 157.850 ;
        RECT 60.680 150.300 60.830 157.850 ;
        RECT 61.280 150.300 61.430 157.850 ;
        RECT 61.880 150.300 62.030 157.850 ;
        RECT 62.480 150.300 62.630 157.850 ;
        RECT 62.780 153.200 63.530 155.000 ;
        RECT 65.930 153.200 66.680 155.000 ;
        RECT 62.780 150.450 66.680 153.200 ;
        RECT 62.780 150.300 63.930 150.450 ;
        RECT 45.530 149.700 63.930 150.300 ;
        RECT 45.530 149.550 46.680 149.700 ;
        RECT 42.780 146.800 46.680 149.550 ;
        RECT 42.780 145.050 43.530 146.800 ;
        RECT 45.930 145.050 46.680 146.800 ;
        RECT 46.830 142.150 46.980 149.700 ;
        RECT 47.430 142.150 47.580 149.700 ;
        RECT 48.030 142.150 48.180 149.700 ;
        RECT 48.630 142.150 48.780 149.700 ;
        RECT 49.230 142.150 49.380 149.700 ;
        RECT 49.830 142.150 49.980 149.700 ;
        RECT 54.230 149.200 55.230 149.700 ;
        RECT 50.880 149.050 58.580 149.200 ;
        RECT 54.230 148.600 55.230 149.050 ;
        RECT 50.880 148.450 58.580 148.600 ;
        RECT 54.230 148.000 55.230 148.450 ;
        RECT 50.880 147.850 58.580 148.000 ;
        RECT 54.230 147.400 55.230 147.850 ;
        RECT 50.880 147.250 58.580 147.400 ;
        RECT 54.230 146.800 55.230 147.250 ;
        RECT 50.880 146.650 58.580 146.800 ;
        RECT 54.230 146.200 55.230 146.650 ;
        RECT 50.880 146.050 58.580 146.200 ;
        RECT 54.230 145.600 55.230 146.050 ;
        RECT 50.880 145.450 58.580 145.600 ;
        RECT 54.230 145.000 55.230 145.450 ;
        RECT 50.880 144.850 58.580 145.000 ;
        RECT 54.230 144.400 55.230 144.850 ;
        RECT 50.880 144.250 58.580 144.400 ;
        RECT 54.230 143.800 55.230 144.250 ;
        RECT 50.880 143.650 58.580 143.800 ;
        RECT 54.230 143.200 55.230 143.650 ;
        RECT 50.880 143.050 58.580 143.200 ;
        RECT 54.230 142.600 55.230 143.050 ;
        RECT 50.880 142.450 58.580 142.600 ;
        RECT 54.230 142.000 55.230 142.450 ;
        RECT 59.480 142.150 59.630 149.700 ;
        RECT 60.080 142.150 60.230 149.700 ;
        RECT 60.680 142.150 60.830 149.700 ;
        RECT 61.280 142.150 61.430 149.700 ;
        RECT 61.880 142.150 62.030 149.700 ;
        RECT 62.480 142.150 62.630 149.700 ;
        RECT 62.780 149.550 63.930 149.700 ;
        RECT 64.580 149.550 64.880 150.450 ;
        RECT 65.530 150.300 66.680 150.450 ;
        RECT 66.830 150.300 66.980 157.850 ;
        RECT 67.430 150.300 67.580 157.850 ;
        RECT 68.030 150.300 68.180 157.850 ;
        RECT 68.630 150.300 68.780 157.850 ;
        RECT 69.230 150.300 69.380 157.850 ;
        RECT 69.830 150.300 69.980 157.850 ;
        RECT 74.230 157.550 75.230 158.000 ;
        RECT 70.880 157.400 78.580 157.550 ;
        RECT 74.230 156.950 75.230 157.400 ;
        RECT 70.880 156.800 78.580 156.950 ;
        RECT 74.230 156.350 75.230 156.800 ;
        RECT 70.880 156.200 78.580 156.350 ;
        RECT 74.230 155.750 75.230 156.200 ;
        RECT 70.880 155.600 78.580 155.750 ;
        RECT 74.230 155.150 75.230 155.600 ;
        RECT 70.880 155.000 78.580 155.150 ;
        RECT 74.230 154.550 75.230 155.000 ;
        RECT 70.880 154.400 78.580 154.550 ;
        RECT 74.230 153.950 75.230 154.400 ;
        RECT 70.880 153.800 78.580 153.950 ;
        RECT 74.230 153.350 75.230 153.800 ;
        RECT 70.880 153.200 78.580 153.350 ;
        RECT 74.230 152.750 75.230 153.200 ;
        RECT 70.880 152.600 78.580 152.750 ;
        RECT 74.230 152.150 75.230 152.600 ;
        RECT 70.880 152.000 78.580 152.150 ;
        RECT 74.230 151.550 75.230 152.000 ;
        RECT 70.880 151.400 78.580 151.550 ;
        RECT 74.230 150.950 75.230 151.400 ;
        RECT 70.880 150.800 78.580 150.950 ;
        RECT 74.230 150.300 75.230 150.800 ;
        RECT 79.480 150.300 79.630 157.850 ;
        RECT 80.080 150.300 80.230 157.850 ;
        RECT 80.680 150.300 80.830 157.850 ;
        RECT 81.280 150.300 81.430 157.850 ;
        RECT 81.880 150.300 82.030 157.850 ;
        RECT 82.480 150.300 82.630 157.850 ;
        RECT 82.780 153.200 83.530 155.000 ;
        RECT 85.930 153.200 86.680 155.000 ;
        RECT 82.780 150.450 86.680 153.200 ;
        RECT 82.780 150.300 83.930 150.450 ;
        RECT 65.530 149.700 83.930 150.300 ;
        RECT 65.530 149.550 66.680 149.700 ;
        RECT 62.780 146.800 66.680 149.550 ;
        RECT 62.780 145.050 63.530 146.800 ;
        RECT 65.930 145.050 66.680 146.800 ;
        RECT 66.830 142.150 66.980 149.700 ;
        RECT 67.430 142.150 67.580 149.700 ;
        RECT 68.030 142.150 68.180 149.700 ;
        RECT 68.630 142.150 68.780 149.700 ;
        RECT 69.230 142.150 69.380 149.700 ;
        RECT 69.830 142.150 69.980 149.700 ;
        RECT 74.230 149.200 75.230 149.700 ;
        RECT 70.880 149.050 78.580 149.200 ;
        RECT 74.230 148.600 75.230 149.050 ;
        RECT 70.880 148.450 78.580 148.600 ;
        RECT 74.230 148.000 75.230 148.450 ;
        RECT 70.880 147.850 78.580 148.000 ;
        RECT 74.230 147.400 75.230 147.850 ;
        RECT 70.880 147.250 78.580 147.400 ;
        RECT 74.230 146.800 75.230 147.250 ;
        RECT 70.880 146.650 78.580 146.800 ;
        RECT 74.230 146.200 75.230 146.650 ;
        RECT 70.880 146.050 78.580 146.200 ;
        RECT 74.230 145.600 75.230 146.050 ;
        RECT 70.880 145.450 78.580 145.600 ;
        RECT 74.230 145.000 75.230 145.450 ;
        RECT 70.880 144.850 78.580 145.000 ;
        RECT 74.230 144.400 75.230 144.850 ;
        RECT 70.880 144.250 78.580 144.400 ;
        RECT 74.230 143.800 75.230 144.250 ;
        RECT 70.880 143.650 78.580 143.800 ;
        RECT 74.230 143.200 75.230 143.650 ;
        RECT 70.880 143.050 78.580 143.200 ;
        RECT 74.230 142.600 75.230 143.050 ;
        RECT 70.880 142.450 78.580 142.600 ;
        RECT 74.230 142.000 75.230 142.450 ;
        RECT 79.480 142.150 79.630 149.700 ;
        RECT 80.080 142.150 80.230 149.700 ;
        RECT 80.680 142.150 80.830 149.700 ;
        RECT 81.280 142.150 81.430 149.700 ;
        RECT 81.880 142.150 82.030 149.700 ;
        RECT 82.480 142.150 82.630 149.700 ;
        RECT 82.780 149.550 83.930 149.700 ;
        RECT 84.580 149.550 84.880 150.450 ;
        RECT 85.530 150.300 86.680 150.450 ;
        RECT 86.830 150.300 86.980 157.850 ;
        RECT 87.430 150.300 87.580 157.850 ;
        RECT 88.030 150.300 88.180 157.850 ;
        RECT 88.630 150.300 88.780 157.850 ;
        RECT 89.230 150.300 89.380 157.850 ;
        RECT 89.830 150.300 89.980 157.850 ;
        RECT 94.230 157.550 95.230 158.000 ;
        RECT 90.880 157.400 98.580 157.550 ;
        RECT 94.230 156.950 95.230 157.400 ;
        RECT 90.880 156.800 98.580 156.950 ;
        RECT 94.230 156.350 95.230 156.800 ;
        RECT 90.880 156.200 98.580 156.350 ;
        RECT 94.230 155.750 95.230 156.200 ;
        RECT 90.880 155.600 98.580 155.750 ;
        RECT 94.230 155.150 95.230 155.600 ;
        RECT 90.880 155.000 98.580 155.150 ;
        RECT 94.230 154.550 95.230 155.000 ;
        RECT 90.880 154.400 98.580 154.550 ;
        RECT 94.230 153.950 95.230 154.400 ;
        RECT 90.880 153.800 98.580 153.950 ;
        RECT 94.230 153.350 95.230 153.800 ;
        RECT 90.880 153.200 98.580 153.350 ;
        RECT 94.230 152.750 95.230 153.200 ;
        RECT 90.880 152.600 98.580 152.750 ;
        RECT 94.230 152.150 95.230 152.600 ;
        RECT 90.880 152.000 98.580 152.150 ;
        RECT 94.230 151.550 95.230 152.000 ;
        RECT 90.880 151.400 98.580 151.550 ;
        RECT 94.230 150.950 95.230 151.400 ;
        RECT 90.880 150.800 98.580 150.950 ;
        RECT 94.230 150.300 95.230 150.800 ;
        RECT 99.480 150.300 99.630 157.850 ;
        RECT 100.080 150.300 100.230 157.850 ;
        RECT 100.680 150.300 100.830 157.850 ;
        RECT 101.280 150.300 101.430 157.850 ;
        RECT 101.880 150.300 102.030 157.850 ;
        RECT 102.480 150.300 102.630 157.850 ;
        RECT 102.780 153.200 103.530 155.000 ;
        RECT 102.780 150.775 104.730 153.200 ;
        RECT 102.780 150.450 111.850 150.775 ;
        RECT 102.780 150.300 103.930 150.450 ;
        RECT 85.530 149.700 103.930 150.300 ;
        RECT 85.530 149.550 86.680 149.700 ;
        RECT 82.780 146.800 86.680 149.550 ;
        RECT 82.780 145.050 83.530 146.800 ;
        RECT 85.930 145.050 86.680 146.800 ;
        RECT 86.830 142.150 86.980 149.700 ;
        RECT 87.430 142.150 87.580 149.700 ;
        RECT 88.030 142.150 88.180 149.700 ;
        RECT 88.630 142.150 88.780 149.700 ;
        RECT 89.230 142.150 89.380 149.700 ;
        RECT 89.830 142.150 89.980 149.700 ;
        RECT 94.230 149.200 95.230 149.700 ;
        RECT 90.880 149.050 98.580 149.200 ;
        RECT 94.230 148.600 95.230 149.050 ;
        RECT 90.880 148.450 98.580 148.600 ;
        RECT 94.230 148.000 95.230 148.450 ;
        RECT 90.880 147.850 98.580 148.000 ;
        RECT 94.230 147.400 95.230 147.850 ;
        RECT 90.880 147.250 98.580 147.400 ;
        RECT 94.230 146.800 95.230 147.250 ;
        RECT 90.880 146.650 98.580 146.800 ;
        RECT 94.230 146.200 95.230 146.650 ;
        RECT 90.880 146.050 98.580 146.200 ;
        RECT 94.230 145.600 95.230 146.050 ;
        RECT 90.880 145.450 98.580 145.600 ;
        RECT 94.230 145.000 95.230 145.450 ;
        RECT 90.880 144.850 98.580 145.000 ;
        RECT 94.230 144.400 95.230 144.850 ;
        RECT 90.880 144.250 98.580 144.400 ;
        RECT 94.230 143.800 95.230 144.250 ;
        RECT 90.880 143.650 98.580 143.800 ;
        RECT 94.230 143.200 95.230 143.650 ;
        RECT 90.880 143.050 98.580 143.200 ;
        RECT 94.230 142.600 95.230 143.050 ;
        RECT 90.880 142.450 98.580 142.600 ;
        RECT 94.230 142.000 95.230 142.450 ;
        RECT 99.480 142.150 99.630 149.700 ;
        RECT 100.080 142.150 100.230 149.700 ;
        RECT 100.680 142.150 100.830 149.700 ;
        RECT 101.280 142.150 101.430 149.700 ;
        RECT 101.880 142.150 102.030 149.700 ;
        RECT 102.480 142.150 102.630 149.700 ;
        RECT 102.780 149.550 103.930 149.700 ;
        RECT 104.580 149.550 111.850 150.450 ;
        RECT 102.780 149.500 111.850 149.550 ;
        RECT 102.780 146.800 104.730 149.500 ;
        RECT 102.780 145.050 103.530 146.800 ;
        RECT 10.880 141.850 18.580 142.000 ;
        RECT 30.880 141.850 38.580 142.000 ;
        RECT 50.880 141.850 58.580 142.000 ;
        RECT 70.880 141.850 78.580 142.000 ;
        RECT 90.880 141.850 98.580 142.000 ;
        RECT 14.230 141.200 15.230 141.850 ;
        RECT 34.230 141.200 35.230 141.850 ;
        RECT 54.230 141.200 55.230 141.850 ;
        RECT 74.230 141.200 75.230 141.850 ;
        RECT 94.230 141.200 95.230 141.850 ;
        RECT 11.530 138.800 17.930 141.200 ;
        RECT 31.530 138.800 37.930 141.200 ;
        RECT 51.530 138.800 57.930 141.200 ;
        RECT 71.530 138.800 77.930 141.200 ;
        RECT 91.530 138.800 97.930 141.200 ;
        RECT 14.230 138.150 15.230 138.800 ;
        RECT 34.230 138.150 35.230 138.800 ;
        RECT 54.230 138.150 55.230 138.800 ;
        RECT 74.230 138.150 75.230 138.800 ;
        RECT 94.230 138.150 95.230 138.800 ;
        RECT 10.880 138.000 18.580 138.150 ;
        RECT 30.880 138.000 38.580 138.150 ;
        RECT 50.880 138.000 58.580 138.150 ;
        RECT 70.880 138.000 78.580 138.150 ;
        RECT 90.880 138.000 98.580 138.150 ;
        RECT 5.930 133.200 6.680 135.000 ;
        RECT 4.730 130.450 6.680 133.200 ;
        RECT 4.730 129.550 4.880 130.450 ;
        RECT 5.530 130.300 6.680 130.450 ;
        RECT 6.830 130.300 6.980 137.850 ;
        RECT 7.430 130.300 7.580 137.850 ;
        RECT 8.030 130.300 8.180 137.850 ;
        RECT 8.630 130.300 8.780 137.850 ;
        RECT 9.230 130.300 9.380 137.850 ;
        RECT 9.830 130.300 9.980 137.850 ;
        RECT 14.230 137.550 15.230 138.000 ;
        RECT 10.880 137.400 18.580 137.550 ;
        RECT 14.230 136.950 15.230 137.400 ;
        RECT 10.880 136.800 18.580 136.950 ;
        RECT 14.230 136.350 15.230 136.800 ;
        RECT 10.880 136.200 18.580 136.350 ;
        RECT 14.230 135.750 15.230 136.200 ;
        RECT 10.880 135.600 18.580 135.750 ;
        RECT 14.230 135.150 15.230 135.600 ;
        RECT 10.880 135.000 18.580 135.150 ;
        RECT 14.230 134.550 15.230 135.000 ;
        RECT 10.880 134.400 18.580 134.550 ;
        RECT 14.230 133.950 15.230 134.400 ;
        RECT 10.880 133.800 18.580 133.950 ;
        RECT 14.230 133.350 15.230 133.800 ;
        RECT 10.880 133.200 18.580 133.350 ;
        RECT 14.230 132.750 15.230 133.200 ;
        RECT 10.880 132.600 18.580 132.750 ;
        RECT 14.230 132.150 15.230 132.600 ;
        RECT 10.880 132.000 18.580 132.150 ;
        RECT 14.230 131.550 15.230 132.000 ;
        RECT 10.880 131.400 18.580 131.550 ;
        RECT 14.230 130.950 15.230 131.400 ;
        RECT 10.880 130.800 18.580 130.950 ;
        RECT 14.230 130.300 15.230 130.800 ;
        RECT 19.480 130.300 19.630 137.850 ;
        RECT 20.080 130.300 20.230 137.850 ;
        RECT 20.680 130.300 20.830 137.850 ;
        RECT 21.280 130.300 21.430 137.850 ;
        RECT 21.880 130.300 22.030 137.850 ;
        RECT 22.480 130.300 22.630 137.850 ;
        RECT 22.780 133.200 23.530 135.000 ;
        RECT 25.930 133.200 26.680 135.000 ;
        RECT 22.780 130.450 26.680 133.200 ;
        RECT 22.780 130.300 23.930 130.450 ;
        RECT 5.530 129.700 23.930 130.300 ;
        RECT 5.530 129.550 6.680 129.700 ;
        RECT 4.730 126.800 6.680 129.550 ;
        RECT 5.930 125.050 6.680 126.800 ;
        RECT 6.830 122.150 6.980 129.700 ;
        RECT 7.430 122.150 7.580 129.700 ;
        RECT 8.030 122.150 8.180 129.700 ;
        RECT 8.630 122.150 8.780 129.700 ;
        RECT 9.230 122.150 9.380 129.700 ;
        RECT 9.830 122.150 9.980 129.700 ;
        RECT 14.230 129.200 15.230 129.700 ;
        RECT 10.880 129.050 18.580 129.200 ;
        RECT 14.230 128.600 15.230 129.050 ;
        RECT 10.880 128.450 18.580 128.600 ;
        RECT 14.230 128.000 15.230 128.450 ;
        RECT 10.880 127.850 18.580 128.000 ;
        RECT 14.230 127.400 15.230 127.850 ;
        RECT 10.880 127.250 18.580 127.400 ;
        RECT 14.230 126.800 15.230 127.250 ;
        RECT 10.880 126.650 18.580 126.800 ;
        RECT 14.230 126.200 15.230 126.650 ;
        RECT 10.880 126.050 18.580 126.200 ;
        RECT 14.230 125.600 15.230 126.050 ;
        RECT 10.880 125.450 18.580 125.600 ;
        RECT 14.230 125.000 15.230 125.450 ;
        RECT 10.880 124.850 18.580 125.000 ;
        RECT 14.230 124.400 15.230 124.850 ;
        RECT 10.880 124.250 18.580 124.400 ;
        RECT 14.230 123.800 15.230 124.250 ;
        RECT 10.880 123.650 18.580 123.800 ;
        RECT 14.230 123.200 15.230 123.650 ;
        RECT 10.880 123.050 18.580 123.200 ;
        RECT 14.230 122.600 15.230 123.050 ;
        RECT 10.880 122.450 18.580 122.600 ;
        RECT 14.230 122.000 15.230 122.450 ;
        RECT 19.480 122.150 19.630 129.700 ;
        RECT 20.080 122.150 20.230 129.700 ;
        RECT 20.680 122.150 20.830 129.700 ;
        RECT 21.280 122.150 21.430 129.700 ;
        RECT 21.880 122.150 22.030 129.700 ;
        RECT 22.480 122.150 22.630 129.700 ;
        RECT 22.780 129.550 23.930 129.700 ;
        RECT 24.580 129.550 24.880 130.450 ;
        RECT 25.530 130.300 26.680 130.450 ;
        RECT 26.830 130.300 26.980 137.850 ;
        RECT 27.430 130.300 27.580 137.850 ;
        RECT 28.030 130.300 28.180 137.850 ;
        RECT 28.630 130.300 28.780 137.850 ;
        RECT 29.230 130.300 29.380 137.850 ;
        RECT 29.830 130.300 29.980 137.850 ;
        RECT 34.230 137.550 35.230 138.000 ;
        RECT 30.880 137.400 38.580 137.550 ;
        RECT 34.230 136.950 35.230 137.400 ;
        RECT 30.880 136.800 38.580 136.950 ;
        RECT 34.230 136.350 35.230 136.800 ;
        RECT 30.880 136.200 38.580 136.350 ;
        RECT 34.230 135.750 35.230 136.200 ;
        RECT 30.880 135.600 38.580 135.750 ;
        RECT 34.230 135.150 35.230 135.600 ;
        RECT 30.880 135.000 38.580 135.150 ;
        RECT 34.230 134.550 35.230 135.000 ;
        RECT 30.880 134.400 38.580 134.550 ;
        RECT 34.230 133.950 35.230 134.400 ;
        RECT 30.880 133.800 38.580 133.950 ;
        RECT 34.230 133.350 35.230 133.800 ;
        RECT 30.880 133.200 38.580 133.350 ;
        RECT 34.230 132.750 35.230 133.200 ;
        RECT 30.880 132.600 38.580 132.750 ;
        RECT 34.230 132.150 35.230 132.600 ;
        RECT 30.880 132.000 38.580 132.150 ;
        RECT 34.230 131.550 35.230 132.000 ;
        RECT 30.880 131.400 38.580 131.550 ;
        RECT 34.230 130.950 35.230 131.400 ;
        RECT 30.880 130.800 38.580 130.950 ;
        RECT 34.230 130.300 35.230 130.800 ;
        RECT 39.480 130.300 39.630 137.850 ;
        RECT 40.080 130.300 40.230 137.850 ;
        RECT 40.680 130.300 40.830 137.850 ;
        RECT 41.280 130.300 41.430 137.850 ;
        RECT 41.880 130.300 42.030 137.850 ;
        RECT 42.480 130.300 42.630 137.850 ;
        RECT 42.780 133.200 43.530 135.000 ;
        RECT 45.930 133.200 46.680 135.000 ;
        RECT 42.780 130.450 46.680 133.200 ;
        RECT 42.780 130.300 43.930 130.450 ;
        RECT 25.530 129.700 43.930 130.300 ;
        RECT 25.530 129.550 26.680 129.700 ;
        RECT 22.780 126.800 26.680 129.550 ;
        RECT 22.780 125.050 23.530 126.800 ;
        RECT 25.930 125.050 26.680 126.800 ;
        RECT 26.830 122.150 26.980 129.700 ;
        RECT 27.430 122.150 27.580 129.700 ;
        RECT 28.030 122.150 28.180 129.700 ;
        RECT 28.630 122.150 28.780 129.700 ;
        RECT 29.230 122.150 29.380 129.700 ;
        RECT 29.830 122.150 29.980 129.700 ;
        RECT 34.230 129.200 35.230 129.700 ;
        RECT 30.880 129.050 38.580 129.200 ;
        RECT 34.230 128.600 35.230 129.050 ;
        RECT 30.880 128.450 38.580 128.600 ;
        RECT 34.230 128.000 35.230 128.450 ;
        RECT 30.880 127.850 38.580 128.000 ;
        RECT 34.230 127.400 35.230 127.850 ;
        RECT 30.880 127.250 38.580 127.400 ;
        RECT 34.230 126.800 35.230 127.250 ;
        RECT 30.880 126.650 38.580 126.800 ;
        RECT 34.230 126.200 35.230 126.650 ;
        RECT 30.880 126.050 38.580 126.200 ;
        RECT 34.230 125.600 35.230 126.050 ;
        RECT 30.880 125.450 38.580 125.600 ;
        RECT 34.230 125.000 35.230 125.450 ;
        RECT 30.880 124.850 38.580 125.000 ;
        RECT 34.230 124.400 35.230 124.850 ;
        RECT 30.880 124.250 38.580 124.400 ;
        RECT 34.230 123.800 35.230 124.250 ;
        RECT 30.880 123.650 38.580 123.800 ;
        RECT 34.230 123.200 35.230 123.650 ;
        RECT 30.880 123.050 38.580 123.200 ;
        RECT 34.230 122.600 35.230 123.050 ;
        RECT 30.880 122.450 38.580 122.600 ;
        RECT 34.230 122.000 35.230 122.450 ;
        RECT 39.480 122.150 39.630 129.700 ;
        RECT 40.080 122.150 40.230 129.700 ;
        RECT 40.680 122.150 40.830 129.700 ;
        RECT 41.280 122.150 41.430 129.700 ;
        RECT 41.880 122.150 42.030 129.700 ;
        RECT 42.480 122.150 42.630 129.700 ;
        RECT 42.780 129.550 43.930 129.700 ;
        RECT 44.580 129.550 44.880 130.450 ;
        RECT 45.530 130.300 46.680 130.450 ;
        RECT 46.830 130.300 46.980 137.850 ;
        RECT 47.430 130.300 47.580 137.850 ;
        RECT 48.030 130.300 48.180 137.850 ;
        RECT 48.630 130.300 48.780 137.850 ;
        RECT 49.230 130.300 49.380 137.850 ;
        RECT 49.830 130.300 49.980 137.850 ;
        RECT 54.230 137.550 55.230 138.000 ;
        RECT 50.880 137.400 58.580 137.550 ;
        RECT 54.230 136.950 55.230 137.400 ;
        RECT 50.880 136.800 58.580 136.950 ;
        RECT 54.230 136.350 55.230 136.800 ;
        RECT 50.880 136.200 58.580 136.350 ;
        RECT 54.230 135.750 55.230 136.200 ;
        RECT 50.880 135.600 58.580 135.750 ;
        RECT 54.230 135.150 55.230 135.600 ;
        RECT 50.880 135.000 58.580 135.150 ;
        RECT 54.230 134.550 55.230 135.000 ;
        RECT 50.880 134.400 58.580 134.550 ;
        RECT 54.230 133.950 55.230 134.400 ;
        RECT 50.880 133.800 58.580 133.950 ;
        RECT 54.230 133.350 55.230 133.800 ;
        RECT 50.880 133.200 58.580 133.350 ;
        RECT 54.230 132.750 55.230 133.200 ;
        RECT 50.880 132.600 58.580 132.750 ;
        RECT 54.230 132.150 55.230 132.600 ;
        RECT 50.880 132.000 58.580 132.150 ;
        RECT 54.230 131.550 55.230 132.000 ;
        RECT 50.880 131.400 58.580 131.550 ;
        RECT 54.230 130.950 55.230 131.400 ;
        RECT 50.880 130.800 58.580 130.950 ;
        RECT 54.230 130.300 55.230 130.800 ;
        RECT 59.480 130.300 59.630 137.850 ;
        RECT 60.080 130.300 60.230 137.850 ;
        RECT 60.680 130.300 60.830 137.850 ;
        RECT 61.280 130.300 61.430 137.850 ;
        RECT 61.880 130.300 62.030 137.850 ;
        RECT 62.480 130.300 62.630 137.850 ;
        RECT 62.780 133.200 63.530 135.000 ;
        RECT 65.930 133.200 66.680 135.000 ;
        RECT 62.780 130.450 66.680 133.200 ;
        RECT 62.780 130.300 63.930 130.450 ;
        RECT 45.530 129.700 63.930 130.300 ;
        RECT 45.530 129.550 46.680 129.700 ;
        RECT 42.780 126.800 46.680 129.550 ;
        RECT 42.780 125.050 43.530 126.800 ;
        RECT 45.930 125.050 46.680 126.800 ;
        RECT 46.830 122.150 46.980 129.700 ;
        RECT 47.430 122.150 47.580 129.700 ;
        RECT 48.030 122.150 48.180 129.700 ;
        RECT 48.630 122.150 48.780 129.700 ;
        RECT 49.230 122.150 49.380 129.700 ;
        RECT 49.830 122.150 49.980 129.700 ;
        RECT 54.230 129.200 55.230 129.700 ;
        RECT 50.880 129.050 58.580 129.200 ;
        RECT 54.230 128.600 55.230 129.050 ;
        RECT 50.880 128.450 58.580 128.600 ;
        RECT 54.230 128.000 55.230 128.450 ;
        RECT 50.880 127.850 58.580 128.000 ;
        RECT 54.230 127.400 55.230 127.850 ;
        RECT 50.880 127.250 58.580 127.400 ;
        RECT 54.230 126.800 55.230 127.250 ;
        RECT 50.880 126.650 58.580 126.800 ;
        RECT 54.230 126.200 55.230 126.650 ;
        RECT 50.880 126.050 58.580 126.200 ;
        RECT 54.230 125.600 55.230 126.050 ;
        RECT 50.880 125.450 58.580 125.600 ;
        RECT 54.230 125.000 55.230 125.450 ;
        RECT 50.880 124.850 58.580 125.000 ;
        RECT 54.230 124.400 55.230 124.850 ;
        RECT 50.880 124.250 58.580 124.400 ;
        RECT 54.230 123.800 55.230 124.250 ;
        RECT 50.880 123.650 58.580 123.800 ;
        RECT 54.230 123.200 55.230 123.650 ;
        RECT 50.880 123.050 58.580 123.200 ;
        RECT 54.230 122.600 55.230 123.050 ;
        RECT 50.880 122.450 58.580 122.600 ;
        RECT 54.230 122.000 55.230 122.450 ;
        RECT 59.480 122.150 59.630 129.700 ;
        RECT 60.080 122.150 60.230 129.700 ;
        RECT 60.680 122.150 60.830 129.700 ;
        RECT 61.280 122.150 61.430 129.700 ;
        RECT 61.880 122.150 62.030 129.700 ;
        RECT 62.480 122.150 62.630 129.700 ;
        RECT 62.780 129.550 63.930 129.700 ;
        RECT 64.580 129.550 64.880 130.450 ;
        RECT 65.530 130.300 66.680 130.450 ;
        RECT 66.830 130.300 66.980 137.850 ;
        RECT 67.430 130.300 67.580 137.850 ;
        RECT 68.030 130.300 68.180 137.850 ;
        RECT 68.630 130.300 68.780 137.850 ;
        RECT 69.230 130.300 69.380 137.850 ;
        RECT 69.830 130.300 69.980 137.850 ;
        RECT 74.230 137.550 75.230 138.000 ;
        RECT 70.880 137.400 78.580 137.550 ;
        RECT 74.230 136.950 75.230 137.400 ;
        RECT 70.880 136.800 78.580 136.950 ;
        RECT 74.230 136.350 75.230 136.800 ;
        RECT 70.880 136.200 78.580 136.350 ;
        RECT 74.230 135.750 75.230 136.200 ;
        RECT 70.880 135.600 78.580 135.750 ;
        RECT 74.230 135.150 75.230 135.600 ;
        RECT 70.880 135.000 78.580 135.150 ;
        RECT 74.230 134.550 75.230 135.000 ;
        RECT 70.880 134.400 78.580 134.550 ;
        RECT 74.230 133.950 75.230 134.400 ;
        RECT 70.880 133.800 78.580 133.950 ;
        RECT 74.230 133.350 75.230 133.800 ;
        RECT 70.880 133.200 78.580 133.350 ;
        RECT 74.230 132.750 75.230 133.200 ;
        RECT 70.880 132.600 78.580 132.750 ;
        RECT 74.230 132.150 75.230 132.600 ;
        RECT 70.880 132.000 78.580 132.150 ;
        RECT 74.230 131.550 75.230 132.000 ;
        RECT 70.880 131.400 78.580 131.550 ;
        RECT 74.230 130.950 75.230 131.400 ;
        RECT 70.880 130.800 78.580 130.950 ;
        RECT 74.230 130.300 75.230 130.800 ;
        RECT 79.480 130.300 79.630 137.850 ;
        RECT 80.080 130.300 80.230 137.850 ;
        RECT 80.680 130.300 80.830 137.850 ;
        RECT 81.280 130.300 81.430 137.850 ;
        RECT 81.880 130.300 82.030 137.850 ;
        RECT 82.480 130.300 82.630 137.850 ;
        RECT 82.780 133.200 83.530 135.000 ;
        RECT 85.930 133.200 86.680 135.000 ;
        RECT 82.780 130.450 86.680 133.200 ;
        RECT 82.780 130.300 83.930 130.450 ;
        RECT 65.530 129.700 83.930 130.300 ;
        RECT 65.530 129.550 66.680 129.700 ;
        RECT 62.780 126.800 66.680 129.550 ;
        RECT 62.780 125.050 63.530 126.800 ;
        RECT 65.930 125.050 66.680 126.800 ;
        RECT 66.830 122.150 66.980 129.700 ;
        RECT 67.430 122.150 67.580 129.700 ;
        RECT 68.030 122.150 68.180 129.700 ;
        RECT 68.630 122.150 68.780 129.700 ;
        RECT 69.230 122.150 69.380 129.700 ;
        RECT 69.830 122.150 69.980 129.700 ;
        RECT 74.230 129.200 75.230 129.700 ;
        RECT 70.880 129.050 78.580 129.200 ;
        RECT 74.230 128.600 75.230 129.050 ;
        RECT 70.880 128.450 78.580 128.600 ;
        RECT 74.230 128.000 75.230 128.450 ;
        RECT 70.880 127.850 78.580 128.000 ;
        RECT 74.230 127.400 75.230 127.850 ;
        RECT 70.880 127.250 78.580 127.400 ;
        RECT 74.230 126.800 75.230 127.250 ;
        RECT 70.880 126.650 78.580 126.800 ;
        RECT 74.230 126.200 75.230 126.650 ;
        RECT 70.880 126.050 78.580 126.200 ;
        RECT 74.230 125.600 75.230 126.050 ;
        RECT 70.880 125.450 78.580 125.600 ;
        RECT 74.230 125.000 75.230 125.450 ;
        RECT 70.880 124.850 78.580 125.000 ;
        RECT 74.230 124.400 75.230 124.850 ;
        RECT 70.880 124.250 78.580 124.400 ;
        RECT 74.230 123.800 75.230 124.250 ;
        RECT 70.880 123.650 78.580 123.800 ;
        RECT 74.230 123.200 75.230 123.650 ;
        RECT 70.880 123.050 78.580 123.200 ;
        RECT 74.230 122.600 75.230 123.050 ;
        RECT 70.880 122.450 78.580 122.600 ;
        RECT 74.230 122.000 75.230 122.450 ;
        RECT 79.480 122.150 79.630 129.700 ;
        RECT 80.080 122.150 80.230 129.700 ;
        RECT 80.680 122.150 80.830 129.700 ;
        RECT 81.280 122.150 81.430 129.700 ;
        RECT 81.880 122.150 82.030 129.700 ;
        RECT 82.480 122.150 82.630 129.700 ;
        RECT 82.780 129.550 83.930 129.700 ;
        RECT 84.580 129.550 84.880 130.450 ;
        RECT 85.530 130.300 86.680 130.450 ;
        RECT 86.830 130.300 86.980 137.850 ;
        RECT 87.430 130.300 87.580 137.850 ;
        RECT 88.030 130.300 88.180 137.850 ;
        RECT 88.630 130.300 88.780 137.850 ;
        RECT 89.230 130.300 89.380 137.850 ;
        RECT 89.830 130.300 89.980 137.850 ;
        RECT 94.230 137.550 95.230 138.000 ;
        RECT 90.880 137.400 98.580 137.550 ;
        RECT 94.230 136.950 95.230 137.400 ;
        RECT 90.880 136.800 98.580 136.950 ;
        RECT 94.230 136.350 95.230 136.800 ;
        RECT 90.880 136.200 98.580 136.350 ;
        RECT 94.230 135.750 95.230 136.200 ;
        RECT 90.880 135.600 98.580 135.750 ;
        RECT 94.230 135.150 95.230 135.600 ;
        RECT 90.880 135.000 98.580 135.150 ;
        RECT 94.230 134.550 95.230 135.000 ;
        RECT 90.880 134.400 98.580 134.550 ;
        RECT 94.230 133.950 95.230 134.400 ;
        RECT 90.880 133.800 98.580 133.950 ;
        RECT 94.230 133.350 95.230 133.800 ;
        RECT 90.880 133.200 98.580 133.350 ;
        RECT 94.230 132.750 95.230 133.200 ;
        RECT 90.880 132.600 98.580 132.750 ;
        RECT 94.230 132.150 95.230 132.600 ;
        RECT 90.880 132.000 98.580 132.150 ;
        RECT 94.230 131.550 95.230 132.000 ;
        RECT 90.880 131.400 98.580 131.550 ;
        RECT 94.230 130.950 95.230 131.400 ;
        RECT 90.880 130.800 98.580 130.950 ;
        RECT 94.230 130.300 95.230 130.800 ;
        RECT 99.480 130.300 99.630 137.850 ;
        RECT 100.080 130.300 100.230 137.850 ;
        RECT 100.680 130.300 100.830 137.850 ;
        RECT 101.280 130.300 101.430 137.850 ;
        RECT 101.880 130.300 102.030 137.850 ;
        RECT 102.480 130.300 102.630 137.850 ;
        RECT 102.780 133.200 103.530 135.000 ;
        RECT 102.780 130.450 104.730 133.200 ;
        RECT 102.780 130.300 103.930 130.450 ;
        RECT 85.530 129.700 103.930 130.300 ;
        RECT 85.530 129.550 86.680 129.700 ;
        RECT 82.780 126.800 86.680 129.550 ;
        RECT 82.780 125.050 83.530 126.800 ;
        RECT 85.930 125.050 86.680 126.800 ;
        RECT 86.830 122.150 86.980 129.700 ;
        RECT 87.430 122.150 87.580 129.700 ;
        RECT 88.030 122.150 88.180 129.700 ;
        RECT 88.630 122.150 88.780 129.700 ;
        RECT 89.230 122.150 89.380 129.700 ;
        RECT 89.830 122.150 89.980 129.700 ;
        RECT 94.230 129.200 95.230 129.700 ;
        RECT 90.880 129.050 98.580 129.200 ;
        RECT 94.230 128.600 95.230 129.050 ;
        RECT 90.880 128.450 98.580 128.600 ;
        RECT 94.230 128.000 95.230 128.450 ;
        RECT 90.880 127.850 98.580 128.000 ;
        RECT 94.230 127.400 95.230 127.850 ;
        RECT 90.880 127.250 98.580 127.400 ;
        RECT 94.230 126.800 95.230 127.250 ;
        RECT 90.880 126.650 98.580 126.800 ;
        RECT 94.230 126.200 95.230 126.650 ;
        RECT 90.880 126.050 98.580 126.200 ;
        RECT 94.230 125.600 95.230 126.050 ;
        RECT 90.880 125.450 98.580 125.600 ;
        RECT 94.230 125.000 95.230 125.450 ;
        RECT 90.880 124.850 98.580 125.000 ;
        RECT 94.230 124.400 95.230 124.850 ;
        RECT 90.880 124.250 98.580 124.400 ;
        RECT 94.230 123.800 95.230 124.250 ;
        RECT 90.880 123.650 98.580 123.800 ;
        RECT 94.230 123.200 95.230 123.650 ;
        RECT 90.880 123.050 98.580 123.200 ;
        RECT 94.230 122.600 95.230 123.050 ;
        RECT 90.880 122.450 98.580 122.600 ;
        RECT 94.230 122.000 95.230 122.450 ;
        RECT 99.480 122.150 99.630 129.700 ;
        RECT 100.080 122.150 100.230 129.700 ;
        RECT 100.680 122.150 100.830 129.700 ;
        RECT 101.280 122.150 101.430 129.700 ;
        RECT 101.880 122.150 102.030 129.700 ;
        RECT 102.480 122.150 102.630 129.700 ;
        RECT 102.780 129.550 103.930 129.700 ;
        RECT 104.580 129.980 104.730 130.450 ;
        RECT 104.580 129.550 111.850 129.980 ;
        RECT 102.780 128.705 111.850 129.550 ;
        RECT 102.780 126.800 104.730 128.705 ;
        RECT 102.780 125.050 103.530 126.800 ;
        RECT 10.880 121.850 18.580 122.000 ;
        RECT 30.880 121.850 38.580 122.000 ;
        RECT 50.880 121.850 58.580 122.000 ;
        RECT 70.880 121.850 78.580 122.000 ;
        RECT 90.880 121.850 98.580 122.000 ;
        RECT 14.230 121.200 15.230 121.850 ;
        RECT 34.230 121.200 35.230 121.850 ;
        RECT 54.230 121.200 55.230 121.850 ;
        RECT 74.230 121.200 75.230 121.850 ;
        RECT 94.230 121.200 95.230 121.850 ;
        RECT 11.530 118.800 17.930 121.200 ;
        RECT 31.530 118.800 37.930 121.200 ;
        RECT 51.530 118.800 57.930 121.200 ;
        RECT 71.530 118.800 77.930 121.200 ;
        RECT 91.530 118.800 97.930 121.200 ;
        RECT 14.230 118.150 15.230 118.800 ;
        RECT 34.230 118.150 35.230 118.800 ;
        RECT 54.230 118.150 55.230 118.800 ;
        RECT 74.230 118.150 75.230 118.800 ;
        RECT 94.230 118.150 95.230 118.800 ;
        RECT 10.880 118.000 18.580 118.150 ;
        RECT 30.880 118.000 38.580 118.150 ;
        RECT 50.880 118.000 58.580 118.150 ;
        RECT 70.880 118.000 78.580 118.150 ;
        RECT 90.880 118.000 98.580 118.150 ;
        RECT 5.930 113.200 6.680 115.000 ;
        RECT 4.730 110.450 6.680 113.200 ;
        RECT 4.730 109.550 4.880 110.450 ;
        RECT 5.530 110.300 6.680 110.450 ;
        RECT 6.830 110.300 6.980 117.850 ;
        RECT 7.430 110.300 7.580 117.850 ;
        RECT 8.030 110.300 8.180 117.850 ;
        RECT 8.630 110.300 8.780 117.850 ;
        RECT 9.230 110.300 9.380 117.850 ;
        RECT 9.830 110.300 9.980 117.850 ;
        RECT 14.230 117.550 15.230 118.000 ;
        RECT 10.880 117.400 18.580 117.550 ;
        RECT 14.230 116.950 15.230 117.400 ;
        RECT 10.880 116.800 18.580 116.950 ;
        RECT 14.230 116.350 15.230 116.800 ;
        RECT 10.880 116.200 18.580 116.350 ;
        RECT 14.230 115.750 15.230 116.200 ;
        RECT 10.880 115.600 18.580 115.750 ;
        RECT 14.230 115.150 15.230 115.600 ;
        RECT 10.880 115.000 18.580 115.150 ;
        RECT 14.230 114.550 15.230 115.000 ;
        RECT 10.880 114.400 18.580 114.550 ;
        RECT 14.230 113.950 15.230 114.400 ;
        RECT 10.880 113.800 18.580 113.950 ;
        RECT 14.230 113.350 15.230 113.800 ;
        RECT 10.880 113.200 18.580 113.350 ;
        RECT 14.230 112.750 15.230 113.200 ;
        RECT 10.880 112.600 18.580 112.750 ;
        RECT 14.230 112.150 15.230 112.600 ;
        RECT 10.880 112.000 18.580 112.150 ;
        RECT 14.230 111.550 15.230 112.000 ;
        RECT 10.880 111.400 18.580 111.550 ;
        RECT 14.230 110.950 15.230 111.400 ;
        RECT 10.880 110.800 18.580 110.950 ;
        RECT 14.230 110.300 15.230 110.800 ;
        RECT 19.480 110.300 19.630 117.850 ;
        RECT 20.080 110.300 20.230 117.850 ;
        RECT 20.680 110.300 20.830 117.850 ;
        RECT 21.280 110.300 21.430 117.850 ;
        RECT 21.880 110.300 22.030 117.850 ;
        RECT 22.480 110.300 22.630 117.850 ;
        RECT 22.780 113.200 23.530 115.000 ;
        RECT 25.930 113.200 26.680 115.000 ;
        RECT 22.780 110.450 26.680 113.200 ;
        RECT 22.780 110.300 23.930 110.450 ;
        RECT 5.530 109.700 23.930 110.300 ;
        RECT 5.530 109.550 6.680 109.700 ;
        RECT 4.730 106.800 6.680 109.550 ;
        RECT 5.930 105.050 6.680 106.800 ;
        RECT 6.830 102.150 6.980 109.700 ;
        RECT 7.430 102.150 7.580 109.700 ;
        RECT 8.030 102.150 8.180 109.700 ;
        RECT 8.630 102.150 8.780 109.700 ;
        RECT 9.230 102.150 9.380 109.700 ;
        RECT 9.830 102.150 9.980 109.700 ;
        RECT 14.230 109.200 15.230 109.700 ;
        RECT 10.880 109.050 18.580 109.200 ;
        RECT 14.230 108.600 15.230 109.050 ;
        RECT 10.880 108.450 18.580 108.600 ;
        RECT 14.230 108.000 15.230 108.450 ;
        RECT 10.880 107.850 18.580 108.000 ;
        RECT 14.230 107.400 15.230 107.850 ;
        RECT 10.880 107.250 18.580 107.400 ;
        RECT 14.230 106.800 15.230 107.250 ;
        RECT 10.880 106.650 18.580 106.800 ;
        RECT 14.230 106.200 15.230 106.650 ;
        RECT 10.880 106.050 18.580 106.200 ;
        RECT 14.230 105.600 15.230 106.050 ;
        RECT 10.880 105.450 18.580 105.600 ;
        RECT 14.230 105.000 15.230 105.450 ;
        RECT 10.880 104.850 18.580 105.000 ;
        RECT 14.230 104.400 15.230 104.850 ;
        RECT 10.880 104.250 18.580 104.400 ;
        RECT 14.230 103.800 15.230 104.250 ;
        RECT 10.880 103.650 18.580 103.800 ;
        RECT 14.230 103.200 15.230 103.650 ;
        RECT 10.880 103.050 18.580 103.200 ;
        RECT 14.230 102.600 15.230 103.050 ;
        RECT 10.880 102.450 18.580 102.600 ;
        RECT 14.230 102.000 15.230 102.450 ;
        RECT 19.480 102.150 19.630 109.700 ;
        RECT 20.080 102.150 20.230 109.700 ;
        RECT 20.680 102.150 20.830 109.700 ;
        RECT 21.280 102.150 21.430 109.700 ;
        RECT 21.880 102.150 22.030 109.700 ;
        RECT 22.480 102.150 22.630 109.700 ;
        RECT 22.780 109.550 23.930 109.700 ;
        RECT 24.580 109.550 24.880 110.450 ;
        RECT 25.530 110.300 26.680 110.450 ;
        RECT 26.830 110.300 26.980 117.850 ;
        RECT 27.430 110.300 27.580 117.850 ;
        RECT 28.030 110.300 28.180 117.850 ;
        RECT 28.630 110.300 28.780 117.850 ;
        RECT 29.230 110.300 29.380 117.850 ;
        RECT 29.830 110.300 29.980 117.850 ;
        RECT 34.230 117.550 35.230 118.000 ;
        RECT 30.880 117.400 38.580 117.550 ;
        RECT 34.230 116.950 35.230 117.400 ;
        RECT 30.880 116.800 38.580 116.950 ;
        RECT 34.230 116.350 35.230 116.800 ;
        RECT 30.880 116.200 38.580 116.350 ;
        RECT 34.230 115.750 35.230 116.200 ;
        RECT 30.880 115.600 38.580 115.750 ;
        RECT 34.230 115.150 35.230 115.600 ;
        RECT 30.880 115.000 38.580 115.150 ;
        RECT 34.230 114.550 35.230 115.000 ;
        RECT 30.880 114.400 38.580 114.550 ;
        RECT 34.230 113.950 35.230 114.400 ;
        RECT 30.880 113.800 38.580 113.950 ;
        RECT 34.230 113.350 35.230 113.800 ;
        RECT 30.880 113.200 38.580 113.350 ;
        RECT 34.230 112.750 35.230 113.200 ;
        RECT 30.880 112.600 38.580 112.750 ;
        RECT 34.230 112.150 35.230 112.600 ;
        RECT 30.880 112.000 38.580 112.150 ;
        RECT 34.230 111.550 35.230 112.000 ;
        RECT 30.880 111.400 38.580 111.550 ;
        RECT 34.230 110.950 35.230 111.400 ;
        RECT 30.880 110.800 38.580 110.950 ;
        RECT 34.230 110.300 35.230 110.800 ;
        RECT 39.480 110.300 39.630 117.850 ;
        RECT 40.080 110.300 40.230 117.850 ;
        RECT 40.680 110.300 40.830 117.850 ;
        RECT 41.280 110.300 41.430 117.850 ;
        RECT 41.880 110.300 42.030 117.850 ;
        RECT 42.480 110.300 42.630 117.850 ;
        RECT 42.780 113.200 43.530 115.000 ;
        RECT 45.930 113.200 46.680 115.000 ;
        RECT 42.780 110.450 46.680 113.200 ;
        RECT 42.780 110.300 43.930 110.450 ;
        RECT 25.530 109.700 43.930 110.300 ;
        RECT 25.530 109.550 26.680 109.700 ;
        RECT 22.780 106.800 26.680 109.550 ;
        RECT 22.780 105.050 23.530 106.800 ;
        RECT 25.930 105.050 26.680 106.800 ;
        RECT 26.830 102.150 26.980 109.700 ;
        RECT 27.430 102.150 27.580 109.700 ;
        RECT 28.030 102.150 28.180 109.700 ;
        RECT 28.630 102.150 28.780 109.700 ;
        RECT 29.230 102.150 29.380 109.700 ;
        RECT 29.830 102.150 29.980 109.700 ;
        RECT 34.230 109.200 35.230 109.700 ;
        RECT 30.880 109.050 38.580 109.200 ;
        RECT 34.230 108.600 35.230 109.050 ;
        RECT 30.880 108.450 38.580 108.600 ;
        RECT 34.230 108.000 35.230 108.450 ;
        RECT 30.880 107.850 38.580 108.000 ;
        RECT 34.230 107.400 35.230 107.850 ;
        RECT 30.880 107.250 38.580 107.400 ;
        RECT 34.230 106.800 35.230 107.250 ;
        RECT 30.880 106.650 38.580 106.800 ;
        RECT 34.230 106.200 35.230 106.650 ;
        RECT 30.880 106.050 38.580 106.200 ;
        RECT 34.230 105.600 35.230 106.050 ;
        RECT 30.880 105.450 38.580 105.600 ;
        RECT 34.230 105.000 35.230 105.450 ;
        RECT 30.880 104.850 38.580 105.000 ;
        RECT 34.230 104.400 35.230 104.850 ;
        RECT 30.880 104.250 38.580 104.400 ;
        RECT 34.230 103.800 35.230 104.250 ;
        RECT 30.880 103.650 38.580 103.800 ;
        RECT 34.230 103.200 35.230 103.650 ;
        RECT 30.880 103.050 38.580 103.200 ;
        RECT 34.230 102.600 35.230 103.050 ;
        RECT 30.880 102.450 38.580 102.600 ;
        RECT 34.230 102.000 35.230 102.450 ;
        RECT 39.480 102.150 39.630 109.700 ;
        RECT 40.080 102.150 40.230 109.700 ;
        RECT 40.680 102.150 40.830 109.700 ;
        RECT 41.280 102.150 41.430 109.700 ;
        RECT 41.880 102.150 42.030 109.700 ;
        RECT 42.480 102.150 42.630 109.700 ;
        RECT 42.780 109.550 43.930 109.700 ;
        RECT 44.580 109.550 44.880 110.450 ;
        RECT 45.530 110.300 46.680 110.450 ;
        RECT 46.830 110.300 46.980 117.850 ;
        RECT 47.430 110.300 47.580 117.850 ;
        RECT 48.030 110.300 48.180 117.850 ;
        RECT 48.630 110.300 48.780 117.850 ;
        RECT 49.230 110.300 49.380 117.850 ;
        RECT 49.830 110.300 49.980 117.850 ;
        RECT 54.230 117.550 55.230 118.000 ;
        RECT 50.880 117.400 58.580 117.550 ;
        RECT 54.230 116.950 55.230 117.400 ;
        RECT 50.880 116.800 58.580 116.950 ;
        RECT 54.230 116.350 55.230 116.800 ;
        RECT 50.880 116.200 58.580 116.350 ;
        RECT 54.230 115.750 55.230 116.200 ;
        RECT 50.880 115.600 58.580 115.750 ;
        RECT 54.230 115.150 55.230 115.600 ;
        RECT 50.880 115.000 58.580 115.150 ;
        RECT 54.230 114.550 55.230 115.000 ;
        RECT 50.880 114.400 58.580 114.550 ;
        RECT 54.230 113.950 55.230 114.400 ;
        RECT 50.880 113.800 58.580 113.950 ;
        RECT 54.230 113.350 55.230 113.800 ;
        RECT 50.880 113.200 58.580 113.350 ;
        RECT 54.230 112.750 55.230 113.200 ;
        RECT 50.880 112.600 58.580 112.750 ;
        RECT 54.230 112.150 55.230 112.600 ;
        RECT 50.880 112.000 58.580 112.150 ;
        RECT 54.230 111.550 55.230 112.000 ;
        RECT 50.880 111.400 58.580 111.550 ;
        RECT 54.230 110.950 55.230 111.400 ;
        RECT 50.880 110.800 58.580 110.950 ;
        RECT 54.230 110.300 55.230 110.800 ;
        RECT 59.480 110.300 59.630 117.850 ;
        RECT 60.080 110.300 60.230 117.850 ;
        RECT 60.680 110.300 60.830 117.850 ;
        RECT 61.280 110.300 61.430 117.850 ;
        RECT 61.880 110.300 62.030 117.850 ;
        RECT 62.480 110.300 62.630 117.850 ;
        RECT 62.780 113.200 63.530 115.000 ;
        RECT 65.930 113.200 66.680 115.000 ;
        RECT 62.780 110.450 66.680 113.200 ;
        RECT 62.780 110.300 63.930 110.450 ;
        RECT 45.530 109.700 63.930 110.300 ;
        RECT 45.530 109.550 46.680 109.700 ;
        RECT 42.780 106.800 46.680 109.550 ;
        RECT 42.780 105.050 43.530 106.800 ;
        RECT 45.930 105.050 46.680 106.800 ;
        RECT 46.830 102.150 46.980 109.700 ;
        RECT 47.430 102.150 47.580 109.700 ;
        RECT 48.030 102.150 48.180 109.700 ;
        RECT 48.630 102.150 48.780 109.700 ;
        RECT 49.230 102.150 49.380 109.700 ;
        RECT 49.830 102.150 49.980 109.700 ;
        RECT 54.230 109.200 55.230 109.700 ;
        RECT 50.880 109.050 58.580 109.200 ;
        RECT 54.230 108.600 55.230 109.050 ;
        RECT 50.880 108.450 58.580 108.600 ;
        RECT 54.230 108.000 55.230 108.450 ;
        RECT 50.880 107.850 58.580 108.000 ;
        RECT 54.230 107.400 55.230 107.850 ;
        RECT 50.880 107.250 58.580 107.400 ;
        RECT 54.230 106.800 55.230 107.250 ;
        RECT 50.880 106.650 58.580 106.800 ;
        RECT 54.230 106.200 55.230 106.650 ;
        RECT 50.880 106.050 58.580 106.200 ;
        RECT 54.230 105.600 55.230 106.050 ;
        RECT 50.880 105.450 58.580 105.600 ;
        RECT 54.230 105.000 55.230 105.450 ;
        RECT 50.880 104.850 58.580 105.000 ;
        RECT 54.230 104.400 55.230 104.850 ;
        RECT 50.880 104.250 58.580 104.400 ;
        RECT 54.230 103.800 55.230 104.250 ;
        RECT 50.880 103.650 58.580 103.800 ;
        RECT 54.230 103.200 55.230 103.650 ;
        RECT 50.880 103.050 58.580 103.200 ;
        RECT 54.230 102.600 55.230 103.050 ;
        RECT 50.880 102.450 58.580 102.600 ;
        RECT 54.230 102.000 55.230 102.450 ;
        RECT 59.480 102.150 59.630 109.700 ;
        RECT 60.080 102.150 60.230 109.700 ;
        RECT 60.680 102.150 60.830 109.700 ;
        RECT 61.280 102.150 61.430 109.700 ;
        RECT 61.880 102.150 62.030 109.700 ;
        RECT 62.480 102.150 62.630 109.700 ;
        RECT 62.780 109.550 63.930 109.700 ;
        RECT 64.580 109.550 64.880 110.450 ;
        RECT 65.530 110.300 66.680 110.450 ;
        RECT 66.830 110.300 66.980 117.850 ;
        RECT 67.430 110.300 67.580 117.850 ;
        RECT 68.030 110.300 68.180 117.850 ;
        RECT 68.630 110.300 68.780 117.850 ;
        RECT 69.230 110.300 69.380 117.850 ;
        RECT 69.830 110.300 69.980 117.850 ;
        RECT 74.230 117.550 75.230 118.000 ;
        RECT 70.880 117.400 78.580 117.550 ;
        RECT 74.230 116.950 75.230 117.400 ;
        RECT 70.880 116.800 78.580 116.950 ;
        RECT 74.230 116.350 75.230 116.800 ;
        RECT 70.880 116.200 78.580 116.350 ;
        RECT 74.230 115.750 75.230 116.200 ;
        RECT 70.880 115.600 78.580 115.750 ;
        RECT 74.230 115.150 75.230 115.600 ;
        RECT 70.880 115.000 78.580 115.150 ;
        RECT 74.230 114.550 75.230 115.000 ;
        RECT 70.880 114.400 78.580 114.550 ;
        RECT 74.230 113.950 75.230 114.400 ;
        RECT 70.880 113.800 78.580 113.950 ;
        RECT 74.230 113.350 75.230 113.800 ;
        RECT 70.880 113.200 78.580 113.350 ;
        RECT 74.230 112.750 75.230 113.200 ;
        RECT 70.880 112.600 78.580 112.750 ;
        RECT 74.230 112.150 75.230 112.600 ;
        RECT 70.880 112.000 78.580 112.150 ;
        RECT 74.230 111.550 75.230 112.000 ;
        RECT 70.880 111.400 78.580 111.550 ;
        RECT 74.230 110.950 75.230 111.400 ;
        RECT 70.880 110.800 78.580 110.950 ;
        RECT 74.230 110.300 75.230 110.800 ;
        RECT 79.480 110.300 79.630 117.850 ;
        RECT 80.080 110.300 80.230 117.850 ;
        RECT 80.680 110.300 80.830 117.850 ;
        RECT 81.280 110.300 81.430 117.850 ;
        RECT 81.880 110.300 82.030 117.850 ;
        RECT 82.480 110.300 82.630 117.850 ;
        RECT 82.780 113.200 83.530 115.000 ;
        RECT 85.930 113.200 86.680 115.000 ;
        RECT 82.780 110.450 86.680 113.200 ;
        RECT 82.780 110.300 83.930 110.450 ;
        RECT 65.530 109.700 83.930 110.300 ;
        RECT 65.530 109.550 66.680 109.700 ;
        RECT 62.780 106.800 66.680 109.550 ;
        RECT 62.780 105.050 63.530 106.800 ;
        RECT 65.930 105.050 66.680 106.800 ;
        RECT 66.830 102.150 66.980 109.700 ;
        RECT 67.430 102.150 67.580 109.700 ;
        RECT 68.030 102.150 68.180 109.700 ;
        RECT 68.630 102.150 68.780 109.700 ;
        RECT 69.230 102.150 69.380 109.700 ;
        RECT 69.830 102.150 69.980 109.700 ;
        RECT 74.230 109.200 75.230 109.700 ;
        RECT 70.880 109.050 78.580 109.200 ;
        RECT 74.230 108.600 75.230 109.050 ;
        RECT 70.880 108.450 78.580 108.600 ;
        RECT 74.230 108.000 75.230 108.450 ;
        RECT 70.880 107.850 78.580 108.000 ;
        RECT 74.230 107.400 75.230 107.850 ;
        RECT 70.880 107.250 78.580 107.400 ;
        RECT 74.230 106.800 75.230 107.250 ;
        RECT 70.880 106.650 78.580 106.800 ;
        RECT 74.230 106.200 75.230 106.650 ;
        RECT 70.880 106.050 78.580 106.200 ;
        RECT 74.230 105.600 75.230 106.050 ;
        RECT 70.880 105.450 78.580 105.600 ;
        RECT 74.230 105.000 75.230 105.450 ;
        RECT 70.880 104.850 78.580 105.000 ;
        RECT 74.230 104.400 75.230 104.850 ;
        RECT 70.880 104.250 78.580 104.400 ;
        RECT 74.230 103.800 75.230 104.250 ;
        RECT 70.880 103.650 78.580 103.800 ;
        RECT 74.230 103.200 75.230 103.650 ;
        RECT 70.880 103.050 78.580 103.200 ;
        RECT 74.230 102.600 75.230 103.050 ;
        RECT 70.880 102.450 78.580 102.600 ;
        RECT 74.230 102.000 75.230 102.450 ;
        RECT 79.480 102.150 79.630 109.700 ;
        RECT 80.080 102.150 80.230 109.700 ;
        RECT 80.680 102.150 80.830 109.700 ;
        RECT 81.280 102.150 81.430 109.700 ;
        RECT 81.880 102.150 82.030 109.700 ;
        RECT 82.480 102.150 82.630 109.700 ;
        RECT 82.780 109.550 83.930 109.700 ;
        RECT 84.580 109.550 84.880 110.450 ;
        RECT 85.530 110.300 86.680 110.450 ;
        RECT 86.830 110.300 86.980 117.850 ;
        RECT 87.430 110.300 87.580 117.850 ;
        RECT 88.030 110.300 88.180 117.850 ;
        RECT 88.630 110.300 88.780 117.850 ;
        RECT 89.230 110.300 89.380 117.850 ;
        RECT 89.830 110.300 89.980 117.850 ;
        RECT 94.230 117.550 95.230 118.000 ;
        RECT 90.880 117.400 98.580 117.550 ;
        RECT 94.230 116.950 95.230 117.400 ;
        RECT 90.880 116.800 98.580 116.950 ;
        RECT 94.230 116.350 95.230 116.800 ;
        RECT 90.880 116.200 98.580 116.350 ;
        RECT 94.230 115.750 95.230 116.200 ;
        RECT 90.880 115.600 98.580 115.750 ;
        RECT 94.230 115.150 95.230 115.600 ;
        RECT 90.880 115.000 98.580 115.150 ;
        RECT 94.230 114.550 95.230 115.000 ;
        RECT 90.880 114.400 98.580 114.550 ;
        RECT 94.230 113.950 95.230 114.400 ;
        RECT 90.880 113.800 98.580 113.950 ;
        RECT 94.230 113.350 95.230 113.800 ;
        RECT 90.880 113.200 98.580 113.350 ;
        RECT 94.230 112.750 95.230 113.200 ;
        RECT 90.880 112.600 98.580 112.750 ;
        RECT 94.230 112.150 95.230 112.600 ;
        RECT 90.880 112.000 98.580 112.150 ;
        RECT 94.230 111.550 95.230 112.000 ;
        RECT 90.880 111.400 98.580 111.550 ;
        RECT 94.230 110.950 95.230 111.400 ;
        RECT 90.880 110.800 98.580 110.950 ;
        RECT 94.230 110.300 95.230 110.800 ;
        RECT 99.480 110.300 99.630 117.850 ;
        RECT 100.080 110.300 100.230 117.850 ;
        RECT 100.680 110.300 100.830 117.850 ;
        RECT 101.280 110.300 101.430 117.850 ;
        RECT 101.880 110.300 102.030 117.850 ;
        RECT 102.480 110.300 102.630 117.850 ;
        RECT 102.780 113.200 103.530 115.000 ;
        RECT 102.780 111.030 104.730 113.200 ;
        RECT 102.780 110.450 111.850 111.030 ;
        RECT 102.780 110.300 103.930 110.450 ;
        RECT 85.530 109.700 103.930 110.300 ;
        RECT 85.530 109.550 86.680 109.700 ;
        RECT 82.780 106.800 86.680 109.550 ;
        RECT 82.780 105.050 83.530 106.800 ;
        RECT 85.930 105.050 86.680 106.800 ;
        RECT 86.830 102.150 86.980 109.700 ;
        RECT 87.430 102.150 87.580 109.700 ;
        RECT 88.030 102.150 88.180 109.700 ;
        RECT 88.630 102.150 88.780 109.700 ;
        RECT 89.230 102.150 89.380 109.700 ;
        RECT 89.830 102.150 89.980 109.700 ;
        RECT 94.230 109.200 95.230 109.700 ;
        RECT 90.880 109.050 98.580 109.200 ;
        RECT 94.230 108.600 95.230 109.050 ;
        RECT 90.880 108.450 98.580 108.600 ;
        RECT 94.230 108.000 95.230 108.450 ;
        RECT 90.880 107.850 98.580 108.000 ;
        RECT 94.230 107.400 95.230 107.850 ;
        RECT 90.880 107.250 98.580 107.400 ;
        RECT 94.230 106.800 95.230 107.250 ;
        RECT 90.880 106.650 98.580 106.800 ;
        RECT 94.230 106.200 95.230 106.650 ;
        RECT 90.880 106.050 98.580 106.200 ;
        RECT 94.230 105.600 95.230 106.050 ;
        RECT 90.880 105.450 98.580 105.600 ;
        RECT 94.230 105.000 95.230 105.450 ;
        RECT 90.880 104.850 98.580 105.000 ;
        RECT 94.230 104.400 95.230 104.850 ;
        RECT 90.880 104.250 98.580 104.400 ;
        RECT 94.230 103.800 95.230 104.250 ;
        RECT 90.880 103.650 98.580 103.800 ;
        RECT 94.230 103.200 95.230 103.650 ;
        RECT 90.880 103.050 98.580 103.200 ;
        RECT 94.230 102.600 95.230 103.050 ;
        RECT 90.880 102.450 98.580 102.600 ;
        RECT 94.230 102.000 95.230 102.450 ;
        RECT 99.480 102.150 99.630 109.700 ;
        RECT 100.080 102.150 100.230 109.700 ;
        RECT 100.680 102.150 100.830 109.700 ;
        RECT 101.280 102.150 101.430 109.700 ;
        RECT 101.880 102.150 102.030 109.700 ;
        RECT 102.480 102.150 102.630 109.700 ;
        RECT 102.780 109.550 103.930 109.700 ;
        RECT 104.580 109.755 111.850 110.450 ;
        RECT 104.580 109.550 104.730 109.755 ;
        RECT 102.780 106.800 104.730 109.550 ;
        RECT 102.780 105.050 103.530 106.800 ;
        RECT 10.880 101.850 18.580 102.000 ;
        RECT 30.880 101.850 38.580 102.000 ;
        RECT 50.880 101.850 58.580 102.000 ;
        RECT 70.880 101.850 78.580 102.000 ;
        RECT 90.880 101.850 98.580 102.000 ;
        RECT 14.230 101.200 15.230 101.850 ;
        RECT 34.230 101.200 35.230 101.850 ;
        RECT 54.230 101.200 55.230 101.850 ;
        RECT 74.230 101.200 75.230 101.850 ;
        RECT 94.230 101.200 95.230 101.850 ;
        RECT 11.530 98.800 17.930 101.200 ;
        RECT 31.530 98.800 37.930 101.200 ;
        RECT 51.530 98.800 57.930 101.200 ;
        RECT 71.530 98.800 77.930 101.200 ;
        RECT 91.530 98.800 97.930 101.200 ;
        RECT 14.230 98.150 15.230 98.800 ;
        RECT 34.230 98.150 35.230 98.800 ;
        RECT 54.230 98.150 55.230 98.800 ;
        RECT 74.230 98.150 75.230 98.800 ;
        RECT 94.230 98.150 95.230 98.800 ;
        RECT 10.880 98.000 18.580 98.150 ;
        RECT 30.880 98.000 38.580 98.150 ;
        RECT 50.880 98.000 58.580 98.150 ;
        RECT 70.880 98.000 78.580 98.150 ;
        RECT 90.880 98.000 98.580 98.150 ;
        RECT 5.930 93.200 6.680 95.000 ;
        RECT 4.730 90.450 6.680 93.200 ;
        RECT 4.730 89.550 4.880 90.450 ;
        RECT 5.530 90.300 6.680 90.450 ;
        RECT 6.830 90.300 6.980 97.850 ;
        RECT 7.430 90.300 7.580 97.850 ;
        RECT 8.030 90.300 8.180 97.850 ;
        RECT 8.630 90.300 8.780 97.850 ;
        RECT 9.230 90.300 9.380 97.850 ;
        RECT 9.830 90.300 9.980 97.850 ;
        RECT 14.230 97.550 15.230 98.000 ;
        RECT 10.880 97.400 18.580 97.550 ;
        RECT 14.230 96.950 15.230 97.400 ;
        RECT 10.880 96.800 18.580 96.950 ;
        RECT 14.230 96.350 15.230 96.800 ;
        RECT 10.880 96.200 18.580 96.350 ;
        RECT 14.230 95.750 15.230 96.200 ;
        RECT 10.880 95.600 18.580 95.750 ;
        RECT 14.230 95.150 15.230 95.600 ;
        RECT 10.880 95.000 18.580 95.150 ;
        RECT 14.230 94.550 15.230 95.000 ;
        RECT 10.880 94.400 18.580 94.550 ;
        RECT 14.230 93.950 15.230 94.400 ;
        RECT 10.880 93.800 18.580 93.950 ;
        RECT 14.230 93.350 15.230 93.800 ;
        RECT 10.880 93.200 18.580 93.350 ;
        RECT 14.230 92.750 15.230 93.200 ;
        RECT 10.880 92.600 18.580 92.750 ;
        RECT 14.230 92.150 15.230 92.600 ;
        RECT 10.880 92.000 18.580 92.150 ;
        RECT 14.230 91.550 15.230 92.000 ;
        RECT 10.880 91.400 18.580 91.550 ;
        RECT 14.230 90.950 15.230 91.400 ;
        RECT 10.880 90.800 18.580 90.950 ;
        RECT 14.230 90.300 15.230 90.800 ;
        RECT 19.480 90.300 19.630 97.850 ;
        RECT 20.080 90.300 20.230 97.850 ;
        RECT 20.680 90.300 20.830 97.850 ;
        RECT 21.280 90.300 21.430 97.850 ;
        RECT 21.880 90.300 22.030 97.850 ;
        RECT 22.480 90.300 22.630 97.850 ;
        RECT 22.780 93.200 23.530 95.000 ;
        RECT 25.930 93.200 26.680 95.000 ;
        RECT 22.780 90.450 26.680 93.200 ;
        RECT 22.780 90.300 23.930 90.450 ;
        RECT 5.530 89.700 23.930 90.300 ;
        RECT 5.530 89.550 6.680 89.700 ;
        RECT 4.730 86.800 6.680 89.550 ;
        RECT 5.930 85.050 6.680 86.800 ;
        RECT 6.830 82.150 6.980 89.700 ;
        RECT 7.430 82.150 7.580 89.700 ;
        RECT 8.030 82.150 8.180 89.700 ;
        RECT 8.630 82.150 8.780 89.700 ;
        RECT 9.230 82.150 9.380 89.700 ;
        RECT 9.830 82.150 9.980 89.700 ;
        RECT 14.230 89.200 15.230 89.700 ;
        RECT 10.880 89.050 18.580 89.200 ;
        RECT 14.230 88.600 15.230 89.050 ;
        RECT 10.880 88.450 18.580 88.600 ;
        RECT 14.230 88.000 15.230 88.450 ;
        RECT 10.880 87.850 18.580 88.000 ;
        RECT 14.230 87.400 15.230 87.850 ;
        RECT 10.880 87.250 18.580 87.400 ;
        RECT 14.230 86.800 15.230 87.250 ;
        RECT 10.880 86.650 18.580 86.800 ;
        RECT 14.230 86.200 15.230 86.650 ;
        RECT 10.880 86.050 18.580 86.200 ;
        RECT 14.230 85.600 15.230 86.050 ;
        RECT 10.880 85.450 18.580 85.600 ;
        RECT 14.230 85.000 15.230 85.450 ;
        RECT 10.880 84.850 18.580 85.000 ;
        RECT 14.230 84.400 15.230 84.850 ;
        RECT 10.880 84.250 18.580 84.400 ;
        RECT 14.230 83.800 15.230 84.250 ;
        RECT 10.880 83.650 18.580 83.800 ;
        RECT 14.230 83.200 15.230 83.650 ;
        RECT 10.880 83.050 18.580 83.200 ;
        RECT 14.230 82.600 15.230 83.050 ;
        RECT 10.880 82.450 18.580 82.600 ;
        RECT 14.230 82.000 15.230 82.450 ;
        RECT 19.480 82.150 19.630 89.700 ;
        RECT 20.080 82.150 20.230 89.700 ;
        RECT 20.680 82.150 20.830 89.700 ;
        RECT 21.280 82.150 21.430 89.700 ;
        RECT 21.880 82.150 22.030 89.700 ;
        RECT 22.480 82.150 22.630 89.700 ;
        RECT 22.780 89.550 23.930 89.700 ;
        RECT 24.580 89.550 24.880 90.450 ;
        RECT 25.530 90.300 26.680 90.450 ;
        RECT 26.830 90.300 26.980 97.850 ;
        RECT 27.430 90.300 27.580 97.850 ;
        RECT 28.030 90.300 28.180 97.850 ;
        RECT 28.630 90.300 28.780 97.850 ;
        RECT 29.230 90.300 29.380 97.850 ;
        RECT 29.830 90.300 29.980 97.850 ;
        RECT 34.230 97.550 35.230 98.000 ;
        RECT 30.880 97.400 38.580 97.550 ;
        RECT 34.230 96.950 35.230 97.400 ;
        RECT 30.880 96.800 38.580 96.950 ;
        RECT 34.230 96.350 35.230 96.800 ;
        RECT 30.880 96.200 38.580 96.350 ;
        RECT 34.230 95.750 35.230 96.200 ;
        RECT 30.880 95.600 38.580 95.750 ;
        RECT 34.230 95.150 35.230 95.600 ;
        RECT 30.880 95.000 38.580 95.150 ;
        RECT 34.230 94.550 35.230 95.000 ;
        RECT 30.880 94.400 38.580 94.550 ;
        RECT 34.230 93.950 35.230 94.400 ;
        RECT 30.880 93.800 38.580 93.950 ;
        RECT 34.230 93.350 35.230 93.800 ;
        RECT 30.880 93.200 38.580 93.350 ;
        RECT 34.230 92.750 35.230 93.200 ;
        RECT 30.880 92.600 38.580 92.750 ;
        RECT 34.230 92.150 35.230 92.600 ;
        RECT 30.880 92.000 38.580 92.150 ;
        RECT 34.230 91.550 35.230 92.000 ;
        RECT 30.880 91.400 38.580 91.550 ;
        RECT 34.230 90.950 35.230 91.400 ;
        RECT 30.880 90.800 38.580 90.950 ;
        RECT 34.230 90.300 35.230 90.800 ;
        RECT 39.480 90.300 39.630 97.850 ;
        RECT 40.080 90.300 40.230 97.850 ;
        RECT 40.680 90.300 40.830 97.850 ;
        RECT 41.280 90.300 41.430 97.850 ;
        RECT 41.880 90.300 42.030 97.850 ;
        RECT 42.480 90.300 42.630 97.850 ;
        RECT 42.780 93.200 43.530 95.000 ;
        RECT 45.930 93.200 46.680 95.000 ;
        RECT 42.780 90.450 46.680 93.200 ;
        RECT 42.780 90.300 43.930 90.450 ;
        RECT 25.530 89.700 43.930 90.300 ;
        RECT 25.530 89.550 26.680 89.700 ;
        RECT 22.780 86.800 26.680 89.550 ;
        RECT 22.780 85.050 23.530 86.800 ;
        RECT 25.930 85.050 26.680 86.800 ;
        RECT 26.830 82.150 26.980 89.700 ;
        RECT 27.430 82.150 27.580 89.700 ;
        RECT 28.030 82.150 28.180 89.700 ;
        RECT 28.630 82.150 28.780 89.700 ;
        RECT 29.230 82.150 29.380 89.700 ;
        RECT 29.830 82.150 29.980 89.700 ;
        RECT 34.230 89.200 35.230 89.700 ;
        RECT 30.880 89.050 38.580 89.200 ;
        RECT 34.230 88.600 35.230 89.050 ;
        RECT 30.880 88.450 38.580 88.600 ;
        RECT 34.230 88.000 35.230 88.450 ;
        RECT 30.880 87.850 38.580 88.000 ;
        RECT 34.230 87.400 35.230 87.850 ;
        RECT 30.880 87.250 38.580 87.400 ;
        RECT 34.230 86.800 35.230 87.250 ;
        RECT 30.880 86.650 38.580 86.800 ;
        RECT 34.230 86.200 35.230 86.650 ;
        RECT 30.880 86.050 38.580 86.200 ;
        RECT 34.230 85.600 35.230 86.050 ;
        RECT 30.880 85.450 38.580 85.600 ;
        RECT 34.230 85.000 35.230 85.450 ;
        RECT 30.880 84.850 38.580 85.000 ;
        RECT 34.230 84.400 35.230 84.850 ;
        RECT 30.880 84.250 38.580 84.400 ;
        RECT 34.230 83.800 35.230 84.250 ;
        RECT 30.880 83.650 38.580 83.800 ;
        RECT 34.230 83.200 35.230 83.650 ;
        RECT 30.880 83.050 38.580 83.200 ;
        RECT 34.230 82.600 35.230 83.050 ;
        RECT 30.880 82.450 38.580 82.600 ;
        RECT 34.230 82.000 35.230 82.450 ;
        RECT 39.480 82.150 39.630 89.700 ;
        RECT 40.080 82.150 40.230 89.700 ;
        RECT 40.680 82.150 40.830 89.700 ;
        RECT 41.280 82.150 41.430 89.700 ;
        RECT 41.880 82.150 42.030 89.700 ;
        RECT 42.480 82.150 42.630 89.700 ;
        RECT 42.780 89.550 43.930 89.700 ;
        RECT 44.580 89.550 44.880 90.450 ;
        RECT 45.530 90.300 46.680 90.450 ;
        RECT 46.830 90.300 46.980 97.850 ;
        RECT 47.430 90.300 47.580 97.850 ;
        RECT 48.030 90.300 48.180 97.850 ;
        RECT 48.630 90.300 48.780 97.850 ;
        RECT 49.230 90.300 49.380 97.850 ;
        RECT 49.830 90.300 49.980 97.850 ;
        RECT 54.230 97.550 55.230 98.000 ;
        RECT 50.880 97.400 58.580 97.550 ;
        RECT 54.230 96.950 55.230 97.400 ;
        RECT 50.880 96.800 58.580 96.950 ;
        RECT 54.230 96.350 55.230 96.800 ;
        RECT 50.880 96.200 58.580 96.350 ;
        RECT 54.230 95.750 55.230 96.200 ;
        RECT 50.880 95.600 58.580 95.750 ;
        RECT 54.230 95.150 55.230 95.600 ;
        RECT 50.880 95.000 58.580 95.150 ;
        RECT 54.230 94.550 55.230 95.000 ;
        RECT 50.880 94.400 58.580 94.550 ;
        RECT 54.230 93.950 55.230 94.400 ;
        RECT 50.880 93.800 58.580 93.950 ;
        RECT 54.230 93.350 55.230 93.800 ;
        RECT 50.880 93.200 58.580 93.350 ;
        RECT 54.230 92.750 55.230 93.200 ;
        RECT 50.880 92.600 58.580 92.750 ;
        RECT 54.230 92.150 55.230 92.600 ;
        RECT 50.880 92.000 58.580 92.150 ;
        RECT 54.230 91.550 55.230 92.000 ;
        RECT 50.880 91.400 58.580 91.550 ;
        RECT 54.230 90.950 55.230 91.400 ;
        RECT 50.880 90.800 58.580 90.950 ;
        RECT 54.230 90.300 55.230 90.800 ;
        RECT 59.480 90.300 59.630 97.850 ;
        RECT 60.080 90.300 60.230 97.850 ;
        RECT 60.680 90.300 60.830 97.850 ;
        RECT 61.280 90.300 61.430 97.850 ;
        RECT 61.880 90.300 62.030 97.850 ;
        RECT 62.480 90.300 62.630 97.850 ;
        RECT 62.780 93.200 63.530 95.000 ;
        RECT 65.930 93.200 66.680 95.000 ;
        RECT 62.780 90.450 66.680 93.200 ;
        RECT 62.780 90.300 63.930 90.450 ;
        RECT 45.530 89.700 63.930 90.300 ;
        RECT 45.530 89.550 46.680 89.700 ;
        RECT 42.780 86.800 46.680 89.550 ;
        RECT 42.780 85.050 43.530 86.800 ;
        RECT 45.930 85.050 46.680 86.800 ;
        RECT 46.830 82.150 46.980 89.700 ;
        RECT 47.430 82.150 47.580 89.700 ;
        RECT 48.030 82.150 48.180 89.700 ;
        RECT 48.630 82.150 48.780 89.700 ;
        RECT 49.230 82.150 49.380 89.700 ;
        RECT 49.830 82.150 49.980 89.700 ;
        RECT 54.230 89.200 55.230 89.700 ;
        RECT 50.880 89.050 58.580 89.200 ;
        RECT 54.230 88.600 55.230 89.050 ;
        RECT 50.880 88.450 58.580 88.600 ;
        RECT 54.230 88.000 55.230 88.450 ;
        RECT 50.880 87.850 58.580 88.000 ;
        RECT 54.230 87.400 55.230 87.850 ;
        RECT 50.880 87.250 58.580 87.400 ;
        RECT 54.230 86.800 55.230 87.250 ;
        RECT 50.880 86.650 58.580 86.800 ;
        RECT 54.230 86.200 55.230 86.650 ;
        RECT 50.880 86.050 58.580 86.200 ;
        RECT 54.230 85.600 55.230 86.050 ;
        RECT 50.880 85.450 58.580 85.600 ;
        RECT 54.230 85.000 55.230 85.450 ;
        RECT 50.880 84.850 58.580 85.000 ;
        RECT 54.230 84.400 55.230 84.850 ;
        RECT 50.880 84.250 58.580 84.400 ;
        RECT 54.230 83.800 55.230 84.250 ;
        RECT 50.880 83.650 58.580 83.800 ;
        RECT 54.230 83.200 55.230 83.650 ;
        RECT 50.880 83.050 58.580 83.200 ;
        RECT 54.230 82.600 55.230 83.050 ;
        RECT 50.880 82.450 58.580 82.600 ;
        RECT 54.230 82.000 55.230 82.450 ;
        RECT 59.480 82.150 59.630 89.700 ;
        RECT 60.080 82.150 60.230 89.700 ;
        RECT 60.680 82.150 60.830 89.700 ;
        RECT 61.280 82.150 61.430 89.700 ;
        RECT 61.880 82.150 62.030 89.700 ;
        RECT 62.480 82.150 62.630 89.700 ;
        RECT 62.780 89.550 63.930 89.700 ;
        RECT 64.580 89.550 64.880 90.450 ;
        RECT 65.530 90.300 66.680 90.450 ;
        RECT 66.830 90.300 66.980 97.850 ;
        RECT 67.430 90.300 67.580 97.850 ;
        RECT 68.030 90.300 68.180 97.850 ;
        RECT 68.630 90.300 68.780 97.850 ;
        RECT 69.230 90.300 69.380 97.850 ;
        RECT 69.830 90.300 69.980 97.850 ;
        RECT 74.230 97.550 75.230 98.000 ;
        RECT 70.880 97.400 78.580 97.550 ;
        RECT 74.230 96.950 75.230 97.400 ;
        RECT 70.880 96.800 78.580 96.950 ;
        RECT 74.230 96.350 75.230 96.800 ;
        RECT 70.880 96.200 78.580 96.350 ;
        RECT 74.230 95.750 75.230 96.200 ;
        RECT 70.880 95.600 78.580 95.750 ;
        RECT 74.230 95.150 75.230 95.600 ;
        RECT 70.880 95.000 78.580 95.150 ;
        RECT 74.230 94.550 75.230 95.000 ;
        RECT 70.880 94.400 78.580 94.550 ;
        RECT 74.230 93.950 75.230 94.400 ;
        RECT 70.880 93.800 78.580 93.950 ;
        RECT 74.230 93.350 75.230 93.800 ;
        RECT 70.880 93.200 78.580 93.350 ;
        RECT 74.230 92.750 75.230 93.200 ;
        RECT 70.880 92.600 78.580 92.750 ;
        RECT 74.230 92.150 75.230 92.600 ;
        RECT 70.880 92.000 78.580 92.150 ;
        RECT 74.230 91.550 75.230 92.000 ;
        RECT 70.880 91.400 78.580 91.550 ;
        RECT 74.230 90.950 75.230 91.400 ;
        RECT 70.880 90.800 78.580 90.950 ;
        RECT 74.230 90.300 75.230 90.800 ;
        RECT 79.480 90.300 79.630 97.850 ;
        RECT 80.080 90.300 80.230 97.850 ;
        RECT 80.680 90.300 80.830 97.850 ;
        RECT 81.280 90.300 81.430 97.850 ;
        RECT 81.880 90.300 82.030 97.850 ;
        RECT 82.480 90.300 82.630 97.850 ;
        RECT 82.780 93.200 83.530 95.000 ;
        RECT 85.930 93.200 86.680 95.000 ;
        RECT 82.780 90.450 86.680 93.200 ;
        RECT 82.780 90.300 83.930 90.450 ;
        RECT 65.530 89.700 83.930 90.300 ;
        RECT 65.530 89.550 66.680 89.700 ;
        RECT 62.780 86.800 66.680 89.550 ;
        RECT 62.780 85.050 63.530 86.800 ;
        RECT 65.930 85.050 66.680 86.800 ;
        RECT 66.830 82.150 66.980 89.700 ;
        RECT 67.430 82.150 67.580 89.700 ;
        RECT 68.030 82.150 68.180 89.700 ;
        RECT 68.630 82.150 68.780 89.700 ;
        RECT 69.230 82.150 69.380 89.700 ;
        RECT 69.830 82.150 69.980 89.700 ;
        RECT 74.230 89.200 75.230 89.700 ;
        RECT 70.880 89.050 78.580 89.200 ;
        RECT 74.230 88.600 75.230 89.050 ;
        RECT 70.880 88.450 78.580 88.600 ;
        RECT 74.230 88.000 75.230 88.450 ;
        RECT 70.880 87.850 78.580 88.000 ;
        RECT 74.230 87.400 75.230 87.850 ;
        RECT 70.880 87.250 78.580 87.400 ;
        RECT 74.230 86.800 75.230 87.250 ;
        RECT 70.880 86.650 78.580 86.800 ;
        RECT 74.230 86.200 75.230 86.650 ;
        RECT 70.880 86.050 78.580 86.200 ;
        RECT 74.230 85.600 75.230 86.050 ;
        RECT 70.880 85.450 78.580 85.600 ;
        RECT 74.230 85.000 75.230 85.450 ;
        RECT 70.880 84.850 78.580 85.000 ;
        RECT 74.230 84.400 75.230 84.850 ;
        RECT 70.880 84.250 78.580 84.400 ;
        RECT 74.230 83.800 75.230 84.250 ;
        RECT 70.880 83.650 78.580 83.800 ;
        RECT 74.230 83.200 75.230 83.650 ;
        RECT 70.880 83.050 78.580 83.200 ;
        RECT 74.230 82.600 75.230 83.050 ;
        RECT 70.880 82.450 78.580 82.600 ;
        RECT 74.230 82.000 75.230 82.450 ;
        RECT 79.480 82.150 79.630 89.700 ;
        RECT 80.080 82.150 80.230 89.700 ;
        RECT 80.680 82.150 80.830 89.700 ;
        RECT 81.280 82.150 81.430 89.700 ;
        RECT 81.880 82.150 82.030 89.700 ;
        RECT 82.480 82.150 82.630 89.700 ;
        RECT 82.780 89.550 83.930 89.700 ;
        RECT 84.580 89.550 84.880 90.450 ;
        RECT 85.530 90.300 86.680 90.450 ;
        RECT 86.830 90.300 86.980 97.850 ;
        RECT 87.430 90.300 87.580 97.850 ;
        RECT 88.030 90.300 88.180 97.850 ;
        RECT 88.630 90.300 88.780 97.850 ;
        RECT 89.230 90.300 89.380 97.850 ;
        RECT 89.830 90.300 89.980 97.850 ;
        RECT 94.230 97.550 95.230 98.000 ;
        RECT 90.880 97.400 98.580 97.550 ;
        RECT 94.230 96.950 95.230 97.400 ;
        RECT 90.880 96.800 98.580 96.950 ;
        RECT 94.230 96.350 95.230 96.800 ;
        RECT 90.880 96.200 98.580 96.350 ;
        RECT 94.230 95.750 95.230 96.200 ;
        RECT 90.880 95.600 98.580 95.750 ;
        RECT 94.230 95.150 95.230 95.600 ;
        RECT 90.880 95.000 98.580 95.150 ;
        RECT 94.230 94.550 95.230 95.000 ;
        RECT 90.880 94.400 98.580 94.550 ;
        RECT 94.230 93.950 95.230 94.400 ;
        RECT 90.880 93.800 98.580 93.950 ;
        RECT 94.230 93.350 95.230 93.800 ;
        RECT 90.880 93.200 98.580 93.350 ;
        RECT 94.230 92.750 95.230 93.200 ;
        RECT 90.880 92.600 98.580 92.750 ;
        RECT 94.230 92.150 95.230 92.600 ;
        RECT 90.880 92.000 98.580 92.150 ;
        RECT 94.230 91.550 95.230 92.000 ;
        RECT 90.880 91.400 98.580 91.550 ;
        RECT 94.230 90.950 95.230 91.400 ;
        RECT 90.880 90.800 98.580 90.950 ;
        RECT 94.230 90.300 95.230 90.800 ;
        RECT 99.480 90.300 99.630 97.850 ;
        RECT 100.080 90.300 100.230 97.850 ;
        RECT 100.680 90.300 100.830 97.850 ;
        RECT 101.280 90.300 101.430 97.850 ;
        RECT 101.880 90.300 102.030 97.850 ;
        RECT 102.480 90.300 102.630 97.850 ;
        RECT 102.780 93.200 103.530 95.000 ;
        RECT 102.780 90.495 104.730 93.200 ;
        RECT 102.780 90.450 111.850 90.495 ;
        RECT 102.780 90.300 103.930 90.450 ;
        RECT 85.530 89.700 103.930 90.300 ;
        RECT 85.530 89.550 86.680 89.700 ;
        RECT 82.780 86.800 86.680 89.550 ;
        RECT 82.780 85.050 83.530 86.800 ;
        RECT 85.930 85.050 86.680 86.800 ;
        RECT 86.830 82.150 86.980 89.700 ;
        RECT 87.430 82.150 87.580 89.700 ;
        RECT 88.030 82.150 88.180 89.700 ;
        RECT 88.630 82.150 88.780 89.700 ;
        RECT 89.230 82.150 89.380 89.700 ;
        RECT 89.830 82.150 89.980 89.700 ;
        RECT 94.230 89.200 95.230 89.700 ;
        RECT 90.880 89.050 98.580 89.200 ;
        RECT 94.230 88.600 95.230 89.050 ;
        RECT 90.880 88.450 98.580 88.600 ;
        RECT 94.230 88.000 95.230 88.450 ;
        RECT 90.880 87.850 98.580 88.000 ;
        RECT 94.230 87.400 95.230 87.850 ;
        RECT 90.880 87.250 98.580 87.400 ;
        RECT 94.230 86.800 95.230 87.250 ;
        RECT 90.880 86.650 98.580 86.800 ;
        RECT 94.230 86.200 95.230 86.650 ;
        RECT 90.880 86.050 98.580 86.200 ;
        RECT 94.230 85.600 95.230 86.050 ;
        RECT 90.880 85.450 98.580 85.600 ;
        RECT 94.230 85.000 95.230 85.450 ;
        RECT 90.880 84.850 98.580 85.000 ;
        RECT 94.230 84.400 95.230 84.850 ;
        RECT 90.880 84.250 98.580 84.400 ;
        RECT 94.230 83.800 95.230 84.250 ;
        RECT 90.880 83.650 98.580 83.800 ;
        RECT 94.230 83.200 95.230 83.650 ;
        RECT 90.880 83.050 98.580 83.200 ;
        RECT 94.230 82.600 95.230 83.050 ;
        RECT 90.880 82.450 98.580 82.600 ;
        RECT 94.230 82.000 95.230 82.450 ;
        RECT 99.480 82.150 99.630 89.700 ;
        RECT 100.080 82.150 100.230 89.700 ;
        RECT 100.680 82.150 100.830 89.700 ;
        RECT 101.280 82.150 101.430 89.700 ;
        RECT 101.880 82.150 102.030 89.700 ;
        RECT 102.480 82.150 102.630 89.700 ;
        RECT 102.780 89.550 103.930 89.700 ;
        RECT 104.580 89.550 111.850 90.450 ;
        RECT 102.780 89.220 111.850 89.550 ;
        RECT 102.780 86.800 104.730 89.220 ;
        RECT 102.780 85.050 103.530 86.800 ;
        RECT 10.880 81.850 18.580 82.000 ;
        RECT 30.880 81.850 38.580 82.000 ;
        RECT 50.880 81.850 58.580 82.000 ;
        RECT 70.880 81.850 78.580 82.000 ;
        RECT 90.880 81.850 98.580 82.000 ;
        RECT 14.230 81.200 15.230 81.850 ;
        RECT 34.230 81.200 35.230 81.850 ;
        RECT 54.230 81.200 55.230 81.850 ;
        RECT 74.230 81.200 75.230 81.850 ;
        RECT 94.230 81.200 95.230 81.850 ;
        RECT 11.530 78.800 17.930 81.200 ;
        RECT 31.530 78.800 37.930 81.200 ;
        RECT 51.530 78.800 57.930 81.200 ;
        RECT 71.530 78.800 77.930 81.200 ;
        RECT 91.530 78.800 97.930 81.200 ;
        RECT 14.230 78.150 15.230 78.800 ;
        RECT 34.230 78.150 35.230 78.800 ;
        RECT 54.230 78.150 55.230 78.800 ;
        RECT 74.230 78.150 75.230 78.800 ;
        RECT 94.230 78.150 95.230 78.800 ;
        RECT 10.880 78.000 18.580 78.150 ;
        RECT 30.880 78.000 38.580 78.150 ;
        RECT 50.880 78.000 58.580 78.150 ;
        RECT 70.880 78.000 78.580 78.150 ;
        RECT 90.880 78.000 98.580 78.150 ;
        RECT 5.930 73.200 6.680 75.000 ;
        RECT 4.730 70.450 6.680 73.200 ;
        RECT 4.730 69.550 4.880 70.450 ;
        RECT 5.530 70.300 6.680 70.450 ;
        RECT 6.830 70.300 6.980 77.850 ;
        RECT 7.430 70.300 7.580 77.850 ;
        RECT 8.030 70.300 8.180 77.850 ;
        RECT 8.630 70.300 8.780 77.850 ;
        RECT 9.230 70.300 9.380 77.850 ;
        RECT 9.830 70.300 9.980 77.850 ;
        RECT 14.230 77.550 15.230 78.000 ;
        RECT 10.880 77.400 18.580 77.550 ;
        RECT 14.230 76.950 15.230 77.400 ;
        RECT 10.880 76.800 18.580 76.950 ;
        RECT 14.230 76.350 15.230 76.800 ;
        RECT 10.880 76.200 18.580 76.350 ;
        RECT 14.230 75.750 15.230 76.200 ;
        RECT 10.880 75.600 18.580 75.750 ;
        RECT 14.230 75.150 15.230 75.600 ;
        RECT 10.880 75.000 18.580 75.150 ;
        RECT 14.230 74.550 15.230 75.000 ;
        RECT 10.880 74.400 18.580 74.550 ;
        RECT 14.230 73.950 15.230 74.400 ;
        RECT 10.880 73.800 18.580 73.950 ;
        RECT 14.230 73.350 15.230 73.800 ;
        RECT 10.880 73.200 18.580 73.350 ;
        RECT 14.230 72.750 15.230 73.200 ;
        RECT 10.880 72.600 18.580 72.750 ;
        RECT 14.230 72.150 15.230 72.600 ;
        RECT 10.880 72.000 18.580 72.150 ;
        RECT 14.230 71.550 15.230 72.000 ;
        RECT 10.880 71.400 18.580 71.550 ;
        RECT 14.230 70.950 15.230 71.400 ;
        RECT 10.880 70.800 18.580 70.950 ;
        RECT 14.230 70.300 15.230 70.800 ;
        RECT 19.480 70.300 19.630 77.850 ;
        RECT 20.080 70.300 20.230 77.850 ;
        RECT 20.680 70.300 20.830 77.850 ;
        RECT 21.280 70.300 21.430 77.850 ;
        RECT 21.880 70.300 22.030 77.850 ;
        RECT 22.480 70.300 22.630 77.850 ;
        RECT 22.780 73.200 23.530 75.000 ;
        RECT 25.930 73.200 26.680 75.000 ;
        RECT 22.780 70.450 26.680 73.200 ;
        RECT 22.780 70.300 23.930 70.450 ;
        RECT 5.530 69.700 23.930 70.300 ;
        RECT 5.530 69.550 6.680 69.700 ;
        RECT 4.730 66.800 6.680 69.550 ;
        RECT 5.930 65.050 6.680 66.800 ;
        RECT 6.830 62.150 6.980 69.700 ;
        RECT 7.430 62.150 7.580 69.700 ;
        RECT 8.030 62.150 8.180 69.700 ;
        RECT 8.630 62.150 8.780 69.700 ;
        RECT 9.230 62.150 9.380 69.700 ;
        RECT 9.830 62.150 9.980 69.700 ;
        RECT 14.230 69.200 15.230 69.700 ;
        RECT 10.880 69.050 18.580 69.200 ;
        RECT 14.230 68.600 15.230 69.050 ;
        RECT 10.880 68.450 18.580 68.600 ;
        RECT 14.230 68.000 15.230 68.450 ;
        RECT 10.880 67.850 18.580 68.000 ;
        RECT 14.230 67.400 15.230 67.850 ;
        RECT 10.880 67.250 18.580 67.400 ;
        RECT 14.230 66.800 15.230 67.250 ;
        RECT 10.880 66.650 18.580 66.800 ;
        RECT 14.230 66.200 15.230 66.650 ;
        RECT 10.880 66.050 18.580 66.200 ;
        RECT 14.230 65.600 15.230 66.050 ;
        RECT 10.880 65.450 18.580 65.600 ;
        RECT 14.230 65.000 15.230 65.450 ;
        RECT 10.880 64.850 18.580 65.000 ;
        RECT 14.230 64.400 15.230 64.850 ;
        RECT 10.880 64.250 18.580 64.400 ;
        RECT 14.230 63.800 15.230 64.250 ;
        RECT 10.880 63.650 18.580 63.800 ;
        RECT 14.230 63.200 15.230 63.650 ;
        RECT 10.880 63.050 18.580 63.200 ;
        RECT 14.230 62.600 15.230 63.050 ;
        RECT 10.880 62.450 18.580 62.600 ;
        RECT 14.230 62.000 15.230 62.450 ;
        RECT 19.480 62.150 19.630 69.700 ;
        RECT 20.080 62.150 20.230 69.700 ;
        RECT 20.680 62.150 20.830 69.700 ;
        RECT 21.280 62.150 21.430 69.700 ;
        RECT 21.880 62.150 22.030 69.700 ;
        RECT 22.480 62.150 22.630 69.700 ;
        RECT 22.780 69.550 23.930 69.700 ;
        RECT 24.580 69.550 24.880 70.450 ;
        RECT 25.530 70.300 26.680 70.450 ;
        RECT 26.830 70.300 26.980 77.850 ;
        RECT 27.430 70.300 27.580 77.850 ;
        RECT 28.030 70.300 28.180 77.850 ;
        RECT 28.630 70.300 28.780 77.850 ;
        RECT 29.230 70.300 29.380 77.850 ;
        RECT 29.830 70.300 29.980 77.850 ;
        RECT 34.230 77.550 35.230 78.000 ;
        RECT 30.880 77.400 38.580 77.550 ;
        RECT 34.230 76.950 35.230 77.400 ;
        RECT 30.880 76.800 38.580 76.950 ;
        RECT 34.230 76.350 35.230 76.800 ;
        RECT 30.880 76.200 38.580 76.350 ;
        RECT 34.230 75.750 35.230 76.200 ;
        RECT 30.880 75.600 38.580 75.750 ;
        RECT 34.230 75.150 35.230 75.600 ;
        RECT 30.880 75.000 38.580 75.150 ;
        RECT 34.230 74.550 35.230 75.000 ;
        RECT 30.880 74.400 38.580 74.550 ;
        RECT 34.230 73.950 35.230 74.400 ;
        RECT 30.880 73.800 38.580 73.950 ;
        RECT 34.230 73.350 35.230 73.800 ;
        RECT 30.880 73.200 38.580 73.350 ;
        RECT 34.230 72.750 35.230 73.200 ;
        RECT 30.880 72.600 38.580 72.750 ;
        RECT 34.230 72.150 35.230 72.600 ;
        RECT 30.880 72.000 38.580 72.150 ;
        RECT 34.230 71.550 35.230 72.000 ;
        RECT 30.880 71.400 38.580 71.550 ;
        RECT 34.230 70.950 35.230 71.400 ;
        RECT 30.880 70.800 38.580 70.950 ;
        RECT 34.230 70.300 35.230 70.800 ;
        RECT 39.480 70.300 39.630 77.850 ;
        RECT 40.080 70.300 40.230 77.850 ;
        RECT 40.680 70.300 40.830 77.850 ;
        RECT 41.280 70.300 41.430 77.850 ;
        RECT 41.880 70.300 42.030 77.850 ;
        RECT 42.480 70.300 42.630 77.850 ;
        RECT 42.780 73.200 43.530 75.000 ;
        RECT 45.930 73.200 46.680 75.000 ;
        RECT 42.780 70.450 46.680 73.200 ;
        RECT 42.780 70.300 43.930 70.450 ;
        RECT 25.530 69.700 43.930 70.300 ;
        RECT 25.530 69.550 26.680 69.700 ;
        RECT 22.780 66.800 26.680 69.550 ;
        RECT 22.780 65.050 23.530 66.800 ;
        RECT 25.930 65.050 26.680 66.800 ;
        RECT 26.830 62.150 26.980 69.700 ;
        RECT 27.430 62.150 27.580 69.700 ;
        RECT 28.030 62.150 28.180 69.700 ;
        RECT 28.630 62.150 28.780 69.700 ;
        RECT 29.230 62.150 29.380 69.700 ;
        RECT 29.830 62.150 29.980 69.700 ;
        RECT 34.230 69.200 35.230 69.700 ;
        RECT 30.880 69.050 38.580 69.200 ;
        RECT 34.230 68.600 35.230 69.050 ;
        RECT 30.880 68.450 38.580 68.600 ;
        RECT 34.230 68.000 35.230 68.450 ;
        RECT 30.880 67.850 38.580 68.000 ;
        RECT 34.230 67.400 35.230 67.850 ;
        RECT 30.880 67.250 38.580 67.400 ;
        RECT 34.230 66.800 35.230 67.250 ;
        RECT 30.880 66.650 38.580 66.800 ;
        RECT 34.230 66.200 35.230 66.650 ;
        RECT 30.880 66.050 38.580 66.200 ;
        RECT 34.230 65.600 35.230 66.050 ;
        RECT 30.880 65.450 38.580 65.600 ;
        RECT 34.230 65.000 35.230 65.450 ;
        RECT 30.880 64.850 38.580 65.000 ;
        RECT 34.230 64.400 35.230 64.850 ;
        RECT 30.880 64.250 38.580 64.400 ;
        RECT 34.230 63.800 35.230 64.250 ;
        RECT 30.880 63.650 38.580 63.800 ;
        RECT 34.230 63.200 35.230 63.650 ;
        RECT 30.880 63.050 38.580 63.200 ;
        RECT 34.230 62.600 35.230 63.050 ;
        RECT 30.880 62.450 38.580 62.600 ;
        RECT 34.230 62.000 35.230 62.450 ;
        RECT 39.480 62.150 39.630 69.700 ;
        RECT 40.080 62.150 40.230 69.700 ;
        RECT 40.680 62.150 40.830 69.700 ;
        RECT 41.280 62.150 41.430 69.700 ;
        RECT 41.880 62.150 42.030 69.700 ;
        RECT 42.480 62.150 42.630 69.700 ;
        RECT 42.780 69.550 43.930 69.700 ;
        RECT 44.580 69.550 44.880 70.450 ;
        RECT 45.530 70.300 46.680 70.450 ;
        RECT 46.830 70.300 46.980 77.850 ;
        RECT 47.430 70.300 47.580 77.850 ;
        RECT 48.030 70.300 48.180 77.850 ;
        RECT 48.630 70.300 48.780 77.850 ;
        RECT 49.230 70.300 49.380 77.850 ;
        RECT 49.830 70.300 49.980 77.850 ;
        RECT 54.230 77.550 55.230 78.000 ;
        RECT 50.880 77.400 58.580 77.550 ;
        RECT 54.230 76.950 55.230 77.400 ;
        RECT 50.880 76.800 58.580 76.950 ;
        RECT 54.230 76.350 55.230 76.800 ;
        RECT 50.880 76.200 58.580 76.350 ;
        RECT 54.230 75.750 55.230 76.200 ;
        RECT 50.880 75.600 58.580 75.750 ;
        RECT 54.230 75.150 55.230 75.600 ;
        RECT 50.880 75.000 58.580 75.150 ;
        RECT 54.230 74.550 55.230 75.000 ;
        RECT 50.880 74.400 58.580 74.550 ;
        RECT 54.230 73.950 55.230 74.400 ;
        RECT 50.880 73.800 58.580 73.950 ;
        RECT 54.230 73.350 55.230 73.800 ;
        RECT 50.880 73.200 58.580 73.350 ;
        RECT 54.230 72.750 55.230 73.200 ;
        RECT 50.880 72.600 58.580 72.750 ;
        RECT 54.230 72.150 55.230 72.600 ;
        RECT 50.880 72.000 58.580 72.150 ;
        RECT 54.230 71.550 55.230 72.000 ;
        RECT 50.880 71.400 58.580 71.550 ;
        RECT 54.230 70.950 55.230 71.400 ;
        RECT 50.880 70.800 58.580 70.950 ;
        RECT 54.230 70.300 55.230 70.800 ;
        RECT 59.480 70.300 59.630 77.850 ;
        RECT 60.080 70.300 60.230 77.850 ;
        RECT 60.680 70.300 60.830 77.850 ;
        RECT 61.280 70.300 61.430 77.850 ;
        RECT 61.880 70.300 62.030 77.850 ;
        RECT 62.480 70.300 62.630 77.850 ;
        RECT 62.780 73.200 63.530 75.000 ;
        RECT 65.930 73.200 66.680 75.000 ;
        RECT 62.780 70.450 66.680 73.200 ;
        RECT 62.780 70.300 63.930 70.450 ;
        RECT 45.530 69.700 63.930 70.300 ;
        RECT 45.530 69.550 46.680 69.700 ;
        RECT 42.780 66.800 46.680 69.550 ;
        RECT 42.780 65.050 43.530 66.800 ;
        RECT 45.930 65.050 46.680 66.800 ;
        RECT 46.830 62.150 46.980 69.700 ;
        RECT 47.430 62.150 47.580 69.700 ;
        RECT 48.030 62.150 48.180 69.700 ;
        RECT 48.630 62.150 48.780 69.700 ;
        RECT 49.230 62.150 49.380 69.700 ;
        RECT 49.830 62.150 49.980 69.700 ;
        RECT 54.230 69.200 55.230 69.700 ;
        RECT 50.880 69.050 58.580 69.200 ;
        RECT 54.230 68.600 55.230 69.050 ;
        RECT 50.880 68.450 58.580 68.600 ;
        RECT 54.230 68.000 55.230 68.450 ;
        RECT 50.880 67.850 58.580 68.000 ;
        RECT 54.230 67.400 55.230 67.850 ;
        RECT 50.880 67.250 58.580 67.400 ;
        RECT 54.230 66.800 55.230 67.250 ;
        RECT 50.880 66.650 58.580 66.800 ;
        RECT 54.230 66.200 55.230 66.650 ;
        RECT 50.880 66.050 58.580 66.200 ;
        RECT 54.230 65.600 55.230 66.050 ;
        RECT 50.880 65.450 58.580 65.600 ;
        RECT 54.230 65.000 55.230 65.450 ;
        RECT 50.880 64.850 58.580 65.000 ;
        RECT 54.230 64.400 55.230 64.850 ;
        RECT 50.880 64.250 58.580 64.400 ;
        RECT 54.230 63.800 55.230 64.250 ;
        RECT 50.880 63.650 58.580 63.800 ;
        RECT 54.230 63.200 55.230 63.650 ;
        RECT 50.880 63.050 58.580 63.200 ;
        RECT 54.230 62.600 55.230 63.050 ;
        RECT 50.880 62.450 58.580 62.600 ;
        RECT 54.230 62.000 55.230 62.450 ;
        RECT 59.480 62.150 59.630 69.700 ;
        RECT 60.080 62.150 60.230 69.700 ;
        RECT 60.680 62.150 60.830 69.700 ;
        RECT 61.280 62.150 61.430 69.700 ;
        RECT 61.880 62.150 62.030 69.700 ;
        RECT 62.480 62.150 62.630 69.700 ;
        RECT 62.780 69.550 63.930 69.700 ;
        RECT 64.580 69.550 64.880 70.450 ;
        RECT 65.530 70.300 66.680 70.450 ;
        RECT 66.830 70.300 66.980 77.850 ;
        RECT 67.430 70.300 67.580 77.850 ;
        RECT 68.030 70.300 68.180 77.850 ;
        RECT 68.630 70.300 68.780 77.850 ;
        RECT 69.230 70.300 69.380 77.850 ;
        RECT 69.830 70.300 69.980 77.850 ;
        RECT 74.230 77.550 75.230 78.000 ;
        RECT 70.880 77.400 78.580 77.550 ;
        RECT 74.230 76.950 75.230 77.400 ;
        RECT 70.880 76.800 78.580 76.950 ;
        RECT 74.230 76.350 75.230 76.800 ;
        RECT 70.880 76.200 78.580 76.350 ;
        RECT 74.230 75.750 75.230 76.200 ;
        RECT 70.880 75.600 78.580 75.750 ;
        RECT 74.230 75.150 75.230 75.600 ;
        RECT 70.880 75.000 78.580 75.150 ;
        RECT 74.230 74.550 75.230 75.000 ;
        RECT 70.880 74.400 78.580 74.550 ;
        RECT 74.230 73.950 75.230 74.400 ;
        RECT 70.880 73.800 78.580 73.950 ;
        RECT 74.230 73.350 75.230 73.800 ;
        RECT 70.880 73.200 78.580 73.350 ;
        RECT 74.230 72.750 75.230 73.200 ;
        RECT 70.880 72.600 78.580 72.750 ;
        RECT 74.230 72.150 75.230 72.600 ;
        RECT 70.880 72.000 78.580 72.150 ;
        RECT 74.230 71.550 75.230 72.000 ;
        RECT 70.880 71.400 78.580 71.550 ;
        RECT 74.230 70.950 75.230 71.400 ;
        RECT 70.880 70.800 78.580 70.950 ;
        RECT 74.230 70.300 75.230 70.800 ;
        RECT 79.480 70.300 79.630 77.850 ;
        RECT 80.080 70.300 80.230 77.850 ;
        RECT 80.680 70.300 80.830 77.850 ;
        RECT 81.280 70.300 81.430 77.850 ;
        RECT 81.880 70.300 82.030 77.850 ;
        RECT 82.480 70.300 82.630 77.850 ;
        RECT 82.780 73.200 83.530 75.000 ;
        RECT 85.930 73.200 86.680 75.000 ;
        RECT 82.780 70.450 86.680 73.200 ;
        RECT 82.780 70.300 83.930 70.450 ;
        RECT 65.530 69.700 83.930 70.300 ;
        RECT 65.530 69.550 66.680 69.700 ;
        RECT 62.780 66.800 66.680 69.550 ;
        RECT 62.780 65.050 63.530 66.800 ;
        RECT 65.930 65.050 66.680 66.800 ;
        RECT 66.830 62.150 66.980 69.700 ;
        RECT 67.430 62.150 67.580 69.700 ;
        RECT 68.030 62.150 68.180 69.700 ;
        RECT 68.630 62.150 68.780 69.700 ;
        RECT 69.230 62.150 69.380 69.700 ;
        RECT 69.830 62.150 69.980 69.700 ;
        RECT 74.230 69.200 75.230 69.700 ;
        RECT 70.880 69.050 78.580 69.200 ;
        RECT 74.230 68.600 75.230 69.050 ;
        RECT 70.880 68.450 78.580 68.600 ;
        RECT 74.230 68.000 75.230 68.450 ;
        RECT 70.880 67.850 78.580 68.000 ;
        RECT 74.230 67.400 75.230 67.850 ;
        RECT 70.880 67.250 78.580 67.400 ;
        RECT 74.230 66.800 75.230 67.250 ;
        RECT 70.880 66.650 78.580 66.800 ;
        RECT 74.230 66.200 75.230 66.650 ;
        RECT 70.880 66.050 78.580 66.200 ;
        RECT 74.230 65.600 75.230 66.050 ;
        RECT 70.880 65.450 78.580 65.600 ;
        RECT 74.230 65.000 75.230 65.450 ;
        RECT 70.880 64.850 78.580 65.000 ;
        RECT 74.230 64.400 75.230 64.850 ;
        RECT 70.880 64.250 78.580 64.400 ;
        RECT 74.230 63.800 75.230 64.250 ;
        RECT 70.880 63.650 78.580 63.800 ;
        RECT 74.230 63.200 75.230 63.650 ;
        RECT 70.880 63.050 78.580 63.200 ;
        RECT 74.230 62.600 75.230 63.050 ;
        RECT 70.880 62.450 78.580 62.600 ;
        RECT 74.230 62.000 75.230 62.450 ;
        RECT 79.480 62.150 79.630 69.700 ;
        RECT 80.080 62.150 80.230 69.700 ;
        RECT 80.680 62.150 80.830 69.700 ;
        RECT 81.280 62.150 81.430 69.700 ;
        RECT 81.880 62.150 82.030 69.700 ;
        RECT 82.480 62.150 82.630 69.700 ;
        RECT 82.780 69.550 83.930 69.700 ;
        RECT 84.580 69.550 84.880 70.450 ;
        RECT 85.530 70.300 86.680 70.450 ;
        RECT 86.830 70.300 86.980 77.850 ;
        RECT 87.430 70.300 87.580 77.850 ;
        RECT 88.030 70.300 88.180 77.850 ;
        RECT 88.630 70.300 88.780 77.850 ;
        RECT 89.230 70.300 89.380 77.850 ;
        RECT 89.830 70.300 89.980 77.850 ;
        RECT 94.230 77.550 95.230 78.000 ;
        RECT 90.880 77.400 98.580 77.550 ;
        RECT 94.230 76.950 95.230 77.400 ;
        RECT 90.880 76.800 98.580 76.950 ;
        RECT 94.230 76.350 95.230 76.800 ;
        RECT 90.880 76.200 98.580 76.350 ;
        RECT 94.230 75.750 95.230 76.200 ;
        RECT 90.880 75.600 98.580 75.750 ;
        RECT 94.230 75.150 95.230 75.600 ;
        RECT 90.880 75.000 98.580 75.150 ;
        RECT 94.230 74.550 95.230 75.000 ;
        RECT 90.880 74.400 98.580 74.550 ;
        RECT 94.230 73.950 95.230 74.400 ;
        RECT 90.880 73.800 98.580 73.950 ;
        RECT 94.230 73.350 95.230 73.800 ;
        RECT 90.880 73.200 98.580 73.350 ;
        RECT 94.230 72.750 95.230 73.200 ;
        RECT 90.880 72.600 98.580 72.750 ;
        RECT 94.230 72.150 95.230 72.600 ;
        RECT 90.880 72.000 98.580 72.150 ;
        RECT 94.230 71.550 95.230 72.000 ;
        RECT 90.880 71.400 98.580 71.550 ;
        RECT 94.230 70.950 95.230 71.400 ;
        RECT 90.880 70.800 98.580 70.950 ;
        RECT 94.230 70.300 95.230 70.800 ;
        RECT 99.480 70.300 99.630 77.850 ;
        RECT 100.080 70.300 100.230 77.850 ;
        RECT 100.680 70.300 100.830 77.850 ;
        RECT 101.280 70.300 101.430 77.850 ;
        RECT 101.880 70.300 102.030 77.850 ;
        RECT 102.480 70.300 102.630 77.850 ;
        RECT 102.780 73.200 103.530 75.000 ;
        RECT 102.780 71.405 104.730 73.200 ;
        RECT 102.780 70.450 111.850 71.405 ;
        RECT 102.780 70.300 103.930 70.450 ;
        RECT 85.530 69.700 103.930 70.300 ;
        RECT 85.530 69.550 86.680 69.700 ;
        RECT 82.780 66.800 86.680 69.550 ;
        RECT 82.780 65.050 83.530 66.800 ;
        RECT 85.930 65.050 86.680 66.800 ;
        RECT 86.830 62.150 86.980 69.700 ;
        RECT 87.430 62.150 87.580 69.700 ;
        RECT 88.030 62.150 88.180 69.700 ;
        RECT 88.630 62.150 88.780 69.700 ;
        RECT 89.230 62.150 89.380 69.700 ;
        RECT 89.830 62.150 89.980 69.700 ;
        RECT 94.230 69.200 95.230 69.700 ;
        RECT 90.880 69.050 98.580 69.200 ;
        RECT 94.230 68.600 95.230 69.050 ;
        RECT 90.880 68.450 98.580 68.600 ;
        RECT 94.230 68.000 95.230 68.450 ;
        RECT 90.880 67.850 98.580 68.000 ;
        RECT 94.230 67.400 95.230 67.850 ;
        RECT 90.880 67.250 98.580 67.400 ;
        RECT 94.230 66.800 95.230 67.250 ;
        RECT 90.880 66.650 98.580 66.800 ;
        RECT 94.230 66.200 95.230 66.650 ;
        RECT 90.880 66.050 98.580 66.200 ;
        RECT 94.230 65.600 95.230 66.050 ;
        RECT 90.880 65.450 98.580 65.600 ;
        RECT 94.230 65.000 95.230 65.450 ;
        RECT 90.880 64.850 98.580 65.000 ;
        RECT 94.230 64.400 95.230 64.850 ;
        RECT 90.880 64.250 98.580 64.400 ;
        RECT 94.230 63.800 95.230 64.250 ;
        RECT 90.880 63.650 98.580 63.800 ;
        RECT 94.230 63.200 95.230 63.650 ;
        RECT 90.880 63.050 98.580 63.200 ;
        RECT 94.230 62.600 95.230 63.050 ;
        RECT 90.880 62.450 98.580 62.600 ;
        RECT 94.230 62.000 95.230 62.450 ;
        RECT 99.480 62.150 99.630 69.700 ;
        RECT 100.080 62.150 100.230 69.700 ;
        RECT 100.680 62.150 100.830 69.700 ;
        RECT 101.280 62.150 101.430 69.700 ;
        RECT 101.880 62.150 102.030 69.700 ;
        RECT 102.480 62.150 102.630 69.700 ;
        RECT 102.780 69.550 103.930 69.700 ;
        RECT 104.580 70.130 111.850 70.450 ;
        RECT 104.580 69.550 104.730 70.130 ;
        RECT 102.780 66.800 104.730 69.550 ;
        RECT 102.780 65.050 103.530 66.800 ;
        RECT 10.880 61.850 18.580 62.000 ;
        RECT 30.880 61.850 38.580 62.000 ;
        RECT 50.880 61.850 58.580 62.000 ;
        RECT 70.880 61.850 78.580 62.000 ;
        RECT 90.880 61.850 98.580 62.000 ;
        RECT 14.230 61.200 15.230 61.850 ;
        RECT 34.230 61.200 35.230 61.850 ;
        RECT 54.230 61.200 55.230 61.850 ;
        RECT 74.230 61.200 75.230 61.850 ;
        RECT 94.230 61.200 95.230 61.850 ;
        RECT 11.530 58.800 17.930 61.200 ;
        RECT 31.530 58.800 37.930 61.200 ;
        RECT 51.530 58.800 57.930 61.200 ;
        RECT 71.530 58.800 77.930 61.200 ;
        RECT 91.530 58.800 97.930 61.200 ;
        RECT 14.230 58.150 15.230 58.800 ;
        RECT 34.230 58.150 35.230 58.800 ;
        RECT 54.230 58.150 55.230 58.800 ;
        RECT 74.230 58.150 75.230 58.800 ;
        RECT 94.230 58.150 95.230 58.800 ;
        RECT 10.880 58.000 18.580 58.150 ;
        RECT 30.880 58.000 38.580 58.150 ;
        RECT 50.880 58.000 58.580 58.150 ;
        RECT 70.880 58.000 78.580 58.150 ;
        RECT 90.880 58.000 98.580 58.150 ;
        RECT 5.930 53.200 6.680 55.000 ;
        RECT 4.730 50.450 6.680 53.200 ;
        RECT 4.730 49.550 4.880 50.450 ;
        RECT 5.530 50.300 6.680 50.450 ;
        RECT 6.830 50.300 6.980 57.850 ;
        RECT 7.430 50.300 7.580 57.850 ;
        RECT 8.030 50.300 8.180 57.850 ;
        RECT 8.630 50.300 8.780 57.850 ;
        RECT 9.230 50.300 9.380 57.850 ;
        RECT 9.830 50.300 9.980 57.850 ;
        RECT 14.230 57.550 15.230 58.000 ;
        RECT 10.880 57.400 18.580 57.550 ;
        RECT 14.230 56.950 15.230 57.400 ;
        RECT 10.880 56.800 18.580 56.950 ;
        RECT 14.230 56.350 15.230 56.800 ;
        RECT 10.880 56.200 18.580 56.350 ;
        RECT 14.230 55.750 15.230 56.200 ;
        RECT 10.880 55.600 18.580 55.750 ;
        RECT 14.230 55.150 15.230 55.600 ;
        RECT 10.880 55.000 18.580 55.150 ;
        RECT 14.230 54.550 15.230 55.000 ;
        RECT 10.880 54.400 18.580 54.550 ;
        RECT 14.230 53.950 15.230 54.400 ;
        RECT 10.880 53.800 18.580 53.950 ;
        RECT 14.230 53.350 15.230 53.800 ;
        RECT 10.880 53.200 18.580 53.350 ;
        RECT 14.230 52.750 15.230 53.200 ;
        RECT 10.880 52.600 18.580 52.750 ;
        RECT 14.230 52.150 15.230 52.600 ;
        RECT 10.880 52.000 18.580 52.150 ;
        RECT 14.230 51.550 15.230 52.000 ;
        RECT 10.880 51.400 18.580 51.550 ;
        RECT 14.230 50.950 15.230 51.400 ;
        RECT 10.880 50.800 18.580 50.950 ;
        RECT 14.230 50.300 15.230 50.800 ;
        RECT 19.480 50.300 19.630 57.850 ;
        RECT 20.080 50.300 20.230 57.850 ;
        RECT 20.680 50.300 20.830 57.850 ;
        RECT 21.280 50.300 21.430 57.850 ;
        RECT 21.880 50.300 22.030 57.850 ;
        RECT 22.480 50.300 22.630 57.850 ;
        RECT 22.780 53.200 23.530 55.000 ;
        RECT 25.930 53.200 26.680 55.000 ;
        RECT 22.780 50.450 26.680 53.200 ;
        RECT 22.780 50.300 23.930 50.450 ;
        RECT 5.530 49.700 23.930 50.300 ;
        RECT 5.530 49.550 6.680 49.700 ;
        RECT 4.730 46.800 6.680 49.550 ;
        RECT 5.930 45.050 6.680 46.800 ;
        RECT 6.830 42.150 6.980 49.700 ;
        RECT 7.430 42.150 7.580 49.700 ;
        RECT 8.030 42.150 8.180 49.700 ;
        RECT 8.630 42.150 8.780 49.700 ;
        RECT 9.230 42.150 9.380 49.700 ;
        RECT 9.830 42.150 9.980 49.700 ;
        RECT 14.230 49.200 15.230 49.700 ;
        RECT 10.880 49.050 18.580 49.200 ;
        RECT 14.230 48.600 15.230 49.050 ;
        RECT 10.880 48.450 18.580 48.600 ;
        RECT 14.230 48.000 15.230 48.450 ;
        RECT 10.880 47.850 18.580 48.000 ;
        RECT 14.230 47.400 15.230 47.850 ;
        RECT 10.880 47.250 18.580 47.400 ;
        RECT 14.230 46.800 15.230 47.250 ;
        RECT 10.880 46.650 18.580 46.800 ;
        RECT 14.230 46.200 15.230 46.650 ;
        RECT 10.880 46.050 18.580 46.200 ;
        RECT 14.230 45.600 15.230 46.050 ;
        RECT 10.880 45.450 18.580 45.600 ;
        RECT 14.230 45.000 15.230 45.450 ;
        RECT 10.880 44.850 18.580 45.000 ;
        RECT 14.230 44.400 15.230 44.850 ;
        RECT 10.880 44.250 18.580 44.400 ;
        RECT 14.230 43.800 15.230 44.250 ;
        RECT 10.880 43.650 18.580 43.800 ;
        RECT 14.230 43.200 15.230 43.650 ;
        RECT 10.880 43.050 18.580 43.200 ;
        RECT 14.230 42.600 15.230 43.050 ;
        RECT 10.880 42.450 18.580 42.600 ;
        RECT 14.230 42.000 15.230 42.450 ;
        RECT 19.480 42.150 19.630 49.700 ;
        RECT 20.080 42.150 20.230 49.700 ;
        RECT 20.680 42.150 20.830 49.700 ;
        RECT 21.280 42.150 21.430 49.700 ;
        RECT 21.880 42.150 22.030 49.700 ;
        RECT 22.480 42.150 22.630 49.700 ;
        RECT 22.780 49.550 23.930 49.700 ;
        RECT 24.580 49.550 24.880 50.450 ;
        RECT 25.530 50.300 26.680 50.450 ;
        RECT 26.830 50.300 26.980 57.850 ;
        RECT 27.430 50.300 27.580 57.850 ;
        RECT 28.030 50.300 28.180 57.850 ;
        RECT 28.630 50.300 28.780 57.850 ;
        RECT 29.230 50.300 29.380 57.850 ;
        RECT 29.830 50.300 29.980 57.850 ;
        RECT 34.230 57.550 35.230 58.000 ;
        RECT 30.880 57.400 38.580 57.550 ;
        RECT 34.230 56.950 35.230 57.400 ;
        RECT 30.880 56.800 38.580 56.950 ;
        RECT 34.230 56.350 35.230 56.800 ;
        RECT 30.880 56.200 38.580 56.350 ;
        RECT 34.230 55.750 35.230 56.200 ;
        RECT 30.880 55.600 38.580 55.750 ;
        RECT 34.230 55.150 35.230 55.600 ;
        RECT 30.880 55.000 38.580 55.150 ;
        RECT 34.230 54.550 35.230 55.000 ;
        RECT 30.880 54.400 38.580 54.550 ;
        RECT 34.230 53.950 35.230 54.400 ;
        RECT 30.880 53.800 38.580 53.950 ;
        RECT 34.230 53.350 35.230 53.800 ;
        RECT 30.880 53.200 38.580 53.350 ;
        RECT 34.230 52.750 35.230 53.200 ;
        RECT 30.880 52.600 38.580 52.750 ;
        RECT 34.230 52.150 35.230 52.600 ;
        RECT 30.880 52.000 38.580 52.150 ;
        RECT 34.230 51.550 35.230 52.000 ;
        RECT 30.880 51.400 38.580 51.550 ;
        RECT 34.230 50.950 35.230 51.400 ;
        RECT 30.880 50.800 38.580 50.950 ;
        RECT 34.230 50.300 35.230 50.800 ;
        RECT 39.480 50.300 39.630 57.850 ;
        RECT 40.080 50.300 40.230 57.850 ;
        RECT 40.680 50.300 40.830 57.850 ;
        RECT 41.280 50.300 41.430 57.850 ;
        RECT 41.880 50.300 42.030 57.850 ;
        RECT 42.480 50.300 42.630 57.850 ;
        RECT 42.780 53.200 43.530 55.000 ;
        RECT 45.930 53.200 46.680 55.000 ;
        RECT 42.780 50.450 46.680 53.200 ;
        RECT 42.780 50.300 43.930 50.450 ;
        RECT 25.530 49.700 43.930 50.300 ;
        RECT 25.530 49.550 26.680 49.700 ;
        RECT 22.780 46.800 26.680 49.550 ;
        RECT 22.780 45.050 23.530 46.800 ;
        RECT 25.930 45.050 26.680 46.800 ;
        RECT 26.830 42.150 26.980 49.700 ;
        RECT 27.430 42.150 27.580 49.700 ;
        RECT 28.030 42.150 28.180 49.700 ;
        RECT 28.630 42.150 28.780 49.700 ;
        RECT 29.230 42.150 29.380 49.700 ;
        RECT 29.830 42.150 29.980 49.700 ;
        RECT 34.230 49.200 35.230 49.700 ;
        RECT 30.880 49.050 38.580 49.200 ;
        RECT 34.230 48.600 35.230 49.050 ;
        RECT 30.880 48.450 38.580 48.600 ;
        RECT 34.230 48.000 35.230 48.450 ;
        RECT 30.880 47.850 38.580 48.000 ;
        RECT 34.230 47.400 35.230 47.850 ;
        RECT 30.880 47.250 38.580 47.400 ;
        RECT 34.230 46.800 35.230 47.250 ;
        RECT 30.880 46.650 38.580 46.800 ;
        RECT 34.230 46.200 35.230 46.650 ;
        RECT 30.880 46.050 38.580 46.200 ;
        RECT 34.230 45.600 35.230 46.050 ;
        RECT 30.880 45.450 38.580 45.600 ;
        RECT 34.230 45.000 35.230 45.450 ;
        RECT 30.880 44.850 38.580 45.000 ;
        RECT 34.230 44.400 35.230 44.850 ;
        RECT 30.880 44.250 38.580 44.400 ;
        RECT 34.230 43.800 35.230 44.250 ;
        RECT 30.880 43.650 38.580 43.800 ;
        RECT 34.230 43.200 35.230 43.650 ;
        RECT 30.880 43.050 38.580 43.200 ;
        RECT 34.230 42.600 35.230 43.050 ;
        RECT 30.880 42.450 38.580 42.600 ;
        RECT 34.230 42.000 35.230 42.450 ;
        RECT 39.480 42.150 39.630 49.700 ;
        RECT 40.080 42.150 40.230 49.700 ;
        RECT 40.680 42.150 40.830 49.700 ;
        RECT 41.280 42.150 41.430 49.700 ;
        RECT 41.880 42.150 42.030 49.700 ;
        RECT 42.480 42.150 42.630 49.700 ;
        RECT 42.780 49.550 43.930 49.700 ;
        RECT 44.580 49.550 44.880 50.450 ;
        RECT 45.530 50.300 46.680 50.450 ;
        RECT 46.830 50.300 46.980 57.850 ;
        RECT 47.430 50.300 47.580 57.850 ;
        RECT 48.030 50.300 48.180 57.850 ;
        RECT 48.630 50.300 48.780 57.850 ;
        RECT 49.230 50.300 49.380 57.850 ;
        RECT 49.830 50.300 49.980 57.850 ;
        RECT 54.230 57.550 55.230 58.000 ;
        RECT 50.880 57.400 58.580 57.550 ;
        RECT 54.230 56.950 55.230 57.400 ;
        RECT 50.880 56.800 58.580 56.950 ;
        RECT 54.230 56.350 55.230 56.800 ;
        RECT 50.880 56.200 58.580 56.350 ;
        RECT 54.230 55.750 55.230 56.200 ;
        RECT 50.880 55.600 58.580 55.750 ;
        RECT 54.230 55.150 55.230 55.600 ;
        RECT 50.880 55.000 58.580 55.150 ;
        RECT 54.230 54.550 55.230 55.000 ;
        RECT 50.880 54.400 58.580 54.550 ;
        RECT 54.230 53.950 55.230 54.400 ;
        RECT 50.880 53.800 58.580 53.950 ;
        RECT 54.230 53.350 55.230 53.800 ;
        RECT 50.880 53.200 58.580 53.350 ;
        RECT 54.230 52.750 55.230 53.200 ;
        RECT 50.880 52.600 58.580 52.750 ;
        RECT 54.230 52.150 55.230 52.600 ;
        RECT 50.880 52.000 58.580 52.150 ;
        RECT 54.230 51.550 55.230 52.000 ;
        RECT 50.880 51.400 58.580 51.550 ;
        RECT 54.230 50.950 55.230 51.400 ;
        RECT 50.880 50.800 58.580 50.950 ;
        RECT 54.230 50.300 55.230 50.800 ;
        RECT 59.480 50.300 59.630 57.850 ;
        RECT 60.080 50.300 60.230 57.850 ;
        RECT 60.680 50.300 60.830 57.850 ;
        RECT 61.280 50.300 61.430 57.850 ;
        RECT 61.880 50.300 62.030 57.850 ;
        RECT 62.480 50.300 62.630 57.850 ;
        RECT 62.780 53.200 63.530 55.000 ;
        RECT 65.930 53.200 66.680 55.000 ;
        RECT 62.780 50.450 66.680 53.200 ;
        RECT 62.780 50.300 63.930 50.450 ;
        RECT 45.530 49.700 63.930 50.300 ;
        RECT 45.530 49.550 46.680 49.700 ;
        RECT 42.780 46.800 46.680 49.550 ;
        RECT 42.780 45.050 43.530 46.800 ;
        RECT 45.930 45.050 46.680 46.800 ;
        RECT 46.830 42.150 46.980 49.700 ;
        RECT 47.430 42.150 47.580 49.700 ;
        RECT 48.030 42.150 48.180 49.700 ;
        RECT 48.630 42.150 48.780 49.700 ;
        RECT 49.230 42.150 49.380 49.700 ;
        RECT 49.830 42.150 49.980 49.700 ;
        RECT 54.230 49.200 55.230 49.700 ;
        RECT 50.880 49.050 58.580 49.200 ;
        RECT 54.230 48.600 55.230 49.050 ;
        RECT 50.880 48.450 58.580 48.600 ;
        RECT 54.230 48.000 55.230 48.450 ;
        RECT 50.880 47.850 58.580 48.000 ;
        RECT 54.230 47.400 55.230 47.850 ;
        RECT 50.880 47.250 58.580 47.400 ;
        RECT 54.230 46.800 55.230 47.250 ;
        RECT 50.880 46.650 58.580 46.800 ;
        RECT 54.230 46.200 55.230 46.650 ;
        RECT 50.880 46.050 58.580 46.200 ;
        RECT 54.230 45.600 55.230 46.050 ;
        RECT 50.880 45.450 58.580 45.600 ;
        RECT 54.230 45.000 55.230 45.450 ;
        RECT 50.880 44.850 58.580 45.000 ;
        RECT 54.230 44.400 55.230 44.850 ;
        RECT 50.880 44.250 58.580 44.400 ;
        RECT 54.230 43.800 55.230 44.250 ;
        RECT 50.880 43.650 58.580 43.800 ;
        RECT 54.230 43.200 55.230 43.650 ;
        RECT 50.880 43.050 58.580 43.200 ;
        RECT 54.230 42.600 55.230 43.050 ;
        RECT 50.880 42.450 58.580 42.600 ;
        RECT 54.230 42.000 55.230 42.450 ;
        RECT 59.480 42.150 59.630 49.700 ;
        RECT 60.080 42.150 60.230 49.700 ;
        RECT 60.680 42.150 60.830 49.700 ;
        RECT 61.280 42.150 61.430 49.700 ;
        RECT 61.880 42.150 62.030 49.700 ;
        RECT 62.480 42.150 62.630 49.700 ;
        RECT 62.780 49.550 63.930 49.700 ;
        RECT 64.580 49.550 64.880 50.450 ;
        RECT 65.530 50.300 66.680 50.450 ;
        RECT 66.830 50.300 66.980 57.850 ;
        RECT 67.430 50.300 67.580 57.850 ;
        RECT 68.030 50.300 68.180 57.850 ;
        RECT 68.630 50.300 68.780 57.850 ;
        RECT 69.230 50.300 69.380 57.850 ;
        RECT 69.830 50.300 69.980 57.850 ;
        RECT 74.230 57.550 75.230 58.000 ;
        RECT 70.880 57.400 78.580 57.550 ;
        RECT 74.230 56.950 75.230 57.400 ;
        RECT 70.880 56.800 78.580 56.950 ;
        RECT 74.230 56.350 75.230 56.800 ;
        RECT 70.880 56.200 78.580 56.350 ;
        RECT 74.230 55.750 75.230 56.200 ;
        RECT 70.880 55.600 78.580 55.750 ;
        RECT 74.230 55.150 75.230 55.600 ;
        RECT 70.880 55.000 78.580 55.150 ;
        RECT 74.230 54.550 75.230 55.000 ;
        RECT 70.880 54.400 78.580 54.550 ;
        RECT 74.230 53.950 75.230 54.400 ;
        RECT 70.880 53.800 78.580 53.950 ;
        RECT 74.230 53.350 75.230 53.800 ;
        RECT 70.880 53.200 78.580 53.350 ;
        RECT 74.230 52.750 75.230 53.200 ;
        RECT 70.880 52.600 78.580 52.750 ;
        RECT 74.230 52.150 75.230 52.600 ;
        RECT 70.880 52.000 78.580 52.150 ;
        RECT 74.230 51.550 75.230 52.000 ;
        RECT 70.880 51.400 78.580 51.550 ;
        RECT 74.230 50.950 75.230 51.400 ;
        RECT 70.880 50.800 78.580 50.950 ;
        RECT 74.230 50.300 75.230 50.800 ;
        RECT 79.480 50.300 79.630 57.850 ;
        RECT 80.080 50.300 80.230 57.850 ;
        RECT 80.680 50.300 80.830 57.850 ;
        RECT 81.280 50.300 81.430 57.850 ;
        RECT 81.880 50.300 82.030 57.850 ;
        RECT 82.480 50.300 82.630 57.850 ;
        RECT 82.780 53.200 83.530 55.000 ;
        RECT 85.930 53.200 86.680 55.000 ;
        RECT 82.780 50.450 86.680 53.200 ;
        RECT 82.780 50.300 83.930 50.450 ;
        RECT 65.530 49.700 83.930 50.300 ;
        RECT 65.530 49.550 66.680 49.700 ;
        RECT 62.780 46.800 66.680 49.550 ;
        RECT 62.780 45.050 63.530 46.800 ;
        RECT 65.930 45.050 66.680 46.800 ;
        RECT 66.830 42.150 66.980 49.700 ;
        RECT 67.430 42.150 67.580 49.700 ;
        RECT 68.030 42.150 68.180 49.700 ;
        RECT 68.630 42.150 68.780 49.700 ;
        RECT 69.230 42.150 69.380 49.700 ;
        RECT 69.830 42.150 69.980 49.700 ;
        RECT 74.230 49.200 75.230 49.700 ;
        RECT 70.880 49.050 78.580 49.200 ;
        RECT 74.230 48.600 75.230 49.050 ;
        RECT 70.880 48.450 78.580 48.600 ;
        RECT 74.230 48.000 75.230 48.450 ;
        RECT 70.880 47.850 78.580 48.000 ;
        RECT 74.230 47.400 75.230 47.850 ;
        RECT 70.880 47.250 78.580 47.400 ;
        RECT 74.230 46.800 75.230 47.250 ;
        RECT 70.880 46.650 78.580 46.800 ;
        RECT 74.230 46.200 75.230 46.650 ;
        RECT 70.880 46.050 78.580 46.200 ;
        RECT 74.230 45.600 75.230 46.050 ;
        RECT 70.880 45.450 78.580 45.600 ;
        RECT 74.230 45.000 75.230 45.450 ;
        RECT 70.880 44.850 78.580 45.000 ;
        RECT 74.230 44.400 75.230 44.850 ;
        RECT 70.880 44.250 78.580 44.400 ;
        RECT 74.230 43.800 75.230 44.250 ;
        RECT 70.880 43.650 78.580 43.800 ;
        RECT 74.230 43.200 75.230 43.650 ;
        RECT 70.880 43.050 78.580 43.200 ;
        RECT 74.230 42.600 75.230 43.050 ;
        RECT 70.880 42.450 78.580 42.600 ;
        RECT 74.230 42.000 75.230 42.450 ;
        RECT 79.480 42.150 79.630 49.700 ;
        RECT 80.080 42.150 80.230 49.700 ;
        RECT 80.680 42.150 80.830 49.700 ;
        RECT 81.280 42.150 81.430 49.700 ;
        RECT 81.880 42.150 82.030 49.700 ;
        RECT 82.480 42.150 82.630 49.700 ;
        RECT 82.780 49.550 83.930 49.700 ;
        RECT 84.580 49.550 84.880 50.450 ;
        RECT 85.530 50.300 86.680 50.450 ;
        RECT 86.830 50.300 86.980 57.850 ;
        RECT 87.430 50.300 87.580 57.850 ;
        RECT 88.030 50.300 88.180 57.850 ;
        RECT 88.630 50.300 88.780 57.850 ;
        RECT 89.230 50.300 89.380 57.850 ;
        RECT 89.830 50.300 89.980 57.850 ;
        RECT 94.230 57.550 95.230 58.000 ;
        RECT 90.880 57.400 98.580 57.550 ;
        RECT 94.230 56.950 95.230 57.400 ;
        RECT 90.880 56.800 98.580 56.950 ;
        RECT 94.230 56.350 95.230 56.800 ;
        RECT 90.880 56.200 98.580 56.350 ;
        RECT 94.230 55.750 95.230 56.200 ;
        RECT 90.880 55.600 98.580 55.750 ;
        RECT 94.230 55.150 95.230 55.600 ;
        RECT 90.880 55.000 98.580 55.150 ;
        RECT 94.230 54.550 95.230 55.000 ;
        RECT 90.880 54.400 98.580 54.550 ;
        RECT 94.230 53.950 95.230 54.400 ;
        RECT 90.880 53.800 98.580 53.950 ;
        RECT 94.230 53.350 95.230 53.800 ;
        RECT 90.880 53.200 98.580 53.350 ;
        RECT 94.230 52.750 95.230 53.200 ;
        RECT 90.880 52.600 98.580 52.750 ;
        RECT 94.230 52.150 95.230 52.600 ;
        RECT 90.880 52.000 98.580 52.150 ;
        RECT 94.230 51.550 95.230 52.000 ;
        RECT 90.880 51.400 98.580 51.550 ;
        RECT 94.230 50.950 95.230 51.400 ;
        RECT 90.880 50.800 98.580 50.950 ;
        RECT 94.230 50.300 95.230 50.800 ;
        RECT 99.480 50.300 99.630 57.850 ;
        RECT 100.080 50.300 100.230 57.850 ;
        RECT 100.680 50.300 100.830 57.850 ;
        RECT 101.280 50.300 101.430 57.850 ;
        RECT 101.880 50.300 102.030 57.850 ;
        RECT 102.480 50.300 102.630 57.850 ;
        RECT 102.780 53.200 103.530 55.000 ;
        RECT 102.780 51.585 104.730 53.200 ;
        RECT 102.780 50.450 111.850 51.585 ;
        RECT 102.780 50.300 103.930 50.450 ;
        RECT 85.530 49.700 103.930 50.300 ;
        RECT 85.530 49.550 86.680 49.700 ;
        RECT 82.780 46.800 86.680 49.550 ;
        RECT 82.780 45.050 83.530 46.800 ;
        RECT 85.930 45.050 86.680 46.800 ;
        RECT 86.830 42.150 86.980 49.700 ;
        RECT 87.430 42.150 87.580 49.700 ;
        RECT 88.030 42.150 88.180 49.700 ;
        RECT 88.630 42.150 88.780 49.700 ;
        RECT 89.230 42.150 89.380 49.700 ;
        RECT 89.830 42.150 89.980 49.700 ;
        RECT 94.230 49.200 95.230 49.700 ;
        RECT 90.880 49.050 98.580 49.200 ;
        RECT 94.230 48.600 95.230 49.050 ;
        RECT 90.880 48.450 98.580 48.600 ;
        RECT 94.230 48.000 95.230 48.450 ;
        RECT 90.880 47.850 98.580 48.000 ;
        RECT 94.230 47.400 95.230 47.850 ;
        RECT 90.880 47.250 98.580 47.400 ;
        RECT 94.230 46.800 95.230 47.250 ;
        RECT 90.880 46.650 98.580 46.800 ;
        RECT 94.230 46.200 95.230 46.650 ;
        RECT 90.880 46.050 98.580 46.200 ;
        RECT 94.230 45.600 95.230 46.050 ;
        RECT 90.880 45.450 98.580 45.600 ;
        RECT 94.230 45.000 95.230 45.450 ;
        RECT 90.880 44.850 98.580 45.000 ;
        RECT 94.230 44.400 95.230 44.850 ;
        RECT 90.880 44.250 98.580 44.400 ;
        RECT 94.230 43.800 95.230 44.250 ;
        RECT 90.880 43.650 98.580 43.800 ;
        RECT 94.230 43.200 95.230 43.650 ;
        RECT 90.880 43.050 98.580 43.200 ;
        RECT 94.230 42.600 95.230 43.050 ;
        RECT 90.880 42.450 98.580 42.600 ;
        RECT 94.230 42.000 95.230 42.450 ;
        RECT 99.480 42.150 99.630 49.700 ;
        RECT 100.080 42.150 100.230 49.700 ;
        RECT 100.680 42.150 100.830 49.700 ;
        RECT 101.280 42.150 101.430 49.700 ;
        RECT 101.880 42.150 102.030 49.700 ;
        RECT 102.480 42.150 102.630 49.700 ;
        RECT 102.780 49.550 103.930 49.700 ;
        RECT 104.580 50.310 111.850 50.450 ;
        RECT 104.580 49.550 104.730 50.310 ;
        RECT 102.780 46.800 104.730 49.550 ;
        RECT 102.780 45.050 103.530 46.800 ;
        RECT 10.880 41.850 18.580 42.000 ;
        RECT 30.880 41.850 38.580 42.000 ;
        RECT 50.880 41.850 58.580 42.000 ;
        RECT 70.880 41.850 78.580 42.000 ;
        RECT 90.880 41.850 98.580 42.000 ;
        RECT 14.230 41.200 15.230 41.850 ;
        RECT 34.230 41.200 35.230 41.850 ;
        RECT 54.230 41.200 55.230 41.850 ;
        RECT 74.230 41.200 75.230 41.850 ;
        RECT 94.230 41.200 95.230 41.850 ;
        RECT 11.530 38.800 17.930 41.200 ;
        RECT 31.530 38.800 37.930 41.200 ;
        RECT 51.530 38.800 57.930 41.200 ;
        RECT 71.530 38.800 77.930 41.200 ;
        RECT 91.530 38.800 97.930 41.200 ;
        RECT 14.230 38.150 15.230 38.800 ;
        RECT 34.230 38.150 35.230 38.800 ;
        RECT 54.230 38.150 55.230 38.800 ;
        RECT 74.230 38.150 75.230 38.800 ;
        RECT 94.230 38.150 95.230 38.800 ;
        RECT 10.880 38.000 18.580 38.150 ;
        RECT 30.880 38.000 38.580 38.150 ;
        RECT 50.880 38.000 58.580 38.150 ;
        RECT 70.880 38.000 78.580 38.150 ;
        RECT 90.880 38.000 98.580 38.150 ;
        RECT 5.930 33.200 6.680 35.000 ;
        RECT 4.730 30.450 6.680 33.200 ;
        RECT 4.730 29.550 4.880 30.450 ;
        RECT 5.530 30.300 6.680 30.450 ;
        RECT 6.830 30.300 6.980 37.850 ;
        RECT 7.430 30.300 7.580 37.850 ;
        RECT 8.030 30.300 8.180 37.850 ;
        RECT 8.630 30.300 8.780 37.850 ;
        RECT 9.230 30.300 9.380 37.850 ;
        RECT 9.830 30.300 9.980 37.850 ;
        RECT 14.230 37.550 15.230 38.000 ;
        RECT 10.880 37.400 18.580 37.550 ;
        RECT 14.230 36.950 15.230 37.400 ;
        RECT 10.880 36.800 18.580 36.950 ;
        RECT 14.230 36.350 15.230 36.800 ;
        RECT 10.880 36.200 18.580 36.350 ;
        RECT 14.230 35.750 15.230 36.200 ;
        RECT 10.880 35.600 18.580 35.750 ;
        RECT 14.230 35.150 15.230 35.600 ;
        RECT 10.880 35.000 18.580 35.150 ;
        RECT 14.230 34.550 15.230 35.000 ;
        RECT 10.880 34.400 18.580 34.550 ;
        RECT 14.230 33.950 15.230 34.400 ;
        RECT 10.880 33.800 18.580 33.950 ;
        RECT 14.230 33.350 15.230 33.800 ;
        RECT 10.880 33.200 18.580 33.350 ;
        RECT 14.230 32.750 15.230 33.200 ;
        RECT 10.880 32.600 18.580 32.750 ;
        RECT 14.230 32.150 15.230 32.600 ;
        RECT 10.880 32.000 18.580 32.150 ;
        RECT 14.230 31.550 15.230 32.000 ;
        RECT 10.880 31.400 18.580 31.550 ;
        RECT 14.230 30.950 15.230 31.400 ;
        RECT 10.880 30.800 18.580 30.950 ;
        RECT 14.230 30.300 15.230 30.800 ;
        RECT 19.480 30.300 19.630 37.850 ;
        RECT 20.080 30.300 20.230 37.850 ;
        RECT 20.680 30.300 20.830 37.850 ;
        RECT 21.280 30.300 21.430 37.850 ;
        RECT 21.880 30.300 22.030 37.850 ;
        RECT 22.480 30.300 22.630 37.850 ;
        RECT 22.780 33.200 23.530 35.000 ;
        RECT 25.930 33.200 26.680 35.000 ;
        RECT 22.780 30.450 26.680 33.200 ;
        RECT 22.780 30.300 23.930 30.450 ;
        RECT 5.530 29.700 23.930 30.300 ;
        RECT 5.530 29.550 6.680 29.700 ;
        RECT 4.730 26.800 6.680 29.550 ;
        RECT 5.930 25.050 6.680 26.800 ;
        RECT 6.830 22.150 6.980 29.700 ;
        RECT 7.430 22.150 7.580 29.700 ;
        RECT 8.030 22.150 8.180 29.700 ;
        RECT 8.630 22.150 8.780 29.700 ;
        RECT 9.230 22.150 9.380 29.700 ;
        RECT 9.830 22.150 9.980 29.700 ;
        RECT 14.230 29.200 15.230 29.700 ;
        RECT 10.880 29.050 18.580 29.200 ;
        RECT 14.230 28.600 15.230 29.050 ;
        RECT 10.880 28.450 18.580 28.600 ;
        RECT 14.230 28.000 15.230 28.450 ;
        RECT 10.880 27.850 18.580 28.000 ;
        RECT 14.230 27.400 15.230 27.850 ;
        RECT 10.880 27.250 18.580 27.400 ;
        RECT 14.230 26.800 15.230 27.250 ;
        RECT 10.880 26.650 18.580 26.800 ;
        RECT 14.230 26.200 15.230 26.650 ;
        RECT 10.880 26.050 18.580 26.200 ;
        RECT 14.230 25.600 15.230 26.050 ;
        RECT 10.880 25.450 18.580 25.600 ;
        RECT 14.230 25.000 15.230 25.450 ;
        RECT 10.880 24.850 18.580 25.000 ;
        RECT 14.230 24.400 15.230 24.850 ;
        RECT 10.880 24.250 18.580 24.400 ;
        RECT 14.230 23.800 15.230 24.250 ;
        RECT 10.880 23.650 18.580 23.800 ;
        RECT 14.230 23.200 15.230 23.650 ;
        RECT 10.880 23.050 18.580 23.200 ;
        RECT 14.230 22.600 15.230 23.050 ;
        RECT 10.880 22.450 18.580 22.600 ;
        RECT 14.230 22.000 15.230 22.450 ;
        RECT 19.480 22.150 19.630 29.700 ;
        RECT 20.080 22.150 20.230 29.700 ;
        RECT 20.680 22.150 20.830 29.700 ;
        RECT 21.280 22.150 21.430 29.700 ;
        RECT 21.880 22.150 22.030 29.700 ;
        RECT 22.480 22.150 22.630 29.700 ;
        RECT 22.780 29.550 23.930 29.700 ;
        RECT 24.580 29.550 24.880 30.450 ;
        RECT 25.530 30.300 26.680 30.450 ;
        RECT 26.830 30.300 26.980 37.850 ;
        RECT 27.430 30.300 27.580 37.850 ;
        RECT 28.030 30.300 28.180 37.850 ;
        RECT 28.630 30.300 28.780 37.850 ;
        RECT 29.230 30.300 29.380 37.850 ;
        RECT 29.830 30.300 29.980 37.850 ;
        RECT 34.230 37.550 35.230 38.000 ;
        RECT 30.880 37.400 38.580 37.550 ;
        RECT 34.230 36.950 35.230 37.400 ;
        RECT 30.880 36.800 38.580 36.950 ;
        RECT 34.230 36.350 35.230 36.800 ;
        RECT 30.880 36.200 38.580 36.350 ;
        RECT 34.230 35.750 35.230 36.200 ;
        RECT 30.880 35.600 38.580 35.750 ;
        RECT 34.230 35.150 35.230 35.600 ;
        RECT 30.880 35.000 38.580 35.150 ;
        RECT 34.230 34.550 35.230 35.000 ;
        RECT 30.880 34.400 38.580 34.550 ;
        RECT 34.230 33.950 35.230 34.400 ;
        RECT 30.880 33.800 38.580 33.950 ;
        RECT 34.230 33.350 35.230 33.800 ;
        RECT 30.880 33.200 38.580 33.350 ;
        RECT 34.230 32.750 35.230 33.200 ;
        RECT 30.880 32.600 38.580 32.750 ;
        RECT 34.230 32.150 35.230 32.600 ;
        RECT 30.880 32.000 38.580 32.150 ;
        RECT 34.230 31.550 35.230 32.000 ;
        RECT 30.880 31.400 38.580 31.550 ;
        RECT 34.230 30.950 35.230 31.400 ;
        RECT 30.880 30.800 38.580 30.950 ;
        RECT 34.230 30.300 35.230 30.800 ;
        RECT 39.480 30.300 39.630 37.850 ;
        RECT 40.080 30.300 40.230 37.850 ;
        RECT 40.680 30.300 40.830 37.850 ;
        RECT 41.280 30.300 41.430 37.850 ;
        RECT 41.880 30.300 42.030 37.850 ;
        RECT 42.480 30.300 42.630 37.850 ;
        RECT 42.780 33.200 43.530 35.000 ;
        RECT 45.930 33.200 46.680 35.000 ;
        RECT 42.780 30.450 46.680 33.200 ;
        RECT 42.780 30.300 43.930 30.450 ;
        RECT 25.530 29.700 43.930 30.300 ;
        RECT 25.530 29.550 26.680 29.700 ;
        RECT 22.780 26.800 26.680 29.550 ;
        RECT 22.780 25.050 23.530 26.800 ;
        RECT 25.930 25.050 26.680 26.800 ;
        RECT 26.830 22.150 26.980 29.700 ;
        RECT 27.430 22.150 27.580 29.700 ;
        RECT 28.030 22.150 28.180 29.700 ;
        RECT 28.630 22.150 28.780 29.700 ;
        RECT 29.230 22.150 29.380 29.700 ;
        RECT 29.830 22.150 29.980 29.700 ;
        RECT 34.230 29.200 35.230 29.700 ;
        RECT 30.880 29.050 38.580 29.200 ;
        RECT 34.230 28.600 35.230 29.050 ;
        RECT 30.880 28.450 38.580 28.600 ;
        RECT 34.230 28.000 35.230 28.450 ;
        RECT 30.880 27.850 38.580 28.000 ;
        RECT 34.230 27.400 35.230 27.850 ;
        RECT 30.880 27.250 38.580 27.400 ;
        RECT 34.230 26.800 35.230 27.250 ;
        RECT 30.880 26.650 38.580 26.800 ;
        RECT 34.230 26.200 35.230 26.650 ;
        RECT 30.880 26.050 38.580 26.200 ;
        RECT 34.230 25.600 35.230 26.050 ;
        RECT 30.880 25.450 38.580 25.600 ;
        RECT 34.230 25.000 35.230 25.450 ;
        RECT 30.880 24.850 38.580 25.000 ;
        RECT 34.230 24.400 35.230 24.850 ;
        RECT 30.880 24.250 38.580 24.400 ;
        RECT 34.230 23.800 35.230 24.250 ;
        RECT 30.880 23.650 38.580 23.800 ;
        RECT 34.230 23.200 35.230 23.650 ;
        RECT 30.880 23.050 38.580 23.200 ;
        RECT 34.230 22.600 35.230 23.050 ;
        RECT 30.880 22.450 38.580 22.600 ;
        RECT 34.230 22.000 35.230 22.450 ;
        RECT 39.480 22.150 39.630 29.700 ;
        RECT 40.080 22.150 40.230 29.700 ;
        RECT 40.680 22.150 40.830 29.700 ;
        RECT 41.280 22.150 41.430 29.700 ;
        RECT 41.880 22.150 42.030 29.700 ;
        RECT 42.480 22.150 42.630 29.700 ;
        RECT 42.780 29.550 43.930 29.700 ;
        RECT 44.580 29.550 44.880 30.450 ;
        RECT 45.530 30.300 46.680 30.450 ;
        RECT 46.830 30.300 46.980 37.850 ;
        RECT 47.430 30.300 47.580 37.850 ;
        RECT 48.030 30.300 48.180 37.850 ;
        RECT 48.630 30.300 48.780 37.850 ;
        RECT 49.230 30.300 49.380 37.850 ;
        RECT 49.830 30.300 49.980 37.850 ;
        RECT 54.230 37.550 55.230 38.000 ;
        RECT 50.880 37.400 58.580 37.550 ;
        RECT 54.230 36.950 55.230 37.400 ;
        RECT 50.880 36.800 58.580 36.950 ;
        RECT 54.230 36.350 55.230 36.800 ;
        RECT 50.880 36.200 58.580 36.350 ;
        RECT 54.230 35.750 55.230 36.200 ;
        RECT 50.880 35.600 58.580 35.750 ;
        RECT 54.230 35.150 55.230 35.600 ;
        RECT 50.880 35.000 58.580 35.150 ;
        RECT 54.230 34.550 55.230 35.000 ;
        RECT 50.880 34.400 58.580 34.550 ;
        RECT 54.230 33.950 55.230 34.400 ;
        RECT 50.880 33.800 58.580 33.950 ;
        RECT 54.230 33.350 55.230 33.800 ;
        RECT 50.880 33.200 58.580 33.350 ;
        RECT 54.230 32.750 55.230 33.200 ;
        RECT 50.880 32.600 58.580 32.750 ;
        RECT 54.230 32.150 55.230 32.600 ;
        RECT 50.880 32.000 58.580 32.150 ;
        RECT 54.230 31.550 55.230 32.000 ;
        RECT 50.880 31.400 58.580 31.550 ;
        RECT 54.230 30.950 55.230 31.400 ;
        RECT 50.880 30.800 58.580 30.950 ;
        RECT 54.230 30.300 55.230 30.800 ;
        RECT 59.480 30.300 59.630 37.850 ;
        RECT 60.080 30.300 60.230 37.850 ;
        RECT 60.680 30.300 60.830 37.850 ;
        RECT 61.280 30.300 61.430 37.850 ;
        RECT 61.880 30.300 62.030 37.850 ;
        RECT 62.480 30.300 62.630 37.850 ;
        RECT 62.780 33.200 63.530 35.000 ;
        RECT 65.930 33.200 66.680 35.000 ;
        RECT 62.780 30.450 66.680 33.200 ;
        RECT 62.780 30.300 63.930 30.450 ;
        RECT 45.530 29.700 63.930 30.300 ;
        RECT 45.530 29.550 46.680 29.700 ;
        RECT 42.780 26.800 46.680 29.550 ;
        RECT 42.780 25.050 43.530 26.800 ;
        RECT 45.930 25.050 46.680 26.800 ;
        RECT 46.830 22.150 46.980 29.700 ;
        RECT 47.430 22.150 47.580 29.700 ;
        RECT 48.030 22.150 48.180 29.700 ;
        RECT 48.630 22.150 48.780 29.700 ;
        RECT 49.230 22.150 49.380 29.700 ;
        RECT 49.830 22.150 49.980 29.700 ;
        RECT 54.230 29.200 55.230 29.700 ;
        RECT 50.880 29.050 58.580 29.200 ;
        RECT 54.230 28.600 55.230 29.050 ;
        RECT 50.880 28.450 58.580 28.600 ;
        RECT 54.230 28.000 55.230 28.450 ;
        RECT 50.880 27.850 58.580 28.000 ;
        RECT 54.230 27.400 55.230 27.850 ;
        RECT 50.880 27.250 58.580 27.400 ;
        RECT 54.230 26.800 55.230 27.250 ;
        RECT 50.880 26.650 58.580 26.800 ;
        RECT 54.230 26.200 55.230 26.650 ;
        RECT 50.880 26.050 58.580 26.200 ;
        RECT 54.230 25.600 55.230 26.050 ;
        RECT 50.880 25.450 58.580 25.600 ;
        RECT 54.230 25.000 55.230 25.450 ;
        RECT 50.880 24.850 58.580 25.000 ;
        RECT 54.230 24.400 55.230 24.850 ;
        RECT 50.880 24.250 58.580 24.400 ;
        RECT 54.230 23.800 55.230 24.250 ;
        RECT 50.880 23.650 58.580 23.800 ;
        RECT 54.230 23.200 55.230 23.650 ;
        RECT 50.880 23.050 58.580 23.200 ;
        RECT 54.230 22.600 55.230 23.050 ;
        RECT 50.880 22.450 58.580 22.600 ;
        RECT 54.230 22.000 55.230 22.450 ;
        RECT 59.480 22.150 59.630 29.700 ;
        RECT 60.080 22.150 60.230 29.700 ;
        RECT 60.680 22.150 60.830 29.700 ;
        RECT 61.280 22.150 61.430 29.700 ;
        RECT 61.880 22.150 62.030 29.700 ;
        RECT 62.480 22.150 62.630 29.700 ;
        RECT 62.780 29.550 63.930 29.700 ;
        RECT 64.580 29.550 64.880 30.450 ;
        RECT 65.530 30.300 66.680 30.450 ;
        RECT 66.830 30.300 66.980 37.850 ;
        RECT 67.430 30.300 67.580 37.850 ;
        RECT 68.030 30.300 68.180 37.850 ;
        RECT 68.630 30.300 68.780 37.850 ;
        RECT 69.230 30.300 69.380 37.850 ;
        RECT 69.830 30.300 69.980 37.850 ;
        RECT 74.230 37.550 75.230 38.000 ;
        RECT 70.880 37.400 78.580 37.550 ;
        RECT 74.230 36.950 75.230 37.400 ;
        RECT 70.880 36.800 78.580 36.950 ;
        RECT 74.230 36.350 75.230 36.800 ;
        RECT 70.880 36.200 78.580 36.350 ;
        RECT 74.230 35.750 75.230 36.200 ;
        RECT 70.880 35.600 78.580 35.750 ;
        RECT 74.230 35.150 75.230 35.600 ;
        RECT 70.880 35.000 78.580 35.150 ;
        RECT 74.230 34.550 75.230 35.000 ;
        RECT 70.880 34.400 78.580 34.550 ;
        RECT 74.230 33.950 75.230 34.400 ;
        RECT 70.880 33.800 78.580 33.950 ;
        RECT 74.230 33.350 75.230 33.800 ;
        RECT 70.880 33.200 78.580 33.350 ;
        RECT 74.230 32.750 75.230 33.200 ;
        RECT 70.880 32.600 78.580 32.750 ;
        RECT 74.230 32.150 75.230 32.600 ;
        RECT 70.880 32.000 78.580 32.150 ;
        RECT 74.230 31.550 75.230 32.000 ;
        RECT 70.880 31.400 78.580 31.550 ;
        RECT 74.230 30.950 75.230 31.400 ;
        RECT 70.880 30.800 78.580 30.950 ;
        RECT 74.230 30.300 75.230 30.800 ;
        RECT 79.480 30.300 79.630 37.850 ;
        RECT 80.080 30.300 80.230 37.850 ;
        RECT 80.680 30.300 80.830 37.850 ;
        RECT 81.280 30.300 81.430 37.850 ;
        RECT 81.880 30.300 82.030 37.850 ;
        RECT 82.480 30.300 82.630 37.850 ;
        RECT 82.780 33.200 83.530 35.000 ;
        RECT 85.930 33.200 86.680 35.000 ;
        RECT 82.780 30.450 86.680 33.200 ;
        RECT 82.780 30.300 83.930 30.450 ;
        RECT 65.530 29.700 83.930 30.300 ;
        RECT 65.530 29.550 66.680 29.700 ;
        RECT 62.780 26.800 66.680 29.550 ;
        RECT 62.780 25.050 63.530 26.800 ;
        RECT 65.930 25.050 66.680 26.800 ;
        RECT 66.830 22.150 66.980 29.700 ;
        RECT 67.430 22.150 67.580 29.700 ;
        RECT 68.030 22.150 68.180 29.700 ;
        RECT 68.630 22.150 68.780 29.700 ;
        RECT 69.230 22.150 69.380 29.700 ;
        RECT 69.830 22.150 69.980 29.700 ;
        RECT 74.230 29.200 75.230 29.700 ;
        RECT 70.880 29.050 78.580 29.200 ;
        RECT 74.230 28.600 75.230 29.050 ;
        RECT 70.880 28.450 78.580 28.600 ;
        RECT 74.230 28.000 75.230 28.450 ;
        RECT 70.880 27.850 78.580 28.000 ;
        RECT 74.230 27.400 75.230 27.850 ;
        RECT 70.880 27.250 78.580 27.400 ;
        RECT 74.230 26.800 75.230 27.250 ;
        RECT 70.880 26.650 78.580 26.800 ;
        RECT 74.230 26.200 75.230 26.650 ;
        RECT 70.880 26.050 78.580 26.200 ;
        RECT 74.230 25.600 75.230 26.050 ;
        RECT 70.880 25.450 78.580 25.600 ;
        RECT 74.230 25.000 75.230 25.450 ;
        RECT 70.880 24.850 78.580 25.000 ;
        RECT 74.230 24.400 75.230 24.850 ;
        RECT 70.880 24.250 78.580 24.400 ;
        RECT 74.230 23.800 75.230 24.250 ;
        RECT 70.880 23.650 78.580 23.800 ;
        RECT 74.230 23.200 75.230 23.650 ;
        RECT 70.880 23.050 78.580 23.200 ;
        RECT 74.230 22.600 75.230 23.050 ;
        RECT 70.880 22.450 78.580 22.600 ;
        RECT 74.230 22.000 75.230 22.450 ;
        RECT 79.480 22.150 79.630 29.700 ;
        RECT 80.080 22.150 80.230 29.700 ;
        RECT 80.680 22.150 80.830 29.700 ;
        RECT 81.280 22.150 81.430 29.700 ;
        RECT 81.880 22.150 82.030 29.700 ;
        RECT 82.480 22.150 82.630 29.700 ;
        RECT 82.780 29.550 83.930 29.700 ;
        RECT 84.580 29.550 84.880 30.450 ;
        RECT 85.530 30.300 86.680 30.450 ;
        RECT 86.830 30.300 86.980 37.850 ;
        RECT 87.430 30.300 87.580 37.850 ;
        RECT 88.030 30.300 88.180 37.850 ;
        RECT 88.630 30.300 88.780 37.850 ;
        RECT 89.230 30.300 89.380 37.850 ;
        RECT 89.830 30.300 89.980 37.850 ;
        RECT 94.230 37.550 95.230 38.000 ;
        RECT 90.880 37.400 98.580 37.550 ;
        RECT 94.230 36.950 95.230 37.400 ;
        RECT 90.880 36.800 98.580 36.950 ;
        RECT 94.230 36.350 95.230 36.800 ;
        RECT 90.880 36.200 98.580 36.350 ;
        RECT 94.230 35.750 95.230 36.200 ;
        RECT 90.880 35.600 98.580 35.750 ;
        RECT 94.230 35.150 95.230 35.600 ;
        RECT 90.880 35.000 98.580 35.150 ;
        RECT 94.230 34.550 95.230 35.000 ;
        RECT 90.880 34.400 98.580 34.550 ;
        RECT 94.230 33.950 95.230 34.400 ;
        RECT 90.880 33.800 98.580 33.950 ;
        RECT 94.230 33.350 95.230 33.800 ;
        RECT 90.880 33.200 98.580 33.350 ;
        RECT 94.230 32.750 95.230 33.200 ;
        RECT 90.880 32.600 98.580 32.750 ;
        RECT 94.230 32.150 95.230 32.600 ;
        RECT 90.880 32.000 98.580 32.150 ;
        RECT 94.230 31.550 95.230 32.000 ;
        RECT 90.880 31.400 98.580 31.550 ;
        RECT 94.230 30.950 95.230 31.400 ;
        RECT 90.880 30.800 98.580 30.950 ;
        RECT 94.230 30.300 95.230 30.800 ;
        RECT 99.480 30.300 99.630 37.850 ;
        RECT 100.080 30.300 100.230 37.850 ;
        RECT 100.680 30.300 100.830 37.850 ;
        RECT 101.280 30.300 101.430 37.850 ;
        RECT 101.880 30.300 102.030 37.850 ;
        RECT 102.480 30.300 102.630 37.850 ;
        RECT 102.780 33.200 103.530 35.000 ;
        RECT 102.780 31.525 104.730 33.200 ;
        RECT 102.780 30.450 111.850 31.525 ;
        RECT 102.780 30.300 103.930 30.450 ;
        RECT 85.530 29.700 103.930 30.300 ;
        RECT 85.530 29.550 86.680 29.700 ;
        RECT 82.780 26.800 86.680 29.550 ;
        RECT 82.780 25.050 83.530 26.800 ;
        RECT 85.930 25.050 86.680 26.800 ;
        RECT 86.830 22.150 86.980 29.700 ;
        RECT 87.430 22.150 87.580 29.700 ;
        RECT 88.030 22.150 88.180 29.700 ;
        RECT 88.630 22.150 88.780 29.700 ;
        RECT 89.230 22.150 89.380 29.700 ;
        RECT 89.830 22.150 89.980 29.700 ;
        RECT 94.230 29.200 95.230 29.700 ;
        RECT 90.880 29.050 98.580 29.200 ;
        RECT 94.230 28.600 95.230 29.050 ;
        RECT 90.880 28.450 98.580 28.600 ;
        RECT 94.230 28.000 95.230 28.450 ;
        RECT 90.880 27.850 98.580 28.000 ;
        RECT 94.230 27.400 95.230 27.850 ;
        RECT 90.880 27.250 98.580 27.400 ;
        RECT 94.230 26.800 95.230 27.250 ;
        RECT 90.880 26.650 98.580 26.800 ;
        RECT 94.230 26.200 95.230 26.650 ;
        RECT 90.880 26.050 98.580 26.200 ;
        RECT 94.230 25.600 95.230 26.050 ;
        RECT 90.880 25.450 98.580 25.600 ;
        RECT 94.230 25.000 95.230 25.450 ;
        RECT 90.880 24.850 98.580 25.000 ;
        RECT 94.230 24.400 95.230 24.850 ;
        RECT 90.880 24.250 98.580 24.400 ;
        RECT 94.230 23.800 95.230 24.250 ;
        RECT 90.880 23.650 98.580 23.800 ;
        RECT 94.230 23.200 95.230 23.650 ;
        RECT 90.880 23.050 98.580 23.200 ;
        RECT 94.230 22.600 95.230 23.050 ;
        RECT 90.880 22.450 98.580 22.600 ;
        RECT 94.230 22.000 95.230 22.450 ;
        RECT 99.480 22.150 99.630 29.700 ;
        RECT 100.080 22.150 100.230 29.700 ;
        RECT 100.680 22.150 100.830 29.700 ;
        RECT 101.280 22.150 101.430 29.700 ;
        RECT 101.880 22.150 102.030 29.700 ;
        RECT 102.480 22.150 102.630 29.700 ;
        RECT 102.780 29.550 103.930 29.700 ;
        RECT 104.580 30.250 111.850 30.450 ;
        RECT 104.580 29.550 104.730 30.250 ;
        RECT 102.780 26.800 104.730 29.550 ;
        RECT 102.780 25.050 103.530 26.800 ;
        RECT 10.880 21.850 18.580 22.000 ;
        RECT 30.880 21.850 38.580 22.000 ;
        RECT 50.880 21.850 58.580 22.000 ;
        RECT 70.880 21.850 78.580 22.000 ;
        RECT 90.880 21.850 98.580 22.000 ;
        RECT 14.230 21.200 15.230 21.850 ;
        RECT 34.230 21.200 35.230 21.850 ;
        RECT 54.230 21.200 55.230 21.850 ;
        RECT 74.230 21.200 75.230 21.850 ;
        RECT 94.230 21.200 95.230 21.850 ;
        RECT 11.530 18.800 17.930 21.200 ;
        RECT 31.530 18.800 37.930 21.200 ;
        RECT 51.530 18.800 57.930 21.200 ;
        RECT 71.530 18.800 77.930 21.200 ;
        RECT 91.530 18.800 97.930 21.200 ;
        RECT 14.230 18.150 15.230 18.800 ;
        RECT 34.230 18.150 35.230 18.800 ;
        RECT 54.230 18.150 55.230 18.800 ;
        RECT 74.230 18.150 75.230 18.800 ;
        RECT 94.230 18.150 95.230 18.800 ;
        RECT 10.880 18.000 18.580 18.150 ;
        RECT 30.880 18.000 38.580 18.150 ;
        RECT 50.880 18.000 58.580 18.150 ;
        RECT 70.880 18.000 78.580 18.150 ;
        RECT 90.880 18.000 98.580 18.150 ;
        RECT 5.930 13.200 6.680 15.000 ;
        RECT 4.730 10.450 6.680 13.200 ;
        RECT 4.730 9.550 4.880 10.450 ;
        RECT 5.530 10.300 6.680 10.450 ;
        RECT 6.830 10.300 6.980 17.850 ;
        RECT 7.430 10.300 7.580 17.850 ;
        RECT 8.030 10.300 8.180 17.850 ;
        RECT 8.630 10.300 8.780 17.850 ;
        RECT 9.230 10.300 9.380 17.850 ;
        RECT 9.830 10.300 9.980 17.850 ;
        RECT 14.230 17.550 15.230 18.000 ;
        RECT 10.880 17.400 18.580 17.550 ;
        RECT 14.230 16.950 15.230 17.400 ;
        RECT 10.880 16.800 18.580 16.950 ;
        RECT 14.230 16.350 15.230 16.800 ;
        RECT 10.880 16.200 18.580 16.350 ;
        RECT 14.230 15.750 15.230 16.200 ;
        RECT 10.880 15.600 18.580 15.750 ;
        RECT 14.230 15.150 15.230 15.600 ;
        RECT 10.880 15.000 18.580 15.150 ;
        RECT 14.230 14.550 15.230 15.000 ;
        RECT 10.880 14.400 18.580 14.550 ;
        RECT 14.230 13.950 15.230 14.400 ;
        RECT 10.880 13.800 18.580 13.950 ;
        RECT 14.230 13.350 15.230 13.800 ;
        RECT 10.880 13.200 18.580 13.350 ;
        RECT 14.230 12.750 15.230 13.200 ;
        RECT 10.880 12.600 18.580 12.750 ;
        RECT 14.230 12.150 15.230 12.600 ;
        RECT 10.880 12.000 18.580 12.150 ;
        RECT 14.230 11.550 15.230 12.000 ;
        RECT 10.880 11.400 18.580 11.550 ;
        RECT 14.230 10.950 15.230 11.400 ;
        RECT 10.880 10.800 18.580 10.950 ;
        RECT 14.230 10.300 15.230 10.800 ;
        RECT 19.480 10.300 19.630 17.850 ;
        RECT 20.080 10.300 20.230 17.850 ;
        RECT 20.680 10.300 20.830 17.850 ;
        RECT 21.280 10.300 21.430 17.850 ;
        RECT 21.880 10.300 22.030 17.850 ;
        RECT 22.480 10.300 22.630 17.850 ;
        RECT 22.780 13.200 23.530 15.000 ;
        RECT 25.930 13.200 26.680 15.000 ;
        RECT 22.780 10.450 26.680 13.200 ;
        RECT 22.780 10.300 23.930 10.450 ;
        RECT 5.530 9.700 23.930 10.300 ;
        RECT 5.530 9.550 6.680 9.700 ;
        RECT 4.730 6.800 6.680 9.550 ;
        RECT 5.930 5.050 6.680 6.800 ;
        RECT 6.830 2.150 6.980 9.700 ;
        RECT 7.430 2.150 7.580 9.700 ;
        RECT 8.030 2.150 8.180 9.700 ;
        RECT 8.630 2.150 8.780 9.700 ;
        RECT 9.230 2.150 9.380 9.700 ;
        RECT 9.830 2.150 9.980 9.700 ;
        RECT 14.230 9.200 15.230 9.700 ;
        RECT 10.880 9.050 18.580 9.200 ;
        RECT 14.230 8.600 15.230 9.050 ;
        RECT 10.880 8.450 18.580 8.600 ;
        RECT 14.230 8.000 15.230 8.450 ;
        RECT 10.880 7.850 18.580 8.000 ;
        RECT 14.230 7.400 15.230 7.850 ;
        RECT 10.880 7.250 18.580 7.400 ;
        RECT 14.230 6.800 15.230 7.250 ;
        RECT 10.880 6.650 18.580 6.800 ;
        RECT 14.230 6.200 15.230 6.650 ;
        RECT 10.880 6.050 18.580 6.200 ;
        RECT 14.230 5.600 15.230 6.050 ;
        RECT 10.880 5.450 18.580 5.600 ;
        RECT 14.230 5.000 15.230 5.450 ;
        RECT 10.880 4.850 18.580 5.000 ;
        RECT 14.230 4.400 15.230 4.850 ;
        RECT 10.880 4.250 18.580 4.400 ;
        RECT 14.230 3.800 15.230 4.250 ;
        RECT 10.880 3.650 18.580 3.800 ;
        RECT 14.230 3.200 15.230 3.650 ;
        RECT 10.880 3.050 18.580 3.200 ;
        RECT 14.230 2.600 15.230 3.050 ;
        RECT 10.880 2.450 18.580 2.600 ;
        RECT 14.230 2.000 15.230 2.450 ;
        RECT 19.480 2.150 19.630 9.700 ;
        RECT 20.080 2.150 20.230 9.700 ;
        RECT 20.680 2.150 20.830 9.700 ;
        RECT 21.280 2.150 21.430 9.700 ;
        RECT 21.880 2.150 22.030 9.700 ;
        RECT 22.480 2.150 22.630 9.700 ;
        RECT 22.780 9.550 23.930 9.700 ;
        RECT 24.580 9.550 24.880 10.450 ;
        RECT 25.530 10.300 26.680 10.450 ;
        RECT 26.830 10.300 26.980 17.850 ;
        RECT 27.430 10.300 27.580 17.850 ;
        RECT 28.030 10.300 28.180 17.850 ;
        RECT 28.630 10.300 28.780 17.850 ;
        RECT 29.230 10.300 29.380 17.850 ;
        RECT 29.830 10.300 29.980 17.850 ;
        RECT 34.230 17.550 35.230 18.000 ;
        RECT 30.880 17.400 38.580 17.550 ;
        RECT 34.230 16.950 35.230 17.400 ;
        RECT 30.880 16.800 38.580 16.950 ;
        RECT 34.230 16.350 35.230 16.800 ;
        RECT 30.880 16.200 38.580 16.350 ;
        RECT 34.230 15.750 35.230 16.200 ;
        RECT 30.880 15.600 38.580 15.750 ;
        RECT 34.230 15.150 35.230 15.600 ;
        RECT 30.880 15.000 38.580 15.150 ;
        RECT 34.230 14.550 35.230 15.000 ;
        RECT 30.880 14.400 38.580 14.550 ;
        RECT 34.230 13.950 35.230 14.400 ;
        RECT 30.880 13.800 38.580 13.950 ;
        RECT 34.230 13.350 35.230 13.800 ;
        RECT 30.880 13.200 38.580 13.350 ;
        RECT 34.230 12.750 35.230 13.200 ;
        RECT 30.880 12.600 38.580 12.750 ;
        RECT 34.230 12.150 35.230 12.600 ;
        RECT 30.880 12.000 38.580 12.150 ;
        RECT 34.230 11.550 35.230 12.000 ;
        RECT 30.880 11.400 38.580 11.550 ;
        RECT 34.230 10.950 35.230 11.400 ;
        RECT 30.880 10.800 38.580 10.950 ;
        RECT 34.230 10.300 35.230 10.800 ;
        RECT 39.480 10.300 39.630 17.850 ;
        RECT 40.080 10.300 40.230 17.850 ;
        RECT 40.680 10.300 40.830 17.850 ;
        RECT 41.280 10.300 41.430 17.850 ;
        RECT 41.880 10.300 42.030 17.850 ;
        RECT 42.480 10.300 42.630 17.850 ;
        RECT 42.780 13.200 43.530 15.000 ;
        RECT 45.930 13.200 46.680 15.000 ;
        RECT 42.780 10.450 46.680 13.200 ;
        RECT 42.780 10.300 43.930 10.450 ;
        RECT 25.530 9.700 43.930 10.300 ;
        RECT 25.530 9.550 26.680 9.700 ;
        RECT 22.780 6.800 26.680 9.550 ;
        RECT 22.780 5.050 23.530 6.800 ;
        RECT 25.930 5.050 26.680 6.800 ;
        RECT 26.830 2.150 26.980 9.700 ;
        RECT 27.430 2.150 27.580 9.700 ;
        RECT 28.030 2.150 28.180 9.700 ;
        RECT 28.630 2.150 28.780 9.700 ;
        RECT 29.230 2.150 29.380 9.700 ;
        RECT 29.830 2.150 29.980 9.700 ;
        RECT 34.230 9.200 35.230 9.700 ;
        RECT 30.880 9.050 38.580 9.200 ;
        RECT 34.230 8.600 35.230 9.050 ;
        RECT 30.880 8.450 38.580 8.600 ;
        RECT 34.230 8.000 35.230 8.450 ;
        RECT 30.880 7.850 38.580 8.000 ;
        RECT 34.230 7.400 35.230 7.850 ;
        RECT 30.880 7.250 38.580 7.400 ;
        RECT 34.230 6.800 35.230 7.250 ;
        RECT 30.880 6.650 38.580 6.800 ;
        RECT 34.230 6.200 35.230 6.650 ;
        RECT 30.880 6.050 38.580 6.200 ;
        RECT 34.230 5.600 35.230 6.050 ;
        RECT 30.880 5.450 38.580 5.600 ;
        RECT 34.230 5.000 35.230 5.450 ;
        RECT 30.880 4.850 38.580 5.000 ;
        RECT 34.230 4.400 35.230 4.850 ;
        RECT 30.880 4.250 38.580 4.400 ;
        RECT 34.230 3.800 35.230 4.250 ;
        RECT 30.880 3.650 38.580 3.800 ;
        RECT 34.230 3.200 35.230 3.650 ;
        RECT 30.880 3.050 38.580 3.200 ;
        RECT 34.230 2.600 35.230 3.050 ;
        RECT 30.880 2.450 38.580 2.600 ;
        RECT 34.230 2.000 35.230 2.450 ;
        RECT 39.480 2.150 39.630 9.700 ;
        RECT 40.080 2.150 40.230 9.700 ;
        RECT 40.680 2.150 40.830 9.700 ;
        RECT 41.280 2.150 41.430 9.700 ;
        RECT 41.880 2.150 42.030 9.700 ;
        RECT 42.480 2.150 42.630 9.700 ;
        RECT 42.780 9.550 43.930 9.700 ;
        RECT 44.580 9.550 44.880 10.450 ;
        RECT 45.530 10.300 46.680 10.450 ;
        RECT 46.830 10.300 46.980 17.850 ;
        RECT 47.430 10.300 47.580 17.850 ;
        RECT 48.030 10.300 48.180 17.850 ;
        RECT 48.630 10.300 48.780 17.850 ;
        RECT 49.230 10.300 49.380 17.850 ;
        RECT 49.830 10.300 49.980 17.850 ;
        RECT 54.230 17.550 55.230 18.000 ;
        RECT 50.880 17.400 58.580 17.550 ;
        RECT 54.230 16.950 55.230 17.400 ;
        RECT 50.880 16.800 58.580 16.950 ;
        RECT 54.230 16.350 55.230 16.800 ;
        RECT 50.880 16.200 58.580 16.350 ;
        RECT 54.230 15.750 55.230 16.200 ;
        RECT 50.880 15.600 58.580 15.750 ;
        RECT 54.230 15.150 55.230 15.600 ;
        RECT 50.880 15.000 58.580 15.150 ;
        RECT 54.230 14.550 55.230 15.000 ;
        RECT 50.880 14.400 58.580 14.550 ;
        RECT 54.230 13.950 55.230 14.400 ;
        RECT 50.880 13.800 58.580 13.950 ;
        RECT 54.230 13.350 55.230 13.800 ;
        RECT 50.880 13.200 58.580 13.350 ;
        RECT 54.230 12.750 55.230 13.200 ;
        RECT 50.880 12.600 58.580 12.750 ;
        RECT 54.230 12.150 55.230 12.600 ;
        RECT 50.880 12.000 58.580 12.150 ;
        RECT 54.230 11.550 55.230 12.000 ;
        RECT 50.880 11.400 58.580 11.550 ;
        RECT 54.230 10.950 55.230 11.400 ;
        RECT 50.880 10.800 58.580 10.950 ;
        RECT 54.230 10.300 55.230 10.800 ;
        RECT 59.480 10.300 59.630 17.850 ;
        RECT 60.080 10.300 60.230 17.850 ;
        RECT 60.680 10.300 60.830 17.850 ;
        RECT 61.280 10.300 61.430 17.850 ;
        RECT 61.880 10.300 62.030 17.850 ;
        RECT 62.480 10.300 62.630 17.850 ;
        RECT 62.780 13.200 63.530 15.000 ;
        RECT 65.930 13.200 66.680 15.000 ;
        RECT 62.780 10.450 66.680 13.200 ;
        RECT 62.780 10.300 63.930 10.450 ;
        RECT 45.530 9.700 63.930 10.300 ;
        RECT 45.530 9.550 46.680 9.700 ;
        RECT 42.780 6.800 46.680 9.550 ;
        RECT 42.780 5.050 43.530 6.800 ;
        RECT 45.930 5.050 46.680 6.800 ;
        RECT 46.830 2.150 46.980 9.700 ;
        RECT 47.430 2.150 47.580 9.700 ;
        RECT 48.030 2.150 48.180 9.700 ;
        RECT 48.630 2.150 48.780 9.700 ;
        RECT 49.230 2.150 49.380 9.700 ;
        RECT 49.830 2.150 49.980 9.700 ;
        RECT 54.230 9.200 55.230 9.700 ;
        RECT 50.880 9.050 58.580 9.200 ;
        RECT 54.230 8.600 55.230 9.050 ;
        RECT 50.880 8.450 58.580 8.600 ;
        RECT 54.230 8.000 55.230 8.450 ;
        RECT 50.880 7.850 58.580 8.000 ;
        RECT 54.230 7.400 55.230 7.850 ;
        RECT 50.880 7.250 58.580 7.400 ;
        RECT 54.230 6.800 55.230 7.250 ;
        RECT 50.880 6.650 58.580 6.800 ;
        RECT 54.230 6.200 55.230 6.650 ;
        RECT 50.880 6.050 58.580 6.200 ;
        RECT 54.230 5.600 55.230 6.050 ;
        RECT 50.880 5.450 58.580 5.600 ;
        RECT 54.230 5.000 55.230 5.450 ;
        RECT 50.880 4.850 58.580 5.000 ;
        RECT 54.230 4.400 55.230 4.850 ;
        RECT 50.880 4.250 58.580 4.400 ;
        RECT 54.230 3.800 55.230 4.250 ;
        RECT 50.880 3.650 58.580 3.800 ;
        RECT 54.230 3.200 55.230 3.650 ;
        RECT 50.880 3.050 58.580 3.200 ;
        RECT 54.230 2.600 55.230 3.050 ;
        RECT 50.880 2.450 58.580 2.600 ;
        RECT 54.230 2.000 55.230 2.450 ;
        RECT 59.480 2.150 59.630 9.700 ;
        RECT 60.080 2.150 60.230 9.700 ;
        RECT 60.680 2.150 60.830 9.700 ;
        RECT 61.280 2.150 61.430 9.700 ;
        RECT 61.880 2.150 62.030 9.700 ;
        RECT 62.480 2.150 62.630 9.700 ;
        RECT 62.780 9.550 63.930 9.700 ;
        RECT 64.580 9.550 64.880 10.450 ;
        RECT 65.530 10.300 66.680 10.450 ;
        RECT 66.830 10.300 66.980 17.850 ;
        RECT 67.430 10.300 67.580 17.850 ;
        RECT 68.030 10.300 68.180 17.850 ;
        RECT 68.630 10.300 68.780 17.850 ;
        RECT 69.230 10.300 69.380 17.850 ;
        RECT 69.830 10.300 69.980 17.850 ;
        RECT 74.230 17.550 75.230 18.000 ;
        RECT 70.880 17.400 78.580 17.550 ;
        RECT 74.230 16.950 75.230 17.400 ;
        RECT 70.880 16.800 78.580 16.950 ;
        RECT 74.230 16.350 75.230 16.800 ;
        RECT 70.880 16.200 78.580 16.350 ;
        RECT 74.230 15.750 75.230 16.200 ;
        RECT 70.880 15.600 78.580 15.750 ;
        RECT 74.230 15.150 75.230 15.600 ;
        RECT 70.880 15.000 78.580 15.150 ;
        RECT 74.230 14.550 75.230 15.000 ;
        RECT 70.880 14.400 78.580 14.550 ;
        RECT 74.230 13.950 75.230 14.400 ;
        RECT 70.880 13.800 78.580 13.950 ;
        RECT 74.230 13.350 75.230 13.800 ;
        RECT 70.880 13.200 78.580 13.350 ;
        RECT 74.230 12.750 75.230 13.200 ;
        RECT 70.880 12.600 78.580 12.750 ;
        RECT 74.230 12.150 75.230 12.600 ;
        RECT 70.880 12.000 78.580 12.150 ;
        RECT 74.230 11.550 75.230 12.000 ;
        RECT 70.880 11.400 78.580 11.550 ;
        RECT 74.230 10.950 75.230 11.400 ;
        RECT 70.880 10.800 78.580 10.950 ;
        RECT 74.230 10.300 75.230 10.800 ;
        RECT 79.480 10.300 79.630 17.850 ;
        RECT 80.080 10.300 80.230 17.850 ;
        RECT 80.680 10.300 80.830 17.850 ;
        RECT 81.280 10.300 81.430 17.850 ;
        RECT 81.880 10.300 82.030 17.850 ;
        RECT 82.480 10.300 82.630 17.850 ;
        RECT 82.780 13.200 83.530 15.000 ;
        RECT 85.930 13.200 86.680 15.000 ;
        RECT 82.780 10.450 86.680 13.200 ;
        RECT 82.780 10.300 83.930 10.450 ;
        RECT 65.530 9.700 83.930 10.300 ;
        RECT 65.530 9.550 66.680 9.700 ;
        RECT 62.780 6.800 66.680 9.550 ;
        RECT 62.780 5.050 63.530 6.800 ;
        RECT 65.930 5.050 66.680 6.800 ;
        RECT 66.830 2.150 66.980 9.700 ;
        RECT 67.430 2.150 67.580 9.700 ;
        RECT 68.030 2.150 68.180 9.700 ;
        RECT 68.630 2.150 68.780 9.700 ;
        RECT 69.230 2.150 69.380 9.700 ;
        RECT 69.830 2.150 69.980 9.700 ;
        RECT 74.230 9.200 75.230 9.700 ;
        RECT 70.880 9.050 78.580 9.200 ;
        RECT 74.230 8.600 75.230 9.050 ;
        RECT 70.880 8.450 78.580 8.600 ;
        RECT 74.230 8.000 75.230 8.450 ;
        RECT 70.880 7.850 78.580 8.000 ;
        RECT 74.230 7.400 75.230 7.850 ;
        RECT 70.880 7.250 78.580 7.400 ;
        RECT 74.230 6.800 75.230 7.250 ;
        RECT 70.880 6.650 78.580 6.800 ;
        RECT 74.230 6.200 75.230 6.650 ;
        RECT 70.880 6.050 78.580 6.200 ;
        RECT 74.230 5.600 75.230 6.050 ;
        RECT 70.880 5.450 78.580 5.600 ;
        RECT 74.230 5.000 75.230 5.450 ;
        RECT 70.880 4.850 78.580 5.000 ;
        RECT 74.230 4.400 75.230 4.850 ;
        RECT 70.880 4.250 78.580 4.400 ;
        RECT 74.230 3.800 75.230 4.250 ;
        RECT 70.880 3.650 78.580 3.800 ;
        RECT 74.230 3.200 75.230 3.650 ;
        RECT 70.880 3.050 78.580 3.200 ;
        RECT 74.230 2.600 75.230 3.050 ;
        RECT 70.880 2.450 78.580 2.600 ;
        RECT 74.230 2.000 75.230 2.450 ;
        RECT 79.480 2.150 79.630 9.700 ;
        RECT 80.080 2.150 80.230 9.700 ;
        RECT 80.680 2.150 80.830 9.700 ;
        RECT 81.280 2.150 81.430 9.700 ;
        RECT 81.880 2.150 82.030 9.700 ;
        RECT 82.480 2.150 82.630 9.700 ;
        RECT 82.780 9.550 83.930 9.700 ;
        RECT 84.580 9.550 84.880 10.450 ;
        RECT 85.530 10.300 86.680 10.450 ;
        RECT 86.830 10.300 86.980 17.850 ;
        RECT 87.430 10.300 87.580 17.850 ;
        RECT 88.030 10.300 88.180 17.850 ;
        RECT 88.630 10.300 88.780 17.850 ;
        RECT 89.230 10.300 89.380 17.850 ;
        RECT 89.830 10.300 89.980 17.850 ;
        RECT 94.230 17.550 95.230 18.000 ;
        RECT 90.880 17.400 98.580 17.550 ;
        RECT 94.230 16.950 95.230 17.400 ;
        RECT 90.880 16.800 98.580 16.950 ;
        RECT 94.230 16.350 95.230 16.800 ;
        RECT 90.880 16.200 98.580 16.350 ;
        RECT 94.230 15.750 95.230 16.200 ;
        RECT 90.880 15.600 98.580 15.750 ;
        RECT 94.230 15.150 95.230 15.600 ;
        RECT 90.880 15.000 98.580 15.150 ;
        RECT 94.230 14.550 95.230 15.000 ;
        RECT 90.880 14.400 98.580 14.550 ;
        RECT 94.230 13.950 95.230 14.400 ;
        RECT 90.880 13.800 98.580 13.950 ;
        RECT 94.230 13.350 95.230 13.800 ;
        RECT 90.880 13.200 98.580 13.350 ;
        RECT 94.230 12.750 95.230 13.200 ;
        RECT 90.880 12.600 98.580 12.750 ;
        RECT 94.230 12.150 95.230 12.600 ;
        RECT 90.880 12.000 98.580 12.150 ;
        RECT 94.230 11.550 95.230 12.000 ;
        RECT 90.880 11.400 98.580 11.550 ;
        RECT 94.230 10.950 95.230 11.400 ;
        RECT 90.880 10.800 98.580 10.950 ;
        RECT 94.230 10.300 95.230 10.800 ;
        RECT 99.480 10.300 99.630 17.850 ;
        RECT 100.080 10.300 100.230 17.850 ;
        RECT 100.680 10.300 100.830 17.850 ;
        RECT 101.280 10.300 101.430 17.850 ;
        RECT 101.880 10.300 102.030 17.850 ;
        RECT 102.480 10.300 102.630 17.850 ;
        RECT 102.780 13.200 103.530 15.000 ;
        RECT 102.780 11.525 104.730 13.200 ;
        RECT 102.780 10.450 111.850 11.525 ;
        RECT 102.780 10.300 103.930 10.450 ;
        RECT 85.530 9.700 103.930 10.300 ;
        RECT 85.530 9.550 86.680 9.700 ;
        RECT 82.780 6.800 86.680 9.550 ;
        RECT 82.780 5.050 83.530 6.800 ;
        RECT 85.930 5.050 86.680 6.800 ;
        RECT 86.830 2.150 86.980 9.700 ;
        RECT 87.430 2.150 87.580 9.700 ;
        RECT 88.030 2.150 88.180 9.700 ;
        RECT 88.630 2.150 88.780 9.700 ;
        RECT 89.230 2.150 89.380 9.700 ;
        RECT 89.830 2.150 89.980 9.700 ;
        RECT 94.230 9.200 95.230 9.700 ;
        RECT 90.880 9.050 98.580 9.200 ;
        RECT 94.230 8.600 95.230 9.050 ;
        RECT 90.880 8.450 98.580 8.600 ;
        RECT 94.230 8.000 95.230 8.450 ;
        RECT 90.880 7.850 98.580 8.000 ;
        RECT 94.230 7.400 95.230 7.850 ;
        RECT 90.880 7.250 98.580 7.400 ;
        RECT 94.230 6.800 95.230 7.250 ;
        RECT 90.880 6.650 98.580 6.800 ;
        RECT 94.230 6.200 95.230 6.650 ;
        RECT 90.880 6.050 98.580 6.200 ;
        RECT 94.230 5.600 95.230 6.050 ;
        RECT 90.880 5.450 98.580 5.600 ;
        RECT 94.230 5.000 95.230 5.450 ;
        RECT 90.880 4.850 98.580 5.000 ;
        RECT 94.230 4.400 95.230 4.850 ;
        RECT 90.880 4.250 98.580 4.400 ;
        RECT 94.230 3.800 95.230 4.250 ;
        RECT 90.880 3.650 98.580 3.800 ;
        RECT 94.230 3.200 95.230 3.650 ;
        RECT 90.880 3.050 98.580 3.200 ;
        RECT 94.230 2.600 95.230 3.050 ;
        RECT 90.880 2.450 98.580 2.600 ;
        RECT 94.230 2.000 95.230 2.450 ;
        RECT 99.480 2.150 99.630 9.700 ;
        RECT 100.080 2.150 100.230 9.700 ;
        RECT 100.680 2.150 100.830 9.700 ;
        RECT 101.280 2.150 101.430 9.700 ;
        RECT 101.880 2.150 102.030 9.700 ;
        RECT 102.480 2.150 102.630 9.700 ;
        RECT 102.780 9.550 103.930 9.700 ;
        RECT 104.580 10.250 111.850 10.450 ;
        RECT 104.580 9.550 104.730 10.250 ;
        RECT 102.780 6.800 104.730 9.550 ;
        RECT 102.780 5.050 103.530 6.800 ;
        RECT 10.880 1.850 18.580 2.000 ;
        RECT 30.880 1.850 38.580 2.000 ;
        RECT 50.880 1.850 58.580 2.000 ;
        RECT 70.880 1.850 78.580 2.000 ;
        RECT 90.880 1.850 98.580 2.000 ;
        RECT 14.230 1.200 15.230 1.850 ;
        RECT 34.230 1.200 35.230 1.850 ;
        RECT 54.230 1.200 55.230 1.850 ;
        RECT 74.230 1.200 75.230 1.850 ;
        RECT 94.230 1.200 95.230 1.850 ;
        RECT 11.530 0.000 17.930 1.200 ;
        RECT 31.530 0.000 37.930 1.200 ;
        RECT 51.530 0.000 57.930 1.200 ;
        RECT 71.530 0.000 77.930 1.200 ;
        RECT 91.530 0.000 97.930 1.200 ;
      LAYER via ;
        RECT 11.630 378.900 12.630 379.900 ;
        RECT 12.780 378.900 13.780 379.900 ;
        RECT 13.930 378.900 15.530 379.900 ;
        RECT 15.680 378.900 16.680 379.900 ;
        RECT 16.830 378.900 17.830 379.900 ;
        RECT 31.630 378.900 32.630 379.900 ;
        RECT 32.780 378.900 33.780 379.900 ;
        RECT 33.930 378.900 35.530 379.900 ;
        RECT 35.680 378.900 36.680 379.900 ;
        RECT 36.830 378.900 37.830 379.900 ;
        RECT 51.630 378.900 52.630 379.900 ;
        RECT 52.780 378.900 53.780 379.900 ;
        RECT 53.930 378.900 55.530 379.900 ;
        RECT 55.680 378.900 56.680 379.900 ;
        RECT 56.830 378.900 57.830 379.900 ;
        RECT 71.630 378.900 72.630 379.900 ;
        RECT 72.780 378.900 73.780 379.900 ;
        RECT 73.930 378.900 75.530 379.900 ;
        RECT 75.680 378.900 76.680 379.900 ;
        RECT 76.830 378.900 77.830 379.900 ;
        RECT 91.630 378.900 92.630 379.900 ;
        RECT 92.780 378.900 93.780 379.900 ;
        RECT 93.930 378.900 95.530 379.900 ;
        RECT 95.680 378.900 96.680 379.900 ;
        RECT 96.830 378.900 97.830 379.900 ;
        RECT 4.830 372.400 5.530 373.100 ;
        RECT 4.830 371.550 5.530 372.250 ;
        RECT 4.830 370.700 5.530 371.400 ;
        RECT 23.930 372.400 24.630 373.100 ;
        RECT 24.830 372.400 25.530 373.100 ;
        RECT 23.930 371.550 24.630 372.250 ;
        RECT 24.830 371.550 25.530 372.250 ;
        RECT 23.930 370.700 24.630 371.400 ;
        RECT 24.830 370.700 25.530 371.400 ;
        RECT 4.830 368.600 5.530 369.300 ;
        RECT 4.830 367.750 5.530 368.450 ;
        RECT 4.830 366.900 5.530 367.600 ;
        RECT 43.930 372.400 44.630 373.100 ;
        RECT 44.830 372.400 45.530 373.100 ;
        RECT 43.930 371.550 44.630 372.250 ;
        RECT 44.830 371.550 45.530 372.250 ;
        RECT 43.930 370.700 44.630 371.400 ;
        RECT 44.830 370.700 45.530 371.400 ;
        RECT 23.930 368.600 24.630 369.300 ;
        RECT 24.830 368.600 25.530 369.300 ;
        RECT 23.930 367.750 24.630 368.450 ;
        RECT 24.830 367.750 25.530 368.450 ;
        RECT 23.930 366.900 24.630 367.600 ;
        RECT 24.830 366.900 25.530 367.600 ;
        RECT 63.930 372.400 64.630 373.100 ;
        RECT 64.830 372.400 65.530 373.100 ;
        RECT 63.930 371.550 64.630 372.250 ;
        RECT 64.830 371.550 65.530 372.250 ;
        RECT 63.930 370.700 64.630 371.400 ;
        RECT 64.830 370.700 65.530 371.400 ;
        RECT 43.930 368.600 44.630 369.300 ;
        RECT 44.830 368.600 45.530 369.300 ;
        RECT 43.930 367.750 44.630 368.450 ;
        RECT 44.830 367.750 45.530 368.450 ;
        RECT 43.930 366.900 44.630 367.600 ;
        RECT 44.830 366.900 45.530 367.600 ;
        RECT 83.930 372.400 84.630 373.100 ;
        RECT 84.830 372.400 85.530 373.100 ;
        RECT 83.930 371.550 84.630 372.250 ;
        RECT 84.830 371.550 85.530 372.250 ;
        RECT 83.930 370.700 84.630 371.400 ;
        RECT 84.830 370.700 85.530 371.400 ;
        RECT 63.930 368.600 64.630 369.300 ;
        RECT 64.830 368.600 65.530 369.300 ;
        RECT 63.930 367.750 64.630 368.450 ;
        RECT 64.830 367.750 65.530 368.450 ;
        RECT 63.930 366.900 64.630 367.600 ;
        RECT 64.830 366.900 65.530 367.600 ;
        RECT 103.930 372.400 104.630 373.100 ;
        RECT 103.930 371.550 104.630 372.250 ;
        RECT 103.930 370.700 104.630 371.400 ;
        RECT 83.930 368.600 84.630 369.300 ;
        RECT 84.830 368.600 85.530 369.300 ;
        RECT 83.930 367.750 84.630 368.450 ;
        RECT 84.830 367.750 85.530 368.450 ;
        RECT 83.930 366.900 84.630 367.600 ;
        RECT 84.830 366.900 85.530 367.600 ;
        RECT 110.050 369.975 110.410 370.355 ;
        RECT 110.680 369.975 111.040 370.355 ;
        RECT 111.280 369.975 111.640 370.355 ;
        RECT 110.050 369.385 110.410 369.765 ;
        RECT 110.680 369.385 111.040 369.765 ;
        RECT 111.280 369.385 111.640 369.765 ;
        RECT 103.930 368.600 104.630 369.300 ;
        RECT 103.930 367.750 104.630 368.450 ;
        RECT 103.930 366.900 104.630 367.600 ;
        RECT 11.630 360.100 12.630 361.100 ;
        RECT 12.730 360.100 13.730 361.100 ;
        RECT 13.880 360.100 15.480 361.100 ;
        RECT 15.680 360.100 16.680 361.100 ;
        RECT 16.830 360.100 17.830 361.100 ;
        RECT 11.630 358.900 12.630 359.900 ;
        RECT 12.780 358.900 13.780 359.900 ;
        RECT 13.930 358.900 15.530 359.900 ;
        RECT 15.680 358.900 16.680 359.900 ;
        RECT 16.830 358.900 17.830 359.900 ;
        RECT 31.630 360.100 32.630 361.100 ;
        RECT 32.730 360.100 33.730 361.100 ;
        RECT 33.880 360.100 35.480 361.100 ;
        RECT 35.680 360.100 36.680 361.100 ;
        RECT 36.830 360.100 37.830 361.100 ;
        RECT 31.630 358.900 32.630 359.900 ;
        RECT 32.780 358.900 33.780 359.900 ;
        RECT 33.930 358.900 35.530 359.900 ;
        RECT 35.680 358.900 36.680 359.900 ;
        RECT 36.830 358.900 37.830 359.900 ;
        RECT 51.630 360.100 52.630 361.100 ;
        RECT 52.730 360.100 53.730 361.100 ;
        RECT 53.880 360.100 55.480 361.100 ;
        RECT 55.680 360.100 56.680 361.100 ;
        RECT 56.830 360.100 57.830 361.100 ;
        RECT 51.630 358.900 52.630 359.900 ;
        RECT 52.780 358.900 53.780 359.900 ;
        RECT 53.930 358.900 55.530 359.900 ;
        RECT 55.680 358.900 56.680 359.900 ;
        RECT 56.830 358.900 57.830 359.900 ;
        RECT 71.630 360.100 72.630 361.100 ;
        RECT 72.730 360.100 73.730 361.100 ;
        RECT 73.880 360.100 75.480 361.100 ;
        RECT 75.680 360.100 76.680 361.100 ;
        RECT 76.830 360.100 77.830 361.100 ;
        RECT 71.630 358.900 72.630 359.900 ;
        RECT 72.780 358.900 73.780 359.900 ;
        RECT 73.930 358.900 75.530 359.900 ;
        RECT 75.680 358.900 76.680 359.900 ;
        RECT 76.830 358.900 77.830 359.900 ;
        RECT 91.630 360.100 92.630 361.100 ;
        RECT 92.730 360.100 93.730 361.100 ;
        RECT 93.880 360.100 95.480 361.100 ;
        RECT 95.680 360.100 96.680 361.100 ;
        RECT 96.830 360.100 97.830 361.100 ;
        RECT 91.630 358.900 92.630 359.900 ;
        RECT 92.780 358.900 93.780 359.900 ;
        RECT 93.930 358.900 95.530 359.900 ;
        RECT 95.680 358.900 96.680 359.900 ;
        RECT 96.830 358.900 97.830 359.900 ;
        RECT 4.830 352.400 5.530 353.100 ;
        RECT 4.830 351.550 5.530 352.250 ;
        RECT 4.830 350.700 5.530 351.400 ;
        RECT 23.930 352.400 24.630 353.100 ;
        RECT 24.830 352.400 25.530 353.100 ;
        RECT 23.930 351.550 24.630 352.250 ;
        RECT 24.830 351.550 25.530 352.250 ;
        RECT 23.930 350.700 24.630 351.400 ;
        RECT 24.830 350.700 25.530 351.400 ;
        RECT 4.830 348.600 5.530 349.300 ;
        RECT 4.830 347.750 5.530 348.450 ;
        RECT 4.830 346.900 5.530 347.600 ;
        RECT 43.930 352.400 44.630 353.100 ;
        RECT 44.830 352.400 45.530 353.100 ;
        RECT 43.930 351.550 44.630 352.250 ;
        RECT 44.830 351.550 45.530 352.250 ;
        RECT 43.930 350.700 44.630 351.400 ;
        RECT 44.830 350.700 45.530 351.400 ;
        RECT 23.930 348.600 24.630 349.300 ;
        RECT 24.830 348.600 25.530 349.300 ;
        RECT 23.930 347.750 24.630 348.450 ;
        RECT 24.830 347.750 25.530 348.450 ;
        RECT 23.930 346.900 24.630 347.600 ;
        RECT 24.830 346.900 25.530 347.600 ;
        RECT 63.930 352.400 64.630 353.100 ;
        RECT 64.830 352.400 65.530 353.100 ;
        RECT 63.930 351.550 64.630 352.250 ;
        RECT 64.830 351.550 65.530 352.250 ;
        RECT 63.930 350.700 64.630 351.400 ;
        RECT 64.830 350.700 65.530 351.400 ;
        RECT 43.930 348.600 44.630 349.300 ;
        RECT 44.830 348.600 45.530 349.300 ;
        RECT 43.930 347.750 44.630 348.450 ;
        RECT 44.830 347.750 45.530 348.450 ;
        RECT 43.930 346.900 44.630 347.600 ;
        RECT 44.830 346.900 45.530 347.600 ;
        RECT 83.930 352.400 84.630 353.100 ;
        RECT 84.830 352.400 85.530 353.100 ;
        RECT 83.930 351.550 84.630 352.250 ;
        RECT 84.830 351.550 85.530 352.250 ;
        RECT 83.930 350.700 84.630 351.400 ;
        RECT 84.830 350.700 85.530 351.400 ;
        RECT 63.930 348.600 64.630 349.300 ;
        RECT 64.830 348.600 65.530 349.300 ;
        RECT 63.930 347.750 64.630 348.450 ;
        RECT 64.830 347.750 65.530 348.450 ;
        RECT 63.930 346.900 64.630 347.600 ;
        RECT 64.830 346.900 65.530 347.600 ;
        RECT 103.930 352.400 104.630 353.100 ;
        RECT 103.930 351.550 104.630 352.250 ;
        RECT 103.930 350.700 104.630 351.400 ;
        RECT 83.930 348.600 84.630 349.300 ;
        RECT 84.830 348.600 85.530 349.300 ;
        RECT 83.930 347.750 84.630 348.450 ;
        RECT 84.830 347.750 85.530 348.450 ;
        RECT 83.930 346.900 84.630 347.600 ;
        RECT 84.830 346.900 85.530 347.600 ;
        RECT 110.050 349.975 110.410 350.355 ;
        RECT 110.680 349.975 111.040 350.355 ;
        RECT 111.280 349.975 111.640 350.355 ;
        RECT 110.050 349.385 110.410 349.765 ;
        RECT 110.680 349.385 111.040 349.765 ;
        RECT 111.280 349.385 111.640 349.765 ;
        RECT 103.930 348.600 104.630 349.300 ;
        RECT 103.930 347.750 104.630 348.450 ;
        RECT 103.930 346.900 104.630 347.600 ;
        RECT 11.630 340.100 12.630 341.100 ;
        RECT 12.730 340.100 13.730 341.100 ;
        RECT 13.880 340.100 15.480 341.100 ;
        RECT 15.680 340.100 16.680 341.100 ;
        RECT 16.830 340.100 17.830 341.100 ;
        RECT 11.630 338.900 12.630 339.900 ;
        RECT 12.780 338.900 13.780 339.900 ;
        RECT 13.930 338.900 15.530 339.900 ;
        RECT 15.680 338.900 16.680 339.900 ;
        RECT 16.830 338.900 17.830 339.900 ;
        RECT 31.630 340.100 32.630 341.100 ;
        RECT 32.730 340.100 33.730 341.100 ;
        RECT 33.880 340.100 35.480 341.100 ;
        RECT 35.680 340.100 36.680 341.100 ;
        RECT 36.830 340.100 37.830 341.100 ;
        RECT 31.630 338.900 32.630 339.900 ;
        RECT 32.780 338.900 33.780 339.900 ;
        RECT 33.930 338.900 35.530 339.900 ;
        RECT 35.680 338.900 36.680 339.900 ;
        RECT 36.830 338.900 37.830 339.900 ;
        RECT 51.630 340.100 52.630 341.100 ;
        RECT 52.730 340.100 53.730 341.100 ;
        RECT 53.880 340.100 55.480 341.100 ;
        RECT 55.680 340.100 56.680 341.100 ;
        RECT 56.830 340.100 57.830 341.100 ;
        RECT 51.630 338.900 52.630 339.900 ;
        RECT 52.780 338.900 53.780 339.900 ;
        RECT 53.930 338.900 55.530 339.900 ;
        RECT 55.680 338.900 56.680 339.900 ;
        RECT 56.830 338.900 57.830 339.900 ;
        RECT 71.630 340.100 72.630 341.100 ;
        RECT 72.730 340.100 73.730 341.100 ;
        RECT 73.880 340.100 75.480 341.100 ;
        RECT 75.680 340.100 76.680 341.100 ;
        RECT 76.830 340.100 77.830 341.100 ;
        RECT 71.630 338.900 72.630 339.900 ;
        RECT 72.780 338.900 73.780 339.900 ;
        RECT 73.930 338.900 75.530 339.900 ;
        RECT 75.680 338.900 76.680 339.900 ;
        RECT 76.830 338.900 77.830 339.900 ;
        RECT 91.630 340.100 92.630 341.100 ;
        RECT 92.730 340.100 93.730 341.100 ;
        RECT 93.880 340.100 95.480 341.100 ;
        RECT 95.680 340.100 96.680 341.100 ;
        RECT 96.830 340.100 97.830 341.100 ;
        RECT 91.630 338.900 92.630 339.900 ;
        RECT 92.780 338.900 93.780 339.900 ;
        RECT 93.930 338.900 95.530 339.900 ;
        RECT 95.680 338.900 96.680 339.900 ;
        RECT 96.830 338.900 97.830 339.900 ;
        RECT 4.830 332.400 5.530 333.100 ;
        RECT 4.830 331.550 5.530 332.250 ;
        RECT 4.830 330.700 5.530 331.400 ;
        RECT 23.930 332.400 24.630 333.100 ;
        RECT 24.830 332.400 25.530 333.100 ;
        RECT 23.930 331.550 24.630 332.250 ;
        RECT 24.830 331.550 25.530 332.250 ;
        RECT 23.930 330.700 24.630 331.400 ;
        RECT 24.830 330.700 25.530 331.400 ;
        RECT 4.830 328.600 5.530 329.300 ;
        RECT 4.830 327.750 5.530 328.450 ;
        RECT 4.830 326.900 5.530 327.600 ;
        RECT 43.930 332.400 44.630 333.100 ;
        RECT 44.830 332.400 45.530 333.100 ;
        RECT 43.930 331.550 44.630 332.250 ;
        RECT 44.830 331.550 45.530 332.250 ;
        RECT 43.930 330.700 44.630 331.400 ;
        RECT 44.830 330.700 45.530 331.400 ;
        RECT 23.930 328.600 24.630 329.300 ;
        RECT 24.830 328.600 25.530 329.300 ;
        RECT 23.930 327.750 24.630 328.450 ;
        RECT 24.830 327.750 25.530 328.450 ;
        RECT 23.930 326.900 24.630 327.600 ;
        RECT 24.830 326.900 25.530 327.600 ;
        RECT 63.930 332.400 64.630 333.100 ;
        RECT 64.830 332.400 65.530 333.100 ;
        RECT 63.930 331.550 64.630 332.250 ;
        RECT 64.830 331.550 65.530 332.250 ;
        RECT 63.930 330.700 64.630 331.400 ;
        RECT 64.830 330.700 65.530 331.400 ;
        RECT 43.930 328.600 44.630 329.300 ;
        RECT 44.830 328.600 45.530 329.300 ;
        RECT 43.930 327.750 44.630 328.450 ;
        RECT 44.830 327.750 45.530 328.450 ;
        RECT 43.930 326.900 44.630 327.600 ;
        RECT 44.830 326.900 45.530 327.600 ;
        RECT 83.930 332.400 84.630 333.100 ;
        RECT 84.830 332.400 85.530 333.100 ;
        RECT 83.930 331.550 84.630 332.250 ;
        RECT 84.830 331.550 85.530 332.250 ;
        RECT 83.930 330.700 84.630 331.400 ;
        RECT 84.830 330.700 85.530 331.400 ;
        RECT 63.930 328.600 64.630 329.300 ;
        RECT 64.830 328.600 65.530 329.300 ;
        RECT 63.930 327.750 64.630 328.450 ;
        RECT 64.830 327.750 65.530 328.450 ;
        RECT 63.930 326.900 64.630 327.600 ;
        RECT 64.830 326.900 65.530 327.600 ;
        RECT 103.930 332.400 104.630 333.100 ;
        RECT 103.930 331.550 104.630 332.250 ;
        RECT 103.930 330.700 104.630 331.400 ;
        RECT 83.930 328.600 84.630 329.300 ;
        RECT 84.830 328.600 85.530 329.300 ;
        RECT 83.930 327.750 84.630 328.450 ;
        RECT 84.830 327.750 85.530 328.450 ;
        RECT 83.930 326.900 84.630 327.600 ;
        RECT 84.830 326.900 85.530 327.600 ;
        RECT 110.050 329.910 110.410 330.290 ;
        RECT 110.680 329.910 111.040 330.290 ;
        RECT 111.280 329.910 111.640 330.290 ;
        RECT 110.050 329.320 110.410 329.700 ;
        RECT 110.680 329.320 111.040 329.700 ;
        RECT 111.280 329.320 111.640 329.700 ;
        RECT 103.930 328.600 104.630 329.300 ;
        RECT 103.930 327.750 104.630 328.450 ;
        RECT 103.930 326.900 104.630 327.600 ;
        RECT 11.630 320.100 12.630 321.100 ;
        RECT 12.730 320.100 13.730 321.100 ;
        RECT 13.880 320.100 15.480 321.100 ;
        RECT 15.680 320.100 16.680 321.100 ;
        RECT 16.830 320.100 17.830 321.100 ;
        RECT 11.630 318.900 12.630 319.900 ;
        RECT 12.780 318.900 13.780 319.900 ;
        RECT 13.930 318.900 15.530 319.900 ;
        RECT 15.680 318.900 16.680 319.900 ;
        RECT 16.830 318.900 17.830 319.900 ;
        RECT 31.630 320.100 32.630 321.100 ;
        RECT 32.730 320.100 33.730 321.100 ;
        RECT 33.880 320.100 35.480 321.100 ;
        RECT 35.680 320.100 36.680 321.100 ;
        RECT 36.830 320.100 37.830 321.100 ;
        RECT 31.630 318.900 32.630 319.900 ;
        RECT 32.780 318.900 33.780 319.900 ;
        RECT 33.930 318.900 35.530 319.900 ;
        RECT 35.680 318.900 36.680 319.900 ;
        RECT 36.830 318.900 37.830 319.900 ;
        RECT 51.630 320.100 52.630 321.100 ;
        RECT 52.730 320.100 53.730 321.100 ;
        RECT 53.880 320.100 55.480 321.100 ;
        RECT 55.680 320.100 56.680 321.100 ;
        RECT 56.830 320.100 57.830 321.100 ;
        RECT 51.630 318.900 52.630 319.900 ;
        RECT 52.780 318.900 53.780 319.900 ;
        RECT 53.930 318.900 55.530 319.900 ;
        RECT 55.680 318.900 56.680 319.900 ;
        RECT 56.830 318.900 57.830 319.900 ;
        RECT 71.630 320.100 72.630 321.100 ;
        RECT 72.730 320.100 73.730 321.100 ;
        RECT 73.880 320.100 75.480 321.100 ;
        RECT 75.680 320.100 76.680 321.100 ;
        RECT 76.830 320.100 77.830 321.100 ;
        RECT 71.630 318.900 72.630 319.900 ;
        RECT 72.780 318.900 73.780 319.900 ;
        RECT 73.930 318.900 75.530 319.900 ;
        RECT 75.680 318.900 76.680 319.900 ;
        RECT 76.830 318.900 77.830 319.900 ;
        RECT 91.630 320.100 92.630 321.100 ;
        RECT 92.730 320.100 93.730 321.100 ;
        RECT 93.880 320.100 95.480 321.100 ;
        RECT 95.680 320.100 96.680 321.100 ;
        RECT 96.830 320.100 97.830 321.100 ;
        RECT 91.630 318.900 92.630 319.900 ;
        RECT 92.780 318.900 93.780 319.900 ;
        RECT 93.930 318.900 95.530 319.900 ;
        RECT 95.680 318.900 96.680 319.900 ;
        RECT 96.830 318.900 97.830 319.900 ;
        RECT 4.830 312.400 5.530 313.100 ;
        RECT 4.830 311.550 5.530 312.250 ;
        RECT 4.830 310.700 5.530 311.400 ;
        RECT 23.930 312.400 24.630 313.100 ;
        RECT 24.830 312.400 25.530 313.100 ;
        RECT 23.930 311.550 24.630 312.250 ;
        RECT 24.830 311.550 25.530 312.250 ;
        RECT 23.930 310.700 24.630 311.400 ;
        RECT 24.830 310.700 25.530 311.400 ;
        RECT 4.830 308.600 5.530 309.300 ;
        RECT 4.830 307.750 5.530 308.450 ;
        RECT 4.830 306.900 5.530 307.600 ;
        RECT 43.930 312.400 44.630 313.100 ;
        RECT 44.830 312.400 45.530 313.100 ;
        RECT 43.930 311.550 44.630 312.250 ;
        RECT 44.830 311.550 45.530 312.250 ;
        RECT 43.930 310.700 44.630 311.400 ;
        RECT 44.830 310.700 45.530 311.400 ;
        RECT 23.930 308.600 24.630 309.300 ;
        RECT 24.830 308.600 25.530 309.300 ;
        RECT 23.930 307.750 24.630 308.450 ;
        RECT 24.830 307.750 25.530 308.450 ;
        RECT 23.930 306.900 24.630 307.600 ;
        RECT 24.830 306.900 25.530 307.600 ;
        RECT 63.930 312.400 64.630 313.100 ;
        RECT 64.830 312.400 65.530 313.100 ;
        RECT 63.930 311.550 64.630 312.250 ;
        RECT 64.830 311.550 65.530 312.250 ;
        RECT 63.930 310.700 64.630 311.400 ;
        RECT 64.830 310.700 65.530 311.400 ;
        RECT 43.930 308.600 44.630 309.300 ;
        RECT 44.830 308.600 45.530 309.300 ;
        RECT 43.930 307.750 44.630 308.450 ;
        RECT 44.830 307.750 45.530 308.450 ;
        RECT 43.930 306.900 44.630 307.600 ;
        RECT 44.830 306.900 45.530 307.600 ;
        RECT 83.930 312.400 84.630 313.100 ;
        RECT 84.830 312.400 85.530 313.100 ;
        RECT 83.930 311.550 84.630 312.250 ;
        RECT 84.830 311.550 85.530 312.250 ;
        RECT 83.930 310.700 84.630 311.400 ;
        RECT 84.830 310.700 85.530 311.400 ;
        RECT 63.930 308.600 64.630 309.300 ;
        RECT 64.830 308.600 65.530 309.300 ;
        RECT 63.930 307.750 64.630 308.450 ;
        RECT 64.830 307.750 65.530 308.450 ;
        RECT 63.930 306.900 64.630 307.600 ;
        RECT 64.830 306.900 65.530 307.600 ;
        RECT 103.930 312.400 104.630 313.100 ;
        RECT 103.930 311.550 104.630 312.250 ;
        RECT 103.930 310.700 104.630 311.400 ;
        RECT 83.930 308.600 84.630 309.300 ;
        RECT 84.830 308.600 85.530 309.300 ;
        RECT 83.930 307.750 84.630 308.450 ;
        RECT 84.830 307.750 85.530 308.450 ;
        RECT 83.930 306.900 84.630 307.600 ;
        RECT 84.830 306.900 85.530 307.600 ;
        RECT 110.050 309.905 110.410 310.285 ;
        RECT 110.680 309.905 111.040 310.285 ;
        RECT 111.280 309.905 111.640 310.285 ;
        RECT 110.050 309.315 110.410 309.695 ;
        RECT 110.680 309.315 111.040 309.695 ;
        RECT 111.280 309.315 111.640 309.695 ;
        RECT 103.930 308.600 104.630 309.300 ;
        RECT 103.930 307.750 104.630 308.450 ;
        RECT 103.930 306.900 104.630 307.600 ;
        RECT 11.630 300.100 12.630 301.100 ;
        RECT 12.730 300.100 13.730 301.100 ;
        RECT 13.880 300.100 15.480 301.100 ;
        RECT 15.680 300.100 16.680 301.100 ;
        RECT 16.830 300.100 17.830 301.100 ;
        RECT 11.630 298.900 12.630 299.900 ;
        RECT 12.780 298.900 13.780 299.900 ;
        RECT 13.930 298.900 15.530 299.900 ;
        RECT 15.680 298.900 16.680 299.900 ;
        RECT 16.830 298.900 17.830 299.900 ;
        RECT 31.630 300.100 32.630 301.100 ;
        RECT 32.730 300.100 33.730 301.100 ;
        RECT 33.880 300.100 35.480 301.100 ;
        RECT 35.680 300.100 36.680 301.100 ;
        RECT 36.830 300.100 37.830 301.100 ;
        RECT 31.630 298.900 32.630 299.900 ;
        RECT 32.780 298.900 33.780 299.900 ;
        RECT 33.930 298.900 35.530 299.900 ;
        RECT 35.680 298.900 36.680 299.900 ;
        RECT 36.830 298.900 37.830 299.900 ;
        RECT 51.630 300.100 52.630 301.100 ;
        RECT 52.730 300.100 53.730 301.100 ;
        RECT 53.880 300.100 55.480 301.100 ;
        RECT 55.680 300.100 56.680 301.100 ;
        RECT 56.830 300.100 57.830 301.100 ;
        RECT 51.630 298.900 52.630 299.900 ;
        RECT 52.780 298.900 53.780 299.900 ;
        RECT 53.930 298.900 55.530 299.900 ;
        RECT 55.680 298.900 56.680 299.900 ;
        RECT 56.830 298.900 57.830 299.900 ;
        RECT 71.630 300.100 72.630 301.100 ;
        RECT 72.730 300.100 73.730 301.100 ;
        RECT 73.880 300.100 75.480 301.100 ;
        RECT 75.680 300.100 76.680 301.100 ;
        RECT 76.830 300.100 77.830 301.100 ;
        RECT 71.630 298.900 72.630 299.900 ;
        RECT 72.780 298.900 73.780 299.900 ;
        RECT 73.930 298.900 75.530 299.900 ;
        RECT 75.680 298.900 76.680 299.900 ;
        RECT 76.830 298.900 77.830 299.900 ;
        RECT 91.630 300.100 92.630 301.100 ;
        RECT 92.730 300.100 93.730 301.100 ;
        RECT 93.880 300.100 95.480 301.100 ;
        RECT 95.680 300.100 96.680 301.100 ;
        RECT 96.830 300.100 97.830 301.100 ;
        RECT 91.630 298.900 92.630 299.900 ;
        RECT 92.780 298.900 93.780 299.900 ;
        RECT 93.930 298.900 95.530 299.900 ;
        RECT 95.680 298.900 96.680 299.900 ;
        RECT 96.830 298.900 97.830 299.900 ;
        RECT 4.830 292.400 5.530 293.100 ;
        RECT 4.830 291.550 5.530 292.250 ;
        RECT 4.830 290.700 5.530 291.400 ;
        RECT 23.930 292.400 24.630 293.100 ;
        RECT 24.830 292.400 25.530 293.100 ;
        RECT 23.930 291.550 24.630 292.250 ;
        RECT 24.830 291.550 25.530 292.250 ;
        RECT 23.930 290.700 24.630 291.400 ;
        RECT 24.830 290.700 25.530 291.400 ;
        RECT 4.830 288.600 5.530 289.300 ;
        RECT 4.830 287.750 5.530 288.450 ;
        RECT 4.830 286.900 5.530 287.600 ;
        RECT 43.930 292.400 44.630 293.100 ;
        RECT 44.830 292.400 45.530 293.100 ;
        RECT 43.930 291.550 44.630 292.250 ;
        RECT 44.830 291.550 45.530 292.250 ;
        RECT 43.930 290.700 44.630 291.400 ;
        RECT 44.830 290.700 45.530 291.400 ;
        RECT 23.930 288.600 24.630 289.300 ;
        RECT 24.830 288.600 25.530 289.300 ;
        RECT 23.930 287.750 24.630 288.450 ;
        RECT 24.830 287.750 25.530 288.450 ;
        RECT 23.930 286.900 24.630 287.600 ;
        RECT 24.830 286.900 25.530 287.600 ;
        RECT 63.930 292.400 64.630 293.100 ;
        RECT 64.830 292.400 65.530 293.100 ;
        RECT 63.930 291.550 64.630 292.250 ;
        RECT 64.830 291.550 65.530 292.250 ;
        RECT 63.930 290.700 64.630 291.400 ;
        RECT 64.830 290.700 65.530 291.400 ;
        RECT 43.930 288.600 44.630 289.300 ;
        RECT 44.830 288.600 45.530 289.300 ;
        RECT 43.930 287.750 44.630 288.450 ;
        RECT 44.830 287.750 45.530 288.450 ;
        RECT 43.930 286.900 44.630 287.600 ;
        RECT 44.830 286.900 45.530 287.600 ;
        RECT 83.930 292.400 84.630 293.100 ;
        RECT 84.830 292.400 85.530 293.100 ;
        RECT 83.930 291.550 84.630 292.250 ;
        RECT 84.830 291.550 85.530 292.250 ;
        RECT 83.930 290.700 84.630 291.400 ;
        RECT 84.830 290.700 85.530 291.400 ;
        RECT 63.930 288.600 64.630 289.300 ;
        RECT 64.830 288.600 65.530 289.300 ;
        RECT 63.930 287.750 64.630 288.450 ;
        RECT 64.830 287.750 65.530 288.450 ;
        RECT 63.930 286.900 64.630 287.600 ;
        RECT 64.830 286.900 65.530 287.600 ;
        RECT 103.930 292.400 104.630 293.100 ;
        RECT 103.930 291.550 104.630 292.250 ;
        RECT 103.930 290.700 104.630 291.400 ;
        RECT 83.930 288.600 84.630 289.300 ;
        RECT 84.830 288.600 85.530 289.300 ;
        RECT 83.930 287.750 84.630 288.450 ;
        RECT 84.830 287.750 85.530 288.450 ;
        RECT 83.930 286.900 84.630 287.600 ;
        RECT 84.830 286.900 85.530 287.600 ;
        RECT 110.050 290.100 110.410 290.480 ;
        RECT 110.680 290.100 111.040 290.480 ;
        RECT 111.280 290.100 111.640 290.480 ;
        RECT 110.050 289.510 110.410 289.890 ;
        RECT 110.680 289.510 111.040 289.890 ;
        RECT 111.280 289.510 111.640 289.890 ;
        RECT 103.930 288.600 104.630 289.300 ;
        RECT 103.930 287.750 104.630 288.450 ;
        RECT 103.930 286.900 104.630 287.600 ;
        RECT 11.630 280.100 12.630 281.100 ;
        RECT 12.730 280.100 13.730 281.100 ;
        RECT 13.880 280.100 15.480 281.100 ;
        RECT 15.680 280.100 16.680 281.100 ;
        RECT 16.830 280.100 17.830 281.100 ;
        RECT 11.630 278.900 12.630 279.900 ;
        RECT 12.780 278.900 13.780 279.900 ;
        RECT 13.930 278.900 15.530 279.900 ;
        RECT 15.680 278.900 16.680 279.900 ;
        RECT 16.830 278.900 17.830 279.900 ;
        RECT 31.630 280.100 32.630 281.100 ;
        RECT 32.730 280.100 33.730 281.100 ;
        RECT 33.880 280.100 35.480 281.100 ;
        RECT 35.680 280.100 36.680 281.100 ;
        RECT 36.830 280.100 37.830 281.100 ;
        RECT 31.630 278.900 32.630 279.900 ;
        RECT 32.780 278.900 33.780 279.900 ;
        RECT 33.930 278.900 35.530 279.900 ;
        RECT 35.680 278.900 36.680 279.900 ;
        RECT 36.830 278.900 37.830 279.900 ;
        RECT 51.630 280.100 52.630 281.100 ;
        RECT 52.730 280.100 53.730 281.100 ;
        RECT 53.880 280.100 55.480 281.100 ;
        RECT 55.680 280.100 56.680 281.100 ;
        RECT 56.830 280.100 57.830 281.100 ;
        RECT 51.630 278.900 52.630 279.900 ;
        RECT 52.780 278.900 53.780 279.900 ;
        RECT 53.930 278.900 55.530 279.900 ;
        RECT 55.680 278.900 56.680 279.900 ;
        RECT 56.830 278.900 57.830 279.900 ;
        RECT 71.630 280.100 72.630 281.100 ;
        RECT 72.730 280.100 73.730 281.100 ;
        RECT 73.880 280.100 75.480 281.100 ;
        RECT 75.680 280.100 76.680 281.100 ;
        RECT 76.830 280.100 77.830 281.100 ;
        RECT 71.630 278.900 72.630 279.900 ;
        RECT 72.780 278.900 73.780 279.900 ;
        RECT 73.930 278.900 75.530 279.900 ;
        RECT 75.680 278.900 76.680 279.900 ;
        RECT 76.830 278.900 77.830 279.900 ;
        RECT 91.630 280.100 92.630 281.100 ;
        RECT 92.730 280.100 93.730 281.100 ;
        RECT 93.880 280.100 95.480 281.100 ;
        RECT 95.680 280.100 96.680 281.100 ;
        RECT 96.830 280.100 97.830 281.100 ;
        RECT 91.630 278.900 92.630 279.900 ;
        RECT 92.780 278.900 93.780 279.900 ;
        RECT 93.930 278.900 95.530 279.900 ;
        RECT 95.680 278.900 96.680 279.900 ;
        RECT 96.830 278.900 97.830 279.900 ;
        RECT 4.830 272.400 5.530 273.100 ;
        RECT 4.830 271.550 5.530 272.250 ;
        RECT 4.830 270.700 5.530 271.400 ;
        RECT 23.930 272.400 24.630 273.100 ;
        RECT 24.830 272.400 25.530 273.100 ;
        RECT 23.930 271.550 24.630 272.250 ;
        RECT 24.830 271.550 25.530 272.250 ;
        RECT 23.930 270.700 24.630 271.400 ;
        RECT 24.830 270.700 25.530 271.400 ;
        RECT 4.830 268.600 5.530 269.300 ;
        RECT 4.830 267.750 5.530 268.450 ;
        RECT 4.830 266.900 5.530 267.600 ;
        RECT 43.930 272.400 44.630 273.100 ;
        RECT 44.830 272.400 45.530 273.100 ;
        RECT 43.930 271.550 44.630 272.250 ;
        RECT 44.830 271.550 45.530 272.250 ;
        RECT 43.930 270.700 44.630 271.400 ;
        RECT 44.830 270.700 45.530 271.400 ;
        RECT 23.930 268.600 24.630 269.300 ;
        RECT 24.830 268.600 25.530 269.300 ;
        RECT 23.930 267.750 24.630 268.450 ;
        RECT 24.830 267.750 25.530 268.450 ;
        RECT 23.930 266.900 24.630 267.600 ;
        RECT 24.830 266.900 25.530 267.600 ;
        RECT 63.930 272.400 64.630 273.100 ;
        RECT 64.830 272.400 65.530 273.100 ;
        RECT 63.930 271.550 64.630 272.250 ;
        RECT 64.830 271.550 65.530 272.250 ;
        RECT 63.930 270.700 64.630 271.400 ;
        RECT 64.830 270.700 65.530 271.400 ;
        RECT 43.930 268.600 44.630 269.300 ;
        RECT 44.830 268.600 45.530 269.300 ;
        RECT 43.930 267.750 44.630 268.450 ;
        RECT 44.830 267.750 45.530 268.450 ;
        RECT 43.930 266.900 44.630 267.600 ;
        RECT 44.830 266.900 45.530 267.600 ;
        RECT 83.930 272.400 84.630 273.100 ;
        RECT 84.830 272.400 85.530 273.100 ;
        RECT 83.930 271.550 84.630 272.250 ;
        RECT 84.830 271.550 85.530 272.250 ;
        RECT 83.930 270.700 84.630 271.400 ;
        RECT 84.830 270.700 85.530 271.400 ;
        RECT 63.930 268.600 64.630 269.300 ;
        RECT 64.830 268.600 65.530 269.300 ;
        RECT 63.930 267.750 64.630 268.450 ;
        RECT 64.830 267.750 65.530 268.450 ;
        RECT 63.930 266.900 64.630 267.600 ;
        RECT 64.830 266.900 65.530 267.600 ;
        RECT 103.930 272.400 104.630 273.100 ;
        RECT 103.930 271.550 104.630 272.250 ;
        RECT 103.930 270.700 104.630 271.400 ;
        RECT 83.930 268.600 84.630 269.300 ;
        RECT 84.830 268.600 85.530 269.300 ;
        RECT 83.930 267.750 84.630 268.450 ;
        RECT 84.830 267.750 85.530 268.450 ;
        RECT 83.930 266.900 84.630 267.600 ;
        RECT 84.830 266.900 85.530 267.600 ;
        RECT 110.050 270.015 110.410 270.395 ;
        RECT 110.680 270.015 111.040 270.395 ;
        RECT 111.280 270.015 111.640 270.395 ;
        RECT 110.050 269.425 110.410 269.805 ;
        RECT 110.680 269.425 111.040 269.805 ;
        RECT 111.280 269.425 111.640 269.805 ;
        RECT 103.930 268.600 104.630 269.300 ;
        RECT 103.930 267.750 104.630 268.450 ;
        RECT 103.930 266.900 104.630 267.600 ;
        RECT 11.630 260.100 12.630 261.100 ;
        RECT 12.730 260.100 13.730 261.100 ;
        RECT 13.880 260.100 15.480 261.100 ;
        RECT 15.680 260.100 16.680 261.100 ;
        RECT 16.830 260.100 17.830 261.100 ;
        RECT 11.630 258.900 12.630 259.900 ;
        RECT 12.780 258.900 13.780 259.900 ;
        RECT 13.930 258.900 15.530 259.900 ;
        RECT 15.680 258.900 16.680 259.900 ;
        RECT 16.830 258.900 17.830 259.900 ;
        RECT 31.630 260.100 32.630 261.100 ;
        RECT 32.730 260.100 33.730 261.100 ;
        RECT 33.880 260.100 35.480 261.100 ;
        RECT 35.680 260.100 36.680 261.100 ;
        RECT 36.830 260.100 37.830 261.100 ;
        RECT 31.630 258.900 32.630 259.900 ;
        RECT 32.780 258.900 33.780 259.900 ;
        RECT 33.930 258.900 35.530 259.900 ;
        RECT 35.680 258.900 36.680 259.900 ;
        RECT 36.830 258.900 37.830 259.900 ;
        RECT 51.630 260.100 52.630 261.100 ;
        RECT 52.730 260.100 53.730 261.100 ;
        RECT 53.880 260.100 55.480 261.100 ;
        RECT 55.680 260.100 56.680 261.100 ;
        RECT 56.830 260.100 57.830 261.100 ;
        RECT 51.630 258.900 52.630 259.900 ;
        RECT 52.780 258.900 53.780 259.900 ;
        RECT 53.930 258.900 55.530 259.900 ;
        RECT 55.680 258.900 56.680 259.900 ;
        RECT 56.830 258.900 57.830 259.900 ;
        RECT 71.630 260.100 72.630 261.100 ;
        RECT 72.730 260.100 73.730 261.100 ;
        RECT 73.880 260.100 75.480 261.100 ;
        RECT 75.680 260.100 76.680 261.100 ;
        RECT 76.830 260.100 77.830 261.100 ;
        RECT 71.630 258.900 72.630 259.900 ;
        RECT 72.780 258.900 73.780 259.900 ;
        RECT 73.930 258.900 75.530 259.900 ;
        RECT 75.680 258.900 76.680 259.900 ;
        RECT 76.830 258.900 77.830 259.900 ;
        RECT 91.630 260.100 92.630 261.100 ;
        RECT 92.730 260.100 93.730 261.100 ;
        RECT 93.880 260.100 95.480 261.100 ;
        RECT 95.680 260.100 96.680 261.100 ;
        RECT 96.830 260.100 97.830 261.100 ;
        RECT 91.630 258.900 92.630 259.900 ;
        RECT 92.780 258.900 93.780 259.900 ;
        RECT 93.930 258.900 95.530 259.900 ;
        RECT 95.680 258.900 96.680 259.900 ;
        RECT 96.830 258.900 97.830 259.900 ;
        RECT 4.830 252.400 5.530 253.100 ;
        RECT 4.830 251.550 5.530 252.250 ;
        RECT 4.830 250.700 5.530 251.400 ;
        RECT 23.930 252.400 24.630 253.100 ;
        RECT 24.830 252.400 25.530 253.100 ;
        RECT 23.930 251.550 24.630 252.250 ;
        RECT 24.830 251.550 25.530 252.250 ;
        RECT 23.930 250.700 24.630 251.400 ;
        RECT 24.830 250.700 25.530 251.400 ;
        RECT 4.830 248.600 5.530 249.300 ;
        RECT 4.830 247.750 5.530 248.450 ;
        RECT 4.830 246.900 5.530 247.600 ;
        RECT 43.930 252.400 44.630 253.100 ;
        RECT 44.830 252.400 45.530 253.100 ;
        RECT 43.930 251.550 44.630 252.250 ;
        RECT 44.830 251.550 45.530 252.250 ;
        RECT 43.930 250.700 44.630 251.400 ;
        RECT 44.830 250.700 45.530 251.400 ;
        RECT 23.930 248.600 24.630 249.300 ;
        RECT 24.830 248.600 25.530 249.300 ;
        RECT 23.930 247.750 24.630 248.450 ;
        RECT 24.830 247.750 25.530 248.450 ;
        RECT 23.930 246.900 24.630 247.600 ;
        RECT 24.830 246.900 25.530 247.600 ;
        RECT 63.930 252.400 64.630 253.100 ;
        RECT 64.830 252.400 65.530 253.100 ;
        RECT 63.930 251.550 64.630 252.250 ;
        RECT 64.830 251.550 65.530 252.250 ;
        RECT 63.930 250.700 64.630 251.400 ;
        RECT 64.830 250.700 65.530 251.400 ;
        RECT 43.930 248.600 44.630 249.300 ;
        RECT 44.830 248.600 45.530 249.300 ;
        RECT 43.930 247.750 44.630 248.450 ;
        RECT 44.830 247.750 45.530 248.450 ;
        RECT 43.930 246.900 44.630 247.600 ;
        RECT 44.830 246.900 45.530 247.600 ;
        RECT 83.930 252.400 84.630 253.100 ;
        RECT 84.830 252.400 85.530 253.100 ;
        RECT 83.930 251.550 84.630 252.250 ;
        RECT 84.830 251.550 85.530 252.250 ;
        RECT 83.930 250.700 84.630 251.400 ;
        RECT 84.830 250.700 85.530 251.400 ;
        RECT 63.930 248.600 64.630 249.300 ;
        RECT 64.830 248.600 65.530 249.300 ;
        RECT 63.930 247.750 64.630 248.450 ;
        RECT 64.830 247.750 65.530 248.450 ;
        RECT 63.930 246.900 64.630 247.600 ;
        RECT 64.830 246.900 65.530 247.600 ;
        RECT 103.930 252.400 104.630 253.100 ;
        RECT 103.930 251.550 104.630 252.250 ;
        RECT 103.930 250.700 104.630 251.400 ;
        RECT 83.930 248.600 84.630 249.300 ;
        RECT 84.830 248.600 85.530 249.300 ;
        RECT 83.930 247.750 84.630 248.450 ;
        RECT 84.830 247.750 85.530 248.450 ;
        RECT 83.930 246.900 84.630 247.600 ;
        RECT 84.830 246.900 85.530 247.600 ;
        RECT 110.050 250.410 110.410 250.790 ;
        RECT 110.680 250.410 111.040 250.790 ;
        RECT 111.280 250.410 111.640 250.790 ;
        RECT 110.050 249.820 110.410 250.200 ;
        RECT 110.680 249.820 111.040 250.200 ;
        RECT 111.280 249.820 111.640 250.200 ;
        RECT 103.930 248.600 104.630 249.300 ;
        RECT 103.930 247.750 104.630 248.450 ;
        RECT 103.930 246.900 104.630 247.600 ;
        RECT 11.630 240.100 12.630 241.100 ;
        RECT 12.730 240.100 13.730 241.100 ;
        RECT 13.880 240.100 15.480 241.100 ;
        RECT 15.680 240.100 16.680 241.100 ;
        RECT 16.830 240.100 17.830 241.100 ;
        RECT 11.630 238.900 12.630 239.900 ;
        RECT 12.780 238.900 13.780 239.900 ;
        RECT 13.930 238.900 15.530 239.900 ;
        RECT 15.680 238.900 16.680 239.900 ;
        RECT 16.830 238.900 17.830 239.900 ;
        RECT 31.630 240.100 32.630 241.100 ;
        RECT 32.730 240.100 33.730 241.100 ;
        RECT 33.880 240.100 35.480 241.100 ;
        RECT 35.680 240.100 36.680 241.100 ;
        RECT 36.830 240.100 37.830 241.100 ;
        RECT 31.630 238.900 32.630 239.900 ;
        RECT 32.780 238.900 33.780 239.900 ;
        RECT 33.930 238.900 35.530 239.900 ;
        RECT 35.680 238.900 36.680 239.900 ;
        RECT 36.830 238.900 37.830 239.900 ;
        RECT 51.630 240.100 52.630 241.100 ;
        RECT 52.730 240.100 53.730 241.100 ;
        RECT 53.880 240.100 55.480 241.100 ;
        RECT 55.680 240.100 56.680 241.100 ;
        RECT 56.830 240.100 57.830 241.100 ;
        RECT 51.630 238.900 52.630 239.900 ;
        RECT 52.780 238.900 53.780 239.900 ;
        RECT 53.930 238.900 55.530 239.900 ;
        RECT 55.680 238.900 56.680 239.900 ;
        RECT 56.830 238.900 57.830 239.900 ;
        RECT 71.630 240.100 72.630 241.100 ;
        RECT 72.730 240.100 73.730 241.100 ;
        RECT 73.880 240.100 75.480 241.100 ;
        RECT 75.680 240.100 76.680 241.100 ;
        RECT 76.830 240.100 77.830 241.100 ;
        RECT 71.630 238.900 72.630 239.900 ;
        RECT 72.780 238.900 73.780 239.900 ;
        RECT 73.930 238.900 75.530 239.900 ;
        RECT 75.680 238.900 76.680 239.900 ;
        RECT 76.830 238.900 77.830 239.900 ;
        RECT 91.630 240.100 92.630 241.100 ;
        RECT 92.730 240.100 93.730 241.100 ;
        RECT 93.880 240.100 95.480 241.100 ;
        RECT 95.680 240.100 96.680 241.100 ;
        RECT 96.830 240.100 97.830 241.100 ;
        RECT 91.630 238.900 92.630 239.900 ;
        RECT 92.780 238.900 93.780 239.900 ;
        RECT 93.930 238.900 95.530 239.900 ;
        RECT 95.680 238.900 96.680 239.900 ;
        RECT 96.830 238.900 97.830 239.900 ;
        RECT 4.830 232.400 5.530 233.100 ;
        RECT 4.830 231.550 5.530 232.250 ;
        RECT 4.830 230.700 5.530 231.400 ;
        RECT 23.930 232.400 24.630 233.100 ;
        RECT 24.830 232.400 25.530 233.100 ;
        RECT 23.930 231.550 24.630 232.250 ;
        RECT 24.830 231.550 25.530 232.250 ;
        RECT 23.930 230.700 24.630 231.400 ;
        RECT 24.830 230.700 25.530 231.400 ;
        RECT 4.830 228.600 5.530 229.300 ;
        RECT 4.830 227.750 5.530 228.450 ;
        RECT 4.830 226.900 5.530 227.600 ;
        RECT 43.930 232.400 44.630 233.100 ;
        RECT 44.830 232.400 45.530 233.100 ;
        RECT 43.930 231.550 44.630 232.250 ;
        RECT 44.830 231.550 45.530 232.250 ;
        RECT 43.930 230.700 44.630 231.400 ;
        RECT 44.830 230.700 45.530 231.400 ;
        RECT 23.930 228.600 24.630 229.300 ;
        RECT 24.830 228.600 25.530 229.300 ;
        RECT 23.930 227.750 24.630 228.450 ;
        RECT 24.830 227.750 25.530 228.450 ;
        RECT 23.930 226.900 24.630 227.600 ;
        RECT 24.830 226.900 25.530 227.600 ;
        RECT 63.930 232.400 64.630 233.100 ;
        RECT 64.830 232.400 65.530 233.100 ;
        RECT 63.930 231.550 64.630 232.250 ;
        RECT 64.830 231.550 65.530 232.250 ;
        RECT 63.930 230.700 64.630 231.400 ;
        RECT 64.830 230.700 65.530 231.400 ;
        RECT 43.930 228.600 44.630 229.300 ;
        RECT 44.830 228.600 45.530 229.300 ;
        RECT 43.930 227.750 44.630 228.450 ;
        RECT 44.830 227.750 45.530 228.450 ;
        RECT 43.930 226.900 44.630 227.600 ;
        RECT 44.830 226.900 45.530 227.600 ;
        RECT 83.930 232.400 84.630 233.100 ;
        RECT 84.830 232.400 85.530 233.100 ;
        RECT 83.930 231.550 84.630 232.250 ;
        RECT 84.830 231.550 85.530 232.250 ;
        RECT 83.930 230.700 84.630 231.400 ;
        RECT 84.830 230.700 85.530 231.400 ;
        RECT 63.930 228.600 64.630 229.300 ;
        RECT 64.830 228.600 65.530 229.300 ;
        RECT 63.930 227.750 64.630 228.450 ;
        RECT 64.830 227.750 65.530 228.450 ;
        RECT 63.930 226.900 64.630 227.600 ;
        RECT 64.830 226.900 65.530 227.600 ;
        RECT 103.930 232.400 104.630 233.100 ;
        RECT 103.930 231.550 104.630 232.250 ;
        RECT 103.930 230.700 104.630 231.400 ;
        RECT 83.930 228.600 84.630 229.300 ;
        RECT 84.830 228.600 85.530 229.300 ;
        RECT 83.930 227.750 84.630 228.450 ;
        RECT 84.830 227.750 85.530 228.450 ;
        RECT 83.930 226.900 84.630 227.600 ;
        RECT 84.830 226.900 85.530 227.600 ;
        RECT 103.930 228.600 104.630 229.300 ;
        RECT 110.050 229.120 110.410 229.500 ;
        RECT 110.680 229.120 111.040 229.500 ;
        RECT 111.280 229.120 111.640 229.500 ;
        RECT 110.050 228.530 110.410 228.910 ;
        RECT 110.680 228.530 111.040 228.910 ;
        RECT 111.280 228.530 111.640 228.910 ;
        RECT 103.930 227.750 104.630 228.450 ;
        RECT 103.930 226.900 104.630 227.600 ;
        RECT 11.630 220.100 12.630 221.100 ;
        RECT 12.730 220.100 13.730 221.100 ;
        RECT 13.880 220.100 15.480 221.100 ;
        RECT 15.680 220.100 16.680 221.100 ;
        RECT 16.830 220.100 17.830 221.100 ;
        RECT 31.630 220.100 32.630 221.100 ;
        RECT 32.730 220.100 33.730 221.100 ;
        RECT 33.880 220.100 35.480 221.100 ;
        RECT 35.680 220.100 36.680 221.100 ;
        RECT 36.830 220.100 37.830 221.100 ;
        RECT 51.630 220.100 52.630 221.100 ;
        RECT 52.730 220.100 53.730 221.100 ;
        RECT 53.880 220.100 55.480 221.100 ;
        RECT 55.680 220.100 56.680 221.100 ;
        RECT 56.830 220.100 57.830 221.100 ;
        RECT 71.630 220.100 72.630 221.100 ;
        RECT 72.730 220.100 73.730 221.100 ;
        RECT 73.880 220.100 75.480 221.100 ;
        RECT 75.680 220.100 76.680 221.100 ;
        RECT 76.830 220.100 77.830 221.100 ;
        RECT 91.630 220.100 92.630 221.100 ;
        RECT 92.730 220.100 93.730 221.100 ;
        RECT 93.880 220.100 95.480 221.100 ;
        RECT 95.680 220.100 96.680 221.100 ;
        RECT 96.830 220.100 97.830 221.100 ;
        RECT 9.425 196.405 10.015 196.975 ;
        RECT 10.205 196.405 10.795 196.975 ;
        RECT 10.985 196.405 11.575 196.975 ;
        RECT 11.630 158.900 12.630 159.900 ;
        RECT 12.780 158.900 13.780 159.900 ;
        RECT 13.930 158.900 15.530 159.900 ;
        RECT 15.680 158.900 16.680 159.900 ;
        RECT 16.830 158.900 17.830 159.900 ;
        RECT 31.630 158.900 32.630 159.900 ;
        RECT 32.780 158.900 33.780 159.900 ;
        RECT 33.930 158.900 35.530 159.900 ;
        RECT 35.680 158.900 36.680 159.900 ;
        RECT 36.830 158.900 37.830 159.900 ;
        RECT 51.630 158.900 52.630 159.900 ;
        RECT 52.780 158.900 53.780 159.900 ;
        RECT 53.930 158.900 55.530 159.900 ;
        RECT 55.680 158.900 56.680 159.900 ;
        RECT 56.830 158.900 57.830 159.900 ;
        RECT 71.630 158.900 72.630 159.900 ;
        RECT 72.780 158.900 73.780 159.900 ;
        RECT 73.930 158.900 75.530 159.900 ;
        RECT 75.680 158.900 76.680 159.900 ;
        RECT 76.830 158.900 77.830 159.900 ;
        RECT 91.630 158.900 92.630 159.900 ;
        RECT 92.780 158.900 93.780 159.900 ;
        RECT 93.930 158.900 95.530 159.900 ;
        RECT 95.680 158.900 96.680 159.900 ;
        RECT 96.830 158.900 97.830 159.900 ;
        RECT 4.830 152.400 5.530 153.100 ;
        RECT 4.830 151.550 5.530 152.250 ;
        RECT 4.830 150.700 5.530 151.400 ;
        RECT 23.930 152.400 24.630 153.100 ;
        RECT 24.830 152.400 25.530 153.100 ;
        RECT 23.930 151.550 24.630 152.250 ;
        RECT 24.830 151.550 25.530 152.250 ;
        RECT 23.930 150.700 24.630 151.400 ;
        RECT 24.830 150.700 25.530 151.400 ;
        RECT 4.830 148.600 5.530 149.300 ;
        RECT 4.830 147.750 5.530 148.450 ;
        RECT 4.830 146.900 5.530 147.600 ;
        RECT 43.930 152.400 44.630 153.100 ;
        RECT 44.830 152.400 45.530 153.100 ;
        RECT 43.930 151.550 44.630 152.250 ;
        RECT 44.830 151.550 45.530 152.250 ;
        RECT 43.930 150.700 44.630 151.400 ;
        RECT 44.830 150.700 45.530 151.400 ;
        RECT 23.930 148.600 24.630 149.300 ;
        RECT 24.830 148.600 25.530 149.300 ;
        RECT 23.930 147.750 24.630 148.450 ;
        RECT 24.830 147.750 25.530 148.450 ;
        RECT 23.930 146.900 24.630 147.600 ;
        RECT 24.830 146.900 25.530 147.600 ;
        RECT 63.930 152.400 64.630 153.100 ;
        RECT 64.830 152.400 65.530 153.100 ;
        RECT 63.930 151.550 64.630 152.250 ;
        RECT 64.830 151.550 65.530 152.250 ;
        RECT 63.930 150.700 64.630 151.400 ;
        RECT 64.830 150.700 65.530 151.400 ;
        RECT 43.930 148.600 44.630 149.300 ;
        RECT 44.830 148.600 45.530 149.300 ;
        RECT 43.930 147.750 44.630 148.450 ;
        RECT 44.830 147.750 45.530 148.450 ;
        RECT 43.930 146.900 44.630 147.600 ;
        RECT 44.830 146.900 45.530 147.600 ;
        RECT 83.930 152.400 84.630 153.100 ;
        RECT 84.830 152.400 85.530 153.100 ;
        RECT 83.930 151.550 84.630 152.250 ;
        RECT 84.830 151.550 85.530 152.250 ;
        RECT 83.930 150.700 84.630 151.400 ;
        RECT 84.830 150.700 85.530 151.400 ;
        RECT 63.930 148.600 64.630 149.300 ;
        RECT 64.830 148.600 65.530 149.300 ;
        RECT 63.930 147.750 64.630 148.450 ;
        RECT 64.830 147.750 65.530 148.450 ;
        RECT 63.930 146.900 64.630 147.600 ;
        RECT 64.830 146.900 65.530 147.600 ;
        RECT 103.930 152.400 104.630 153.100 ;
        RECT 103.930 151.550 104.630 152.250 ;
        RECT 103.930 150.700 104.630 151.400 ;
        RECT 83.930 148.600 84.630 149.300 ;
        RECT 84.830 148.600 85.530 149.300 ;
        RECT 83.930 147.750 84.630 148.450 ;
        RECT 84.830 147.750 85.530 148.450 ;
        RECT 83.930 146.900 84.630 147.600 ;
        RECT 84.830 146.900 85.530 147.600 ;
        RECT 110.050 150.270 110.410 150.650 ;
        RECT 110.680 150.270 111.040 150.650 ;
        RECT 111.280 150.270 111.640 150.650 ;
        RECT 110.050 149.680 110.410 150.060 ;
        RECT 110.680 149.680 111.040 150.060 ;
        RECT 111.280 149.680 111.640 150.060 ;
        RECT 103.930 148.600 104.630 149.300 ;
        RECT 103.930 147.750 104.630 148.450 ;
        RECT 103.930 146.900 104.630 147.600 ;
        RECT 11.630 140.100 12.630 141.100 ;
        RECT 12.730 140.100 13.730 141.100 ;
        RECT 13.880 140.100 15.480 141.100 ;
        RECT 15.680 140.100 16.680 141.100 ;
        RECT 16.830 140.100 17.830 141.100 ;
        RECT 11.630 138.900 12.630 139.900 ;
        RECT 12.780 138.900 13.780 139.900 ;
        RECT 13.930 138.900 15.530 139.900 ;
        RECT 15.680 138.900 16.680 139.900 ;
        RECT 16.830 138.900 17.830 139.900 ;
        RECT 31.630 140.100 32.630 141.100 ;
        RECT 32.730 140.100 33.730 141.100 ;
        RECT 33.880 140.100 35.480 141.100 ;
        RECT 35.680 140.100 36.680 141.100 ;
        RECT 36.830 140.100 37.830 141.100 ;
        RECT 31.630 138.900 32.630 139.900 ;
        RECT 32.780 138.900 33.780 139.900 ;
        RECT 33.930 138.900 35.530 139.900 ;
        RECT 35.680 138.900 36.680 139.900 ;
        RECT 36.830 138.900 37.830 139.900 ;
        RECT 51.630 140.100 52.630 141.100 ;
        RECT 52.730 140.100 53.730 141.100 ;
        RECT 53.880 140.100 55.480 141.100 ;
        RECT 55.680 140.100 56.680 141.100 ;
        RECT 56.830 140.100 57.830 141.100 ;
        RECT 51.630 138.900 52.630 139.900 ;
        RECT 52.780 138.900 53.780 139.900 ;
        RECT 53.930 138.900 55.530 139.900 ;
        RECT 55.680 138.900 56.680 139.900 ;
        RECT 56.830 138.900 57.830 139.900 ;
        RECT 71.630 140.100 72.630 141.100 ;
        RECT 72.730 140.100 73.730 141.100 ;
        RECT 73.880 140.100 75.480 141.100 ;
        RECT 75.680 140.100 76.680 141.100 ;
        RECT 76.830 140.100 77.830 141.100 ;
        RECT 71.630 138.900 72.630 139.900 ;
        RECT 72.780 138.900 73.780 139.900 ;
        RECT 73.930 138.900 75.530 139.900 ;
        RECT 75.680 138.900 76.680 139.900 ;
        RECT 76.830 138.900 77.830 139.900 ;
        RECT 91.630 140.100 92.630 141.100 ;
        RECT 92.730 140.100 93.730 141.100 ;
        RECT 93.880 140.100 95.480 141.100 ;
        RECT 95.680 140.100 96.680 141.100 ;
        RECT 96.830 140.100 97.830 141.100 ;
        RECT 91.630 138.900 92.630 139.900 ;
        RECT 92.780 138.900 93.780 139.900 ;
        RECT 93.930 138.900 95.530 139.900 ;
        RECT 95.680 138.900 96.680 139.900 ;
        RECT 96.830 138.900 97.830 139.900 ;
        RECT 4.830 132.400 5.530 133.100 ;
        RECT 4.830 131.550 5.530 132.250 ;
        RECT 4.830 130.700 5.530 131.400 ;
        RECT 23.930 132.400 24.630 133.100 ;
        RECT 24.830 132.400 25.530 133.100 ;
        RECT 23.930 131.550 24.630 132.250 ;
        RECT 24.830 131.550 25.530 132.250 ;
        RECT 23.930 130.700 24.630 131.400 ;
        RECT 24.830 130.700 25.530 131.400 ;
        RECT 4.830 128.600 5.530 129.300 ;
        RECT 4.830 127.750 5.530 128.450 ;
        RECT 4.830 126.900 5.530 127.600 ;
        RECT 43.930 132.400 44.630 133.100 ;
        RECT 44.830 132.400 45.530 133.100 ;
        RECT 43.930 131.550 44.630 132.250 ;
        RECT 44.830 131.550 45.530 132.250 ;
        RECT 43.930 130.700 44.630 131.400 ;
        RECT 44.830 130.700 45.530 131.400 ;
        RECT 23.930 128.600 24.630 129.300 ;
        RECT 24.830 128.600 25.530 129.300 ;
        RECT 23.930 127.750 24.630 128.450 ;
        RECT 24.830 127.750 25.530 128.450 ;
        RECT 23.930 126.900 24.630 127.600 ;
        RECT 24.830 126.900 25.530 127.600 ;
        RECT 63.930 132.400 64.630 133.100 ;
        RECT 64.830 132.400 65.530 133.100 ;
        RECT 63.930 131.550 64.630 132.250 ;
        RECT 64.830 131.550 65.530 132.250 ;
        RECT 63.930 130.700 64.630 131.400 ;
        RECT 64.830 130.700 65.530 131.400 ;
        RECT 43.930 128.600 44.630 129.300 ;
        RECT 44.830 128.600 45.530 129.300 ;
        RECT 43.930 127.750 44.630 128.450 ;
        RECT 44.830 127.750 45.530 128.450 ;
        RECT 43.930 126.900 44.630 127.600 ;
        RECT 44.830 126.900 45.530 127.600 ;
        RECT 83.930 132.400 84.630 133.100 ;
        RECT 84.830 132.400 85.530 133.100 ;
        RECT 83.930 131.550 84.630 132.250 ;
        RECT 84.830 131.550 85.530 132.250 ;
        RECT 83.930 130.700 84.630 131.400 ;
        RECT 84.830 130.700 85.530 131.400 ;
        RECT 63.930 128.600 64.630 129.300 ;
        RECT 64.830 128.600 65.530 129.300 ;
        RECT 63.930 127.750 64.630 128.450 ;
        RECT 64.830 127.750 65.530 128.450 ;
        RECT 63.930 126.900 64.630 127.600 ;
        RECT 64.830 126.900 65.530 127.600 ;
        RECT 103.930 132.400 104.630 133.100 ;
        RECT 103.930 131.550 104.630 132.250 ;
        RECT 103.930 130.700 104.630 131.400 ;
        RECT 83.930 128.600 84.630 129.300 ;
        RECT 84.830 128.600 85.530 129.300 ;
        RECT 83.930 127.750 84.630 128.450 ;
        RECT 84.830 127.750 85.530 128.450 ;
        RECT 83.930 126.900 84.630 127.600 ;
        RECT 84.830 126.900 85.530 127.600 ;
        RECT 110.050 129.475 110.410 129.855 ;
        RECT 110.680 129.475 111.040 129.855 ;
        RECT 111.280 129.475 111.640 129.855 ;
        RECT 103.930 128.600 104.630 129.300 ;
        RECT 110.050 128.885 110.410 129.265 ;
        RECT 110.680 128.885 111.040 129.265 ;
        RECT 111.280 128.885 111.640 129.265 ;
        RECT 103.930 127.750 104.630 128.450 ;
        RECT 103.930 126.900 104.630 127.600 ;
        RECT 11.630 120.100 12.630 121.100 ;
        RECT 12.730 120.100 13.730 121.100 ;
        RECT 13.880 120.100 15.480 121.100 ;
        RECT 15.680 120.100 16.680 121.100 ;
        RECT 16.830 120.100 17.830 121.100 ;
        RECT 11.630 118.900 12.630 119.900 ;
        RECT 12.780 118.900 13.780 119.900 ;
        RECT 13.930 118.900 15.530 119.900 ;
        RECT 15.680 118.900 16.680 119.900 ;
        RECT 16.830 118.900 17.830 119.900 ;
        RECT 31.630 120.100 32.630 121.100 ;
        RECT 32.730 120.100 33.730 121.100 ;
        RECT 33.880 120.100 35.480 121.100 ;
        RECT 35.680 120.100 36.680 121.100 ;
        RECT 36.830 120.100 37.830 121.100 ;
        RECT 31.630 118.900 32.630 119.900 ;
        RECT 32.780 118.900 33.780 119.900 ;
        RECT 33.930 118.900 35.530 119.900 ;
        RECT 35.680 118.900 36.680 119.900 ;
        RECT 36.830 118.900 37.830 119.900 ;
        RECT 51.630 120.100 52.630 121.100 ;
        RECT 52.730 120.100 53.730 121.100 ;
        RECT 53.880 120.100 55.480 121.100 ;
        RECT 55.680 120.100 56.680 121.100 ;
        RECT 56.830 120.100 57.830 121.100 ;
        RECT 51.630 118.900 52.630 119.900 ;
        RECT 52.780 118.900 53.780 119.900 ;
        RECT 53.930 118.900 55.530 119.900 ;
        RECT 55.680 118.900 56.680 119.900 ;
        RECT 56.830 118.900 57.830 119.900 ;
        RECT 71.630 120.100 72.630 121.100 ;
        RECT 72.730 120.100 73.730 121.100 ;
        RECT 73.880 120.100 75.480 121.100 ;
        RECT 75.680 120.100 76.680 121.100 ;
        RECT 76.830 120.100 77.830 121.100 ;
        RECT 71.630 118.900 72.630 119.900 ;
        RECT 72.780 118.900 73.780 119.900 ;
        RECT 73.930 118.900 75.530 119.900 ;
        RECT 75.680 118.900 76.680 119.900 ;
        RECT 76.830 118.900 77.830 119.900 ;
        RECT 91.630 120.100 92.630 121.100 ;
        RECT 92.730 120.100 93.730 121.100 ;
        RECT 93.880 120.100 95.480 121.100 ;
        RECT 95.680 120.100 96.680 121.100 ;
        RECT 96.830 120.100 97.830 121.100 ;
        RECT 91.630 118.900 92.630 119.900 ;
        RECT 92.780 118.900 93.780 119.900 ;
        RECT 93.930 118.900 95.530 119.900 ;
        RECT 95.680 118.900 96.680 119.900 ;
        RECT 96.830 118.900 97.830 119.900 ;
        RECT 4.830 112.400 5.530 113.100 ;
        RECT 4.830 111.550 5.530 112.250 ;
        RECT 4.830 110.700 5.530 111.400 ;
        RECT 23.930 112.400 24.630 113.100 ;
        RECT 24.830 112.400 25.530 113.100 ;
        RECT 23.930 111.550 24.630 112.250 ;
        RECT 24.830 111.550 25.530 112.250 ;
        RECT 23.930 110.700 24.630 111.400 ;
        RECT 24.830 110.700 25.530 111.400 ;
        RECT 4.830 108.600 5.530 109.300 ;
        RECT 4.830 107.750 5.530 108.450 ;
        RECT 4.830 106.900 5.530 107.600 ;
        RECT 43.930 112.400 44.630 113.100 ;
        RECT 44.830 112.400 45.530 113.100 ;
        RECT 43.930 111.550 44.630 112.250 ;
        RECT 44.830 111.550 45.530 112.250 ;
        RECT 43.930 110.700 44.630 111.400 ;
        RECT 44.830 110.700 45.530 111.400 ;
        RECT 23.930 108.600 24.630 109.300 ;
        RECT 24.830 108.600 25.530 109.300 ;
        RECT 23.930 107.750 24.630 108.450 ;
        RECT 24.830 107.750 25.530 108.450 ;
        RECT 23.930 106.900 24.630 107.600 ;
        RECT 24.830 106.900 25.530 107.600 ;
        RECT 63.930 112.400 64.630 113.100 ;
        RECT 64.830 112.400 65.530 113.100 ;
        RECT 63.930 111.550 64.630 112.250 ;
        RECT 64.830 111.550 65.530 112.250 ;
        RECT 63.930 110.700 64.630 111.400 ;
        RECT 64.830 110.700 65.530 111.400 ;
        RECT 43.930 108.600 44.630 109.300 ;
        RECT 44.830 108.600 45.530 109.300 ;
        RECT 43.930 107.750 44.630 108.450 ;
        RECT 44.830 107.750 45.530 108.450 ;
        RECT 43.930 106.900 44.630 107.600 ;
        RECT 44.830 106.900 45.530 107.600 ;
        RECT 83.930 112.400 84.630 113.100 ;
        RECT 84.830 112.400 85.530 113.100 ;
        RECT 83.930 111.550 84.630 112.250 ;
        RECT 84.830 111.550 85.530 112.250 ;
        RECT 83.930 110.700 84.630 111.400 ;
        RECT 84.830 110.700 85.530 111.400 ;
        RECT 63.930 108.600 64.630 109.300 ;
        RECT 64.830 108.600 65.530 109.300 ;
        RECT 63.930 107.750 64.630 108.450 ;
        RECT 64.830 107.750 65.530 108.450 ;
        RECT 63.930 106.900 64.630 107.600 ;
        RECT 64.830 106.900 65.530 107.600 ;
        RECT 103.930 112.400 104.630 113.100 ;
        RECT 103.930 111.550 104.630 112.250 ;
        RECT 103.930 110.700 104.630 111.400 ;
        RECT 110.050 110.525 110.410 110.905 ;
        RECT 110.680 110.525 111.040 110.905 ;
        RECT 111.280 110.525 111.640 110.905 ;
        RECT 83.930 108.600 84.630 109.300 ;
        RECT 84.830 108.600 85.530 109.300 ;
        RECT 83.930 107.750 84.630 108.450 ;
        RECT 84.830 107.750 85.530 108.450 ;
        RECT 83.930 106.900 84.630 107.600 ;
        RECT 84.830 106.900 85.530 107.600 ;
        RECT 110.050 109.935 110.410 110.315 ;
        RECT 110.680 109.935 111.040 110.315 ;
        RECT 111.280 109.935 111.640 110.315 ;
        RECT 103.930 108.600 104.630 109.300 ;
        RECT 103.930 107.750 104.630 108.450 ;
        RECT 103.930 106.900 104.630 107.600 ;
        RECT 11.630 100.100 12.630 101.100 ;
        RECT 12.730 100.100 13.730 101.100 ;
        RECT 13.880 100.100 15.480 101.100 ;
        RECT 15.680 100.100 16.680 101.100 ;
        RECT 16.830 100.100 17.830 101.100 ;
        RECT 11.630 98.900 12.630 99.900 ;
        RECT 12.780 98.900 13.780 99.900 ;
        RECT 13.930 98.900 15.530 99.900 ;
        RECT 15.680 98.900 16.680 99.900 ;
        RECT 16.830 98.900 17.830 99.900 ;
        RECT 31.630 100.100 32.630 101.100 ;
        RECT 32.730 100.100 33.730 101.100 ;
        RECT 33.880 100.100 35.480 101.100 ;
        RECT 35.680 100.100 36.680 101.100 ;
        RECT 36.830 100.100 37.830 101.100 ;
        RECT 31.630 98.900 32.630 99.900 ;
        RECT 32.780 98.900 33.780 99.900 ;
        RECT 33.930 98.900 35.530 99.900 ;
        RECT 35.680 98.900 36.680 99.900 ;
        RECT 36.830 98.900 37.830 99.900 ;
        RECT 51.630 100.100 52.630 101.100 ;
        RECT 52.730 100.100 53.730 101.100 ;
        RECT 53.880 100.100 55.480 101.100 ;
        RECT 55.680 100.100 56.680 101.100 ;
        RECT 56.830 100.100 57.830 101.100 ;
        RECT 51.630 98.900 52.630 99.900 ;
        RECT 52.780 98.900 53.780 99.900 ;
        RECT 53.930 98.900 55.530 99.900 ;
        RECT 55.680 98.900 56.680 99.900 ;
        RECT 56.830 98.900 57.830 99.900 ;
        RECT 71.630 100.100 72.630 101.100 ;
        RECT 72.730 100.100 73.730 101.100 ;
        RECT 73.880 100.100 75.480 101.100 ;
        RECT 75.680 100.100 76.680 101.100 ;
        RECT 76.830 100.100 77.830 101.100 ;
        RECT 71.630 98.900 72.630 99.900 ;
        RECT 72.780 98.900 73.780 99.900 ;
        RECT 73.930 98.900 75.530 99.900 ;
        RECT 75.680 98.900 76.680 99.900 ;
        RECT 76.830 98.900 77.830 99.900 ;
        RECT 91.630 100.100 92.630 101.100 ;
        RECT 92.730 100.100 93.730 101.100 ;
        RECT 93.880 100.100 95.480 101.100 ;
        RECT 95.680 100.100 96.680 101.100 ;
        RECT 96.830 100.100 97.830 101.100 ;
        RECT 91.630 98.900 92.630 99.900 ;
        RECT 92.780 98.900 93.780 99.900 ;
        RECT 93.930 98.900 95.530 99.900 ;
        RECT 95.680 98.900 96.680 99.900 ;
        RECT 96.830 98.900 97.830 99.900 ;
        RECT 4.830 92.400 5.530 93.100 ;
        RECT 4.830 91.550 5.530 92.250 ;
        RECT 4.830 90.700 5.530 91.400 ;
        RECT 23.930 92.400 24.630 93.100 ;
        RECT 24.830 92.400 25.530 93.100 ;
        RECT 23.930 91.550 24.630 92.250 ;
        RECT 24.830 91.550 25.530 92.250 ;
        RECT 23.930 90.700 24.630 91.400 ;
        RECT 24.830 90.700 25.530 91.400 ;
        RECT 4.830 88.600 5.530 89.300 ;
        RECT 4.830 87.750 5.530 88.450 ;
        RECT 4.830 86.900 5.530 87.600 ;
        RECT 43.930 92.400 44.630 93.100 ;
        RECT 44.830 92.400 45.530 93.100 ;
        RECT 43.930 91.550 44.630 92.250 ;
        RECT 44.830 91.550 45.530 92.250 ;
        RECT 43.930 90.700 44.630 91.400 ;
        RECT 44.830 90.700 45.530 91.400 ;
        RECT 23.930 88.600 24.630 89.300 ;
        RECT 24.830 88.600 25.530 89.300 ;
        RECT 23.930 87.750 24.630 88.450 ;
        RECT 24.830 87.750 25.530 88.450 ;
        RECT 23.930 86.900 24.630 87.600 ;
        RECT 24.830 86.900 25.530 87.600 ;
        RECT 63.930 92.400 64.630 93.100 ;
        RECT 64.830 92.400 65.530 93.100 ;
        RECT 63.930 91.550 64.630 92.250 ;
        RECT 64.830 91.550 65.530 92.250 ;
        RECT 63.930 90.700 64.630 91.400 ;
        RECT 64.830 90.700 65.530 91.400 ;
        RECT 43.930 88.600 44.630 89.300 ;
        RECT 44.830 88.600 45.530 89.300 ;
        RECT 43.930 87.750 44.630 88.450 ;
        RECT 44.830 87.750 45.530 88.450 ;
        RECT 43.930 86.900 44.630 87.600 ;
        RECT 44.830 86.900 45.530 87.600 ;
        RECT 83.930 92.400 84.630 93.100 ;
        RECT 84.830 92.400 85.530 93.100 ;
        RECT 83.930 91.550 84.630 92.250 ;
        RECT 84.830 91.550 85.530 92.250 ;
        RECT 83.930 90.700 84.630 91.400 ;
        RECT 84.830 90.700 85.530 91.400 ;
        RECT 63.930 88.600 64.630 89.300 ;
        RECT 64.830 88.600 65.530 89.300 ;
        RECT 63.930 87.750 64.630 88.450 ;
        RECT 64.830 87.750 65.530 88.450 ;
        RECT 63.930 86.900 64.630 87.600 ;
        RECT 64.830 86.900 65.530 87.600 ;
        RECT 103.930 92.400 104.630 93.100 ;
        RECT 103.930 91.550 104.630 92.250 ;
        RECT 103.930 90.700 104.630 91.400 ;
        RECT 83.930 88.600 84.630 89.300 ;
        RECT 84.830 88.600 85.530 89.300 ;
        RECT 83.930 87.750 84.630 88.450 ;
        RECT 84.830 87.750 85.530 88.450 ;
        RECT 83.930 86.900 84.630 87.600 ;
        RECT 84.830 86.900 85.530 87.600 ;
        RECT 110.050 89.990 110.410 90.370 ;
        RECT 110.680 89.990 111.040 90.370 ;
        RECT 111.280 89.990 111.640 90.370 ;
        RECT 110.050 89.400 110.410 89.780 ;
        RECT 110.680 89.400 111.040 89.780 ;
        RECT 111.280 89.400 111.640 89.780 ;
        RECT 103.930 88.600 104.630 89.300 ;
        RECT 103.930 87.750 104.630 88.450 ;
        RECT 103.930 86.900 104.630 87.600 ;
        RECT 11.630 80.100 12.630 81.100 ;
        RECT 12.730 80.100 13.730 81.100 ;
        RECT 13.880 80.100 15.480 81.100 ;
        RECT 15.680 80.100 16.680 81.100 ;
        RECT 16.830 80.100 17.830 81.100 ;
        RECT 11.630 78.900 12.630 79.900 ;
        RECT 12.780 78.900 13.780 79.900 ;
        RECT 13.930 78.900 15.530 79.900 ;
        RECT 15.680 78.900 16.680 79.900 ;
        RECT 16.830 78.900 17.830 79.900 ;
        RECT 31.630 80.100 32.630 81.100 ;
        RECT 32.730 80.100 33.730 81.100 ;
        RECT 33.880 80.100 35.480 81.100 ;
        RECT 35.680 80.100 36.680 81.100 ;
        RECT 36.830 80.100 37.830 81.100 ;
        RECT 31.630 78.900 32.630 79.900 ;
        RECT 32.780 78.900 33.780 79.900 ;
        RECT 33.930 78.900 35.530 79.900 ;
        RECT 35.680 78.900 36.680 79.900 ;
        RECT 36.830 78.900 37.830 79.900 ;
        RECT 51.630 80.100 52.630 81.100 ;
        RECT 52.730 80.100 53.730 81.100 ;
        RECT 53.880 80.100 55.480 81.100 ;
        RECT 55.680 80.100 56.680 81.100 ;
        RECT 56.830 80.100 57.830 81.100 ;
        RECT 51.630 78.900 52.630 79.900 ;
        RECT 52.780 78.900 53.780 79.900 ;
        RECT 53.930 78.900 55.530 79.900 ;
        RECT 55.680 78.900 56.680 79.900 ;
        RECT 56.830 78.900 57.830 79.900 ;
        RECT 71.630 80.100 72.630 81.100 ;
        RECT 72.730 80.100 73.730 81.100 ;
        RECT 73.880 80.100 75.480 81.100 ;
        RECT 75.680 80.100 76.680 81.100 ;
        RECT 76.830 80.100 77.830 81.100 ;
        RECT 71.630 78.900 72.630 79.900 ;
        RECT 72.780 78.900 73.780 79.900 ;
        RECT 73.930 78.900 75.530 79.900 ;
        RECT 75.680 78.900 76.680 79.900 ;
        RECT 76.830 78.900 77.830 79.900 ;
        RECT 91.630 80.100 92.630 81.100 ;
        RECT 92.730 80.100 93.730 81.100 ;
        RECT 93.880 80.100 95.480 81.100 ;
        RECT 95.680 80.100 96.680 81.100 ;
        RECT 96.830 80.100 97.830 81.100 ;
        RECT 91.630 78.900 92.630 79.900 ;
        RECT 92.780 78.900 93.780 79.900 ;
        RECT 93.930 78.900 95.530 79.900 ;
        RECT 95.680 78.900 96.680 79.900 ;
        RECT 96.830 78.900 97.830 79.900 ;
        RECT 4.830 72.400 5.530 73.100 ;
        RECT 4.830 71.550 5.530 72.250 ;
        RECT 4.830 70.700 5.530 71.400 ;
        RECT 23.930 72.400 24.630 73.100 ;
        RECT 24.830 72.400 25.530 73.100 ;
        RECT 23.930 71.550 24.630 72.250 ;
        RECT 24.830 71.550 25.530 72.250 ;
        RECT 23.930 70.700 24.630 71.400 ;
        RECT 24.830 70.700 25.530 71.400 ;
        RECT 4.830 68.600 5.530 69.300 ;
        RECT 4.830 67.750 5.530 68.450 ;
        RECT 4.830 66.900 5.530 67.600 ;
        RECT 43.930 72.400 44.630 73.100 ;
        RECT 44.830 72.400 45.530 73.100 ;
        RECT 43.930 71.550 44.630 72.250 ;
        RECT 44.830 71.550 45.530 72.250 ;
        RECT 43.930 70.700 44.630 71.400 ;
        RECT 44.830 70.700 45.530 71.400 ;
        RECT 23.930 68.600 24.630 69.300 ;
        RECT 24.830 68.600 25.530 69.300 ;
        RECT 23.930 67.750 24.630 68.450 ;
        RECT 24.830 67.750 25.530 68.450 ;
        RECT 23.930 66.900 24.630 67.600 ;
        RECT 24.830 66.900 25.530 67.600 ;
        RECT 63.930 72.400 64.630 73.100 ;
        RECT 64.830 72.400 65.530 73.100 ;
        RECT 63.930 71.550 64.630 72.250 ;
        RECT 64.830 71.550 65.530 72.250 ;
        RECT 63.930 70.700 64.630 71.400 ;
        RECT 64.830 70.700 65.530 71.400 ;
        RECT 43.930 68.600 44.630 69.300 ;
        RECT 44.830 68.600 45.530 69.300 ;
        RECT 43.930 67.750 44.630 68.450 ;
        RECT 44.830 67.750 45.530 68.450 ;
        RECT 43.930 66.900 44.630 67.600 ;
        RECT 44.830 66.900 45.530 67.600 ;
        RECT 83.930 72.400 84.630 73.100 ;
        RECT 84.830 72.400 85.530 73.100 ;
        RECT 83.930 71.550 84.630 72.250 ;
        RECT 84.830 71.550 85.530 72.250 ;
        RECT 83.930 70.700 84.630 71.400 ;
        RECT 84.830 70.700 85.530 71.400 ;
        RECT 63.930 68.600 64.630 69.300 ;
        RECT 64.830 68.600 65.530 69.300 ;
        RECT 63.930 67.750 64.630 68.450 ;
        RECT 64.830 67.750 65.530 68.450 ;
        RECT 63.930 66.900 64.630 67.600 ;
        RECT 64.830 66.900 65.530 67.600 ;
        RECT 103.930 72.400 104.630 73.100 ;
        RECT 103.930 71.550 104.630 72.250 ;
        RECT 103.930 70.700 104.630 71.400 ;
        RECT 110.050 70.900 110.410 71.280 ;
        RECT 110.680 70.900 111.040 71.280 ;
        RECT 111.280 70.900 111.640 71.280 ;
        RECT 83.930 68.600 84.630 69.300 ;
        RECT 84.830 68.600 85.530 69.300 ;
        RECT 83.930 67.750 84.630 68.450 ;
        RECT 84.830 67.750 85.530 68.450 ;
        RECT 83.930 66.900 84.630 67.600 ;
        RECT 84.830 66.900 85.530 67.600 ;
        RECT 110.050 70.310 110.410 70.690 ;
        RECT 110.680 70.310 111.040 70.690 ;
        RECT 111.280 70.310 111.640 70.690 ;
        RECT 103.930 68.600 104.630 69.300 ;
        RECT 103.930 67.750 104.630 68.450 ;
        RECT 103.930 66.900 104.630 67.600 ;
        RECT 11.630 60.100 12.630 61.100 ;
        RECT 12.730 60.100 13.730 61.100 ;
        RECT 13.880 60.100 15.480 61.100 ;
        RECT 15.680 60.100 16.680 61.100 ;
        RECT 16.830 60.100 17.830 61.100 ;
        RECT 11.630 58.900 12.630 59.900 ;
        RECT 12.780 58.900 13.780 59.900 ;
        RECT 13.930 58.900 15.530 59.900 ;
        RECT 15.680 58.900 16.680 59.900 ;
        RECT 16.830 58.900 17.830 59.900 ;
        RECT 31.630 60.100 32.630 61.100 ;
        RECT 32.730 60.100 33.730 61.100 ;
        RECT 33.880 60.100 35.480 61.100 ;
        RECT 35.680 60.100 36.680 61.100 ;
        RECT 36.830 60.100 37.830 61.100 ;
        RECT 31.630 58.900 32.630 59.900 ;
        RECT 32.780 58.900 33.780 59.900 ;
        RECT 33.930 58.900 35.530 59.900 ;
        RECT 35.680 58.900 36.680 59.900 ;
        RECT 36.830 58.900 37.830 59.900 ;
        RECT 51.630 60.100 52.630 61.100 ;
        RECT 52.730 60.100 53.730 61.100 ;
        RECT 53.880 60.100 55.480 61.100 ;
        RECT 55.680 60.100 56.680 61.100 ;
        RECT 56.830 60.100 57.830 61.100 ;
        RECT 51.630 58.900 52.630 59.900 ;
        RECT 52.780 58.900 53.780 59.900 ;
        RECT 53.930 58.900 55.530 59.900 ;
        RECT 55.680 58.900 56.680 59.900 ;
        RECT 56.830 58.900 57.830 59.900 ;
        RECT 71.630 60.100 72.630 61.100 ;
        RECT 72.730 60.100 73.730 61.100 ;
        RECT 73.880 60.100 75.480 61.100 ;
        RECT 75.680 60.100 76.680 61.100 ;
        RECT 76.830 60.100 77.830 61.100 ;
        RECT 71.630 58.900 72.630 59.900 ;
        RECT 72.780 58.900 73.780 59.900 ;
        RECT 73.930 58.900 75.530 59.900 ;
        RECT 75.680 58.900 76.680 59.900 ;
        RECT 76.830 58.900 77.830 59.900 ;
        RECT 91.630 60.100 92.630 61.100 ;
        RECT 92.730 60.100 93.730 61.100 ;
        RECT 93.880 60.100 95.480 61.100 ;
        RECT 95.680 60.100 96.680 61.100 ;
        RECT 96.830 60.100 97.830 61.100 ;
        RECT 91.630 58.900 92.630 59.900 ;
        RECT 92.780 58.900 93.780 59.900 ;
        RECT 93.930 58.900 95.530 59.900 ;
        RECT 95.680 58.900 96.680 59.900 ;
        RECT 96.830 58.900 97.830 59.900 ;
        RECT 4.830 52.400 5.530 53.100 ;
        RECT 4.830 51.550 5.530 52.250 ;
        RECT 4.830 50.700 5.530 51.400 ;
        RECT 23.930 52.400 24.630 53.100 ;
        RECT 24.830 52.400 25.530 53.100 ;
        RECT 23.930 51.550 24.630 52.250 ;
        RECT 24.830 51.550 25.530 52.250 ;
        RECT 23.930 50.700 24.630 51.400 ;
        RECT 24.830 50.700 25.530 51.400 ;
        RECT 4.830 48.600 5.530 49.300 ;
        RECT 4.830 47.750 5.530 48.450 ;
        RECT 4.830 46.900 5.530 47.600 ;
        RECT 43.930 52.400 44.630 53.100 ;
        RECT 44.830 52.400 45.530 53.100 ;
        RECT 43.930 51.550 44.630 52.250 ;
        RECT 44.830 51.550 45.530 52.250 ;
        RECT 43.930 50.700 44.630 51.400 ;
        RECT 44.830 50.700 45.530 51.400 ;
        RECT 23.930 48.600 24.630 49.300 ;
        RECT 24.830 48.600 25.530 49.300 ;
        RECT 23.930 47.750 24.630 48.450 ;
        RECT 24.830 47.750 25.530 48.450 ;
        RECT 23.930 46.900 24.630 47.600 ;
        RECT 24.830 46.900 25.530 47.600 ;
        RECT 63.930 52.400 64.630 53.100 ;
        RECT 64.830 52.400 65.530 53.100 ;
        RECT 63.930 51.550 64.630 52.250 ;
        RECT 64.830 51.550 65.530 52.250 ;
        RECT 63.930 50.700 64.630 51.400 ;
        RECT 64.830 50.700 65.530 51.400 ;
        RECT 43.930 48.600 44.630 49.300 ;
        RECT 44.830 48.600 45.530 49.300 ;
        RECT 43.930 47.750 44.630 48.450 ;
        RECT 44.830 47.750 45.530 48.450 ;
        RECT 43.930 46.900 44.630 47.600 ;
        RECT 44.830 46.900 45.530 47.600 ;
        RECT 83.930 52.400 84.630 53.100 ;
        RECT 84.830 52.400 85.530 53.100 ;
        RECT 83.930 51.550 84.630 52.250 ;
        RECT 84.830 51.550 85.530 52.250 ;
        RECT 83.930 50.700 84.630 51.400 ;
        RECT 84.830 50.700 85.530 51.400 ;
        RECT 63.930 48.600 64.630 49.300 ;
        RECT 64.830 48.600 65.530 49.300 ;
        RECT 63.930 47.750 64.630 48.450 ;
        RECT 64.830 47.750 65.530 48.450 ;
        RECT 63.930 46.900 64.630 47.600 ;
        RECT 64.830 46.900 65.530 47.600 ;
        RECT 103.930 52.400 104.630 53.100 ;
        RECT 103.930 51.550 104.630 52.250 ;
        RECT 103.930 50.700 104.630 51.400 ;
        RECT 110.050 51.080 110.410 51.460 ;
        RECT 110.680 51.080 111.040 51.460 ;
        RECT 111.280 51.080 111.640 51.460 ;
        RECT 110.050 50.490 110.410 50.870 ;
        RECT 110.680 50.490 111.040 50.870 ;
        RECT 111.280 50.490 111.640 50.870 ;
        RECT 83.930 48.600 84.630 49.300 ;
        RECT 84.830 48.600 85.530 49.300 ;
        RECT 83.930 47.750 84.630 48.450 ;
        RECT 84.830 47.750 85.530 48.450 ;
        RECT 83.930 46.900 84.630 47.600 ;
        RECT 84.830 46.900 85.530 47.600 ;
        RECT 103.930 48.600 104.630 49.300 ;
        RECT 103.930 47.750 104.630 48.450 ;
        RECT 103.930 46.900 104.630 47.600 ;
        RECT 11.630 40.100 12.630 41.100 ;
        RECT 12.730 40.100 13.730 41.100 ;
        RECT 13.880 40.100 15.480 41.100 ;
        RECT 15.680 40.100 16.680 41.100 ;
        RECT 16.830 40.100 17.830 41.100 ;
        RECT 11.630 38.900 12.630 39.900 ;
        RECT 12.780 38.900 13.780 39.900 ;
        RECT 13.930 38.900 15.530 39.900 ;
        RECT 15.680 38.900 16.680 39.900 ;
        RECT 16.830 38.900 17.830 39.900 ;
        RECT 31.630 40.100 32.630 41.100 ;
        RECT 32.730 40.100 33.730 41.100 ;
        RECT 33.880 40.100 35.480 41.100 ;
        RECT 35.680 40.100 36.680 41.100 ;
        RECT 36.830 40.100 37.830 41.100 ;
        RECT 31.630 38.900 32.630 39.900 ;
        RECT 32.780 38.900 33.780 39.900 ;
        RECT 33.930 38.900 35.530 39.900 ;
        RECT 35.680 38.900 36.680 39.900 ;
        RECT 36.830 38.900 37.830 39.900 ;
        RECT 51.630 40.100 52.630 41.100 ;
        RECT 52.730 40.100 53.730 41.100 ;
        RECT 53.880 40.100 55.480 41.100 ;
        RECT 55.680 40.100 56.680 41.100 ;
        RECT 56.830 40.100 57.830 41.100 ;
        RECT 51.630 38.900 52.630 39.900 ;
        RECT 52.780 38.900 53.780 39.900 ;
        RECT 53.930 38.900 55.530 39.900 ;
        RECT 55.680 38.900 56.680 39.900 ;
        RECT 56.830 38.900 57.830 39.900 ;
        RECT 71.630 40.100 72.630 41.100 ;
        RECT 72.730 40.100 73.730 41.100 ;
        RECT 73.880 40.100 75.480 41.100 ;
        RECT 75.680 40.100 76.680 41.100 ;
        RECT 76.830 40.100 77.830 41.100 ;
        RECT 71.630 38.900 72.630 39.900 ;
        RECT 72.780 38.900 73.780 39.900 ;
        RECT 73.930 38.900 75.530 39.900 ;
        RECT 75.680 38.900 76.680 39.900 ;
        RECT 76.830 38.900 77.830 39.900 ;
        RECT 91.630 40.100 92.630 41.100 ;
        RECT 92.730 40.100 93.730 41.100 ;
        RECT 93.880 40.100 95.480 41.100 ;
        RECT 95.680 40.100 96.680 41.100 ;
        RECT 96.830 40.100 97.830 41.100 ;
        RECT 91.630 38.900 92.630 39.900 ;
        RECT 92.780 38.900 93.780 39.900 ;
        RECT 93.930 38.900 95.530 39.900 ;
        RECT 95.680 38.900 96.680 39.900 ;
        RECT 96.830 38.900 97.830 39.900 ;
        RECT 4.830 32.400 5.530 33.100 ;
        RECT 4.830 31.550 5.530 32.250 ;
        RECT 4.830 30.700 5.530 31.400 ;
        RECT 23.930 32.400 24.630 33.100 ;
        RECT 24.830 32.400 25.530 33.100 ;
        RECT 23.930 31.550 24.630 32.250 ;
        RECT 24.830 31.550 25.530 32.250 ;
        RECT 23.930 30.700 24.630 31.400 ;
        RECT 24.830 30.700 25.530 31.400 ;
        RECT 4.830 28.600 5.530 29.300 ;
        RECT 4.830 27.750 5.530 28.450 ;
        RECT 4.830 26.900 5.530 27.600 ;
        RECT 43.930 32.400 44.630 33.100 ;
        RECT 44.830 32.400 45.530 33.100 ;
        RECT 43.930 31.550 44.630 32.250 ;
        RECT 44.830 31.550 45.530 32.250 ;
        RECT 43.930 30.700 44.630 31.400 ;
        RECT 44.830 30.700 45.530 31.400 ;
        RECT 23.930 28.600 24.630 29.300 ;
        RECT 24.830 28.600 25.530 29.300 ;
        RECT 23.930 27.750 24.630 28.450 ;
        RECT 24.830 27.750 25.530 28.450 ;
        RECT 23.930 26.900 24.630 27.600 ;
        RECT 24.830 26.900 25.530 27.600 ;
        RECT 63.930 32.400 64.630 33.100 ;
        RECT 64.830 32.400 65.530 33.100 ;
        RECT 63.930 31.550 64.630 32.250 ;
        RECT 64.830 31.550 65.530 32.250 ;
        RECT 63.930 30.700 64.630 31.400 ;
        RECT 64.830 30.700 65.530 31.400 ;
        RECT 43.930 28.600 44.630 29.300 ;
        RECT 44.830 28.600 45.530 29.300 ;
        RECT 43.930 27.750 44.630 28.450 ;
        RECT 44.830 27.750 45.530 28.450 ;
        RECT 43.930 26.900 44.630 27.600 ;
        RECT 44.830 26.900 45.530 27.600 ;
        RECT 83.930 32.400 84.630 33.100 ;
        RECT 84.830 32.400 85.530 33.100 ;
        RECT 83.930 31.550 84.630 32.250 ;
        RECT 84.830 31.550 85.530 32.250 ;
        RECT 83.930 30.700 84.630 31.400 ;
        RECT 84.830 30.700 85.530 31.400 ;
        RECT 63.930 28.600 64.630 29.300 ;
        RECT 64.830 28.600 65.530 29.300 ;
        RECT 63.930 27.750 64.630 28.450 ;
        RECT 64.830 27.750 65.530 28.450 ;
        RECT 63.930 26.900 64.630 27.600 ;
        RECT 64.830 26.900 65.530 27.600 ;
        RECT 103.930 32.400 104.630 33.100 ;
        RECT 103.930 31.550 104.630 32.250 ;
        RECT 103.930 30.700 104.630 31.400 ;
        RECT 110.050 31.020 110.410 31.400 ;
        RECT 110.680 31.020 111.040 31.400 ;
        RECT 111.280 31.020 111.640 31.400 ;
        RECT 83.930 28.600 84.630 29.300 ;
        RECT 84.830 28.600 85.530 29.300 ;
        RECT 83.930 27.750 84.630 28.450 ;
        RECT 84.830 27.750 85.530 28.450 ;
        RECT 83.930 26.900 84.630 27.600 ;
        RECT 84.830 26.900 85.530 27.600 ;
        RECT 110.050 30.430 110.410 30.810 ;
        RECT 110.680 30.430 111.040 30.810 ;
        RECT 111.280 30.430 111.640 30.810 ;
        RECT 103.930 28.600 104.630 29.300 ;
        RECT 103.930 27.750 104.630 28.450 ;
        RECT 103.930 26.900 104.630 27.600 ;
        RECT 11.630 20.100 12.630 21.100 ;
        RECT 12.730 20.100 13.730 21.100 ;
        RECT 13.880 20.100 15.480 21.100 ;
        RECT 15.680 20.100 16.680 21.100 ;
        RECT 16.830 20.100 17.830 21.100 ;
        RECT 11.630 18.900 12.630 19.900 ;
        RECT 12.780 18.900 13.780 19.900 ;
        RECT 13.930 18.900 15.530 19.900 ;
        RECT 15.680 18.900 16.680 19.900 ;
        RECT 16.830 18.900 17.830 19.900 ;
        RECT 31.630 20.100 32.630 21.100 ;
        RECT 32.730 20.100 33.730 21.100 ;
        RECT 33.880 20.100 35.480 21.100 ;
        RECT 35.680 20.100 36.680 21.100 ;
        RECT 36.830 20.100 37.830 21.100 ;
        RECT 31.630 18.900 32.630 19.900 ;
        RECT 32.780 18.900 33.780 19.900 ;
        RECT 33.930 18.900 35.530 19.900 ;
        RECT 35.680 18.900 36.680 19.900 ;
        RECT 36.830 18.900 37.830 19.900 ;
        RECT 51.630 20.100 52.630 21.100 ;
        RECT 52.730 20.100 53.730 21.100 ;
        RECT 53.880 20.100 55.480 21.100 ;
        RECT 55.680 20.100 56.680 21.100 ;
        RECT 56.830 20.100 57.830 21.100 ;
        RECT 51.630 18.900 52.630 19.900 ;
        RECT 52.780 18.900 53.780 19.900 ;
        RECT 53.930 18.900 55.530 19.900 ;
        RECT 55.680 18.900 56.680 19.900 ;
        RECT 56.830 18.900 57.830 19.900 ;
        RECT 71.630 20.100 72.630 21.100 ;
        RECT 72.730 20.100 73.730 21.100 ;
        RECT 73.880 20.100 75.480 21.100 ;
        RECT 75.680 20.100 76.680 21.100 ;
        RECT 76.830 20.100 77.830 21.100 ;
        RECT 71.630 18.900 72.630 19.900 ;
        RECT 72.780 18.900 73.780 19.900 ;
        RECT 73.930 18.900 75.530 19.900 ;
        RECT 75.680 18.900 76.680 19.900 ;
        RECT 76.830 18.900 77.830 19.900 ;
        RECT 91.630 20.100 92.630 21.100 ;
        RECT 92.730 20.100 93.730 21.100 ;
        RECT 93.880 20.100 95.480 21.100 ;
        RECT 95.680 20.100 96.680 21.100 ;
        RECT 96.830 20.100 97.830 21.100 ;
        RECT 91.630 18.900 92.630 19.900 ;
        RECT 92.780 18.900 93.780 19.900 ;
        RECT 93.930 18.900 95.530 19.900 ;
        RECT 95.680 18.900 96.680 19.900 ;
        RECT 96.830 18.900 97.830 19.900 ;
        RECT 4.830 12.400 5.530 13.100 ;
        RECT 4.830 11.550 5.530 12.250 ;
        RECT 4.830 10.700 5.530 11.400 ;
        RECT 23.930 12.400 24.630 13.100 ;
        RECT 24.830 12.400 25.530 13.100 ;
        RECT 23.930 11.550 24.630 12.250 ;
        RECT 24.830 11.550 25.530 12.250 ;
        RECT 23.930 10.700 24.630 11.400 ;
        RECT 24.830 10.700 25.530 11.400 ;
        RECT 4.830 8.600 5.530 9.300 ;
        RECT 4.830 7.750 5.530 8.450 ;
        RECT 4.830 6.900 5.530 7.600 ;
        RECT 43.930 12.400 44.630 13.100 ;
        RECT 44.830 12.400 45.530 13.100 ;
        RECT 43.930 11.550 44.630 12.250 ;
        RECT 44.830 11.550 45.530 12.250 ;
        RECT 43.930 10.700 44.630 11.400 ;
        RECT 44.830 10.700 45.530 11.400 ;
        RECT 23.930 8.600 24.630 9.300 ;
        RECT 24.830 8.600 25.530 9.300 ;
        RECT 23.930 7.750 24.630 8.450 ;
        RECT 24.830 7.750 25.530 8.450 ;
        RECT 23.930 6.900 24.630 7.600 ;
        RECT 24.830 6.900 25.530 7.600 ;
        RECT 63.930 12.400 64.630 13.100 ;
        RECT 64.830 12.400 65.530 13.100 ;
        RECT 63.930 11.550 64.630 12.250 ;
        RECT 64.830 11.550 65.530 12.250 ;
        RECT 63.930 10.700 64.630 11.400 ;
        RECT 64.830 10.700 65.530 11.400 ;
        RECT 43.930 8.600 44.630 9.300 ;
        RECT 44.830 8.600 45.530 9.300 ;
        RECT 43.930 7.750 44.630 8.450 ;
        RECT 44.830 7.750 45.530 8.450 ;
        RECT 43.930 6.900 44.630 7.600 ;
        RECT 44.830 6.900 45.530 7.600 ;
        RECT 83.930 12.400 84.630 13.100 ;
        RECT 84.830 12.400 85.530 13.100 ;
        RECT 83.930 11.550 84.630 12.250 ;
        RECT 84.830 11.550 85.530 12.250 ;
        RECT 83.930 10.700 84.630 11.400 ;
        RECT 84.830 10.700 85.530 11.400 ;
        RECT 63.930 8.600 64.630 9.300 ;
        RECT 64.830 8.600 65.530 9.300 ;
        RECT 63.930 7.750 64.630 8.450 ;
        RECT 64.830 7.750 65.530 8.450 ;
        RECT 63.930 6.900 64.630 7.600 ;
        RECT 64.830 6.900 65.530 7.600 ;
        RECT 103.930 12.400 104.630 13.100 ;
        RECT 103.930 11.550 104.630 12.250 ;
        RECT 103.930 10.700 104.630 11.400 ;
        RECT 110.050 11.020 110.410 11.400 ;
        RECT 110.680 11.020 111.040 11.400 ;
        RECT 111.280 11.020 111.640 11.400 ;
        RECT 83.930 8.600 84.630 9.300 ;
        RECT 84.830 8.600 85.530 9.300 ;
        RECT 83.930 7.750 84.630 8.450 ;
        RECT 84.830 7.750 85.530 8.450 ;
        RECT 83.930 6.900 84.630 7.600 ;
        RECT 84.830 6.900 85.530 7.600 ;
        RECT 110.050 10.430 110.410 10.810 ;
        RECT 110.680 10.430 111.040 10.810 ;
        RECT 111.280 10.430 111.640 10.810 ;
        RECT 103.930 8.600 104.630 9.300 ;
        RECT 103.930 7.750 104.630 8.450 ;
        RECT 103.930 6.900 104.630 7.600 ;
        RECT 11.630 0.100 12.630 1.100 ;
        RECT 12.730 0.100 13.730 1.100 ;
        RECT 13.880 0.100 15.480 1.100 ;
        RECT 15.680 0.100 16.680 1.100 ;
        RECT 16.830 0.100 17.830 1.100 ;
        RECT 31.630 0.100 32.630 1.100 ;
        RECT 32.730 0.100 33.730 1.100 ;
        RECT 33.880 0.100 35.480 1.100 ;
        RECT 35.680 0.100 36.680 1.100 ;
        RECT 36.830 0.100 37.830 1.100 ;
        RECT 51.630 0.100 52.630 1.100 ;
        RECT 52.730 0.100 53.730 1.100 ;
        RECT 53.880 0.100 55.480 1.100 ;
        RECT 55.680 0.100 56.680 1.100 ;
        RECT 56.830 0.100 57.830 1.100 ;
        RECT 71.630 0.100 72.630 1.100 ;
        RECT 72.730 0.100 73.730 1.100 ;
        RECT 73.880 0.100 75.480 1.100 ;
        RECT 75.680 0.100 76.680 1.100 ;
        RECT 76.830 0.100 77.830 1.100 ;
        RECT 91.630 0.100 92.630 1.100 ;
        RECT 92.730 0.100 93.730 1.100 ;
        RECT 93.880 0.100 95.480 1.100 ;
        RECT 95.680 0.100 96.680 1.100 ;
        RECT 96.830 0.100 97.830 1.100 ;
      LAYER met2 ;
        RECT 11.530 379.100 17.930 380.000 ;
        RECT 31.530 379.100 37.930 380.000 ;
        RECT 51.530 379.100 57.930 380.000 ;
        RECT 71.530 379.100 77.930 380.000 ;
        RECT 91.530 379.100 97.930 380.000 ;
        RECT 9.630 378.600 19.830 379.100 ;
        RECT 29.630 378.600 39.830 379.100 ;
        RECT 49.630 378.600 59.830 379.100 ;
        RECT 69.630 378.600 79.830 379.100 ;
        RECT 89.630 378.600 99.830 379.100 ;
        RECT 6.530 378.550 22.930 378.600 ;
        RECT 6.530 378.000 10.330 378.550 ;
        RECT 10.030 377.550 10.330 378.000 ;
        RECT 6.480 377.400 10.330 377.550 ;
        RECT 10.030 376.950 10.330 377.400 ;
        RECT 6.480 376.800 10.330 376.950 ;
        RECT 10.030 376.350 10.330 376.800 ;
        RECT 6.480 376.200 10.330 376.350 ;
        RECT 10.030 375.750 10.330 376.200 ;
        RECT 6.480 375.600 10.330 375.750 ;
        RECT 10.030 375.150 10.330 375.600 ;
        RECT 6.480 375.000 10.330 375.150 ;
        RECT 10.030 374.550 10.330 375.000 ;
        RECT 6.480 374.400 10.330 374.550 ;
        RECT 10.030 373.950 10.330 374.400 ;
        RECT 6.480 373.800 10.330 373.950 ;
        RECT 10.030 373.350 10.330 373.800 ;
        RECT 6.480 373.200 10.330 373.350 ;
        RECT 4.730 366.800 5.630 373.200 ;
        RECT 10.030 372.750 10.330 373.200 ;
        RECT 6.480 372.600 10.330 372.750 ;
        RECT 10.030 372.150 10.330 372.600 ;
        RECT 6.480 372.000 10.330 372.150 ;
        RECT 10.030 371.550 10.330 372.000 ;
        RECT 6.480 371.400 10.330 371.550 ;
        RECT 10.030 370.950 10.330 371.400 ;
        RECT 6.480 370.800 10.330 370.950 ;
        RECT 10.030 370.350 10.330 370.800 ;
        RECT 10.780 370.350 10.930 378.550 ;
        RECT 11.380 370.350 11.530 378.550 ;
        RECT 11.980 370.350 12.130 378.550 ;
        RECT 12.580 370.350 12.730 378.550 ;
        RECT 13.180 370.350 13.330 378.550 ;
        RECT 13.780 370.350 13.930 378.550 ;
        RECT 10.030 369.200 10.330 369.650 ;
        RECT 6.480 369.050 10.330 369.200 ;
        RECT 10.030 368.600 10.330 369.050 ;
        RECT 6.480 368.450 10.330 368.600 ;
        RECT 10.030 368.000 10.330 368.450 ;
        RECT 6.480 367.850 10.330 368.000 ;
        RECT 10.030 367.400 10.330 367.850 ;
        RECT 6.480 367.250 10.330 367.400 ;
        RECT 10.030 366.800 10.330 367.250 ;
        RECT 6.480 366.650 10.330 366.800 ;
        RECT 10.030 366.200 10.330 366.650 ;
        RECT 6.480 366.050 10.330 366.200 ;
        RECT 10.030 365.600 10.330 366.050 ;
        RECT 6.480 365.450 10.330 365.600 ;
        RECT 10.030 365.000 10.330 365.450 ;
        RECT 6.480 364.850 10.330 365.000 ;
        RECT 10.030 364.400 10.330 364.850 ;
        RECT 6.480 364.250 10.330 364.400 ;
        RECT 10.030 363.800 10.330 364.250 ;
        RECT 6.480 363.650 10.330 363.800 ;
        RECT 10.030 363.200 10.330 363.650 ;
        RECT 6.480 363.050 10.330 363.200 ;
        RECT 10.030 362.600 10.330 363.050 ;
        RECT 6.480 362.450 10.330 362.600 ;
        RECT 10.030 362.000 10.330 362.450 ;
        RECT 6.530 361.450 10.330 362.000 ;
        RECT 10.780 361.450 10.930 369.650 ;
        RECT 11.380 361.450 11.530 369.650 ;
        RECT 11.980 361.450 12.130 369.650 ;
        RECT 12.580 361.450 12.730 369.650 ;
        RECT 13.180 361.450 13.330 369.650 ;
        RECT 13.780 361.450 13.930 369.650 ;
        RECT 14.380 361.450 15.080 378.550 ;
        RECT 15.530 370.350 15.680 378.550 ;
        RECT 16.130 370.350 16.280 378.550 ;
        RECT 16.730 370.350 16.880 378.550 ;
        RECT 17.330 370.350 17.480 378.550 ;
        RECT 17.930 370.350 18.080 378.550 ;
        RECT 18.530 370.350 18.680 378.550 ;
        RECT 19.130 378.000 22.930 378.550 ;
        RECT 26.530 378.550 42.930 378.600 ;
        RECT 26.530 378.000 30.330 378.550 ;
        RECT 19.130 377.550 19.430 378.000 ;
        RECT 30.030 377.550 30.330 378.000 ;
        RECT 19.130 377.400 22.980 377.550 ;
        RECT 26.480 377.400 30.330 377.550 ;
        RECT 19.130 376.950 19.430 377.400 ;
        RECT 30.030 376.950 30.330 377.400 ;
        RECT 19.130 376.800 22.980 376.950 ;
        RECT 26.480 376.800 30.330 376.950 ;
        RECT 19.130 376.350 19.430 376.800 ;
        RECT 30.030 376.350 30.330 376.800 ;
        RECT 19.130 376.200 22.980 376.350 ;
        RECT 26.480 376.200 30.330 376.350 ;
        RECT 19.130 375.750 19.430 376.200 ;
        RECT 30.030 375.750 30.330 376.200 ;
        RECT 19.130 375.600 22.980 375.750 ;
        RECT 26.480 375.600 30.330 375.750 ;
        RECT 19.130 375.150 19.430 375.600 ;
        RECT 30.030 375.150 30.330 375.600 ;
        RECT 19.130 375.000 22.980 375.150 ;
        RECT 26.480 375.000 30.330 375.150 ;
        RECT 19.130 374.550 19.430 375.000 ;
        RECT 30.030 374.550 30.330 375.000 ;
        RECT 19.130 374.400 22.980 374.550 ;
        RECT 26.480 374.400 30.330 374.550 ;
        RECT 19.130 373.950 19.430 374.400 ;
        RECT 30.030 373.950 30.330 374.400 ;
        RECT 19.130 373.800 22.980 373.950 ;
        RECT 26.480 373.800 30.330 373.950 ;
        RECT 19.130 373.350 19.430 373.800 ;
        RECT 30.030 373.350 30.330 373.800 ;
        RECT 19.130 373.200 22.980 373.350 ;
        RECT 26.480 373.200 30.330 373.350 ;
        RECT 19.130 372.750 19.430 373.200 ;
        RECT 19.130 372.600 22.980 372.750 ;
        RECT 19.130 372.150 19.430 372.600 ;
        RECT 19.130 372.000 22.980 372.150 ;
        RECT 19.130 371.550 19.430 372.000 ;
        RECT 19.130 371.400 22.980 371.550 ;
        RECT 19.130 370.950 19.430 371.400 ;
        RECT 19.130 370.800 22.980 370.950 ;
        RECT 19.130 370.350 19.430 370.800 ;
        RECT 15.530 361.450 15.680 369.650 ;
        RECT 16.130 361.450 16.280 369.650 ;
        RECT 16.730 361.450 16.880 369.650 ;
        RECT 17.330 361.450 17.480 369.650 ;
        RECT 17.930 361.450 18.080 369.650 ;
        RECT 18.530 361.450 18.680 369.650 ;
        RECT 19.130 369.200 19.430 369.650 ;
        RECT 19.130 369.050 22.980 369.200 ;
        RECT 19.130 368.600 19.430 369.050 ;
        RECT 19.130 368.450 22.980 368.600 ;
        RECT 19.130 368.000 19.430 368.450 ;
        RECT 19.130 367.850 22.980 368.000 ;
        RECT 19.130 367.400 19.430 367.850 ;
        RECT 19.130 367.250 22.980 367.400 ;
        RECT 19.130 366.800 19.430 367.250 ;
        RECT 23.830 366.800 25.630 373.200 ;
        RECT 30.030 372.750 30.330 373.200 ;
        RECT 26.480 372.600 30.330 372.750 ;
        RECT 30.030 372.150 30.330 372.600 ;
        RECT 26.480 372.000 30.330 372.150 ;
        RECT 30.030 371.550 30.330 372.000 ;
        RECT 26.480 371.400 30.330 371.550 ;
        RECT 30.030 370.950 30.330 371.400 ;
        RECT 26.480 370.800 30.330 370.950 ;
        RECT 30.030 370.350 30.330 370.800 ;
        RECT 30.780 370.350 30.930 378.550 ;
        RECT 31.380 370.350 31.530 378.550 ;
        RECT 31.980 370.350 32.130 378.550 ;
        RECT 32.580 370.350 32.730 378.550 ;
        RECT 33.180 370.350 33.330 378.550 ;
        RECT 33.780 370.350 33.930 378.550 ;
        RECT 30.030 369.200 30.330 369.650 ;
        RECT 26.480 369.050 30.330 369.200 ;
        RECT 30.030 368.600 30.330 369.050 ;
        RECT 26.480 368.450 30.330 368.600 ;
        RECT 30.030 368.000 30.330 368.450 ;
        RECT 26.480 367.850 30.330 368.000 ;
        RECT 30.030 367.400 30.330 367.850 ;
        RECT 26.480 367.250 30.330 367.400 ;
        RECT 30.030 366.800 30.330 367.250 ;
        RECT 19.130 366.650 22.980 366.800 ;
        RECT 26.480 366.650 30.330 366.800 ;
        RECT 19.130 366.200 19.430 366.650 ;
        RECT 30.030 366.200 30.330 366.650 ;
        RECT 19.130 366.050 22.980 366.200 ;
        RECT 26.480 366.050 30.330 366.200 ;
        RECT 19.130 365.600 19.430 366.050 ;
        RECT 30.030 365.600 30.330 366.050 ;
        RECT 19.130 365.450 22.980 365.600 ;
        RECT 26.480 365.450 30.330 365.600 ;
        RECT 19.130 365.000 19.430 365.450 ;
        RECT 30.030 365.000 30.330 365.450 ;
        RECT 19.130 364.850 22.980 365.000 ;
        RECT 26.480 364.850 30.330 365.000 ;
        RECT 19.130 364.400 19.430 364.850 ;
        RECT 30.030 364.400 30.330 364.850 ;
        RECT 19.130 364.250 22.980 364.400 ;
        RECT 26.480 364.250 30.330 364.400 ;
        RECT 19.130 363.800 19.430 364.250 ;
        RECT 30.030 363.800 30.330 364.250 ;
        RECT 19.130 363.650 22.980 363.800 ;
        RECT 26.480 363.650 30.330 363.800 ;
        RECT 19.130 363.200 19.430 363.650 ;
        RECT 30.030 363.200 30.330 363.650 ;
        RECT 19.130 363.050 22.980 363.200 ;
        RECT 26.480 363.050 30.330 363.200 ;
        RECT 19.130 362.600 19.430 363.050 ;
        RECT 30.030 362.600 30.330 363.050 ;
        RECT 19.130 362.450 22.980 362.600 ;
        RECT 26.480 362.450 30.330 362.600 ;
        RECT 19.130 362.000 19.430 362.450 ;
        RECT 30.030 362.000 30.330 362.450 ;
        RECT 19.130 361.450 22.930 362.000 ;
        RECT 6.530 361.400 22.930 361.450 ;
        RECT 26.530 361.450 30.330 362.000 ;
        RECT 30.780 361.450 30.930 369.650 ;
        RECT 31.380 361.450 31.530 369.650 ;
        RECT 31.980 361.450 32.130 369.650 ;
        RECT 32.580 361.450 32.730 369.650 ;
        RECT 33.180 361.450 33.330 369.650 ;
        RECT 33.780 361.450 33.930 369.650 ;
        RECT 34.380 361.450 35.080 378.550 ;
        RECT 35.530 370.350 35.680 378.550 ;
        RECT 36.130 370.350 36.280 378.550 ;
        RECT 36.730 370.350 36.880 378.550 ;
        RECT 37.330 370.350 37.480 378.550 ;
        RECT 37.930 370.350 38.080 378.550 ;
        RECT 38.530 370.350 38.680 378.550 ;
        RECT 39.130 378.000 42.930 378.550 ;
        RECT 46.530 378.550 62.930 378.600 ;
        RECT 46.530 378.000 50.330 378.550 ;
        RECT 39.130 377.550 39.430 378.000 ;
        RECT 50.030 377.550 50.330 378.000 ;
        RECT 39.130 377.400 42.980 377.550 ;
        RECT 46.480 377.400 50.330 377.550 ;
        RECT 39.130 376.950 39.430 377.400 ;
        RECT 50.030 376.950 50.330 377.400 ;
        RECT 39.130 376.800 42.980 376.950 ;
        RECT 46.480 376.800 50.330 376.950 ;
        RECT 39.130 376.350 39.430 376.800 ;
        RECT 50.030 376.350 50.330 376.800 ;
        RECT 39.130 376.200 42.980 376.350 ;
        RECT 46.480 376.200 50.330 376.350 ;
        RECT 39.130 375.750 39.430 376.200 ;
        RECT 50.030 375.750 50.330 376.200 ;
        RECT 39.130 375.600 42.980 375.750 ;
        RECT 46.480 375.600 50.330 375.750 ;
        RECT 39.130 375.150 39.430 375.600 ;
        RECT 50.030 375.150 50.330 375.600 ;
        RECT 39.130 375.000 42.980 375.150 ;
        RECT 46.480 375.000 50.330 375.150 ;
        RECT 39.130 374.550 39.430 375.000 ;
        RECT 50.030 374.550 50.330 375.000 ;
        RECT 39.130 374.400 42.980 374.550 ;
        RECT 46.480 374.400 50.330 374.550 ;
        RECT 39.130 373.950 39.430 374.400 ;
        RECT 50.030 373.950 50.330 374.400 ;
        RECT 39.130 373.800 42.980 373.950 ;
        RECT 46.480 373.800 50.330 373.950 ;
        RECT 39.130 373.350 39.430 373.800 ;
        RECT 50.030 373.350 50.330 373.800 ;
        RECT 39.130 373.200 42.980 373.350 ;
        RECT 46.480 373.200 50.330 373.350 ;
        RECT 39.130 372.750 39.430 373.200 ;
        RECT 39.130 372.600 42.980 372.750 ;
        RECT 39.130 372.150 39.430 372.600 ;
        RECT 39.130 372.000 42.980 372.150 ;
        RECT 39.130 371.550 39.430 372.000 ;
        RECT 39.130 371.400 42.980 371.550 ;
        RECT 39.130 370.950 39.430 371.400 ;
        RECT 39.130 370.800 42.980 370.950 ;
        RECT 39.130 370.350 39.430 370.800 ;
        RECT 35.530 361.450 35.680 369.650 ;
        RECT 36.130 361.450 36.280 369.650 ;
        RECT 36.730 361.450 36.880 369.650 ;
        RECT 37.330 361.450 37.480 369.650 ;
        RECT 37.930 361.450 38.080 369.650 ;
        RECT 38.530 361.450 38.680 369.650 ;
        RECT 39.130 369.200 39.430 369.650 ;
        RECT 39.130 369.050 42.980 369.200 ;
        RECT 39.130 368.600 39.430 369.050 ;
        RECT 39.130 368.450 42.980 368.600 ;
        RECT 39.130 368.000 39.430 368.450 ;
        RECT 39.130 367.850 42.980 368.000 ;
        RECT 39.130 367.400 39.430 367.850 ;
        RECT 39.130 367.250 42.980 367.400 ;
        RECT 39.130 366.800 39.430 367.250 ;
        RECT 43.830 366.800 45.630 373.200 ;
        RECT 50.030 372.750 50.330 373.200 ;
        RECT 46.480 372.600 50.330 372.750 ;
        RECT 50.030 372.150 50.330 372.600 ;
        RECT 46.480 372.000 50.330 372.150 ;
        RECT 50.030 371.550 50.330 372.000 ;
        RECT 46.480 371.400 50.330 371.550 ;
        RECT 50.030 370.950 50.330 371.400 ;
        RECT 46.480 370.800 50.330 370.950 ;
        RECT 50.030 370.350 50.330 370.800 ;
        RECT 50.780 370.350 50.930 378.550 ;
        RECT 51.380 370.350 51.530 378.550 ;
        RECT 51.980 370.350 52.130 378.550 ;
        RECT 52.580 370.350 52.730 378.550 ;
        RECT 53.180 370.350 53.330 378.550 ;
        RECT 53.780 370.350 53.930 378.550 ;
        RECT 50.030 369.200 50.330 369.650 ;
        RECT 46.480 369.050 50.330 369.200 ;
        RECT 50.030 368.600 50.330 369.050 ;
        RECT 46.480 368.450 50.330 368.600 ;
        RECT 50.030 368.000 50.330 368.450 ;
        RECT 46.480 367.850 50.330 368.000 ;
        RECT 50.030 367.400 50.330 367.850 ;
        RECT 46.480 367.250 50.330 367.400 ;
        RECT 50.030 366.800 50.330 367.250 ;
        RECT 39.130 366.650 42.980 366.800 ;
        RECT 46.480 366.650 50.330 366.800 ;
        RECT 39.130 366.200 39.430 366.650 ;
        RECT 50.030 366.200 50.330 366.650 ;
        RECT 39.130 366.050 42.980 366.200 ;
        RECT 46.480 366.050 50.330 366.200 ;
        RECT 39.130 365.600 39.430 366.050 ;
        RECT 50.030 365.600 50.330 366.050 ;
        RECT 39.130 365.450 42.980 365.600 ;
        RECT 46.480 365.450 50.330 365.600 ;
        RECT 39.130 365.000 39.430 365.450 ;
        RECT 50.030 365.000 50.330 365.450 ;
        RECT 39.130 364.850 42.980 365.000 ;
        RECT 46.480 364.850 50.330 365.000 ;
        RECT 39.130 364.400 39.430 364.850 ;
        RECT 50.030 364.400 50.330 364.850 ;
        RECT 39.130 364.250 42.980 364.400 ;
        RECT 46.480 364.250 50.330 364.400 ;
        RECT 39.130 363.800 39.430 364.250 ;
        RECT 50.030 363.800 50.330 364.250 ;
        RECT 39.130 363.650 42.980 363.800 ;
        RECT 46.480 363.650 50.330 363.800 ;
        RECT 39.130 363.200 39.430 363.650 ;
        RECT 50.030 363.200 50.330 363.650 ;
        RECT 39.130 363.050 42.980 363.200 ;
        RECT 46.480 363.050 50.330 363.200 ;
        RECT 39.130 362.600 39.430 363.050 ;
        RECT 50.030 362.600 50.330 363.050 ;
        RECT 39.130 362.450 42.980 362.600 ;
        RECT 46.480 362.450 50.330 362.600 ;
        RECT 39.130 362.000 39.430 362.450 ;
        RECT 50.030 362.000 50.330 362.450 ;
        RECT 39.130 361.450 42.930 362.000 ;
        RECT 26.530 361.400 42.930 361.450 ;
        RECT 46.530 361.450 50.330 362.000 ;
        RECT 50.780 361.450 50.930 369.650 ;
        RECT 51.380 361.450 51.530 369.650 ;
        RECT 51.980 361.450 52.130 369.650 ;
        RECT 52.580 361.450 52.730 369.650 ;
        RECT 53.180 361.450 53.330 369.650 ;
        RECT 53.780 361.450 53.930 369.650 ;
        RECT 54.380 361.450 55.080 378.550 ;
        RECT 55.530 370.350 55.680 378.550 ;
        RECT 56.130 370.350 56.280 378.550 ;
        RECT 56.730 370.350 56.880 378.550 ;
        RECT 57.330 370.350 57.480 378.550 ;
        RECT 57.930 370.350 58.080 378.550 ;
        RECT 58.530 370.350 58.680 378.550 ;
        RECT 59.130 378.000 62.930 378.550 ;
        RECT 66.530 378.550 82.930 378.600 ;
        RECT 66.530 378.000 70.330 378.550 ;
        RECT 59.130 377.550 59.430 378.000 ;
        RECT 70.030 377.550 70.330 378.000 ;
        RECT 59.130 377.400 62.980 377.550 ;
        RECT 66.480 377.400 70.330 377.550 ;
        RECT 59.130 376.950 59.430 377.400 ;
        RECT 70.030 376.950 70.330 377.400 ;
        RECT 59.130 376.800 62.980 376.950 ;
        RECT 66.480 376.800 70.330 376.950 ;
        RECT 59.130 376.350 59.430 376.800 ;
        RECT 70.030 376.350 70.330 376.800 ;
        RECT 59.130 376.200 62.980 376.350 ;
        RECT 66.480 376.200 70.330 376.350 ;
        RECT 59.130 375.750 59.430 376.200 ;
        RECT 70.030 375.750 70.330 376.200 ;
        RECT 59.130 375.600 62.980 375.750 ;
        RECT 66.480 375.600 70.330 375.750 ;
        RECT 59.130 375.150 59.430 375.600 ;
        RECT 70.030 375.150 70.330 375.600 ;
        RECT 59.130 375.000 62.980 375.150 ;
        RECT 66.480 375.000 70.330 375.150 ;
        RECT 59.130 374.550 59.430 375.000 ;
        RECT 70.030 374.550 70.330 375.000 ;
        RECT 59.130 374.400 62.980 374.550 ;
        RECT 66.480 374.400 70.330 374.550 ;
        RECT 59.130 373.950 59.430 374.400 ;
        RECT 70.030 373.950 70.330 374.400 ;
        RECT 59.130 373.800 62.980 373.950 ;
        RECT 66.480 373.800 70.330 373.950 ;
        RECT 59.130 373.350 59.430 373.800 ;
        RECT 70.030 373.350 70.330 373.800 ;
        RECT 59.130 373.200 62.980 373.350 ;
        RECT 66.480 373.200 70.330 373.350 ;
        RECT 59.130 372.750 59.430 373.200 ;
        RECT 59.130 372.600 62.980 372.750 ;
        RECT 59.130 372.150 59.430 372.600 ;
        RECT 59.130 372.000 62.980 372.150 ;
        RECT 59.130 371.550 59.430 372.000 ;
        RECT 59.130 371.400 62.980 371.550 ;
        RECT 59.130 370.950 59.430 371.400 ;
        RECT 59.130 370.800 62.980 370.950 ;
        RECT 59.130 370.350 59.430 370.800 ;
        RECT 55.530 361.450 55.680 369.650 ;
        RECT 56.130 361.450 56.280 369.650 ;
        RECT 56.730 361.450 56.880 369.650 ;
        RECT 57.330 361.450 57.480 369.650 ;
        RECT 57.930 361.450 58.080 369.650 ;
        RECT 58.530 361.450 58.680 369.650 ;
        RECT 59.130 369.200 59.430 369.650 ;
        RECT 59.130 369.050 62.980 369.200 ;
        RECT 59.130 368.600 59.430 369.050 ;
        RECT 59.130 368.450 62.980 368.600 ;
        RECT 59.130 368.000 59.430 368.450 ;
        RECT 59.130 367.850 62.980 368.000 ;
        RECT 59.130 367.400 59.430 367.850 ;
        RECT 59.130 367.250 62.980 367.400 ;
        RECT 59.130 366.800 59.430 367.250 ;
        RECT 63.830 366.800 65.630 373.200 ;
        RECT 70.030 372.750 70.330 373.200 ;
        RECT 66.480 372.600 70.330 372.750 ;
        RECT 70.030 372.150 70.330 372.600 ;
        RECT 66.480 372.000 70.330 372.150 ;
        RECT 70.030 371.550 70.330 372.000 ;
        RECT 66.480 371.400 70.330 371.550 ;
        RECT 70.030 370.950 70.330 371.400 ;
        RECT 66.480 370.800 70.330 370.950 ;
        RECT 70.030 370.350 70.330 370.800 ;
        RECT 70.780 370.350 70.930 378.550 ;
        RECT 71.380 370.350 71.530 378.550 ;
        RECT 71.980 370.350 72.130 378.550 ;
        RECT 72.580 370.350 72.730 378.550 ;
        RECT 73.180 370.350 73.330 378.550 ;
        RECT 73.780 370.350 73.930 378.550 ;
        RECT 70.030 369.200 70.330 369.650 ;
        RECT 66.480 369.050 70.330 369.200 ;
        RECT 70.030 368.600 70.330 369.050 ;
        RECT 66.480 368.450 70.330 368.600 ;
        RECT 70.030 368.000 70.330 368.450 ;
        RECT 66.480 367.850 70.330 368.000 ;
        RECT 70.030 367.400 70.330 367.850 ;
        RECT 66.480 367.250 70.330 367.400 ;
        RECT 70.030 366.800 70.330 367.250 ;
        RECT 59.130 366.650 62.980 366.800 ;
        RECT 66.480 366.650 70.330 366.800 ;
        RECT 59.130 366.200 59.430 366.650 ;
        RECT 70.030 366.200 70.330 366.650 ;
        RECT 59.130 366.050 62.980 366.200 ;
        RECT 66.480 366.050 70.330 366.200 ;
        RECT 59.130 365.600 59.430 366.050 ;
        RECT 70.030 365.600 70.330 366.050 ;
        RECT 59.130 365.450 62.980 365.600 ;
        RECT 66.480 365.450 70.330 365.600 ;
        RECT 59.130 365.000 59.430 365.450 ;
        RECT 70.030 365.000 70.330 365.450 ;
        RECT 59.130 364.850 62.980 365.000 ;
        RECT 66.480 364.850 70.330 365.000 ;
        RECT 59.130 364.400 59.430 364.850 ;
        RECT 70.030 364.400 70.330 364.850 ;
        RECT 59.130 364.250 62.980 364.400 ;
        RECT 66.480 364.250 70.330 364.400 ;
        RECT 59.130 363.800 59.430 364.250 ;
        RECT 70.030 363.800 70.330 364.250 ;
        RECT 59.130 363.650 62.980 363.800 ;
        RECT 66.480 363.650 70.330 363.800 ;
        RECT 59.130 363.200 59.430 363.650 ;
        RECT 70.030 363.200 70.330 363.650 ;
        RECT 59.130 363.050 62.980 363.200 ;
        RECT 66.480 363.050 70.330 363.200 ;
        RECT 59.130 362.600 59.430 363.050 ;
        RECT 70.030 362.600 70.330 363.050 ;
        RECT 59.130 362.450 62.980 362.600 ;
        RECT 66.480 362.450 70.330 362.600 ;
        RECT 59.130 362.000 59.430 362.450 ;
        RECT 70.030 362.000 70.330 362.450 ;
        RECT 59.130 361.450 62.930 362.000 ;
        RECT 46.530 361.400 62.930 361.450 ;
        RECT 66.530 361.450 70.330 362.000 ;
        RECT 70.780 361.450 70.930 369.650 ;
        RECT 71.380 361.450 71.530 369.650 ;
        RECT 71.980 361.450 72.130 369.650 ;
        RECT 72.580 361.450 72.730 369.650 ;
        RECT 73.180 361.450 73.330 369.650 ;
        RECT 73.780 361.450 73.930 369.650 ;
        RECT 74.380 361.450 75.080 378.550 ;
        RECT 75.530 370.350 75.680 378.550 ;
        RECT 76.130 370.350 76.280 378.550 ;
        RECT 76.730 370.350 76.880 378.550 ;
        RECT 77.330 370.350 77.480 378.550 ;
        RECT 77.930 370.350 78.080 378.550 ;
        RECT 78.530 370.350 78.680 378.550 ;
        RECT 79.130 378.000 82.930 378.550 ;
        RECT 86.530 378.550 102.930 378.600 ;
        RECT 86.530 378.000 90.330 378.550 ;
        RECT 79.130 377.550 79.430 378.000 ;
        RECT 90.030 377.550 90.330 378.000 ;
        RECT 79.130 377.400 82.980 377.550 ;
        RECT 86.480 377.400 90.330 377.550 ;
        RECT 79.130 376.950 79.430 377.400 ;
        RECT 90.030 376.950 90.330 377.400 ;
        RECT 79.130 376.800 82.980 376.950 ;
        RECT 86.480 376.800 90.330 376.950 ;
        RECT 79.130 376.350 79.430 376.800 ;
        RECT 90.030 376.350 90.330 376.800 ;
        RECT 79.130 376.200 82.980 376.350 ;
        RECT 86.480 376.200 90.330 376.350 ;
        RECT 79.130 375.750 79.430 376.200 ;
        RECT 90.030 375.750 90.330 376.200 ;
        RECT 79.130 375.600 82.980 375.750 ;
        RECT 86.480 375.600 90.330 375.750 ;
        RECT 79.130 375.150 79.430 375.600 ;
        RECT 90.030 375.150 90.330 375.600 ;
        RECT 79.130 375.000 82.980 375.150 ;
        RECT 86.480 375.000 90.330 375.150 ;
        RECT 79.130 374.550 79.430 375.000 ;
        RECT 90.030 374.550 90.330 375.000 ;
        RECT 79.130 374.400 82.980 374.550 ;
        RECT 86.480 374.400 90.330 374.550 ;
        RECT 79.130 373.950 79.430 374.400 ;
        RECT 90.030 373.950 90.330 374.400 ;
        RECT 79.130 373.800 82.980 373.950 ;
        RECT 86.480 373.800 90.330 373.950 ;
        RECT 79.130 373.350 79.430 373.800 ;
        RECT 90.030 373.350 90.330 373.800 ;
        RECT 79.130 373.200 82.980 373.350 ;
        RECT 86.480 373.200 90.330 373.350 ;
        RECT 79.130 372.750 79.430 373.200 ;
        RECT 79.130 372.600 82.980 372.750 ;
        RECT 79.130 372.150 79.430 372.600 ;
        RECT 79.130 372.000 82.980 372.150 ;
        RECT 79.130 371.550 79.430 372.000 ;
        RECT 79.130 371.400 82.980 371.550 ;
        RECT 79.130 370.950 79.430 371.400 ;
        RECT 79.130 370.800 82.980 370.950 ;
        RECT 79.130 370.350 79.430 370.800 ;
        RECT 75.530 361.450 75.680 369.650 ;
        RECT 76.130 361.450 76.280 369.650 ;
        RECT 76.730 361.450 76.880 369.650 ;
        RECT 77.330 361.450 77.480 369.650 ;
        RECT 77.930 361.450 78.080 369.650 ;
        RECT 78.530 361.450 78.680 369.650 ;
        RECT 79.130 369.200 79.430 369.650 ;
        RECT 79.130 369.050 82.980 369.200 ;
        RECT 79.130 368.600 79.430 369.050 ;
        RECT 79.130 368.450 82.980 368.600 ;
        RECT 79.130 368.000 79.430 368.450 ;
        RECT 79.130 367.850 82.980 368.000 ;
        RECT 79.130 367.400 79.430 367.850 ;
        RECT 79.130 367.250 82.980 367.400 ;
        RECT 79.130 366.800 79.430 367.250 ;
        RECT 83.830 366.800 85.630 373.200 ;
        RECT 90.030 372.750 90.330 373.200 ;
        RECT 86.480 372.600 90.330 372.750 ;
        RECT 90.030 372.150 90.330 372.600 ;
        RECT 86.480 372.000 90.330 372.150 ;
        RECT 90.030 371.550 90.330 372.000 ;
        RECT 86.480 371.400 90.330 371.550 ;
        RECT 90.030 370.950 90.330 371.400 ;
        RECT 86.480 370.800 90.330 370.950 ;
        RECT 90.030 370.350 90.330 370.800 ;
        RECT 90.780 370.350 90.930 378.550 ;
        RECT 91.380 370.350 91.530 378.550 ;
        RECT 91.980 370.350 92.130 378.550 ;
        RECT 92.580 370.350 92.730 378.550 ;
        RECT 93.180 370.350 93.330 378.550 ;
        RECT 93.780 370.350 93.930 378.550 ;
        RECT 90.030 369.200 90.330 369.650 ;
        RECT 86.480 369.050 90.330 369.200 ;
        RECT 90.030 368.600 90.330 369.050 ;
        RECT 86.480 368.450 90.330 368.600 ;
        RECT 90.030 368.000 90.330 368.450 ;
        RECT 86.480 367.850 90.330 368.000 ;
        RECT 90.030 367.400 90.330 367.850 ;
        RECT 86.480 367.250 90.330 367.400 ;
        RECT 90.030 366.800 90.330 367.250 ;
        RECT 79.130 366.650 82.980 366.800 ;
        RECT 86.480 366.650 90.330 366.800 ;
        RECT 79.130 366.200 79.430 366.650 ;
        RECT 90.030 366.200 90.330 366.650 ;
        RECT 79.130 366.050 82.980 366.200 ;
        RECT 86.480 366.050 90.330 366.200 ;
        RECT 79.130 365.600 79.430 366.050 ;
        RECT 90.030 365.600 90.330 366.050 ;
        RECT 79.130 365.450 82.980 365.600 ;
        RECT 86.480 365.450 90.330 365.600 ;
        RECT 79.130 365.000 79.430 365.450 ;
        RECT 90.030 365.000 90.330 365.450 ;
        RECT 79.130 364.850 82.980 365.000 ;
        RECT 86.480 364.850 90.330 365.000 ;
        RECT 79.130 364.400 79.430 364.850 ;
        RECT 90.030 364.400 90.330 364.850 ;
        RECT 79.130 364.250 82.980 364.400 ;
        RECT 86.480 364.250 90.330 364.400 ;
        RECT 79.130 363.800 79.430 364.250 ;
        RECT 90.030 363.800 90.330 364.250 ;
        RECT 79.130 363.650 82.980 363.800 ;
        RECT 86.480 363.650 90.330 363.800 ;
        RECT 79.130 363.200 79.430 363.650 ;
        RECT 90.030 363.200 90.330 363.650 ;
        RECT 79.130 363.050 82.980 363.200 ;
        RECT 86.480 363.050 90.330 363.200 ;
        RECT 79.130 362.600 79.430 363.050 ;
        RECT 90.030 362.600 90.330 363.050 ;
        RECT 79.130 362.450 82.980 362.600 ;
        RECT 86.480 362.450 90.330 362.600 ;
        RECT 79.130 362.000 79.430 362.450 ;
        RECT 90.030 362.000 90.330 362.450 ;
        RECT 79.130 361.450 82.930 362.000 ;
        RECT 66.530 361.400 82.930 361.450 ;
        RECT 86.530 361.450 90.330 362.000 ;
        RECT 90.780 361.450 90.930 369.650 ;
        RECT 91.380 361.450 91.530 369.650 ;
        RECT 91.980 361.450 92.130 369.650 ;
        RECT 92.580 361.450 92.730 369.650 ;
        RECT 93.180 361.450 93.330 369.650 ;
        RECT 93.780 361.450 93.930 369.650 ;
        RECT 94.380 361.450 95.080 378.550 ;
        RECT 95.530 370.350 95.680 378.550 ;
        RECT 96.130 370.350 96.280 378.550 ;
        RECT 96.730 370.350 96.880 378.550 ;
        RECT 97.330 370.350 97.480 378.550 ;
        RECT 97.930 370.350 98.080 378.550 ;
        RECT 98.530 370.350 98.680 378.550 ;
        RECT 99.130 378.000 102.930 378.550 ;
        RECT 99.130 377.550 99.430 378.000 ;
        RECT 99.130 377.400 102.980 377.550 ;
        RECT 99.130 376.950 99.430 377.400 ;
        RECT 99.130 376.800 102.980 376.950 ;
        RECT 99.130 376.350 99.430 376.800 ;
        RECT 99.130 376.200 102.980 376.350 ;
        RECT 99.130 375.750 99.430 376.200 ;
        RECT 99.130 375.600 102.980 375.750 ;
        RECT 99.130 375.150 99.430 375.600 ;
        RECT 99.130 375.000 102.980 375.150 ;
        RECT 99.130 374.550 99.430 375.000 ;
        RECT 99.130 374.400 102.980 374.550 ;
        RECT 99.130 373.950 99.430 374.400 ;
        RECT 99.130 373.800 102.980 373.950 ;
        RECT 99.130 373.350 99.430 373.800 ;
        RECT 99.130 373.200 102.980 373.350 ;
        RECT 99.130 372.750 99.430 373.200 ;
        RECT 99.130 372.600 102.980 372.750 ;
        RECT 99.130 372.150 99.430 372.600 ;
        RECT 99.130 372.000 102.980 372.150 ;
        RECT 99.130 371.550 99.430 372.000 ;
        RECT 99.130 371.400 102.980 371.550 ;
        RECT 99.130 370.950 99.430 371.400 ;
        RECT 99.130 370.800 102.980 370.950 ;
        RECT 99.130 370.350 99.430 370.800 ;
        RECT 95.530 361.450 95.680 369.650 ;
        RECT 96.130 361.450 96.280 369.650 ;
        RECT 96.730 361.450 96.880 369.650 ;
        RECT 97.330 361.450 97.480 369.650 ;
        RECT 97.930 361.450 98.080 369.650 ;
        RECT 98.530 361.450 98.680 369.650 ;
        RECT 99.130 369.200 99.430 369.650 ;
        RECT 99.130 369.050 102.980 369.200 ;
        RECT 99.130 368.600 99.430 369.050 ;
        RECT 99.130 368.450 102.980 368.600 ;
        RECT 99.130 368.000 99.430 368.450 ;
        RECT 99.130 367.850 102.980 368.000 ;
        RECT 99.130 367.400 99.430 367.850 ;
        RECT 99.130 367.250 102.980 367.400 ;
        RECT 99.130 366.800 99.430 367.250 ;
        RECT 103.830 366.800 104.730 373.200 ;
        RECT 109.850 369.205 111.850 370.480 ;
        RECT 99.130 366.650 102.980 366.800 ;
        RECT 99.130 366.200 99.430 366.650 ;
        RECT 99.130 366.050 102.980 366.200 ;
        RECT 99.130 365.600 99.430 366.050 ;
        RECT 99.130 365.450 102.980 365.600 ;
        RECT 99.130 365.000 99.430 365.450 ;
        RECT 99.130 364.850 102.980 365.000 ;
        RECT 99.130 364.400 99.430 364.850 ;
        RECT 99.130 364.250 102.980 364.400 ;
        RECT 99.130 363.800 99.430 364.250 ;
        RECT 99.130 363.650 102.980 363.800 ;
        RECT 99.130 363.200 99.430 363.650 ;
        RECT 99.130 363.050 102.980 363.200 ;
        RECT 99.130 362.600 99.430 363.050 ;
        RECT 99.130 362.450 102.980 362.600 ;
        RECT 99.130 362.000 99.430 362.450 ;
        RECT 99.130 361.450 102.930 362.000 ;
        RECT 86.530 361.400 102.930 361.450 ;
        RECT 9.630 360.900 19.830 361.400 ;
        RECT 29.630 360.900 39.830 361.400 ;
        RECT 49.630 360.900 59.830 361.400 ;
        RECT 69.630 360.900 79.830 361.400 ;
        RECT 89.630 360.900 99.830 361.400 ;
        RECT 11.530 359.100 17.930 360.900 ;
        RECT 31.530 359.100 37.930 360.900 ;
        RECT 51.530 359.100 57.930 360.900 ;
        RECT 71.530 359.100 77.930 360.900 ;
        RECT 91.530 359.100 97.930 360.900 ;
        RECT 9.630 358.600 19.830 359.100 ;
        RECT 29.630 358.600 39.830 359.100 ;
        RECT 49.630 358.600 59.830 359.100 ;
        RECT 69.630 358.600 79.830 359.100 ;
        RECT 89.630 358.600 99.830 359.100 ;
        RECT 6.530 358.550 22.930 358.600 ;
        RECT 6.530 358.000 10.330 358.550 ;
        RECT 10.030 357.550 10.330 358.000 ;
        RECT 6.480 357.400 10.330 357.550 ;
        RECT 10.030 356.950 10.330 357.400 ;
        RECT 6.480 356.800 10.330 356.950 ;
        RECT 10.030 356.350 10.330 356.800 ;
        RECT 6.480 356.200 10.330 356.350 ;
        RECT 10.030 355.750 10.330 356.200 ;
        RECT 6.480 355.600 10.330 355.750 ;
        RECT 10.030 355.150 10.330 355.600 ;
        RECT 6.480 355.000 10.330 355.150 ;
        RECT 10.030 354.550 10.330 355.000 ;
        RECT 6.480 354.400 10.330 354.550 ;
        RECT 10.030 353.950 10.330 354.400 ;
        RECT 6.480 353.800 10.330 353.950 ;
        RECT 10.030 353.350 10.330 353.800 ;
        RECT 6.480 353.200 10.330 353.350 ;
        RECT 4.730 346.800 5.630 353.200 ;
        RECT 10.030 352.750 10.330 353.200 ;
        RECT 6.480 352.600 10.330 352.750 ;
        RECT 10.030 352.150 10.330 352.600 ;
        RECT 6.480 352.000 10.330 352.150 ;
        RECT 10.030 351.550 10.330 352.000 ;
        RECT 6.480 351.400 10.330 351.550 ;
        RECT 10.030 350.950 10.330 351.400 ;
        RECT 6.480 350.800 10.330 350.950 ;
        RECT 10.030 350.350 10.330 350.800 ;
        RECT 10.780 350.350 10.930 358.550 ;
        RECT 11.380 350.350 11.530 358.550 ;
        RECT 11.980 350.350 12.130 358.550 ;
        RECT 12.580 350.350 12.730 358.550 ;
        RECT 13.180 350.350 13.330 358.550 ;
        RECT 13.780 350.350 13.930 358.550 ;
        RECT 10.030 349.200 10.330 349.650 ;
        RECT 6.480 349.050 10.330 349.200 ;
        RECT 10.030 348.600 10.330 349.050 ;
        RECT 6.480 348.450 10.330 348.600 ;
        RECT 10.030 348.000 10.330 348.450 ;
        RECT 6.480 347.850 10.330 348.000 ;
        RECT 10.030 347.400 10.330 347.850 ;
        RECT 6.480 347.250 10.330 347.400 ;
        RECT 10.030 346.800 10.330 347.250 ;
        RECT 6.480 346.650 10.330 346.800 ;
        RECT 10.030 346.200 10.330 346.650 ;
        RECT 6.480 346.050 10.330 346.200 ;
        RECT 10.030 345.600 10.330 346.050 ;
        RECT 6.480 345.450 10.330 345.600 ;
        RECT 10.030 345.000 10.330 345.450 ;
        RECT 6.480 344.850 10.330 345.000 ;
        RECT 10.030 344.400 10.330 344.850 ;
        RECT 6.480 344.250 10.330 344.400 ;
        RECT 10.030 343.800 10.330 344.250 ;
        RECT 6.480 343.650 10.330 343.800 ;
        RECT 10.030 343.200 10.330 343.650 ;
        RECT 6.480 343.050 10.330 343.200 ;
        RECT 10.030 342.600 10.330 343.050 ;
        RECT 6.480 342.450 10.330 342.600 ;
        RECT 10.030 342.000 10.330 342.450 ;
        RECT 6.530 341.450 10.330 342.000 ;
        RECT 10.780 341.450 10.930 349.650 ;
        RECT 11.380 341.450 11.530 349.650 ;
        RECT 11.980 341.450 12.130 349.650 ;
        RECT 12.580 341.450 12.730 349.650 ;
        RECT 13.180 341.450 13.330 349.650 ;
        RECT 13.780 341.450 13.930 349.650 ;
        RECT 14.380 341.450 15.080 358.550 ;
        RECT 15.530 350.350 15.680 358.550 ;
        RECT 16.130 350.350 16.280 358.550 ;
        RECT 16.730 350.350 16.880 358.550 ;
        RECT 17.330 350.350 17.480 358.550 ;
        RECT 17.930 350.350 18.080 358.550 ;
        RECT 18.530 350.350 18.680 358.550 ;
        RECT 19.130 358.000 22.930 358.550 ;
        RECT 26.530 358.550 42.930 358.600 ;
        RECT 26.530 358.000 30.330 358.550 ;
        RECT 19.130 357.550 19.430 358.000 ;
        RECT 30.030 357.550 30.330 358.000 ;
        RECT 19.130 357.400 22.980 357.550 ;
        RECT 26.480 357.400 30.330 357.550 ;
        RECT 19.130 356.950 19.430 357.400 ;
        RECT 30.030 356.950 30.330 357.400 ;
        RECT 19.130 356.800 22.980 356.950 ;
        RECT 26.480 356.800 30.330 356.950 ;
        RECT 19.130 356.350 19.430 356.800 ;
        RECT 30.030 356.350 30.330 356.800 ;
        RECT 19.130 356.200 22.980 356.350 ;
        RECT 26.480 356.200 30.330 356.350 ;
        RECT 19.130 355.750 19.430 356.200 ;
        RECT 30.030 355.750 30.330 356.200 ;
        RECT 19.130 355.600 22.980 355.750 ;
        RECT 26.480 355.600 30.330 355.750 ;
        RECT 19.130 355.150 19.430 355.600 ;
        RECT 30.030 355.150 30.330 355.600 ;
        RECT 19.130 355.000 22.980 355.150 ;
        RECT 26.480 355.000 30.330 355.150 ;
        RECT 19.130 354.550 19.430 355.000 ;
        RECT 30.030 354.550 30.330 355.000 ;
        RECT 19.130 354.400 22.980 354.550 ;
        RECT 26.480 354.400 30.330 354.550 ;
        RECT 19.130 353.950 19.430 354.400 ;
        RECT 30.030 353.950 30.330 354.400 ;
        RECT 19.130 353.800 22.980 353.950 ;
        RECT 26.480 353.800 30.330 353.950 ;
        RECT 19.130 353.350 19.430 353.800 ;
        RECT 30.030 353.350 30.330 353.800 ;
        RECT 19.130 353.200 22.980 353.350 ;
        RECT 26.480 353.200 30.330 353.350 ;
        RECT 19.130 352.750 19.430 353.200 ;
        RECT 19.130 352.600 22.980 352.750 ;
        RECT 19.130 352.150 19.430 352.600 ;
        RECT 19.130 352.000 22.980 352.150 ;
        RECT 19.130 351.550 19.430 352.000 ;
        RECT 19.130 351.400 22.980 351.550 ;
        RECT 19.130 350.950 19.430 351.400 ;
        RECT 19.130 350.800 22.980 350.950 ;
        RECT 19.130 350.350 19.430 350.800 ;
        RECT 15.530 341.450 15.680 349.650 ;
        RECT 16.130 341.450 16.280 349.650 ;
        RECT 16.730 341.450 16.880 349.650 ;
        RECT 17.330 341.450 17.480 349.650 ;
        RECT 17.930 341.450 18.080 349.650 ;
        RECT 18.530 341.450 18.680 349.650 ;
        RECT 19.130 349.200 19.430 349.650 ;
        RECT 19.130 349.050 22.980 349.200 ;
        RECT 19.130 348.600 19.430 349.050 ;
        RECT 19.130 348.450 22.980 348.600 ;
        RECT 19.130 348.000 19.430 348.450 ;
        RECT 19.130 347.850 22.980 348.000 ;
        RECT 19.130 347.400 19.430 347.850 ;
        RECT 19.130 347.250 22.980 347.400 ;
        RECT 19.130 346.800 19.430 347.250 ;
        RECT 23.830 346.800 25.630 353.200 ;
        RECT 30.030 352.750 30.330 353.200 ;
        RECT 26.480 352.600 30.330 352.750 ;
        RECT 30.030 352.150 30.330 352.600 ;
        RECT 26.480 352.000 30.330 352.150 ;
        RECT 30.030 351.550 30.330 352.000 ;
        RECT 26.480 351.400 30.330 351.550 ;
        RECT 30.030 350.950 30.330 351.400 ;
        RECT 26.480 350.800 30.330 350.950 ;
        RECT 30.030 350.350 30.330 350.800 ;
        RECT 30.780 350.350 30.930 358.550 ;
        RECT 31.380 350.350 31.530 358.550 ;
        RECT 31.980 350.350 32.130 358.550 ;
        RECT 32.580 350.350 32.730 358.550 ;
        RECT 33.180 350.350 33.330 358.550 ;
        RECT 33.780 350.350 33.930 358.550 ;
        RECT 30.030 349.200 30.330 349.650 ;
        RECT 26.480 349.050 30.330 349.200 ;
        RECT 30.030 348.600 30.330 349.050 ;
        RECT 26.480 348.450 30.330 348.600 ;
        RECT 30.030 348.000 30.330 348.450 ;
        RECT 26.480 347.850 30.330 348.000 ;
        RECT 30.030 347.400 30.330 347.850 ;
        RECT 26.480 347.250 30.330 347.400 ;
        RECT 30.030 346.800 30.330 347.250 ;
        RECT 19.130 346.650 22.980 346.800 ;
        RECT 26.480 346.650 30.330 346.800 ;
        RECT 19.130 346.200 19.430 346.650 ;
        RECT 30.030 346.200 30.330 346.650 ;
        RECT 19.130 346.050 22.980 346.200 ;
        RECT 26.480 346.050 30.330 346.200 ;
        RECT 19.130 345.600 19.430 346.050 ;
        RECT 30.030 345.600 30.330 346.050 ;
        RECT 19.130 345.450 22.980 345.600 ;
        RECT 26.480 345.450 30.330 345.600 ;
        RECT 19.130 345.000 19.430 345.450 ;
        RECT 30.030 345.000 30.330 345.450 ;
        RECT 19.130 344.850 22.980 345.000 ;
        RECT 26.480 344.850 30.330 345.000 ;
        RECT 19.130 344.400 19.430 344.850 ;
        RECT 30.030 344.400 30.330 344.850 ;
        RECT 19.130 344.250 22.980 344.400 ;
        RECT 26.480 344.250 30.330 344.400 ;
        RECT 19.130 343.800 19.430 344.250 ;
        RECT 30.030 343.800 30.330 344.250 ;
        RECT 19.130 343.650 22.980 343.800 ;
        RECT 26.480 343.650 30.330 343.800 ;
        RECT 19.130 343.200 19.430 343.650 ;
        RECT 30.030 343.200 30.330 343.650 ;
        RECT 19.130 343.050 22.980 343.200 ;
        RECT 26.480 343.050 30.330 343.200 ;
        RECT 19.130 342.600 19.430 343.050 ;
        RECT 30.030 342.600 30.330 343.050 ;
        RECT 19.130 342.450 22.980 342.600 ;
        RECT 26.480 342.450 30.330 342.600 ;
        RECT 19.130 342.000 19.430 342.450 ;
        RECT 30.030 342.000 30.330 342.450 ;
        RECT 19.130 341.450 22.930 342.000 ;
        RECT 6.530 341.400 22.930 341.450 ;
        RECT 26.530 341.450 30.330 342.000 ;
        RECT 30.780 341.450 30.930 349.650 ;
        RECT 31.380 341.450 31.530 349.650 ;
        RECT 31.980 341.450 32.130 349.650 ;
        RECT 32.580 341.450 32.730 349.650 ;
        RECT 33.180 341.450 33.330 349.650 ;
        RECT 33.780 341.450 33.930 349.650 ;
        RECT 34.380 341.450 35.080 358.550 ;
        RECT 35.530 350.350 35.680 358.550 ;
        RECT 36.130 350.350 36.280 358.550 ;
        RECT 36.730 350.350 36.880 358.550 ;
        RECT 37.330 350.350 37.480 358.550 ;
        RECT 37.930 350.350 38.080 358.550 ;
        RECT 38.530 350.350 38.680 358.550 ;
        RECT 39.130 358.000 42.930 358.550 ;
        RECT 46.530 358.550 62.930 358.600 ;
        RECT 46.530 358.000 50.330 358.550 ;
        RECT 39.130 357.550 39.430 358.000 ;
        RECT 50.030 357.550 50.330 358.000 ;
        RECT 39.130 357.400 42.980 357.550 ;
        RECT 46.480 357.400 50.330 357.550 ;
        RECT 39.130 356.950 39.430 357.400 ;
        RECT 50.030 356.950 50.330 357.400 ;
        RECT 39.130 356.800 42.980 356.950 ;
        RECT 46.480 356.800 50.330 356.950 ;
        RECT 39.130 356.350 39.430 356.800 ;
        RECT 50.030 356.350 50.330 356.800 ;
        RECT 39.130 356.200 42.980 356.350 ;
        RECT 46.480 356.200 50.330 356.350 ;
        RECT 39.130 355.750 39.430 356.200 ;
        RECT 50.030 355.750 50.330 356.200 ;
        RECT 39.130 355.600 42.980 355.750 ;
        RECT 46.480 355.600 50.330 355.750 ;
        RECT 39.130 355.150 39.430 355.600 ;
        RECT 50.030 355.150 50.330 355.600 ;
        RECT 39.130 355.000 42.980 355.150 ;
        RECT 46.480 355.000 50.330 355.150 ;
        RECT 39.130 354.550 39.430 355.000 ;
        RECT 50.030 354.550 50.330 355.000 ;
        RECT 39.130 354.400 42.980 354.550 ;
        RECT 46.480 354.400 50.330 354.550 ;
        RECT 39.130 353.950 39.430 354.400 ;
        RECT 50.030 353.950 50.330 354.400 ;
        RECT 39.130 353.800 42.980 353.950 ;
        RECT 46.480 353.800 50.330 353.950 ;
        RECT 39.130 353.350 39.430 353.800 ;
        RECT 50.030 353.350 50.330 353.800 ;
        RECT 39.130 353.200 42.980 353.350 ;
        RECT 46.480 353.200 50.330 353.350 ;
        RECT 39.130 352.750 39.430 353.200 ;
        RECT 39.130 352.600 42.980 352.750 ;
        RECT 39.130 352.150 39.430 352.600 ;
        RECT 39.130 352.000 42.980 352.150 ;
        RECT 39.130 351.550 39.430 352.000 ;
        RECT 39.130 351.400 42.980 351.550 ;
        RECT 39.130 350.950 39.430 351.400 ;
        RECT 39.130 350.800 42.980 350.950 ;
        RECT 39.130 350.350 39.430 350.800 ;
        RECT 35.530 341.450 35.680 349.650 ;
        RECT 36.130 341.450 36.280 349.650 ;
        RECT 36.730 341.450 36.880 349.650 ;
        RECT 37.330 341.450 37.480 349.650 ;
        RECT 37.930 341.450 38.080 349.650 ;
        RECT 38.530 341.450 38.680 349.650 ;
        RECT 39.130 349.200 39.430 349.650 ;
        RECT 39.130 349.050 42.980 349.200 ;
        RECT 39.130 348.600 39.430 349.050 ;
        RECT 39.130 348.450 42.980 348.600 ;
        RECT 39.130 348.000 39.430 348.450 ;
        RECT 39.130 347.850 42.980 348.000 ;
        RECT 39.130 347.400 39.430 347.850 ;
        RECT 39.130 347.250 42.980 347.400 ;
        RECT 39.130 346.800 39.430 347.250 ;
        RECT 43.830 346.800 45.630 353.200 ;
        RECT 50.030 352.750 50.330 353.200 ;
        RECT 46.480 352.600 50.330 352.750 ;
        RECT 50.030 352.150 50.330 352.600 ;
        RECT 46.480 352.000 50.330 352.150 ;
        RECT 50.030 351.550 50.330 352.000 ;
        RECT 46.480 351.400 50.330 351.550 ;
        RECT 50.030 350.950 50.330 351.400 ;
        RECT 46.480 350.800 50.330 350.950 ;
        RECT 50.030 350.350 50.330 350.800 ;
        RECT 50.780 350.350 50.930 358.550 ;
        RECT 51.380 350.350 51.530 358.550 ;
        RECT 51.980 350.350 52.130 358.550 ;
        RECT 52.580 350.350 52.730 358.550 ;
        RECT 53.180 350.350 53.330 358.550 ;
        RECT 53.780 350.350 53.930 358.550 ;
        RECT 50.030 349.200 50.330 349.650 ;
        RECT 46.480 349.050 50.330 349.200 ;
        RECT 50.030 348.600 50.330 349.050 ;
        RECT 46.480 348.450 50.330 348.600 ;
        RECT 50.030 348.000 50.330 348.450 ;
        RECT 46.480 347.850 50.330 348.000 ;
        RECT 50.030 347.400 50.330 347.850 ;
        RECT 46.480 347.250 50.330 347.400 ;
        RECT 50.030 346.800 50.330 347.250 ;
        RECT 39.130 346.650 42.980 346.800 ;
        RECT 46.480 346.650 50.330 346.800 ;
        RECT 39.130 346.200 39.430 346.650 ;
        RECT 50.030 346.200 50.330 346.650 ;
        RECT 39.130 346.050 42.980 346.200 ;
        RECT 46.480 346.050 50.330 346.200 ;
        RECT 39.130 345.600 39.430 346.050 ;
        RECT 50.030 345.600 50.330 346.050 ;
        RECT 39.130 345.450 42.980 345.600 ;
        RECT 46.480 345.450 50.330 345.600 ;
        RECT 39.130 345.000 39.430 345.450 ;
        RECT 50.030 345.000 50.330 345.450 ;
        RECT 39.130 344.850 42.980 345.000 ;
        RECT 46.480 344.850 50.330 345.000 ;
        RECT 39.130 344.400 39.430 344.850 ;
        RECT 50.030 344.400 50.330 344.850 ;
        RECT 39.130 344.250 42.980 344.400 ;
        RECT 46.480 344.250 50.330 344.400 ;
        RECT 39.130 343.800 39.430 344.250 ;
        RECT 50.030 343.800 50.330 344.250 ;
        RECT 39.130 343.650 42.980 343.800 ;
        RECT 46.480 343.650 50.330 343.800 ;
        RECT 39.130 343.200 39.430 343.650 ;
        RECT 50.030 343.200 50.330 343.650 ;
        RECT 39.130 343.050 42.980 343.200 ;
        RECT 46.480 343.050 50.330 343.200 ;
        RECT 39.130 342.600 39.430 343.050 ;
        RECT 50.030 342.600 50.330 343.050 ;
        RECT 39.130 342.450 42.980 342.600 ;
        RECT 46.480 342.450 50.330 342.600 ;
        RECT 39.130 342.000 39.430 342.450 ;
        RECT 50.030 342.000 50.330 342.450 ;
        RECT 39.130 341.450 42.930 342.000 ;
        RECT 26.530 341.400 42.930 341.450 ;
        RECT 46.530 341.450 50.330 342.000 ;
        RECT 50.780 341.450 50.930 349.650 ;
        RECT 51.380 341.450 51.530 349.650 ;
        RECT 51.980 341.450 52.130 349.650 ;
        RECT 52.580 341.450 52.730 349.650 ;
        RECT 53.180 341.450 53.330 349.650 ;
        RECT 53.780 341.450 53.930 349.650 ;
        RECT 54.380 341.450 55.080 358.550 ;
        RECT 55.530 350.350 55.680 358.550 ;
        RECT 56.130 350.350 56.280 358.550 ;
        RECT 56.730 350.350 56.880 358.550 ;
        RECT 57.330 350.350 57.480 358.550 ;
        RECT 57.930 350.350 58.080 358.550 ;
        RECT 58.530 350.350 58.680 358.550 ;
        RECT 59.130 358.000 62.930 358.550 ;
        RECT 66.530 358.550 82.930 358.600 ;
        RECT 66.530 358.000 70.330 358.550 ;
        RECT 59.130 357.550 59.430 358.000 ;
        RECT 70.030 357.550 70.330 358.000 ;
        RECT 59.130 357.400 62.980 357.550 ;
        RECT 66.480 357.400 70.330 357.550 ;
        RECT 59.130 356.950 59.430 357.400 ;
        RECT 70.030 356.950 70.330 357.400 ;
        RECT 59.130 356.800 62.980 356.950 ;
        RECT 66.480 356.800 70.330 356.950 ;
        RECT 59.130 356.350 59.430 356.800 ;
        RECT 70.030 356.350 70.330 356.800 ;
        RECT 59.130 356.200 62.980 356.350 ;
        RECT 66.480 356.200 70.330 356.350 ;
        RECT 59.130 355.750 59.430 356.200 ;
        RECT 70.030 355.750 70.330 356.200 ;
        RECT 59.130 355.600 62.980 355.750 ;
        RECT 66.480 355.600 70.330 355.750 ;
        RECT 59.130 355.150 59.430 355.600 ;
        RECT 70.030 355.150 70.330 355.600 ;
        RECT 59.130 355.000 62.980 355.150 ;
        RECT 66.480 355.000 70.330 355.150 ;
        RECT 59.130 354.550 59.430 355.000 ;
        RECT 70.030 354.550 70.330 355.000 ;
        RECT 59.130 354.400 62.980 354.550 ;
        RECT 66.480 354.400 70.330 354.550 ;
        RECT 59.130 353.950 59.430 354.400 ;
        RECT 70.030 353.950 70.330 354.400 ;
        RECT 59.130 353.800 62.980 353.950 ;
        RECT 66.480 353.800 70.330 353.950 ;
        RECT 59.130 353.350 59.430 353.800 ;
        RECT 70.030 353.350 70.330 353.800 ;
        RECT 59.130 353.200 62.980 353.350 ;
        RECT 66.480 353.200 70.330 353.350 ;
        RECT 59.130 352.750 59.430 353.200 ;
        RECT 59.130 352.600 62.980 352.750 ;
        RECT 59.130 352.150 59.430 352.600 ;
        RECT 59.130 352.000 62.980 352.150 ;
        RECT 59.130 351.550 59.430 352.000 ;
        RECT 59.130 351.400 62.980 351.550 ;
        RECT 59.130 350.950 59.430 351.400 ;
        RECT 59.130 350.800 62.980 350.950 ;
        RECT 59.130 350.350 59.430 350.800 ;
        RECT 55.530 341.450 55.680 349.650 ;
        RECT 56.130 341.450 56.280 349.650 ;
        RECT 56.730 341.450 56.880 349.650 ;
        RECT 57.330 341.450 57.480 349.650 ;
        RECT 57.930 341.450 58.080 349.650 ;
        RECT 58.530 341.450 58.680 349.650 ;
        RECT 59.130 349.200 59.430 349.650 ;
        RECT 59.130 349.050 62.980 349.200 ;
        RECT 59.130 348.600 59.430 349.050 ;
        RECT 59.130 348.450 62.980 348.600 ;
        RECT 59.130 348.000 59.430 348.450 ;
        RECT 59.130 347.850 62.980 348.000 ;
        RECT 59.130 347.400 59.430 347.850 ;
        RECT 59.130 347.250 62.980 347.400 ;
        RECT 59.130 346.800 59.430 347.250 ;
        RECT 63.830 346.800 65.630 353.200 ;
        RECT 70.030 352.750 70.330 353.200 ;
        RECT 66.480 352.600 70.330 352.750 ;
        RECT 70.030 352.150 70.330 352.600 ;
        RECT 66.480 352.000 70.330 352.150 ;
        RECT 70.030 351.550 70.330 352.000 ;
        RECT 66.480 351.400 70.330 351.550 ;
        RECT 70.030 350.950 70.330 351.400 ;
        RECT 66.480 350.800 70.330 350.950 ;
        RECT 70.030 350.350 70.330 350.800 ;
        RECT 70.780 350.350 70.930 358.550 ;
        RECT 71.380 350.350 71.530 358.550 ;
        RECT 71.980 350.350 72.130 358.550 ;
        RECT 72.580 350.350 72.730 358.550 ;
        RECT 73.180 350.350 73.330 358.550 ;
        RECT 73.780 350.350 73.930 358.550 ;
        RECT 70.030 349.200 70.330 349.650 ;
        RECT 66.480 349.050 70.330 349.200 ;
        RECT 70.030 348.600 70.330 349.050 ;
        RECT 66.480 348.450 70.330 348.600 ;
        RECT 70.030 348.000 70.330 348.450 ;
        RECT 66.480 347.850 70.330 348.000 ;
        RECT 70.030 347.400 70.330 347.850 ;
        RECT 66.480 347.250 70.330 347.400 ;
        RECT 70.030 346.800 70.330 347.250 ;
        RECT 59.130 346.650 62.980 346.800 ;
        RECT 66.480 346.650 70.330 346.800 ;
        RECT 59.130 346.200 59.430 346.650 ;
        RECT 70.030 346.200 70.330 346.650 ;
        RECT 59.130 346.050 62.980 346.200 ;
        RECT 66.480 346.050 70.330 346.200 ;
        RECT 59.130 345.600 59.430 346.050 ;
        RECT 70.030 345.600 70.330 346.050 ;
        RECT 59.130 345.450 62.980 345.600 ;
        RECT 66.480 345.450 70.330 345.600 ;
        RECT 59.130 345.000 59.430 345.450 ;
        RECT 70.030 345.000 70.330 345.450 ;
        RECT 59.130 344.850 62.980 345.000 ;
        RECT 66.480 344.850 70.330 345.000 ;
        RECT 59.130 344.400 59.430 344.850 ;
        RECT 70.030 344.400 70.330 344.850 ;
        RECT 59.130 344.250 62.980 344.400 ;
        RECT 66.480 344.250 70.330 344.400 ;
        RECT 59.130 343.800 59.430 344.250 ;
        RECT 70.030 343.800 70.330 344.250 ;
        RECT 59.130 343.650 62.980 343.800 ;
        RECT 66.480 343.650 70.330 343.800 ;
        RECT 59.130 343.200 59.430 343.650 ;
        RECT 70.030 343.200 70.330 343.650 ;
        RECT 59.130 343.050 62.980 343.200 ;
        RECT 66.480 343.050 70.330 343.200 ;
        RECT 59.130 342.600 59.430 343.050 ;
        RECT 70.030 342.600 70.330 343.050 ;
        RECT 59.130 342.450 62.980 342.600 ;
        RECT 66.480 342.450 70.330 342.600 ;
        RECT 59.130 342.000 59.430 342.450 ;
        RECT 70.030 342.000 70.330 342.450 ;
        RECT 59.130 341.450 62.930 342.000 ;
        RECT 46.530 341.400 62.930 341.450 ;
        RECT 66.530 341.450 70.330 342.000 ;
        RECT 70.780 341.450 70.930 349.650 ;
        RECT 71.380 341.450 71.530 349.650 ;
        RECT 71.980 341.450 72.130 349.650 ;
        RECT 72.580 341.450 72.730 349.650 ;
        RECT 73.180 341.450 73.330 349.650 ;
        RECT 73.780 341.450 73.930 349.650 ;
        RECT 74.380 341.450 75.080 358.550 ;
        RECT 75.530 350.350 75.680 358.550 ;
        RECT 76.130 350.350 76.280 358.550 ;
        RECT 76.730 350.350 76.880 358.550 ;
        RECT 77.330 350.350 77.480 358.550 ;
        RECT 77.930 350.350 78.080 358.550 ;
        RECT 78.530 350.350 78.680 358.550 ;
        RECT 79.130 358.000 82.930 358.550 ;
        RECT 86.530 358.550 102.930 358.600 ;
        RECT 86.530 358.000 90.330 358.550 ;
        RECT 79.130 357.550 79.430 358.000 ;
        RECT 90.030 357.550 90.330 358.000 ;
        RECT 79.130 357.400 82.980 357.550 ;
        RECT 86.480 357.400 90.330 357.550 ;
        RECT 79.130 356.950 79.430 357.400 ;
        RECT 90.030 356.950 90.330 357.400 ;
        RECT 79.130 356.800 82.980 356.950 ;
        RECT 86.480 356.800 90.330 356.950 ;
        RECT 79.130 356.350 79.430 356.800 ;
        RECT 90.030 356.350 90.330 356.800 ;
        RECT 79.130 356.200 82.980 356.350 ;
        RECT 86.480 356.200 90.330 356.350 ;
        RECT 79.130 355.750 79.430 356.200 ;
        RECT 90.030 355.750 90.330 356.200 ;
        RECT 79.130 355.600 82.980 355.750 ;
        RECT 86.480 355.600 90.330 355.750 ;
        RECT 79.130 355.150 79.430 355.600 ;
        RECT 90.030 355.150 90.330 355.600 ;
        RECT 79.130 355.000 82.980 355.150 ;
        RECT 86.480 355.000 90.330 355.150 ;
        RECT 79.130 354.550 79.430 355.000 ;
        RECT 90.030 354.550 90.330 355.000 ;
        RECT 79.130 354.400 82.980 354.550 ;
        RECT 86.480 354.400 90.330 354.550 ;
        RECT 79.130 353.950 79.430 354.400 ;
        RECT 90.030 353.950 90.330 354.400 ;
        RECT 79.130 353.800 82.980 353.950 ;
        RECT 86.480 353.800 90.330 353.950 ;
        RECT 79.130 353.350 79.430 353.800 ;
        RECT 90.030 353.350 90.330 353.800 ;
        RECT 79.130 353.200 82.980 353.350 ;
        RECT 86.480 353.200 90.330 353.350 ;
        RECT 79.130 352.750 79.430 353.200 ;
        RECT 79.130 352.600 82.980 352.750 ;
        RECT 79.130 352.150 79.430 352.600 ;
        RECT 79.130 352.000 82.980 352.150 ;
        RECT 79.130 351.550 79.430 352.000 ;
        RECT 79.130 351.400 82.980 351.550 ;
        RECT 79.130 350.950 79.430 351.400 ;
        RECT 79.130 350.800 82.980 350.950 ;
        RECT 79.130 350.350 79.430 350.800 ;
        RECT 75.530 341.450 75.680 349.650 ;
        RECT 76.130 341.450 76.280 349.650 ;
        RECT 76.730 341.450 76.880 349.650 ;
        RECT 77.330 341.450 77.480 349.650 ;
        RECT 77.930 341.450 78.080 349.650 ;
        RECT 78.530 341.450 78.680 349.650 ;
        RECT 79.130 349.200 79.430 349.650 ;
        RECT 79.130 349.050 82.980 349.200 ;
        RECT 79.130 348.600 79.430 349.050 ;
        RECT 79.130 348.450 82.980 348.600 ;
        RECT 79.130 348.000 79.430 348.450 ;
        RECT 79.130 347.850 82.980 348.000 ;
        RECT 79.130 347.400 79.430 347.850 ;
        RECT 79.130 347.250 82.980 347.400 ;
        RECT 79.130 346.800 79.430 347.250 ;
        RECT 83.830 346.800 85.630 353.200 ;
        RECT 90.030 352.750 90.330 353.200 ;
        RECT 86.480 352.600 90.330 352.750 ;
        RECT 90.030 352.150 90.330 352.600 ;
        RECT 86.480 352.000 90.330 352.150 ;
        RECT 90.030 351.550 90.330 352.000 ;
        RECT 86.480 351.400 90.330 351.550 ;
        RECT 90.030 350.950 90.330 351.400 ;
        RECT 86.480 350.800 90.330 350.950 ;
        RECT 90.030 350.350 90.330 350.800 ;
        RECT 90.780 350.350 90.930 358.550 ;
        RECT 91.380 350.350 91.530 358.550 ;
        RECT 91.980 350.350 92.130 358.550 ;
        RECT 92.580 350.350 92.730 358.550 ;
        RECT 93.180 350.350 93.330 358.550 ;
        RECT 93.780 350.350 93.930 358.550 ;
        RECT 90.030 349.200 90.330 349.650 ;
        RECT 86.480 349.050 90.330 349.200 ;
        RECT 90.030 348.600 90.330 349.050 ;
        RECT 86.480 348.450 90.330 348.600 ;
        RECT 90.030 348.000 90.330 348.450 ;
        RECT 86.480 347.850 90.330 348.000 ;
        RECT 90.030 347.400 90.330 347.850 ;
        RECT 86.480 347.250 90.330 347.400 ;
        RECT 90.030 346.800 90.330 347.250 ;
        RECT 79.130 346.650 82.980 346.800 ;
        RECT 86.480 346.650 90.330 346.800 ;
        RECT 79.130 346.200 79.430 346.650 ;
        RECT 90.030 346.200 90.330 346.650 ;
        RECT 79.130 346.050 82.980 346.200 ;
        RECT 86.480 346.050 90.330 346.200 ;
        RECT 79.130 345.600 79.430 346.050 ;
        RECT 90.030 345.600 90.330 346.050 ;
        RECT 79.130 345.450 82.980 345.600 ;
        RECT 86.480 345.450 90.330 345.600 ;
        RECT 79.130 345.000 79.430 345.450 ;
        RECT 90.030 345.000 90.330 345.450 ;
        RECT 79.130 344.850 82.980 345.000 ;
        RECT 86.480 344.850 90.330 345.000 ;
        RECT 79.130 344.400 79.430 344.850 ;
        RECT 90.030 344.400 90.330 344.850 ;
        RECT 79.130 344.250 82.980 344.400 ;
        RECT 86.480 344.250 90.330 344.400 ;
        RECT 79.130 343.800 79.430 344.250 ;
        RECT 90.030 343.800 90.330 344.250 ;
        RECT 79.130 343.650 82.980 343.800 ;
        RECT 86.480 343.650 90.330 343.800 ;
        RECT 79.130 343.200 79.430 343.650 ;
        RECT 90.030 343.200 90.330 343.650 ;
        RECT 79.130 343.050 82.980 343.200 ;
        RECT 86.480 343.050 90.330 343.200 ;
        RECT 79.130 342.600 79.430 343.050 ;
        RECT 90.030 342.600 90.330 343.050 ;
        RECT 79.130 342.450 82.980 342.600 ;
        RECT 86.480 342.450 90.330 342.600 ;
        RECT 79.130 342.000 79.430 342.450 ;
        RECT 90.030 342.000 90.330 342.450 ;
        RECT 79.130 341.450 82.930 342.000 ;
        RECT 66.530 341.400 82.930 341.450 ;
        RECT 86.530 341.450 90.330 342.000 ;
        RECT 90.780 341.450 90.930 349.650 ;
        RECT 91.380 341.450 91.530 349.650 ;
        RECT 91.980 341.450 92.130 349.650 ;
        RECT 92.580 341.450 92.730 349.650 ;
        RECT 93.180 341.450 93.330 349.650 ;
        RECT 93.780 341.450 93.930 349.650 ;
        RECT 94.380 341.450 95.080 358.550 ;
        RECT 95.530 350.350 95.680 358.550 ;
        RECT 96.130 350.350 96.280 358.550 ;
        RECT 96.730 350.350 96.880 358.550 ;
        RECT 97.330 350.350 97.480 358.550 ;
        RECT 97.930 350.350 98.080 358.550 ;
        RECT 98.530 350.350 98.680 358.550 ;
        RECT 99.130 358.000 102.930 358.550 ;
        RECT 99.130 357.550 99.430 358.000 ;
        RECT 99.130 357.400 102.980 357.550 ;
        RECT 99.130 356.950 99.430 357.400 ;
        RECT 99.130 356.800 102.980 356.950 ;
        RECT 99.130 356.350 99.430 356.800 ;
        RECT 99.130 356.200 102.980 356.350 ;
        RECT 99.130 355.750 99.430 356.200 ;
        RECT 99.130 355.600 102.980 355.750 ;
        RECT 99.130 355.150 99.430 355.600 ;
        RECT 99.130 355.000 102.980 355.150 ;
        RECT 99.130 354.550 99.430 355.000 ;
        RECT 99.130 354.400 102.980 354.550 ;
        RECT 99.130 353.950 99.430 354.400 ;
        RECT 99.130 353.800 102.980 353.950 ;
        RECT 99.130 353.350 99.430 353.800 ;
        RECT 99.130 353.200 102.980 353.350 ;
        RECT 99.130 352.750 99.430 353.200 ;
        RECT 99.130 352.600 102.980 352.750 ;
        RECT 99.130 352.150 99.430 352.600 ;
        RECT 99.130 352.000 102.980 352.150 ;
        RECT 99.130 351.550 99.430 352.000 ;
        RECT 99.130 351.400 102.980 351.550 ;
        RECT 99.130 350.950 99.430 351.400 ;
        RECT 99.130 350.800 102.980 350.950 ;
        RECT 99.130 350.350 99.430 350.800 ;
        RECT 95.530 341.450 95.680 349.650 ;
        RECT 96.130 341.450 96.280 349.650 ;
        RECT 96.730 341.450 96.880 349.650 ;
        RECT 97.330 341.450 97.480 349.650 ;
        RECT 97.930 341.450 98.080 349.650 ;
        RECT 98.530 341.450 98.680 349.650 ;
        RECT 99.130 349.200 99.430 349.650 ;
        RECT 99.130 349.050 102.980 349.200 ;
        RECT 99.130 348.600 99.430 349.050 ;
        RECT 99.130 348.450 102.980 348.600 ;
        RECT 99.130 348.000 99.430 348.450 ;
        RECT 99.130 347.850 102.980 348.000 ;
        RECT 99.130 347.400 99.430 347.850 ;
        RECT 99.130 347.250 102.980 347.400 ;
        RECT 99.130 346.800 99.430 347.250 ;
        RECT 103.830 346.800 104.730 353.200 ;
        RECT 109.850 349.205 111.850 350.480 ;
        RECT 99.130 346.650 102.980 346.800 ;
        RECT 99.130 346.200 99.430 346.650 ;
        RECT 99.130 346.050 102.980 346.200 ;
        RECT 99.130 345.600 99.430 346.050 ;
        RECT 99.130 345.450 102.980 345.600 ;
        RECT 99.130 345.000 99.430 345.450 ;
        RECT 99.130 344.850 102.980 345.000 ;
        RECT 99.130 344.400 99.430 344.850 ;
        RECT 99.130 344.250 102.980 344.400 ;
        RECT 99.130 343.800 99.430 344.250 ;
        RECT 99.130 343.650 102.980 343.800 ;
        RECT 99.130 343.200 99.430 343.650 ;
        RECT 99.130 343.050 102.980 343.200 ;
        RECT 99.130 342.600 99.430 343.050 ;
        RECT 99.130 342.450 102.980 342.600 ;
        RECT 99.130 342.000 99.430 342.450 ;
        RECT 99.130 341.450 102.930 342.000 ;
        RECT 86.530 341.400 102.930 341.450 ;
        RECT 9.630 340.900 19.830 341.400 ;
        RECT 29.630 340.900 39.830 341.400 ;
        RECT 49.630 340.900 59.830 341.400 ;
        RECT 69.630 340.900 79.830 341.400 ;
        RECT 89.630 340.900 99.830 341.400 ;
        RECT 11.530 339.100 17.930 340.900 ;
        RECT 31.530 339.100 37.930 340.900 ;
        RECT 51.530 339.100 57.930 340.900 ;
        RECT 71.530 339.100 77.930 340.900 ;
        RECT 91.530 339.100 97.930 340.900 ;
        RECT 9.630 338.600 19.830 339.100 ;
        RECT 29.630 338.600 39.830 339.100 ;
        RECT 49.630 338.600 59.830 339.100 ;
        RECT 69.630 338.600 79.830 339.100 ;
        RECT 89.630 338.600 99.830 339.100 ;
        RECT 6.530 338.550 22.930 338.600 ;
        RECT 6.530 338.000 10.330 338.550 ;
        RECT 10.030 337.550 10.330 338.000 ;
        RECT 6.480 337.400 10.330 337.550 ;
        RECT 10.030 336.950 10.330 337.400 ;
        RECT 6.480 336.800 10.330 336.950 ;
        RECT 10.030 336.350 10.330 336.800 ;
        RECT 6.480 336.200 10.330 336.350 ;
        RECT 10.030 335.750 10.330 336.200 ;
        RECT 6.480 335.600 10.330 335.750 ;
        RECT 10.030 335.150 10.330 335.600 ;
        RECT 6.480 335.000 10.330 335.150 ;
        RECT 10.030 334.550 10.330 335.000 ;
        RECT 6.480 334.400 10.330 334.550 ;
        RECT 10.030 333.950 10.330 334.400 ;
        RECT 6.480 333.800 10.330 333.950 ;
        RECT 10.030 333.350 10.330 333.800 ;
        RECT 6.480 333.200 10.330 333.350 ;
        RECT 4.730 326.800 5.630 333.200 ;
        RECT 10.030 332.750 10.330 333.200 ;
        RECT 6.480 332.600 10.330 332.750 ;
        RECT 10.030 332.150 10.330 332.600 ;
        RECT 6.480 332.000 10.330 332.150 ;
        RECT 10.030 331.550 10.330 332.000 ;
        RECT 6.480 331.400 10.330 331.550 ;
        RECT 10.030 330.950 10.330 331.400 ;
        RECT 6.480 330.800 10.330 330.950 ;
        RECT 10.030 330.350 10.330 330.800 ;
        RECT 10.780 330.350 10.930 338.550 ;
        RECT 11.380 330.350 11.530 338.550 ;
        RECT 11.980 330.350 12.130 338.550 ;
        RECT 12.580 330.350 12.730 338.550 ;
        RECT 13.180 330.350 13.330 338.550 ;
        RECT 13.780 330.350 13.930 338.550 ;
        RECT 10.030 329.200 10.330 329.650 ;
        RECT 6.480 329.050 10.330 329.200 ;
        RECT 10.030 328.600 10.330 329.050 ;
        RECT 6.480 328.450 10.330 328.600 ;
        RECT 10.030 328.000 10.330 328.450 ;
        RECT 6.480 327.850 10.330 328.000 ;
        RECT 10.030 327.400 10.330 327.850 ;
        RECT 6.480 327.250 10.330 327.400 ;
        RECT 10.030 326.800 10.330 327.250 ;
        RECT 6.480 326.650 10.330 326.800 ;
        RECT 10.030 326.200 10.330 326.650 ;
        RECT 6.480 326.050 10.330 326.200 ;
        RECT 10.030 325.600 10.330 326.050 ;
        RECT 6.480 325.450 10.330 325.600 ;
        RECT 10.030 325.000 10.330 325.450 ;
        RECT 6.480 324.850 10.330 325.000 ;
        RECT 10.030 324.400 10.330 324.850 ;
        RECT 6.480 324.250 10.330 324.400 ;
        RECT 10.030 323.800 10.330 324.250 ;
        RECT 6.480 323.650 10.330 323.800 ;
        RECT 10.030 323.200 10.330 323.650 ;
        RECT 6.480 323.050 10.330 323.200 ;
        RECT 10.030 322.600 10.330 323.050 ;
        RECT 6.480 322.450 10.330 322.600 ;
        RECT 10.030 322.000 10.330 322.450 ;
        RECT 6.530 321.450 10.330 322.000 ;
        RECT 10.780 321.450 10.930 329.650 ;
        RECT 11.380 321.450 11.530 329.650 ;
        RECT 11.980 321.450 12.130 329.650 ;
        RECT 12.580 321.450 12.730 329.650 ;
        RECT 13.180 321.450 13.330 329.650 ;
        RECT 13.780 321.450 13.930 329.650 ;
        RECT 14.380 321.450 15.080 338.550 ;
        RECT 15.530 330.350 15.680 338.550 ;
        RECT 16.130 330.350 16.280 338.550 ;
        RECT 16.730 330.350 16.880 338.550 ;
        RECT 17.330 330.350 17.480 338.550 ;
        RECT 17.930 330.350 18.080 338.550 ;
        RECT 18.530 330.350 18.680 338.550 ;
        RECT 19.130 338.000 22.930 338.550 ;
        RECT 26.530 338.550 42.930 338.600 ;
        RECT 26.530 338.000 30.330 338.550 ;
        RECT 19.130 337.550 19.430 338.000 ;
        RECT 30.030 337.550 30.330 338.000 ;
        RECT 19.130 337.400 22.980 337.550 ;
        RECT 26.480 337.400 30.330 337.550 ;
        RECT 19.130 336.950 19.430 337.400 ;
        RECT 30.030 336.950 30.330 337.400 ;
        RECT 19.130 336.800 22.980 336.950 ;
        RECT 26.480 336.800 30.330 336.950 ;
        RECT 19.130 336.350 19.430 336.800 ;
        RECT 30.030 336.350 30.330 336.800 ;
        RECT 19.130 336.200 22.980 336.350 ;
        RECT 26.480 336.200 30.330 336.350 ;
        RECT 19.130 335.750 19.430 336.200 ;
        RECT 30.030 335.750 30.330 336.200 ;
        RECT 19.130 335.600 22.980 335.750 ;
        RECT 26.480 335.600 30.330 335.750 ;
        RECT 19.130 335.150 19.430 335.600 ;
        RECT 30.030 335.150 30.330 335.600 ;
        RECT 19.130 335.000 22.980 335.150 ;
        RECT 26.480 335.000 30.330 335.150 ;
        RECT 19.130 334.550 19.430 335.000 ;
        RECT 30.030 334.550 30.330 335.000 ;
        RECT 19.130 334.400 22.980 334.550 ;
        RECT 26.480 334.400 30.330 334.550 ;
        RECT 19.130 333.950 19.430 334.400 ;
        RECT 30.030 333.950 30.330 334.400 ;
        RECT 19.130 333.800 22.980 333.950 ;
        RECT 26.480 333.800 30.330 333.950 ;
        RECT 19.130 333.350 19.430 333.800 ;
        RECT 30.030 333.350 30.330 333.800 ;
        RECT 19.130 333.200 22.980 333.350 ;
        RECT 26.480 333.200 30.330 333.350 ;
        RECT 19.130 332.750 19.430 333.200 ;
        RECT 19.130 332.600 22.980 332.750 ;
        RECT 19.130 332.150 19.430 332.600 ;
        RECT 19.130 332.000 22.980 332.150 ;
        RECT 19.130 331.550 19.430 332.000 ;
        RECT 19.130 331.400 22.980 331.550 ;
        RECT 19.130 330.950 19.430 331.400 ;
        RECT 19.130 330.800 22.980 330.950 ;
        RECT 19.130 330.350 19.430 330.800 ;
        RECT 15.530 321.450 15.680 329.650 ;
        RECT 16.130 321.450 16.280 329.650 ;
        RECT 16.730 321.450 16.880 329.650 ;
        RECT 17.330 321.450 17.480 329.650 ;
        RECT 17.930 321.450 18.080 329.650 ;
        RECT 18.530 321.450 18.680 329.650 ;
        RECT 19.130 329.200 19.430 329.650 ;
        RECT 19.130 329.050 22.980 329.200 ;
        RECT 19.130 328.600 19.430 329.050 ;
        RECT 19.130 328.450 22.980 328.600 ;
        RECT 19.130 328.000 19.430 328.450 ;
        RECT 19.130 327.850 22.980 328.000 ;
        RECT 19.130 327.400 19.430 327.850 ;
        RECT 19.130 327.250 22.980 327.400 ;
        RECT 19.130 326.800 19.430 327.250 ;
        RECT 23.830 326.800 25.630 333.200 ;
        RECT 30.030 332.750 30.330 333.200 ;
        RECT 26.480 332.600 30.330 332.750 ;
        RECT 30.030 332.150 30.330 332.600 ;
        RECT 26.480 332.000 30.330 332.150 ;
        RECT 30.030 331.550 30.330 332.000 ;
        RECT 26.480 331.400 30.330 331.550 ;
        RECT 30.030 330.950 30.330 331.400 ;
        RECT 26.480 330.800 30.330 330.950 ;
        RECT 30.030 330.350 30.330 330.800 ;
        RECT 30.780 330.350 30.930 338.550 ;
        RECT 31.380 330.350 31.530 338.550 ;
        RECT 31.980 330.350 32.130 338.550 ;
        RECT 32.580 330.350 32.730 338.550 ;
        RECT 33.180 330.350 33.330 338.550 ;
        RECT 33.780 330.350 33.930 338.550 ;
        RECT 30.030 329.200 30.330 329.650 ;
        RECT 26.480 329.050 30.330 329.200 ;
        RECT 30.030 328.600 30.330 329.050 ;
        RECT 26.480 328.450 30.330 328.600 ;
        RECT 30.030 328.000 30.330 328.450 ;
        RECT 26.480 327.850 30.330 328.000 ;
        RECT 30.030 327.400 30.330 327.850 ;
        RECT 26.480 327.250 30.330 327.400 ;
        RECT 30.030 326.800 30.330 327.250 ;
        RECT 19.130 326.650 22.980 326.800 ;
        RECT 26.480 326.650 30.330 326.800 ;
        RECT 19.130 326.200 19.430 326.650 ;
        RECT 30.030 326.200 30.330 326.650 ;
        RECT 19.130 326.050 22.980 326.200 ;
        RECT 26.480 326.050 30.330 326.200 ;
        RECT 19.130 325.600 19.430 326.050 ;
        RECT 30.030 325.600 30.330 326.050 ;
        RECT 19.130 325.450 22.980 325.600 ;
        RECT 26.480 325.450 30.330 325.600 ;
        RECT 19.130 325.000 19.430 325.450 ;
        RECT 30.030 325.000 30.330 325.450 ;
        RECT 19.130 324.850 22.980 325.000 ;
        RECT 26.480 324.850 30.330 325.000 ;
        RECT 19.130 324.400 19.430 324.850 ;
        RECT 30.030 324.400 30.330 324.850 ;
        RECT 19.130 324.250 22.980 324.400 ;
        RECT 26.480 324.250 30.330 324.400 ;
        RECT 19.130 323.800 19.430 324.250 ;
        RECT 30.030 323.800 30.330 324.250 ;
        RECT 19.130 323.650 22.980 323.800 ;
        RECT 26.480 323.650 30.330 323.800 ;
        RECT 19.130 323.200 19.430 323.650 ;
        RECT 30.030 323.200 30.330 323.650 ;
        RECT 19.130 323.050 22.980 323.200 ;
        RECT 26.480 323.050 30.330 323.200 ;
        RECT 19.130 322.600 19.430 323.050 ;
        RECT 30.030 322.600 30.330 323.050 ;
        RECT 19.130 322.450 22.980 322.600 ;
        RECT 26.480 322.450 30.330 322.600 ;
        RECT 19.130 322.000 19.430 322.450 ;
        RECT 30.030 322.000 30.330 322.450 ;
        RECT 19.130 321.450 22.930 322.000 ;
        RECT 6.530 321.400 22.930 321.450 ;
        RECT 26.530 321.450 30.330 322.000 ;
        RECT 30.780 321.450 30.930 329.650 ;
        RECT 31.380 321.450 31.530 329.650 ;
        RECT 31.980 321.450 32.130 329.650 ;
        RECT 32.580 321.450 32.730 329.650 ;
        RECT 33.180 321.450 33.330 329.650 ;
        RECT 33.780 321.450 33.930 329.650 ;
        RECT 34.380 321.450 35.080 338.550 ;
        RECT 35.530 330.350 35.680 338.550 ;
        RECT 36.130 330.350 36.280 338.550 ;
        RECT 36.730 330.350 36.880 338.550 ;
        RECT 37.330 330.350 37.480 338.550 ;
        RECT 37.930 330.350 38.080 338.550 ;
        RECT 38.530 330.350 38.680 338.550 ;
        RECT 39.130 338.000 42.930 338.550 ;
        RECT 46.530 338.550 62.930 338.600 ;
        RECT 46.530 338.000 50.330 338.550 ;
        RECT 39.130 337.550 39.430 338.000 ;
        RECT 50.030 337.550 50.330 338.000 ;
        RECT 39.130 337.400 42.980 337.550 ;
        RECT 46.480 337.400 50.330 337.550 ;
        RECT 39.130 336.950 39.430 337.400 ;
        RECT 50.030 336.950 50.330 337.400 ;
        RECT 39.130 336.800 42.980 336.950 ;
        RECT 46.480 336.800 50.330 336.950 ;
        RECT 39.130 336.350 39.430 336.800 ;
        RECT 50.030 336.350 50.330 336.800 ;
        RECT 39.130 336.200 42.980 336.350 ;
        RECT 46.480 336.200 50.330 336.350 ;
        RECT 39.130 335.750 39.430 336.200 ;
        RECT 50.030 335.750 50.330 336.200 ;
        RECT 39.130 335.600 42.980 335.750 ;
        RECT 46.480 335.600 50.330 335.750 ;
        RECT 39.130 335.150 39.430 335.600 ;
        RECT 50.030 335.150 50.330 335.600 ;
        RECT 39.130 335.000 42.980 335.150 ;
        RECT 46.480 335.000 50.330 335.150 ;
        RECT 39.130 334.550 39.430 335.000 ;
        RECT 50.030 334.550 50.330 335.000 ;
        RECT 39.130 334.400 42.980 334.550 ;
        RECT 46.480 334.400 50.330 334.550 ;
        RECT 39.130 333.950 39.430 334.400 ;
        RECT 50.030 333.950 50.330 334.400 ;
        RECT 39.130 333.800 42.980 333.950 ;
        RECT 46.480 333.800 50.330 333.950 ;
        RECT 39.130 333.350 39.430 333.800 ;
        RECT 50.030 333.350 50.330 333.800 ;
        RECT 39.130 333.200 42.980 333.350 ;
        RECT 46.480 333.200 50.330 333.350 ;
        RECT 39.130 332.750 39.430 333.200 ;
        RECT 39.130 332.600 42.980 332.750 ;
        RECT 39.130 332.150 39.430 332.600 ;
        RECT 39.130 332.000 42.980 332.150 ;
        RECT 39.130 331.550 39.430 332.000 ;
        RECT 39.130 331.400 42.980 331.550 ;
        RECT 39.130 330.950 39.430 331.400 ;
        RECT 39.130 330.800 42.980 330.950 ;
        RECT 39.130 330.350 39.430 330.800 ;
        RECT 35.530 321.450 35.680 329.650 ;
        RECT 36.130 321.450 36.280 329.650 ;
        RECT 36.730 321.450 36.880 329.650 ;
        RECT 37.330 321.450 37.480 329.650 ;
        RECT 37.930 321.450 38.080 329.650 ;
        RECT 38.530 321.450 38.680 329.650 ;
        RECT 39.130 329.200 39.430 329.650 ;
        RECT 39.130 329.050 42.980 329.200 ;
        RECT 39.130 328.600 39.430 329.050 ;
        RECT 39.130 328.450 42.980 328.600 ;
        RECT 39.130 328.000 39.430 328.450 ;
        RECT 39.130 327.850 42.980 328.000 ;
        RECT 39.130 327.400 39.430 327.850 ;
        RECT 39.130 327.250 42.980 327.400 ;
        RECT 39.130 326.800 39.430 327.250 ;
        RECT 43.830 326.800 45.630 333.200 ;
        RECT 50.030 332.750 50.330 333.200 ;
        RECT 46.480 332.600 50.330 332.750 ;
        RECT 50.030 332.150 50.330 332.600 ;
        RECT 46.480 332.000 50.330 332.150 ;
        RECT 50.030 331.550 50.330 332.000 ;
        RECT 46.480 331.400 50.330 331.550 ;
        RECT 50.030 330.950 50.330 331.400 ;
        RECT 46.480 330.800 50.330 330.950 ;
        RECT 50.030 330.350 50.330 330.800 ;
        RECT 50.780 330.350 50.930 338.550 ;
        RECT 51.380 330.350 51.530 338.550 ;
        RECT 51.980 330.350 52.130 338.550 ;
        RECT 52.580 330.350 52.730 338.550 ;
        RECT 53.180 330.350 53.330 338.550 ;
        RECT 53.780 330.350 53.930 338.550 ;
        RECT 50.030 329.200 50.330 329.650 ;
        RECT 46.480 329.050 50.330 329.200 ;
        RECT 50.030 328.600 50.330 329.050 ;
        RECT 46.480 328.450 50.330 328.600 ;
        RECT 50.030 328.000 50.330 328.450 ;
        RECT 46.480 327.850 50.330 328.000 ;
        RECT 50.030 327.400 50.330 327.850 ;
        RECT 46.480 327.250 50.330 327.400 ;
        RECT 50.030 326.800 50.330 327.250 ;
        RECT 39.130 326.650 42.980 326.800 ;
        RECT 46.480 326.650 50.330 326.800 ;
        RECT 39.130 326.200 39.430 326.650 ;
        RECT 50.030 326.200 50.330 326.650 ;
        RECT 39.130 326.050 42.980 326.200 ;
        RECT 46.480 326.050 50.330 326.200 ;
        RECT 39.130 325.600 39.430 326.050 ;
        RECT 50.030 325.600 50.330 326.050 ;
        RECT 39.130 325.450 42.980 325.600 ;
        RECT 46.480 325.450 50.330 325.600 ;
        RECT 39.130 325.000 39.430 325.450 ;
        RECT 50.030 325.000 50.330 325.450 ;
        RECT 39.130 324.850 42.980 325.000 ;
        RECT 46.480 324.850 50.330 325.000 ;
        RECT 39.130 324.400 39.430 324.850 ;
        RECT 50.030 324.400 50.330 324.850 ;
        RECT 39.130 324.250 42.980 324.400 ;
        RECT 46.480 324.250 50.330 324.400 ;
        RECT 39.130 323.800 39.430 324.250 ;
        RECT 50.030 323.800 50.330 324.250 ;
        RECT 39.130 323.650 42.980 323.800 ;
        RECT 46.480 323.650 50.330 323.800 ;
        RECT 39.130 323.200 39.430 323.650 ;
        RECT 50.030 323.200 50.330 323.650 ;
        RECT 39.130 323.050 42.980 323.200 ;
        RECT 46.480 323.050 50.330 323.200 ;
        RECT 39.130 322.600 39.430 323.050 ;
        RECT 50.030 322.600 50.330 323.050 ;
        RECT 39.130 322.450 42.980 322.600 ;
        RECT 46.480 322.450 50.330 322.600 ;
        RECT 39.130 322.000 39.430 322.450 ;
        RECT 50.030 322.000 50.330 322.450 ;
        RECT 39.130 321.450 42.930 322.000 ;
        RECT 26.530 321.400 42.930 321.450 ;
        RECT 46.530 321.450 50.330 322.000 ;
        RECT 50.780 321.450 50.930 329.650 ;
        RECT 51.380 321.450 51.530 329.650 ;
        RECT 51.980 321.450 52.130 329.650 ;
        RECT 52.580 321.450 52.730 329.650 ;
        RECT 53.180 321.450 53.330 329.650 ;
        RECT 53.780 321.450 53.930 329.650 ;
        RECT 54.380 321.450 55.080 338.550 ;
        RECT 55.530 330.350 55.680 338.550 ;
        RECT 56.130 330.350 56.280 338.550 ;
        RECT 56.730 330.350 56.880 338.550 ;
        RECT 57.330 330.350 57.480 338.550 ;
        RECT 57.930 330.350 58.080 338.550 ;
        RECT 58.530 330.350 58.680 338.550 ;
        RECT 59.130 338.000 62.930 338.550 ;
        RECT 66.530 338.550 82.930 338.600 ;
        RECT 66.530 338.000 70.330 338.550 ;
        RECT 59.130 337.550 59.430 338.000 ;
        RECT 70.030 337.550 70.330 338.000 ;
        RECT 59.130 337.400 62.980 337.550 ;
        RECT 66.480 337.400 70.330 337.550 ;
        RECT 59.130 336.950 59.430 337.400 ;
        RECT 70.030 336.950 70.330 337.400 ;
        RECT 59.130 336.800 62.980 336.950 ;
        RECT 66.480 336.800 70.330 336.950 ;
        RECT 59.130 336.350 59.430 336.800 ;
        RECT 70.030 336.350 70.330 336.800 ;
        RECT 59.130 336.200 62.980 336.350 ;
        RECT 66.480 336.200 70.330 336.350 ;
        RECT 59.130 335.750 59.430 336.200 ;
        RECT 70.030 335.750 70.330 336.200 ;
        RECT 59.130 335.600 62.980 335.750 ;
        RECT 66.480 335.600 70.330 335.750 ;
        RECT 59.130 335.150 59.430 335.600 ;
        RECT 70.030 335.150 70.330 335.600 ;
        RECT 59.130 335.000 62.980 335.150 ;
        RECT 66.480 335.000 70.330 335.150 ;
        RECT 59.130 334.550 59.430 335.000 ;
        RECT 70.030 334.550 70.330 335.000 ;
        RECT 59.130 334.400 62.980 334.550 ;
        RECT 66.480 334.400 70.330 334.550 ;
        RECT 59.130 333.950 59.430 334.400 ;
        RECT 70.030 333.950 70.330 334.400 ;
        RECT 59.130 333.800 62.980 333.950 ;
        RECT 66.480 333.800 70.330 333.950 ;
        RECT 59.130 333.350 59.430 333.800 ;
        RECT 70.030 333.350 70.330 333.800 ;
        RECT 59.130 333.200 62.980 333.350 ;
        RECT 66.480 333.200 70.330 333.350 ;
        RECT 59.130 332.750 59.430 333.200 ;
        RECT 59.130 332.600 62.980 332.750 ;
        RECT 59.130 332.150 59.430 332.600 ;
        RECT 59.130 332.000 62.980 332.150 ;
        RECT 59.130 331.550 59.430 332.000 ;
        RECT 59.130 331.400 62.980 331.550 ;
        RECT 59.130 330.950 59.430 331.400 ;
        RECT 59.130 330.800 62.980 330.950 ;
        RECT 59.130 330.350 59.430 330.800 ;
        RECT 55.530 321.450 55.680 329.650 ;
        RECT 56.130 321.450 56.280 329.650 ;
        RECT 56.730 321.450 56.880 329.650 ;
        RECT 57.330 321.450 57.480 329.650 ;
        RECT 57.930 321.450 58.080 329.650 ;
        RECT 58.530 321.450 58.680 329.650 ;
        RECT 59.130 329.200 59.430 329.650 ;
        RECT 59.130 329.050 62.980 329.200 ;
        RECT 59.130 328.600 59.430 329.050 ;
        RECT 59.130 328.450 62.980 328.600 ;
        RECT 59.130 328.000 59.430 328.450 ;
        RECT 59.130 327.850 62.980 328.000 ;
        RECT 59.130 327.400 59.430 327.850 ;
        RECT 59.130 327.250 62.980 327.400 ;
        RECT 59.130 326.800 59.430 327.250 ;
        RECT 63.830 326.800 65.630 333.200 ;
        RECT 70.030 332.750 70.330 333.200 ;
        RECT 66.480 332.600 70.330 332.750 ;
        RECT 70.030 332.150 70.330 332.600 ;
        RECT 66.480 332.000 70.330 332.150 ;
        RECT 70.030 331.550 70.330 332.000 ;
        RECT 66.480 331.400 70.330 331.550 ;
        RECT 70.030 330.950 70.330 331.400 ;
        RECT 66.480 330.800 70.330 330.950 ;
        RECT 70.030 330.350 70.330 330.800 ;
        RECT 70.780 330.350 70.930 338.550 ;
        RECT 71.380 330.350 71.530 338.550 ;
        RECT 71.980 330.350 72.130 338.550 ;
        RECT 72.580 330.350 72.730 338.550 ;
        RECT 73.180 330.350 73.330 338.550 ;
        RECT 73.780 330.350 73.930 338.550 ;
        RECT 70.030 329.200 70.330 329.650 ;
        RECT 66.480 329.050 70.330 329.200 ;
        RECT 70.030 328.600 70.330 329.050 ;
        RECT 66.480 328.450 70.330 328.600 ;
        RECT 70.030 328.000 70.330 328.450 ;
        RECT 66.480 327.850 70.330 328.000 ;
        RECT 70.030 327.400 70.330 327.850 ;
        RECT 66.480 327.250 70.330 327.400 ;
        RECT 70.030 326.800 70.330 327.250 ;
        RECT 59.130 326.650 62.980 326.800 ;
        RECT 66.480 326.650 70.330 326.800 ;
        RECT 59.130 326.200 59.430 326.650 ;
        RECT 70.030 326.200 70.330 326.650 ;
        RECT 59.130 326.050 62.980 326.200 ;
        RECT 66.480 326.050 70.330 326.200 ;
        RECT 59.130 325.600 59.430 326.050 ;
        RECT 70.030 325.600 70.330 326.050 ;
        RECT 59.130 325.450 62.980 325.600 ;
        RECT 66.480 325.450 70.330 325.600 ;
        RECT 59.130 325.000 59.430 325.450 ;
        RECT 70.030 325.000 70.330 325.450 ;
        RECT 59.130 324.850 62.980 325.000 ;
        RECT 66.480 324.850 70.330 325.000 ;
        RECT 59.130 324.400 59.430 324.850 ;
        RECT 70.030 324.400 70.330 324.850 ;
        RECT 59.130 324.250 62.980 324.400 ;
        RECT 66.480 324.250 70.330 324.400 ;
        RECT 59.130 323.800 59.430 324.250 ;
        RECT 70.030 323.800 70.330 324.250 ;
        RECT 59.130 323.650 62.980 323.800 ;
        RECT 66.480 323.650 70.330 323.800 ;
        RECT 59.130 323.200 59.430 323.650 ;
        RECT 70.030 323.200 70.330 323.650 ;
        RECT 59.130 323.050 62.980 323.200 ;
        RECT 66.480 323.050 70.330 323.200 ;
        RECT 59.130 322.600 59.430 323.050 ;
        RECT 70.030 322.600 70.330 323.050 ;
        RECT 59.130 322.450 62.980 322.600 ;
        RECT 66.480 322.450 70.330 322.600 ;
        RECT 59.130 322.000 59.430 322.450 ;
        RECT 70.030 322.000 70.330 322.450 ;
        RECT 59.130 321.450 62.930 322.000 ;
        RECT 46.530 321.400 62.930 321.450 ;
        RECT 66.530 321.450 70.330 322.000 ;
        RECT 70.780 321.450 70.930 329.650 ;
        RECT 71.380 321.450 71.530 329.650 ;
        RECT 71.980 321.450 72.130 329.650 ;
        RECT 72.580 321.450 72.730 329.650 ;
        RECT 73.180 321.450 73.330 329.650 ;
        RECT 73.780 321.450 73.930 329.650 ;
        RECT 74.380 321.450 75.080 338.550 ;
        RECT 75.530 330.350 75.680 338.550 ;
        RECT 76.130 330.350 76.280 338.550 ;
        RECT 76.730 330.350 76.880 338.550 ;
        RECT 77.330 330.350 77.480 338.550 ;
        RECT 77.930 330.350 78.080 338.550 ;
        RECT 78.530 330.350 78.680 338.550 ;
        RECT 79.130 338.000 82.930 338.550 ;
        RECT 86.530 338.550 102.930 338.600 ;
        RECT 86.530 338.000 90.330 338.550 ;
        RECT 79.130 337.550 79.430 338.000 ;
        RECT 90.030 337.550 90.330 338.000 ;
        RECT 79.130 337.400 82.980 337.550 ;
        RECT 86.480 337.400 90.330 337.550 ;
        RECT 79.130 336.950 79.430 337.400 ;
        RECT 90.030 336.950 90.330 337.400 ;
        RECT 79.130 336.800 82.980 336.950 ;
        RECT 86.480 336.800 90.330 336.950 ;
        RECT 79.130 336.350 79.430 336.800 ;
        RECT 90.030 336.350 90.330 336.800 ;
        RECT 79.130 336.200 82.980 336.350 ;
        RECT 86.480 336.200 90.330 336.350 ;
        RECT 79.130 335.750 79.430 336.200 ;
        RECT 90.030 335.750 90.330 336.200 ;
        RECT 79.130 335.600 82.980 335.750 ;
        RECT 86.480 335.600 90.330 335.750 ;
        RECT 79.130 335.150 79.430 335.600 ;
        RECT 90.030 335.150 90.330 335.600 ;
        RECT 79.130 335.000 82.980 335.150 ;
        RECT 86.480 335.000 90.330 335.150 ;
        RECT 79.130 334.550 79.430 335.000 ;
        RECT 90.030 334.550 90.330 335.000 ;
        RECT 79.130 334.400 82.980 334.550 ;
        RECT 86.480 334.400 90.330 334.550 ;
        RECT 79.130 333.950 79.430 334.400 ;
        RECT 90.030 333.950 90.330 334.400 ;
        RECT 79.130 333.800 82.980 333.950 ;
        RECT 86.480 333.800 90.330 333.950 ;
        RECT 79.130 333.350 79.430 333.800 ;
        RECT 90.030 333.350 90.330 333.800 ;
        RECT 79.130 333.200 82.980 333.350 ;
        RECT 86.480 333.200 90.330 333.350 ;
        RECT 79.130 332.750 79.430 333.200 ;
        RECT 79.130 332.600 82.980 332.750 ;
        RECT 79.130 332.150 79.430 332.600 ;
        RECT 79.130 332.000 82.980 332.150 ;
        RECT 79.130 331.550 79.430 332.000 ;
        RECT 79.130 331.400 82.980 331.550 ;
        RECT 79.130 330.950 79.430 331.400 ;
        RECT 79.130 330.800 82.980 330.950 ;
        RECT 79.130 330.350 79.430 330.800 ;
        RECT 75.530 321.450 75.680 329.650 ;
        RECT 76.130 321.450 76.280 329.650 ;
        RECT 76.730 321.450 76.880 329.650 ;
        RECT 77.330 321.450 77.480 329.650 ;
        RECT 77.930 321.450 78.080 329.650 ;
        RECT 78.530 321.450 78.680 329.650 ;
        RECT 79.130 329.200 79.430 329.650 ;
        RECT 79.130 329.050 82.980 329.200 ;
        RECT 79.130 328.600 79.430 329.050 ;
        RECT 79.130 328.450 82.980 328.600 ;
        RECT 79.130 328.000 79.430 328.450 ;
        RECT 79.130 327.850 82.980 328.000 ;
        RECT 79.130 327.400 79.430 327.850 ;
        RECT 79.130 327.250 82.980 327.400 ;
        RECT 79.130 326.800 79.430 327.250 ;
        RECT 83.830 326.800 85.630 333.200 ;
        RECT 90.030 332.750 90.330 333.200 ;
        RECT 86.480 332.600 90.330 332.750 ;
        RECT 90.030 332.150 90.330 332.600 ;
        RECT 86.480 332.000 90.330 332.150 ;
        RECT 90.030 331.550 90.330 332.000 ;
        RECT 86.480 331.400 90.330 331.550 ;
        RECT 90.030 330.950 90.330 331.400 ;
        RECT 86.480 330.800 90.330 330.950 ;
        RECT 90.030 330.350 90.330 330.800 ;
        RECT 90.780 330.350 90.930 338.550 ;
        RECT 91.380 330.350 91.530 338.550 ;
        RECT 91.980 330.350 92.130 338.550 ;
        RECT 92.580 330.350 92.730 338.550 ;
        RECT 93.180 330.350 93.330 338.550 ;
        RECT 93.780 330.350 93.930 338.550 ;
        RECT 90.030 329.200 90.330 329.650 ;
        RECT 86.480 329.050 90.330 329.200 ;
        RECT 90.030 328.600 90.330 329.050 ;
        RECT 86.480 328.450 90.330 328.600 ;
        RECT 90.030 328.000 90.330 328.450 ;
        RECT 86.480 327.850 90.330 328.000 ;
        RECT 90.030 327.400 90.330 327.850 ;
        RECT 86.480 327.250 90.330 327.400 ;
        RECT 90.030 326.800 90.330 327.250 ;
        RECT 79.130 326.650 82.980 326.800 ;
        RECT 86.480 326.650 90.330 326.800 ;
        RECT 79.130 326.200 79.430 326.650 ;
        RECT 90.030 326.200 90.330 326.650 ;
        RECT 79.130 326.050 82.980 326.200 ;
        RECT 86.480 326.050 90.330 326.200 ;
        RECT 79.130 325.600 79.430 326.050 ;
        RECT 90.030 325.600 90.330 326.050 ;
        RECT 79.130 325.450 82.980 325.600 ;
        RECT 86.480 325.450 90.330 325.600 ;
        RECT 79.130 325.000 79.430 325.450 ;
        RECT 90.030 325.000 90.330 325.450 ;
        RECT 79.130 324.850 82.980 325.000 ;
        RECT 86.480 324.850 90.330 325.000 ;
        RECT 79.130 324.400 79.430 324.850 ;
        RECT 90.030 324.400 90.330 324.850 ;
        RECT 79.130 324.250 82.980 324.400 ;
        RECT 86.480 324.250 90.330 324.400 ;
        RECT 79.130 323.800 79.430 324.250 ;
        RECT 90.030 323.800 90.330 324.250 ;
        RECT 79.130 323.650 82.980 323.800 ;
        RECT 86.480 323.650 90.330 323.800 ;
        RECT 79.130 323.200 79.430 323.650 ;
        RECT 90.030 323.200 90.330 323.650 ;
        RECT 79.130 323.050 82.980 323.200 ;
        RECT 86.480 323.050 90.330 323.200 ;
        RECT 79.130 322.600 79.430 323.050 ;
        RECT 90.030 322.600 90.330 323.050 ;
        RECT 79.130 322.450 82.980 322.600 ;
        RECT 86.480 322.450 90.330 322.600 ;
        RECT 79.130 322.000 79.430 322.450 ;
        RECT 90.030 322.000 90.330 322.450 ;
        RECT 79.130 321.450 82.930 322.000 ;
        RECT 66.530 321.400 82.930 321.450 ;
        RECT 86.530 321.450 90.330 322.000 ;
        RECT 90.780 321.450 90.930 329.650 ;
        RECT 91.380 321.450 91.530 329.650 ;
        RECT 91.980 321.450 92.130 329.650 ;
        RECT 92.580 321.450 92.730 329.650 ;
        RECT 93.180 321.450 93.330 329.650 ;
        RECT 93.780 321.450 93.930 329.650 ;
        RECT 94.380 321.450 95.080 338.550 ;
        RECT 95.530 330.350 95.680 338.550 ;
        RECT 96.130 330.350 96.280 338.550 ;
        RECT 96.730 330.350 96.880 338.550 ;
        RECT 97.330 330.350 97.480 338.550 ;
        RECT 97.930 330.350 98.080 338.550 ;
        RECT 98.530 330.350 98.680 338.550 ;
        RECT 99.130 338.000 102.930 338.550 ;
        RECT 99.130 337.550 99.430 338.000 ;
        RECT 99.130 337.400 102.980 337.550 ;
        RECT 99.130 336.950 99.430 337.400 ;
        RECT 99.130 336.800 102.980 336.950 ;
        RECT 99.130 336.350 99.430 336.800 ;
        RECT 99.130 336.200 102.980 336.350 ;
        RECT 99.130 335.750 99.430 336.200 ;
        RECT 99.130 335.600 102.980 335.750 ;
        RECT 99.130 335.150 99.430 335.600 ;
        RECT 99.130 335.000 102.980 335.150 ;
        RECT 99.130 334.550 99.430 335.000 ;
        RECT 99.130 334.400 102.980 334.550 ;
        RECT 99.130 333.950 99.430 334.400 ;
        RECT 99.130 333.800 102.980 333.950 ;
        RECT 99.130 333.350 99.430 333.800 ;
        RECT 99.130 333.200 102.980 333.350 ;
        RECT 99.130 332.750 99.430 333.200 ;
        RECT 99.130 332.600 102.980 332.750 ;
        RECT 99.130 332.150 99.430 332.600 ;
        RECT 99.130 332.000 102.980 332.150 ;
        RECT 99.130 331.550 99.430 332.000 ;
        RECT 99.130 331.400 102.980 331.550 ;
        RECT 99.130 330.950 99.430 331.400 ;
        RECT 99.130 330.800 102.980 330.950 ;
        RECT 99.130 330.350 99.430 330.800 ;
        RECT 95.530 321.450 95.680 329.650 ;
        RECT 96.130 321.450 96.280 329.650 ;
        RECT 96.730 321.450 96.880 329.650 ;
        RECT 97.330 321.450 97.480 329.650 ;
        RECT 97.930 321.450 98.080 329.650 ;
        RECT 98.530 321.450 98.680 329.650 ;
        RECT 99.130 329.200 99.430 329.650 ;
        RECT 99.130 329.050 102.980 329.200 ;
        RECT 99.130 328.600 99.430 329.050 ;
        RECT 99.130 328.450 102.980 328.600 ;
        RECT 99.130 328.000 99.430 328.450 ;
        RECT 99.130 327.850 102.980 328.000 ;
        RECT 99.130 327.400 99.430 327.850 ;
        RECT 99.130 327.250 102.980 327.400 ;
        RECT 99.130 326.800 99.430 327.250 ;
        RECT 103.830 326.800 104.730 333.200 ;
        RECT 109.850 329.140 111.850 330.415 ;
        RECT 99.130 326.650 102.980 326.800 ;
        RECT 99.130 326.200 99.430 326.650 ;
        RECT 99.130 326.050 102.980 326.200 ;
        RECT 99.130 325.600 99.430 326.050 ;
        RECT 99.130 325.450 102.980 325.600 ;
        RECT 99.130 325.000 99.430 325.450 ;
        RECT 99.130 324.850 102.980 325.000 ;
        RECT 99.130 324.400 99.430 324.850 ;
        RECT 99.130 324.250 102.980 324.400 ;
        RECT 99.130 323.800 99.430 324.250 ;
        RECT 99.130 323.650 102.980 323.800 ;
        RECT 99.130 323.200 99.430 323.650 ;
        RECT 99.130 323.050 102.980 323.200 ;
        RECT 99.130 322.600 99.430 323.050 ;
        RECT 99.130 322.450 102.980 322.600 ;
        RECT 99.130 322.000 99.430 322.450 ;
        RECT 99.130 321.450 102.930 322.000 ;
        RECT 86.530 321.400 102.930 321.450 ;
        RECT 9.630 320.900 19.830 321.400 ;
        RECT 29.630 320.900 39.830 321.400 ;
        RECT 49.630 320.900 59.830 321.400 ;
        RECT 69.630 320.900 79.830 321.400 ;
        RECT 89.630 320.900 99.830 321.400 ;
        RECT 11.530 319.100 17.930 320.900 ;
        RECT 31.530 319.100 37.930 320.900 ;
        RECT 51.530 319.100 57.930 320.900 ;
        RECT 71.530 319.100 77.930 320.900 ;
        RECT 91.530 319.100 97.930 320.900 ;
        RECT 9.630 318.600 19.830 319.100 ;
        RECT 29.630 318.600 39.830 319.100 ;
        RECT 49.630 318.600 59.830 319.100 ;
        RECT 69.630 318.600 79.830 319.100 ;
        RECT 89.630 318.600 99.830 319.100 ;
        RECT 6.530 318.550 22.930 318.600 ;
        RECT 6.530 318.000 10.330 318.550 ;
        RECT 10.030 317.550 10.330 318.000 ;
        RECT 6.480 317.400 10.330 317.550 ;
        RECT 10.030 316.950 10.330 317.400 ;
        RECT 6.480 316.800 10.330 316.950 ;
        RECT 10.030 316.350 10.330 316.800 ;
        RECT 6.480 316.200 10.330 316.350 ;
        RECT 10.030 315.750 10.330 316.200 ;
        RECT 6.480 315.600 10.330 315.750 ;
        RECT 10.030 315.150 10.330 315.600 ;
        RECT 6.480 315.000 10.330 315.150 ;
        RECT 10.030 314.550 10.330 315.000 ;
        RECT 6.480 314.400 10.330 314.550 ;
        RECT 10.030 313.950 10.330 314.400 ;
        RECT 6.480 313.800 10.330 313.950 ;
        RECT 10.030 313.350 10.330 313.800 ;
        RECT 6.480 313.200 10.330 313.350 ;
        RECT 4.730 306.800 5.630 313.200 ;
        RECT 10.030 312.750 10.330 313.200 ;
        RECT 6.480 312.600 10.330 312.750 ;
        RECT 10.030 312.150 10.330 312.600 ;
        RECT 6.480 312.000 10.330 312.150 ;
        RECT 10.030 311.550 10.330 312.000 ;
        RECT 6.480 311.400 10.330 311.550 ;
        RECT 10.030 310.950 10.330 311.400 ;
        RECT 6.480 310.800 10.330 310.950 ;
        RECT 10.030 310.350 10.330 310.800 ;
        RECT 10.780 310.350 10.930 318.550 ;
        RECT 11.380 310.350 11.530 318.550 ;
        RECT 11.980 310.350 12.130 318.550 ;
        RECT 12.580 310.350 12.730 318.550 ;
        RECT 13.180 310.350 13.330 318.550 ;
        RECT 13.780 310.350 13.930 318.550 ;
        RECT 10.030 309.200 10.330 309.650 ;
        RECT 6.480 309.050 10.330 309.200 ;
        RECT 10.030 308.600 10.330 309.050 ;
        RECT 6.480 308.450 10.330 308.600 ;
        RECT 10.030 308.000 10.330 308.450 ;
        RECT 6.480 307.850 10.330 308.000 ;
        RECT 10.030 307.400 10.330 307.850 ;
        RECT 6.480 307.250 10.330 307.400 ;
        RECT 10.030 306.800 10.330 307.250 ;
        RECT 6.480 306.650 10.330 306.800 ;
        RECT 10.030 306.200 10.330 306.650 ;
        RECT 6.480 306.050 10.330 306.200 ;
        RECT 10.030 305.600 10.330 306.050 ;
        RECT 6.480 305.450 10.330 305.600 ;
        RECT 10.030 305.000 10.330 305.450 ;
        RECT 6.480 304.850 10.330 305.000 ;
        RECT 10.030 304.400 10.330 304.850 ;
        RECT 6.480 304.250 10.330 304.400 ;
        RECT 10.030 303.800 10.330 304.250 ;
        RECT 6.480 303.650 10.330 303.800 ;
        RECT 10.030 303.200 10.330 303.650 ;
        RECT 6.480 303.050 10.330 303.200 ;
        RECT 10.030 302.600 10.330 303.050 ;
        RECT 6.480 302.450 10.330 302.600 ;
        RECT 10.030 302.000 10.330 302.450 ;
        RECT 6.530 301.450 10.330 302.000 ;
        RECT 10.780 301.450 10.930 309.650 ;
        RECT 11.380 301.450 11.530 309.650 ;
        RECT 11.980 301.450 12.130 309.650 ;
        RECT 12.580 301.450 12.730 309.650 ;
        RECT 13.180 301.450 13.330 309.650 ;
        RECT 13.780 301.450 13.930 309.650 ;
        RECT 14.380 301.450 15.080 318.550 ;
        RECT 15.530 310.350 15.680 318.550 ;
        RECT 16.130 310.350 16.280 318.550 ;
        RECT 16.730 310.350 16.880 318.550 ;
        RECT 17.330 310.350 17.480 318.550 ;
        RECT 17.930 310.350 18.080 318.550 ;
        RECT 18.530 310.350 18.680 318.550 ;
        RECT 19.130 318.000 22.930 318.550 ;
        RECT 26.530 318.550 42.930 318.600 ;
        RECT 26.530 318.000 30.330 318.550 ;
        RECT 19.130 317.550 19.430 318.000 ;
        RECT 30.030 317.550 30.330 318.000 ;
        RECT 19.130 317.400 22.980 317.550 ;
        RECT 26.480 317.400 30.330 317.550 ;
        RECT 19.130 316.950 19.430 317.400 ;
        RECT 30.030 316.950 30.330 317.400 ;
        RECT 19.130 316.800 22.980 316.950 ;
        RECT 26.480 316.800 30.330 316.950 ;
        RECT 19.130 316.350 19.430 316.800 ;
        RECT 30.030 316.350 30.330 316.800 ;
        RECT 19.130 316.200 22.980 316.350 ;
        RECT 26.480 316.200 30.330 316.350 ;
        RECT 19.130 315.750 19.430 316.200 ;
        RECT 30.030 315.750 30.330 316.200 ;
        RECT 19.130 315.600 22.980 315.750 ;
        RECT 26.480 315.600 30.330 315.750 ;
        RECT 19.130 315.150 19.430 315.600 ;
        RECT 30.030 315.150 30.330 315.600 ;
        RECT 19.130 315.000 22.980 315.150 ;
        RECT 26.480 315.000 30.330 315.150 ;
        RECT 19.130 314.550 19.430 315.000 ;
        RECT 30.030 314.550 30.330 315.000 ;
        RECT 19.130 314.400 22.980 314.550 ;
        RECT 26.480 314.400 30.330 314.550 ;
        RECT 19.130 313.950 19.430 314.400 ;
        RECT 30.030 313.950 30.330 314.400 ;
        RECT 19.130 313.800 22.980 313.950 ;
        RECT 26.480 313.800 30.330 313.950 ;
        RECT 19.130 313.350 19.430 313.800 ;
        RECT 30.030 313.350 30.330 313.800 ;
        RECT 19.130 313.200 22.980 313.350 ;
        RECT 26.480 313.200 30.330 313.350 ;
        RECT 19.130 312.750 19.430 313.200 ;
        RECT 19.130 312.600 22.980 312.750 ;
        RECT 19.130 312.150 19.430 312.600 ;
        RECT 19.130 312.000 22.980 312.150 ;
        RECT 19.130 311.550 19.430 312.000 ;
        RECT 19.130 311.400 22.980 311.550 ;
        RECT 19.130 310.950 19.430 311.400 ;
        RECT 19.130 310.800 22.980 310.950 ;
        RECT 19.130 310.350 19.430 310.800 ;
        RECT 15.530 301.450 15.680 309.650 ;
        RECT 16.130 301.450 16.280 309.650 ;
        RECT 16.730 301.450 16.880 309.650 ;
        RECT 17.330 301.450 17.480 309.650 ;
        RECT 17.930 301.450 18.080 309.650 ;
        RECT 18.530 301.450 18.680 309.650 ;
        RECT 19.130 309.200 19.430 309.650 ;
        RECT 19.130 309.050 22.980 309.200 ;
        RECT 19.130 308.600 19.430 309.050 ;
        RECT 19.130 308.450 22.980 308.600 ;
        RECT 19.130 308.000 19.430 308.450 ;
        RECT 19.130 307.850 22.980 308.000 ;
        RECT 19.130 307.400 19.430 307.850 ;
        RECT 19.130 307.250 22.980 307.400 ;
        RECT 19.130 306.800 19.430 307.250 ;
        RECT 23.830 306.800 25.630 313.200 ;
        RECT 30.030 312.750 30.330 313.200 ;
        RECT 26.480 312.600 30.330 312.750 ;
        RECT 30.030 312.150 30.330 312.600 ;
        RECT 26.480 312.000 30.330 312.150 ;
        RECT 30.030 311.550 30.330 312.000 ;
        RECT 26.480 311.400 30.330 311.550 ;
        RECT 30.030 310.950 30.330 311.400 ;
        RECT 26.480 310.800 30.330 310.950 ;
        RECT 30.030 310.350 30.330 310.800 ;
        RECT 30.780 310.350 30.930 318.550 ;
        RECT 31.380 310.350 31.530 318.550 ;
        RECT 31.980 310.350 32.130 318.550 ;
        RECT 32.580 310.350 32.730 318.550 ;
        RECT 33.180 310.350 33.330 318.550 ;
        RECT 33.780 310.350 33.930 318.550 ;
        RECT 30.030 309.200 30.330 309.650 ;
        RECT 26.480 309.050 30.330 309.200 ;
        RECT 30.030 308.600 30.330 309.050 ;
        RECT 26.480 308.450 30.330 308.600 ;
        RECT 30.030 308.000 30.330 308.450 ;
        RECT 26.480 307.850 30.330 308.000 ;
        RECT 30.030 307.400 30.330 307.850 ;
        RECT 26.480 307.250 30.330 307.400 ;
        RECT 30.030 306.800 30.330 307.250 ;
        RECT 19.130 306.650 22.980 306.800 ;
        RECT 26.480 306.650 30.330 306.800 ;
        RECT 19.130 306.200 19.430 306.650 ;
        RECT 30.030 306.200 30.330 306.650 ;
        RECT 19.130 306.050 22.980 306.200 ;
        RECT 26.480 306.050 30.330 306.200 ;
        RECT 19.130 305.600 19.430 306.050 ;
        RECT 30.030 305.600 30.330 306.050 ;
        RECT 19.130 305.450 22.980 305.600 ;
        RECT 26.480 305.450 30.330 305.600 ;
        RECT 19.130 305.000 19.430 305.450 ;
        RECT 30.030 305.000 30.330 305.450 ;
        RECT 19.130 304.850 22.980 305.000 ;
        RECT 26.480 304.850 30.330 305.000 ;
        RECT 19.130 304.400 19.430 304.850 ;
        RECT 30.030 304.400 30.330 304.850 ;
        RECT 19.130 304.250 22.980 304.400 ;
        RECT 26.480 304.250 30.330 304.400 ;
        RECT 19.130 303.800 19.430 304.250 ;
        RECT 30.030 303.800 30.330 304.250 ;
        RECT 19.130 303.650 22.980 303.800 ;
        RECT 26.480 303.650 30.330 303.800 ;
        RECT 19.130 303.200 19.430 303.650 ;
        RECT 30.030 303.200 30.330 303.650 ;
        RECT 19.130 303.050 22.980 303.200 ;
        RECT 26.480 303.050 30.330 303.200 ;
        RECT 19.130 302.600 19.430 303.050 ;
        RECT 30.030 302.600 30.330 303.050 ;
        RECT 19.130 302.450 22.980 302.600 ;
        RECT 26.480 302.450 30.330 302.600 ;
        RECT 19.130 302.000 19.430 302.450 ;
        RECT 30.030 302.000 30.330 302.450 ;
        RECT 19.130 301.450 22.930 302.000 ;
        RECT 6.530 301.400 22.930 301.450 ;
        RECT 26.530 301.450 30.330 302.000 ;
        RECT 30.780 301.450 30.930 309.650 ;
        RECT 31.380 301.450 31.530 309.650 ;
        RECT 31.980 301.450 32.130 309.650 ;
        RECT 32.580 301.450 32.730 309.650 ;
        RECT 33.180 301.450 33.330 309.650 ;
        RECT 33.780 301.450 33.930 309.650 ;
        RECT 34.380 301.450 35.080 318.550 ;
        RECT 35.530 310.350 35.680 318.550 ;
        RECT 36.130 310.350 36.280 318.550 ;
        RECT 36.730 310.350 36.880 318.550 ;
        RECT 37.330 310.350 37.480 318.550 ;
        RECT 37.930 310.350 38.080 318.550 ;
        RECT 38.530 310.350 38.680 318.550 ;
        RECT 39.130 318.000 42.930 318.550 ;
        RECT 46.530 318.550 62.930 318.600 ;
        RECT 46.530 318.000 50.330 318.550 ;
        RECT 39.130 317.550 39.430 318.000 ;
        RECT 50.030 317.550 50.330 318.000 ;
        RECT 39.130 317.400 42.980 317.550 ;
        RECT 46.480 317.400 50.330 317.550 ;
        RECT 39.130 316.950 39.430 317.400 ;
        RECT 50.030 316.950 50.330 317.400 ;
        RECT 39.130 316.800 42.980 316.950 ;
        RECT 46.480 316.800 50.330 316.950 ;
        RECT 39.130 316.350 39.430 316.800 ;
        RECT 50.030 316.350 50.330 316.800 ;
        RECT 39.130 316.200 42.980 316.350 ;
        RECT 46.480 316.200 50.330 316.350 ;
        RECT 39.130 315.750 39.430 316.200 ;
        RECT 50.030 315.750 50.330 316.200 ;
        RECT 39.130 315.600 42.980 315.750 ;
        RECT 46.480 315.600 50.330 315.750 ;
        RECT 39.130 315.150 39.430 315.600 ;
        RECT 50.030 315.150 50.330 315.600 ;
        RECT 39.130 315.000 42.980 315.150 ;
        RECT 46.480 315.000 50.330 315.150 ;
        RECT 39.130 314.550 39.430 315.000 ;
        RECT 50.030 314.550 50.330 315.000 ;
        RECT 39.130 314.400 42.980 314.550 ;
        RECT 46.480 314.400 50.330 314.550 ;
        RECT 39.130 313.950 39.430 314.400 ;
        RECT 50.030 313.950 50.330 314.400 ;
        RECT 39.130 313.800 42.980 313.950 ;
        RECT 46.480 313.800 50.330 313.950 ;
        RECT 39.130 313.350 39.430 313.800 ;
        RECT 50.030 313.350 50.330 313.800 ;
        RECT 39.130 313.200 42.980 313.350 ;
        RECT 46.480 313.200 50.330 313.350 ;
        RECT 39.130 312.750 39.430 313.200 ;
        RECT 39.130 312.600 42.980 312.750 ;
        RECT 39.130 312.150 39.430 312.600 ;
        RECT 39.130 312.000 42.980 312.150 ;
        RECT 39.130 311.550 39.430 312.000 ;
        RECT 39.130 311.400 42.980 311.550 ;
        RECT 39.130 310.950 39.430 311.400 ;
        RECT 39.130 310.800 42.980 310.950 ;
        RECT 39.130 310.350 39.430 310.800 ;
        RECT 35.530 301.450 35.680 309.650 ;
        RECT 36.130 301.450 36.280 309.650 ;
        RECT 36.730 301.450 36.880 309.650 ;
        RECT 37.330 301.450 37.480 309.650 ;
        RECT 37.930 301.450 38.080 309.650 ;
        RECT 38.530 301.450 38.680 309.650 ;
        RECT 39.130 309.200 39.430 309.650 ;
        RECT 39.130 309.050 42.980 309.200 ;
        RECT 39.130 308.600 39.430 309.050 ;
        RECT 39.130 308.450 42.980 308.600 ;
        RECT 39.130 308.000 39.430 308.450 ;
        RECT 39.130 307.850 42.980 308.000 ;
        RECT 39.130 307.400 39.430 307.850 ;
        RECT 39.130 307.250 42.980 307.400 ;
        RECT 39.130 306.800 39.430 307.250 ;
        RECT 43.830 306.800 45.630 313.200 ;
        RECT 50.030 312.750 50.330 313.200 ;
        RECT 46.480 312.600 50.330 312.750 ;
        RECT 50.030 312.150 50.330 312.600 ;
        RECT 46.480 312.000 50.330 312.150 ;
        RECT 50.030 311.550 50.330 312.000 ;
        RECT 46.480 311.400 50.330 311.550 ;
        RECT 50.030 310.950 50.330 311.400 ;
        RECT 46.480 310.800 50.330 310.950 ;
        RECT 50.030 310.350 50.330 310.800 ;
        RECT 50.780 310.350 50.930 318.550 ;
        RECT 51.380 310.350 51.530 318.550 ;
        RECT 51.980 310.350 52.130 318.550 ;
        RECT 52.580 310.350 52.730 318.550 ;
        RECT 53.180 310.350 53.330 318.550 ;
        RECT 53.780 310.350 53.930 318.550 ;
        RECT 50.030 309.200 50.330 309.650 ;
        RECT 46.480 309.050 50.330 309.200 ;
        RECT 50.030 308.600 50.330 309.050 ;
        RECT 46.480 308.450 50.330 308.600 ;
        RECT 50.030 308.000 50.330 308.450 ;
        RECT 46.480 307.850 50.330 308.000 ;
        RECT 50.030 307.400 50.330 307.850 ;
        RECT 46.480 307.250 50.330 307.400 ;
        RECT 50.030 306.800 50.330 307.250 ;
        RECT 39.130 306.650 42.980 306.800 ;
        RECT 46.480 306.650 50.330 306.800 ;
        RECT 39.130 306.200 39.430 306.650 ;
        RECT 50.030 306.200 50.330 306.650 ;
        RECT 39.130 306.050 42.980 306.200 ;
        RECT 46.480 306.050 50.330 306.200 ;
        RECT 39.130 305.600 39.430 306.050 ;
        RECT 50.030 305.600 50.330 306.050 ;
        RECT 39.130 305.450 42.980 305.600 ;
        RECT 46.480 305.450 50.330 305.600 ;
        RECT 39.130 305.000 39.430 305.450 ;
        RECT 50.030 305.000 50.330 305.450 ;
        RECT 39.130 304.850 42.980 305.000 ;
        RECT 46.480 304.850 50.330 305.000 ;
        RECT 39.130 304.400 39.430 304.850 ;
        RECT 50.030 304.400 50.330 304.850 ;
        RECT 39.130 304.250 42.980 304.400 ;
        RECT 46.480 304.250 50.330 304.400 ;
        RECT 39.130 303.800 39.430 304.250 ;
        RECT 50.030 303.800 50.330 304.250 ;
        RECT 39.130 303.650 42.980 303.800 ;
        RECT 46.480 303.650 50.330 303.800 ;
        RECT 39.130 303.200 39.430 303.650 ;
        RECT 50.030 303.200 50.330 303.650 ;
        RECT 39.130 303.050 42.980 303.200 ;
        RECT 46.480 303.050 50.330 303.200 ;
        RECT 39.130 302.600 39.430 303.050 ;
        RECT 50.030 302.600 50.330 303.050 ;
        RECT 39.130 302.450 42.980 302.600 ;
        RECT 46.480 302.450 50.330 302.600 ;
        RECT 39.130 302.000 39.430 302.450 ;
        RECT 50.030 302.000 50.330 302.450 ;
        RECT 39.130 301.450 42.930 302.000 ;
        RECT 26.530 301.400 42.930 301.450 ;
        RECT 46.530 301.450 50.330 302.000 ;
        RECT 50.780 301.450 50.930 309.650 ;
        RECT 51.380 301.450 51.530 309.650 ;
        RECT 51.980 301.450 52.130 309.650 ;
        RECT 52.580 301.450 52.730 309.650 ;
        RECT 53.180 301.450 53.330 309.650 ;
        RECT 53.780 301.450 53.930 309.650 ;
        RECT 54.380 301.450 55.080 318.550 ;
        RECT 55.530 310.350 55.680 318.550 ;
        RECT 56.130 310.350 56.280 318.550 ;
        RECT 56.730 310.350 56.880 318.550 ;
        RECT 57.330 310.350 57.480 318.550 ;
        RECT 57.930 310.350 58.080 318.550 ;
        RECT 58.530 310.350 58.680 318.550 ;
        RECT 59.130 318.000 62.930 318.550 ;
        RECT 66.530 318.550 82.930 318.600 ;
        RECT 66.530 318.000 70.330 318.550 ;
        RECT 59.130 317.550 59.430 318.000 ;
        RECT 70.030 317.550 70.330 318.000 ;
        RECT 59.130 317.400 62.980 317.550 ;
        RECT 66.480 317.400 70.330 317.550 ;
        RECT 59.130 316.950 59.430 317.400 ;
        RECT 70.030 316.950 70.330 317.400 ;
        RECT 59.130 316.800 62.980 316.950 ;
        RECT 66.480 316.800 70.330 316.950 ;
        RECT 59.130 316.350 59.430 316.800 ;
        RECT 70.030 316.350 70.330 316.800 ;
        RECT 59.130 316.200 62.980 316.350 ;
        RECT 66.480 316.200 70.330 316.350 ;
        RECT 59.130 315.750 59.430 316.200 ;
        RECT 70.030 315.750 70.330 316.200 ;
        RECT 59.130 315.600 62.980 315.750 ;
        RECT 66.480 315.600 70.330 315.750 ;
        RECT 59.130 315.150 59.430 315.600 ;
        RECT 70.030 315.150 70.330 315.600 ;
        RECT 59.130 315.000 62.980 315.150 ;
        RECT 66.480 315.000 70.330 315.150 ;
        RECT 59.130 314.550 59.430 315.000 ;
        RECT 70.030 314.550 70.330 315.000 ;
        RECT 59.130 314.400 62.980 314.550 ;
        RECT 66.480 314.400 70.330 314.550 ;
        RECT 59.130 313.950 59.430 314.400 ;
        RECT 70.030 313.950 70.330 314.400 ;
        RECT 59.130 313.800 62.980 313.950 ;
        RECT 66.480 313.800 70.330 313.950 ;
        RECT 59.130 313.350 59.430 313.800 ;
        RECT 70.030 313.350 70.330 313.800 ;
        RECT 59.130 313.200 62.980 313.350 ;
        RECT 66.480 313.200 70.330 313.350 ;
        RECT 59.130 312.750 59.430 313.200 ;
        RECT 59.130 312.600 62.980 312.750 ;
        RECT 59.130 312.150 59.430 312.600 ;
        RECT 59.130 312.000 62.980 312.150 ;
        RECT 59.130 311.550 59.430 312.000 ;
        RECT 59.130 311.400 62.980 311.550 ;
        RECT 59.130 310.950 59.430 311.400 ;
        RECT 59.130 310.800 62.980 310.950 ;
        RECT 59.130 310.350 59.430 310.800 ;
        RECT 55.530 301.450 55.680 309.650 ;
        RECT 56.130 301.450 56.280 309.650 ;
        RECT 56.730 301.450 56.880 309.650 ;
        RECT 57.330 301.450 57.480 309.650 ;
        RECT 57.930 301.450 58.080 309.650 ;
        RECT 58.530 301.450 58.680 309.650 ;
        RECT 59.130 309.200 59.430 309.650 ;
        RECT 59.130 309.050 62.980 309.200 ;
        RECT 59.130 308.600 59.430 309.050 ;
        RECT 59.130 308.450 62.980 308.600 ;
        RECT 59.130 308.000 59.430 308.450 ;
        RECT 59.130 307.850 62.980 308.000 ;
        RECT 59.130 307.400 59.430 307.850 ;
        RECT 59.130 307.250 62.980 307.400 ;
        RECT 59.130 306.800 59.430 307.250 ;
        RECT 63.830 306.800 65.630 313.200 ;
        RECT 70.030 312.750 70.330 313.200 ;
        RECT 66.480 312.600 70.330 312.750 ;
        RECT 70.030 312.150 70.330 312.600 ;
        RECT 66.480 312.000 70.330 312.150 ;
        RECT 70.030 311.550 70.330 312.000 ;
        RECT 66.480 311.400 70.330 311.550 ;
        RECT 70.030 310.950 70.330 311.400 ;
        RECT 66.480 310.800 70.330 310.950 ;
        RECT 70.030 310.350 70.330 310.800 ;
        RECT 70.780 310.350 70.930 318.550 ;
        RECT 71.380 310.350 71.530 318.550 ;
        RECT 71.980 310.350 72.130 318.550 ;
        RECT 72.580 310.350 72.730 318.550 ;
        RECT 73.180 310.350 73.330 318.550 ;
        RECT 73.780 310.350 73.930 318.550 ;
        RECT 70.030 309.200 70.330 309.650 ;
        RECT 66.480 309.050 70.330 309.200 ;
        RECT 70.030 308.600 70.330 309.050 ;
        RECT 66.480 308.450 70.330 308.600 ;
        RECT 70.030 308.000 70.330 308.450 ;
        RECT 66.480 307.850 70.330 308.000 ;
        RECT 70.030 307.400 70.330 307.850 ;
        RECT 66.480 307.250 70.330 307.400 ;
        RECT 70.030 306.800 70.330 307.250 ;
        RECT 59.130 306.650 62.980 306.800 ;
        RECT 66.480 306.650 70.330 306.800 ;
        RECT 59.130 306.200 59.430 306.650 ;
        RECT 70.030 306.200 70.330 306.650 ;
        RECT 59.130 306.050 62.980 306.200 ;
        RECT 66.480 306.050 70.330 306.200 ;
        RECT 59.130 305.600 59.430 306.050 ;
        RECT 70.030 305.600 70.330 306.050 ;
        RECT 59.130 305.450 62.980 305.600 ;
        RECT 66.480 305.450 70.330 305.600 ;
        RECT 59.130 305.000 59.430 305.450 ;
        RECT 70.030 305.000 70.330 305.450 ;
        RECT 59.130 304.850 62.980 305.000 ;
        RECT 66.480 304.850 70.330 305.000 ;
        RECT 59.130 304.400 59.430 304.850 ;
        RECT 70.030 304.400 70.330 304.850 ;
        RECT 59.130 304.250 62.980 304.400 ;
        RECT 66.480 304.250 70.330 304.400 ;
        RECT 59.130 303.800 59.430 304.250 ;
        RECT 70.030 303.800 70.330 304.250 ;
        RECT 59.130 303.650 62.980 303.800 ;
        RECT 66.480 303.650 70.330 303.800 ;
        RECT 59.130 303.200 59.430 303.650 ;
        RECT 70.030 303.200 70.330 303.650 ;
        RECT 59.130 303.050 62.980 303.200 ;
        RECT 66.480 303.050 70.330 303.200 ;
        RECT 59.130 302.600 59.430 303.050 ;
        RECT 70.030 302.600 70.330 303.050 ;
        RECT 59.130 302.450 62.980 302.600 ;
        RECT 66.480 302.450 70.330 302.600 ;
        RECT 59.130 302.000 59.430 302.450 ;
        RECT 70.030 302.000 70.330 302.450 ;
        RECT 59.130 301.450 62.930 302.000 ;
        RECT 46.530 301.400 62.930 301.450 ;
        RECT 66.530 301.450 70.330 302.000 ;
        RECT 70.780 301.450 70.930 309.650 ;
        RECT 71.380 301.450 71.530 309.650 ;
        RECT 71.980 301.450 72.130 309.650 ;
        RECT 72.580 301.450 72.730 309.650 ;
        RECT 73.180 301.450 73.330 309.650 ;
        RECT 73.780 301.450 73.930 309.650 ;
        RECT 74.380 301.450 75.080 318.550 ;
        RECT 75.530 310.350 75.680 318.550 ;
        RECT 76.130 310.350 76.280 318.550 ;
        RECT 76.730 310.350 76.880 318.550 ;
        RECT 77.330 310.350 77.480 318.550 ;
        RECT 77.930 310.350 78.080 318.550 ;
        RECT 78.530 310.350 78.680 318.550 ;
        RECT 79.130 318.000 82.930 318.550 ;
        RECT 86.530 318.550 102.930 318.600 ;
        RECT 86.530 318.000 90.330 318.550 ;
        RECT 79.130 317.550 79.430 318.000 ;
        RECT 90.030 317.550 90.330 318.000 ;
        RECT 79.130 317.400 82.980 317.550 ;
        RECT 86.480 317.400 90.330 317.550 ;
        RECT 79.130 316.950 79.430 317.400 ;
        RECT 90.030 316.950 90.330 317.400 ;
        RECT 79.130 316.800 82.980 316.950 ;
        RECT 86.480 316.800 90.330 316.950 ;
        RECT 79.130 316.350 79.430 316.800 ;
        RECT 90.030 316.350 90.330 316.800 ;
        RECT 79.130 316.200 82.980 316.350 ;
        RECT 86.480 316.200 90.330 316.350 ;
        RECT 79.130 315.750 79.430 316.200 ;
        RECT 90.030 315.750 90.330 316.200 ;
        RECT 79.130 315.600 82.980 315.750 ;
        RECT 86.480 315.600 90.330 315.750 ;
        RECT 79.130 315.150 79.430 315.600 ;
        RECT 90.030 315.150 90.330 315.600 ;
        RECT 79.130 315.000 82.980 315.150 ;
        RECT 86.480 315.000 90.330 315.150 ;
        RECT 79.130 314.550 79.430 315.000 ;
        RECT 90.030 314.550 90.330 315.000 ;
        RECT 79.130 314.400 82.980 314.550 ;
        RECT 86.480 314.400 90.330 314.550 ;
        RECT 79.130 313.950 79.430 314.400 ;
        RECT 90.030 313.950 90.330 314.400 ;
        RECT 79.130 313.800 82.980 313.950 ;
        RECT 86.480 313.800 90.330 313.950 ;
        RECT 79.130 313.350 79.430 313.800 ;
        RECT 90.030 313.350 90.330 313.800 ;
        RECT 79.130 313.200 82.980 313.350 ;
        RECT 86.480 313.200 90.330 313.350 ;
        RECT 79.130 312.750 79.430 313.200 ;
        RECT 79.130 312.600 82.980 312.750 ;
        RECT 79.130 312.150 79.430 312.600 ;
        RECT 79.130 312.000 82.980 312.150 ;
        RECT 79.130 311.550 79.430 312.000 ;
        RECT 79.130 311.400 82.980 311.550 ;
        RECT 79.130 310.950 79.430 311.400 ;
        RECT 79.130 310.800 82.980 310.950 ;
        RECT 79.130 310.350 79.430 310.800 ;
        RECT 75.530 301.450 75.680 309.650 ;
        RECT 76.130 301.450 76.280 309.650 ;
        RECT 76.730 301.450 76.880 309.650 ;
        RECT 77.330 301.450 77.480 309.650 ;
        RECT 77.930 301.450 78.080 309.650 ;
        RECT 78.530 301.450 78.680 309.650 ;
        RECT 79.130 309.200 79.430 309.650 ;
        RECT 79.130 309.050 82.980 309.200 ;
        RECT 79.130 308.600 79.430 309.050 ;
        RECT 79.130 308.450 82.980 308.600 ;
        RECT 79.130 308.000 79.430 308.450 ;
        RECT 79.130 307.850 82.980 308.000 ;
        RECT 79.130 307.400 79.430 307.850 ;
        RECT 79.130 307.250 82.980 307.400 ;
        RECT 79.130 306.800 79.430 307.250 ;
        RECT 83.830 306.800 85.630 313.200 ;
        RECT 90.030 312.750 90.330 313.200 ;
        RECT 86.480 312.600 90.330 312.750 ;
        RECT 90.030 312.150 90.330 312.600 ;
        RECT 86.480 312.000 90.330 312.150 ;
        RECT 90.030 311.550 90.330 312.000 ;
        RECT 86.480 311.400 90.330 311.550 ;
        RECT 90.030 310.950 90.330 311.400 ;
        RECT 86.480 310.800 90.330 310.950 ;
        RECT 90.030 310.350 90.330 310.800 ;
        RECT 90.780 310.350 90.930 318.550 ;
        RECT 91.380 310.350 91.530 318.550 ;
        RECT 91.980 310.350 92.130 318.550 ;
        RECT 92.580 310.350 92.730 318.550 ;
        RECT 93.180 310.350 93.330 318.550 ;
        RECT 93.780 310.350 93.930 318.550 ;
        RECT 90.030 309.200 90.330 309.650 ;
        RECT 86.480 309.050 90.330 309.200 ;
        RECT 90.030 308.600 90.330 309.050 ;
        RECT 86.480 308.450 90.330 308.600 ;
        RECT 90.030 308.000 90.330 308.450 ;
        RECT 86.480 307.850 90.330 308.000 ;
        RECT 90.030 307.400 90.330 307.850 ;
        RECT 86.480 307.250 90.330 307.400 ;
        RECT 90.030 306.800 90.330 307.250 ;
        RECT 79.130 306.650 82.980 306.800 ;
        RECT 86.480 306.650 90.330 306.800 ;
        RECT 79.130 306.200 79.430 306.650 ;
        RECT 90.030 306.200 90.330 306.650 ;
        RECT 79.130 306.050 82.980 306.200 ;
        RECT 86.480 306.050 90.330 306.200 ;
        RECT 79.130 305.600 79.430 306.050 ;
        RECT 90.030 305.600 90.330 306.050 ;
        RECT 79.130 305.450 82.980 305.600 ;
        RECT 86.480 305.450 90.330 305.600 ;
        RECT 79.130 305.000 79.430 305.450 ;
        RECT 90.030 305.000 90.330 305.450 ;
        RECT 79.130 304.850 82.980 305.000 ;
        RECT 86.480 304.850 90.330 305.000 ;
        RECT 79.130 304.400 79.430 304.850 ;
        RECT 90.030 304.400 90.330 304.850 ;
        RECT 79.130 304.250 82.980 304.400 ;
        RECT 86.480 304.250 90.330 304.400 ;
        RECT 79.130 303.800 79.430 304.250 ;
        RECT 90.030 303.800 90.330 304.250 ;
        RECT 79.130 303.650 82.980 303.800 ;
        RECT 86.480 303.650 90.330 303.800 ;
        RECT 79.130 303.200 79.430 303.650 ;
        RECT 90.030 303.200 90.330 303.650 ;
        RECT 79.130 303.050 82.980 303.200 ;
        RECT 86.480 303.050 90.330 303.200 ;
        RECT 79.130 302.600 79.430 303.050 ;
        RECT 90.030 302.600 90.330 303.050 ;
        RECT 79.130 302.450 82.980 302.600 ;
        RECT 86.480 302.450 90.330 302.600 ;
        RECT 79.130 302.000 79.430 302.450 ;
        RECT 90.030 302.000 90.330 302.450 ;
        RECT 79.130 301.450 82.930 302.000 ;
        RECT 66.530 301.400 82.930 301.450 ;
        RECT 86.530 301.450 90.330 302.000 ;
        RECT 90.780 301.450 90.930 309.650 ;
        RECT 91.380 301.450 91.530 309.650 ;
        RECT 91.980 301.450 92.130 309.650 ;
        RECT 92.580 301.450 92.730 309.650 ;
        RECT 93.180 301.450 93.330 309.650 ;
        RECT 93.780 301.450 93.930 309.650 ;
        RECT 94.380 301.450 95.080 318.550 ;
        RECT 95.530 310.350 95.680 318.550 ;
        RECT 96.130 310.350 96.280 318.550 ;
        RECT 96.730 310.350 96.880 318.550 ;
        RECT 97.330 310.350 97.480 318.550 ;
        RECT 97.930 310.350 98.080 318.550 ;
        RECT 98.530 310.350 98.680 318.550 ;
        RECT 99.130 318.000 102.930 318.550 ;
        RECT 99.130 317.550 99.430 318.000 ;
        RECT 99.130 317.400 102.980 317.550 ;
        RECT 99.130 316.950 99.430 317.400 ;
        RECT 99.130 316.800 102.980 316.950 ;
        RECT 99.130 316.350 99.430 316.800 ;
        RECT 99.130 316.200 102.980 316.350 ;
        RECT 99.130 315.750 99.430 316.200 ;
        RECT 99.130 315.600 102.980 315.750 ;
        RECT 99.130 315.150 99.430 315.600 ;
        RECT 99.130 315.000 102.980 315.150 ;
        RECT 99.130 314.550 99.430 315.000 ;
        RECT 99.130 314.400 102.980 314.550 ;
        RECT 99.130 313.950 99.430 314.400 ;
        RECT 99.130 313.800 102.980 313.950 ;
        RECT 99.130 313.350 99.430 313.800 ;
        RECT 99.130 313.200 102.980 313.350 ;
        RECT 99.130 312.750 99.430 313.200 ;
        RECT 99.130 312.600 102.980 312.750 ;
        RECT 99.130 312.150 99.430 312.600 ;
        RECT 99.130 312.000 102.980 312.150 ;
        RECT 99.130 311.550 99.430 312.000 ;
        RECT 99.130 311.400 102.980 311.550 ;
        RECT 99.130 310.950 99.430 311.400 ;
        RECT 99.130 310.800 102.980 310.950 ;
        RECT 99.130 310.350 99.430 310.800 ;
        RECT 95.530 301.450 95.680 309.650 ;
        RECT 96.130 301.450 96.280 309.650 ;
        RECT 96.730 301.450 96.880 309.650 ;
        RECT 97.330 301.450 97.480 309.650 ;
        RECT 97.930 301.450 98.080 309.650 ;
        RECT 98.530 301.450 98.680 309.650 ;
        RECT 99.130 309.200 99.430 309.650 ;
        RECT 99.130 309.050 102.980 309.200 ;
        RECT 99.130 308.600 99.430 309.050 ;
        RECT 99.130 308.450 102.980 308.600 ;
        RECT 99.130 308.000 99.430 308.450 ;
        RECT 99.130 307.850 102.980 308.000 ;
        RECT 99.130 307.400 99.430 307.850 ;
        RECT 99.130 307.250 102.980 307.400 ;
        RECT 99.130 306.800 99.430 307.250 ;
        RECT 103.830 306.800 104.730 313.200 ;
        RECT 109.850 309.135 111.850 310.410 ;
        RECT 99.130 306.650 102.980 306.800 ;
        RECT 99.130 306.200 99.430 306.650 ;
        RECT 99.130 306.050 102.980 306.200 ;
        RECT 99.130 305.600 99.430 306.050 ;
        RECT 99.130 305.450 102.980 305.600 ;
        RECT 99.130 305.000 99.430 305.450 ;
        RECT 99.130 304.850 102.980 305.000 ;
        RECT 99.130 304.400 99.430 304.850 ;
        RECT 99.130 304.250 102.980 304.400 ;
        RECT 99.130 303.800 99.430 304.250 ;
        RECT 99.130 303.650 102.980 303.800 ;
        RECT 99.130 303.200 99.430 303.650 ;
        RECT 99.130 303.050 102.980 303.200 ;
        RECT 99.130 302.600 99.430 303.050 ;
        RECT 99.130 302.450 102.980 302.600 ;
        RECT 99.130 302.000 99.430 302.450 ;
        RECT 99.130 301.450 102.930 302.000 ;
        RECT 86.530 301.400 102.930 301.450 ;
        RECT 9.630 300.900 19.830 301.400 ;
        RECT 29.630 300.900 39.830 301.400 ;
        RECT 49.630 300.900 59.830 301.400 ;
        RECT 69.630 300.900 79.830 301.400 ;
        RECT 89.630 300.900 99.830 301.400 ;
        RECT 11.530 299.100 17.930 300.900 ;
        RECT 31.530 299.100 37.930 300.900 ;
        RECT 51.530 299.100 57.930 300.900 ;
        RECT 71.530 299.100 77.930 300.900 ;
        RECT 91.530 299.100 97.930 300.900 ;
        RECT 9.630 298.600 19.830 299.100 ;
        RECT 29.630 298.600 39.830 299.100 ;
        RECT 49.630 298.600 59.830 299.100 ;
        RECT 69.630 298.600 79.830 299.100 ;
        RECT 89.630 298.600 99.830 299.100 ;
        RECT 6.530 298.550 22.930 298.600 ;
        RECT 6.530 298.000 10.330 298.550 ;
        RECT 10.030 297.550 10.330 298.000 ;
        RECT 6.480 297.400 10.330 297.550 ;
        RECT 10.030 296.950 10.330 297.400 ;
        RECT 6.480 296.800 10.330 296.950 ;
        RECT 10.030 296.350 10.330 296.800 ;
        RECT 6.480 296.200 10.330 296.350 ;
        RECT 10.030 295.750 10.330 296.200 ;
        RECT 6.480 295.600 10.330 295.750 ;
        RECT 10.030 295.150 10.330 295.600 ;
        RECT 6.480 295.000 10.330 295.150 ;
        RECT 10.030 294.550 10.330 295.000 ;
        RECT 6.480 294.400 10.330 294.550 ;
        RECT 10.030 293.950 10.330 294.400 ;
        RECT 6.480 293.800 10.330 293.950 ;
        RECT 10.030 293.350 10.330 293.800 ;
        RECT 6.480 293.200 10.330 293.350 ;
        RECT 4.730 286.800 5.630 293.200 ;
        RECT 10.030 292.750 10.330 293.200 ;
        RECT 6.480 292.600 10.330 292.750 ;
        RECT 10.030 292.150 10.330 292.600 ;
        RECT 6.480 292.000 10.330 292.150 ;
        RECT 10.030 291.550 10.330 292.000 ;
        RECT 6.480 291.400 10.330 291.550 ;
        RECT 10.030 290.950 10.330 291.400 ;
        RECT 6.480 290.800 10.330 290.950 ;
        RECT 10.030 290.350 10.330 290.800 ;
        RECT 10.780 290.350 10.930 298.550 ;
        RECT 11.380 290.350 11.530 298.550 ;
        RECT 11.980 290.350 12.130 298.550 ;
        RECT 12.580 290.350 12.730 298.550 ;
        RECT 13.180 290.350 13.330 298.550 ;
        RECT 13.780 290.350 13.930 298.550 ;
        RECT 10.030 289.200 10.330 289.650 ;
        RECT 6.480 289.050 10.330 289.200 ;
        RECT 10.030 288.600 10.330 289.050 ;
        RECT 6.480 288.450 10.330 288.600 ;
        RECT 10.030 288.000 10.330 288.450 ;
        RECT 6.480 287.850 10.330 288.000 ;
        RECT 10.030 287.400 10.330 287.850 ;
        RECT 6.480 287.250 10.330 287.400 ;
        RECT 10.030 286.800 10.330 287.250 ;
        RECT 6.480 286.650 10.330 286.800 ;
        RECT 10.030 286.200 10.330 286.650 ;
        RECT 6.480 286.050 10.330 286.200 ;
        RECT 10.030 285.600 10.330 286.050 ;
        RECT 6.480 285.450 10.330 285.600 ;
        RECT 10.030 285.000 10.330 285.450 ;
        RECT 6.480 284.850 10.330 285.000 ;
        RECT 10.030 284.400 10.330 284.850 ;
        RECT 6.480 284.250 10.330 284.400 ;
        RECT 10.030 283.800 10.330 284.250 ;
        RECT 6.480 283.650 10.330 283.800 ;
        RECT 10.030 283.200 10.330 283.650 ;
        RECT 6.480 283.050 10.330 283.200 ;
        RECT 10.030 282.600 10.330 283.050 ;
        RECT 6.480 282.450 10.330 282.600 ;
        RECT 10.030 282.000 10.330 282.450 ;
        RECT 6.530 281.450 10.330 282.000 ;
        RECT 10.780 281.450 10.930 289.650 ;
        RECT 11.380 281.450 11.530 289.650 ;
        RECT 11.980 281.450 12.130 289.650 ;
        RECT 12.580 281.450 12.730 289.650 ;
        RECT 13.180 281.450 13.330 289.650 ;
        RECT 13.780 281.450 13.930 289.650 ;
        RECT 14.380 281.450 15.080 298.550 ;
        RECT 15.530 290.350 15.680 298.550 ;
        RECT 16.130 290.350 16.280 298.550 ;
        RECT 16.730 290.350 16.880 298.550 ;
        RECT 17.330 290.350 17.480 298.550 ;
        RECT 17.930 290.350 18.080 298.550 ;
        RECT 18.530 290.350 18.680 298.550 ;
        RECT 19.130 298.000 22.930 298.550 ;
        RECT 26.530 298.550 42.930 298.600 ;
        RECT 26.530 298.000 30.330 298.550 ;
        RECT 19.130 297.550 19.430 298.000 ;
        RECT 30.030 297.550 30.330 298.000 ;
        RECT 19.130 297.400 22.980 297.550 ;
        RECT 26.480 297.400 30.330 297.550 ;
        RECT 19.130 296.950 19.430 297.400 ;
        RECT 30.030 296.950 30.330 297.400 ;
        RECT 19.130 296.800 22.980 296.950 ;
        RECT 26.480 296.800 30.330 296.950 ;
        RECT 19.130 296.350 19.430 296.800 ;
        RECT 30.030 296.350 30.330 296.800 ;
        RECT 19.130 296.200 22.980 296.350 ;
        RECT 26.480 296.200 30.330 296.350 ;
        RECT 19.130 295.750 19.430 296.200 ;
        RECT 30.030 295.750 30.330 296.200 ;
        RECT 19.130 295.600 22.980 295.750 ;
        RECT 26.480 295.600 30.330 295.750 ;
        RECT 19.130 295.150 19.430 295.600 ;
        RECT 30.030 295.150 30.330 295.600 ;
        RECT 19.130 295.000 22.980 295.150 ;
        RECT 26.480 295.000 30.330 295.150 ;
        RECT 19.130 294.550 19.430 295.000 ;
        RECT 30.030 294.550 30.330 295.000 ;
        RECT 19.130 294.400 22.980 294.550 ;
        RECT 26.480 294.400 30.330 294.550 ;
        RECT 19.130 293.950 19.430 294.400 ;
        RECT 30.030 293.950 30.330 294.400 ;
        RECT 19.130 293.800 22.980 293.950 ;
        RECT 26.480 293.800 30.330 293.950 ;
        RECT 19.130 293.350 19.430 293.800 ;
        RECT 30.030 293.350 30.330 293.800 ;
        RECT 19.130 293.200 22.980 293.350 ;
        RECT 26.480 293.200 30.330 293.350 ;
        RECT 19.130 292.750 19.430 293.200 ;
        RECT 19.130 292.600 22.980 292.750 ;
        RECT 19.130 292.150 19.430 292.600 ;
        RECT 19.130 292.000 22.980 292.150 ;
        RECT 19.130 291.550 19.430 292.000 ;
        RECT 19.130 291.400 22.980 291.550 ;
        RECT 19.130 290.950 19.430 291.400 ;
        RECT 19.130 290.800 22.980 290.950 ;
        RECT 19.130 290.350 19.430 290.800 ;
        RECT 15.530 281.450 15.680 289.650 ;
        RECT 16.130 281.450 16.280 289.650 ;
        RECT 16.730 281.450 16.880 289.650 ;
        RECT 17.330 281.450 17.480 289.650 ;
        RECT 17.930 281.450 18.080 289.650 ;
        RECT 18.530 281.450 18.680 289.650 ;
        RECT 19.130 289.200 19.430 289.650 ;
        RECT 19.130 289.050 22.980 289.200 ;
        RECT 19.130 288.600 19.430 289.050 ;
        RECT 19.130 288.450 22.980 288.600 ;
        RECT 19.130 288.000 19.430 288.450 ;
        RECT 19.130 287.850 22.980 288.000 ;
        RECT 19.130 287.400 19.430 287.850 ;
        RECT 19.130 287.250 22.980 287.400 ;
        RECT 19.130 286.800 19.430 287.250 ;
        RECT 23.830 286.800 25.630 293.200 ;
        RECT 30.030 292.750 30.330 293.200 ;
        RECT 26.480 292.600 30.330 292.750 ;
        RECT 30.030 292.150 30.330 292.600 ;
        RECT 26.480 292.000 30.330 292.150 ;
        RECT 30.030 291.550 30.330 292.000 ;
        RECT 26.480 291.400 30.330 291.550 ;
        RECT 30.030 290.950 30.330 291.400 ;
        RECT 26.480 290.800 30.330 290.950 ;
        RECT 30.030 290.350 30.330 290.800 ;
        RECT 30.780 290.350 30.930 298.550 ;
        RECT 31.380 290.350 31.530 298.550 ;
        RECT 31.980 290.350 32.130 298.550 ;
        RECT 32.580 290.350 32.730 298.550 ;
        RECT 33.180 290.350 33.330 298.550 ;
        RECT 33.780 290.350 33.930 298.550 ;
        RECT 30.030 289.200 30.330 289.650 ;
        RECT 26.480 289.050 30.330 289.200 ;
        RECT 30.030 288.600 30.330 289.050 ;
        RECT 26.480 288.450 30.330 288.600 ;
        RECT 30.030 288.000 30.330 288.450 ;
        RECT 26.480 287.850 30.330 288.000 ;
        RECT 30.030 287.400 30.330 287.850 ;
        RECT 26.480 287.250 30.330 287.400 ;
        RECT 30.030 286.800 30.330 287.250 ;
        RECT 19.130 286.650 22.980 286.800 ;
        RECT 26.480 286.650 30.330 286.800 ;
        RECT 19.130 286.200 19.430 286.650 ;
        RECT 30.030 286.200 30.330 286.650 ;
        RECT 19.130 286.050 22.980 286.200 ;
        RECT 26.480 286.050 30.330 286.200 ;
        RECT 19.130 285.600 19.430 286.050 ;
        RECT 30.030 285.600 30.330 286.050 ;
        RECT 19.130 285.450 22.980 285.600 ;
        RECT 26.480 285.450 30.330 285.600 ;
        RECT 19.130 285.000 19.430 285.450 ;
        RECT 30.030 285.000 30.330 285.450 ;
        RECT 19.130 284.850 22.980 285.000 ;
        RECT 26.480 284.850 30.330 285.000 ;
        RECT 19.130 284.400 19.430 284.850 ;
        RECT 30.030 284.400 30.330 284.850 ;
        RECT 19.130 284.250 22.980 284.400 ;
        RECT 26.480 284.250 30.330 284.400 ;
        RECT 19.130 283.800 19.430 284.250 ;
        RECT 30.030 283.800 30.330 284.250 ;
        RECT 19.130 283.650 22.980 283.800 ;
        RECT 26.480 283.650 30.330 283.800 ;
        RECT 19.130 283.200 19.430 283.650 ;
        RECT 30.030 283.200 30.330 283.650 ;
        RECT 19.130 283.050 22.980 283.200 ;
        RECT 26.480 283.050 30.330 283.200 ;
        RECT 19.130 282.600 19.430 283.050 ;
        RECT 30.030 282.600 30.330 283.050 ;
        RECT 19.130 282.450 22.980 282.600 ;
        RECT 26.480 282.450 30.330 282.600 ;
        RECT 19.130 282.000 19.430 282.450 ;
        RECT 30.030 282.000 30.330 282.450 ;
        RECT 19.130 281.450 22.930 282.000 ;
        RECT 6.530 281.400 22.930 281.450 ;
        RECT 26.530 281.450 30.330 282.000 ;
        RECT 30.780 281.450 30.930 289.650 ;
        RECT 31.380 281.450 31.530 289.650 ;
        RECT 31.980 281.450 32.130 289.650 ;
        RECT 32.580 281.450 32.730 289.650 ;
        RECT 33.180 281.450 33.330 289.650 ;
        RECT 33.780 281.450 33.930 289.650 ;
        RECT 34.380 281.450 35.080 298.550 ;
        RECT 35.530 290.350 35.680 298.550 ;
        RECT 36.130 290.350 36.280 298.550 ;
        RECT 36.730 290.350 36.880 298.550 ;
        RECT 37.330 290.350 37.480 298.550 ;
        RECT 37.930 290.350 38.080 298.550 ;
        RECT 38.530 290.350 38.680 298.550 ;
        RECT 39.130 298.000 42.930 298.550 ;
        RECT 46.530 298.550 62.930 298.600 ;
        RECT 46.530 298.000 50.330 298.550 ;
        RECT 39.130 297.550 39.430 298.000 ;
        RECT 50.030 297.550 50.330 298.000 ;
        RECT 39.130 297.400 42.980 297.550 ;
        RECT 46.480 297.400 50.330 297.550 ;
        RECT 39.130 296.950 39.430 297.400 ;
        RECT 50.030 296.950 50.330 297.400 ;
        RECT 39.130 296.800 42.980 296.950 ;
        RECT 46.480 296.800 50.330 296.950 ;
        RECT 39.130 296.350 39.430 296.800 ;
        RECT 50.030 296.350 50.330 296.800 ;
        RECT 39.130 296.200 42.980 296.350 ;
        RECT 46.480 296.200 50.330 296.350 ;
        RECT 39.130 295.750 39.430 296.200 ;
        RECT 50.030 295.750 50.330 296.200 ;
        RECT 39.130 295.600 42.980 295.750 ;
        RECT 46.480 295.600 50.330 295.750 ;
        RECT 39.130 295.150 39.430 295.600 ;
        RECT 50.030 295.150 50.330 295.600 ;
        RECT 39.130 295.000 42.980 295.150 ;
        RECT 46.480 295.000 50.330 295.150 ;
        RECT 39.130 294.550 39.430 295.000 ;
        RECT 50.030 294.550 50.330 295.000 ;
        RECT 39.130 294.400 42.980 294.550 ;
        RECT 46.480 294.400 50.330 294.550 ;
        RECT 39.130 293.950 39.430 294.400 ;
        RECT 50.030 293.950 50.330 294.400 ;
        RECT 39.130 293.800 42.980 293.950 ;
        RECT 46.480 293.800 50.330 293.950 ;
        RECT 39.130 293.350 39.430 293.800 ;
        RECT 50.030 293.350 50.330 293.800 ;
        RECT 39.130 293.200 42.980 293.350 ;
        RECT 46.480 293.200 50.330 293.350 ;
        RECT 39.130 292.750 39.430 293.200 ;
        RECT 39.130 292.600 42.980 292.750 ;
        RECT 39.130 292.150 39.430 292.600 ;
        RECT 39.130 292.000 42.980 292.150 ;
        RECT 39.130 291.550 39.430 292.000 ;
        RECT 39.130 291.400 42.980 291.550 ;
        RECT 39.130 290.950 39.430 291.400 ;
        RECT 39.130 290.800 42.980 290.950 ;
        RECT 39.130 290.350 39.430 290.800 ;
        RECT 35.530 281.450 35.680 289.650 ;
        RECT 36.130 281.450 36.280 289.650 ;
        RECT 36.730 281.450 36.880 289.650 ;
        RECT 37.330 281.450 37.480 289.650 ;
        RECT 37.930 281.450 38.080 289.650 ;
        RECT 38.530 281.450 38.680 289.650 ;
        RECT 39.130 289.200 39.430 289.650 ;
        RECT 39.130 289.050 42.980 289.200 ;
        RECT 39.130 288.600 39.430 289.050 ;
        RECT 39.130 288.450 42.980 288.600 ;
        RECT 39.130 288.000 39.430 288.450 ;
        RECT 39.130 287.850 42.980 288.000 ;
        RECT 39.130 287.400 39.430 287.850 ;
        RECT 39.130 287.250 42.980 287.400 ;
        RECT 39.130 286.800 39.430 287.250 ;
        RECT 43.830 286.800 45.630 293.200 ;
        RECT 50.030 292.750 50.330 293.200 ;
        RECT 46.480 292.600 50.330 292.750 ;
        RECT 50.030 292.150 50.330 292.600 ;
        RECT 46.480 292.000 50.330 292.150 ;
        RECT 50.030 291.550 50.330 292.000 ;
        RECT 46.480 291.400 50.330 291.550 ;
        RECT 50.030 290.950 50.330 291.400 ;
        RECT 46.480 290.800 50.330 290.950 ;
        RECT 50.030 290.350 50.330 290.800 ;
        RECT 50.780 290.350 50.930 298.550 ;
        RECT 51.380 290.350 51.530 298.550 ;
        RECT 51.980 290.350 52.130 298.550 ;
        RECT 52.580 290.350 52.730 298.550 ;
        RECT 53.180 290.350 53.330 298.550 ;
        RECT 53.780 290.350 53.930 298.550 ;
        RECT 50.030 289.200 50.330 289.650 ;
        RECT 46.480 289.050 50.330 289.200 ;
        RECT 50.030 288.600 50.330 289.050 ;
        RECT 46.480 288.450 50.330 288.600 ;
        RECT 50.030 288.000 50.330 288.450 ;
        RECT 46.480 287.850 50.330 288.000 ;
        RECT 50.030 287.400 50.330 287.850 ;
        RECT 46.480 287.250 50.330 287.400 ;
        RECT 50.030 286.800 50.330 287.250 ;
        RECT 39.130 286.650 42.980 286.800 ;
        RECT 46.480 286.650 50.330 286.800 ;
        RECT 39.130 286.200 39.430 286.650 ;
        RECT 50.030 286.200 50.330 286.650 ;
        RECT 39.130 286.050 42.980 286.200 ;
        RECT 46.480 286.050 50.330 286.200 ;
        RECT 39.130 285.600 39.430 286.050 ;
        RECT 50.030 285.600 50.330 286.050 ;
        RECT 39.130 285.450 42.980 285.600 ;
        RECT 46.480 285.450 50.330 285.600 ;
        RECT 39.130 285.000 39.430 285.450 ;
        RECT 50.030 285.000 50.330 285.450 ;
        RECT 39.130 284.850 42.980 285.000 ;
        RECT 46.480 284.850 50.330 285.000 ;
        RECT 39.130 284.400 39.430 284.850 ;
        RECT 50.030 284.400 50.330 284.850 ;
        RECT 39.130 284.250 42.980 284.400 ;
        RECT 46.480 284.250 50.330 284.400 ;
        RECT 39.130 283.800 39.430 284.250 ;
        RECT 50.030 283.800 50.330 284.250 ;
        RECT 39.130 283.650 42.980 283.800 ;
        RECT 46.480 283.650 50.330 283.800 ;
        RECT 39.130 283.200 39.430 283.650 ;
        RECT 50.030 283.200 50.330 283.650 ;
        RECT 39.130 283.050 42.980 283.200 ;
        RECT 46.480 283.050 50.330 283.200 ;
        RECT 39.130 282.600 39.430 283.050 ;
        RECT 50.030 282.600 50.330 283.050 ;
        RECT 39.130 282.450 42.980 282.600 ;
        RECT 46.480 282.450 50.330 282.600 ;
        RECT 39.130 282.000 39.430 282.450 ;
        RECT 50.030 282.000 50.330 282.450 ;
        RECT 39.130 281.450 42.930 282.000 ;
        RECT 26.530 281.400 42.930 281.450 ;
        RECT 46.530 281.450 50.330 282.000 ;
        RECT 50.780 281.450 50.930 289.650 ;
        RECT 51.380 281.450 51.530 289.650 ;
        RECT 51.980 281.450 52.130 289.650 ;
        RECT 52.580 281.450 52.730 289.650 ;
        RECT 53.180 281.450 53.330 289.650 ;
        RECT 53.780 281.450 53.930 289.650 ;
        RECT 54.380 281.450 55.080 298.550 ;
        RECT 55.530 290.350 55.680 298.550 ;
        RECT 56.130 290.350 56.280 298.550 ;
        RECT 56.730 290.350 56.880 298.550 ;
        RECT 57.330 290.350 57.480 298.550 ;
        RECT 57.930 290.350 58.080 298.550 ;
        RECT 58.530 290.350 58.680 298.550 ;
        RECT 59.130 298.000 62.930 298.550 ;
        RECT 66.530 298.550 82.930 298.600 ;
        RECT 66.530 298.000 70.330 298.550 ;
        RECT 59.130 297.550 59.430 298.000 ;
        RECT 70.030 297.550 70.330 298.000 ;
        RECT 59.130 297.400 62.980 297.550 ;
        RECT 66.480 297.400 70.330 297.550 ;
        RECT 59.130 296.950 59.430 297.400 ;
        RECT 70.030 296.950 70.330 297.400 ;
        RECT 59.130 296.800 62.980 296.950 ;
        RECT 66.480 296.800 70.330 296.950 ;
        RECT 59.130 296.350 59.430 296.800 ;
        RECT 70.030 296.350 70.330 296.800 ;
        RECT 59.130 296.200 62.980 296.350 ;
        RECT 66.480 296.200 70.330 296.350 ;
        RECT 59.130 295.750 59.430 296.200 ;
        RECT 70.030 295.750 70.330 296.200 ;
        RECT 59.130 295.600 62.980 295.750 ;
        RECT 66.480 295.600 70.330 295.750 ;
        RECT 59.130 295.150 59.430 295.600 ;
        RECT 70.030 295.150 70.330 295.600 ;
        RECT 59.130 295.000 62.980 295.150 ;
        RECT 66.480 295.000 70.330 295.150 ;
        RECT 59.130 294.550 59.430 295.000 ;
        RECT 70.030 294.550 70.330 295.000 ;
        RECT 59.130 294.400 62.980 294.550 ;
        RECT 66.480 294.400 70.330 294.550 ;
        RECT 59.130 293.950 59.430 294.400 ;
        RECT 70.030 293.950 70.330 294.400 ;
        RECT 59.130 293.800 62.980 293.950 ;
        RECT 66.480 293.800 70.330 293.950 ;
        RECT 59.130 293.350 59.430 293.800 ;
        RECT 70.030 293.350 70.330 293.800 ;
        RECT 59.130 293.200 62.980 293.350 ;
        RECT 66.480 293.200 70.330 293.350 ;
        RECT 59.130 292.750 59.430 293.200 ;
        RECT 59.130 292.600 62.980 292.750 ;
        RECT 59.130 292.150 59.430 292.600 ;
        RECT 59.130 292.000 62.980 292.150 ;
        RECT 59.130 291.550 59.430 292.000 ;
        RECT 59.130 291.400 62.980 291.550 ;
        RECT 59.130 290.950 59.430 291.400 ;
        RECT 59.130 290.800 62.980 290.950 ;
        RECT 59.130 290.350 59.430 290.800 ;
        RECT 55.530 281.450 55.680 289.650 ;
        RECT 56.130 281.450 56.280 289.650 ;
        RECT 56.730 281.450 56.880 289.650 ;
        RECT 57.330 281.450 57.480 289.650 ;
        RECT 57.930 281.450 58.080 289.650 ;
        RECT 58.530 281.450 58.680 289.650 ;
        RECT 59.130 289.200 59.430 289.650 ;
        RECT 59.130 289.050 62.980 289.200 ;
        RECT 59.130 288.600 59.430 289.050 ;
        RECT 59.130 288.450 62.980 288.600 ;
        RECT 59.130 288.000 59.430 288.450 ;
        RECT 59.130 287.850 62.980 288.000 ;
        RECT 59.130 287.400 59.430 287.850 ;
        RECT 59.130 287.250 62.980 287.400 ;
        RECT 59.130 286.800 59.430 287.250 ;
        RECT 63.830 286.800 65.630 293.200 ;
        RECT 70.030 292.750 70.330 293.200 ;
        RECT 66.480 292.600 70.330 292.750 ;
        RECT 70.030 292.150 70.330 292.600 ;
        RECT 66.480 292.000 70.330 292.150 ;
        RECT 70.030 291.550 70.330 292.000 ;
        RECT 66.480 291.400 70.330 291.550 ;
        RECT 70.030 290.950 70.330 291.400 ;
        RECT 66.480 290.800 70.330 290.950 ;
        RECT 70.030 290.350 70.330 290.800 ;
        RECT 70.780 290.350 70.930 298.550 ;
        RECT 71.380 290.350 71.530 298.550 ;
        RECT 71.980 290.350 72.130 298.550 ;
        RECT 72.580 290.350 72.730 298.550 ;
        RECT 73.180 290.350 73.330 298.550 ;
        RECT 73.780 290.350 73.930 298.550 ;
        RECT 70.030 289.200 70.330 289.650 ;
        RECT 66.480 289.050 70.330 289.200 ;
        RECT 70.030 288.600 70.330 289.050 ;
        RECT 66.480 288.450 70.330 288.600 ;
        RECT 70.030 288.000 70.330 288.450 ;
        RECT 66.480 287.850 70.330 288.000 ;
        RECT 70.030 287.400 70.330 287.850 ;
        RECT 66.480 287.250 70.330 287.400 ;
        RECT 70.030 286.800 70.330 287.250 ;
        RECT 59.130 286.650 62.980 286.800 ;
        RECT 66.480 286.650 70.330 286.800 ;
        RECT 59.130 286.200 59.430 286.650 ;
        RECT 70.030 286.200 70.330 286.650 ;
        RECT 59.130 286.050 62.980 286.200 ;
        RECT 66.480 286.050 70.330 286.200 ;
        RECT 59.130 285.600 59.430 286.050 ;
        RECT 70.030 285.600 70.330 286.050 ;
        RECT 59.130 285.450 62.980 285.600 ;
        RECT 66.480 285.450 70.330 285.600 ;
        RECT 59.130 285.000 59.430 285.450 ;
        RECT 70.030 285.000 70.330 285.450 ;
        RECT 59.130 284.850 62.980 285.000 ;
        RECT 66.480 284.850 70.330 285.000 ;
        RECT 59.130 284.400 59.430 284.850 ;
        RECT 70.030 284.400 70.330 284.850 ;
        RECT 59.130 284.250 62.980 284.400 ;
        RECT 66.480 284.250 70.330 284.400 ;
        RECT 59.130 283.800 59.430 284.250 ;
        RECT 70.030 283.800 70.330 284.250 ;
        RECT 59.130 283.650 62.980 283.800 ;
        RECT 66.480 283.650 70.330 283.800 ;
        RECT 59.130 283.200 59.430 283.650 ;
        RECT 70.030 283.200 70.330 283.650 ;
        RECT 59.130 283.050 62.980 283.200 ;
        RECT 66.480 283.050 70.330 283.200 ;
        RECT 59.130 282.600 59.430 283.050 ;
        RECT 70.030 282.600 70.330 283.050 ;
        RECT 59.130 282.450 62.980 282.600 ;
        RECT 66.480 282.450 70.330 282.600 ;
        RECT 59.130 282.000 59.430 282.450 ;
        RECT 70.030 282.000 70.330 282.450 ;
        RECT 59.130 281.450 62.930 282.000 ;
        RECT 46.530 281.400 62.930 281.450 ;
        RECT 66.530 281.450 70.330 282.000 ;
        RECT 70.780 281.450 70.930 289.650 ;
        RECT 71.380 281.450 71.530 289.650 ;
        RECT 71.980 281.450 72.130 289.650 ;
        RECT 72.580 281.450 72.730 289.650 ;
        RECT 73.180 281.450 73.330 289.650 ;
        RECT 73.780 281.450 73.930 289.650 ;
        RECT 74.380 281.450 75.080 298.550 ;
        RECT 75.530 290.350 75.680 298.550 ;
        RECT 76.130 290.350 76.280 298.550 ;
        RECT 76.730 290.350 76.880 298.550 ;
        RECT 77.330 290.350 77.480 298.550 ;
        RECT 77.930 290.350 78.080 298.550 ;
        RECT 78.530 290.350 78.680 298.550 ;
        RECT 79.130 298.000 82.930 298.550 ;
        RECT 86.530 298.550 102.930 298.600 ;
        RECT 86.530 298.000 90.330 298.550 ;
        RECT 79.130 297.550 79.430 298.000 ;
        RECT 90.030 297.550 90.330 298.000 ;
        RECT 79.130 297.400 82.980 297.550 ;
        RECT 86.480 297.400 90.330 297.550 ;
        RECT 79.130 296.950 79.430 297.400 ;
        RECT 90.030 296.950 90.330 297.400 ;
        RECT 79.130 296.800 82.980 296.950 ;
        RECT 86.480 296.800 90.330 296.950 ;
        RECT 79.130 296.350 79.430 296.800 ;
        RECT 90.030 296.350 90.330 296.800 ;
        RECT 79.130 296.200 82.980 296.350 ;
        RECT 86.480 296.200 90.330 296.350 ;
        RECT 79.130 295.750 79.430 296.200 ;
        RECT 90.030 295.750 90.330 296.200 ;
        RECT 79.130 295.600 82.980 295.750 ;
        RECT 86.480 295.600 90.330 295.750 ;
        RECT 79.130 295.150 79.430 295.600 ;
        RECT 90.030 295.150 90.330 295.600 ;
        RECT 79.130 295.000 82.980 295.150 ;
        RECT 86.480 295.000 90.330 295.150 ;
        RECT 79.130 294.550 79.430 295.000 ;
        RECT 90.030 294.550 90.330 295.000 ;
        RECT 79.130 294.400 82.980 294.550 ;
        RECT 86.480 294.400 90.330 294.550 ;
        RECT 79.130 293.950 79.430 294.400 ;
        RECT 90.030 293.950 90.330 294.400 ;
        RECT 79.130 293.800 82.980 293.950 ;
        RECT 86.480 293.800 90.330 293.950 ;
        RECT 79.130 293.350 79.430 293.800 ;
        RECT 90.030 293.350 90.330 293.800 ;
        RECT 79.130 293.200 82.980 293.350 ;
        RECT 86.480 293.200 90.330 293.350 ;
        RECT 79.130 292.750 79.430 293.200 ;
        RECT 79.130 292.600 82.980 292.750 ;
        RECT 79.130 292.150 79.430 292.600 ;
        RECT 79.130 292.000 82.980 292.150 ;
        RECT 79.130 291.550 79.430 292.000 ;
        RECT 79.130 291.400 82.980 291.550 ;
        RECT 79.130 290.950 79.430 291.400 ;
        RECT 79.130 290.800 82.980 290.950 ;
        RECT 79.130 290.350 79.430 290.800 ;
        RECT 75.530 281.450 75.680 289.650 ;
        RECT 76.130 281.450 76.280 289.650 ;
        RECT 76.730 281.450 76.880 289.650 ;
        RECT 77.330 281.450 77.480 289.650 ;
        RECT 77.930 281.450 78.080 289.650 ;
        RECT 78.530 281.450 78.680 289.650 ;
        RECT 79.130 289.200 79.430 289.650 ;
        RECT 79.130 289.050 82.980 289.200 ;
        RECT 79.130 288.600 79.430 289.050 ;
        RECT 79.130 288.450 82.980 288.600 ;
        RECT 79.130 288.000 79.430 288.450 ;
        RECT 79.130 287.850 82.980 288.000 ;
        RECT 79.130 287.400 79.430 287.850 ;
        RECT 79.130 287.250 82.980 287.400 ;
        RECT 79.130 286.800 79.430 287.250 ;
        RECT 83.830 286.800 85.630 293.200 ;
        RECT 90.030 292.750 90.330 293.200 ;
        RECT 86.480 292.600 90.330 292.750 ;
        RECT 90.030 292.150 90.330 292.600 ;
        RECT 86.480 292.000 90.330 292.150 ;
        RECT 90.030 291.550 90.330 292.000 ;
        RECT 86.480 291.400 90.330 291.550 ;
        RECT 90.030 290.950 90.330 291.400 ;
        RECT 86.480 290.800 90.330 290.950 ;
        RECT 90.030 290.350 90.330 290.800 ;
        RECT 90.780 290.350 90.930 298.550 ;
        RECT 91.380 290.350 91.530 298.550 ;
        RECT 91.980 290.350 92.130 298.550 ;
        RECT 92.580 290.350 92.730 298.550 ;
        RECT 93.180 290.350 93.330 298.550 ;
        RECT 93.780 290.350 93.930 298.550 ;
        RECT 90.030 289.200 90.330 289.650 ;
        RECT 86.480 289.050 90.330 289.200 ;
        RECT 90.030 288.600 90.330 289.050 ;
        RECT 86.480 288.450 90.330 288.600 ;
        RECT 90.030 288.000 90.330 288.450 ;
        RECT 86.480 287.850 90.330 288.000 ;
        RECT 90.030 287.400 90.330 287.850 ;
        RECT 86.480 287.250 90.330 287.400 ;
        RECT 90.030 286.800 90.330 287.250 ;
        RECT 79.130 286.650 82.980 286.800 ;
        RECT 86.480 286.650 90.330 286.800 ;
        RECT 79.130 286.200 79.430 286.650 ;
        RECT 90.030 286.200 90.330 286.650 ;
        RECT 79.130 286.050 82.980 286.200 ;
        RECT 86.480 286.050 90.330 286.200 ;
        RECT 79.130 285.600 79.430 286.050 ;
        RECT 90.030 285.600 90.330 286.050 ;
        RECT 79.130 285.450 82.980 285.600 ;
        RECT 86.480 285.450 90.330 285.600 ;
        RECT 79.130 285.000 79.430 285.450 ;
        RECT 90.030 285.000 90.330 285.450 ;
        RECT 79.130 284.850 82.980 285.000 ;
        RECT 86.480 284.850 90.330 285.000 ;
        RECT 79.130 284.400 79.430 284.850 ;
        RECT 90.030 284.400 90.330 284.850 ;
        RECT 79.130 284.250 82.980 284.400 ;
        RECT 86.480 284.250 90.330 284.400 ;
        RECT 79.130 283.800 79.430 284.250 ;
        RECT 90.030 283.800 90.330 284.250 ;
        RECT 79.130 283.650 82.980 283.800 ;
        RECT 86.480 283.650 90.330 283.800 ;
        RECT 79.130 283.200 79.430 283.650 ;
        RECT 90.030 283.200 90.330 283.650 ;
        RECT 79.130 283.050 82.980 283.200 ;
        RECT 86.480 283.050 90.330 283.200 ;
        RECT 79.130 282.600 79.430 283.050 ;
        RECT 90.030 282.600 90.330 283.050 ;
        RECT 79.130 282.450 82.980 282.600 ;
        RECT 86.480 282.450 90.330 282.600 ;
        RECT 79.130 282.000 79.430 282.450 ;
        RECT 90.030 282.000 90.330 282.450 ;
        RECT 79.130 281.450 82.930 282.000 ;
        RECT 66.530 281.400 82.930 281.450 ;
        RECT 86.530 281.450 90.330 282.000 ;
        RECT 90.780 281.450 90.930 289.650 ;
        RECT 91.380 281.450 91.530 289.650 ;
        RECT 91.980 281.450 92.130 289.650 ;
        RECT 92.580 281.450 92.730 289.650 ;
        RECT 93.180 281.450 93.330 289.650 ;
        RECT 93.780 281.450 93.930 289.650 ;
        RECT 94.380 281.450 95.080 298.550 ;
        RECT 95.530 290.350 95.680 298.550 ;
        RECT 96.130 290.350 96.280 298.550 ;
        RECT 96.730 290.350 96.880 298.550 ;
        RECT 97.330 290.350 97.480 298.550 ;
        RECT 97.930 290.350 98.080 298.550 ;
        RECT 98.530 290.350 98.680 298.550 ;
        RECT 99.130 298.000 102.930 298.550 ;
        RECT 99.130 297.550 99.430 298.000 ;
        RECT 99.130 297.400 102.980 297.550 ;
        RECT 99.130 296.950 99.430 297.400 ;
        RECT 99.130 296.800 102.980 296.950 ;
        RECT 99.130 296.350 99.430 296.800 ;
        RECT 99.130 296.200 102.980 296.350 ;
        RECT 99.130 295.750 99.430 296.200 ;
        RECT 99.130 295.600 102.980 295.750 ;
        RECT 99.130 295.150 99.430 295.600 ;
        RECT 99.130 295.000 102.980 295.150 ;
        RECT 99.130 294.550 99.430 295.000 ;
        RECT 99.130 294.400 102.980 294.550 ;
        RECT 99.130 293.950 99.430 294.400 ;
        RECT 99.130 293.800 102.980 293.950 ;
        RECT 99.130 293.350 99.430 293.800 ;
        RECT 99.130 293.200 102.980 293.350 ;
        RECT 99.130 292.750 99.430 293.200 ;
        RECT 99.130 292.600 102.980 292.750 ;
        RECT 99.130 292.150 99.430 292.600 ;
        RECT 99.130 292.000 102.980 292.150 ;
        RECT 99.130 291.550 99.430 292.000 ;
        RECT 99.130 291.400 102.980 291.550 ;
        RECT 99.130 290.950 99.430 291.400 ;
        RECT 99.130 290.800 102.980 290.950 ;
        RECT 99.130 290.350 99.430 290.800 ;
        RECT 95.530 281.450 95.680 289.650 ;
        RECT 96.130 281.450 96.280 289.650 ;
        RECT 96.730 281.450 96.880 289.650 ;
        RECT 97.330 281.450 97.480 289.650 ;
        RECT 97.930 281.450 98.080 289.650 ;
        RECT 98.530 281.450 98.680 289.650 ;
        RECT 99.130 289.200 99.430 289.650 ;
        RECT 99.130 289.050 102.980 289.200 ;
        RECT 99.130 288.600 99.430 289.050 ;
        RECT 99.130 288.450 102.980 288.600 ;
        RECT 99.130 288.000 99.430 288.450 ;
        RECT 99.130 287.850 102.980 288.000 ;
        RECT 99.130 287.400 99.430 287.850 ;
        RECT 99.130 287.250 102.980 287.400 ;
        RECT 99.130 286.800 99.430 287.250 ;
        RECT 103.830 286.800 104.730 293.200 ;
        RECT 109.850 289.330 111.850 290.605 ;
        RECT 99.130 286.650 102.980 286.800 ;
        RECT 99.130 286.200 99.430 286.650 ;
        RECT 99.130 286.050 102.980 286.200 ;
        RECT 99.130 285.600 99.430 286.050 ;
        RECT 99.130 285.450 102.980 285.600 ;
        RECT 99.130 285.000 99.430 285.450 ;
        RECT 99.130 284.850 102.980 285.000 ;
        RECT 99.130 284.400 99.430 284.850 ;
        RECT 99.130 284.250 102.980 284.400 ;
        RECT 99.130 283.800 99.430 284.250 ;
        RECT 99.130 283.650 102.980 283.800 ;
        RECT 99.130 283.200 99.430 283.650 ;
        RECT 99.130 283.050 102.980 283.200 ;
        RECT 99.130 282.600 99.430 283.050 ;
        RECT 99.130 282.450 102.980 282.600 ;
        RECT 99.130 282.000 99.430 282.450 ;
        RECT 99.130 281.450 102.930 282.000 ;
        RECT 86.530 281.400 102.930 281.450 ;
        RECT 9.630 280.900 19.830 281.400 ;
        RECT 29.630 280.900 39.830 281.400 ;
        RECT 49.630 280.900 59.830 281.400 ;
        RECT 69.630 280.900 79.830 281.400 ;
        RECT 89.630 280.900 99.830 281.400 ;
        RECT 11.530 279.100 17.930 280.900 ;
        RECT 31.530 279.100 37.930 280.900 ;
        RECT 51.530 279.100 57.930 280.900 ;
        RECT 71.530 279.100 77.930 280.900 ;
        RECT 91.530 279.100 97.930 280.900 ;
        RECT 9.630 278.600 19.830 279.100 ;
        RECT 29.630 278.600 39.830 279.100 ;
        RECT 49.630 278.600 59.830 279.100 ;
        RECT 69.630 278.600 79.830 279.100 ;
        RECT 89.630 278.600 99.830 279.100 ;
        RECT 6.530 278.550 22.930 278.600 ;
        RECT 6.530 278.000 10.330 278.550 ;
        RECT 10.030 277.550 10.330 278.000 ;
        RECT 6.480 277.400 10.330 277.550 ;
        RECT 10.030 276.950 10.330 277.400 ;
        RECT 6.480 276.800 10.330 276.950 ;
        RECT 10.030 276.350 10.330 276.800 ;
        RECT 6.480 276.200 10.330 276.350 ;
        RECT 10.030 275.750 10.330 276.200 ;
        RECT 6.480 275.600 10.330 275.750 ;
        RECT 10.030 275.150 10.330 275.600 ;
        RECT 6.480 275.000 10.330 275.150 ;
        RECT 10.030 274.550 10.330 275.000 ;
        RECT 6.480 274.400 10.330 274.550 ;
        RECT 10.030 273.950 10.330 274.400 ;
        RECT 6.480 273.800 10.330 273.950 ;
        RECT 10.030 273.350 10.330 273.800 ;
        RECT 6.480 273.200 10.330 273.350 ;
        RECT 4.730 266.800 5.630 273.200 ;
        RECT 10.030 272.750 10.330 273.200 ;
        RECT 6.480 272.600 10.330 272.750 ;
        RECT 10.030 272.150 10.330 272.600 ;
        RECT 6.480 272.000 10.330 272.150 ;
        RECT 10.030 271.550 10.330 272.000 ;
        RECT 6.480 271.400 10.330 271.550 ;
        RECT 10.030 270.950 10.330 271.400 ;
        RECT 6.480 270.800 10.330 270.950 ;
        RECT 10.030 270.350 10.330 270.800 ;
        RECT 10.780 270.350 10.930 278.550 ;
        RECT 11.380 270.350 11.530 278.550 ;
        RECT 11.980 270.350 12.130 278.550 ;
        RECT 12.580 270.350 12.730 278.550 ;
        RECT 13.180 270.350 13.330 278.550 ;
        RECT 13.780 270.350 13.930 278.550 ;
        RECT 10.030 269.200 10.330 269.650 ;
        RECT 6.480 269.050 10.330 269.200 ;
        RECT 10.030 268.600 10.330 269.050 ;
        RECT 6.480 268.450 10.330 268.600 ;
        RECT 10.030 268.000 10.330 268.450 ;
        RECT 6.480 267.850 10.330 268.000 ;
        RECT 10.030 267.400 10.330 267.850 ;
        RECT 6.480 267.250 10.330 267.400 ;
        RECT 10.030 266.800 10.330 267.250 ;
        RECT 6.480 266.650 10.330 266.800 ;
        RECT 10.030 266.200 10.330 266.650 ;
        RECT 6.480 266.050 10.330 266.200 ;
        RECT 10.030 265.600 10.330 266.050 ;
        RECT 6.480 265.450 10.330 265.600 ;
        RECT 10.030 265.000 10.330 265.450 ;
        RECT 6.480 264.850 10.330 265.000 ;
        RECT 10.030 264.400 10.330 264.850 ;
        RECT 6.480 264.250 10.330 264.400 ;
        RECT 10.030 263.800 10.330 264.250 ;
        RECT 6.480 263.650 10.330 263.800 ;
        RECT 10.030 263.200 10.330 263.650 ;
        RECT 6.480 263.050 10.330 263.200 ;
        RECT 10.030 262.600 10.330 263.050 ;
        RECT 6.480 262.450 10.330 262.600 ;
        RECT 10.030 262.000 10.330 262.450 ;
        RECT 6.530 261.450 10.330 262.000 ;
        RECT 10.780 261.450 10.930 269.650 ;
        RECT 11.380 261.450 11.530 269.650 ;
        RECT 11.980 261.450 12.130 269.650 ;
        RECT 12.580 261.450 12.730 269.650 ;
        RECT 13.180 261.450 13.330 269.650 ;
        RECT 13.780 261.450 13.930 269.650 ;
        RECT 14.380 261.450 15.080 278.550 ;
        RECT 15.530 270.350 15.680 278.550 ;
        RECT 16.130 270.350 16.280 278.550 ;
        RECT 16.730 270.350 16.880 278.550 ;
        RECT 17.330 270.350 17.480 278.550 ;
        RECT 17.930 270.350 18.080 278.550 ;
        RECT 18.530 270.350 18.680 278.550 ;
        RECT 19.130 278.000 22.930 278.550 ;
        RECT 26.530 278.550 42.930 278.600 ;
        RECT 26.530 278.000 30.330 278.550 ;
        RECT 19.130 277.550 19.430 278.000 ;
        RECT 30.030 277.550 30.330 278.000 ;
        RECT 19.130 277.400 22.980 277.550 ;
        RECT 26.480 277.400 30.330 277.550 ;
        RECT 19.130 276.950 19.430 277.400 ;
        RECT 30.030 276.950 30.330 277.400 ;
        RECT 19.130 276.800 22.980 276.950 ;
        RECT 26.480 276.800 30.330 276.950 ;
        RECT 19.130 276.350 19.430 276.800 ;
        RECT 30.030 276.350 30.330 276.800 ;
        RECT 19.130 276.200 22.980 276.350 ;
        RECT 26.480 276.200 30.330 276.350 ;
        RECT 19.130 275.750 19.430 276.200 ;
        RECT 30.030 275.750 30.330 276.200 ;
        RECT 19.130 275.600 22.980 275.750 ;
        RECT 26.480 275.600 30.330 275.750 ;
        RECT 19.130 275.150 19.430 275.600 ;
        RECT 30.030 275.150 30.330 275.600 ;
        RECT 19.130 275.000 22.980 275.150 ;
        RECT 26.480 275.000 30.330 275.150 ;
        RECT 19.130 274.550 19.430 275.000 ;
        RECT 30.030 274.550 30.330 275.000 ;
        RECT 19.130 274.400 22.980 274.550 ;
        RECT 26.480 274.400 30.330 274.550 ;
        RECT 19.130 273.950 19.430 274.400 ;
        RECT 30.030 273.950 30.330 274.400 ;
        RECT 19.130 273.800 22.980 273.950 ;
        RECT 26.480 273.800 30.330 273.950 ;
        RECT 19.130 273.350 19.430 273.800 ;
        RECT 30.030 273.350 30.330 273.800 ;
        RECT 19.130 273.200 22.980 273.350 ;
        RECT 26.480 273.200 30.330 273.350 ;
        RECT 19.130 272.750 19.430 273.200 ;
        RECT 19.130 272.600 22.980 272.750 ;
        RECT 19.130 272.150 19.430 272.600 ;
        RECT 19.130 272.000 22.980 272.150 ;
        RECT 19.130 271.550 19.430 272.000 ;
        RECT 19.130 271.400 22.980 271.550 ;
        RECT 19.130 270.950 19.430 271.400 ;
        RECT 19.130 270.800 22.980 270.950 ;
        RECT 19.130 270.350 19.430 270.800 ;
        RECT 15.530 261.450 15.680 269.650 ;
        RECT 16.130 261.450 16.280 269.650 ;
        RECT 16.730 261.450 16.880 269.650 ;
        RECT 17.330 261.450 17.480 269.650 ;
        RECT 17.930 261.450 18.080 269.650 ;
        RECT 18.530 261.450 18.680 269.650 ;
        RECT 19.130 269.200 19.430 269.650 ;
        RECT 19.130 269.050 22.980 269.200 ;
        RECT 19.130 268.600 19.430 269.050 ;
        RECT 19.130 268.450 22.980 268.600 ;
        RECT 19.130 268.000 19.430 268.450 ;
        RECT 19.130 267.850 22.980 268.000 ;
        RECT 19.130 267.400 19.430 267.850 ;
        RECT 19.130 267.250 22.980 267.400 ;
        RECT 19.130 266.800 19.430 267.250 ;
        RECT 23.830 266.800 25.630 273.200 ;
        RECT 30.030 272.750 30.330 273.200 ;
        RECT 26.480 272.600 30.330 272.750 ;
        RECT 30.030 272.150 30.330 272.600 ;
        RECT 26.480 272.000 30.330 272.150 ;
        RECT 30.030 271.550 30.330 272.000 ;
        RECT 26.480 271.400 30.330 271.550 ;
        RECT 30.030 270.950 30.330 271.400 ;
        RECT 26.480 270.800 30.330 270.950 ;
        RECT 30.030 270.350 30.330 270.800 ;
        RECT 30.780 270.350 30.930 278.550 ;
        RECT 31.380 270.350 31.530 278.550 ;
        RECT 31.980 270.350 32.130 278.550 ;
        RECT 32.580 270.350 32.730 278.550 ;
        RECT 33.180 270.350 33.330 278.550 ;
        RECT 33.780 270.350 33.930 278.550 ;
        RECT 30.030 269.200 30.330 269.650 ;
        RECT 26.480 269.050 30.330 269.200 ;
        RECT 30.030 268.600 30.330 269.050 ;
        RECT 26.480 268.450 30.330 268.600 ;
        RECT 30.030 268.000 30.330 268.450 ;
        RECT 26.480 267.850 30.330 268.000 ;
        RECT 30.030 267.400 30.330 267.850 ;
        RECT 26.480 267.250 30.330 267.400 ;
        RECT 30.030 266.800 30.330 267.250 ;
        RECT 19.130 266.650 22.980 266.800 ;
        RECT 26.480 266.650 30.330 266.800 ;
        RECT 19.130 266.200 19.430 266.650 ;
        RECT 30.030 266.200 30.330 266.650 ;
        RECT 19.130 266.050 22.980 266.200 ;
        RECT 26.480 266.050 30.330 266.200 ;
        RECT 19.130 265.600 19.430 266.050 ;
        RECT 30.030 265.600 30.330 266.050 ;
        RECT 19.130 265.450 22.980 265.600 ;
        RECT 26.480 265.450 30.330 265.600 ;
        RECT 19.130 265.000 19.430 265.450 ;
        RECT 30.030 265.000 30.330 265.450 ;
        RECT 19.130 264.850 22.980 265.000 ;
        RECT 26.480 264.850 30.330 265.000 ;
        RECT 19.130 264.400 19.430 264.850 ;
        RECT 30.030 264.400 30.330 264.850 ;
        RECT 19.130 264.250 22.980 264.400 ;
        RECT 26.480 264.250 30.330 264.400 ;
        RECT 19.130 263.800 19.430 264.250 ;
        RECT 30.030 263.800 30.330 264.250 ;
        RECT 19.130 263.650 22.980 263.800 ;
        RECT 26.480 263.650 30.330 263.800 ;
        RECT 19.130 263.200 19.430 263.650 ;
        RECT 30.030 263.200 30.330 263.650 ;
        RECT 19.130 263.050 22.980 263.200 ;
        RECT 26.480 263.050 30.330 263.200 ;
        RECT 19.130 262.600 19.430 263.050 ;
        RECT 30.030 262.600 30.330 263.050 ;
        RECT 19.130 262.450 22.980 262.600 ;
        RECT 26.480 262.450 30.330 262.600 ;
        RECT 19.130 262.000 19.430 262.450 ;
        RECT 30.030 262.000 30.330 262.450 ;
        RECT 19.130 261.450 22.930 262.000 ;
        RECT 6.530 261.400 22.930 261.450 ;
        RECT 26.530 261.450 30.330 262.000 ;
        RECT 30.780 261.450 30.930 269.650 ;
        RECT 31.380 261.450 31.530 269.650 ;
        RECT 31.980 261.450 32.130 269.650 ;
        RECT 32.580 261.450 32.730 269.650 ;
        RECT 33.180 261.450 33.330 269.650 ;
        RECT 33.780 261.450 33.930 269.650 ;
        RECT 34.380 261.450 35.080 278.550 ;
        RECT 35.530 270.350 35.680 278.550 ;
        RECT 36.130 270.350 36.280 278.550 ;
        RECT 36.730 270.350 36.880 278.550 ;
        RECT 37.330 270.350 37.480 278.550 ;
        RECT 37.930 270.350 38.080 278.550 ;
        RECT 38.530 270.350 38.680 278.550 ;
        RECT 39.130 278.000 42.930 278.550 ;
        RECT 46.530 278.550 62.930 278.600 ;
        RECT 46.530 278.000 50.330 278.550 ;
        RECT 39.130 277.550 39.430 278.000 ;
        RECT 50.030 277.550 50.330 278.000 ;
        RECT 39.130 277.400 42.980 277.550 ;
        RECT 46.480 277.400 50.330 277.550 ;
        RECT 39.130 276.950 39.430 277.400 ;
        RECT 50.030 276.950 50.330 277.400 ;
        RECT 39.130 276.800 42.980 276.950 ;
        RECT 46.480 276.800 50.330 276.950 ;
        RECT 39.130 276.350 39.430 276.800 ;
        RECT 50.030 276.350 50.330 276.800 ;
        RECT 39.130 276.200 42.980 276.350 ;
        RECT 46.480 276.200 50.330 276.350 ;
        RECT 39.130 275.750 39.430 276.200 ;
        RECT 50.030 275.750 50.330 276.200 ;
        RECT 39.130 275.600 42.980 275.750 ;
        RECT 46.480 275.600 50.330 275.750 ;
        RECT 39.130 275.150 39.430 275.600 ;
        RECT 50.030 275.150 50.330 275.600 ;
        RECT 39.130 275.000 42.980 275.150 ;
        RECT 46.480 275.000 50.330 275.150 ;
        RECT 39.130 274.550 39.430 275.000 ;
        RECT 50.030 274.550 50.330 275.000 ;
        RECT 39.130 274.400 42.980 274.550 ;
        RECT 46.480 274.400 50.330 274.550 ;
        RECT 39.130 273.950 39.430 274.400 ;
        RECT 50.030 273.950 50.330 274.400 ;
        RECT 39.130 273.800 42.980 273.950 ;
        RECT 46.480 273.800 50.330 273.950 ;
        RECT 39.130 273.350 39.430 273.800 ;
        RECT 50.030 273.350 50.330 273.800 ;
        RECT 39.130 273.200 42.980 273.350 ;
        RECT 46.480 273.200 50.330 273.350 ;
        RECT 39.130 272.750 39.430 273.200 ;
        RECT 39.130 272.600 42.980 272.750 ;
        RECT 39.130 272.150 39.430 272.600 ;
        RECT 39.130 272.000 42.980 272.150 ;
        RECT 39.130 271.550 39.430 272.000 ;
        RECT 39.130 271.400 42.980 271.550 ;
        RECT 39.130 270.950 39.430 271.400 ;
        RECT 39.130 270.800 42.980 270.950 ;
        RECT 39.130 270.350 39.430 270.800 ;
        RECT 35.530 261.450 35.680 269.650 ;
        RECT 36.130 261.450 36.280 269.650 ;
        RECT 36.730 261.450 36.880 269.650 ;
        RECT 37.330 261.450 37.480 269.650 ;
        RECT 37.930 261.450 38.080 269.650 ;
        RECT 38.530 261.450 38.680 269.650 ;
        RECT 39.130 269.200 39.430 269.650 ;
        RECT 39.130 269.050 42.980 269.200 ;
        RECT 39.130 268.600 39.430 269.050 ;
        RECT 39.130 268.450 42.980 268.600 ;
        RECT 39.130 268.000 39.430 268.450 ;
        RECT 39.130 267.850 42.980 268.000 ;
        RECT 39.130 267.400 39.430 267.850 ;
        RECT 39.130 267.250 42.980 267.400 ;
        RECT 39.130 266.800 39.430 267.250 ;
        RECT 43.830 266.800 45.630 273.200 ;
        RECT 50.030 272.750 50.330 273.200 ;
        RECT 46.480 272.600 50.330 272.750 ;
        RECT 50.030 272.150 50.330 272.600 ;
        RECT 46.480 272.000 50.330 272.150 ;
        RECT 50.030 271.550 50.330 272.000 ;
        RECT 46.480 271.400 50.330 271.550 ;
        RECT 50.030 270.950 50.330 271.400 ;
        RECT 46.480 270.800 50.330 270.950 ;
        RECT 50.030 270.350 50.330 270.800 ;
        RECT 50.780 270.350 50.930 278.550 ;
        RECT 51.380 270.350 51.530 278.550 ;
        RECT 51.980 270.350 52.130 278.550 ;
        RECT 52.580 270.350 52.730 278.550 ;
        RECT 53.180 270.350 53.330 278.550 ;
        RECT 53.780 270.350 53.930 278.550 ;
        RECT 50.030 269.200 50.330 269.650 ;
        RECT 46.480 269.050 50.330 269.200 ;
        RECT 50.030 268.600 50.330 269.050 ;
        RECT 46.480 268.450 50.330 268.600 ;
        RECT 50.030 268.000 50.330 268.450 ;
        RECT 46.480 267.850 50.330 268.000 ;
        RECT 50.030 267.400 50.330 267.850 ;
        RECT 46.480 267.250 50.330 267.400 ;
        RECT 50.030 266.800 50.330 267.250 ;
        RECT 39.130 266.650 42.980 266.800 ;
        RECT 46.480 266.650 50.330 266.800 ;
        RECT 39.130 266.200 39.430 266.650 ;
        RECT 50.030 266.200 50.330 266.650 ;
        RECT 39.130 266.050 42.980 266.200 ;
        RECT 46.480 266.050 50.330 266.200 ;
        RECT 39.130 265.600 39.430 266.050 ;
        RECT 50.030 265.600 50.330 266.050 ;
        RECT 39.130 265.450 42.980 265.600 ;
        RECT 46.480 265.450 50.330 265.600 ;
        RECT 39.130 265.000 39.430 265.450 ;
        RECT 50.030 265.000 50.330 265.450 ;
        RECT 39.130 264.850 42.980 265.000 ;
        RECT 46.480 264.850 50.330 265.000 ;
        RECT 39.130 264.400 39.430 264.850 ;
        RECT 50.030 264.400 50.330 264.850 ;
        RECT 39.130 264.250 42.980 264.400 ;
        RECT 46.480 264.250 50.330 264.400 ;
        RECT 39.130 263.800 39.430 264.250 ;
        RECT 50.030 263.800 50.330 264.250 ;
        RECT 39.130 263.650 42.980 263.800 ;
        RECT 46.480 263.650 50.330 263.800 ;
        RECT 39.130 263.200 39.430 263.650 ;
        RECT 50.030 263.200 50.330 263.650 ;
        RECT 39.130 263.050 42.980 263.200 ;
        RECT 46.480 263.050 50.330 263.200 ;
        RECT 39.130 262.600 39.430 263.050 ;
        RECT 50.030 262.600 50.330 263.050 ;
        RECT 39.130 262.450 42.980 262.600 ;
        RECT 46.480 262.450 50.330 262.600 ;
        RECT 39.130 262.000 39.430 262.450 ;
        RECT 50.030 262.000 50.330 262.450 ;
        RECT 39.130 261.450 42.930 262.000 ;
        RECT 26.530 261.400 42.930 261.450 ;
        RECT 46.530 261.450 50.330 262.000 ;
        RECT 50.780 261.450 50.930 269.650 ;
        RECT 51.380 261.450 51.530 269.650 ;
        RECT 51.980 261.450 52.130 269.650 ;
        RECT 52.580 261.450 52.730 269.650 ;
        RECT 53.180 261.450 53.330 269.650 ;
        RECT 53.780 261.450 53.930 269.650 ;
        RECT 54.380 261.450 55.080 278.550 ;
        RECT 55.530 270.350 55.680 278.550 ;
        RECT 56.130 270.350 56.280 278.550 ;
        RECT 56.730 270.350 56.880 278.550 ;
        RECT 57.330 270.350 57.480 278.550 ;
        RECT 57.930 270.350 58.080 278.550 ;
        RECT 58.530 270.350 58.680 278.550 ;
        RECT 59.130 278.000 62.930 278.550 ;
        RECT 66.530 278.550 82.930 278.600 ;
        RECT 66.530 278.000 70.330 278.550 ;
        RECT 59.130 277.550 59.430 278.000 ;
        RECT 70.030 277.550 70.330 278.000 ;
        RECT 59.130 277.400 62.980 277.550 ;
        RECT 66.480 277.400 70.330 277.550 ;
        RECT 59.130 276.950 59.430 277.400 ;
        RECT 70.030 276.950 70.330 277.400 ;
        RECT 59.130 276.800 62.980 276.950 ;
        RECT 66.480 276.800 70.330 276.950 ;
        RECT 59.130 276.350 59.430 276.800 ;
        RECT 70.030 276.350 70.330 276.800 ;
        RECT 59.130 276.200 62.980 276.350 ;
        RECT 66.480 276.200 70.330 276.350 ;
        RECT 59.130 275.750 59.430 276.200 ;
        RECT 70.030 275.750 70.330 276.200 ;
        RECT 59.130 275.600 62.980 275.750 ;
        RECT 66.480 275.600 70.330 275.750 ;
        RECT 59.130 275.150 59.430 275.600 ;
        RECT 70.030 275.150 70.330 275.600 ;
        RECT 59.130 275.000 62.980 275.150 ;
        RECT 66.480 275.000 70.330 275.150 ;
        RECT 59.130 274.550 59.430 275.000 ;
        RECT 70.030 274.550 70.330 275.000 ;
        RECT 59.130 274.400 62.980 274.550 ;
        RECT 66.480 274.400 70.330 274.550 ;
        RECT 59.130 273.950 59.430 274.400 ;
        RECT 70.030 273.950 70.330 274.400 ;
        RECT 59.130 273.800 62.980 273.950 ;
        RECT 66.480 273.800 70.330 273.950 ;
        RECT 59.130 273.350 59.430 273.800 ;
        RECT 70.030 273.350 70.330 273.800 ;
        RECT 59.130 273.200 62.980 273.350 ;
        RECT 66.480 273.200 70.330 273.350 ;
        RECT 59.130 272.750 59.430 273.200 ;
        RECT 59.130 272.600 62.980 272.750 ;
        RECT 59.130 272.150 59.430 272.600 ;
        RECT 59.130 272.000 62.980 272.150 ;
        RECT 59.130 271.550 59.430 272.000 ;
        RECT 59.130 271.400 62.980 271.550 ;
        RECT 59.130 270.950 59.430 271.400 ;
        RECT 59.130 270.800 62.980 270.950 ;
        RECT 59.130 270.350 59.430 270.800 ;
        RECT 55.530 261.450 55.680 269.650 ;
        RECT 56.130 261.450 56.280 269.650 ;
        RECT 56.730 261.450 56.880 269.650 ;
        RECT 57.330 261.450 57.480 269.650 ;
        RECT 57.930 261.450 58.080 269.650 ;
        RECT 58.530 261.450 58.680 269.650 ;
        RECT 59.130 269.200 59.430 269.650 ;
        RECT 59.130 269.050 62.980 269.200 ;
        RECT 59.130 268.600 59.430 269.050 ;
        RECT 59.130 268.450 62.980 268.600 ;
        RECT 59.130 268.000 59.430 268.450 ;
        RECT 59.130 267.850 62.980 268.000 ;
        RECT 59.130 267.400 59.430 267.850 ;
        RECT 59.130 267.250 62.980 267.400 ;
        RECT 59.130 266.800 59.430 267.250 ;
        RECT 63.830 266.800 65.630 273.200 ;
        RECT 70.030 272.750 70.330 273.200 ;
        RECT 66.480 272.600 70.330 272.750 ;
        RECT 70.030 272.150 70.330 272.600 ;
        RECT 66.480 272.000 70.330 272.150 ;
        RECT 70.030 271.550 70.330 272.000 ;
        RECT 66.480 271.400 70.330 271.550 ;
        RECT 70.030 270.950 70.330 271.400 ;
        RECT 66.480 270.800 70.330 270.950 ;
        RECT 70.030 270.350 70.330 270.800 ;
        RECT 70.780 270.350 70.930 278.550 ;
        RECT 71.380 270.350 71.530 278.550 ;
        RECT 71.980 270.350 72.130 278.550 ;
        RECT 72.580 270.350 72.730 278.550 ;
        RECT 73.180 270.350 73.330 278.550 ;
        RECT 73.780 270.350 73.930 278.550 ;
        RECT 70.030 269.200 70.330 269.650 ;
        RECT 66.480 269.050 70.330 269.200 ;
        RECT 70.030 268.600 70.330 269.050 ;
        RECT 66.480 268.450 70.330 268.600 ;
        RECT 70.030 268.000 70.330 268.450 ;
        RECT 66.480 267.850 70.330 268.000 ;
        RECT 70.030 267.400 70.330 267.850 ;
        RECT 66.480 267.250 70.330 267.400 ;
        RECT 70.030 266.800 70.330 267.250 ;
        RECT 59.130 266.650 62.980 266.800 ;
        RECT 66.480 266.650 70.330 266.800 ;
        RECT 59.130 266.200 59.430 266.650 ;
        RECT 70.030 266.200 70.330 266.650 ;
        RECT 59.130 266.050 62.980 266.200 ;
        RECT 66.480 266.050 70.330 266.200 ;
        RECT 59.130 265.600 59.430 266.050 ;
        RECT 70.030 265.600 70.330 266.050 ;
        RECT 59.130 265.450 62.980 265.600 ;
        RECT 66.480 265.450 70.330 265.600 ;
        RECT 59.130 265.000 59.430 265.450 ;
        RECT 70.030 265.000 70.330 265.450 ;
        RECT 59.130 264.850 62.980 265.000 ;
        RECT 66.480 264.850 70.330 265.000 ;
        RECT 59.130 264.400 59.430 264.850 ;
        RECT 70.030 264.400 70.330 264.850 ;
        RECT 59.130 264.250 62.980 264.400 ;
        RECT 66.480 264.250 70.330 264.400 ;
        RECT 59.130 263.800 59.430 264.250 ;
        RECT 70.030 263.800 70.330 264.250 ;
        RECT 59.130 263.650 62.980 263.800 ;
        RECT 66.480 263.650 70.330 263.800 ;
        RECT 59.130 263.200 59.430 263.650 ;
        RECT 70.030 263.200 70.330 263.650 ;
        RECT 59.130 263.050 62.980 263.200 ;
        RECT 66.480 263.050 70.330 263.200 ;
        RECT 59.130 262.600 59.430 263.050 ;
        RECT 70.030 262.600 70.330 263.050 ;
        RECT 59.130 262.450 62.980 262.600 ;
        RECT 66.480 262.450 70.330 262.600 ;
        RECT 59.130 262.000 59.430 262.450 ;
        RECT 70.030 262.000 70.330 262.450 ;
        RECT 59.130 261.450 62.930 262.000 ;
        RECT 46.530 261.400 62.930 261.450 ;
        RECT 66.530 261.450 70.330 262.000 ;
        RECT 70.780 261.450 70.930 269.650 ;
        RECT 71.380 261.450 71.530 269.650 ;
        RECT 71.980 261.450 72.130 269.650 ;
        RECT 72.580 261.450 72.730 269.650 ;
        RECT 73.180 261.450 73.330 269.650 ;
        RECT 73.780 261.450 73.930 269.650 ;
        RECT 74.380 261.450 75.080 278.550 ;
        RECT 75.530 270.350 75.680 278.550 ;
        RECT 76.130 270.350 76.280 278.550 ;
        RECT 76.730 270.350 76.880 278.550 ;
        RECT 77.330 270.350 77.480 278.550 ;
        RECT 77.930 270.350 78.080 278.550 ;
        RECT 78.530 270.350 78.680 278.550 ;
        RECT 79.130 278.000 82.930 278.550 ;
        RECT 86.530 278.550 102.930 278.600 ;
        RECT 86.530 278.000 90.330 278.550 ;
        RECT 79.130 277.550 79.430 278.000 ;
        RECT 90.030 277.550 90.330 278.000 ;
        RECT 79.130 277.400 82.980 277.550 ;
        RECT 86.480 277.400 90.330 277.550 ;
        RECT 79.130 276.950 79.430 277.400 ;
        RECT 90.030 276.950 90.330 277.400 ;
        RECT 79.130 276.800 82.980 276.950 ;
        RECT 86.480 276.800 90.330 276.950 ;
        RECT 79.130 276.350 79.430 276.800 ;
        RECT 90.030 276.350 90.330 276.800 ;
        RECT 79.130 276.200 82.980 276.350 ;
        RECT 86.480 276.200 90.330 276.350 ;
        RECT 79.130 275.750 79.430 276.200 ;
        RECT 90.030 275.750 90.330 276.200 ;
        RECT 79.130 275.600 82.980 275.750 ;
        RECT 86.480 275.600 90.330 275.750 ;
        RECT 79.130 275.150 79.430 275.600 ;
        RECT 90.030 275.150 90.330 275.600 ;
        RECT 79.130 275.000 82.980 275.150 ;
        RECT 86.480 275.000 90.330 275.150 ;
        RECT 79.130 274.550 79.430 275.000 ;
        RECT 90.030 274.550 90.330 275.000 ;
        RECT 79.130 274.400 82.980 274.550 ;
        RECT 86.480 274.400 90.330 274.550 ;
        RECT 79.130 273.950 79.430 274.400 ;
        RECT 90.030 273.950 90.330 274.400 ;
        RECT 79.130 273.800 82.980 273.950 ;
        RECT 86.480 273.800 90.330 273.950 ;
        RECT 79.130 273.350 79.430 273.800 ;
        RECT 90.030 273.350 90.330 273.800 ;
        RECT 79.130 273.200 82.980 273.350 ;
        RECT 86.480 273.200 90.330 273.350 ;
        RECT 79.130 272.750 79.430 273.200 ;
        RECT 79.130 272.600 82.980 272.750 ;
        RECT 79.130 272.150 79.430 272.600 ;
        RECT 79.130 272.000 82.980 272.150 ;
        RECT 79.130 271.550 79.430 272.000 ;
        RECT 79.130 271.400 82.980 271.550 ;
        RECT 79.130 270.950 79.430 271.400 ;
        RECT 79.130 270.800 82.980 270.950 ;
        RECT 79.130 270.350 79.430 270.800 ;
        RECT 75.530 261.450 75.680 269.650 ;
        RECT 76.130 261.450 76.280 269.650 ;
        RECT 76.730 261.450 76.880 269.650 ;
        RECT 77.330 261.450 77.480 269.650 ;
        RECT 77.930 261.450 78.080 269.650 ;
        RECT 78.530 261.450 78.680 269.650 ;
        RECT 79.130 269.200 79.430 269.650 ;
        RECT 79.130 269.050 82.980 269.200 ;
        RECT 79.130 268.600 79.430 269.050 ;
        RECT 79.130 268.450 82.980 268.600 ;
        RECT 79.130 268.000 79.430 268.450 ;
        RECT 79.130 267.850 82.980 268.000 ;
        RECT 79.130 267.400 79.430 267.850 ;
        RECT 79.130 267.250 82.980 267.400 ;
        RECT 79.130 266.800 79.430 267.250 ;
        RECT 83.830 266.800 85.630 273.200 ;
        RECT 90.030 272.750 90.330 273.200 ;
        RECT 86.480 272.600 90.330 272.750 ;
        RECT 90.030 272.150 90.330 272.600 ;
        RECT 86.480 272.000 90.330 272.150 ;
        RECT 90.030 271.550 90.330 272.000 ;
        RECT 86.480 271.400 90.330 271.550 ;
        RECT 90.030 270.950 90.330 271.400 ;
        RECT 86.480 270.800 90.330 270.950 ;
        RECT 90.030 270.350 90.330 270.800 ;
        RECT 90.780 270.350 90.930 278.550 ;
        RECT 91.380 270.350 91.530 278.550 ;
        RECT 91.980 270.350 92.130 278.550 ;
        RECT 92.580 270.350 92.730 278.550 ;
        RECT 93.180 270.350 93.330 278.550 ;
        RECT 93.780 270.350 93.930 278.550 ;
        RECT 90.030 269.200 90.330 269.650 ;
        RECT 86.480 269.050 90.330 269.200 ;
        RECT 90.030 268.600 90.330 269.050 ;
        RECT 86.480 268.450 90.330 268.600 ;
        RECT 90.030 268.000 90.330 268.450 ;
        RECT 86.480 267.850 90.330 268.000 ;
        RECT 90.030 267.400 90.330 267.850 ;
        RECT 86.480 267.250 90.330 267.400 ;
        RECT 90.030 266.800 90.330 267.250 ;
        RECT 79.130 266.650 82.980 266.800 ;
        RECT 86.480 266.650 90.330 266.800 ;
        RECT 79.130 266.200 79.430 266.650 ;
        RECT 90.030 266.200 90.330 266.650 ;
        RECT 79.130 266.050 82.980 266.200 ;
        RECT 86.480 266.050 90.330 266.200 ;
        RECT 79.130 265.600 79.430 266.050 ;
        RECT 90.030 265.600 90.330 266.050 ;
        RECT 79.130 265.450 82.980 265.600 ;
        RECT 86.480 265.450 90.330 265.600 ;
        RECT 79.130 265.000 79.430 265.450 ;
        RECT 90.030 265.000 90.330 265.450 ;
        RECT 79.130 264.850 82.980 265.000 ;
        RECT 86.480 264.850 90.330 265.000 ;
        RECT 79.130 264.400 79.430 264.850 ;
        RECT 90.030 264.400 90.330 264.850 ;
        RECT 79.130 264.250 82.980 264.400 ;
        RECT 86.480 264.250 90.330 264.400 ;
        RECT 79.130 263.800 79.430 264.250 ;
        RECT 90.030 263.800 90.330 264.250 ;
        RECT 79.130 263.650 82.980 263.800 ;
        RECT 86.480 263.650 90.330 263.800 ;
        RECT 79.130 263.200 79.430 263.650 ;
        RECT 90.030 263.200 90.330 263.650 ;
        RECT 79.130 263.050 82.980 263.200 ;
        RECT 86.480 263.050 90.330 263.200 ;
        RECT 79.130 262.600 79.430 263.050 ;
        RECT 90.030 262.600 90.330 263.050 ;
        RECT 79.130 262.450 82.980 262.600 ;
        RECT 86.480 262.450 90.330 262.600 ;
        RECT 79.130 262.000 79.430 262.450 ;
        RECT 90.030 262.000 90.330 262.450 ;
        RECT 79.130 261.450 82.930 262.000 ;
        RECT 66.530 261.400 82.930 261.450 ;
        RECT 86.530 261.450 90.330 262.000 ;
        RECT 90.780 261.450 90.930 269.650 ;
        RECT 91.380 261.450 91.530 269.650 ;
        RECT 91.980 261.450 92.130 269.650 ;
        RECT 92.580 261.450 92.730 269.650 ;
        RECT 93.180 261.450 93.330 269.650 ;
        RECT 93.780 261.450 93.930 269.650 ;
        RECT 94.380 261.450 95.080 278.550 ;
        RECT 95.530 270.350 95.680 278.550 ;
        RECT 96.130 270.350 96.280 278.550 ;
        RECT 96.730 270.350 96.880 278.550 ;
        RECT 97.330 270.350 97.480 278.550 ;
        RECT 97.930 270.350 98.080 278.550 ;
        RECT 98.530 270.350 98.680 278.550 ;
        RECT 99.130 278.000 102.930 278.550 ;
        RECT 99.130 277.550 99.430 278.000 ;
        RECT 99.130 277.400 102.980 277.550 ;
        RECT 99.130 276.950 99.430 277.400 ;
        RECT 99.130 276.800 102.980 276.950 ;
        RECT 99.130 276.350 99.430 276.800 ;
        RECT 99.130 276.200 102.980 276.350 ;
        RECT 99.130 275.750 99.430 276.200 ;
        RECT 99.130 275.600 102.980 275.750 ;
        RECT 99.130 275.150 99.430 275.600 ;
        RECT 99.130 275.000 102.980 275.150 ;
        RECT 99.130 274.550 99.430 275.000 ;
        RECT 99.130 274.400 102.980 274.550 ;
        RECT 99.130 273.950 99.430 274.400 ;
        RECT 99.130 273.800 102.980 273.950 ;
        RECT 99.130 273.350 99.430 273.800 ;
        RECT 99.130 273.200 102.980 273.350 ;
        RECT 99.130 272.750 99.430 273.200 ;
        RECT 99.130 272.600 102.980 272.750 ;
        RECT 99.130 272.150 99.430 272.600 ;
        RECT 99.130 272.000 102.980 272.150 ;
        RECT 99.130 271.550 99.430 272.000 ;
        RECT 99.130 271.400 102.980 271.550 ;
        RECT 99.130 270.950 99.430 271.400 ;
        RECT 99.130 270.800 102.980 270.950 ;
        RECT 99.130 270.350 99.430 270.800 ;
        RECT 95.530 261.450 95.680 269.650 ;
        RECT 96.130 261.450 96.280 269.650 ;
        RECT 96.730 261.450 96.880 269.650 ;
        RECT 97.330 261.450 97.480 269.650 ;
        RECT 97.930 261.450 98.080 269.650 ;
        RECT 98.530 261.450 98.680 269.650 ;
        RECT 99.130 269.200 99.430 269.650 ;
        RECT 99.130 269.050 102.980 269.200 ;
        RECT 99.130 268.600 99.430 269.050 ;
        RECT 99.130 268.450 102.980 268.600 ;
        RECT 99.130 268.000 99.430 268.450 ;
        RECT 99.130 267.850 102.980 268.000 ;
        RECT 99.130 267.400 99.430 267.850 ;
        RECT 99.130 267.250 102.980 267.400 ;
        RECT 99.130 266.800 99.430 267.250 ;
        RECT 103.830 266.800 104.730 273.200 ;
        RECT 109.850 269.245 111.850 270.520 ;
        RECT 99.130 266.650 102.980 266.800 ;
        RECT 99.130 266.200 99.430 266.650 ;
        RECT 99.130 266.050 102.980 266.200 ;
        RECT 99.130 265.600 99.430 266.050 ;
        RECT 99.130 265.450 102.980 265.600 ;
        RECT 99.130 265.000 99.430 265.450 ;
        RECT 99.130 264.850 102.980 265.000 ;
        RECT 99.130 264.400 99.430 264.850 ;
        RECT 99.130 264.250 102.980 264.400 ;
        RECT 99.130 263.800 99.430 264.250 ;
        RECT 99.130 263.650 102.980 263.800 ;
        RECT 99.130 263.200 99.430 263.650 ;
        RECT 99.130 263.050 102.980 263.200 ;
        RECT 99.130 262.600 99.430 263.050 ;
        RECT 99.130 262.450 102.980 262.600 ;
        RECT 99.130 262.000 99.430 262.450 ;
        RECT 99.130 261.450 102.930 262.000 ;
        RECT 86.530 261.400 102.930 261.450 ;
        RECT 9.630 260.900 19.830 261.400 ;
        RECT 29.630 260.900 39.830 261.400 ;
        RECT 49.630 260.900 59.830 261.400 ;
        RECT 69.630 260.900 79.830 261.400 ;
        RECT 89.630 260.900 99.830 261.400 ;
        RECT 11.530 259.100 17.930 260.900 ;
        RECT 31.530 259.100 37.930 260.900 ;
        RECT 51.530 259.100 57.930 260.900 ;
        RECT 71.530 259.100 77.930 260.900 ;
        RECT 91.530 259.100 97.930 260.900 ;
        RECT 9.630 258.600 19.830 259.100 ;
        RECT 29.630 258.600 39.830 259.100 ;
        RECT 49.630 258.600 59.830 259.100 ;
        RECT 69.630 258.600 79.830 259.100 ;
        RECT 89.630 258.600 99.830 259.100 ;
        RECT 6.530 258.550 22.930 258.600 ;
        RECT 6.530 258.000 10.330 258.550 ;
        RECT 10.030 257.550 10.330 258.000 ;
        RECT 6.480 257.400 10.330 257.550 ;
        RECT 10.030 256.950 10.330 257.400 ;
        RECT 6.480 256.800 10.330 256.950 ;
        RECT 10.030 256.350 10.330 256.800 ;
        RECT 6.480 256.200 10.330 256.350 ;
        RECT 10.030 255.750 10.330 256.200 ;
        RECT 6.480 255.600 10.330 255.750 ;
        RECT 10.030 255.150 10.330 255.600 ;
        RECT 6.480 255.000 10.330 255.150 ;
        RECT 10.030 254.550 10.330 255.000 ;
        RECT 6.480 254.400 10.330 254.550 ;
        RECT 10.030 253.950 10.330 254.400 ;
        RECT 6.480 253.800 10.330 253.950 ;
        RECT 10.030 253.350 10.330 253.800 ;
        RECT 6.480 253.200 10.330 253.350 ;
        RECT 4.730 246.800 5.630 253.200 ;
        RECT 10.030 252.750 10.330 253.200 ;
        RECT 6.480 252.600 10.330 252.750 ;
        RECT 10.030 252.150 10.330 252.600 ;
        RECT 6.480 252.000 10.330 252.150 ;
        RECT 10.030 251.550 10.330 252.000 ;
        RECT 6.480 251.400 10.330 251.550 ;
        RECT 10.030 250.950 10.330 251.400 ;
        RECT 6.480 250.800 10.330 250.950 ;
        RECT 10.030 250.350 10.330 250.800 ;
        RECT 10.780 250.350 10.930 258.550 ;
        RECT 11.380 250.350 11.530 258.550 ;
        RECT 11.980 250.350 12.130 258.550 ;
        RECT 12.580 250.350 12.730 258.550 ;
        RECT 13.180 250.350 13.330 258.550 ;
        RECT 13.780 250.350 13.930 258.550 ;
        RECT 10.030 249.200 10.330 249.650 ;
        RECT 6.480 249.050 10.330 249.200 ;
        RECT 10.030 248.600 10.330 249.050 ;
        RECT 6.480 248.450 10.330 248.600 ;
        RECT 10.030 248.000 10.330 248.450 ;
        RECT 6.480 247.850 10.330 248.000 ;
        RECT 10.030 247.400 10.330 247.850 ;
        RECT 6.480 247.250 10.330 247.400 ;
        RECT 10.030 246.800 10.330 247.250 ;
        RECT 6.480 246.650 10.330 246.800 ;
        RECT 10.030 246.200 10.330 246.650 ;
        RECT 6.480 246.050 10.330 246.200 ;
        RECT 10.030 245.600 10.330 246.050 ;
        RECT 6.480 245.450 10.330 245.600 ;
        RECT 10.030 245.000 10.330 245.450 ;
        RECT 6.480 244.850 10.330 245.000 ;
        RECT 10.030 244.400 10.330 244.850 ;
        RECT 6.480 244.250 10.330 244.400 ;
        RECT 10.030 243.800 10.330 244.250 ;
        RECT 6.480 243.650 10.330 243.800 ;
        RECT 10.030 243.200 10.330 243.650 ;
        RECT 6.480 243.050 10.330 243.200 ;
        RECT 10.030 242.600 10.330 243.050 ;
        RECT 6.480 242.450 10.330 242.600 ;
        RECT 10.030 242.000 10.330 242.450 ;
        RECT 6.530 241.450 10.330 242.000 ;
        RECT 10.780 241.450 10.930 249.650 ;
        RECT 11.380 241.450 11.530 249.650 ;
        RECT 11.980 241.450 12.130 249.650 ;
        RECT 12.580 241.450 12.730 249.650 ;
        RECT 13.180 241.450 13.330 249.650 ;
        RECT 13.780 241.450 13.930 249.650 ;
        RECT 14.380 241.450 15.080 258.550 ;
        RECT 15.530 250.350 15.680 258.550 ;
        RECT 16.130 250.350 16.280 258.550 ;
        RECT 16.730 250.350 16.880 258.550 ;
        RECT 17.330 250.350 17.480 258.550 ;
        RECT 17.930 250.350 18.080 258.550 ;
        RECT 18.530 250.350 18.680 258.550 ;
        RECT 19.130 258.000 22.930 258.550 ;
        RECT 26.530 258.550 42.930 258.600 ;
        RECT 26.530 258.000 30.330 258.550 ;
        RECT 19.130 257.550 19.430 258.000 ;
        RECT 30.030 257.550 30.330 258.000 ;
        RECT 19.130 257.400 22.980 257.550 ;
        RECT 26.480 257.400 30.330 257.550 ;
        RECT 19.130 256.950 19.430 257.400 ;
        RECT 30.030 256.950 30.330 257.400 ;
        RECT 19.130 256.800 22.980 256.950 ;
        RECT 26.480 256.800 30.330 256.950 ;
        RECT 19.130 256.350 19.430 256.800 ;
        RECT 30.030 256.350 30.330 256.800 ;
        RECT 19.130 256.200 22.980 256.350 ;
        RECT 26.480 256.200 30.330 256.350 ;
        RECT 19.130 255.750 19.430 256.200 ;
        RECT 30.030 255.750 30.330 256.200 ;
        RECT 19.130 255.600 22.980 255.750 ;
        RECT 26.480 255.600 30.330 255.750 ;
        RECT 19.130 255.150 19.430 255.600 ;
        RECT 30.030 255.150 30.330 255.600 ;
        RECT 19.130 255.000 22.980 255.150 ;
        RECT 26.480 255.000 30.330 255.150 ;
        RECT 19.130 254.550 19.430 255.000 ;
        RECT 30.030 254.550 30.330 255.000 ;
        RECT 19.130 254.400 22.980 254.550 ;
        RECT 26.480 254.400 30.330 254.550 ;
        RECT 19.130 253.950 19.430 254.400 ;
        RECT 30.030 253.950 30.330 254.400 ;
        RECT 19.130 253.800 22.980 253.950 ;
        RECT 26.480 253.800 30.330 253.950 ;
        RECT 19.130 253.350 19.430 253.800 ;
        RECT 30.030 253.350 30.330 253.800 ;
        RECT 19.130 253.200 22.980 253.350 ;
        RECT 26.480 253.200 30.330 253.350 ;
        RECT 19.130 252.750 19.430 253.200 ;
        RECT 19.130 252.600 22.980 252.750 ;
        RECT 19.130 252.150 19.430 252.600 ;
        RECT 19.130 252.000 22.980 252.150 ;
        RECT 19.130 251.550 19.430 252.000 ;
        RECT 19.130 251.400 22.980 251.550 ;
        RECT 19.130 250.950 19.430 251.400 ;
        RECT 19.130 250.800 22.980 250.950 ;
        RECT 19.130 250.350 19.430 250.800 ;
        RECT 15.530 241.450 15.680 249.650 ;
        RECT 16.130 241.450 16.280 249.650 ;
        RECT 16.730 241.450 16.880 249.650 ;
        RECT 17.330 241.450 17.480 249.650 ;
        RECT 17.930 241.450 18.080 249.650 ;
        RECT 18.530 241.450 18.680 249.650 ;
        RECT 19.130 249.200 19.430 249.650 ;
        RECT 19.130 249.050 22.980 249.200 ;
        RECT 19.130 248.600 19.430 249.050 ;
        RECT 19.130 248.450 22.980 248.600 ;
        RECT 19.130 248.000 19.430 248.450 ;
        RECT 19.130 247.850 22.980 248.000 ;
        RECT 19.130 247.400 19.430 247.850 ;
        RECT 19.130 247.250 22.980 247.400 ;
        RECT 19.130 246.800 19.430 247.250 ;
        RECT 23.830 246.800 25.630 253.200 ;
        RECT 30.030 252.750 30.330 253.200 ;
        RECT 26.480 252.600 30.330 252.750 ;
        RECT 30.030 252.150 30.330 252.600 ;
        RECT 26.480 252.000 30.330 252.150 ;
        RECT 30.030 251.550 30.330 252.000 ;
        RECT 26.480 251.400 30.330 251.550 ;
        RECT 30.030 250.950 30.330 251.400 ;
        RECT 26.480 250.800 30.330 250.950 ;
        RECT 30.030 250.350 30.330 250.800 ;
        RECT 30.780 250.350 30.930 258.550 ;
        RECT 31.380 250.350 31.530 258.550 ;
        RECT 31.980 250.350 32.130 258.550 ;
        RECT 32.580 250.350 32.730 258.550 ;
        RECT 33.180 250.350 33.330 258.550 ;
        RECT 33.780 250.350 33.930 258.550 ;
        RECT 30.030 249.200 30.330 249.650 ;
        RECT 26.480 249.050 30.330 249.200 ;
        RECT 30.030 248.600 30.330 249.050 ;
        RECT 26.480 248.450 30.330 248.600 ;
        RECT 30.030 248.000 30.330 248.450 ;
        RECT 26.480 247.850 30.330 248.000 ;
        RECT 30.030 247.400 30.330 247.850 ;
        RECT 26.480 247.250 30.330 247.400 ;
        RECT 30.030 246.800 30.330 247.250 ;
        RECT 19.130 246.650 22.980 246.800 ;
        RECT 26.480 246.650 30.330 246.800 ;
        RECT 19.130 246.200 19.430 246.650 ;
        RECT 30.030 246.200 30.330 246.650 ;
        RECT 19.130 246.050 22.980 246.200 ;
        RECT 26.480 246.050 30.330 246.200 ;
        RECT 19.130 245.600 19.430 246.050 ;
        RECT 30.030 245.600 30.330 246.050 ;
        RECT 19.130 245.450 22.980 245.600 ;
        RECT 26.480 245.450 30.330 245.600 ;
        RECT 19.130 245.000 19.430 245.450 ;
        RECT 30.030 245.000 30.330 245.450 ;
        RECT 19.130 244.850 22.980 245.000 ;
        RECT 26.480 244.850 30.330 245.000 ;
        RECT 19.130 244.400 19.430 244.850 ;
        RECT 30.030 244.400 30.330 244.850 ;
        RECT 19.130 244.250 22.980 244.400 ;
        RECT 26.480 244.250 30.330 244.400 ;
        RECT 19.130 243.800 19.430 244.250 ;
        RECT 30.030 243.800 30.330 244.250 ;
        RECT 19.130 243.650 22.980 243.800 ;
        RECT 26.480 243.650 30.330 243.800 ;
        RECT 19.130 243.200 19.430 243.650 ;
        RECT 30.030 243.200 30.330 243.650 ;
        RECT 19.130 243.050 22.980 243.200 ;
        RECT 26.480 243.050 30.330 243.200 ;
        RECT 19.130 242.600 19.430 243.050 ;
        RECT 30.030 242.600 30.330 243.050 ;
        RECT 19.130 242.450 22.980 242.600 ;
        RECT 26.480 242.450 30.330 242.600 ;
        RECT 19.130 242.000 19.430 242.450 ;
        RECT 30.030 242.000 30.330 242.450 ;
        RECT 19.130 241.450 22.930 242.000 ;
        RECT 6.530 241.400 22.930 241.450 ;
        RECT 26.530 241.450 30.330 242.000 ;
        RECT 30.780 241.450 30.930 249.650 ;
        RECT 31.380 241.450 31.530 249.650 ;
        RECT 31.980 241.450 32.130 249.650 ;
        RECT 32.580 241.450 32.730 249.650 ;
        RECT 33.180 241.450 33.330 249.650 ;
        RECT 33.780 241.450 33.930 249.650 ;
        RECT 34.380 241.450 35.080 258.550 ;
        RECT 35.530 250.350 35.680 258.550 ;
        RECT 36.130 250.350 36.280 258.550 ;
        RECT 36.730 250.350 36.880 258.550 ;
        RECT 37.330 250.350 37.480 258.550 ;
        RECT 37.930 250.350 38.080 258.550 ;
        RECT 38.530 250.350 38.680 258.550 ;
        RECT 39.130 258.000 42.930 258.550 ;
        RECT 46.530 258.550 62.930 258.600 ;
        RECT 46.530 258.000 50.330 258.550 ;
        RECT 39.130 257.550 39.430 258.000 ;
        RECT 50.030 257.550 50.330 258.000 ;
        RECT 39.130 257.400 42.980 257.550 ;
        RECT 46.480 257.400 50.330 257.550 ;
        RECT 39.130 256.950 39.430 257.400 ;
        RECT 50.030 256.950 50.330 257.400 ;
        RECT 39.130 256.800 42.980 256.950 ;
        RECT 46.480 256.800 50.330 256.950 ;
        RECT 39.130 256.350 39.430 256.800 ;
        RECT 50.030 256.350 50.330 256.800 ;
        RECT 39.130 256.200 42.980 256.350 ;
        RECT 46.480 256.200 50.330 256.350 ;
        RECT 39.130 255.750 39.430 256.200 ;
        RECT 50.030 255.750 50.330 256.200 ;
        RECT 39.130 255.600 42.980 255.750 ;
        RECT 46.480 255.600 50.330 255.750 ;
        RECT 39.130 255.150 39.430 255.600 ;
        RECT 50.030 255.150 50.330 255.600 ;
        RECT 39.130 255.000 42.980 255.150 ;
        RECT 46.480 255.000 50.330 255.150 ;
        RECT 39.130 254.550 39.430 255.000 ;
        RECT 50.030 254.550 50.330 255.000 ;
        RECT 39.130 254.400 42.980 254.550 ;
        RECT 46.480 254.400 50.330 254.550 ;
        RECT 39.130 253.950 39.430 254.400 ;
        RECT 50.030 253.950 50.330 254.400 ;
        RECT 39.130 253.800 42.980 253.950 ;
        RECT 46.480 253.800 50.330 253.950 ;
        RECT 39.130 253.350 39.430 253.800 ;
        RECT 50.030 253.350 50.330 253.800 ;
        RECT 39.130 253.200 42.980 253.350 ;
        RECT 46.480 253.200 50.330 253.350 ;
        RECT 39.130 252.750 39.430 253.200 ;
        RECT 39.130 252.600 42.980 252.750 ;
        RECT 39.130 252.150 39.430 252.600 ;
        RECT 39.130 252.000 42.980 252.150 ;
        RECT 39.130 251.550 39.430 252.000 ;
        RECT 39.130 251.400 42.980 251.550 ;
        RECT 39.130 250.950 39.430 251.400 ;
        RECT 39.130 250.800 42.980 250.950 ;
        RECT 39.130 250.350 39.430 250.800 ;
        RECT 35.530 241.450 35.680 249.650 ;
        RECT 36.130 241.450 36.280 249.650 ;
        RECT 36.730 241.450 36.880 249.650 ;
        RECT 37.330 241.450 37.480 249.650 ;
        RECT 37.930 241.450 38.080 249.650 ;
        RECT 38.530 241.450 38.680 249.650 ;
        RECT 39.130 249.200 39.430 249.650 ;
        RECT 39.130 249.050 42.980 249.200 ;
        RECT 39.130 248.600 39.430 249.050 ;
        RECT 39.130 248.450 42.980 248.600 ;
        RECT 39.130 248.000 39.430 248.450 ;
        RECT 39.130 247.850 42.980 248.000 ;
        RECT 39.130 247.400 39.430 247.850 ;
        RECT 39.130 247.250 42.980 247.400 ;
        RECT 39.130 246.800 39.430 247.250 ;
        RECT 43.830 246.800 45.630 253.200 ;
        RECT 50.030 252.750 50.330 253.200 ;
        RECT 46.480 252.600 50.330 252.750 ;
        RECT 50.030 252.150 50.330 252.600 ;
        RECT 46.480 252.000 50.330 252.150 ;
        RECT 50.030 251.550 50.330 252.000 ;
        RECT 46.480 251.400 50.330 251.550 ;
        RECT 50.030 250.950 50.330 251.400 ;
        RECT 46.480 250.800 50.330 250.950 ;
        RECT 50.030 250.350 50.330 250.800 ;
        RECT 50.780 250.350 50.930 258.550 ;
        RECT 51.380 250.350 51.530 258.550 ;
        RECT 51.980 250.350 52.130 258.550 ;
        RECT 52.580 250.350 52.730 258.550 ;
        RECT 53.180 250.350 53.330 258.550 ;
        RECT 53.780 250.350 53.930 258.550 ;
        RECT 50.030 249.200 50.330 249.650 ;
        RECT 46.480 249.050 50.330 249.200 ;
        RECT 50.030 248.600 50.330 249.050 ;
        RECT 46.480 248.450 50.330 248.600 ;
        RECT 50.030 248.000 50.330 248.450 ;
        RECT 46.480 247.850 50.330 248.000 ;
        RECT 50.030 247.400 50.330 247.850 ;
        RECT 46.480 247.250 50.330 247.400 ;
        RECT 50.030 246.800 50.330 247.250 ;
        RECT 39.130 246.650 42.980 246.800 ;
        RECT 46.480 246.650 50.330 246.800 ;
        RECT 39.130 246.200 39.430 246.650 ;
        RECT 50.030 246.200 50.330 246.650 ;
        RECT 39.130 246.050 42.980 246.200 ;
        RECT 46.480 246.050 50.330 246.200 ;
        RECT 39.130 245.600 39.430 246.050 ;
        RECT 50.030 245.600 50.330 246.050 ;
        RECT 39.130 245.450 42.980 245.600 ;
        RECT 46.480 245.450 50.330 245.600 ;
        RECT 39.130 245.000 39.430 245.450 ;
        RECT 50.030 245.000 50.330 245.450 ;
        RECT 39.130 244.850 42.980 245.000 ;
        RECT 46.480 244.850 50.330 245.000 ;
        RECT 39.130 244.400 39.430 244.850 ;
        RECT 50.030 244.400 50.330 244.850 ;
        RECT 39.130 244.250 42.980 244.400 ;
        RECT 46.480 244.250 50.330 244.400 ;
        RECT 39.130 243.800 39.430 244.250 ;
        RECT 50.030 243.800 50.330 244.250 ;
        RECT 39.130 243.650 42.980 243.800 ;
        RECT 46.480 243.650 50.330 243.800 ;
        RECT 39.130 243.200 39.430 243.650 ;
        RECT 50.030 243.200 50.330 243.650 ;
        RECT 39.130 243.050 42.980 243.200 ;
        RECT 46.480 243.050 50.330 243.200 ;
        RECT 39.130 242.600 39.430 243.050 ;
        RECT 50.030 242.600 50.330 243.050 ;
        RECT 39.130 242.450 42.980 242.600 ;
        RECT 46.480 242.450 50.330 242.600 ;
        RECT 39.130 242.000 39.430 242.450 ;
        RECT 50.030 242.000 50.330 242.450 ;
        RECT 39.130 241.450 42.930 242.000 ;
        RECT 26.530 241.400 42.930 241.450 ;
        RECT 46.530 241.450 50.330 242.000 ;
        RECT 50.780 241.450 50.930 249.650 ;
        RECT 51.380 241.450 51.530 249.650 ;
        RECT 51.980 241.450 52.130 249.650 ;
        RECT 52.580 241.450 52.730 249.650 ;
        RECT 53.180 241.450 53.330 249.650 ;
        RECT 53.780 241.450 53.930 249.650 ;
        RECT 54.380 241.450 55.080 258.550 ;
        RECT 55.530 250.350 55.680 258.550 ;
        RECT 56.130 250.350 56.280 258.550 ;
        RECT 56.730 250.350 56.880 258.550 ;
        RECT 57.330 250.350 57.480 258.550 ;
        RECT 57.930 250.350 58.080 258.550 ;
        RECT 58.530 250.350 58.680 258.550 ;
        RECT 59.130 258.000 62.930 258.550 ;
        RECT 66.530 258.550 82.930 258.600 ;
        RECT 66.530 258.000 70.330 258.550 ;
        RECT 59.130 257.550 59.430 258.000 ;
        RECT 70.030 257.550 70.330 258.000 ;
        RECT 59.130 257.400 62.980 257.550 ;
        RECT 66.480 257.400 70.330 257.550 ;
        RECT 59.130 256.950 59.430 257.400 ;
        RECT 70.030 256.950 70.330 257.400 ;
        RECT 59.130 256.800 62.980 256.950 ;
        RECT 66.480 256.800 70.330 256.950 ;
        RECT 59.130 256.350 59.430 256.800 ;
        RECT 70.030 256.350 70.330 256.800 ;
        RECT 59.130 256.200 62.980 256.350 ;
        RECT 66.480 256.200 70.330 256.350 ;
        RECT 59.130 255.750 59.430 256.200 ;
        RECT 70.030 255.750 70.330 256.200 ;
        RECT 59.130 255.600 62.980 255.750 ;
        RECT 66.480 255.600 70.330 255.750 ;
        RECT 59.130 255.150 59.430 255.600 ;
        RECT 70.030 255.150 70.330 255.600 ;
        RECT 59.130 255.000 62.980 255.150 ;
        RECT 66.480 255.000 70.330 255.150 ;
        RECT 59.130 254.550 59.430 255.000 ;
        RECT 70.030 254.550 70.330 255.000 ;
        RECT 59.130 254.400 62.980 254.550 ;
        RECT 66.480 254.400 70.330 254.550 ;
        RECT 59.130 253.950 59.430 254.400 ;
        RECT 70.030 253.950 70.330 254.400 ;
        RECT 59.130 253.800 62.980 253.950 ;
        RECT 66.480 253.800 70.330 253.950 ;
        RECT 59.130 253.350 59.430 253.800 ;
        RECT 70.030 253.350 70.330 253.800 ;
        RECT 59.130 253.200 62.980 253.350 ;
        RECT 66.480 253.200 70.330 253.350 ;
        RECT 59.130 252.750 59.430 253.200 ;
        RECT 59.130 252.600 62.980 252.750 ;
        RECT 59.130 252.150 59.430 252.600 ;
        RECT 59.130 252.000 62.980 252.150 ;
        RECT 59.130 251.550 59.430 252.000 ;
        RECT 59.130 251.400 62.980 251.550 ;
        RECT 59.130 250.950 59.430 251.400 ;
        RECT 59.130 250.800 62.980 250.950 ;
        RECT 59.130 250.350 59.430 250.800 ;
        RECT 55.530 241.450 55.680 249.650 ;
        RECT 56.130 241.450 56.280 249.650 ;
        RECT 56.730 241.450 56.880 249.650 ;
        RECT 57.330 241.450 57.480 249.650 ;
        RECT 57.930 241.450 58.080 249.650 ;
        RECT 58.530 241.450 58.680 249.650 ;
        RECT 59.130 249.200 59.430 249.650 ;
        RECT 59.130 249.050 62.980 249.200 ;
        RECT 59.130 248.600 59.430 249.050 ;
        RECT 59.130 248.450 62.980 248.600 ;
        RECT 59.130 248.000 59.430 248.450 ;
        RECT 59.130 247.850 62.980 248.000 ;
        RECT 59.130 247.400 59.430 247.850 ;
        RECT 59.130 247.250 62.980 247.400 ;
        RECT 59.130 246.800 59.430 247.250 ;
        RECT 63.830 246.800 65.630 253.200 ;
        RECT 70.030 252.750 70.330 253.200 ;
        RECT 66.480 252.600 70.330 252.750 ;
        RECT 70.030 252.150 70.330 252.600 ;
        RECT 66.480 252.000 70.330 252.150 ;
        RECT 70.030 251.550 70.330 252.000 ;
        RECT 66.480 251.400 70.330 251.550 ;
        RECT 70.030 250.950 70.330 251.400 ;
        RECT 66.480 250.800 70.330 250.950 ;
        RECT 70.030 250.350 70.330 250.800 ;
        RECT 70.780 250.350 70.930 258.550 ;
        RECT 71.380 250.350 71.530 258.550 ;
        RECT 71.980 250.350 72.130 258.550 ;
        RECT 72.580 250.350 72.730 258.550 ;
        RECT 73.180 250.350 73.330 258.550 ;
        RECT 73.780 250.350 73.930 258.550 ;
        RECT 70.030 249.200 70.330 249.650 ;
        RECT 66.480 249.050 70.330 249.200 ;
        RECT 70.030 248.600 70.330 249.050 ;
        RECT 66.480 248.450 70.330 248.600 ;
        RECT 70.030 248.000 70.330 248.450 ;
        RECT 66.480 247.850 70.330 248.000 ;
        RECT 70.030 247.400 70.330 247.850 ;
        RECT 66.480 247.250 70.330 247.400 ;
        RECT 70.030 246.800 70.330 247.250 ;
        RECT 59.130 246.650 62.980 246.800 ;
        RECT 66.480 246.650 70.330 246.800 ;
        RECT 59.130 246.200 59.430 246.650 ;
        RECT 70.030 246.200 70.330 246.650 ;
        RECT 59.130 246.050 62.980 246.200 ;
        RECT 66.480 246.050 70.330 246.200 ;
        RECT 59.130 245.600 59.430 246.050 ;
        RECT 70.030 245.600 70.330 246.050 ;
        RECT 59.130 245.450 62.980 245.600 ;
        RECT 66.480 245.450 70.330 245.600 ;
        RECT 59.130 245.000 59.430 245.450 ;
        RECT 70.030 245.000 70.330 245.450 ;
        RECT 59.130 244.850 62.980 245.000 ;
        RECT 66.480 244.850 70.330 245.000 ;
        RECT 59.130 244.400 59.430 244.850 ;
        RECT 70.030 244.400 70.330 244.850 ;
        RECT 59.130 244.250 62.980 244.400 ;
        RECT 66.480 244.250 70.330 244.400 ;
        RECT 59.130 243.800 59.430 244.250 ;
        RECT 70.030 243.800 70.330 244.250 ;
        RECT 59.130 243.650 62.980 243.800 ;
        RECT 66.480 243.650 70.330 243.800 ;
        RECT 59.130 243.200 59.430 243.650 ;
        RECT 70.030 243.200 70.330 243.650 ;
        RECT 59.130 243.050 62.980 243.200 ;
        RECT 66.480 243.050 70.330 243.200 ;
        RECT 59.130 242.600 59.430 243.050 ;
        RECT 70.030 242.600 70.330 243.050 ;
        RECT 59.130 242.450 62.980 242.600 ;
        RECT 66.480 242.450 70.330 242.600 ;
        RECT 59.130 242.000 59.430 242.450 ;
        RECT 70.030 242.000 70.330 242.450 ;
        RECT 59.130 241.450 62.930 242.000 ;
        RECT 46.530 241.400 62.930 241.450 ;
        RECT 66.530 241.450 70.330 242.000 ;
        RECT 70.780 241.450 70.930 249.650 ;
        RECT 71.380 241.450 71.530 249.650 ;
        RECT 71.980 241.450 72.130 249.650 ;
        RECT 72.580 241.450 72.730 249.650 ;
        RECT 73.180 241.450 73.330 249.650 ;
        RECT 73.780 241.450 73.930 249.650 ;
        RECT 74.380 241.450 75.080 258.550 ;
        RECT 75.530 250.350 75.680 258.550 ;
        RECT 76.130 250.350 76.280 258.550 ;
        RECT 76.730 250.350 76.880 258.550 ;
        RECT 77.330 250.350 77.480 258.550 ;
        RECT 77.930 250.350 78.080 258.550 ;
        RECT 78.530 250.350 78.680 258.550 ;
        RECT 79.130 258.000 82.930 258.550 ;
        RECT 86.530 258.550 102.930 258.600 ;
        RECT 86.530 258.000 90.330 258.550 ;
        RECT 79.130 257.550 79.430 258.000 ;
        RECT 90.030 257.550 90.330 258.000 ;
        RECT 79.130 257.400 82.980 257.550 ;
        RECT 86.480 257.400 90.330 257.550 ;
        RECT 79.130 256.950 79.430 257.400 ;
        RECT 90.030 256.950 90.330 257.400 ;
        RECT 79.130 256.800 82.980 256.950 ;
        RECT 86.480 256.800 90.330 256.950 ;
        RECT 79.130 256.350 79.430 256.800 ;
        RECT 90.030 256.350 90.330 256.800 ;
        RECT 79.130 256.200 82.980 256.350 ;
        RECT 86.480 256.200 90.330 256.350 ;
        RECT 79.130 255.750 79.430 256.200 ;
        RECT 90.030 255.750 90.330 256.200 ;
        RECT 79.130 255.600 82.980 255.750 ;
        RECT 86.480 255.600 90.330 255.750 ;
        RECT 79.130 255.150 79.430 255.600 ;
        RECT 90.030 255.150 90.330 255.600 ;
        RECT 79.130 255.000 82.980 255.150 ;
        RECT 86.480 255.000 90.330 255.150 ;
        RECT 79.130 254.550 79.430 255.000 ;
        RECT 90.030 254.550 90.330 255.000 ;
        RECT 79.130 254.400 82.980 254.550 ;
        RECT 86.480 254.400 90.330 254.550 ;
        RECT 79.130 253.950 79.430 254.400 ;
        RECT 90.030 253.950 90.330 254.400 ;
        RECT 79.130 253.800 82.980 253.950 ;
        RECT 86.480 253.800 90.330 253.950 ;
        RECT 79.130 253.350 79.430 253.800 ;
        RECT 90.030 253.350 90.330 253.800 ;
        RECT 79.130 253.200 82.980 253.350 ;
        RECT 86.480 253.200 90.330 253.350 ;
        RECT 79.130 252.750 79.430 253.200 ;
        RECT 79.130 252.600 82.980 252.750 ;
        RECT 79.130 252.150 79.430 252.600 ;
        RECT 79.130 252.000 82.980 252.150 ;
        RECT 79.130 251.550 79.430 252.000 ;
        RECT 79.130 251.400 82.980 251.550 ;
        RECT 79.130 250.950 79.430 251.400 ;
        RECT 79.130 250.800 82.980 250.950 ;
        RECT 79.130 250.350 79.430 250.800 ;
        RECT 75.530 241.450 75.680 249.650 ;
        RECT 76.130 241.450 76.280 249.650 ;
        RECT 76.730 241.450 76.880 249.650 ;
        RECT 77.330 241.450 77.480 249.650 ;
        RECT 77.930 241.450 78.080 249.650 ;
        RECT 78.530 241.450 78.680 249.650 ;
        RECT 79.130 249.200 79.430 249.650 ;
        RECT 79.130 249.050 82.980 249.200 ;
        RECT 79.130 248.600 79.430 249.050 ;
        RECT 79.130 248.450 82.980 248.600 ;
        RECT 79.130 248.000 79.430 248.450 ;
        RECT 79.130 247.850 82.980 248.000 ;
        RECT 79.130 247.400 79.430 247.850 ;
        RECT 79.130 247.250 82.980 247.400 ;
        RECT 79.130 246.800 79.430 247.250 ;
        RECT 83.830 246.800 85.630 253.200 ;
        RECT 90.030 252.750 90.330 253.200 ;
        RECT 86.480 252.600 90.330 252.750 ;
        RECT 90.030 252.150 90.330 252.600 ;
        RECT 86.480 252.000 90.330 252.150 ;
        RECT 90.030 251.550 90.330 252.000 ;
        RECT 86.480 251.400 90.330 251.550 ;
        RECT 90.030 250.950 90.330 251.400 ;
        RECT 86.480 250.800 90.330 250.950 ;
        RECT 90.030 250.350 90.330 250.800 ;
        RECT 90.780 250.350 90.930 258.550 ;
        RECT 91.380 250.350 91.530 258.550 ;
        RECT 91.980 250.350 92.130 258.550 ;
        RECT 92.580 250.350 92.730 258.550 ;
        RECT 93.180 250.350 93.330 258.550 ;
        RECT 93.780 250.350 93.930 258.550 ;
        RECT 90.030 249.200 90.330 249.650 ;
        RECT 86.480 249.050 90.330 249.200 ;
        RECT 90.030 248.600 90.330 249.050 ;
        RECT 86.480 248.450 90.330 248.600 ;
        RECT 90.030 248.000 90.330 248.450 ;
        RECT 86.480 247.850 90.330 248.000 ;
        RECT 90.030 247.400 90.330 247.850 ;
        RECT 86.480 247.250 90.330 247.400 ;
        RECT 90.030 246.800 90.330 247.250 ;
        RECT 79.130 246.650 82.980 246.800 ;
        RECT 86.480 246.650 90.330 246.800 ;
        RECT 79.130 246.200 79.430 246.650 ;
        RECT 90.030 246.200 90.330 246.650 ;
        RECT 79.130 246.050 82.980 246.200 ;
        RECT 86.480 246.050 90.330 246.200 ;
        RECT 79.130 245.600 79.430 246.050 ;
        RECT 90.030 245.600 90.330 246.050 ;
        RECT 79.130 245.450 82.980 245.600 ;
        RECT 86.480 245.450 90.330 245.600 ;
        RECT 79.130 245.000 79.430 245.450 ;
        RECT 90.030 245.000 90.330 245.450 ;
        RECT 79.130 244.850 82.980 245.000 ;
        RECT 86.480 244.850 90.330 245.000 ;
        RECT 79.130 244.400 79.430 244.850 ;
        RECT 90.030 244.400 90.330 244.850 ;
        RECT 79.130 244.250 82.980 244.400 ;
        RECT 86.480 244.250 90.330 244.400 ;
        RECT 79.130 243.800 79.430 244.250 ;
        RECT 90.030 243.800 90.330 244.250 ;
        RECT 79.130 243.650 82.980 243.800 ;
        RECT 86.480 243.650 90.330 243.800 ;
        RECT 79.130 243.200 79.430 243.650 ;
        RECT 90.030 243.200 90.330 243.650 ;
        RECT 79.130 243.050 82.980 243.200 ;
        RECT 86.480 243.050 90.330 243.200 ;
        RECT 79.130 242.600 79.430 243.050 ;
        RECT 90.030 242.600 90.330 243.050 ;
        RECT 79.130 242.450 82.980 242.600 ;
        RECT 86.480 242.450 90.330 242.600 ;
        RECT 79.130 242.000 79.430 242.450 ;
        RECT 90.030 242.000 90.330 242.450 ;
        RECT 79.130 241.450 82.930 242.000 ;
        RECT 66.530 241.400 82.930 241.450 ;
        RECT 86.530 241.450 90.330 242.000 ;
        RECT 90.780 241.450 90.930 249.650 ;
        RECT 91.380 241.450 91.530 249.650 ;
        RECT 91.980 241.450 92.130 249.650 ;
        RECT 92.580 241.450 92.730 249.650 ;
        RECT 93.180 241.450 93.330 249.650 ;
        RECT 93.780 241.450 93.930 249.650 ;
        RECT 94.380 241.450 95.080 258.550 ;
        RECT 95.530 250.350 95.680 258.550 ;
        RECT 96.130 250.350 96.280 258.550 ;
        RECT 96.730 250.350 96.880 258.550 ;
        RECT 97.330 250.350 97.480 258.550 ;
        RECT 97.930 250.350 98.080 258.550 ;
        RECT 98.530 250.350 98.680 258.550 ;
        RECT 99.130 258.000 102.930 258.550 ;
        RECT 99.130 257.550 99.430 258.000 ;
        RECT 99.130 257.400 102.980 257.550 ;
        RECT 99.130 256.950 99.430 257.400 ;
        RECT 99.130 256.800 102.980 256.950 ;
        RECT 99.130 256.350 99.430 256.800 ;
        RECT 99.130 256.200 102.980 256.350 ;
        RECT 99.130 255.750 99.430 256.200 ;
        RECT 99.130 255.600 102.980 255.750 ;
        RECT 99.130 255.150 99.430 255.600 ;
        RECT 99.130 255.000 102.980 255.150 ;
        RECT 99.130 254.550 99.430 255.000 ;
        RECT 99.130 254.400 102.980 254.550 ;
        RECT 99.130 253.950 99.430 254.400 ;
        RECT 99.130 253.800 102.980 253.950 ;
        RECT 99.130 253.350 99.430 253.800 ;
        RECT 99.130 253.200 102.980 253.350 ;
        RECT 99.130 252.750 99.430 253.200 ;
        RECT 99.130 252.600 102.980 252.750 ;
        RECT 99.130 252.150 99.430 252.600 ;
        RECT 99.130 252.000 102.980 252.150 ;
        RECT 99.130 251.550 99.430 252.000 ;
        RECT 99.130 251.400 102.980 251.550 ;
        RECT 99.130 250.950 99.430 251.400 ;
        RECT 99.130 250.800 102.980 250.950 ;
        RECT 99.130 250.350 99.430 250.800 ;
        RECT 95.530 241.450 95.680 249.650 ;
        RECT 96.130 241.450 96.280 249.650 ;
        RECT 96.730 241.450 96.880 249.650 ;
        RECT 97.330 241.450 97.480 249.650 ;
        RECT 97.930 241.450 98.080 249.650 ;
        RECT 98.530 241.450 98.680 249.650 ;
        RECT 99.130 249.200 99.430 249.650 ;
        RECT 99.130 249.050 102.980 249.200 ;
        RECT 99.130 248.600 99.430 249.050 ;
        RECT 99.130 248.450 102.980 248.600 ;
        RECT 99.130 248.000 99.430 248.450 ;
        RECT 99.130 247.850 102.980 248.000 ;
        RECT 99.130 247.400 99.430 247.850 ;
        RECT 99.130 247.250 102.980 247.400 ;
        RECT 99.130 246.800 99.430 247.250 ;
        RECT 103.830 246.800 104.730 253.200 ;
        RECT 109.850 249.640 111.850 250.915 ;
        RECT 99.130 246.650 102.980 246.800 ;
        RECT 99.130 246.200 99.430 246.650 ;
        RECT 99.130 246.050 102.980 246.200 ;
        RECT 99.130 245.600 99.430 246.050 ;
        RECT 99.130 245.450 102.980 245.600 ;
        RECT 99.130 245.000 99.430 245.450 ;
        RECT 99.130 244.850 102.980 245.000 ;
        RECT 99.130 244.400 99.430 244.850 ;
        RECT 99.130 244.250 102.980 244.400 ;
        RECT 99.130 243.800 99.430 244.250 ;
        RECT 99.130 243.650 102.980 243.800 ;
        RECT 99.130 243.200 99.430 243.650 ;
        RECT 99.130 243.050 102.980 243.200 ;
        RECT 99.130 242.600 99.430 243.050 ;
        RECT 99.130 242.450 102.980 242.600 ;
        RECT 99.130 242.000 99.430 242.450 ;
        RECT 99.130 241.450 102.930 242.000 ;
        RECT 86.530 241.400 102.930 241.450 ;
        RECT 9.630 240.900 19.830 241.400 ;
        RECT 29.630 240.900 39.830 241.400 ;
        RECT 49.630 240.900 59.830 241.400 ;
        RECT 69.630 240.900 79.830 241.400 ;
        RECT 89.630 240.900 99.830 241.400 ;
        RECT 11.530 239.100 17.930 240.900 ;
        RECT 31.530 239.100 37.930 240.900 ;
        RECT 51.530 239.100 57.930 240.900 ;
        RECT 71.530 239.100 77.930 240.900 ;
        RECT 91.530 239.100 97.930 240.900 ;
        RECT 9.630 238.600 19.830 239.100 ;
        RECT 29.630 238.600 39.830 239.100 ;
        RECT 49.630 238.600 59.830 239.100 ;
        RECT 69.630 238.600 79.830 239.100 ;
        RECT 89.630 238.600 99.830 239.100 ;
        RECT 6.530 238.550 22.930 238.600 ;
        RECT 6.530 238.000 10.330 238.550 ;
        RECT 10.030 237.550 10.330 238.000 ;
        RECT 6.480 237.400 10.330 237.550 ;
        RECT 10.030 236.950 10.330 237.400 ;
        RECT 6.480 236.800 10.330 236.950 ;
        RECT 10.030 236.350 10.330 236.800 ;
        RECT 6.480 236.200 10.330 236.350 ;
        RECT 10.030 235.750 10.330 236.200 ;
        RECT 6.480 235.600 10.330 235.750 ;
        RECT 10.030 235.150 10.330 235.600 ;
        RECT 6.480 235.000 10.330 235.150 ;
        RECT 10.030 234.550 10.330 235.000 ;
        RECT 6.480 234.400 10.330 234.550 ;
        RECT 10.030 233.950 10.330 234.400 ;
        RECT 6.480 233.800 10.330 233.950 ;
        RECT 10.030 233.350 10.330 233.800 ;
        RECT 6.480 233.200 10.330 233.350 ;
        RECT 4.730 226.800 5.630 233.200 ;
        RECT 10.030 232.750 10.330 233.200 ;
        RECT 6.480 232.600 10.330 232.750 ;
        RECT 10.030 232.150 10.330 232.600 ;
        RECT 6.480 232.000 10.330 232.150 ;
        RECT 10.030 231.550 10.330 232.000 ;
        RECT 6.480 231.400 10.330 231.550 ;
        RECT 10.030 230.950 10.330 231.400 ;
        RECT 6.480 230.800 10.330 230.950 ;
        RECT 10.030 230.350 10.330 230.800 ;
        RECT 10.780 230.350 10.930 238.550 ;
        RECT 11.380 230.350 11.530 238.550 ;
        RECT 11.980 230.350 12.130 238.550 ;
        RECT 12.580 230.350 12.730 238.550 ;
        RECT 13.180 230.350 13.330 238.550 ;
        RECT 13.780 230.350 13.930 238.550 ;
        RECT 10.030 229.200 10.330 229.650 ;
        RECT 6.480 229.050 10.330 229.200 ;
        RECT 10.030 228.600 10.330 229.050 ;
        RECT 6.480 228.450 10.330 228.600 ;
        RECT 10.030 228.000 10.330 228.450 ;
        RECT 6.480 227.850 10.330 228.000 ;
        RECT 10.030 227.400 10.330 227.850 ;
        RECT 6.480 227.250 10.330 227.400 ;
        RECT 10.030 226.800 10.330 227.250 ;
        RECT 6.480 226.650 10.330 226.800 ;
        RECT 10.030 226.200 10.330 226.650 ;
        RECT 6.480 226.050 10.330 226.200 ;
        RECT 10.030 225.600 10.330 226.050 ;
        RECT 6.480 225.450 10.330 225.600 ;
        RECT 10.030 225.000 10.330 225.450 ;
        RECT 6.480 224.850 10.330 225.000 ;
        RECT 10.030 224.400 10.330 224.850 ;
        RECT 6.480 224.250 10.330 224.400 ;
        RECT 10.030 223.800 10.330 224.250 ;
        RECT 6.480 223.650 10.330 223.800 ;
        RECT 10.030 223.200 10.330 223.650 ;
        RECT 6.480 223.050 10.330 223.200 ;
        RECT 10.030 222.600 10.330 223.050 ;
        RECT 6.480 222.450 10.330 222.600 ;
        RECT 10.030 222.000 10.330 222.450 ;
        RECT 6.530 221.450 10.330 222.000 ;
        RECT 10.780 221.450 10.930 229.650 ;
        RECT 11.380 221.450 11.530 229.650 ;
        RECT 11.980 221.450 12.130 229.650 ;
        RECT 12.580 221.450 12.730 229.650 ;
        RECT 13.180 221.450 13.330 229.650 ;
        RECT 13.780 221.450 13.930 229.650 ;
        RECT 14.380 221.450 15.080 238.550 ;
        RECT 15.530 230.350 15.680 238.550 ;
        RECT 16.130 230.350 16.280 238.550 ;
        RECT 16.730 230.350 16.880 238.550 ;
        RECT 17.330 230.350 17.480 238.550 ;
        RECT 17.930 230.350 18.080 238.550 ;
        RECT 18.530 230.350 18.680 238.550 ;
        RECT 19.130 238.000 22.930 238.550 ;
        RECT 26.530 238.550 42.930 238.600 ;
        RECT 26.530 238.000 30.330 238.550 ;
        RECT 19.130 237.550 19.430 238.000 ;
        RECT 30.030 237.550 30.330 238.000 ;
        RECT 19.130 237.400 22.980 237.550 ;
        RECT 26.480 237.400 30.330 237.550 ;
        RECT 19.130 236.950 19.430 237.400 ;
        RECT 30.030 236.950 30.330 237.400 ;
        RECT 19.130 236.800 22.980 236.950 ;
        RECT 26.480 236.800 30.330 236.950 ;
        RECT 19.130 236.350 19.430 236.800 ;
        RECT 30.030 236.350 30.330 236.800 ;
        RECT 19.130 236.200 22.980 236.350 ;
        RECT 26.480 236.200 30.330 236.350 ;
        RECT 19.130 235.750 19.430 236.200 ;
        RECT 30.030 235.750 30.330 236.200 ;
        RECT 19.130 235.600 22.980 235.750 ;
        RECT 26.480 235.600 30.330 235.750 ;
        RECT 19.130 235.150 19.430 235.600 ;
        RECT 30.030 235.150 30.330 235.600 ;
        RECT 19.130 235.000 22.980 235.150 ;
        RECT 26.480 235.000 30.330 235.150 ;
        RECT 19.130 234.550 19.430 235.000 ;
        RECT 30.030 234.550 30.330 235.000 ;
        RECT 19.130 234.400 22.980 234.550 ;
        RECT 26.480 234.400 30.330 234.550 ;
        RECT 19.130 233.950 19.430 234.400 ;
        RECT 30.030 233.950 30.330 234.400 ;
        RECT 19.130 233.800 22.980 233.950 ;
        RECT 26.480 233.800 30.330 233.950 ;
        RECT 19.130 233.350 19.430 233.800 ;
        RECT 30.030 233.350 30.330 233.800 ;
        RECT 19.130 233.200 22.980 233.350 ;
        RECT 26.480 233.200 30.330 233.350 ;
        RECT 19.130 232.750 19.430 233.200 ;
        RECT 19.130 232.600 22.980 232.750 ;
        RECT 19.130 232.150 19.430 232.600 ;
        RECT 19.130 232.000 22.980 232.150 ;
        RECT 19.130 231.550 19.430 232.000 ;
        RECT 19.130 231.400 22.980 231.550 ;
        RECT 19.130 230.950 19.430 231.400 ;
        RECT 19.130 230.800 22.980 230.950 ;
        RECT 19.130 230.350 19.430 230.800 ;
        RECT 15.530 221.450 15.680 229.650 ;
        RECT 16.130 221.450 16.280 229.650 ;
        RECT 16.730 221.450 16.880 229.650 ;
        RECT 17.330 221.450 17.480 229.650 ;
        RECT 17.930 221.450 18.080 229.650 ;
        RECT 18.530 221.450 18.680 229.650 ;
        RECT 19.130 229.200 19.430 229.650 ;
        RECT 19.130 229.050 22.980 229.200 ;
        RECT 19.130 228.600 19.430 229.050 ;
        RECT 19.130 228.450 22.980 228.600 ;
        RECT 19.130 228.000 19.430 228.450 ;
        RECT 19.130 227.850 22.980 228.000 ;
        RECT 19.130 227.400 19.430 227.850 ;
        RECT 19.130 227.250 22.980 227.400 ;
        RECT 19.130 226.800 19.430 227.250 ;
        RECT 23.830 226.800 25.630 233.200 ;
        RECT 30.030 232.750 30.330 233.200 ;
        RECT 26.480 232.600 30.330 232.750 ;
        RECT 30.030 232.150 30.330 232.600 ;
        RECT 26.480 232.000 30.330 232.150 ;
        RECT 30.030 231.550 30.330 232.000 ;
        RECT 26.480 231.400 30.330 231.550 ;
        RECT 30.030 230.950 30.330 231.400 ;
        RECT 26.480 230.800 30.330 230.950 ;
        RECT 30.030 230.350 30.330 230.800 ;
        RECT 30.780 230.350 30.930 238.550 ;
        RECT 31.380 230.350 31.530 238.550 ;
        RECT 31.980 230.350 32.130 238.550 ;
        RECT 32.580 230.350 32.730 238.550 ;
        RECT 33.180 230.350 33.330 238.550 ;
        RECT 33.780 230.350 33.930 238.550 ;
        RECT 30.030 229.200 30.330 229.650 ;
        RECT 26.480 229.050 30.330 229.200 ;
        RECT 30.030 228.600 30.330 229.050 ;
        RECT 26.480 228.450 30.330 228.600 ;
        RECT 30.030 228.000 30.330 228.450 ;
        RECT 26.480 227.850 30.330 228.000 ;
        RECT 30.030 227.400 30.330 227.850 ;
        RECT 26.480 227.250 30.330 227.400 ;
        RECT 30.030 226.800 30.330 227.250 ;
        RECT 19.130 226.650 22.980 226.800 ;
        RECT 26.480 226.650 30.330 226.800 ;
        RECT 19.130 226.200 19.430 226.650 ;
        RECT 30.030 226.200 30.330 226.650 ;
        RECT 19.130 226.050 22.980 226.200 ;
        RECT 26.480 226.050 30.330 226.200 ;
        RECT 19.130 225.600 19.430 226.050 ;
        RECT 30.030 225.600 30.330 226.050 ;
        RECT 19.130 225.450 22.980 225.600 ;
        RECT 26.480 225.450 30.330 225.600 ;
        RECT 19.130 225.000 19.430 225.450 ;
        RECT 30.030 225.000 30.330 225.450 ;
        RECT 19.130 224.850 22.980 225.000 ;
        RECT 26.480 224.850 30.330 225.000 ;
        RECT 19.130 224.400 19.430 224.850 ;
        RECT 30.030 224.400 30.330 224.850 ;
        RECT 19.130 224.250 22.980 224.400 ;
        RECT 26.480 224.250 30.330 224.400 ;
        RECT 19.130 223.800 19.430 224.250 ;
        RECT 30.030 223.800 30.330 224.250 ;
        RECT 19.130 223.650 22.980 223.800 ;
        RECT 26.480 223.650 30.330 223.800 ;
        RECT 19.130 223.200 19.430 223.650 ;
        RECT 30.030 223.200 30.330 223.650 ;
        RECT 19.130 223.050 22.980 223.200 ;
        RECT 26.480 223.050 30.330 223.200 ;
        RECT 19.130 222.600 19.430 223.050 ;
        RECT 30.030 222.600 30.330 223.050 ;
        RECT 19.130 222.450 22.980 222.600 ;
        RECT 26.480 222.450 30.330 222.600 ;
        RECT 19.130 222.000 19.430 222.450 ;
        RECT 30.030 222.000 30.330 222.450 ;
        RECT 19.130 221.450 22.930 222.000 ;
        RECT 6.530 221.400 22.930 221.450 ;
        RECT 26.530 221.450 30.330 222.000 ;
        RECT 30.780 221.450 30.930 229.650 ;
        RECT 31.380 221.450 31.530 229.650 ;
        RECT 31.980 221.450 32.130 229.650 ;
        RECT 32.580 221.450 32.730 229.650 ;
        RECT 33.180 221.450 33.330 229.650 ;
        RECT 33.780 221.450 33.930 229.650 ;
        RECT 34.380 221.450 35.080 238.550 ;
        RECT 35.530 230.350 35.680 238.550 ;
        RECT 36.130 230.350 36.280 238.550 ;
        RECT 36.730 230.350 36.880 238.550 ;
        RECT 37.330 230.350 37.480 238.550 ;
        RECT 37.930 230.350 38.080 238.550 ;
        RECT 38.530 230.350 38.680 238.550 ;
        RECT 39.130 238.000 42.930 238.550 ;
        RECT 46.530 238.550 62.930 238.600 ;
        RECT 46.530 238.000 50.330 238.550 ;
        RECT 39.130 237.550 39.430 238.000 ;
        RECT 50.030 237.550 50.330 238.000 ;
        RECT 39.130 237.400 42.980 237.550 ;
        RECT 46.480 237.400 50.330 237.550 ;
        RECT 39.130 236.950 39.430 237.400 ;
        RECT 50.030 236.950 50.330 237.400 ;
        RECT 39.130 236.800 42.980 236.950 ;
        RECT 46.480 236.800 50.330 236.950 ;
        RECT 39.130 236.350 39.430 236.800 ;
        RECT 50.030 236.350 50.330 236.800 ;
        RECT 39.130 236.200 42.980 236.350 ;
        RECT 46.480 236.200 50.330 236.350 ;
        RECT 39.130 235.750 39.430 236.200 ;
        RECT 50.030 235.750 50.330 236.200 ;
        RECT 39.130 235.600 42.980 235.750 ;
        RECT 46.480 235.600 50.330 235.750 ;
        RECT 39.130 235.150 39.430 235.600 ;
        RECT 50.030 235.150 50.330 235.600 ;
        RECT 39.130 235.000 42.980 235.150 ;
        RECT 46.480 235.000 50.330 235.150 ;
        RECT 39.130 234.550 39.430 235.000 ;
        RECT 50.030 234.550 50.330 235.000 ;
        RECT 39.130 234.400 42.980 234.550 ;
        RECT 46.480 234.400 50.330 234.550 ;
        RECT 39.130 233.950 39.430 234.400 ;
        RECT 50.030 233.950 50.330 234.400 ;
        RECT 39.130 233.800 42.980 233.950 ;
        RECT 46.480 233.800 50.330 233.950 ;
        RECT 39.130 233.350 39.430 233.800 ;
        RECT 50.030 233.350 50.330 233.800 ;
        RECT 39.130 233.200 42.980 233.350 ;
        RECT 46.480 233.200 50.330 233.350 ;
        RECT 39.130 232.750 39.430 233.200 ;
        RECT 39.130 232.600 42.980 232.750 ;
        RECT 39.130 232.150 39.430 232.600 ;
        RECT 39.130 232.000 42.980 232.150 ;
        RECT 39.130 231.550 39.430 232.000 ;
        RECT 39.130 231.400 42.980 231.550 ;
        RECT 39.130 230.950 39.430 231.400 ;
        RECT 39.130 230.800 42.980 230.950 ;
        RECT 39.130 230.350 39.430 230.800 ;
        RECT 35.530 221.450 35.680 229.650 ;
        RECT 36.130 221.450 36.280 229.650 ;
        RECT 36.730 221.450 36.880 229.650 ;
        RECT 37.330 221.450 37.480 229.650 ;
        RECT 37.930 221.450 38.080 229.650 ;
        RECT 38.530 221.450 38.680 229.650 ;
        RECT 39.130 229.200 39.430 229.650 ;
        RECT 39.130 229.050 42.980 229.200 ;
        RECT 39.130 228.600 39.430 229.050 ;
        RECT 39.130 228.450 42.980 228.600 ;
        RECT 39.130 228.000 39.430 228.450 ;
        RECT 39.130 227.850 42.980 228.000 ;
        RECT 39.130 227.400 39.430 227.850 ;
        RECT 39.130 227.250 42.980 227.400 ;
        RECT 39.130 226.800 39.430 227.250 ;
        RECT 43.830 226.800 45.630 233.200 ;
        RECT 50.030 232.750 50.330 233.200 ;
        RECT 46.480 232.600 50.330 232.750 ;
        RECT 50.030 232.150 50.330 232.600 ;
        RECT 46.480 232.000 50.330 232.150 ;
        RECT 50.030 231.550 50.330 232.000 ;
        RECT 46.480 231.400 50.330 231.550 ;
        RECT 50.030 230.950 50.330 231.400 ;
        RECT 46.480 230.800 50.330 230.950 ;
        RECT 50.030 230.350 50.330 230.800 ;
        RECT 50.780 230.350 50.930 238.550 ;
        RECT 51.380 230.350 51.530 238.550 ;
        RECT 51.980 230.350 52.130 238.550 ;
        RECT 52.580 230.350 52.730 238.550 ;
        RECT 53.180 230.350 53.330 238.550 ;
        RECT 53.780 230.350 53.930 238.550 ;
        RECT 50.030 229.200 50.330 229.650 ;
        RECT 46.480 229.050 50.330 229.200 ;
        RECT 50.030 228.600 50.330 229.050 ;
        RECT 46.480 228.450 50.330 228.600 ;
        RECT 50.030 228.000 50.330 228.450 ;
        RECT 46.480 227.850 50.330 228.000 ;
        RECT 50.030 227.400 50.330 227.850 ;
        RECT 46.480 227.250 50.330 227.400 ;
        RECT 50.030 226.800 50.330 227.250 ;
        RECT 39.130 226.650 42.980 226.800 ;
        RECT 46.480 226.650 50.330 226.800 ;
        RECT 39.130 226.200 39.430 226.650 ;
        RECT 50.030 226.200 50.330 226.650 ;
        RECT 39.130 226.050 42.980 226.200 ;
        RECT 46.480 226.050 50.330 226.200 ;
        RECT 39.130 225.600 39.430 226.050 ;
        RECT 50.030 225.600 50.330 226.050 ;
        RECT 39.130 225.450 42.980 225.600 ;
        RECT 46.480 225.450 50.330 225.600 ;
        RECT 39.130 225.000 39.430 225.450 ;
        RECT 50.030 225.000 50.330 225.450 ;
        RECT 39.130 224.850 42.980 225.000 ;
        RECT 46.480 224.850 50.330 225.000 ;
        RECT 39.130 224.400 39.430 224.850 ;
        RECT 50.030 224.400 50.330 224.850 ;
        RECT 39.130 224.250 42.980 224.400 ;
        RECT 46.480 224.250 50.330 224.400 ;
        RECT 39.130 223.800 39.430 224.250 ;
        RECT 50.030 223.800 50.330 224.250 ;
        RECT 39.130 223.650 42.980 223.800 ;
        RECT 46.480 223.650 50.330 223.800 ;
        RECT 39.130 223.200 39.430 223.650 ;
        RECT 50.030 223.200 50.330 223.650 ;
        RECT 39.130 223.050 42.980 223.200 ;
        RECT 46.480 223.050 50.330 223.200 ;
        RECT 39.130 222.600 39.430 223.050 ;
        RECT 50.030 222.600 50.330 223.050 ;
        RECT 39.130 222.450 42.980 222.600 ;
        RECT 46.480 222.450 50.330 222.600 ;
        RECT 39.130 222.000 39.430 222.450 ;
        RECT 50.030 222.000 50.330 222.450 ;
        RECT 39.130 221.450 42.930 222.000 ;
        RECT 26.530 221.400 42.930 221.450 ;
        RECT 46.530 221.450 50.330 222.000 ;
        RECT 50.780 221.450 50.930 229.650 ;
        RECT 51.380 221.450 51.530 229.650 ;
        RECT 51.980 221.450 52.130 229.650 ;
        RECT 52.580 221.450 52.730 229.650 ;
        RECT 53.180 221.450 53.330 229.650 ;
        RECT 53.780 221.450 53.930 229.650 ;
        RECT 54.380 221.450 55.080 238.550 ;
        RECT 55.530 230.350 55.680 238.550 ;
        RECT 56.130 230.350 56.280 238.550 ;
        RECT 56.730 230.350 56.880 238.550 ;
        RECT 57.330 230.350 57.480 238.550 ;
        RECT 57.930 230.350 58.080 238.550 ;
        RECT 58.530 230.350 58.680 238.550 ;
        RECT 59.130 238.000 62.930 238.550 ;
        RECT 66.530 238.550 82.930 238.600 ;
        RECT 66.530 238.000 70.330 238.550 ;
        RECT 59.130 237.550 59.430 238.000 ;
        RECT 70.030 237.550 70.330 238.000 ;
        RECT 59.130 237.400 62.980 237.550 ;
        RECT 66.480 237.400 70.330 237.550 ;
        RECT 59.130 236.950 59.430 237.400 ;
        RECT 70.030 236.950 70.330 237.400 ;
        RECT 59.130 236.800 62.980 236.950 ;
        RECT 66.480 236.800 70.330 236.950 ;
        RECT 59.130 236.350 59.430 236.800 ;
        RECT 70.030 236.350 70.330 236.800 ;
        RECT 59.130 236.200 62.980 236.350 ;
        RECT 66.480 236.200 70.330 236.350 ;
        RECT 59.130 235.750 59.430 236.200 ;
        RECT 70.030 235.750 70.330 236.200 ;
        RECT 59.130 235.600 62.980 235.750 ;
        RECT 66.480 235.600 70.330 235.750 ;
        RECT 59.130 235.150 59.430 235.600 ;
        RECT 70.030 235.150 70.330 235.600 ;
        RECT 59.130 235.000 62.980 235.150 ;
        RECT 66.480 235.000 70.330 235.150 ;
        RECT 59.130 234.550 59.430 235.000 ;
        RECT 70.030 234.550 70.330 235.000 ;
        RECT 59.130 234.400 62.980 234.550 ;
        RECT 66.480 234.400 70.330 234.550 ;
        RECT 59.130 233.950 59.430 234.400 ;
        RECT 70.030 233.950 70.330 234.400 ;
        RECT 59.130 233.800 62.980 233.950 ;
        RECT 66.480 233.800 70.330 233.950 ;
        RECT 59.130 233.350 59.430 233.800 ;
        RECT 70.030 233.350 70.330 233.800 ;
        RECT 59.130 233.200 62.980 233.350 ;
        RECT 66.480 233.200 70.330 233.350 ;
        RECT 59.130 232.750 59.430 233.200 ;
        RECT 59.130 232.600 62.980 232.750 ;
        RECT 59.130 232.150 59.430 232.600 ;
        RECT 59.130 232.000 62.980 232.150 ;
        RECT 59.130 231.550 59.430 232.000 ;
        RECT 59.130 231.400 62.980 231.550 ;
        RECT 59.130 230.950 59.430 231.400 ;
        RECT 59.130 230.800 62.980 230.950 ;
        RECT 59.130 230.350 59.430 230.800 ;
        RECT 55.530 221.450 55.680 229.650 ;
        RECT 56.130 221.450 56.280 229.650 ;
        RECT 56.730 221.450 56.880 229.650 ;
        RECT 57.330 221.450 57.480 229.650 ;
        RECT 57.930 221.450 58.080 229.650 ;
        RECT 58.530 221.450 58.680 229.650 ;
        RECT 59.130 229.200 59.430 229.650 ;
        RECT 59.130 229.050 62.980 229.200 ;
        RECT 59.130 228.600 59.430 229.050 ;
        RECT 59.130 228.450 62.980 228.600 ;
        RECT 59.130 228.000 59.430 228.450 ;
        RECT 59.130 227.850 62.980 228.000 ;
        RECT 59.130 227.400 59.430 227.850 ;
        RECT 59.130 227.250 62.980 227.400 ;
        RECT 59.130 226.800 59.430 227.250 ;
        RECT 63.830 226.800 65.630 233.200 ;
        RECT 70.030 232.750 70.330 233.200 ;
        RECT 66.480 232.600 70.330 232.750 ;
        RECT 70.030 232.150 70.330 232.600 ;
        RECT 66.480 232.000 70.330 232.150 ;
        RECT 70.030 231.550 70.330 232.000 ;
        RECT 66.480 231.400 70.330 231.550 ;
        RECT 70.030 230.950 70.330 231.400 ;
        RECT 66.480 230.800 70.330 230.950 ;
        RECT 70.030 230.350 70.330 230.800 ;
        RECT 70.780 230.350 70.930 238.550 ;
        RECT 71.380 230.350 71.530 238.550 ;
        RECT 71.980 230.350 72.130 238.550 ;
        RECT 72.580 230.350 72.730 238.550 ;
        RECT 73.180 230.350 73.330 238.550 ;
        RECT 73.780 230.350 73.930 238.550 ;
        RECT 70.030 229.200 70.330 229.650 ;
        RECT 66.480 229.050 70.330 229.200 ;
        RECT 70.030 228.600 70.330 229.050 ;
        RECT 66.480 228.450 70.330 228.600 ;
        RECT 70.030 228.000 70.330 228.450 ;
        RECT 66.480 227.850 70.330 228.000 ;
        RECT 70.030 227.400 70.330 227.850 ;
        RECT 66.480 227.250 70.330 227.400 ;
        RECT 70.030 226.800 70.330 227.250 ;
        RECT 59.130 226.650 62.980 226.800 ;
        RECT 66.480 226.650 70.330 226.800 ;
        RECT 59.130 226.200 59.430 226.650 ;
        RECT 70.030 226.200 70.330 226.650 ;
        RECT 59.130 226.050 62.980 226.200 ;
        RECT 66.480 226.050 70.330 226.200 ;
        RECT 59.130 225.600 59.430 226.050 ;
        RECT 70.030 225.600 70.330 226.050 ;
        RECT 59.130 225.450 62.980 225.600 ;
        RECT 66.480 225.450 70.330 225.600 ;
        RECT 59.130 225.000 59.430 225.450 ;
        RECT 70.030 225.000 70.330 225.450 ;
        RECT 59.130 224.850 62.980 225.000 ;
        RECT 66.480 224.850 70.330 225.000 ;
        RECT 59.130 224.400 59.430 224.850 ;
        RECT 70.030 224.400 70.330 224.850 ;
        RECT 59.130 224.250 62.980 224.400 ;
        RECT 66.480 224.250 70.330 224.400 ;
        RECT 59.130 223.800 59.430 224.250 ;
        RECT 70.030 223.800 70.330 224.250 ;
        RECT 59.130 223.650 62.980 223.800 ;
        RECT 66.480 223.650 70.330 223.800 ;
        RECT 59.130 223.200 59.430 223.650 ;
        RECT 70.030 223.200 70.330 223.650 ;
        RECT 59.130 223.050 62.980 223.200 ;
        RECT 66.480 223.050 70.330 223.200 ;
        RECT 59.130 222.600 59.430 223.050 ;
        RECT 70.030 222.600 70.330 223.050 ;
        RECT 59.130 222.450 62.980 222.600 ;
        RECT 66.480 222.450 70.330 222.600 ;
        RECT 59.130 222.000 59.430 222.450 ;
        RECT 70.030 222.000 70.330 222.450 ;
        RECT 59.130 221.450 62.930 222.000 ;
        RECT 46.530 221.400 62.930 221.450 ;
        RECT 66.530 221.450 70.330 222.000 ;
        RECT 70.780 221.450 70.930 229.650 ;
        RECT 71.380 221.450 71.530 229.650 ;
        RECT 71.980 221.450 72.130 229.650 ;
        RECT 72.580 221.450 72.730 229.650 ;
        RECT 73.180 221.450 73.330 229.650 ;
        RECT 73.780 221.450 73.930 229.650 ;
        RECT 74.380 221.450 75.080 238.550 ;
        RECT 75.530 230.350 75.680 238.550 ;
        RECT 76.130 230.350 76.280 238.550 ;
        RECT 76.730 230.350 76.880 238.550 ;
        RECT 77.330 230.350 77.480 238.550 ;
        RECT 77.930 230.350 78.080 238.550 ;
        RECT 78.530 230.350 78.680 238.550 ;
        RECT 79.130 238.000 82.930 238.550 ;
        RECT 86.530 238.550 102.930 238.600 ;
        RECT 86.530 238.000 90.330 238.550 ;
        RECT 79.130 237.550 79.430 238.000 ;
        RECT 90.030 237.550 90.330 238.000 ;
        RECT 79.130 237.400 82.980 237.550 ;
        RECT 86.480 237.400 90.330 237.550 ;
        RECT 79.130 236.950 79.430 237.400 ;
        RECT 90.030 236.950 90.330 237.400 ;
        RECT 79.130 236.800 82.980 236.950 ;
        RECT 86.480 236.800 90.330 236.950 ;
        RECT 79.130 236.350 79.430 236.800 ;
        RECT 90.030 236.350 90.330 236.800 ;
        RECT 79.130 236.200 82.980 236.350 ;
        RECT 86.480 236.200 90.330 236.350 ;
        RECT 79.130 235.750 79.430 236.200 ;
        RECT 90.030 235.750 90.330 236.200 ;
        RECT 79.130 235.600 82.980 235.750 ;
        RECT 86.480 235.600 90.330 235.750 ;
        RECT 79.130 235.150 79.430 235.600 ;
        RECT 90.030 235.150 90.330 235.600 ;
        RECT 79.130 235.000 82.980 235.150 ;
        RECT 86.480 235.000 90.330 235.150 ;
        RECT 79.130 234.550 79.430 235.000 ;
        RECT 90.030 234.550 90.330 235.000 ;
        RECT 79.130 234.400 82.980 234.550 ;
        RECT 86.480 234.400 90.330 234.550 ;
        RECT 79.130 233.950 79.430 234.400 ;
        RECT 90.030 233.950 90.330 234.400 ;
        RECT 79.130 233.800 82.980 233.950 ;
        RECT 86.480 233.800 90.330 233.950 ;
        RECT 79.130 233.350 79.430 233.800 ;
        RECT 90.030 233.350 90.330 233.800 ;
        RECT 79.130 233.200 82.980 233.350 ;
        RECT 86.480 233.200 90.330 233.350 ;
        RECT 79.130 232.750 79.430 233.200 ;
        RECT 79.130 232.600 82.980 232.750 ;
        RECT 79.130 232.150 79.430 232.600 ;
        RECT 79.130 232.000 82.980 232.150 ;
        RECT 79.130 231.550 79.430 232.000 ;
        RECT 79.130 231.400 82.980 231.550 ;
        RECT 79.130 230.950 79.430 231.400 ;
        RECT 79.130 230.800 82.980 230.950 ;
        RECT 79.130 230.350 79.430 230.800 ;
        RECT 75.530 221.450 75.680 229.650 ;
        RECT 76.130 221.450 76.280 229.650 ;
        RECT 76.730 221.450 76.880 229.650 ;
        RECT 77.330 221.450 77.480 229.650 ;
        RECT 77.930 221.450 78.080 229.650 ;
        RECT 78.530 221.450 78.680 229.650 ;
        RECT 79.130 229.200 79.430 229.650 ;
        RECT 79.130 229.050 82.980 229.200 ;
        RECT 79.130 228.600 79.430 229.050 ;
        RECT 79.130 228.450 82.980 228.600 ;
        RECT 79.130 228.000 79.430 228.450 ;
        RECT 79.130 227.850 82.980 228.000 ;
        RECT 79.130 227.400 79.430 227.850 ;
        RECT 79.130 227.250 82.980 227.400 ;
        RECT 79.130 226.800 79.430 227.250 ;
        RECT 83.830 226.800 85.630 233.200 ;
        RECT 90.030 232.750 90.330 233.200 ;
        RECT 86.480 232.600 90.330 232.750 ;
        RECT 90.030 232.150 90.330 232.600 ;
        RECT 86.480 232.000 90.330 232.150 ;
        RECT 90.030 231.550 90.330 232.000 ;
        RECT 86.480 231.400 90.330 231.550 ;
        RECT 90.030 230.950 90.330 231.400 ;
        RECT 86.480 230.800 90.330 230.950 ;
        RECT 90.030 230.350 90.330 230.800 ;
        RECT 90.780 230.350 90.930 238.550 ;
        RECT 91.380 230.350 91.530 238.550 ;
        RECT 91.980 230.350 92.130 238.550 ;
        RECT 92.580 230.350 92.730 238.550 ;
        RECT 93.180 230.350 93.330 238.550 ;
        RECT 93.780 230.350 93.930 238.550 ;
        RECT 90.030 229.200 90.330 229.650 ;
        RECT 86.480 229.050 90.330 229.200 ;
        RECT 90.030 228.600 90.330 229.050 ;
        RECT 86.480 228.450 90.330 228.600 ;
        RECT 90.030 228.000 90.330 228.450 ;
        RECT 86.480 227.850 90.330 228.000 ;
        RECT 90.030 227.400 90.330 227.850 ;
        RECT 86.480 227.250 90.330 227.400 ;
        RECT 90.030 226.800 90.330 227.250 ;
        RECT 79.130 226.650 82.980 226.800 ;
        RECT 86.480 226.650 90.330 226.800 ;
        RECT 79.130 226.200 79.430 226.650 ;
        RECT 90.030 226.200 90.330 226.650 ;
        RECT 79.130 226.050 82.980 226.200 ;
        RECT 86.480 226.050 90.330 226.200 ;
        RECT 79.130 225.600 79.430 226.050 ;
        RECT 90.030 225.600 90.330 226.050 ;
        RECT 79.130 225.450 82.980 225.600 ;
        RECT 86.480 225.450 90.330 225.600 ;
        RECT 79.130 225.000 79.430 225.450 ;
        RECT 90.030 225.000 90.330 225.450 ;
        RECT 79.130 224.850 82.980 225.000 ;
        RECT 86.480 224.850 90.330 225.000 ;
        RECT 79.130 224.400 79.430 224.850 ;
        RECT 90.030 224.400 90.330 224.850 ;
        RECT 79.130 224.250 82.980 224.400 ;
        RECT 86.480 224.250 90.330 224.400 ;
        RECT 79.130 223.800 79.430 224.250 ;
        RECT 90.030 223.800 90.330 224.250 ;
        RECT 79.130 223.650 82.980 223.800 ;
        RECT 86.480 223.650 90.330 223.800 ;
        RECT 79.130 223.200 79.430 223.650 ;
        RECT 90.030 223.200 90.330 223.650 ;
        RECT 79.130 223.050 82.980 223.200 ;
        RECT 86.480 223.050 90.330 223.200 ;
        RECT 79.130 222.600 79.430 223.050 ;
        RECT 90.030 222.600 90.330 223.050 ;
        RECT 79.130 222.450 82.980 222.600 ;
        RECT 86.480 222.450 90.330 222.600 ;
        RECT 79.130 222.000 79.430 222.450 ;
        RECT 90.030 222.000 90.330 222.450 ;
        RECT 79.130 221.450 82.930 222.000 ;
        RECT 66.530 221.400 82.930 221.450 ;
        RECT 86.530 221.450 90.330 222.000 ;
        RECT 90.780 221.450 90.930 229.650 ;
        RECT 91.380 221.450 91.530 229.650 ;
        RECT 91.980 221.450 92.130 229.650 ;
        RECT 92.580 221.450 92.730 229.650 ;
        RECT 93.180 221.450 93.330 229.650 ;
        RECT 93.780 221.450 93.930 229.650 ;
        RECT 94.380 221.450 95.080 238.550 ;
        RECT 95.530 230.350 95.680 238.550 ;
        RECT 96.130 230.350 96.280 238.550 ;
        RECT 96.730 230.350 96.880 238.550 ;
        RECT 97.330 230.350 97.480 238.550 ;
        RECT 97.930 230.350 98.080 238.550 ;
        RECT 98.530 230.350 98.680 238.550 ;
        RECT 99.130 238.000 102.930 238.550 ;
        RECT 99.130 237.550 99.430 238.000 ;
        RECT 99.130 237.400 102.980 237.550 ;
        RECT 99.130 236.950 99.430 237.400 ;
        RECT 99.130 236.800 102.980 236.950 ;
        RECT 99.130 236.350 99.430 236.800 ;
        RECT 99.130 236.200 102.980 236.350 ;
        RECT 99.130 235.750 99.430 236.200 ;
        RECT 99.130 235.600 102.980 235.750 ;
        RECT 99.130 235.150 99.430 235.600 ;
        RECT 99.130 235.000 102.980 235.150 ;
        RECT 99.130 234.550 99.430 235.000 ;
        RECT 99.130 234.400 102.980 234.550 ;
        RECT 99.130 233.950 99.430 234.400 ;
        RECT 99.130 233.800 102.980 233.950 ;
        RECT 99.130 233.350 99.430 233.800 ;
        RECT 99.130 233.200 102.980 233.350 ;
        RECT 99.130 232.750 99.430 233.200 ;
        RECT 99.130 232.600 102.980 232.750 ;
        RECT 99.130 232.150 99.430 232.600 ;
        RECT 99.130 232.000 102.980 232.150 ;
        RECT 99.130 231.550 99.430 232.000 ;
        RECT 99.130 231.400 102.980 231.550 ;
        RECT 99.130 230.950 99.430 231.400 ;
        RECT 99.130 230.800 102.980 230.950 ;
        RECT 99.130 230.350 99.430 230.800 ;
        RECT 95.530 221.450 95.680 229.650 ;
        RECT 96.130 221.450 96.280 229.650 ;
        RECT 96.730 221.450 96.880 229.650 ;
        RECT 97.330 221.450 97.480 229.650 ;
        RECT 97.930 221.450 98.080 229.650 ;
        RECT 98.530 221.450 98.680 229.650 ;
        RECT 99.130 229.200 99.430 229.650 ;
        RECT 99.130 229.050 102.980 229.200 ;
        RECT 99.130 228.600 99.430 229.050 ;
        RECT 99.130 228.450 102.980 228.600 ;
        RECT 99.130 228.000 99.430 228.450 ;
        RECT 99.130 227.850 102.980 228.000 ;
        RECT 99.130 227.400 99.430 227.850 ;
        RECT 99.130 227.250 102.980 227.400 ;
        RECT 99.130 226.800 99.430 227.250 ;
        RECT 103.830 226.800 104.730 233.200 ;
        RECT 109.850 228.350 111.850 229.625 ;
        RECT 99.130 226.650 102.980 226.800 ;
        RECT 99.130 226.200 99.430 226.650 ;
        RECT 99.130 226.050 102.980 226.200 ;
        RECT 99.130 225.600 99.430 226.050 ;
        RECT 99.130 225.450 102.980 225.600 ;
        RECT 99.130 225.000 99.430 225.450 ;
        RECT 99.130 224.850 102.980 225.000 ;
        RECT 99.130 224.400 99.430 224.850 ;
        RECT 99.130 224.250 102.980 224.400 ;
        RECT 99.130 223.800 99.430 224.250 ;
        RECT 99.130 223.650 102.980 223.800 ;
        RECT 99.130 223.200 99.430 223.650 ;
        RECT 99.130 223.050 102.980 223.200 ;
        RECT 99.130 222.600 99.430 223.050 ;
        RECT 99.130 222.450 102.980 222.600 ;
        RECT 99.130 222.000 99.430 222.450 ;
        RECT 99.130 221.450 102.930 222.000 ;
        RECT 86.530 221.400 102.930 221.450 ;
        RECT 9.630 220.900 19.830 221.400 ;
        RECT 29.630 220.900 39.830 221.400 ;
        RECT 49.630 220.900 59.830 221.400 ;
        RECT 69.630 220.900 79.830 221.400 ;
        RECT 89.630 220.900 99.830 221.400 ;
        RECT 11.530 220.000 17.930 220.900 ;
        RECT 31.530 220.000 37.930 220.900 ;
        RECT 51.530 220.000 57.930 220.900 ;
        RECT 71.530 220.000 77.930 220.900 ;
        RECT 91.530 220.000 97.930 220.900 ;
        RECT 12.340 198.555 14.335 220.000 ;
        RECT 109.850 217.400 111.850 219.350 ;
        RECT 9.335 197.190 14.340 198.555 ;
        RECT 9.340 197.050 11.335 197.190 ;
        RECT 9.340 196.350 11.675 197.050 ;
        RECT 9.340 164.680 11.335 196.350 ;
        RECT 109.850 182.980 111.850 184.930 ;
        RECT 9.340 163.550 13.710 164.680 ;
        RECT 9.330 162.425 13.710 163.550 ;
        RECT 11.530 160.000 13.710 162.425 ;
        RECT 11.530 159.100 17.930 160.000 ;
        RECT 31.530 159.100 37.930 160.000 ;
        RECT 51.530 159.100 57.930 160.000 ;
        RECT 71.530 159.100 77.930 160.000 ;
        RECT 91.530 159.100 97.930 160.000 ;
        RECT 9.630 158.600 19.830 159.100 ;
        RECT 29.630 158.600 39.830 159.100 ;
        RECT 49.630 158.600 59.830 159.100 ;
        RECT 69.630 158.600 79.830 159.100 ;
        RECT 89.630 158.600 99.830 159.100 ;
        RECT 6.530 158.550 22.930 158.600 ;
        RECT 6.530 158.000 10.330 158.550 ;
        RECT 10.030 157.550 10.330 158.000 ;
        RECT 6.480 157.400 10.330 157.550 ;
        RECT 10.030 156.950 10.330 157.400 ;
        RECT 6.480 156.800 10.330 156.950 ;
        RECT 10.030 156.350 10.330 156.800 ;
        RECT 6.480 156.200 10.330 156.350 ;
        RECT 10.030 155.750 10.330 156.200 ;
        RECT 6.480 155.600 10.330 155.750 ;
        RECT 10.030 155.150 10.330 155.600 ;
        RECT 6.480 155.000 10.330 155.150 ;
        RECT 10.030 154.550 10.330 155.000 ;
        RECT 6.480 154.400 10.330 154.550 ;
        RECT 10.030 153.950 10.330 154.400 ;
        RECT 6.480 153.800 10.330 153.950 ;
        RECT 10.030 153.350 10.330 153.800 ;
        RECT 6.480 153.200 10.330 153.350 ;
        RECT 4.730 146.800 5.630 153.200 ;
        RECT 10.030 152.750 10.330 153.200 ;
        RECT 6.480 152.600 10.330 152.750 ;
        RECT 10.030 152.150 10.330 152.600 ;
        RECT 6.480 152.000 10.330 152.150 ;
        RECT 10.030 151.550 10.330 152.000 ;
        RECT 6.480 151.400 10.330 151.550 ;
        RECT 10.030 150.950 10.330 151.400 ;
        RECT 6.480 150.800 10.330 150.950 ;
        RECT 10.030 150.350 10.330 150.800 ;
        RECT 10.780 150.350 10.930 158.550 ;
        RECT 11.380 150.350 11.530 158.550 ;
        RECT 11.980 150.350 12.130 158.550 ;
        RECT 12.580 150.350 12.730 158.550 ;
        RECT 13.180 150.350 13.330 158.550 ;
        RECT 13.780 150.350 13.930 158.550 ;
        RECT 10.030 149.200 10.330 149.650 ;
        RECT 6.480 149.050 10.330 149.200 ;
        RECT 10.030 148.600 10.330 149.050 ;
        RECT 6.480 148.450 10.330 148.600 ;
        RECT 10.030 148.000 10.330 148.450 ;
        RECT 6.480 147.850 10.330 148.000 ;
        RECT 10.030 147.400 10.330 147.850 ;
        RECT 6.480 147.250 10.330 147.400 ;
        RECT 10.030 146.800 10.330 147.250 ;
        RECT 6.480 146.650 10.330 146.800 ;
        RECT 10.030 146.200 10.330 146.650 ;
        RECT 6.480 146.050 10.330 146.200 ;
        RECT 10.030 145.600 10.330 146.050 ;
        RECT 6.480 145.450 10.330 145.600 ;
        RECT 10.030 145.000 10.330 145.450 ;
        RECT 6.480 144.850 10.330 145.000 ;
        RECT 10.030 144.400 10.330 144.850 ;
        RECT 6.480 144.250 10.330 144.400 ;
        RECT 10.030 143.800 10.330 144.250 ;
        RECT 6.480 143.650 10.330 143.800 ;
        RECT 10.030 143.200 10.330 143.650 ;
        RECT 6.480 143.050 10.330 143.200 ;
        RECT 10.030 142.600 10.330 143.050 ;
        RECT 6.480 142.450 10.330 142.600 ;
        RECT 10.030 142.000 10.330 142.450 ;
        RECT 6.530 141.450 10.330 142.000 ;
        RECT 10.780 141.450 10.930 149.650 ;
        RECT 11.380 141.450 11.530 149.650 ;
        RECT 11.980 141.450 12.130 149.650 ;
        RECT 12.580 141.450 12.730 149.650 ;
        RECT 13.180 141.450 13.330 149.650 ;
        RECT 13.780 141.450 13.930 149.650 ;
        RECT 14.380 141.450 15.080 158.550 ;
        RECT 15.530 150.350 15.680 158.550 ;
        RECT 16.130 150.350 16.280 158.550 ;
        RECT 16.730 150.350 16.880 158.550 ;
        RECT 17.330 150.350 17.480 158.550 ;
        RECT 17.930 150.350 18.080 158.550 ;
        RECT 18.530 150.350 18.680 158.550 ;
        RECT 19.130 158.000 22.930 158.550 ;
        RECT 26.530 158.550 42.930 158.600 ;
        RECT 26.530 158.000 30.330 158.550 ;
        RECT 19.130 157.550 19.430 158.000 ;
        RECT 30.030 157.550 30.330 158.000 ;
        RECT 19.130 157.400 22.980 157.550 ;
        RECT 26.480 157.400 30.330 157.550 ;
        RECT 19.130 156.950 19.430 157.400 ;
        RECT 30.030 156.950 30.330 157.400 ;
        RECT 19.130 156.800 22.980 156.950 ;
        RECT 26.480 156.800 30.330 156.950 ;
        RECT 19.130 156.350 19.430 156.800 ;
        RECT 30.030 156.350 30.330 156.800 ;
        RECT 19.130 156.200 22.980 156.350 ;
        RECT 26.480 156.200 30.330 156.350 ;
        RECT 19.130 155.750 19.430 156.200 ;
        RECT 30.030 155.750 30.330 156.200 ;
        RECT 19.130 155.600 22.980 155.750 ;
        RECT 26.480 155.600 30.330 155.750 ;
        RECT 19.130 155.150 19.430 155.600 ;
        RECT 30.030 155.150 30.330 155.600 ;
        RECT 19.130 155.000 22.980 155.150 ;
        RECT 26.480 155.000 30.330 155.150 ;
        RECT 19.130 154.550 19.430 155.000 ;
        RECT 30.030 154.550 30.330 155.000 ;
        RECT 19.130 154.400 22.980 154.550 ;
        RECT 26.480 154.400 30.330 154.550 ;
        RECT 19.130 153.950 19.430 154.400 ;
        RECT 30.030 153.950 30.330 154.400 ;
        RECT 19.130 153.800 22.980 153.950 ;
        RECT 26.480 153.800 30.330 153.950 ;
        RECT 19.130 153.350 19.430 153.800 ;
        RECT 30.030 153.350 30.330 153.800 ;
        RECT 19.130 153.200 22.980 153.350 ;
        RECT 26.480 153.200 30.330 153.350 ;
        RECT 19.130 152.750 19.430 153.200 ;
        RECT 19.130 152.600 22.980 152.750 ;
        RECT 19.130 152.150 19.430 152.600 ;
        RECT 19.130 152.000 22.980 152.150 ;
        RECT 19.130 151.550 19.430 152.000 ;
        RECT 19.130 151.400 22.980 151.550 ;
        RECT 19.130 150.950 19.430 151.400 ;
        RECT 19.130 150.800 22.980 150.950 ;
        RECT 19.130 150.350 19.430 150.800 ;
        RECT 15.530 141.450 15.680 149.650 ;
        RECT 16.130 141.450 16.280 149.650 ;
        RECT 16.730 141.450 16.880 149.650 ;
        RECT 17.330 141.450 17.480 149.650 ;
        RECT 17.930 141.450 18.080 149.650 ;
        RECT 18.530 141.450 18.680 149.650 ;
        RECT 19.130 149.200 19.430 149.650 ;
        RECT 19.130 149.050 22.980 149.200 ;
        RECT 19.130 148.600 19.430 149.050 ;
        RECT 19.130 148.450 22.980 148.600 ;
        RECT 19.130 148.000 19.430 148.450 ;
        RECT 19.130 147.850 22.980 148.000 ;
        RECT 19.130 147.400 19.430 147.850 ;
        RECT 19.130 147.250 22.980 147.400 ;
        RECT 19.130 146.800 19.430 147.250 ;
        RECT 23.830 146.800 25.630 153.200 ;
        RECT 30.030 152.750 30.330 153.200 ;
        RECT 26.480 152.600 30.330 152.750 ;
        RECT 30.030 152.150 30.330 152.600 ;
        RECT 26.480 152.000 30.330 152.150 ;
        RECT 30.030 151.550 30.330 152.000 ;
        RECT 26.480 151.400 30.330 151.550 ;
        RECT 30.030 150.950 30.330 151.400 ;
        RECT 26.480 150.800 30.330 150.950 ;
        RECT 30.030 150.350 30.330 150.800 ;
        RECT 30.780 150.350 30.930 158.550 ;
        RECT 31.380 150.350 31.530 158.550 ;
        RECT 31.980 150.350 32.130 158.550 ;
        RECT 32.580 150.350 32.730 158.550 ;
        RECT 33.180 150.350 33.330 158.550 ;
        RECT 33.780 150.350 33.930 158.550 ;
        RECT 30.030 149.200 30.330 149.650 ;
        RECT 26.480 149.050 30.330 149.200 ;
        RECT 30.030 148.600 30.330 149.050 ;
        RECT 26.480 148.450 30.330 148.600 ;
        RECT 30.030 148.000 30.330 148.450 ;
        RECT 26.480 147.850 30.330 148.000 ;
        RECT 30.030 147.400 30.330 147.850 ;
        RECT 26.480 147.250 30.330 147.400 ;
        RECT 30.030 146.800 30.330 147.250 ;
        RECT 19.130 146.650 22.980 146.800 ;
        RECT 26.480 146.650 30.330 146.800 ;
        RECT 19.130 146.200 19.430 146.650 ;
        RECT 30.030 146.200 30.330 146.650 ;
        RECT 19.130 146.050 22.980 146.200 ;
        RECT 26.480 146.050 30.330 146.200 ;
        RECT 19.130 145.600 19.430 146.050 ;
        RECT 30.030 145.600 30.330 146.050 ;
        RECT 19.130 145.450 22.980 145.600 ;
        RECT 26.480 145.450 30.330 145.600 ;
        RECT 19.130 145.000 19.430 145.450 ;
        RECT 30.030 145.000 30.330 145.450 ;
        RECT 19.130 144.850 22.980 145.000 ;
        RECT 26.480 144.850 30.330 145.000 ;
        RECT 19.130 144.400 19.430 144.850 ;
        RECT 30.030 144.400 30.330 144.850 ;
        RECT 19.130 144.250 22.980 144.400 ;
        RECT 26.480 144.250 30.330 144.400 ;
        RECT 19.130 143.800 19.430 144.250 ;
        RECT 30.030 143.800 30.330 144.250 ;
        RECT 19.130 143.650 22.980 143.800 ;
        RECT 26.480 143.650 30.330 143.800 ;
        RECT 19.130 143.200 19.430 143.650 ;
        RECT 30.030 143.200 30.330 143.650 ;
        RECT 19.130 143.050 22.980 143.200 ;
        RECT 26.480 143.050 30.330 143.200 ;
        RECT 19.130 142.600 19.430 143.050 ;
        RECT 30.030 142.600 30.330 143.050 ;
        RECT 19.130 142.450 22.980 142.600 ;
        RECT 26.480 142.450 30.330 142.600 ;
        RECT 19.130 142.000 19.430 142.450 ;
        RECT 30.030 142.000 30.330 142.450 ;
        RECT 19.130 141.450 22.930 142.000 ;
        RECT 6.530 141.400 22.930 141.450 ;
        RECT 26.530 141.450 30.330 142.000 ;
        RECT 30.780 141.450 30.930 149.650 ;
        RECT 31.380 141.450 31.530 149.650 ;
        RECT 31.980 141.450 32.130 149.650 ;
        RECT 32.580 141.450 32.730 149.650 ;
        RECT 33.180 141.450 33.330 149.650 ;
        RECT 33.780 141.450 33.930 149.650 ;
        RECT 34.380 141.450 35.080 158.550 ;
        RECT 35.530 150.350 35.680 158.550 ;
        RECT 36.130 150.350 36.280 158.550 ;
        RECT 36.730 150.350 36.880 158.550 ;
        RECT 37.330 150.350 37.480 158.550 ;
        RECT 37.930 150.350 38.080 158.550 ;
        RECT 38.530 150.350 38.680 158.550 ;
        RECT 39.130 158.000 42.930 158.550 ;
        RECT 46.530 158.550 62.930 158.600 ;
        RECT 46.530 158.000 50.330 158.550 ;
        RECT 39.130 157.550 39.430 158.000 ;
        RECT 50.030 157.550 50.330 158.000 ;
        RECT 39.130 157.400 42.980 157.550 ;
        RECT 46.480 157.400 50.330 157.550 ;
        RECT 39.130 156.950 39.430 157.400 ;
        RECT 50.030 156.950 50.330 157.400 ;
        RECT 39.130 156.800 42.980 156.950 ;
        RECT 46.480 156.800 50.330 156.950 ;
        RECT 39.130 156.350 39.430 156.800 ;
        RECT 50.030 156.350 50.330 156.800 ;
        RECT 39.130 156.200 42.980 156.350 ;
        RECT 46.480 156.200 50.330 156.350 ;
        RECT 39.130 155.750 39.430 156.200 ;
        RECT 50.030 155.750 50.330 156.200 ;
        RECT 39.130 155.600 42.980 155.750 ;
        RECT 46.480 155.600 50.330 155.750 ;
        RECT 39.130 155.150 39.430 155.600 ;
        RECT 50.030 155.150 50.330 155.600 ;
        RECT 39.130 155.000 42.980 155.150 ;
        RECT 46.480 155.000 50.330 155.150 ;
        RECT 39.130 154.550 39.430 155.000 ;
        RECT 50.030 154.550 50.330 155.000 ;
        RECT 39.130 154.400 42.980 154.550 ;
        RECT 46.480 154.400 50.330 154.550 ;
        RECT 39.130 153.950 39.430 154.400 ;
        RECT 50.030 153.950 50.330 154.400 ;
        RECT 39.130 153.800 42.980 153.950 ;
        RECT 46.480 153.800 50.330 153.950 ;
        RECT 39.130 153.350 39.430 153.800 ;
        RECT 50.030 153.350 50.330 153.800 ;
        RECT 39.130 153.200 42.980 153.350 ;
        RECT 46.480 153.200 50.330 153.350 ;
        RECT 39.130 152.750 39.430 153.200 ;
        RECT 39.130 152.600 42.980 152.750 ;
        RECT 39.130 152.150 39.430 152.600 ;
        RECT 39.130 152.000 42.980 152.150 ;
        RECT 39.130 151.550 39.430 152.000 ;
        RECT 39.130 151.400 42.980 151.550 ;
        RECT 39.130 150.950 39.430 151.400 ;
        RECT 39.130 150.800 42.980 150.950 ;
        RECT 39.130 150.350 39.430 150.800 ;
        RECT 35.530 141.450 35.680 149.650 ;
        RECT 36.130 141.450 36.280 149.650 ;
        RECT 36.730 141.450 36.880 149.650 ;
        RECT 37.330 141.450 37.480 149.650 ;
        RECT 37.930 141.450 38.080 149.650 ;
        RECT 38.530 141.450 38.680 149.650 ;
        RECT 39.130 149.200 39.430 149.650 ;
        RECT 39.130 149.050 42.980 149.200 ;
        RECT 39.130 148.600 39.430 149.050 ;
        RECT 39.130 148.450 42.980 148.600 ;
        RECT 39.130 148.000 39.430 148.450 ;
        RECT 39.130 147.850 42.980 148.000 ;
        RECT 39.130 147.400 39.430 147.850 ;
        RECT 39.130 147.250 42.980 147.400 ;
        RECT 39.130 146.800 39.430 147.250 ;
        RECT 43.830 146.800 45.630 153.200 ;
        RECT 50.030 152.750 50.330 153.200 ;
        RECT 46.480 152.600 50.330 152.750 ;
        RECT 50.030 152.150 50.330 152.600 ;
        RECT 46.480 152.000 50.330 152.150 ;
        RECT 50.030 151.550 50.330 152.000 ;
        RECT 46.480 151.400 50.330 151.550 ;
        RECT 50.030 150.950 50.330 151.400 ;
        RECT 46.480 150.800 50.330 150.950 ;
        RECT 50.030 150.350 50.330 150.800 ;
        RECT 50.780 150.350 50.930 158.550 ;
        RECT 51.380 150.350 51.530 158.550 ;
        RECT 51.980 150.350 52.130 158.550 ;
        RECT 52.580 150.350 52.730 158.550 ;
        RECT 53.180 150.350 53.330 158.550 ;
        RECT 53.780 150.350 53.930 158.550 ;
        RECT 50.030 149.200 50.330 149.650 ;
        RECT 46.480 149.050 50.330 149.200 ;
        RECT 50.030 148.600 50.330 149.050 ;
        RECT 46.480 148.450 50.330 148.600 ;
        RECT 50.030 148.000 50.330 148.450 ;
        RECT 46.480 147.850 50.330 148.000 ;
        RECT 50.030 147.400 50.330 147.850 ;
        RECT 46.480 147.250 50.330 147.400 ;
        RECT 50.030 146.800 50.330 147.250 ;
        RECT 39.130 146.650 42.980 146.800 ;
        RECT 46.480 146.650 50.330 146.800 ;
        RECT 39.130 146.200 39.430 146.650 ;
        RECT 50.030 146.200 50.330 146.650 ;
        RECT 39.130 146.050 42.980 146.200 ;
        RECT 46.480 146.050 50.330 146.200 ;
        RECT 39.130 145.600 39.430 146.050 ;
        RECT 50.030 145.600 50.330 146.050 ;
        RECT 39.130 145.450 42.980 145.600 ;
        RECT 46.480 145.450 50.330 145.600 ;
        RECT 39.130 145.000 39.430 145.450 ;
        RECT 50.030 145.000 50.330 145.450 ;
        RECT 39.130 144.850 42.980 145.000 ;
        RECT 46.480 144.850 50.330 145.000 ;
        RECT 39.130 144.400 39.430 144.850 ;
        RECT 50.030 144.400 50.330 144.850 ;
        RECT 39.130 144.250 42.980 144.400 ;
        RECT 46.480 144.250 50.330 144.400 ;
        RECT 39.130 143.800 39.430 144.250 ;
        RECT 50.030 143.800 50.330 144.250 ;
        RECT 39.130 143.650 42.980 143.800 ;
        RECT 46.480 143.650 50.330 143.800 ;
        RECT 39.130 143.200 39.430 143.650 ;
        RECT 50.030 143.200 50.330 143.650 ;
        RECT 39.130 143.050 42.980 143.200 ;
        RECT 46.480 143.050 50.330 143.200 ;
        RECT 39.130 142.600 39.430 143.050 ;
        RECT 50.030 142.600 50.330 143.050 ;
        RECT 39.130 142.450 42.980 142.600 ;
        RECT 46.480 142.450 50.330 142.600 ;
        RECT 39.130 142.000 39.430 142.450 ;
        RECT 50.030 142.000 50.330 142.450 ;
        RECT 39.130 141.450 42.930 142.000 ;
        RECT 26.530 141.400 42.930 141.450 ;
        RECT 46.530 141.450 50.330 142.000 ;
        RECT 50.780 141.450 50.930 149.650 ;
        RECT 51.380 141.450 51.530 149.650 ;
        RECT 51.980 141.450 52.130 149.650 ;
        RECT 52.580 141.450 52.730 149.650 ;
        RECT 53.180 141.450 53.330 149.650 ;
        RECT 53.780 141.450 53.930 149.650 ;
        RECT 54.380 141.450 55.080 158.550 ;
        RECT 55.530 150.350 55.680 158.550 ;
        RECT 56.130 150.350 56.280 158.550 ;
        RECT 56.730 150.350 56.880 158.550 ;
        RECT 57.330 150.350 57.480 158.550 ;
        RECT 57.930 150.350 58.080 158.550 ;
        RECT 58.530 150.350 58.680 158.550 ;
        RECT 59.130 158.000 62.930 158.550 ;
        RECT 66.530 158.550 82.930 158.600 ;
        RECT 66.530 158.000 70.330 158.550 ;
        RECT 59.130 157.550 59.430 158.000 ;
        RECT 70.030 157.550 70.330 158.000 ;
        RECT 59.130 157.400 62.980 157.550 ;
        RECT 66.480 157.400 70.330 157.550 ;
        RECT 59.130 156.950 59.430 157.400 ;
        RECT 70.030 156.950 70.330 157.400 ;
        RECT 59.130 156.800 62.980 156.950 ;
        RECT 66.480 156.800 70.330 156.950 ;
        RECT 59.130 156.350 59.430 156.800 ;
        RECT 70.030 156.350 70.330 156.800 ;
        RECT 59.130 156.200 62.980 156.350 ;
        RECT 66.480 156.200 70.330 156.350 ;
        RECT 59.130 155.750 59.430 156.200 ;
        RECT 70.030 155.750 70.330 156.200 ;
        RECT 59.130 155.600 62.980 155.750 ;
        RECT 66.480 155.600 70.330 155.750 ;
        RECT 59.130 155.150 59.430 155.600 ;
        RECT 70.030 155.150 70.330 155.600 ;
        RECT 59.130 155.000 62.980 155.150 ;
        RECT 66.480 155.000 70.330 155.150 ;
        RECT 59.130 154.550 59.430 155.000 ;
        RECT 70.030 154.550 70.330 155.000 ;
        RECT 59.130 154.400 62.980 154.550 ;
        RECT 66.480 154.400 70.330 154.550 ;
        RECT 59.130 153.950 59.430 154.400 ;
        RECT 70.030 153.950 70.330 154.400 ;
        RECT 59.130 153.800 62.980 153.950 ;
        RECT 66.480 153.800 70.330 153.950 ;
        RECT 59.130 153.350 59.430 153.800 ;
        RECT 70.030 153.350 70.330 153.800 ;
        RECT 59.130 153.200 62.980 153.350 ;
        RECT 66.480 153.200 70.330 153.350 ;
        RECT 59.130 152.750 59.430 153.200 ;
        RECT 59.130 152.600 62.980 152.750 ;
        RECT 59.130 152.150 59.430 152.600 ;
        RECT 59.130 152.000 62.980 152.150 ;
        RECT 59.130 151.550 59.430 152.000 ;
        RECT 59.130 151.400 62.980 151.550 ;
        RECT 59.130 150.950 59.430 151.400 ;
        RECT 59.130 150.800 62.980 150.950 ;
        RECT 59.130 150.350 59.430 150.800 ;
        RECT 55.530 141.450 55.680 149.650 ;
        RECT 56.130 141.450 56.280 149.650 ;
        RECT 56.730 141.450 56.880 149.650 ;
        RECT 57.330 141.450 57.480 149.650 ;
        RECT 57.930 141.450 58.080 149.650 ;
        RECT 58.530 141.450 58.680 149.650 ;
        RECT 59.130 149.200 59.430 149.650 ;
        RECT 59.130 149.050 62.980 149.200 ;
        RECT 59.130 148.600 59.430 149.050 ;
        RECT 59.130 148.450 62.980 148.600 ;
        RECT 59.130 148.000 59.430 148.450 ;
        RECT 59.130 147.850 62.980 148.000 ;
        RECT 59.130 147.400 59.430 147.850 ;
        RECT 59.130 147.250 62.980 147.400 ;
        RECT 59.130 146.800 59.430 147.250 ;
        RECT 63.830 146.800 65.630 153.200 ;
        RECT 70.030 152.750 70.330 153.200 ;
        RECT 66.480 152.600 70.330 152.750 ;
        RECT 70.030 152.150 70.330 152.600 ;
        RECT 66.480 152.000 70.330 152.150 ;
        RECT 70.030 151.550 70.330 152.000 ;
        RECT 66.480 151.400 70.330 151.550 ;
        RECT 70.030 150.950 70.330 151.400 ;
        RECT 66.480 150.800 70.330 150.950 ;
        RECT 70.030 150.350 70.330 150.800 ;
        RECT 70.780 150.350 70.930 158.550 ;
        RECT 71.380 150.350 71.530 158.550 ;
        RECT 71.980 150.350 72.130 158.550 ;
        RECT 72.580 150.350 72.730 158.550 ;
        RECT 73.180 150.350 73.330 158.550 ;
        RECT 73.780 150.350 73.930 158.550 ;
        RECT 70.030 149.200 70.330 149.650 ;
        RECT 66.480 149.050 70.330 149.200 ;
        RECT 70.030 148.600 70.330 149.050 ;
        RECT 66.480 148.450 70.330 148.600 ;
        RECT 70.030 148.000 70.330 148.450 ;
        RECT 66.480 147.850 70.330 148.000 ;
        RECT 70.030 147.400 70.330 147.850 ;
        RECT 66.480 147.250 70.330 147.400 ;
        RECT 70.030 146.800 70.330 147.250 ;
        RECT 59.130 146.650 62.980 146.800 ;
        RECT 66.480 146.650 70.330 146.800 ;
        RECT 59.130 146.200 59.430 146.650 ;
        RECT 70.030 146.200 70.330 146.650 ;
        RECT 59.130 146.050 62.980 146.200 ;
        RECT 66.480 146.050 70.330 146.200 ;
        RECT 59.130 145.600 59.430 146.050 ;
        RECT 70.030 145.600 70.330 146.050 ;
        RECT 59.130 145.450 62.980 145.600 ;
        RECT 66.480 145.450 70.330 145.600 ;
        RECT 59.130 145.000 59.430 145.450 ;
        RECT 70.030 145.000 70.330 145.450 ;
        RECT 59.130 144.850 62.980 145.000 ;
        RECT 66.480 144.850 70.330 145.000 ;
        RECT 59.130 144.400 59.430 144.850 ;
        RECT 70.030 144.400 70.330 144.850 ;
        RECT 59.130 144.250 62.980 144.400 ;
        RECT 66.480 144.250 70.330 144.400 ;
        RECT 59.130 143.800 59.430 144.250 ;
        RECT 70.030 143.800 70.330 144.250 ;
        RECT 59.130 143.650 62.980 143.800 ;
        RECT 66.480 143.650 70.330 143.800 ;
        RECT 59.130 143.200 59.430 143.650 ;
        RECT 70.030 143.200 70.330 143.650 ;
        RECT 59.130 143.050 62.980 143.200 ;
        RECT 66.480 143.050 70.330 143.200 ;
        RECT 59.130 142.600 59.430 143.050 ;
        RECT 70.030 142.600 70.330 143.050 ;
        RECT 59.130 142.450 62.980 142.600 ;
        RECT 66.480 142.450 70.330 142.600 ;
        RECT 59.130 142.000 59.430 142.450 ;
        RECT 70.030 142.000 70.330 142.450 ;
        RECT 59.130 141.450 62.930 142.000 ;
        RECT 46.530 141.400 62.930 141.450 ;
        RECT 66.530 141.450 70.330 142.000 ;
        RECT 70.780 141.450 70.930 149.650 ;
        RECT 71.380 141.450 71.530 149.650 ;
        RECT 71.980 141.450 72.130 149.650 ;
        RECT 72.580 141.450 72.730 149.650 ;
        RECT 73.180 141.450 73.330 149.650 ;
        RECT 73.780 141.450 73.930 149.650 ;
        RECT 74.380 141.450 75.080 158.550 ;
        RECT 75.530 150.350 75.680 158.550 ;
        RECT 76.130 150.350 76.280 158.550 ;
        RECT 76.730 150.350 76.880 158.550 ;
        RECT 77.330 150.350 77.480 158.550 ;
        RECT 77.930 150.350 78.080 158.550 ;
        RECT 78.530 150.350 78.680 158.550 ;
        RECT 79.130 158.000 82.930 158.550 ;
        RECT 86.530 158.550 102.930 158.600 ;
        RECT 86.530 158.000 90.330 158.550 ;
        RECT 79.130 157.550 79.430 158.000 ;
        RECT 90.030 157.550 90.330 158.000 ;
        RECT 79.130 157.400 82.980 157.550 ;
        RECT 86.480 157.400 90.330 157.550 ;
        RECT 79.130 156.950 79.430 157.400 ;
        RECT 90.030 156.950 90.330 157.400 ;
        RECT 79.130 156.800 82.980 156.950 ;
        RECT 86.480 156.800 90.330 156.950 ;
        RECT 79.130 156.350 79.430 156.800 ;
        RECT 90.030 156.350 90.330 156.800 ;
        RECT 79.130 156.200 82.980 156.350 ;
        RECT 86.480 156.200 90.330 156.350 ;
        RECT 79.130 155.750 79.430 156.200 ;
        RECT 90.030 155.750 90.330 156.200 ;
        RECT 79.130 155.600 82.980 155.750 ;
        RECT 86.480 155.600 90.330 155.750 ;
        RECT 79.130 155.150 79.430 155.600 ;
        RECT 90.030 155.150 90.330 155.600 ;
        RECT 79.130 155.000 82.980 155.150 ;
        RECT 86.480 155.000 90.330 155.150 ;
        RECT 79.130 154.550 79.430 155.000 ;
        RECT 90.030 154.550 90.330 155.000 ;
        RECT 79.130 154.400 82.980 154.550 ;
        RECT 86.480 154.400 90.330 154.550 ;
        RECT 79.130 153.950 79.430 154.400 ;
        RECT 90.030 153.950 90.330 154.400 ;
        RECT 79.130 153.800 82.980 153.950 ;
        RECT 86.480 153.800 90.330 153.950 ;
        RECT 79.130 153.350 79.430 153.800 ;
        RECT 90.030 153.350 90.330 153.800 ;
        RECT 79.130 153.200 82.980 153.350 ;
        RECT 86.480 153.200 90.330 153.350 ;
        RECT 79.130 152.750 79.430 153.200 ;
        RECT 79.130 152.600 82.980 152.750 ;
        RECT 79.130 152.150 79.430 152.600 ;
        RECT 79.130 152.000 82.980 152.150 ;
        RECT 79.130 151.550 79.430 152.000 ;
        RECT 79.130 151.400 82.980 151.550 ;
        RECT 79.130 150.950 79.430 151.400 ;
        RECT 79.130 150.800 82.980 150.950 ;
        RECT 79.130 150.350 79.430 150.800 ;
        RECT 75.530 141.450 75.680 149.650 ;
        RECT 76.130 141.450 76.280 149.650 ;
        RECT 76.730 141.450 76.880 149.650 ;
        RECT 77.330 141.450 77.480 149.650 ;
        RECT 77.930 141.450 78.080 149.650 ;
        RECT 78.530 141.450 78.680 149.650 ;
        RECT 79.130 149.200 79.430 149.650 ;
        RECT 79.130 149.050 82.980 149.200 ;
        RECT 79.130 148.600 79.430 149.050 ;
        RECT 79.130 148.450 82.980 148.600 ;
        RECT 79.130 148.000 79.430 148.450 ;
        RECT 79.130 147.850 82.980 148.000 ;
        RECT 79.130 147.400 79.430 147.850 ;
        RECT 79.130 147.250 82.980 147.400 ;
        RECT 79.130 146.800 79.430 147.250 ;
        RECT 83.830 146.800 85.630 153.200 ;
        RECT 90.030 152.750 90.330 153.200 ;
        RECT 86.480 152.600 90.330 152.750 ;
        RECT 90.030 152.150 90.330 152.600 ;
        RECT 86.480 152.000 90.330 152.150 ;
        RECT 90.030 151.550 90.330 152.000 ;
        RECT 86.480 151.400 90.330 151.550 ;
        RECT 90.030 150.950 90.330 151.400 ;
        RECT 86.480 150.800 90.330 150.950 ;
        RECT 90.030 150.350 90.330 150.800 ;
        RECT 90.780 150.350 90.930 158.550 ;
        RECT 91.380 150.350 91.530 158.550 ;
        RECT 91.980 150.350 92.130 158.550 ;
        RECT 92.580 150.350 92.730 158.550 ;
        RECT 93.180 150.350 93.330 158.550 ;
        RECT 93.780 150.350 93.930 158.550 ;
        RECT 90.030 149.200 90.330 149.650 ;
        RECT 86.480 149.050 90.330 149.200 ;
        RECT 90.030 148.600 90.330 149.050 ;
        RECT 86.480 148.450 90.330 148.600 ;
        RECT 90.030 148.000 90.330 148.450 ;
        RECT 86.480 147.850 90.330 148.000 ;
        RECT 90.030 147.400 90.330 147.850 ;
        RECT 86.480 147.250 90.330 147.400 ;
        RECT 90.030 146.800 90.330 147.250 ;
        RECT 79.130 146.650 82.980 146.800 ;
        RECT 86.480 146.650 90.330 146.800 ;
        RECT 79.130 146.200 79.430 146.650 ;
        RECT 90.030 146.200 90.330 146.650 ;
        RECT 79.130 146.050 82.980 146.200 ;
        RECT 86.480 146.050 90.330 146.200 ;
        RECT 79.130 145.600 79.430 146.050 ;
        RECT 90.030 145.600 90.330 146.050 ;
        RECT 79.130 145.450 82.980 145.600 ;
        RECT 86.480 145.450 90.330 145.600 ;
        RECT 79.130 145.000 79.430 145.450 ;
        RECT 90.030 145.000 90.330 145.450 ;
        RECT 79.130 144.850 82.980 145.000 ;
        RECT 86.480 144.850 90.330 145.000 ;
        RECT 79.130 144.400 79.430 144.850 ;
        RECT 90.030 144.400 90.330 144.850 ;
        RECT 79.130 144.250 82.980 144.400 ;
        RECT 86.480 144.250 90.330 144.400 ;
        RECT 79.130 143.800 79.430 144.250 ;
        RECT 90.030 143.800 90.330 144.250 ;
        RECT 79.130 143.650 82.980 143.800 ;
        RECT 86.480 143.650 90.330 143.800 ;
        RECT 79.130 143.200 79.430 143.650 ;
        RECT 90.030 143.200 90.330 143.650 ;
        RECT 79.130 143.050 82.980 143.200 ;
        RECT 86.480 143.050 90.330 143.200 ;
        RECT 79.130 142.600 79.430 143.050 ;
        RECT 90.030 142.600 90.330 143.050 ;
        RECT 79.130 142.450 82.980 142.600 ;
        RECT 86.480 142.450 90.330 142.600 ;
        RECT 79.130 142.000 79.430 142.450 ;
        RECT 90.030 142.000 90.330 142.450 ;
        RECT 79.130 141.450 82.930 142.000 ;
        RECT 66.530 141.400 82.930 141.450 ;
        RECT 86.530 141.450 90.330 142.000 ;
        RECT 90.780 141.450 90.930 149.650 ;
        RECT 91.380 141.450 91.530 149.650 ;
        RECT 91.980 141.450 92.130 149.650 ;
        RECT 92.580 141.450 92.730 149.650 ;
        RECT 93.180 141.450 93.330 149.650 ;
        RECT 93.780 141.450 93.930 149.650 ;
        RECT 94.380 141.450 95.080 158.550 ;
        RECT 95.530 150.350 95.680 158.550 ;
        RECT 96.130 150.350 96.280 158.550 ;
        RECT 96.730 150.350 96.880 158.550 ;
        RECT 97.330 150.350 97.480 158.550 ;
        RECT 97.930 150.350 98.080 158.550 ;
        RECT 98.530 150.350 98.680 158.550 ;
        RECT 99.130 158.000 102.930 158.550 ;
        RECT 99.130 157.550 99.430 158.000 ;
        RECT 99.130 157.400 102.980 157.550 ;
        RECT 99.130 156.950 99.430 157.400 ;
        RECT 99.130 156.800 102.980 156.950 ;
        RECT 99.130 156.350 99.430 156.800 ;
        RECT 99.130 156.200 102.980 156.350 ;
        RECT 99.130 155.750 99.430 156.200 ;
        RECT 99.130 155.600 102.980 155.750 ;
        RECT 99.130 155.150 99.430 155.600 ;
        RECT 99.130 155.000 102.980 155.150 ;
        RECT 99.130 154.550 99.430 155.000 ;
        RECT 99.130 154.400 102.980 154.550 ;
        RECT 99.130 153.950 99.430 154.400 ;
        RECT 99.130 153.800 102.980 153.950 ;
        RECT 99.130 153.350 99.430 153.800 ;
        RECT 99.130 153.200 102.980 153.350 ;
        RECT 99.130 152.750 99.430 153.200 ;
        RECT 99.130 152.600 102.980 152.750 ;
        RECT 99.130 152.150 99.430 152.600 ;
        RECT 99.130 152.000 102.980 152.150 ;
        RECT 99.130 151.550 99.430 152.000 ;
        RECT 99.130 151.400 102.980 151.550 ;
        RECT 99.130 150.950 99.430 151.400 ;
        RECT 99.130 150.800 102.980 150.950 ;
        RECT 99.130 150.350 99.430 150.800 ;
        RECT 95.530 141.450 95.680 149.650 ;
        RECT 96.130 141.450 96.280 149.650 ;
        RECT 96.730 141.450 96.880 149.650 ;
        RECT 97.330 141.450 97.480 149.650 ;
        RECT 97.930 141.450 98.080 149.650 ;
        RECT 98.530 141.450 98.680 149.650 ;
        RECT 99.130 149.200 99.430 149.650 ;
        RECT 99.130 149.050 102.980 149.200 ;
        RECT 99.130 148.600 99.430 149.050 ;
        RECT 99.130 148.450 102.980 148.600 ;
        RECT 99.130 148.000 99.430 148.450 ;
        RECT 99.130 147.850 102.980 148.000 ;
        RECT 99.130 147.400 99.430 147.850 ;
        RECT 99.130 147.250 102.980 147.400 ;
        RECT 99.130 146.800 99.430 147.250 ;
        RECT 103.830 146.800 104.730 153.200 ;
        RECT 109.850 149.500 111.850 150.775 ;
        RECT 99.130 146.650 102.980 146.800 ;
        RECT 99.130 146.200 99.430 146.650 ;
        RECT 99.130 146.050 102.980 146.200 ;
        RECT 99.130 145.600 99.430 146.050 ;
        RECT 99.130 145.450 102.980 145.600 ;
        RECT 99.130 145.000 99.430 145.450 ;
        RECT 99.130 144.850 102.980 145.000 ;
        RECT 99.130 144.400 99.430 144.850 ;
        RECT 99.130 144.250 102.980 144.400 ;
        RECT 99.130 143.800 99.430 144.250 ;
        RECT 99.130 143.650 102.980 143.800 ;
        RECT 99.130 143.200 99.430 143.650 ;
        RECT 99.130 143.050 102.980 143.200 ;
        RECT 99.130 142.600 99.430 143.050 ;
        RECT 99.130 142.450 102.980 142.600 ;
        RECT 99.130 142.000 99.430 142.450 ;
        RECT 99.130 141.450 102.930 142.000 ;
        RECT 86.530 141.400 102.930 141.450 ;
        RECT 9.630 140.900 19.830 141.400 ;
        RECT 29.630 140.900 39.830 141.400 ;
        RECT 49.630 140.900 59.830 141.400 ;
        RECT 69.630 140.900 79.830 141.400 ;
        RECT 89.630 140.900 99.830 141.400 ;
        RECT 11.530 139.100 17.930 140.900 ;
        RECT 31.530 139.100 37.930 140.900 ;
        RECT 51.530 139.100 57.930 140.900 ;
        RECT 71.530 139.100 77.930 140.900 ;
        RECT 91.530 139.100 97.930 140.900 ;
        RECT 9.630 138.600 19.830 139.100 ;
        RECT 29.630 138.600 39.830 139.100 ;
        RECT 49.630 138.600 59.830 139.100 ;
        RECT 69.630 138.600 79.830 139.100 ;
        RECT 89.630 138.600 99.830 139.100 ;
        RECT 6.530 138.550 22.930 138.600 ;
        RECT 6.530 138.000 10.330 138.550 ;
        RECT 10.030 137.550 10.330 138.000 ;
        RECT 6.480 137.400 10.330 137.550 ;
        RECT 10.030 136.950 10.330 137.400 ;
        RECT 6.480 136.800 10.330 136.950 ;
        RECT 10.030 136.350 10.330 136.800 ;
        RECT 6.480 136.200 10.330 136.350 ;
        RECT 10.030 135.750 10.330 136.200 ;
        RECT 6.480 135.600 10.330 135.750 ;
        RECT 10.030 135.150 10.330 135.600 ;
        RECT 6.480 135.000 10.330 135.150 ;
        RECT 10.030 134.550 10.330 135.000 ;
        RECT 6.480 134.400 10.330 134.550 ;
        RECT 10.030 133.950 10.330 134.400 ;
        RECT 6.480 133.800 10.330 133.950 ;
        RECT 10.030 133.350 10.330 133.800 ;
        RECT 6.480 133.200 10.330 133.350 ;
        RECT 4.730 126.800 5.630 133.200 ;
        RECT 10.030 132.750 10.330 133.200 ;
        RECT 6.480 132.600 10.330 132.750 ;
        RECT 10.030 132.150 10.330 132.600 ;
        RECT 6.480 132.000 10.330 132.150 ;
        RECT 10.030 131.550 10.330 132.000 ;
        RECT 6.480 131.400 10.330 131.550 ;
        RECT 10.030 130.950 10.330 131.400 ;
        RECT 6.480 130.800 10.330 130.950 ;
        RECT 10.030 130.350 10.330 130.800 ;
        RECT 10.780 130.350 10.930 138.550 ;
        RECT 11.380 130.350 11.530 138.550 ;
        RECT 11.980 130.350 12.130 138.550 ;
        RECT 12.580 130.350 12.730 138.550 ;
        RECT 13.180 130.350 13.330 138.550 ;
        RECT 13.780 130.350 13.930 138.550 ;
        RECT 10.030 129.200 10.330 129.650 ;
        RECT 6.480 129.050 10.330 129.200 ;
        RECT 10.030 128.600 10.330 129.050 ;
        RECT 6.480 128.450 10.330 128.600 ;
        RECT 10.030 128.000 10.330 128.450 ;
        RECT 6.480 127.850 10.330 128.000 ;
        RECT 10.030 127.400 10.330 127.850 ;
        RECT 6.480 127.250 10.330 127.400 ;
        RECT 10.030 126.800 10.330 127.250 ;
        RECT 6.480 126.650 10.330 126.800 ;
        RECT 10.030 126.200 10.330 126.650 ;
        RECT 6.480 126.050 10.330 126.200 ;
        RECT 10.030 125.600 10.330 126.050 ;
        RECT 6.480 125.450 10.330 125.600 ;
        RECT 10.030 125.000 10.330 125.450 ;
        RECT 6.480 124.850 10.330 125.000 ;
        RECT 10.030 124.400 10.330 124.850 ;
        RECT 6.480 124.250 10.330 124.400 ;
        RECT 10.030 123.800 10.330 124.250 ;
        RECT 6.480 123.650 10.330 123.800 ;
        RECT 10.030 123.200 10.330 123.650 ;
        RECT 6.480 123.050 10.330 123.200 ;
        RECT 10.030 122.600 10.330 123.050 ;
        RECT 6.480 122.450 10.330 122.600 ;
        RECT 10.030 122.000 10.330 122.450 ;
        RECT 6.530 121.450 10.330 122.000 ;
        RECT 10.780 121.450 10.930 129.650 ;
        RECT 11.380 121.450 11.530 129.650 ;
        RECT 11.980 121.450 12.130 129.650 ;
        RECT 12.580 121.450 12.730 129.650 ;
        RECT 13.180 121.450 13.330 129.650 ;
        RECT 13.780 121.450 13.930 129.650 ;
        RECT 14.380 121.450 15.080 138.550 ;
        RECT 15.530 130.350 15.680 138.550 ;
        RECT 16.130 130.350 16.280 138.550 ;
        RECT 16.730 130.350 16.880 138.550 ;
        RECT 17.330 130.350 17.480 138.550 ;
        RECT 17.930 130.350 18.080 138.550 ;
        RECT 18.530 130.350 18.680 138.550 ;
        RECT 19.130 138.000 22.930 138.550 ;
        RECT 26.530 138.550 42.930 138.600 ;
        RECT 26.530 138.000 30.330 138.550 ;
        RECT 19.130 137.550 19.430 138.000 ;
        RECT 30.030 137.550 30.330 138.000 ;
        RECT 19.130 137.400 22.980 137.550 ;
        RECT 26.480 137.400 30.330 137.550 ;
        RECT 19.130 136.950 19.430 137.400 ;
        RECT 30.030 136.950 30.330 137.400 ;
        RECT 19.130 136.800 22.980 136.950 ;
        RECT 26.480 136.800 30.330 136.950 ;
        RECT 19.130 136.350 19.430 136.800 ;
        RECT 30.030 136.350 30.330 136.800 ;
        RECT 19.130 136.200 22.980 136.350 ;
        RECT 26.480 136.200 30.330 136.350 ;
        RECT 19.130 135.750 19.430 136.200 ;
        RECT 30.030 135.750 30.330 136.200 ;
        RECT 19.130 135.600 22.980 135.750 ;
        RECT 26.480 135.600 30.330 135.750 ;
        RECT 19.130 135.150 19.430 135.600 ;
        RECT 30.030 135.150 30.330 135.600 ;
        RECT 19.130 135.000 22.980 135.150 ;
        RECT 26.480 135.000 30.330 135.150 ;
        RECT 19.130 134.550 19.430 135.000 ;
        RECT 30.030 134.550 30.330 135.000 ;
        RECT 19.130 134.400 22.980 134.550 ;
        RECT 26.480 134.400 30.330 134.550 ;
        RECT 19.130 133.950 19.430 134.400 ;
        RECT 30.030 133.950 30.330 134.400 ;
        RECT 19.130 133.800 22.980 133.950 ;
        RECT 26.480 133.800 30.330 133.950 ;
        RECT 19.130 133.350 19.430 133.800 ;
        RECT 30.030 133.350 30.330 133.800 ;
        RECT 19.130 133.200 22.980 133.350 ;
        RECT 26.480 133.200 30.330 133.350 ;
        RECT 19.130 132.750 19.430 133.200 ;
        RECT 19.130 132.600 22.980 132.750 ;
        RECT 19.130 132.150 19.430 132.600 ;
        RECT 19.130 132.000 22.980 132.150 ;
        RECT 19.130 131.550 19.430 132.000 ;
        RECT 19.130 131.400 22.980 131.550 ;
        RECT 19.130 130.950 19.430 131.400 ;
        RECT 19.130 130.800 22.980 130.950 ;
        RECT 19.130 130.350 19.430 130.800 ;
        RECT 15.530 121.450 15.680 129.650 ;
        RECT 16.130 121.450 16.280 129.650 ;
        RECT 16.730 121.450 16.880 129.650 ;
        RECT 17.330 121.450 17.480 129.650 ;
        RECT 17.930 121.450 18.080 129.650 ;
        RECT 18.530 121.450 18.680 129.650 ;
        RECT 19.130 129.200 19.430 129.650 ;
        RECT 19.130 129.050 22.980 129.200 ;
        RECT 19.130 128.600 19.430 129.050 ;
        RECT 19.130 128.450 22.980 128.600 ;
        RECT 19.130 128.000 19.430 128.450 ;
        RECT 19.130 127.850 22.980 128.000 ;
        RECT 19.130 127.400 19.430 127.850 ;
        RECT 19.130 127.250 22.980 127.400 ;
        RECT 19.130 126.800 19.430 127.250 ;
        RECT 23.830 126.800 25.630 133.200 ;
        RECT 30.030 132.750 30.330 133.200 ;
        RECT 26.480 132.600 30.330 132.750 ;
        RECT 30.030 132.150 30.330 132.600 ;
        RECT 26.480 132.000 30.330 132.150 ;
        RECT 30.030 131.550 30.330 132.000 ;
        RECT 26.480 131.400 30.330 131.550 ;
        RECT 30.030 130.950 30.330 131.400 ;
        RECT 26.480 130.800 30.330 130.950 ;
        RECT 30.030 130.350 30.330 130.800 ;
        RECT 30.780 130.350 30.930 138.550 ;
        RECT 31.380 130.350 31.530 138.550 ;
        RECT 31.980 130.350 32.130 138.550 ;
        RECT 32.580 130.350 32.730 138.550 ;
        RECT 33.180 130.350 33.330 138.550 ;
        RECT 33.780 130.350 33.930 138.550 ;
        RECT 30.030 129.200 30.330 129.650 ;
        RECT 26.480 129.050 30.330 129.200 ;
        RECT 30.030 128.600 30.330 129.050 ;
        RECT 26.480 128.450 30.330 128.600 ;
        RECT 30.030 128.000 30.330 128.450 ;
        RECT 26.480 127.850 30.330 128.000 ;
        RECT 30.030 127.400 30.330 127.850 ;
        RECT 26.480 127.250 30.330 127.400 ;
        RECT 30.030 126.800 30.330 127.250 ;
        RECT 19.130 126.650 22.980 126.800 ;
        RECT 26.480 126.650 30.330 126.800 ;
        RECT 19.130 126.200 19.430 126.650 ;
        RECT 30.030 126.200 30.330 126.650 ;
        RECT 19.130 126.050 22.980 126.200 ;
        RECT 26.480 126.050 30.330 126.200 ;
        RECT 19.130 125.600 19.430 126.050 ;
        RECT 30.030 125.600 30.330 126.050 ;
        RECT 19.130 125.450 22.980 125.600 ;
        RECT 26.480 125.450 30.330 125.600 ;
        RECT 19.130 125.000 19.430 125.450 ;
        RECT 30.030 125.000 30.330 125.450 ;
        RECT 19.130 124.850 22.980 125.000 ;
        RECT 26.480 124.850 30.330 125.000 ;
        RECT 19.130 124.400 19.430 124.850 ;
        RECT 30.030 124.400 30.330 124.850 ;
        RECT 19.130 124.250 22.980 124.400 ;
        RECT 26.480 124.250 30.330 124.400 ;
        RECT 19.130 123.800 19.430 124.250 ;
        RECT 30.030 123.800 30.330 124.250 ;
        RECT 19.130 123.650 22.980 123.800 ;
        RECT 26.480 123.650 30.330 123.800 ;
        RECT 19.130 123.200 19.430 123.650 ;
        RECT 30.030 123.200 30.330 123.650 ;
        RECT 19.130 123.050 22.980 123.200 ;
        RECT 26.480 123.050 30.330 123.200 ;
        RECT 19.130 122.600 19.430 123.050 ;
        RECT 30.030 122.600 30.330 123.050 ;
        RECT 19.130 122.450 22.980 122.600 ;
        RECT 26.480 122.450 30.330 122.600 ;
        RECT 19.130 122.000 19.430 122.450 ;
        RECT 30.030 122.000 30.330 122.450 ;
        RECT 19.130 121.450 22.930 122.000 ;
        RECT 6.530 121.400 22.930 121.450 ;
        RECT 26.530 121.450 30.330 122.000 ;
        RECT 30.780 121.450 30.930 129.650 ;
        RECT 31.380 121.450 31.530 129.650 ;
        RECT 31.980 121.450 32.130 129.650 ;
        RECT 32.580 121.450 32.730 129.650 ;
        RECT 33.180 121.450 33.330 129.650 ;
        RECT 33.780 121.450 33.930 129.650 ;
        RECT 34.380 121.450 35.080 138.550 ;
        RECT 35.530 130.350 35.680 138.550 ;
        RECT 36.130 130.350 36.280 138.550 ;
        RECT 36.730 130.350 36.880 138.550 ;
        RECT 37.330 130.350 37.480 138.550 ;
        RECT 37.930 130.350 38.080 138.550 ;
        RECT 38.530 130.350 38.680 138.550 ;
        RECT 39.130 138.000 42.930 138.550 ;
        RECT 46.530 138.550 62.930 138.600 ;
        RECT 46.530 138.000 50.330 138.550 ;
        RECT 39.130 137.550 39.430 138.000 ;
        RECT 50.030 137.550 50.330 138.000 ;
        RECT 39.130 137.400 42.980 137.550 ;
        RECT 46.480 137.400 50.330 137.550 ;
        RECT 39.130 136.950 39.430 137.400 ;
        RECT 50.030 136.950 50.330 137.400 ;
        RECT 39.130 136.800 42.980 136.950 ;
        RECT 46.480 136.800 50.330 136.950 ;
        RECT 39.130 136.350 39.430 136.800 ;
        RECT 50.030 136.350 50.330 136.800 ;
        RECT 39.130 136.200 42.980 136.350 ;
        RECT 46.480 136.200 50.330 136.350 ;
        RECT 39.130 135.750 39.430 136.200 ;
        RECT 50.030 135.750 50.330 136.200 ;
        RECT 39.130 135.600 42.980 135.750 ;
        RECT 46.480 135.600 50.330 135.750 ;
        RECT 39.130 135.150 39.430 135.600 ;
        RECT 50.030 135.150 50.330 135.600 ;
        RECT 39.130 135.000 42.980 135.150 ;
        RECT 46.480 135.000 50.330 135.150 ;
        RECT 39.130 134.550 39.430 135.000 ;
        RECT 50.030 134.550 50.330 135.000 ;
        RECT 39.130 134.400 42.980 134.550 ;
        RECT 46.480 134.400 50.330 134.550 ;
        RECT 39.130 133.950 39.430 134.400 ;
        RECT 50.030 133.950 50.330 134.400 ;
        RECT 39.130 133.800 42.980 133.950 ;
        RECT 46.480 133.800 50.330 133.950 ;
        RECT 39.130 133.350 39.430 133.800 ;
        RECT 50.030 133.350 50.330 133.800 ;
        RECT 39.130 133.200 42.980 133.350 ;
        RECT 46.480 133.200 50.330 133.350 ;
        RECT 39.130 132.750 39.430 133.200 ;
        RECT 39.130 132.600 42.980 132.750 ;
        RECT 39.130 132.150 39.430 132.600 ;
        RECT 39.130 132.000 42.980 132.150 ;
        RECT 39.130 131.550 39.430 132.000 ;
        RECT 39.130 131.400 42.980 131.550 ;
        RECT 39.130 130.950 39.430 131.400 ;
        RECT 39.130 130.800 42.980 130.950 ;
        RECT 39.130 130.350 39.430 130.800 ;
        RECT 35.530 121.450 35.680 129.650 ;
        RECT 36.130 121.450 36.280 129.650 ;
        RECT 36.730 121.450 36.880 129.650 ;
        RECT 37.330 121.450 37.480 129.650 ;
        RECT 37.930 121.450 38.080 129.650 ;
        RECT 38.530 121.450 38.680 129.650 ;
        RECT 39.130 129.200 39.430 129.650 ;
        RECT 39.130 129.050 42.980 129.200 ;
        RECT 39.130 128.600 39.430 129.050 ;
        RECT 39.130 128.450 42.980 128.600 ;
        RECT 39.130 128.000 39.430 128.450 ;
        RECT 39.130 127.850 42.980 128.000 ;
        RECT 39.130 127.400 39.430 127.850 ;
        RECT 39.130 127.250 42.980 127.400 ;
        RECT 39.130 126.800 39.430 127.250 ;
        RECT 43.830 126.800 45.630 133.200 ;
        RECT 50.030 132.750 50.330 133.200 ;
        RECT 46.480 132.600 50.330 132.750 ;
        RECT 50.030 132.150 50.330 132.600 ;
        RECT 46.480 132.000 50.330 132.150 ;
        RECT 50.030 131.550 50.330 132.000 ;
        RECT 46.480 131.400 50.330 131.550 ;
        RECT 50.030 130.950 50.330 131.400 ;
        RECT 46.480 130.800 50.330 130.950 ;
        RECT 50.030 130.350 50.330 130.800 ;
        RECT 50.780 130.350 50.930 138.550 ;
        RECT 51.380 130.350 51.530 138.550 ;
        RECT 51.980 130.350 52.130 138.550 ;
        RECT 52.580 130.350 52.730 138.550 ;
        RECT 53.180 130.350 53.330 138.550 ;
        RECT 53.780 130.350 53.930 138.550 ;
        RECT 50.030 129.200 50.330 129.650 ;
        RECT 46.480 129.050 50.330 129.200 ;
        RECT 50.030 128.600 50.330 129.050 ;
        RECT 46.480 128.450 50.330 128.600 ;
        RECT 50.030 128.000 50.330 128.450 ;
        RECT 46.480 127.850 50.330 128.000 ;
        RECT 50.030 127.400 50.330 127.850 ;
        RECT 46.480 127.250 50.330 127.400 ;
        RECT 50.030 126.800 50.330 127.250 ;
        RECT 39.130 126.650 42.980 126.800 ;
        RECT 46.480 126.650 50.330 126.800 ;
        RECT 39.130 126.200 39.430 126.650 ;
        RECT 50.030 126.200 50.330 126.650 ;
        RECT 39.130 126.050 42.980 126.200 ;
        RECT 46.480 126.050 50.330 126.200 ;
        RECT 39.130 125.600 39.430 126.050 ;
        RECT 50.030 125.600 50.330 126.050 ;
        RECT 39.130 125.450 42.980 125.600 ;
        RECT 46.480 125.450 50.330 125.600 ;
        RECT 39.130 125.000 39.430 125.450 ;
        RECT 50.030 125.000 50.330 125.450 ;
        RECT 39.130 124.850 42.980 125.000 ;
        RECT 46.480 124.850 50.330 125.000 ;
        RECT 39.130 124.400 39.430 124.850 ;
        RECT 50.030 124.400 50.330 124.850 ;
        RECT 39.130 124.250 42.980 124.400 ;
        RECT 46.480 124.250 50.330 124.400 ;
        RECT 39.130 123.800 39.430 124.250 ;
        RECT 50.030 123.800 50.330 124.250 ;
        RECT 39.130 123.650 42.980 123.800 ;
        RECT 46.480 123.650 50.330 123.800 ;
        RECT 39.130 123.200 39.430 123.650 ;
        RECT 50.030 123.200 50.330 123.650 ;
        RECT 39.130 123.050 42.980 123.200 ;
        RECT 46.480 123.050 50.330 123.200 ;
        RECT 39.130 122.600 39.430 123.050 ;
        RECT 50.030 122.600 50.330 123.050 ;
        RECT 39.130 122.450 42.980 122.600 ;
        RECT 46.480 122.450 50.330 122.600 ;
        RECT 39.130 122.000 39.430 122.450 ;
        RECT 50.030 122.000 50.330 122.450 ;
        RECT 39.130 121.450 42.930 122.000 ;
        RECT 26.530 121.400 42.930 121.450 ;
        RECT 46.530 121.450 50.330 122.000 ;
        RECT 50.780 121.450 50.930 129.650 ;
        RECT 51.380 121.450 51.530 129.650 ;
        RECT 51.980 121.450 52.130 129.650 ;
        RECT 52.580 121.450 52.730 129.650 ;
        RECT 53.180 121.450 53.330 129.650 ;
        RECT 53.780 121.450 53.930 129.650 ;
        RECT 54.380 121.450 55.080 138.550 ;
        RECT 55.530 130.350 55.680 138.550 ;
        RECT 56.130 130.350 56.280 138.550 ;
        RECT 56.730 130.350 56.880 138.550 ;
        RECT 57.330 130.350 57.480 138.550 ;
        RECT 57.930 130.350 58.080 138.550 ;
        RECT 58.530 130.350 58.680 138.550 ;
        RECT 59.130 138.000 62.930 138.550 ;
        RECT 66.530 138.550 82.930 138.600 ;
        RECT 66.530 138.000 70.330 138.550 ;
        RECT 59.130 137.550 59.430 138.000 ;
        RECT 70.030 137.550 70.330 138.000 ;
        RECT 59.130 137.400 62.980 137.550 ;
        RECT 66.480 137.400 70.330 137.550 ;
        RECT 59.130 136.950 59.430 137.400 ;
        RECT 70.030 136.950 70.330 137.400 ;
        RECT 59.130 136.800 62.980 136.950 ;
        RECT 66.480 136.800 70.330 136.950 ;
        RECT 59.130 136.350 59.430 136.800 ;
        RECT 70.030 136.350 70.330 136.800 ;
        RECT 59.130 136.200 62.980 136.350 ;
        RECT 66.480 136.200 70.330 136.350 ;
        RECT 59.130 135.750 59.430 136.200 ;
        RECT 70.030 135.750 70.330 136.200 ;
        RECT 59.130 135.600 62.980 135.750 ;
        RECT 66.480 135.600 70.330 135.750 ;
        RECT 59.130 135.150 59.430 135.600 ;
        RECT 70.030 135.150 70.330 135.600 ;
        RECT 59.130 135.000 62.980 135.150 ;
        RECT 66.480 135.000 70.330 135.150 ;
        RECT 59.130 134.550 59.430 135.000 ;
        RECT 70.030 134.550 70.330 135.000 ;
        RECT 59.130 134.400 62.980 134.550 ;
        RECT 66.480 134.400 70.330 134.550 ;
        RECT 59.130 133.950 59.430 134.400 ;
        RECT 70.030 133.950 70.330 134.400 ;
        RECT 59.130 133.800 62.980 133.950 ;
        RECT 66.480 133.800 70.330 133.950 ;
        RECT 59.130 133.350 59.430 133.800 ;
        RECT 70.030 133.350 70.330 133.800 ;
        RECT 59.130 133.200 62.980 133.350 ;
        RECT 66.480 133.200 70.330 133.350 ;
        RECT 59.130 132.750 59.430 133.200 ;
        RECT 59.130 132.600 62.980 132.750 ;
        RECT 59.130 132.150 59.430 132.600 ;
        RECT 59.130 132.000 62.980 132.150 ;
        RECT 59.130 131.550 59.430 132.000 ;
        RECT 59.130 131.400 62.980 131.550 ;
        RECT 59.130 130.950 59.430 131.400 ;
        RECT 59.130 130.800 62.980 130.950 ;
        RECT 59.130 130.350 59.430 130.800 ;
        RECT 55.530 121.450 55.680 129.650 ;
        RECT 56.130 121.450 56.280 129.650 ;
        RECT 56.730 121.450 56.880 129.650 ;
        RECT 57.330 121.450 57.480 129.650 ;
        RECT 57.930 121.450 58.080 129.650 ;
        RECT 58.530 121.450 58.680 129.650 ;
        RECT 59.130 129.200 59.430 129.650 ;
        RECT 59.130 129.050 62.980 129.200 ;
        RECT 59.130 128.600 59.430 129.050 ;
        RECT 59.130 128.450 62.980 128.600 ;
        RECT 59.130 128.000 59.430 128.450 ;
        RECT 59.130 127.850 62.980 128.000 ;
        RECT 59.130 127.400 59.430 127.850 ;
        RECT 59.130 127.250 62.980 127.400 ;
        RECT 59.130 126.800 59.430 127.250 ;
        RECT 63.830 126.800 65.630 133.200 ;
        RECT 70.030 132.750 70.330 133.200 ;
        RECT 66.480 132.600 70.330 132.750 ;
        RECT 70.030 132.150 70.330 132.600 ;
        RECT 66.480 132.000 70.330 132.150 ;
        RECT 70.030 131.550 70.330 132.000 ;
        RECT 66.480 131.400 70.330 131.550 ;
        RECT 70.030 130.950 70.330 131.400 ;
        RECT 66.480 130.800 70.330 130.950 ;
        RECT 70.030 130.350 70.330 130.800 ;
        RECT 70.780 130.350 70.930 138.550 ;
        RECT 71.380 130.350 71.530 138.550 ;
        RECT 71.980 130.350 72.130 138.550 ;
        RECT 72.580 130.350 72.730 138.550 ;
        RECT 73.180 130.350 73.330 138.550 ;
        RECT 73.780 130.350 73.930 138.550 ;
        RECT 70.030 129.200 70.330 129.650 ;
        RECT 66.480 129.050 70.330 129.200 ;
        RECT 70.030 128.600 70.330 129.050 ;
        RECT 66.480 128.450 70.330 128.600 ;
        RECT 70.030 128.000 70.330 128.450 ;
        RECT 66.480 127.850 70.330 128.000 ;
        RECT 70.030 127.400 70.330 127.850 ;
        RECT 66.480 127.250 70.330 127.400 ;
        RECT 70.030 126.800 70.330 127.250 ;
        RECT 59.130 126.650 62.980 126.800 ;
        RECT 66.480 126.650 70.330 126.800 ;
        RECT 59.130 126.200 59.430 126.650 ;
        RECT 70.030 126.200 70.330 126.650 ;
        RECT 59.130 126.050 62.980 126.200 ;
        RECT 66.480 126.050 70.330 126.200 ;
        RECT 59.130 125.600 59.430 126.050 ;
        RECT 70.030 125.600 70.330 126.050 ;
        RECT 59.130 125.450 62.980 125.600 ;
        RECT 66.480 125.450 70.330 125.600 ;
        RECT 59.130 125.000 59.430 125.450 ;
        RECT 70.030 125.000 70.330 125.450 ;
        RECT 59.130 124.850 62.980 125.000 ;
        RECT 66.480 124.850 70.330 125.000 ;
        RECT 59.130 124.400 59.430 124.850 ;
        RECT 70.030 124.400 70.330 124.850 ;
        RECT 59.130 124.250 62.980 124.400 ;
        RECT 66.480 124.250 70.330 124.400 ;
        RECT 59.130 123.800 59.430 124.250 ;
        RECT 70.030 123.800 70.330 124.250 ;
        RECT 59.130 123.650 62.980 123.800 ;
        RECT 66.480 123.650 70.330 123.800 ;
        RECT 59.130 123.200 59.430 123.650 ;
        RECT 70.030 123.200 70.330 123.650 ;
        RECT 59.130 123.050 62.980 123.200 ;
        RECT 66.480 123.050 70.330 123.200 ;
        RECT 59.130 122.600 59.430 123.050 ;
        RECT 70.030 122.600 70.330 123.050 ;
        RECT 59.130 122.450 62.980 122.600 ;
        RECT 66.480 122.450 70.330 122.600 ;
        RECT 59.130 122.000 59.430 122.450 ;
        RECT 70.030 122.000 70.330 122.450 ;
        RECT 59.130 121.450 62.930 122.000 ;
        RECT 46.530 121.400 62.930 121.450 ;
        RECT 66.530 121.450 70.330 122.000 ;
        RECT 70.780 121.450 70.930 129.650 ;
        RECT 71.380 121.450 71.530 129.650 ;
        RECT 71.980 121.450 72.130 129.650 ;
        RECT 72.580 121.450 72.730 129.650 ;
        RECT 73.180 121.450 73.330 129.650 ;
        RECT 73.780 121.450 73.930 129.650 ;
        RECT 74.380 121.450 75.080 138.550 ;
        RECT 75.530 130.350 75.680 138.550 ;
        RECT 76.130 130.350 76.280 138.550 ;
        RECT 76.730 130.350 76.880 138.550 ;
        RECT 77.330 130.350 77.480 138.550 ;
        RECT 77.930 130.350 78.080 138.550 ;
        RECT 78.530 130.350 78.680 138.550 ;
        RECT 79.130 138.000 82.930 138.550 ;
        RECT 86.530 138.550 102.930 138.600 ;
        RECT 86.530 138.000 90.330 138.550 ;
        RECT 79.130 137.550 79.430 138.000 ;
        RECT 90.030 137.550 90.330 138.000 ;
        RECT 79.130 137.400 82.980 137.550 ;
        RECT 86.480 137.400 90.330 137.550 ;
        RECT 79.130 136.950 79.430 137.400 ;
        RECT 90.030 136.950 90.330 137.400 ;
        RECT 79.130 136.800 82.980 136.950 ;
        RECT 86.480 136.800 90.330 136.950 ;
        RECT 79.130 136.350 79.430 136.800 ;
        RECT 90.030 136.350 90.330 136.800 ;
        RECT 79.130 136.200 82.980 136.350 ;
        RECT 86.480 136.200 90.330 136.350 ;
        RECT 79.130 135.750 79.430 136.200 ;
        RECT 90.030 135.750 90.330 136.200 ;
        RECT 79.130 135.600 82.980 135.750 ;
        RECT 86.480 135.600 90.330 135.750 ;
        RECT 79.130 135.150 79.430 135.600 ;
        RECT 90.030 135.150 90.330 135.600 ;
        RECT 79.130 135.000 82.980 135.150 ;
        RECT 86.480 135.000 90.330 135.150 ;
        RECT 79.130 134.550 79.430 135.000 ;
        RECT 90.030 134.550 90.330 135.000 ;
        RECT 79.130 134.400 82.980 134.550 ;
        RECT 86.480 134.400 90.330 134.550 ;
        RECT 79.130 133.950 79.430 134.400 ;
        RECT 90.030 133.950 90.330 134.400 ;
        RECT 79.130 133.800 82.980 133.950 ;
        RECT 86.480 133.800 90.330 133.950 ;
        RECT 79.130 133.350 79.430 133.800 ;
        RECT 90.030 133.350 90.330 133.800 ;
        RECT 79.130 133.200 82.980 133.350 ;
        RECT 86.480 133.200 90.330 133.350 ;
        RECT 79.130 132.750 79.430 133.200 ;
        RECT 79.130 132.600 82.980 132.750 ;
        RECT 79.130 132.150 79.430 132.600 ;
        RECT 79.130 132.000 82.980 132.150 ;
        RECT 79.130 131.550 79.430 132.000 ;
        RECT 79.130 131.400 82.980 131.550 ;
        RECT 79.130 130.950 79.430 131.400 ;
        RECT 79.130 130.800 82.980 130.950 ;
        RECT 79.130 130.350 79.430 130.800 ;
        RECT 75.530 121.450 75.680 129.650 ;
        RECT 76.130 121.450 76.280 129.650 ;
        RECT 76.730 121.450 76.880 129.650 ;
        RECT 77.330 121.450 77.480 129.650 ;
        RECT 77.930 121.450 78.080 129.650 ;
        RECT 78.530 121.450 78.680 129.650 ;
        RECT 79.130 129.200 79.430 129.650 ;
        RECT 79.130 129.050 82.980 129.200 ;
        RECT 79.130 128.600 79.430 129.050 ;
        RECT 79.130 128.450 82.980 128.600 ;
        RECT 79.130 128.000 79.430 128.450 ;
        RECT 79.130 127.850 82.980 128.000 ;
        RECT 79.130 127.400 79.430 127.850 ;
        RECT 79.130 127.250 82.980 127.400 ;
        RECT 79.130 126.800 79.430 127.250 ;
        RECT 83.830 126.800 85.630 133.200 ;
        RECT 90.030 132.750 90.330 133.200 ;
        RECT 86.480 132.600 90.330 132.750 ;
        RECT 90.030 132.150 90.330 132.600 ;
        RECT 86.480 132.000 90.330 132.150 ;
        RECT 90.030 131.550 90.330 132.000 ;
        RECT 86.480 131.400 90.330 131.550 ;
        RECT 90.030 130.950 90.330 131.400 ;
        RECT 86.480 130.800 90.330 130.950 ;
        RECT 90.030 130.350 90.330 130.800 ;
        RECT 90.780 130.350 90.930 138.550 ;
        RECT 91.380 130.350 91.530 138.550 ;
        RECT 91.980 130.350 92.130 138.550 ;
        RECT 92.580 130.350 92.730 138.550 ;
        RECT 93.180 130.350 93.330 138.550 ;
        RECT 93.780 130.350 93.930 138.550 ;
        RECT 90.030 129.200 90.330 129.650 ;
        RECT 86.480 129.050 90.330 129.200 ;
        RECT 90.030 128.600 90.330 129.050 ;
        RECT 86.480 128.450 90.330 128.600 ;
        RECT 90.030 128.000 90.330 128.450 ;
        RECT 86.480 127.850 90.330 128.000 ;
        RECT 90.030 127.400 90.330 127.850 ;
        RECT 86.480 127.250 90.330 127.400 ;
        RECT 90.030 126.800 90.330 127.250 ;
        RECT 79.130 126.650 82.980 126.800 ;
        RECT 86.480 126.650 90.330 126.800 ;
        RECT 79.130 126.200 79.430 126.650 ;
        RECT 90.030 126.200 90.330 126.650 ;
        RECT 79.130 126.050 82.980 126.200 ;
        RECT 86.480 126.050 90.330 126.200 ;
        RECT 79.130 125.600 79.430 126.050 ;
        RECT 90.030 125.600 90.330 126.050 ;
        RECT 79.130 125.450 82.980 125.600 ;
        RECT 86.480 125.450 90.330 125.600 ;
        RECT 79.130 125.000 79.430 125.450 ;
        RECT 90.030 125.000 90.330 125.450 ;
        RECT 79.130 124.850 82.980 125.000 ;
        RECT 86.480 124.850 90.330 125.000 ;
        RECT 79.130 124.400 79.430 124.850 ;
        RECT 90.030 124.400 90.330 124.850 ;
        RECT 79.130 124.250 82.980 124.400 ;
        RECT 86.480 124.250 90.330 124.400 ;
        RECT 79.130 123.800 79.430 124.250 ;
        RECT 90.030 123.800 90.330 124.250 ;
        RECT 79.130 123.650 82.980 123.800 ;
        RECT 86.480 123.650 90.330 123.800 ;
        RECT 79.130 123.200 79.430 123.650 ;
        RECT 90.030 123.200 90.330 123.650 ;
        RECT 79.130 123.050 82.980 123.200 ;
        RECT 86.480 123.050 90.330 123.200 ;
        RECT 79.130 122.600 79.430 123.050 ;
        RECT 90.030 122.600 90.330 123.050 ;
        RECT 79.130 122.450 82.980 122.600 ;
        RECT 86.480 122.450 90.330 122.600 ;
        RECT 79.130 122.000 79.430 122.450 ;
        RECT 90.030 122.000 90.330 122.450 ;
        RECT 79.130 121.450 82.930 122.000 ;
        RECT 66.530 121.400 82.930 121.450 ;
        RECT 86.530 121.450 90.330 122.000 ;
        RECT 90.780 121.450 90.930 129.650 ;
        RECT 91.380 121.450 91.530 129.650 ;
        RECT 91.980 121.450 92.130 129.650 ;
        RECT 92.580 121.450 92.730 129.650 ;
        RECT 93.180 121.450 93.330 129.650 ;
        RECT 93.780 121.450 93.930 129.650 ;
        RECT 94.380 121.450 95.080 138.550 ;
        RECT 95.530 130.350 95.680 138.550 ;
        RECT 96.130 130.350 96.280 138.550 ;
        RECT 96.730 130.350 96.880 138.550 ;
        RECT 97.330 130.350 97.480 138.550 ;
        RECT 97.930 130.350 98.080 138.550 ;
        RECT 98.530 130.350 98.680 138.550 ;
        RECT 99.130 138.000 102.930 138.550 ;
        RECT 99.130 137.550 99.430 138.000 ;
        RECT 99.130 137.400 102.980 137.550 ;
        RECT 99.130 136.950 99.430 137.400 ;
        RECT 99.130 136.800 102.980 136.950 ;
        RECT 99.130 136.350 99.430 136.800 ;
        RECT 99.130 136.200 102.980 136.350 ;
        RECT 99.130 135.750 99.430 136.200 ;
        RECT 99.130 135.600 102.980 135.750 ;
        RECT 99.130 135.150 99.430 135.600 ;
        RECT 99.130 135.000 102.980 135.150 ;
        RECT 99.130 134.550 99.430 135.000 ;
        RECT 99.130 134.400 102.980 134.550 ;
        RECT 99.130 133.950 99.430 134.400 ;
        RECT 99.130 133.800 102.980 133.950 ;
        RECT 99.130 133.350 99.430 133.800 ;
        RECT 99.130 133.200 102.980 133.350 ;
        RECT 99.130 132.750 99.430 133.200 ;
        RECT 99.130 132.600 102.980 132.750 ;
        RECT 99.130 132.150 99.430 132.600 ;
        RECT 99.130 132.000 102.980 132.150 ;
        RECT 99.130 131.550 99.430 132.000 ;
        RECT 99.130 131.400 102.980 131.550 ;
        RECT 99.130 130.950 99.430 131.400 ;
        RECT 99.130 130.800 102.980 130.950 ;
        RECT 99.130 130.350 99.430 130.800 ;
        RECT 95.530 121.450 95.680 129.650 ;
        RECT 96.130 121.450 96.280 129.650 ;
        RECT 96.730 121.450 96.880 129.650 ;
        RECT 97.330 121.450 97.480 129.650 ;
        RECT 97.930 121.450 98.080 129.650 ;
        RECT 98.530 121.450 98.680 129.650 ;
        RECT 99.130 129.200 99.430 129.650 ;
        RECT 99.130 129.050 102.980 129.200 ;
        RECT 99.130 128.600 99.430 129.050 ;
        RECT 99.130 128.450 102.980 128.600 ;
        RECT 99.130 128.000 99.430 128.450 ;
        RECT 99.130 127.850 102.980 128.000 ;
        RECT 99.130 127.400 99.430 127.850 ;
        RECT 99.130 127.250 102.980 127.400 ;
        RECT 99.130 126.800 99.430 127.250 ;
        RECT 103.830 126.800 104.730 133.200 ;
        RECT 109.850 128.705 111.850 129.980 ;
        RECT 99.130 126.650 102.980 126.800 ;
        RECT 99.130 126.200 99.430 126.650 ;
        RECT 99.130 126.050 102.980 126.200 ;
        RECT 99.130 125.600 99.430 126.050 ;
        RECT 99.130 125.450 102.980 125.600 ;
        RECT 99.130 125.000 99.430 125.450 ;
        RECT 99.130 124.850 102.980 125.000 ;
        RECT 99.130 124.400 99.430 124.850 ;
        RECT 99.130 124.250 102.980 124.400 ;
        RECT 99.130 123.800 99.430 124.250 ;
        RECT 99.130 123.650 102.980 123.800 ;
        RECT 99.130 123.200 99.430 123.650 ;
        RECT 99.130 123.050 102.980 123.200 ;
        RECT 99.130 122.600 99.430 123.050 ;
        RECT 99.130 122.450 102.980 122.600 ;
        RECT 99.130 122.000 99.430 122.450 ;
        RECT 99.130 121.450 102.930 122.000 ;
        RECT 86.530 121.400 102.930 121.450 ;
        RECT 9.630 120.900 19.830 121.400 ;
        RECT 29.630 120.900 39.830 121.400 ;
        RECT 49.630 120.900 59.830 121.400 ;
        RECT 69.630 120.900 79.830 121.400 ;
        RECT 89.630 120.900 99.830 121.400 ;
        RECT 11.530 119.100 17.930 120.900 ;
        RECT 31.530 119.100 37.930 120.900 ;
        RECT 51.530 119.100 57.930 120.900 ;
        RECT 71.530 119.100 77.930 120.900 ;
        RECT 91.530 119.100 97.930 120.900 ;
        RECT 9.630 118.600 19.830 119.100 ;
        RECT 29.630 118.600 39.830 119.100 ;
        RECT 49.630 118.600 59.830 119.100 ;
        RECT 69.630 118.600 79.830 119.100 ;
        RECT 89.630 118.600 99.830 119.100 ;
        RECT 6.530 118.550 22.930 118.600 ;
        RECT 6.530 118.000 10.330 118.550 ;
        RECT 10.030 117.550 10.330 118.000 ;
        RECT 6.480 117.400 10.330 117.550 ;
        RECT 10.030 116.950 10.330 117.400 ;
        RECT 6.480 116.800 10.330 116.950 ;
        RECT 10.030 116.350 10.330 116.800 ;
        RECT 6.480 116.200 10.330 116.350 ;
        RECT 10.030 115.750 10.330 116.200 ;
        RECT 6.480 115.600 10.330 115.750 ;
        RECT 10.030 115.150 10.330 115.600 ;
        RECT 6.480 115.000 10.330 115.150 ;
        RECT 10.030 114.550 10.330 115.000 ;
        RECT 6.480 114.400 10.330 114.550 ;
        RECT 10.030 113.950 10.330 114.400 ;
        RECT 6.480 113.800 10.330 113.950 ;
        RECT 10.030 113.350 10.330 113.800 ;
        RECT 6.480 113.200 10.330 113.350 ;
        RECT 4.730 106.800 5.630 113.200 ;
        RECT 10.030 112.750 10.330 113.200 ;
        RECT 6.480 112.600 10.330 112.750 ;
        RECT 10.030 112.150 10.330 112.600 ;
        RECT 6.480 112.000 10.330 112.150 ;
        RECT 10.030 111.550 10.330 112.000 ;
        RECT 6.480 111.400 10.330 111.550 ;
        RECT 10.030 110.950 10.330 111.400 ;
        RECT 6.480 110.800 10.330 110.950 ;
        RECT 10.030 110.350 10.330 110.800 ;
        RECT 10.780 110.350 10.930 118.550 ;
        RECT 11.380 110.350 11.530 118.550 ;
        RECT 11.980 110.350 12.130 118.550 ;
        RECT 12.580 110.350 12.730 118.550 ;
        RECT 13.180 110.350 13.330 118.550 ;
        RECT 13.780 110.350 13.930 118.550 ;
        RECT 10.030 109.200 10.330 109.650 ;
        RECT 6.480 109.050 10.330 109.200 ;
        RECT 10.030 108.600 10.330 109.050 ;
        RECT 6.480 108.450 10.330 108.600 ;
        RECT 10.030 108.000 10.330 108.450 ;
        RECT 6.480 107.850 10.330 108.000 ;
        RECT 10.030 107.400 10.330 107.850 ;
        RECT 6.480 107.250 10.330 107.400 ;
        RECT 10.030 106.800 10.330 107.250 ;
        RECT 6.480 106.650 10.330 106.800 ;
        RECT 10.030 106.200 10.330 106.650 ;
        RECT 6.480 106.050 10.330 106.200 ;
        RECT 10.030 105.600 10.330 106.050 ;
        RECT 6.480 105.450 10.330 105.600 ;
        RECT 10.030 105.000 10.330 105.450 ;
        RECT 6.480 104.850 10.330 105.000 ;
        RECT 10.030 104.400 10.330 104.850 ;
        RECT 6.480 104.250 10.330 104.400 ;
        RECT 10.030 103.800 10.330 104.250 ;
        RECT 6.480 103.650 10.330 103.800 ;
        RECT 10.030 103.200 10.330 103.650 ;
        RECT 6.480 103.050 10.330 103.200 ;
        RECT 10.030 102.600 10.330 103.050 ;
        RECT 6.480 102.450 10.330 102.600 ;
        RECT 10.030 102.000 10.330 102.450 ;
        RECT 6.530 101.450 10.330 102.000 ;
        RECT 10.780 101.450 10.930 109.650 ;
        RECT 11.380 101.450 11.530 109.650 ;
        RECT 11.980 101.450 12.130 109.650 ;
        RECT 12.580 101.450 12.730 109.650 ;
        RECT 13.180 101.450 13.330 109.650 ;
        RECT 13.780 101.450 13.930 109.650 ;
        RECT 14.380 101.450 15.080 118.550 ;
        RECT 15.530 110.350 15.680 118.550 ;
        RECT 16.130 110.350 16.280 118.550 ;
        RECT 16.730 110.350 16.880 118.550 ;
        RECT 17.330 110.350 17.480 118.550 ;
        RECT 17.930 110.350 18.080 118.550 ;
        RECT 18.530 110.350 18.680 118.550 ;
        RECT 19.130 118.000 22.930 118.550 ;
        RECT 26.530 118.550 42.930 118.600 ;
        RECT 26.530 118.000 30.330 118.550 ;
        RECT 19.130 117.550 19.430 118.000 ;
        RECT 30.030 117.550 30.330 118.000 ;
        RECT 19.130 117.400 22.980 117.550 ;
        RECT 26.480 117.400 30.330 117.550 ;
        RECT 19.130 116.950 19.430 117.400 ;
        RECT 30.030 116.950 30.330 117.400 ;
        RECT 19.130 116.800 22.980 116.950 ;
        RECT 26.480 116.800 30.330 116.950 ;
        RECT 19.130 116.350 19.430 116.800 ;
        RECT 30.030 116.350 30.330 116.800 ;
        RECT 19.130 116.200 22.980 116.350 ;
        RECT 26.480 116.200 30.330 116.350 ;
        RECT 19.130 115.750 19.430 116.200 ;
        RECT 30.030 115.750 30.330 116.200 ;
        RECT 19.130 115.600 22.980 115.750 ;
        RECT 26.480 115.600 30.330 115.750 ;
        RECT 19.130 115.150 19.430 115.600 ;
        RECT 30.030 115.150 30.330 115.600 ;
        RECT 19.130 115.000 22.980 115.150 ;
        RECT 26.480 115.000 30.330 115.150 ;
        RECT 19.130 114.550 19.430 115.000 ;
        RECT 30.030 114.550 30.330 115.000 ;
        RECT 19.130 114.400 22.980 114.550 ;
        RECT 26.480 114.400 30.330 114.550 ;
        RECT 19.130 113.950 19.430 114.400 ;
        RECT 30.030 113.950 30.330 114.400 ;
        RECT 19.130 113.800 22.980 113.950 ;
        RECT 26.480 113.800 30.330 113.950 ;
        RECT 19.130 113.350 19.430 113.800 ;
        RECT 30.030 113.350 30.330 113.800 ;
        RECT 19.130 113.200 22.980 113.350 ;
        RECT 26.480 113.200 30.330 113.350 ;
        RECT 19.130 112.750 19.430 113.200 ;
        RECT 19.130 112.600 22.980 112.750 ;
        RECT 19.130 112.150 19.430 112.600 ;
        RECT 19.130 112.000 22.980 112.150 ;
        RECT 19.130 111.550 19.430 112.000 ;
        RECT 19.130 111.400 22.980 111.550 ;
        RECT 19.130 110.950 19.430 111.400 ;
        RECT 19.130 110.800 22.980 110.950 ;
        RECT 19.130 110.350 19.430 110.800 ;
        RECT 15.530 101.450 15.680 109.650 ;
        RECT 16.130 101.450 16.280 109.650 ;
        RECT 16.730 101.450 16.880 109.650 ;
        RECT 17.330 101.450 17.480 109.650 ;
        RECT 17.930 101.450 18.080 109.650 ;
        RECT 18.530 101.450 18.680 109.650 ;
        RECT 19.130 109.200 19.430 109.650 ;
        RECT 19.130 109.050 22.980 109.200 ;
        RECT 19.130 108.600 19.430 109.050 ;
        RECT 19.130 108.450 22.980 108.600 ;
        RECT 19.130 108.000 19.430 108.450 ;
        RECT 19.130 107.850 22.980 108.000 ;
        RECT 19.130 107.400 19.430 107.850 ;
        RECT 19.130 107.250 22.980 107.400 ;
        RECT 19.130 106.800 19.430 107.250 ;
        RECT 23.830 106.800 25.630 113.200 ;
        RECT 30.030 112.750 30.330 113.200 ;
        RECT 26.480 112.600 30.330 112.750 ;
        RECT 30.030 112.150 30.330 112.600 ;
        RECT 26.480 112.000 30.330 112.150 ;
        RECT 30.030 111.550 30.330 112.000 ;
        RECT 26.480 111.400 30.330 111.550 ;
        RECT 30.030 110.950 30.330 111.400 ;
        RECT 26.480 110.800 30.330 110.950 ;
        RECT 30.030 110.350 30.330 110.800 ;
        RECT 30.780 110.350 30.930 118.550 ;
        RECT 31.380 110.350 31.530 118.550 ;
        RECT 31.980 110.350 32.130 118.550 ;
        RECT 32.580 110.350 32.730 118.550 ;
        RECT 33.180 110.350 33.330 118.550 ;
        RECT 33.780 110.350 33.930 118.550 ;
        RECT 30.030 109.200 30.330 109.650 ;
        RECT 26.480 109.050 30.330 109.200 ;
        RECT 30.030 108.600 30.330 109.050 ;
        RECT 26.480 108.450 30.330 108.600 ;
        RECT 30.030 108.000 30.330 108.450 ;
        RECT 26.480 107.850 30.330 108.000 ;
        RECT 30.030 107.400 30.330 107.850 ;
        RECT 26.480 107.250 30.330 107.400 ;
        RECT 30.030 106.800 30.330 107.250 ;
        RECT 19.130 106.650 22.980 106.800 ;
        RECT 26.480 106.650 30.330 106.800 ;
        RECT 19.130 106.200 19.430 106.650 ;
        RECT 30.030 106.200 30.330 106.650 ;
        RECT 19.130 106.050 22.980 106.200 ;
        RECT 26.480 106.050 30.330 106.200 ;
        RECT 19.130 105.600 19.430 106.050 ;
        RECT 30.030 105.600 30.330 106.050 ;
        RECT 19.130 105.450 22.980 105.600 ;
        RECT 26.480 105.450 30.330 105.600 ;
        RECT 19.130 105.000 19.430 105.450 ;
        RECT 30.030 105.000 30.330 105.450 ;
        RECT 19.130 104.850 22.980 105.000 ;
        RECT 26.480 104.850 30.330 105.000 ;
        RECT 19.130 104.400 19.430 104.850 ;
        RECT 30.030 104.400 30.330 104.850 ;
        RECT 19.130 104.250 22.980 104.400 ;
        RECT 26.480 104.250 30.330 104.400 ;
        RECT 19.130 103.800 19.430 104.250 ;
        RECT 30.030 103.800 30.330 104.250 ;
        RECT 19.130 103.650 22.980 103.800 ;
        RECT 26.480 103.650 30.330 103.800 ;
        RECT 19.130 103.200 19.430 103.650 ;
        RECT 30.030 103.200 30.330 103.650 ;
        RECT 19.130 103.050 22.980 103.200 ;
        RECT 26.480 103.050 30.330 103.200 ;
        RECT 19.130 102.600 19.430 103.050 ;
        RECT 30.030 102.600 30.330 103.050 ;
        RECT 19.130 102.450 22.980 102.600 ;
        RECT 26.480 102.450 30.330 102.600 ;
        RECT 19.130 102.000 19.430 102.450 ;
        RECT 30.030 102.000 30.330 102.450 ;
        RECT 19.130 101.450 22.930 102.000 ;
        RECT 6.530 101.400 22.930 101.450 ;
        RECT 26.530 101.450 30.330 102.000 ;
        RECT 30.780 101.450 30.930 109.650 ;
        RECT 31.380 101.450 31.530 109.650 ;
        RECT 31.980 101.450 32.130 109.650 ;
        RECT 32.580 101.450 32.730 109.650 ;
        RECT 33.180 101.450 33.330 109.650 ;
        RECT 33.780 101.450 33.930 109.650 ;
        RECT 34.380 101.450 35.080 118.550 ;
        RECT 35.530 110.350 35.680 118.550 ;
        RECT 36.130 110.350 36.280 118.550 ;
        RECT 36.730 110.350 36.880 118.550 ;
        RECT 37.330 110.350 37.480 118.550 ;
        RECT 37.930 110.350 38.080 118.550 ;
        RECT 38.530 110.350 38.680 118.550 ;
        RECT 39.130 118.000 42.930 118.550 ;
        RECT 46.530 118.550 62.930 118.600 ;
        RECT 46.530 118.000 50.330 118.550 ;
        RECT 39.130 117.550 39.430 118.000 ;
        RECT 50.030 117.550 50.330 118.000 ;
        RECT 39.130 117.400 42.980 117.550 ;
        RECT 46.480 117.400 50.330 117.550 ;
        RECT 39.130 116.950 39.430 117.400 ;
        RECT 50.030 116.950 50.330 117.400 ;
        RECT 39.130 116.800 42.980 116.950 ;
        RECT 46.480 116.800 50.330 116.950 ;
        RECT 39.130 116.350 39.430 116.800 ;
        RECT 50.030 116.350 50.330 116.800 ;
        RECT 39.130 116.200 42.980 116.350 ;
        RECT 46.480 116.200 50.330 116.350 ;
        RECT 39.130 115.750 39.430 116.200 ;
        RECT 50.030 115.750 50.330 116.200 ;
        RECT 39.130 115.600 42.980 115.750 ;
        RECT 46.480 115.600 50.330 115.750 ;
        RECT 39.130 115.150 39.430 115.600 ;
        RECT 50.030 115.150 50.330 115.600 ;
        RECT 39.130 115.000 42.980 115.150 ;
        RECT 46.480 115.000 50.330 115.150 ;
        RECT 39.130 114.550 39.430 115.000 ;
        RECT 50.030 114.550 50.330 115.000 ;
        RECT 39.130 114.400 42.980 114.550 ;
        RECT 46.480 114.400 50.330 114.550 ;
        RECT 39.130 113.950 39.430 114.400 ;
        RECT 50.030 113.950 50.330 114.400 ;
        RECT 39.130 113.800 42.980 113.950 ;
        RECT 46.480 113.800 50.330 113.950 ;
        RECT 39.130 113.350 39.430 113.800 ;
        RECT 50.030 113.350 50.330 113.800 ;
        RECT 39.130 113.200 42.980 113.350 ;
        RECT 46.480 113.200 50.330 113.350 ;
        RECT 39.130 112.750 39.430 113.200 ;
        RECT 39.130 112.600 42.980 112.750 ;
        RECT 39.130 112.150 39.430 112.600 ;
        RECT 39.130 112.000 42.980 112.150 ;
        RECT 39.130 111.550 39.430 112.000 ;
        RECT 39.130 111.400 42.980 111.550 ;
        RECT 39.130 110.950 39.430 111.400 ;
        RECT 39.130 110.800 42.980 110.950 ;
        RECT 39.130 110.350 39.430 110.800 ;
        RECT 35.530 101.450 35.680 109.650 ;
        RECT 36.130 101.450 36.280 109.650 ;
        RECT 36.730 101.450 36.880 109.650 ;
        RECT 37.330 101.450 37.480 109.650 ;
        RECT 37.930 101.450 38.080 109.650 ;
        RECT 38.530 101.450 38.680 109.650 ;
        RECT 39.130 109.200 39.430 109.650 ;
        RECT 39.130 109.050 42.980 109.200 ;
        RECT 39.130 108.600 39.430 109.050 ;
        RECT 39.130 108.450 42.980 108.600 ;
        RECT 39.130 108.000 39.430 108.450 ;
        RECT 39.130 107.850 42.980 108.000 ;
        RECT 39.130 107.400 39.430 107.850 ;
        RECT 39.130 107.250 42.980 107.400 ;
        RECT 39.130 106.800 39.430 107.250 ;
        RECT 43.830 106.800 45.630 113.200 ;
        RECT 50.030 112.750 50.330 113.200 ;
        RECT 46.480 112.600 50.330 112.750 ;
        RECT 50.030 112.150 50.330 112.600 ;
        RECT 46.480 112.000 50.330 112.150 ;
        RECT 50.030 111.550 50.330 112.000 ;
        RECT 46.480 111.400 50.330 111.550 ;
        RECT 50.030 110.950 50.330 111.400 ;
        RECT 46.480 110.800 50.330 110.950 ;
        RECT 50.030 110.350 50.330 110.800 ;
        RECT 50.780 110.350 50.930 118.550 ;
        RECT 51.380 110.350 51.530 118.550 ;
        RECT 51.980 110.350 52.130 118.550 ;
        RECT 52.580 110.350 52.730 118.550 ;
        RECT 53.180 110.350 53.330 118.550 ;
        RECT 53.780 110.350 53.930 118.550 ;
        RECT 50.030 109.200 50.330 109.650 ;
        RECT 46.480 109.050 50.330 109.200 ;
        RECT 50.030 108.600 50.330 109.050 ;
        RECT 46.480 108.450 50.330 108.600 ;
        RECT 50.030 108.000 50.330 108.450 ;
        RECT 46.480 107.850 50.330 108.000 ;
        RECT 50.030 107.400 50.330 107.850 ;
        RECT 46.480 107.250 50.330 107.400 ;
        RECT 50.030 106.800 50.330 107.250 ;
        RECT 39.130 106.650 42.980 106.800 ;
        RECT 46.480 106.650 50.330 106.800 ;
        RECT 39.130 106.200 39.430 106.650 ;
        RECT 50.030 106.200 50.330 106.650 ;
        RECT 39.130 106.050 42.980 106.200 ;
        RECT 46.480 106.050 50.330 106.200 ;
        RECT 39.130 105.600 39.430 106.050 ;
        RECT 50.030 105.600 50.330 106.050 ;
        RECT 39.130 105.450 42.980 105.600 ;
        RECT 46.480 105.450 50.330 105.600 ;
        RECT 39.130 105.000 39.430 105.450 ;
        RECT 50.030 105.000 50.330 105.450 ;
        RECT 39.130 104.850 42.980 105.000 ;
        RECT 46.480 104.850 50.330 105.000 ;
        RECT 39.130 104.400 39.430 104.850 ;
        RECT 50.030 104.400 50.330 104.850 ;
        RECT 39.130 104.250 42.980 104.400 ;
        RECT 46.480 104.250 50.330 104.400 ;
        RECT 39.130 103.800 39.430 104.250 ;
        RECT 50.030 103.800 50.330 104.250 ;
        RECT 39.130 103.650 42.980 103.800 ;
        RECT 46.480 103.650 50.330 103.800 ;
        RECT 39.130 103.200 39.430 103.650 ;
        RECT 50.030 103.200 50.330 103.650 ;
        RECT 39.130 103.050 42.980 103.200 ;
        RECT 46.480 103.050 50.330 103.200 ;
        RECT 39.130 102.600 39.430 103.050 ;
        RECT 50.030 102.600 50.330 103.050 ;
        RECT 39.130 102.450 42.980 102.600 ;
        RECT 46.480 102.450 50.330 102.600 ;
        RECT 39.130 102.000 39.430 102.450 ;
        RECT 50.030 102.000 50.330 102.450 ;
        RECT 39.130 101.450 42.930 102.000 ;
        RECT 26.530 101.400 42.930 101.450 ;
        RECT 46.530 101.450 50.330 102.000 ;
        RECT 50.780 101.450 50.930 109.650 ;
        RECT 51.380 101.450 51.530 109.650 ;
        RECT 51.980 101.450 52.130 109.650 ;
        RECT 52.580 101.450 52.730 109.650 ;
        RECT 53.180 101.450 53.330 109.650 ;
        RECT 53.780 101.450 53.930 109.650 ;
        RECT 54.380 101.450 55.080 118.550 ;
        RECT 55.530 110.350 55.680 118.550 ;
        RECT 56.130 110.350 56.280 118.550 ;
        RECT 56.730 110.350 56.880 118.550 ;
        RECT 57.330 110.350 57.480 118.550 ;
        RECT 57.930 110.350 58.080 118.550 ;
        RECT 58.530 110.350 58.680 118.550 ;
        RECT 59.130 118.000 62.930 118.550 ;
        RECT 66.530 118.550 82.930 118.600 ;
        RECT 66.530 118.000 70.330 118.550 ;
        RECT 59.130 117.550 59.430 118.000 ;
        RECT 70.030 117.550 70.330 118.000 ;
        RECT 59.130 117.400 62.980 117.550 ;
        RECT 66.480 117.400 70.330 117.550 ;
        RECT 59.130 116.950 59.430 117.400 ;
        RECT 70.030 116.950 70.330 117.400 ;
        RECT 59.130 116.800 62.980 116.950 ;
        RECT 66.480 116.800 70.330 116.950 ;
        RECT 59.130 116.350 59.430 116.800 ;
        RECT 70.030 116.350 70.330 116.800 ;
        RECT 59.130 116.200 62.980 116.350 ;
        RECT 66.480 116.200 70.330 116.350 ;
        RECT 59.130 115.750 59.430 116.200 ;
        RECT 70.030 115.750 70.330 116.200 ;
        RECT 59.130 115.600 62.980 115.750 ;
        RECT 66.480 115.600 70.330 115.750 ;
        RECT 59.130 115.150 59.430 115.600 ;
        RECT 70.030 115.150 70.330 115.600 ;
        RECT 59.130 115.000 62.980 115.150 ;
        RECT 66.480 115.000 70.330 115.150 ;
        RECT 59.130 114.550 59.430 115.000 ;
        RECT 70.030 114.550 70.330 115.000 ;
        RECT 59.130 114.400 62.980 114.550 ;
        RECT 66.480 114.400 70.330 114.550 ;
        RECT 59.130 113.950 59.430 114.400 ;
        RECT 70.030 113.950 70.330 114.400 ;
        RECT 59.130 113.800 62.980 113.950 ;
        RECT 66.480 113.800 70.330 113.950 ;
        RECT 59.130 113.350 59.430 113.800 ;
        RECT 70.030 113.350 70.330 113.800 ;
        RECT 59.130 113.200 62.980 113.350 ;
        RECT 66.480 113.200 70.330 113.350 ;
        RECT 59.130 112.750 59.430 113.200 ;
        RECT 59.130 112.600 62.980 112.750 ;
        RECT 59.130 112.150 59.430 112.600 ;
        RECT 59.130 112.000 62.980 112.150 ;
        RECT 59.130 111.550 59.430 112.000 ;
        RECT 59.130 111.400 62.980 111.550 ;
        RECT 59.130 110.950 59.430 111.400 ;
        RECT 59.130 110.800 62.980 110.950 ;
        RECT 59.130 110.350 59.430 110.800 ;
        RECT 55.530 101.450 55.680 109.650 ;
        RECT 56.130 101.450 56.280 109.650 ;
        RECT 56.730 101.450 56.880 109.650 ;
        RECT 57.330 101.450 57.480 109.650 ;
        RECT 57.930 101.450 58.080 109.650 ;
        RECT 58.530 101.450 58.680 109.650 ;
        RECT 59.130 109.200 59.430 109.650 ;
        RECT 59.130 109.050 62.980 109.200 ;
        RECT 59.130 108.600 59.430 109.050 ;
        RECT 59.130 108.450 62.980 108.600 ;
        RECT 59.130 108.000 59.430 108.450 ;
        RECT 59.130 107.850 62.980 108.000 ;
        RECT 59.130 107.400 59.430 107.850 ;
        RECT 59.130 107.250 62.980 107.400 ;
        RECT 59.130 106.800 59.430 107.250 ;
        RECT 63.830 106.800 65.630 113.200 ;
        RECT 70.030 112.750 70.330 113.200 ;
        RECT 66.480 112.600 70.330 112.750 ;
        RECT 70.030 112.150 70.330 112.600 ;
        RECT 66.480 112.000 70.330 112.150 ;
        RECT 70.030 111.550 70.330 112.000 ;
        RECT 66.480 111.400 70.330 111.550 ;
        RECT 70.030 110.950 70.330 111.400 ;
        RECT 66.480 110.800 70.330 110.950 ;
        RECT 70.030 110.350 70.330 110.800 ;
        RECT 70.780 110.350 70.930 118.550 ;
        RECT 71.380 110.350 71.530 118.550 ;
        RECT 71.980 110.350 72.130 118.550 ;
        RECT 72.580 110.350 72.730 118.550 ;
        RECT 73.180 110.350 73.330 118.550 ;
        RECT 73.780 110.350 73.930 118.550 ;
        RECT 70.030 109.200 70.330 109.650 ;
        RECT 66.480 109.050 70.330 109.200 ;
        RECT 70.030 108.600 70.330 109.050 ;
        RECT 66.480 108.450 70.330 108.600 ;
        RECT 70.030 108.000 70.330 108.450 ;
        RECT 66.480 107.850 70.330 108.000 ;
        RECT 70.030 107.400 70.330 107.850 ;
        RECT 66.480 107.250 70.330 107.400 ;
        RECT 70.030 106.800 70.330 107.250 ;
        RECT 59.130 106.650 62.980 106.800 ;
        RECT 66.480 106.650 70.330 106.800 ;
        RECT 59.130 106.200 59.430 106.650 ;
        RECT 70.030 106.200 70.330 106.650 ;
        RECT 59.130 106.050 62.980 106.200 ;
        RECT 66.480 106.050 70.330 106.200 ;
        RECT 59.130 105.600 59.430 106.050 ;
        RECT 70.030 105.600 70.330 106.050 ;
        RECT 59.130 105.450 62.980 105.600 ;
        RECT 66.480 105.450 70.330 105.600 ;
        RECT 59.130 105.000 59.430 105.450 ;
        RECT 70.030 105.000 70.330 105.450 ;
        RECT 59.130 104.850 62.980 105.000 ;
        RECT 66.480 104.850 70.330 105.000 ;
        RECT 59.130 104.400 59.430 104.850 ;
        RECT 70.030 104.400 70.330 104.850 ;
        RECT 59.130 104.250 62.980 104.400 ;
        RECT 66.480 104.250 70.330 104.400 ;
        RECT 59.130 103.800 59.430 104.250 ;
        RECT 70.030 103.800 70.330 104.250 ;
        RECT 59.130 103.650 62.980 103.800 ;
        RECT 66.480 103.650 70.330 103.800 ;
        RECT 59.130 103.200 59.430 103.650 ;
        RECT 70.030 103.200 70.330 103.650 ;
        RECT 59.130 103.050 62.980 103.200 ;
        RECT 66.480 103.050 70.330 103.200 ;
        RECT 59.130 102.600 59.430 103.050 ;
        RECT 70.030 102.600 70.330 103.050 ;
        RECT 59.130 102.450 62.980 102.600 ;
        RECT 66.480 102.450 70.330 102.600 ;
        RECT 59.130 102.000 59.430 102.450 ;
        RECT 70.030 102.000 70.330 102.450 ;
        RECT 59.130 101.450 62.930 102.000 ;
        RECT 46.530 101.400 62.930 101.450 ;
        RECT 66.530 101.450 70.330 102.000 ;
        RECT 70.780 101.450 70.930 109.650 ;
        RECT 71.380 101.450 71.530 109.650 ;
        RECT 71.980 101.450 72.130 109.650 ;
        RECT 72.580 101.450 72.730 109.650 ;
        RECT 73.180 101.450 73.330 109.650 ;
        RECT 73.780 101.450 73.930 109.650 ;
        RECT 74.380 101.450 75.080 118.550 ;
        RECT 75.530 110.350 75.680 118.550 ;
        RECT 76.130 110.350 76.280 118.550 ;
        RECT 76.730 110.350 76.880 118.550 ;
        RECT 77.330 110.350 77.480 118.550 ;
        RECT 77.930 110.350 78.080 118.550 ;
        RECT 78.530 110.350 78.680 118.550 ;
        RECT 79.130 118.000 82.930 118.550 ;
        RECT 86.530 118.550 102.930 118.600 ;
        RECT 86.530 118.000 90.330 118.550 ;
        RECT 79.130 117.550 79.430 118.000 ;
        RECT 90.030 117.550 90.330 118.000 ;
        RECT 79.130 117.400 82.980 117.550 ;
        RECT 86.480 117.400 90.330 117.550 ;
        RECT 79.130 116.950 79.430 117.400 ;
        RECT 90.030 116.950 90.330 117.400 ;
        RECT 79.130 116.800 82.980 116.950 ;
        RECT 86.480 116.800 90.330 116.950 ;
        RECT 79.130 116.350 79.430 116.800 ;
        RECT 90.030 116.350 90.330 116.800 ;
        RECT 79.130 116.200 82.980 116.350 ;
        RECT 86.480 116.200 90.330 116.350 ;
        RECT 79.130 115.750 79.430 116.200 ;
        RECT 90.030 115.750 90.330 116.200 ;
        RECT 79.130 115.600 82.980 115.750 ;
        RECT 86.480 115.600 90.330 115.750 ;
        RECT 79.130 115.150 79.430 115.600 ;
        RECT 90.030 115.150 90.330 115.600 ;
        RECT 79.130 115.000 82.980 115.150 ;
        RECT 86.480 115.000 90.330 115.150 ;
        RECT 79.130 114.550 79.430 115.000 ;
        RECT 90.030 114.550 90.330 115.000 ;
        RECT 79.130 114.400 82.980 114.550 ;
        RECT 86.480 114.400 90.330 114.550 ;
        RECT 79.130 113.950 79.430 114.400 ;
        RECT 90.030 113.950 90.330 114.400 ;
        RECT 79.130 113.800 82.980 113.950 ;
        RECT 86.480 113.800 90.330 113.950 ;
        RECT 79.130 113.350 79.430 113.800 ;
        RECT 90.030 113.350 90.330 113.800 ;
        RECT 79.130 113.200 82.980 113.350 ;
        RECT 86.480 113.200 90.330 113.350 ;
        RECT 79.130 112.750 79.430 113.200 ;
        RECT 79.130 112.600 82.980 112.750 ;
        RECT 79.130 112.150 79.430 112.600 ;
        RECT 79.130 112.000 82.980 112.150 ;
        RECT 79.130 111.550 79.430 112.000 ;
        RECT 79.130 111.400 82.980 111.550 ;
        RECT 79.130 110.950 79.430 111.400 ;
        RECT 79.130 110.800 82.980 110.950 ;
        RECT 79.130 110.350 79.430 110.800 ;
        RECT 75.530 101.450 75.680 109.650 ;
        RECT 76.130 101.450 76.280 109.650 ;
        RECT 76.730 101.450 76.880 109.650 ;
        RECT 77.330 101.450 77.480 109.650 ;
        RECT 77.930 101.450 78.080 109.650 ;
        RECT 78.530 101.450 78.680 109.650 ;
        RECT 79.130 109.200 79.430 109.650 ;
        RECT 79.130 109.050 82.980 109.200 ;
        RECT 79.130 108.600 79.430 109.050 ;
        RECT 79.130 108.450 82.980 108.600 ;
        RECT 79.130 108.000 79.430 108.450 ;
        RECT 79.130 107.850 82.980 108.000 ;
        RECT 79.130 107.400 79.430 107.850 ;
        RECT 79.130 107.250 82.980 107.400 ;
        RECT 79.130 106.800 79.430 107.250 ;
        RECT 83.830 106.800 85.630 113.200 ;
        RECT 90.030 112.750 90.330 113.200 ;
        RECT 86.480 112.600 90.330 112.750 ;
        RECT 90.030 112.150 90.330 112.600 ;
        RECT 86.480 112.000 90.330 112.150 ;
        RECT 90.030 111.550 90.330 112.000 ;
        RECT 86.480 111.400 90.330 111.550 ;
        RECT 90.030 110.950 90.330 111.400 ;
        RECT 86.480 110.800 90.330 110.950 ;
        RECT 90.030 110.350 90.330 110.800 ;
        RECT 90.780 110.350 90.930 118.550 ;
        RECT 91.380 110.350 91.530 118.550 ;
        RECT 91.980 110.350 92.130 118.550 ;
        RECT 92.580 110.350 92.730 118.550 ;
        RECT 93.180 110.350 93.330 118.550 ;
        RECT 93.780 110.350 93.930 118.550 ;
        RECT 90.030 109.200 90.330 109.650 ;
        RECT 86.480 109.050 90.330 109.200 ;
        RECT 90.030 108.600 90.330 109.050 ;
        RECT 86.480 108.450 90.330 108.600 ;
        RECT 90.030 108.000 90.330 108.450 ;
        RECT 86.480 107.850 90.330 108.000 ;
        RECT 90.030 107.400 90.330 107.850 ;
        RECT 86.480 107.250 90.330 107.400 ;
        RECT 90.030 106.800 90.330 107.250 ;
        RECT 79.130 106.650 82.980 106.800 ;
        RECT 86.480 106.650 90.330 106.800 ;
        RECT 79.130 106.200 79.430 106.650 ;
        RECT 90.030 106.200 90.330 106.650 ;
        RECT 79.130 106.050 82.980 106.200 ;
        RECT 86.480 106.050 90.330 106.200 ;
        RECT 79.130 105.600 79.430 106.050 ;
        RECT 90.030 105.600 90.330 106.050 ;
        RECT 79.130 105.450 82.980 105.600 ;
        RECT 86.480 105.450 90.330 105.600 ;
        RECT 79.130 105.000 79.430 105.450 ;
        RECT 90.030 105.000 90.330 105.450 ;
        RECT 79.130 104.850 82.980 105.000 ;
        RECT 86.480 104.850 90.330 105.000 ;
        RECT 79.130 104.400 79.430 104.850 ;
        RECT 90.030 104.400 90.330 104.850 ;
        RECT 79.130 104.250 82.980 104.400 ;
        RECT 86.480 104.250 90.330 104.400 ;
        RECT 79.130 103.800 79.430 104.250 ;
        RECT 90.030 103.800 90.330 104.250 ;
        RECT 79.130 103.650 82.980 103.800 ;
        RECT 86.480 103.650 90.330 103.800 ;
        RECT 79.130 103.200 79.430 103.650 ;
        RECT 90.030 103.200 90.330 103.650 ;
        RECT 79.130 103.050 82.980 103.200 ;
        RECT 86.480 103.050 90.330 103.200 ;
        RECT 79.130 102.600 79.430 103.050 ;
        RECT 90.030 102.600 90.330 103.050 ;
        RECT 79.130 102.450 82.980 102.600 ;
        RECT 86.480 102.450 90.330 102.600 ;
        RECT 79.130 102.000 79.430 102.450 ;
        RECT 90.030 102.000 90.330 102.450 ;
        RECT 79.130 101.450 82.930 102.000 ;
        RECT 66.530 101.400 82.930 101.450 ;
        RECT 86.530 101.450 90.330 102.000 ;
        RECT 90.780 101.450 90.930 109.650 ;
        RECT 91.380 101.450 91.530 109.650 ;
        RECT 91.980 101.450 92.130 109.650 ;
        RECT 92.580 101.450 92.730 109.650 ;
        RECT 93.180 101.450 93.330 109.650 ;
        RECT 93.780 101.450 93.930 109.650 ;
        RECT 94.380 101.450 95.080 118.550 ;
        RECT 95.530 110.350 95.680 118.550 ;
        RECT 96.130 110.350 96.280 118.550 ;
        RECT 96.730 110.350 96.880 118.550 ;
        RECT 97.330 110.350 97.480 118.550 ;
        RECT 97.930 110.350 98.080 118.550 ;
        RECT 98.530 110.350 98.680 118.550 ;
        RECT 99.130 118.000 102.930 118.550 ;
        RECT 99.130 117.550 99.430 118.000 ;
        RECT 99.130 117.400 102.980 117.550 ;
        RECT 99.130 116.950 99.430 117.400 ;
        RECT 99.130 116.800 102.980 116.950 ;
        RECT 99.130 116.350 99.430 116.800 ;
        RECT 99.130 116.200 102.980 116.350 ;
        RECT 99.130 115.750 99.430 116.200 ;
        RECT 99.130 115.600 102.980 115.750 ;
        RECT 99.130 115.150 99.430 115.600 ;
        RECT 99.130 115.000 102.980 115.150 ;
        RECT 99.130 114.550 99.430 115.000 ;
        RECT 99.130 114.400 102.980 114.550 ;
        RECT 99.130 113.950 99.430 114.400 ;
        RECT 99.130 113.800 102.980 113.950 ;
        RECT 99.130 113.350 99.430 113.800 ;
        RECT 99.130 113.200 102.980 113.350 ;
        RECT 99.130 112.750 99.430 113.200 ;
        RECT 99.130 112.600 102.980 112.750 ;
        RECT 99.130 112.150 99.430 112.600 ;
        RECT 99.130 112.000 102.980 112.150 ;
        RECT 99.130 111.550 99.430 112.000 ;
        RECT 99.130 111.400 102.980 111.550 ;
        RECT 99.130 110.950 99.430 111.400 ;
        RECT 99.130 110.800 102.980 110.950 ;
        RECT 99.130 110.350 99.430 110.800 ;
        RECT 95.530 101.450 95.680 109.650 ;
        RECT 96.130 101.450 96.280 109.650 ;
        RECT 96.730 101.450 96.880 109.650 ;
        RECT 97.330 101.450 97.480 109.650 ;
        RECT 97.930 101.450 98.080 109.650 ;
        RECT 98.530 101.450 98.680 109.650 ;
        RECT 99.130 109.200 99.430 109.650 ;
        RECT 99.130 109.050 102.980 109.200 ;
        RECT 99.130 108.600 99.430 109.050 ;
        RECT 99.130 108.450 102.980 108.600 ;
        RECT 99.130 108.000 99.430 108.450 ;
        RECT 99.130 107.850 102.980 108.000 ;
        RECT 99.130 107.400 99.430 107.850 ;
        RECT 99.130 107.250 102.980 107.400 ;
        RECT 99.130 106.800 99.430 107.250 ;
        RECT 103.830 106.800 104.730 113.200 ;
        RECT 109.850 109.755 111.850 111.030 ;
        RECT 99.130 106.650 102.980 106.800 ;
        RECT 99.130 106.200 99.430 106.650 ;
        RECT 99.130 106.050 102.980 106.200 ;
        RECT 99.130 105.600 99.430 106.050 ;
        RECT 99.130 105.450 102.980 105.600 ;
        RECT 99.130 105.000 99.430 105.450 ;
        RECT 99.130 104.850 102.980 105.000 ;
        RECT 99.130 104.400 99.430 104.850 ;
        RECT 99.130 104.250 102.980 104.400 ;
        RECT 99.130 103.800 99.430 104.250 ;
        RECT 99.130 103.650 102.980 103.800 ;
        RECT 99.130 103.200 99.430 103.650 ;
        RECT 99.130 103.050 102.980 103.200 ;
        RECT 99.130 102.600 99.430 103.050 ;
        RECT 99.130 102.450 102.980 102.600 ;
        RECT 99.130 102.000 99.430 102.450 ;
        RECT 99.130 101.450 102.930 102.000 ;
        RECT 86.530 101.400 102.930 101.450 ;
        RECT 9.630 100.900 19.830 101.400 ;
        RECT 29.630 100.900 39.830 101.400 ;
        RECT 49.630 100.900 59.830 101.400 ;
        RECT 69.630 100.900 79.830 101.400 ;
        RECT 89.630 100.900 99.830 101.400 ;
        RECT 11.530 99.100 17.930 100.900 ;
        RECT 31.530 99.100 37.930 100.900 ;
        RECT 51.530 99.100 57.930 100.900 ;
        RECT 71.530 99.100 77.930 100.900 ;
        RECT 91.530 99.100 97.930 100.900 ;
        RECT 9.630 98.600 19.830 99.100 ;
        RECT 29.630 98.600 39.830 99.100 ;
        RECT 49.630 98.600 59.830 99.100 ;
        RECT 69.630 98.600 79.830 99.100 ;
        RECT 89.630 98.600 99.830 99.100 ;
        RECT 6.530 98.550 22.930 98.600 ;
        RECT 6.530 98.000 10.330 98.550 ;
        RECT 10.030 97.550 10.330 98.000 ;
        RECT 6.480 97.400 10.330 97.550 ;
        RECT 10.030 96.950 10.330 97.400 ;
        RECT 6.480 96.800 10.330 96.950 ;
        RECT 10.030 96.350 10.330 96.800 ;
        RECT 6.480 96.200 10.330 96.350 ;
        RECT 10.030 95.750 10.330 96.200 ;
        RECT 6.480 95.600 10.330 95.750 ;
        RECT 10.030 95.150 10.330 95.600 ;
        RECT 6.480 95.000 10.330 95.150 ;
        RECT 10.030 94.550 10.330 95.000 ;
        RECT 6.480 94.400 10.330 94.550 ;
        RECT 10.030 93.950 10.330 94.400 ;
        RECT 6.480 93.800 10.330 93.950 ;
        RECT 10.030 93.350 10.330 93.800 ;
        RECT 6.480 93.200 10.330 93.350 ;
        RECT 4.730 86.800 5.630 93.200 ;
        RECT 10.030 92.750 10.330 93.200 ;
        RECT 6.480 92.600 10.330 92.750 ;
        RECT 10.030 92.150 10.330 92.600 ;
        RECT 6.480 92.000 10.330 92.150 ;
        RECT 10.030 91.550 10.330 92.000 ;
        RECT 6.480 91.400 10.330 91.550 ;
        RECT 10.030 90.950 10.330 91.400 ;
        RECT 6.480 90.800 10.330 90.950 ;
        RECT 10.030 90.350 10.330 90.800 ;
        RECT 10.780 90.350 10.930 98.550 ;
        RECT 11.380 90.350 11.530 98.550 ;
        RECT 11.980 90.350 12.130 98.550 ;
        RECT 12.580 90.350 12.730 98.550 ;
        RECT 13.180 90.350 13.330 98.550 ;
        RECT 13.780 90.350 13.930 98.550 ;
        RECT 10.030 89.200 10.330 89.650 ;
        RECT 6.480 89.050 10.330 89.200 ;
        RECT 10.030 88.600 10.330 89.050 ;
        RECT 6.480 88.450 10.330 88.600 ;
        RECT 10.030 88.000 10.330 88.450 ;
        RECT 6.480 87.850 10.330 88.000 ;
        RECT 10.030 87.400 10.330 87.850 ;
        RECT 6.480 87.250 10.330 87.400 ;
        RECT 10.030 86.800 10.330 87.250 ;
        RECT 6.480 86.650 10.330 86.800 ;
        RECT 10.030 86.200 10.330 86.650 ;
        RECT 6.480 86.050 10.330 86.200 ;
        RECT 10.030 85.600 10.330 86.050 ;
        RECT 6.480 85.450 10.330 85.600 ;
        RECT 10.030 85.000 10.330 85.450 ;
        RECT 6.480 84.850 10.330 85.000 ;
        RECT 10.030 84.400 10.330 84.850 ;
        RECT 6.480 84.250 10.330 84.400 ;
        RECT 10.030 83.800 10.330 84.250 ;
        RECT 6.480 83.650 10.330 83.800 ;
        RECT 10.030 83.200 10.330 83.650 ;
        RECT 6.480 83.050 10.330 83.200 ;
        RECT 10.030 82.600 10.330 83.050 ;
        RECT 6.480 82.450 10.330 82.600 ;
        RECT 10.030 82.000 10.330 82.450 ;
        RECT 6.530 81.450 10.330 82.000 ;
        RECT 10.780 81.450 10.930 89.650 ;
        RECT 11.380 81.450 11.530 89.650 ;
        RECT 11.980 81.450 12.130 89.650 ;
        RECT 12.580 81.450 12.730 89.650 ;
        RECT 13.180 81.450 13.330 89.650 ;
        RECT 13.780 81.450 13.930 89.650 ;
        RECT 14.380 81.450 15.080 98.550 ;
        RECT 15.530 90.350 15.680 98.550 ;
        RECT 16.130 90.350 16.280 98.550 ;
        RECT 16.730 90.350 16.880 98.550 ;
        RECT 17.330 90.350 17.480 98.550 ;
        RECT 17.930 90.350 18.080 98.550 ;
        RECT 18.530 90.350 18.680 98.550 ;
        RECT 19.130 98.000 22.930 98.550 ;
        RECT 26.530 98.550 42.930 98.600 ;
        RECT 26.530 98.000 30.330 98.550 ;
        RECT 19.130 97.550 19.430 98.000 ;
        RECT 30.030 97.550 30.330 98.000 ;
        RECT 19.130 97.400 22.980 97.550 ;
        RECT 26.480 97.400 30.330 97.550 ;
        RECT 19.130 96.950 19.430 97.400 ;
        RECT 30.030 96.950 30.330 97.400 ;
        RECT 19.130 96.800 22.980 96.950 ;
        RECT 26.480 96.800 30.330 96.950 ;
        RECT 19.130 96.350 19.430 96.800 ;
        RECT 30.030 96.350 30.330 96.800 ;
        RECT 19.130 96.200 22.980 96.350 ;
        RECT 26.480 96.200 30.330 96.350 ;
        RECT 19.130 95.750 19.430 96.200 ;
        RECT 30.030 95.750 30.330 96.200 ;
        RECT 19.130 95.600 22.980 95.750 ;
        RECT 26.480 95.600 30.330 95.750 ;
        RECT 19.130 95.150 19.430 95.600 ;
        RECT 30.030 95.150 30.330 95.600 ;
        RECT 19.130 95.000 22.980 95.150 ;
        RECT 26.480 95.000 30.330 95.150 ;
        RECT 19.130 94.550 19.430 95.000 ;
        RECT 30.030 94.550 30.330 95.000 ;
        RECT 19.130 94.400 22.980 94.550 ;
        RECT 26.480 94.400 30.330 94.550 ;
        RECT 19.130 93.950 19.430 94.400 ;
        RECT 30.030 93.950 30.330 94.400 ;
        RECT 19.130 93.800 22.980 93.950 ;
        RECT 26.480 93.800 30.330 93.950 ;
        RECT 19.130 93.350 19.430 93.800 ;
        RECT 30.030 93.350 30.330 93.800 ;
        RECT 19.130 93.200 22.980 93.350 ;
        RECT 26.480 93.200 30.330 93.350 ;
        RECT 19.130 92.750 19.430 93.200 ;
        RECT 19.130 92.600 22.980 92.750 ;
        RECT 19.130 92.150 19.430 92.600 ;
        RECT 19.130 92.000 22.980 92.150 ;
        RECT 19.130 91.550 19.430 92.000 ;
        RECT 19.130 91.400 22.980 91.550 ;
        RECT 19.130 90.950 19.430 91.400 ;
        RECT 19.130 90.800 22.980 90.950 ;
        RECT 19.130 90.350 19.430 90.800 ;
        RECT 15.530 81.450 15.680 89.650 ;
        RECT 16.130 81.450 16.280 89.650 ;
        RECT 16.730 81.450 16.880 89.650 ;
        RECT 17.330 81.450 17.480 89.650 ;
        RECT 17.930 81.450 18.080 89.650 ;
        RECT 18.530 81.450 18.680 89.650 ;
        RECT 19.130 89.200 19.430 89.650 ;
        RECT 19.130 89.050 22.980 89.200 ;
        RECT 19.130 88.600 19.430 89.050 ;
        RECT 19.130 88.450 22.980 88.600 ;
        RECT 19.130 88.000 19.430 88.450 ;
        RECT 19.130 87.850 22.980 88.000 ;
        RECT 19.130 87.400 19.430 87.850 ;
        RECT 19.130 87.250 22.980 87.400 ;
        RECT 19.130 86.800 19.430 87.250 ;
        RECT 23.830 86.800 25.630 93.200 ;
        RECT 30.030 92.750 30.330 93.200 ;
        RECT 26.480 92.600 30.330 92.750 ;
        RECT 30.030 92.150 30.330 92.600 ;
        RECT 26.480 92.000 30.330 92.150 ;
        RECT 30.030 91.550 30.330 92.000 ;
        RECT 26.480 91.400 30.330 91.550 ;
        RECT 30.030 90.950 30.330 91.400 ;
        RECT 26.480 90.800 30.330 90.950 ;
        RECT 30.030 90.350 30.330 90.800 ;
        RECT 30.780 90.350 30.930 98.550 ;
        RECT 31.380 90.350 31.530 98.550 ;
        RECT 31.980 90.350 32.130 98.550 ;
        RECT 32.580 90.350 32.730 98.550 ;
        RECT 33.180 90.350 33.330 98.550 ;
        RECT 33.780 90.350 33.930 98.550 ;
        RECT 30.030 89.200 30.330 89.650 ;
        RECT 26.480 89.050 30.330 89.200 ;
        RECT 30.030 88.600 30.330 89.050 ;
        RECT 26.480 88.450 30.330 88.600 ;
        RECT 30.030 88.000 30.330 88.450 ;
        RECT 26.480 87.850 30.330 88.000 ;
        RECT 30.030 87.400 30.330 87.850 ;
        RECT 26.480 87.250 30.330 87.400 ;
        RECT 30.030 86.800 30.330 87.250 ;
        RECT 19.130 86.650 22.980 86.800 ;
        RECT 26.480 86.650 30.330 86.800 ;
        RECT 19.130 86.200 19.430 86.650 ;
        RECT 30.030 86.200 30.330 86.650 ;
        RECT 19.130 86.050 22.980 86.200 ;
        RECT 26.480 86.050 30.330 86.200 ;
        RECT 19.130 85.600 19.430 86.050 ;
        RECT 30.030 85.600 30.330 86.050 ;
        RECT 19.130 85.450 22.980 85.600 ;
        RECT 26.480 85.450 30.330 85.600 ;
        RECT 19.130 85.000 19.430 85.450 ;
        RECT 30.030 85.000 30.330 85.450 ;
        RECT 19.130 84.850 22.980 85.000 ;
        RECT 26.480 84.850 30.330 85.000 ;
        RECT 19.130 84.400 19.430 84.850 ;
        RECT 30.030 84.400 30.330 84.850 ;
        RECT 19.130 84.250 22.980 84.400 ;
        RECT 26.480 84.250 30.330 84.400 ;
        RECT 19.130 83.800 19.430 84.250 ;
        RECT 30.030 83.800 30.330 84.250 ;
        RECT 19.130 83.650 22.980 83.800 ;
        RECT 26.480 83.650 30.330 83.800 ;
        RECT 19.130 83.200 19.430 83.650 ;
        RECT 30.030 83.200 30.330 83.650 ;
        RECT 19.130 83.050 22.980 83.200 ;
        RECT 26.480 83.050 30.330 83.200 ;
        RECT 19.130 82.600 19.430 83.050 ;
        RECT 30.030 82.600 30.330 83.050 ;
        RECT 19.130 82.450 22.980 82.600 ;
        RECT 26.480 82.450 30.330 82.600 ;
        RECT 19.130 82.000 19.430 82.450 ;
        RECT 30.030 82.000 30.330 82.450 ;
        RECT 19.130 81.450 22.930 82.000 ;
        RECT 6.530 81.400 22.930 81.450 ;
        RECT 26.530 81.450 30.330 82.000 ;
        RECT 30.780 81.450 30.930 89.650 ;
        RECT 31.380 81.450 31.530 89.650 ;
        RECT 31.980 81.450 32.130 89.650 ;
        RECT 32.580 81.450 32.730 89.650 ;
        RECT 33.180 81.450 33.330 89.650 ;
        RECT 33.780 81.450 33.930 89.650 ;
        RECT 34.380 81.450 35.080 98.550 ;
        RECT 35.530 90.350 35.680 98.550 ;
        RECT 36.130 90.350 36.280 98.550 ;
        RECT 36.730 90.350 36.880 98.550 ;
        RECT 37.330 90.350 37.480 98.550 ;
        RECT 37.930 90.350 38.080 98.550 ;
        RECT 38.530 90.350 38.680 98.550 ;
        RECT 39.130 98.000 42.930 98.550 ;
        RECT 46.530 98.550 62.930 98.600 ;
        RECT 46.530 98.000 50.330 98.550 ;
        RECT 39.130 97.550 39.430 98.000 ;
        RECT 50.030 97.550 50.330 98.000 ;
        RECT 39.130 97.400 42.980 97.550 ;
        RECT 46.480 97.400 50.330 97.550 ;
        RECT 39.130 96.950 39.430 97.400 ;
        RECT 50.030 96.950 50.330 97.400 ;
        RECT 39.130 96.800 42.980 96.950 ;
        RECT 46.480 96.800 50.330 96.950 ;
        RECT 39.130 96.350 39.430 96.800 ;
        RECT 50.030 96.350 50.330 96.800 ;
        RECT 39.130 96.200 42.980 96.350 ;
        RECT 46.480 96.200 50.330 96.350 ;
        RECT 39.130 95.750 39.430 96.200 ;
        RECT 50.030 95.750 50.330 96.200 ;
        RECT 39.130 95.600 42.980 95.750 ;
        RECT 46.480 95.600 50.330 95.750 ;
        RECT 39.130 95.150 39.430 95.600 ;
        RECT 50.030 95.150 50.330 95.600 ;
        RECT 39.130 95.000 42.980 95.150 ;
        RECT 46.480 95.000 50.330 95.150 ;
        RECT 39.130 94.550 39.430 95.000 ;
        RECT 50.030 94.550 50.330 95.000 ;
        RECT 39.130 94.400 42.980 94.550 ;
        RECT 46.480 94.400 50.330 94.550 ;
        RECT 39.130 93.950 39.430 94.400 ;
        RECT 50.030 93.950 50.330 94.400 ;
        RECT 39.130 93.800 42.980 93.950 ;
        RECT 46.480 93.800 50.330 93.950 ;
        RECT 39.130 93.350 39.430 93.800 ;
        RECT 50.030 93.350 50.330 93.800 ;
        RECT 39.130 93.200 42.980 93.350 ;
        RECT 46.480 93.200 50.330 93.350 ;
        RECT 39.130 92.750 39.430 93.200 ;
        RECT 39.130 92.600 42.980 92.750 ;
        RECT 39.130 92.150 39.430 92.600 ;
        RECT 39.130 92.000 42.980 92.150 ;
        RECT 39.130 91.550 39.430 92.000 ;
        RECT 39.130 91.400 42.980 91.550 ;
        RECT 39.130 90.950 39.430 91.400 ;
        RECT 39.130 90.800 42.980 90.950 ;
        RECT 39.130 90.350 39.430 90.800 ;
        RECT 35.530 81.450 35.680 89.650 ;
        RECT 36.130 81.450 36.280 89.650 ;
        RECT 36.730 81.450 36.880 89.650 ;
        RECT 37.330 81.450 37.480 89.650 ;
        RECT 37.930 81.450 38.080 89.650 ;
        RECT 38.530 81.450 38.680 89.650 ;
        RECT 39.130 89.200 39.430 89.650 ;
        RECT 39.130 89.050 42.980 89.200 ;
        RECT 39.130 88.600 39.430 89.050 ;
        RECT 39.130 88.450 42.980 88.600 ;
        RECT 39.130 88.000 39.430 88.450 ;
        RECT 39.130 87.850 42.980 88.000 ;
        RECT 39.130 87.400 39.430 87.850 ;
        RECT 39.130 87.250 42.980 87.400 ;
        RECT 39.130 86.800 39.430 87.250 ;
        RECT 43.830 86.800 45.630 93.200 ;
        RECT 50.030 92.750 50.330 93.200 ;
        RECT 46.480 92.600 50.330 92.750 ;
        RECT 50.030 92.150 50.330 92.600 ;
        RECT 46.480 92.000 50.330 92.150 ;
        RECT 50.030 91.550 50.330 92.000 ;
        RECT 46.480 91.400 50.330 91.550 ;
        RECT 50.030 90.950 50.330 91.400 ;
        RECT 46.480 90.800 50.330 90.950 ;
        RECT 50.030 90.350 50.330 90.800 ;
        RECT 50.780 90.350 50.930 98.550 ;
        RECT 51.380 90.350 51.530 98.550 ;
        RECT 51.980 90.350 52.130 98.550 ;
        RECT 52.580 90.350 52.730 98.550 ;
        RECT 53.180 90.350 53.330 98.550 ;
        RECT 53.780 90.350 53.930 98.550 ;
        RECT 50.030 89.200 50.330 89.650 ;
        RECT 46.480 89.050 50.330 89.200 ;
        RECT 50.030 88.600 50.330 89.050 ;
        RECT 46.480 88.450 50.330 88.600 ;
        RECT 50.030 88.000 50.330 88.450 ;
        RECT 46.480 87.850 50.330 88.000 ;
        RECT 50.030 87.400 50.330 87.850 ;
        RECT 46.480 87.250 50.330 87.400 ;
        RECT 50.030 86.800 50.330 87.250 ;
        RECT 39.130 86.650 42.980 86.800 ;
        RECT 46.480 86.650 50.330 86.800 ;
        RECT 39.130 86.200 39.430 86.650 ;
        RECT 50.030 86.200 50.330 86.650 ;
        RECT 39.130 86.050 42.980 86.200 ;
        RECT 46.480 86.050 50.330 86.200 ;
        RECT 39.130 85.600 39.430 86.050 ;
        RECT 50.030 85.600 50.330 86.050 ;
        RECT 39.130 85.450 42.980 85.600 ;
        RECT 46.480 85.450 50.330 85.600 ;
        RECT 39.130 85.000 39.430 85.450 ;
        RECT 50.030 85.000 50.330 85.450 ;
        RECT 39.130 84.850 42.980 85.000 ;
        RECT 46.480 84.850 50.330 85.000 ;
        RECT 39.130 84.400 39.430 84.850 ;
        RECT 50.030 84.400 50.330 84.850 ;
        RECT 39.130 84.250 42.980 84.400 ;
        RECT 46.480 84.250 50.330 84.400 ;
        RECT 39.130 83.800 39.430 84.250 ;
        RECT 50.030 83.800 50.330 84.250 ;
        RECT 39.130 83.650 42.980 83.800 ;
        RECT 46.480 83.650 50.330 83.800 ;
        RECT 39.130 83.200 39.430 83.650 ;
        RECT 50.030 83.200 50.330 83.650 ;
        RECT 39.130 83.050 42.980 83.200 ;
        RECT 46.480 83.050 50.330 83.200 ;
        RECT 39.130 82.600 39.430 83.050 ;
        RECT 50.030 82.600 50.330 83.050 ;
        RECT 39.130 82.450 42.980 82.600 ;
        RECT 46.480 82.450 50.330 82.600 ;
        RECT 39.130 82.000 39.430 82.450 ;
        RECT 50.030 82.000 50.330 82.450 ;
        RECT 39.130 81.450 42.930 82.000 ;
        RECT 26.530 81.400 42.930 81.450 ;
        RECT 46.530 81.450 50.330 82.000 ;
        RECT 50.780 81.450 50.930 89.650 ;
        RECT 51.380 81.450 51.530 89.650 ;
        RECT 51.980 81.450 52.130 89.650 ;
        RECT 52.580 81.450 52.730 89.650 ;
        RECT 53.180 81.450 53.330 89.650 ;
        RECT 53.780 81.450 53.930 89.650 ;
        RECT 54.380 81.450 55.080 98.550 ;
        RECT 55.530 90.350 55.680 98.550 ;
        RECT 56.130 90.350 56.280 98.550 ;
        RECT 56.730 90.350 56.880 98.550 ;
        RECT 57.330 90.350 57.480 98.550 ;
        RECT 57.930 90.350 58.080 98.550 ;
        RECT 58.530 90.350 58.680 98.550 ;
        RECT 59.130 98.000 62.930 98.550 ;
        RECT 66.530 98.550 82.930 98.600 ;
        RECT 66.530 98.000 70.330 98.550 ;
        RECT 59.130 97.550 59.430 98.000 ;
        RECT 70.030 97.550 70.330 98.000 ;
        RECT 59.130 97.400 62.980 97.550 ;
        RECT 66.480 97.400 70.330 97.550 ;
        RECT 59.130 96.950 59.430 97.400 ;
        RECT 70.030 96.950 70.330 97.400 ;
        RECT 59.130 96.800 62.980 96.950 ;
        RECT 66.480 96.800 70.330 96.950 ;
        RECT 59.130 96.350 59.430 96.800 ;
        RECT 70.030 96.350 70.330 96.800 ;
        RECT 59.130 96.200 62.980 96.350 ;
        RECT 66.480 96.200 70.330 96.350 ;
        RECT 59.130 95.750 59.430 96.200 ;
        RECT 70.030 95.750 70.330 96.200 ;
        RECT 59.130 95.600 62.980 95.750 ;
        RECT 66.480 95.600 70.330 95.750 ;
        RECT 59.130 95.150 59.430 95.600 ;
        RECT 70.030 95.150 70.330 95.600 ;
        RECT 59.130 95.000 62.980 95.150 ;
        RECT 66.480 95.000 70.330 95.150 ;
        RECT 59.130 94.550 59.430 95.000 ;
        RECT 70.030 94.550 70.330 95.000 ;
        RECT 59.130 94.400 62.980 94.550 ;
        RECT 66.480 94.400 70.330 94.550 ;
        RECT 59.130 93.950 59.430 94.400 ;
        RECT 70.030 93.950 70.330 94.400 ;
        RECT 59.130 93.800 62.980 93.950 ;
        RECT 66.480 93.800 70.330 93.950 ;
        RECT 59.130 93.350 59.430 93.800 ;
        RECT 70.030 93.350 70.330 93.800 ;
        RECT 59.130 93.200 62.980 93.350 ;
        RECT 66.480 93.200 70.330 93.350 ;
        RECT 59.130 92.750 59.430 93.200 ;
        RECT 59.130 92.600 62.980 92.750 ;
        RECT 59.130 92.150 59.430 92.600 ;
        RECT 59.130 92.000 62.980 92.150 ;
        RECT 59.130 91.550 59.430 92.000 ;
        RECT 59.130 91.400 62.980 91.550 ;
        RECT 59.130 90.950 59.430 91.400 ;
        RECT 59.130 90.800 62.980 90.950 ;
        RECT 59.130 90.350 59.430 90.800 ;
        RECT 55.530 81.450 55.680 89.650 ;
        RECT 56.130 81.450 56.280 89.650 ;
        RECT 56.730 81.450 56.880 89.650 ;
        RECT 57.330 81.450 57.480 89.650 ;
        RECT 57.930 81.450 58.080 89.650 ;
        RECT 58.530 81.450 58.680 89.650 ;
        RECT 59.130 89.200 59.430 89.650 ;
        RECT 59.130 89.050 62.980 89.200 ;
        RECT 59.130 88.600 59.430 89.050 ;
        RECT 59.130 88.450 62.980 88.600 ;
        RECT 59.130 88.000 59.430 88.450 ;
        RECT 59.130 87.850 62.980 88.000 ;
        RECT 59.130 87.400 59.430 87.850 ;
        RECT 59.130 87.250 62.980 87.400 ;
        RECT 59.130 86.800 59.430 87.250 ;
        RECT 63.830 86.800 65.630 93.200 ;
        RECT 70.030 92.750 70.330 93.200 ;
        RECT 66.480 92.600 70.330 92.750 ;
        RECT 70.030 92.150 70.330 92.600 ;
        RECT 66.480 92.000 70.330 92.150 ;
        RECT 70.030 91.550 70.330 92.000 ;
        RECT 66.480 91.400 70.330 91.550 ;
        RECT 70.030 90.950 70.330 91.400 ;
        RECT 66.480 90.800 70.330 90.950 ;
        RECT 70.030 90.350 70.330 90.800 ;
        RECT 70.780 90.350 70.930 98.550 ;
        RECT 71.380 90.350 71.530 98.550 ;
        RECT 71.980 90.350 72.130 98.550 ;
        RECT 72.580 90.350 72.730 98.550 ;
        RECT 73.180 90.350 73.330 98.550 ;
        RECT 73.780 90.350 73.930 98.550 ;
        RECT 70.030 89.200 70.330 89.650 ;
        RECT 66.480 89.050 70.330 89.200 ;
        RECT 70.030 88.600 70.330 89.050 ;
        RECT 66.480 88.450 70.330 88.600 ;
        RECT 70.030 88.000 70.330 88.450 ;
        RECT 66.480 87.850 70.330 88.000 ;
        RECT 70.030 87.400 70.330 87.850 ;
        RECT 66.480 87.250 70.330 87.400 ;
        RECT 70.030 86.800 70.330 87.250 ;
        RECT 59.130 86.650 62.980 86.800 ;
        RECT 66.480 86.650 70.330 86.800 ;
        RECT 59.130 86.200 59.430 86.650 ;
        RECT 70.030 86.200 70.330 86.650 ;
        RECT 59.130 86.050 62.980 86.200 ;
        RECT 66.480 86.050 70.330 86.200 ;
        RECT 59.130 85.600 59.430 86.050 ;
        RECT 70.030 85.600 70.330 86.050 ;
        RECT 59.130 85.450 62.980 85.600 ;
        RECT 66.480 85.450 70.330 85.600 ;
        RECT 59.130 85.000 59.430 85.450 ;
        RECT 70.030 85.000 70.330 85.450 ;
        RECT 59.130 84.850 62.980 85.000 ;
        RECT 66.480 84.850 70.330 85.000 ;
        RECT 59.130 84.400 59.430 84.850 ;
        RECT 70.030 84.400 70.330 84.850 ;
        RECT 59.130 84.250 62.980 84.400 ;
        RECT 66.480 84.250 70.330 84.400 ;
        RECT 59.130 83.800 59.430 84.250 ;
        RECT 70.030 83.800 70.330 84.250 ;
        RECT 59.130 83.650 62.980 83.800 ;
        RECT 66.480 83.650 70.330 83.800 ;
        RECT 59.130 83.200 59.430 83.650 ;
        RECT 70.030 83.200 70.330 83.650 ;
        RECT 59.130 83.050 62.980 83.200 ;
        RECT 66.480 83.050 70.330 83.200 ;
        RECT 59.130 82.600 59.430 83.050 ;
        RECT 70.030 82.600 70.330 83.050 ;
        RECT 59.130 82.450 62.980 82.600 ;
        RECT 66.480 82.450 70.330 82.600 ;
        RECT 59.130 82.000 59.430 82.450 ;
        RECT 70.030 82.000 70.330 82.450 ;
        RECT 59.130 81.450 62.930 82.000 ;
        RECT 46.530 81.400 62.930 81.450 ;
        RECT 66.530 81.450 70.330 82.000 ;
        RECT 70.780 81.450 70.930 89.650 ;
        RECT 71.380 81.450 71.530 89.650 ;
        RECT 71.980 81.450 72.130 89.650 ;
        RECT 72.580 81.450 72.730 89.650 ;
        RECT 73.180 81.450 73.330 89.650 ;
        RECT 73.780 81.450 73.930 89.650 ;
        RECT 74.380 81.450 75.080 98.550 ;
        RECT 75.530 90.350 75.680 98.550 ;
        RECT 76.130 90.350 76.280 98.550 ;
        RECT 76.730 90.350 76.880 98.550 ;
        RECT 77.330 90.350 77.480 98.550 ;
        RECT 77.930 90.350 78.080 98.550 ;
        RECT 78.530 90.350 78.680 98.550 ;
        RECT 79.130 98.000 82.930 98.550 ;
        RECT 86.530 98.550 102.930 98.600 ;
        RECT 86.530 98.000 90.330 98.550 ;
        RECT 79.130 97.550 79.430 98.000 ;
        RECT 90.030 97.550 90.330 98.000 ;
        RECT 79.130 97.400 82.980 97.550 ;
        RECT 86.480 97.400 90.330 97.550 ;
        RECT 79.130 96.950 79.430 97.400 ;
        RECT 90.030 96.950 90.330 97.400 ;
        RECT 79.130 96.800 82.980 96.950 ;
        RECT 86.480 96.800 90.330 96.950 ;
        RECT 79.130 96.350 79.430 96.800 ;
        RECT 90.030 96.350 90.330 96.800 ;
        RECT 79.130 96.200 82.980 96.350 ;
        RECT 86.480 96.200 90.330 96.350 ;
        RECT 79.130 95.750 79.430 96.200 ;
        RECT 90.030 95.750 90.330 96.200 ;
        RECT 79.130 95.600 82.980 95.750 ;
        RECT 86.480 95.600 90.330 95.750 ;
        RECT 79.130 95.150 79.430 95.600 ;
        RECT 90.030 95.150 90.330 95.600 ;
        RECT 79.130 95.000 82.980 95.150 ;
        RECT 86.480 95.000 90.330 95.150 ;
        RECT 79.130 94.550 79.430 95.000 ;
        RECT 90.030 94.550 90.330 95.000 ;
        RECT 79.130 94.400 82.980 94.550 ;
        RECT 86.480 94.400 90.330 94.550 ;
        RECT 79.130 93.950 79.430 94.400 ;
        RECT 90.030 93.950 90.330 94.400 ;
        RECT 79.130 93.800 82.980 93.950 ;
        RECT 86.480 93.800 90.330 93.950 ;
        RECT 79.130 93.350 79.430 93.800 ;
        RECT 90.030 93.350 90.330 93.800 ;
        RECT 79.130 93.200 82.980 93.350 ;
        RECT 86.480 93.200 90.330 93.350 ;
        RECT 79.130 92.750 79.430 93.200 ;
        RECT 79.130 92.600 82.980 92.750 ;
        RECT 79.130 92.150 79.430 92.600 ;
        RECT 79.130 92.000 82.980 92.150 ;
        RECT 79.130 91.550 79.430 92.000 ;
        RECT 79.130 91.400 82.980 91.550 ;
        RECT 79.130 90.950 79.430 91.400 ;
        RECT 79.130 90.800 82.980 90.950 ;
        RECT 79.130 90.350 79.430 90.800 ;
        RECT 75.530 81.450 75.680 89.650 ;
        RECT 76.130 81.450 76.280 89.650 ;
        RECT 76.730 81.450 76.880 89.650 ;
        RECT 77.330 81.450 77.480 89.650 ;
        RECT 77.930 81.450 78.080 89.650 ;
        RECT 78.530 81.450 78.680 89.650 ;
        RECT 79.130 89.200 79.430 89.650 ;
        RECT 79.130 89.050 82.980 89.200 ;
        RECT 79.130 88.600 79.430 89.050 ;
        RECT 79.130 88.450 82.980 88.600 ;
        RECT 79.130 88.000 79.430 88.450 ;
        RECT 79.130 87.850 82.980 88.000 ;
        RECT 79.130 87.400 79.430 87.850 ;
        RECT 79.130 87.250 82.980 87.400 ;
        RECT 79.130 86.800 79.430 87.250 ;
        RECT 83.830 86.800 85.630 93.200 ;
        RECT 90.030 92.750 90.330 93.200 ;
        RECT 86.480 92.600 90.330 92.750 ;
        RECT 90.030 92.150 90.330 92.600 ;
        RECT 86.480 92.000 90.330 92.150 ;
        RECT 90.030 91.550 90.330 92.000 ;
        RECT 86.480 91.400 90.330 91.550 ;
        RECT 90.030 90.950 90.330 91.400 ;
        RECT 86.480 90.800 90.330 90.950 ;
        RECT 90.030 90.350 90.330 90.800 ;
        RECT 90.780 90.350 90.930 98.550 ;
        RECT 91.380 90.350 91.530 98.550 ;
        RECT 91.980 90.350 92.130 98.550 ;
        RECT 92.580 90.350 92.730 98.550 ;
        RECT 93.180 90.350 93.330 98.550 ;
        RECT 93.780 90.350 93.930 98.550 ;
        RECT 90.030 89.200 90.330 89.650 ;
        RECT 86.480 89.050 90.330 89.200 ;
        RECT 90.030 88.600 90.330 89.050 ;
        RECT 86.480 88.450 90.330 88.600 ;
        RECT 90.030 88.000 90.330 88.450 ;
        RECT 86.480 87.850 90.330 88.000 ;
        RECT 90.030 87.400 90.330 87.850 ;
        RECT 86.480 87.250 90.330 87.400 ;
        RECT 90.030 86.800 90.330 87.250 ;
        RECT 79.130 86.650 82.980 86.800 ;
        RECT 86.480 86.650 90.330 86.800 ;
        RECT 79.130 86.200 79.430 86.650 ;
        RECT 90.030 86.200 90.330 86.650 ;
        RECT 79.130 86.050 82.980 86.200 ;
        RECT 86.480 86.050 90.330 86.200 ;
        RECT 79.130 85.600 79.430 86.050 ;
        RECT 90.030 85.600 90.330 86.050 ;
        RECT 79.130 85.450 82.980 85.600 ;
        RECT 86.480 85.450 90.330 85.600 ;
        RECT 79.130 85.000 79.430 85.450 ;
        RECT 90.030 85.000 90.330 85.450 ;
        RECT 79.130 84.850 82.980 85.000 ;
        RECT 86.480 84.850 90.330 85.000 ;
        RECT 79.130 84.400 79.430 84.850 ;
        RECT 90.030 84.400 90.330 84.850 ;
        RECT 79.130 84.250 82.980 84.400 ;
        RECT 86.480 84.250 90.330 84.400 ;
        RECT 79.130 83.800 79.430 84.250 ;
        RECT 90.030 83.800 90.330 84.250 ;
        RECT 79.130 83.650 82.980 83.800 ;
        RECT 86.480 83.650 90.330 83.800 ;
        RECT 79.130 83.200 79.430 83.650 ;
        RECT 90.030 83.200 90.330 83.650 ;
        RECT 79.130 83.050 82.980 83.200 ;
        RECT 86.480 83.050 90.330 83.200 ;
        RECT 79.130 82.600 79.430 83.050 ;
        RECT 90.030 82.600 90.330 83.050 ;
        RECT 79.130 82.450 82.980 82.600 ;
        RECT 86.480 82.450 90.330 82.600 ;
        RECT 79.130 82.000 79.430 82.450 ;
        RECT 90.030 82.000 90.330 82.450 ;
        RECT 79.130 81.450 82.930 82.000 ;
        RECT 66.530 81.400 82.930 81.450 ;
        RECT 86.530 81.450 90.330 82.000 ;
        RECT 90.780 81.450 90.930 89.650 ;
        RECT 91.380 81.450 91.530 89.650 ;
        RECT 91.980 81.450 92.130 89.650 ;
        RECT 92.580 81.450 92.730 89.650 ;
        RECT 93.180 81.450 93.330 89.650 ;
        RECT 93.780 81.450 93.930 89.650 ;
        RECT 94.380 81.450 95.080 98.550 ;
        RECT 95.530 90.350 95.680 98.550 ;
        RECT 96.130 90.350 96.280 98.550 ;
        RECT 96.730 90.350 96.880 98.550 ;
        RECT 97.330 90.350 97.480 98.550 ;
        RECT 97.930 90.350 98.080 98.550 ;
        RECT 98.530 90.350 98.680 98.550 ;
        RECT 99.130 98.000 102.930 98.550 ;
        RECT 99.130 97.550 99.430 98.000 ;
        RECT 99.130 97.400 102.980 97.550 ;
        RECT 99.130 96.950 99.430 97.400 ;
        RECT 99.130 96.800 102.980 96.950 ;
        RECT 99.130 96.350 99.430 96.800 ;
        RECT 99.130 96.200 102.980 96.350 ;
        RECT 99.130 95.750 99.430 96.200 ;
        RECT 99.130 95.600 102.980 95.750 ;
        RECT 99.130 95.150 99.430 95.600 ;
        RECT 99.130 95.000 102.980 95.150 ;
        RECT 99.130 94.550 99.430 95.000 ;
        RECT 99.130 94.400 102.980 94.550 ;
        RECT 99.130 93.950 99.430 94.400 ;
        RECT 99.130 93.800 102.980 93.950 ;
        RECT 99.130 93.350 99.430 93.800 ;
        RECT 99.130 93.200 102.980 93.350 ;
        RECT 99.130 92.750 99.430 93.200 ;
        RECT 99.130 92.600 102.980 92.750 ;
        RECT 99.130 92.150 99.430 92.600 ;
        RECT 99.130 92.000 102.980 92.150 ;
        RECT 99.130 91.550 99.430 92.000 ;
        RECT 99.130 91.400 102.980 91.550 ;
        RECT 99.130 90.950 99.430 91.400 ;
        RECT 99.130 90.800 102.980 90.950 ;
        RECT 99.130 90.350 99.430 90.800 ;
        RECT 95.530 81.450 95.680 89.650 ;
        RECT 96.130 81.450 96.280 89.650 ;
        RECT 96.730 81.450 96.880 89.650 ;
        RECT 97.330 81.450 97.480 89.650 ;
        RECT 97.930 81.450 98.080 89.650 ;
        RECT 98.530 81.450 98.680 89.650 ;
        RECT 99.130 89.200 99.430 89.650 ;
        RECT 99.130 89.050 102.980 89.200 ;
        RECT 99.130 88.600 99.430 89.050 ;
        RECT 99.130 88.450 102.980 88.600 ;
        RECT 99.130 88.000 99.430 88.450 ;
        RECT 99.130 87.850 102.980 88.000 ;
        RECT 99.130 87.400 99.430 87.850 ;
        RECT 99.130 87.250 102.980 87.400 ;
        RECT 99.130 86.800 99.430 87.250 ;
        RECT 103.830 86.800 104.730 93.200 ;
        RECT 109.850 89.220 111.850 90.495 ;
        RECT 99.130 86.650 102.980 86.800 ;
        RECT 99.130 86.200 99.430 86.650 ;
        RECT 99.130 86.050 102.980 86.200 ;
        RECT 99.130 85.600 99.430 86.050 ;
        RECT 99.130 85.450 102.980 85.600 ;
        RECT 99.130 85.000 99.430 85.450 ;
        RECT 99.130 84.850 102.980 85.000 ;
        RECT 99.130 84.400 99.430 84.850 ;
        RECT 99.130 84.250 102.980 84.400 ;
        RECT 99.130 83.800 99.430 84.250 ;
        RECT 99.130 83.650 102.980 83.800 ;
        RECT 99.130 83.200 99.430 83.650 ;
        RECT 99.130 83.050 102.980 83.200 ;
        RECT 99.130 82.600 99.430 83.050 ;
        RECT 99.130 82.450 102.980 82.600 ;
        RECT 99.130 82.000 99.430 82.450 ;
        RECT 99.130 81.450 102.930 82.000 ;
        RECT 86.530 81.400 102.930 81.450 ;
        RECT 9.630 80.900 19.830 81.400 ;
        RECT 29.630 80.900 39.830 81.400 ;
        RECT 49.630 80.900 59.830 81.400 ;
        RECT 69.630 80.900 79.830 81.400 ;
        RECT 89.630 80.900 99.830 81.400 ;
        RECT 11.530 79.100 17.930 80.900 ;
        RECT 31.530 79.100 37.930 80.900 ;
        RECT 51.530 79.100 57.930 80.900 ;
        RECT 71.530 79.100 77.930 80.900 ;
        RECT 91.530 79.100 97.930 80.900 ;
        RECT 9.630 78.600 19.830 79.100 ;
        RECT 29.630 78.600 39.830 79.100 ;
        RECT 49.630 78.600 59.830 79.100 ;
        RECT 69.630 78.600 79.830 79.100 ;
        RECT 89.630 78.600 99.830 79.100 ;
        RECT 6.530 78.550 22.930 78.600 ;
        RECT 6.530 78.000 10.330 78.550 ;
        RECT 10.030 77.550 10.330 78.000 ;
        RECT 6.480 77.400 10.330 77.550 ;
        RECT 10.030 76.950 10.330 77.400 ;
        RECT 6.480 76.800 10.330 76.950 ;
        RECT 10.030 76.350 10.330 76.800 ;
        RECT 6.480 76.200 10.330 76.350 ;
        RECT 10.030 75.750 10.330 76.200 ;
        RECT 6.480 75.600 10.330 75.750 ;
        RECT 10.030 75.150 10.330 75.600 ;
        RECT 6.480 75.000 10.330 75.150 ;
        RECT 10.030 74.550 10.330 75.000 ;
        RECT 6.480 74.400 10.330 74.550 ;
        RECT 10.030 73.950 10.330 74.400 ;
        RECT 6.480 73.800 10.330 73.950 ;
        RECT 10.030 73.350 10.330 73.800 ;
        RECT 6.480 73.200 10.330 73.350 ;
        RECT 4.730 66.800 5.630 73.200 ;
        RECT 10.030 72.750 10.330 73.200 ;
        RECT 6.480 72.600 10.330 72.750 ;
        RECT 10.030 72.150 10.330 72.600 ;
        RECT 6.480 72.000 10.330 72.150 ;
        RECT 10.030 71.550 10.330 72.000 ;
        RECT 6.480 71.400 10.330 71.550 ;
        RECT 10.030 70.950 10.330 71.400 ;
        RECT 6.480 70.800 10.330 70.950 ;
        RECT 10.030 70.350 10.330 70.800 ;
        RECT 10.780 70.350 10.930 78.550 ;
        RECT 11.380 70.350 11.530 78.550 ;
        RECT 11.980 70.350 12.130 78.550 ;
        RECT 12.580 70.350 12.730 78.550 ;
        RECT 13.180 70.350 13.330 78.550 ;
        RECT 13.780 70.350 13.930 78.550 ;
        RECT 10.030 69.200 10.330 69.650 ;
        RECT 6.480 69.050 10.330 69.200 ;
        RECT 10.030 68.600 10.330 69.050 ;
        RECT 6.480 68.450 10.330 68.600 ;
        RECT 10.030 68.000 10.330 68.450 ;
        RECT 6.480 67.850 10.330 68.000 ;
        RECT 10.030 67.400 10.330 67.850 ;
        RECT 6.480 67.250 10.330 67.400 ;
        RECT 10.030 66.800 10.330 67.250 ;
        RECT 6.480 66.650 10.330 66.800 ;
        RECT 10.030 66.200 10.330 66.650 ;
        RECT 6.480 66.050 10.330 66.200 ;
        RECT 10.030 65.600 10.330 66.050 ;
        RECT 6.480 65.450 10.330 65.600 ;
        RECT 10.030 65.000 10.330 65.450 ;
        RECT 6.480 64.850 10.330 65.000 ;
        RECT 10.030 64.400 10.330 64.850 ;
        RECT 6.480 64.250 10.330 64.400 ;
        RECT 10.030 63.800 10.330 64.250 ;
        RECT 6.480 63.650 10.330 63.800 ;
        RECT 10.030 63.200 10.330 63.650 ;
        RECT 6.480 63.050 10.330 63.200 ;
        RECT 10.030 62.600 10.330 63.050 ;
        RECT 6.480 62.450 10.330 62.600 ;
        RECT 10.030 62.000 10.330 62.450 ;
        RECT 6.530 61.450 10.330 62.000 ;
        RECT 10.780 61.450 10.930 69.650 ;
        RECT 11.380 61.450 11.530 69.650 ;
        RECT 11.980 61.450 12.130 69.650 ;
        RECT 12.580 61.450 12.730 69.650 ;
        RECT 13.180 61.450 13.330 69.650 ;
        RECT 13.780 61.450 13.930 69.650 ;
        RECT 14.380 61.450 15.080 78.550 ;
        RECT 15.530 70.350 15.680 78.550 ;
        RECT 16.130 70.350 16.280 78.550 ;
        RECT 16.730 70.350 16.880 78.550 ;
        RECT 17.330 70.350 17.480 78.550 ;
        RECT 17.930 70.350 18.080 78.550 ;
        RECT 18.530 70.350 18.680 78.550 ;
        RECT 19.130 78.000 22.930 78.550 ;
        RECT 26.530 78.550 42.930 78.600 ;
        RECT 26.530 78.000 30.330 78.550 ;
        RECT 19.130 77.550 19.430 78.000 ;
        RECT 30.030 77.550 30.330 78.000 ;
        RECT 19.130 77.400 22.980 77.550 ;
        RECT 26.480 77.400 30.330 77.550 ;
        RECT 19.130 76.950 19.430 77.400 ;
        RECT 30.030 76.950 30.330 77.400 ;
        RECT 19.130 76.800 22.980 76.950 ;
        RECT 26.480 76.800 30.330 76.950 ;
        RECT 19.130 76.350 19.430 76.800 ;
        RECT 30.030 76.350 30.330 76.800 ;
        RECT 19.130 76.200 22.980 76.350 ;
        RECT 26.480 76.200 30.330 76.350 ;
        RECT 19.130 75.750 19.430 76.200 ;
        RECT 30.030 75.750 30.330 76.200 ;
        RECT 19.130 75.600 22.980 75.750 ;
        RECT 26.480 75.600 30.330 75.750 ;
        RECT 19.130 75.150 19.430 75.600 ;
        RECT 30.030 75.150 30.330 75.600 ;
        RECT 19.130 75.000 22.980 75.150 ;
        RECT 26.480 75.000 30.330 75.150 ;
        RECT 19.130 74.550 19.430 75.000 ;
        RECT 30.030 74.550 30.330 75.000 ;
        RECT 19.130 74.400 22.980 74.550 ;
        RECT 26.480 74.400 30.330 74.550 ;
        RECT 19.130 73.950 19.430 74.400 ;
        RECT 30.030 73.950 30.330 74.400 ;
        RECT 19.130 73.800 22.980 73.950 ;
        RECT 26.480 73.800 30.330 73.950 ;
        RECT 19.130 73.350 19.430 73.800 ;
        RECT 30.030 73.350 30.330 73.800 ;
        RECT 19.130 73.200 22.980 73.350 ;
        RECT 26.480 73.200 30.330 73.350 ;
        RECT 19.130 72.750 19.430 73.200 ;
        RECT 19.130 72.600 22.980 72.750 ;
        RECT 19.130 72.150 19.430 72.600 ;
        RECT 19.130 72.000 22.980 72.150 ;
        RECT 19.130 71.550 19.430 72.000 ;
        RECT 19.130 71.400 22.980 71.550 ;
        RECT 19.130 70.950 19.430 71.400 ;
        RECT 19.130 70.800 22.980 70.950 ;
        RECT 19.130 70.350 19.430 70.800 ;
        RECT 15.530 61.450 15.680 69.650 ;
        RECT 16.130 61.450 16.280 69.650 ;
        RECT 16.730 61.450 16.880 69.650 ;
        RECT 17.330 61.450 17.480 69.650 ;
        RECT 17.930 61.450 18.080 69.650 ;
        RECT 18.530 61.450 18.680 69.650 ;
        RECT 19.130 69.200 19.430 69.650 ;
        RECT 19.130 69.050 22.980 69.200 ;
        RECT 19.130 68.600 19.430 69.050 ;
        RECT 19.130 68.450 22.980 68.600 ;
        RECT 19.130 68.000 19.430 68.450 ;
        RECT 19.130 67.850 22.980 68.000 ;
        RECT 19.130 67.400 19.430 67.850 ;
        RECT 19.130 67.250 22.980 67.400 ;
        RECT 19.130 66.800 19.430 67.250 ;
        RECT 23.830 66.800 25.630 73.200 ;
        RECT 30.030 72.750 30.330 73.200 ;
        RECT 26.480 72.600 30.330 72.750 ;
        RECT 30.030 72.150 30.330 72.600 ;
        RECT 26.480 72.000 30.330 72.150 ;
        RECT 30.030 71.550 30.330 72.000 ;
        RECT 26.480 71.400 30.330 71.550 ;
        RECT 30.030 70.950 30.330 71.400 ;
        RECT 26.480 70.800 30.330 70.950 ;
        RECT 30.030 70.350 30.330 70.800 ;
        RECT 30.780 70.350 30.930 78.550 ;
        RECT 31.380 70.350 31.530 78.550 ;
        RECT 31.980 70.350 32.130 78.550 ;
        RECT 32.580 70.350 32.730 78.550 ;
        RECT 33.180 70.350 33.330 78.550 ;
        RECT 33.780 70.350 33.930 78.550 ;
        RECT 30.030 69.200 30.330 69.650 ;
        RECT 26.480 69.050 30.330 69.200 ;
        RECT 30.030 68.600 30.330 69.050 ;
        RECT 26.480 68.450 30.330 68.600 ;
        RECT 30.030 68.000 30.330 68.450 ;
        RECT 26.480 67.850 30.330 68.000 ;
        RECT 30.030 67.400 30.330 67.850 ;
        RECT 26.480 67.250 30.330 67.400 ;
        RECT 30.030 66.800 30.330 67.250 ;
        RECT 19.130 66.650 22.980 66.800 ;
        RECT 26.480 66.650 30.330 66.800 ;
        RECT 19.130 66.200 19.430 66.650 ;
        RECT 30.030 66.200 30.330 66.650 ;
        RECT 19.130 66.050 22.980 66.200 ;
        RECT 26.480 66.050 30.330 66.200 ;
        RECT 19.130 65.600 19.430 66.050 ;
        RECT 30.030 65.600 30.330 66.050 ;
        RECT 19.130 65.450 22.980 65.600 ;
        RECT 26.480 65.450 30.330 65.600 ;
        RECT 19.130 65.000 19.430 65.450 ;
        RECT 30.030 65.000 30.330 65.450 ;
        RECT 19.130 64.850 22.980 65.000 ;
        RECT 26.480 64.850 30.330 65.000 ;
        RECT 19.130 64.400 19.430 64.850 ;
        RECT 30.030 64.400 30.330 64.850 ;
        RECT 19.130 64.250 22.980 64.400 ;
        RECT 26.480 64.250 30.330 64.400 ;
        RECT 19.130 63.800 19.430 64.250 ;
        RECT 30.030 63.800 30.330 64.250 ;
        RECT 19.130 63.650 22.980 63.800 ;
        RECT 26.480 63.650 30.330 63.800 ;
        RECT 19.130 63.200 19.430 63.650 ;
        RECT 30.030 63.200 30.330 63.650 ;
        RECT 19.130 63.050 22.980 63.200 ;
        RECT 26.480 63.050 30.330 63.200 ;
        RECT 19.130 62.600 19.430 63.050 ;
        RECT 30.030 62.600 30.330 63.050 ;
        RECT 19.130 62.450 22.980 62.600 ;
        RECT 26.480 62.450 30.330 62.600 ;
        RECT 19.130 62.000 19.430 62.450 ;
        RECT 30.030 62.000 30.330 62.450 ;
        RECT 19.130 61.450 22.930 62.000 ;
        RECT 6.530 61.400 22.930 61.450 ;
        RECT 26.530 61.450 30.330 62.000 ;
        RECT 30.780 61.450 30.930 69.650 ;
        RECT 31.380 61.450 31.530 69.650 ;
        RECT 31.980 61.450 32.130 69.650 ;
        RECT 32.580 61.450 32.730 69.650 ;
        RECT 33.180 61.450 33.330 69.650 ;
        RECT 33.780 61.450 33.930 69.650 ;
        RECT 34.380 61.450 35.080 78.550 ;
        RECT 35.530 70.350 35.680 78.550 ;
        RECT 36.130 70.350 36.280 78.550 ;
        RECT 36.730 70.350 36.880 78.550 ;
        RECT 37.330 70.350 37.480 78.550 ;
        RECT 37.930 70.350 38.080 78.550 ;
        RECT 38.530 70.350 38.680 78.550 ;
        RECT 39.130 78.000 42.930 78.550 ;
        RECT 46.530 78.550 62.930 78.600 ;
        RECT 46.530 78.000 50.330 78.550 ;
        RECT 39.130 77.550 39.430 78.000 ;
        RECT 50.030 77.550 50.330 78.000 ;
        RECT 39.130 77.400 42.980 77.550 ;
        RECT 46.480 77.400 50.330 77.550 ;
        RECT 39.130 76.950 39.430 77.400 ;
        RECT 50.030 76.950 50.330 77.400 ;
        RECT 39.130 76.800 42.980 76.950 ;
        RECT 46.480 76.800 50.330 76.950 ;
        RECT 39.130 76.350 39.430 76.800 ;
        RECT 50.030 76.350 50.330 76.800 ;
        RECT 39.130 76.200 42.980 76.350 ;
        RECT 46.480 76.200 50.330 76.350 ;
        RECT 39.130 75.750 39.430 76.200 ;
        RECT 50.030 75.750 50.330 76.200 ;
        RECT 39.130 75.600 42.980 75.750 ;
        RECT 46.480 75.600 50.330 75.750 ;
        RECT 39.130 75.150 39.430 75.600 ;
        RECT 50.030 75.150 50.330 75.600 ;
        RECT 39.130 75.000 42.980 75.150 ;
        RECT 46.480 75.000 50.330 75.150 ;
        RECT 39.130 74.550 39.430 75.000 ;
        RECT 50.030 74.550 50.330 75.000 ;
        RECT 39.130 74.400 42.980 74.550 ;
        RECT 46.480 74.400 50.330 74.550 ;
        RECT 39.130 73.950 39.430 74.400 ;
        RECT 50.030 73.950 50.330 74.400 ;
        RECT 39.130 73.800 42.980 73.950 ;
        RECT 46.480 73.800 50.330 73.950 ;
        RECT 39.130 73.350 39.430 73.800 ;
        RECT 50.030 73.350 50.330 73.800 ;
        RECT 39.130 73.200 42.980 73.350 ;
        RECT 46.480 73.200 50.330 73.350 ;
        RECT 39.130 72.750 39.430 73.200 ;
        RECT 39.130 72.600 42.980 72.750 ;
        RECT 39.130 72.150 39.430 72.600 ;
        RECT 39.130 72.000 42.980 72.150 ;
        RECT 39.130 71.550 39.430 72.000 ;
        RECT 39.130 71.400 42.980 71.550 ;
        RECT 39.130 70.950 39.430 71.400 ;
        RECT 39.130 70.800 42.980 70.950 ;
        RECT 39.130 70.350 39.430 70.800 ;
        RECT 35.530 61.450 35.680 69.650 ;
        RECT 36.130 61.450 36.280 69.650 ;
        RECT 36.730 61.450 36.880 69.650 ;
        RECT 37.330 61.450 37.480 69.650 ;
        RECT 37.930 61.450 38.080 69.650 ;
        RECT 38.530 61.450 38.680 69.650 ;
        RECT 39.130 69.200 39.430 69.650 ;
        RECT 39.130 69.050 42.980 69.200 ;
        RECT 39.130 68.600 39.430 69.050 ;
        RECT 39.130 68.450 42.980 68.600 ;
        RECT 39.130 68.000 39.430 68.450 ;
        RECT 39.130 67.850 42.980 68.000 ;
        RECT 39.130 67.400 39.430 67.850 ;
        RECT 39.130 67.250 42.980 67.400 ;
        RECT 39.130 66.800 39.430 67.250 ;
        RECT 43.830 66.800 45.630 73.200 ;
        RECT 50.030 72.750 50.330 73.200 ;
        RECT 46.480 72.600 50.330 72.750 ;
        RECT 50.030 72.150 50.330 72.600 ;
        RECT 46.480 72.000 50.330 72.150 ;
        RECT 50.030 71.550 50.330 72.000 ;
        RECT 46.480 71.400 50.330 71.550 ;
        RECT 50.030 70.950 50.330 71.400 ;
        RECT 46.480 70.800 50.330 70.950 ;
        RECT 50.030 70.350 50.330 70.800 ;
        RECT 50.780 70.350 50.930 78.550 ;
        RECT 51.380 70.350 51.530 78.550 ;
        RECT 51.980 70.350 52.130 78.550 ;
        RECT 52.580 70.350 52.730 78.550 ;
        RECT 53.180 70.350 53.330 78.550 ;
        RECT 53.780 70.350 53.930 78.550 ;
        RECT 50.030 69.200 50.330 69.650 ;
        RECT 46.480 69.050 50.330 69.200 ;
        RECT 50.030 68.600 50.330 69.050 ;
        RECT 46.480 68.450 50.330 68.600 ;
        RECT 50.030 68.000 50.330 68.450 ;
        RECT 46.480 67.850 50.330 68.000 ;
        RECT 50.030 67.400 50.330 67.850 ;
        RECT 46.480 67.250 50.330 67.400 ;
        RECT 50.030 66.800 50.330 67.250 ;
        RECT 39.130 66.650 42.980 66.800 ;
        RECT 46.480 66.650 50.330 66.800 ;
        RECT 39.130 66.200 39.430 66.650 ;
        RECT 50.030 66.200 50.330 66.650 ;
        RECT 39.130 66.050 42.980 66.200 ;
        RECT 46.480 66.050 50.330 66.200 ;
        RECT 39.130 65.600 39.430 66.050 ;
        RECT 50.030 65.600 50.330 66.050 ;
        RECT 39.130 65.450 42.980 65.600 ;
        RECT 46.480 65.450 50.330 65.600 ;
        RECT 39.130 65.000 39.430 65.450 ;
        RECT 50.030 65.000 50.330 65.450 ;
        RECT 39.130 64.850 42.980 65.000 ;
        RECT 46.480 64.850 50.330 65.000 ;
        RECT 39.130 64.400 39.430 64.850 ;
        RECT 50.030 64.400 50.330 64.850 ;
        RECT 39.130 64.250 42.980 64.400 ;
        RECT 46.480 64.250 50.330 64.400 ;
        RECT 39.130 63.800 39.430 64.250 ;
        RECT 50.030 63.800 50.330 64.250 ;
        RECT 39.130 63.650 42.980 63.800 ;
        RECT 46.480 63.650 50.330 63.800 ;
        RECT 39.130 63.200 39.430 63.650 ;
        RECT 50.030 63.200 50.330 63.650 ;
        RECT 39.130 63.050 42.980 63.200 ;
        RECT 46.480 63.050 50.330 63.200 ;
        RECT 39.130 62.600 39.430 63.050 ;
        RECT 50.030 62.600 50.330 63.050 ;
        RECT 39.130 62.450 42.980 62.600 ;
        RECT 46.480 62.450 50.330 62.600 ;
        RECT 39.130 62.000 39.430 62.450 ;
        RECT 50.030 62.000 50.330 62.450 ;
        RECT 39.130 61.450 42.930 62.000 ;
        RECT 26.530 61.400 42.930 61.450 ;
        RECT 46.530 61.450 50.330 62.000 ;
        RECT 50.780 61.450 50.930 69.650 ;
        RECT 51.380 61.450 51.530 69.650 ;
        RECT 51.980 61.450 52.130 69.650 ;
        RECT 52.580 61.450 52.730 69.650 ;
        RECT 53.180 61.450 53.330 69.650 ;
        RECT 53.780 61.450 53.930 69.650 ;
        RECT 54.380 61.450 55.080 78.550 ;
        RECT 55.530 70.350 55.680 78.550 ;
        RECT 56.130 70.350 56.280 78.550 ;
        RECT 56.730 70.350 56.880 78.550 ;
        RECT 57.330 70.350 57.480 78.550 ;
        RECT 57.930 70.350 58.080 78.550 ;
        RECT 58.530 70.350 58.680 78.550 ;
        RECT 59.130 78.000 62.930 78.550 ;
        RECT 66.530 78.550 82.930 78.600 ;
        RECT 66.530 78.000 70.330 78.550 ;
        RECT 59.130 77.550 59.430 78.000 ;
        RECT 70.030 77.550 70.330 78.000 ;
        RECT 59.130 77.400 62.980 77.550 ;
        RECT 66.480 77.400 70.330 77.550 ;
        RECT 59.130 76.950 59.430 77.400 ;
        RECT 70.030 76.950 70.330 77.400 ;
        RECT 59.130 76.800 62.980 76.950 ;
        RECT 66.480 76.800 70.330 76.950 ;
        RECT 59.130 76.350 59.430 76.800 ;
        RECT 70.030 76.350 70.330 76.800 ;
        RECT 59.130 76.200 62.980 76.350 ;
        RECT 66.480 76.200 70.330 76.350 ;
        RECT 59.130 75.750 59.430 76.200 ;
        RECT 70.030 75.750 70.330 76.200 ;
        RECT 59.130 75.600 62.980 75.750 ;
        RECT 66.480 75.600 70.330 75.750 ;
        RECT 59.130 75.150 59.430 75.600 ;
        RECT 70.030 75.150 70.330 75.600 ;
        RECT 59.130 75.000 62.980 75.150 ;
        RECT 66.480 75.000 70.330 75.150 ;
        RECT 59.130 74.550 59.430 75.000 ;
        RECT 70.030 74.550 70.330 75.000 ;
        RECT 59.130 74.400 62.980 74.550 ;
        RECT 66.480 74.400 70.330 74.550 ;
        RECT 59.130 73.950 59.430 74.400 ;
        RECT 70.030 73.950 70.330 74.400 ;
        RECT 59.130 73.800 62.980 73.950 ;
        RECT 66.480 73.800 70.330 73.950 ;
        RECT 59.130 73.350 59.430 73.800 ;
        RECT 70.030 73.350 70.330 73.800 ;
        RECT 59.130 73.200 62.980 73.350 ;
        RECT 66.480 73.200 70.330 73.350 ;
        RECT 59.130 72.750 59.430 73.200 ;
        RECT 59.130 72.600 62.980 72.750 ;
        RECT 59.130 72.150 59.430 72.600 ;
        RECT 59.130 72.000 62.980 72.150 ;
        RECT 59.130 71.550 59.430 72.000 ;
        RECT 59.130 71.400 62.980 71.550 ;
        RECT 59.130 70.950 59.430 71.400 ;
        RECT 59.130 70.800 62.980 70.950 ;
        RECT 59.130 70.350 59.430 70.800 ;
        RECT 55.530 61.450 55.680 69.650 ;
        RECT 56.130 61.450 56.280 69.650 ;
        RECT 56.730 61.450 56.880 69.650 ;
        RECT 57.330 61.450 57.480 69.650 ;
        RECT 57.930 61.450 58.080 69.650 ;
        RECT 58.530 61.450 58.680 69.650 ;
        RECT 59.130 69.200 59.430 69.650 ;
        RECT 59.130 69.050 62.980 69.200 ;
        RECT 59.130 68.600 59.430 69.050 ;
        RECT 59.130 68.450 62.980 68.600 ;
        RECT 59.130 68.000 59.430 68.450 ;
        RECT 59.130 67.850 62.980 68.000 ;
        RECT 59.130 67.400 59.430 67.850 ;
        RECT 59.130 67.250 62.980 67.400 ;
        RECT 59.130 66.800 59.430 67.250 ;
        RECT 63.830 66.800 65.630 73.200 ;
        RECT 70.030 72.750 70.330 73.200 ;
        RECT 66.480 72.600 70.330 72.750 ;
        RECT 70.030 72.150 70.330 72.600 ;
        RECT 66.480 72.000 70.330 72.150 ;
        RECT 70.030 71.550 70.330 72.000 ;
        RECT 66.480 71.400 70.330 71.550 ;
        RECT 70.030 70.950 70.330 71.400 ;
        RECT 66.480 70.800 70.330 70.950 ;
        RECT 70.030 70.350 70.330 70.800 ;
        RECT 70.780 70.350 70.930 78.550 ;
        RECT 71.380 70.350 71.530 78.550 ;
        RECT 71.980 70.350 72.130 78.550 ;
        RECT 72.580 70.350 72.730 78.550 ;
        RECT 73.180 70.350 73.330 78.550 ;
        RECT 73.780 70.350 73.930 78.550 ;
        RECT 70.030 69.200 70.330 69.650 ;
        RECT 66.480 69.050 70.330 69.200 ;
        RECT 70.030 68.600 70.330 69.050 ;
        RECT 66.480 68.450 70.330 68.600 ;
        RECT 70.030 68.000 70.330 68.450 ;
        RECT 66.480 67.850 70.330 68.000 ;
        RECT 70.030 67.400 70.330 67.850 ;
        RECT 66.480 67.250 70.330 67.400 ;
        RECT 70.030 66.800 70.330 67.250 ;
        RECT 59.130 66.650 62.980 66.800 ;
        RECT 66.480 66.650 70.330 66.800 ;
        RECT 59.130 66.200 59.430 66.650 ;
        RECT 70.030 66.200 70.330 66.650 ;
        RECT 59.130 66.050 62.980 66.200 ;
        RECT 66.480 66.050 70.330 66.200 ;
        RECT 59.130 65.600 59.430 66.050 ;
        RECT 70.030 65.600 70.330 66.050 ;
        RECT 59.130 65.450 62.980 65.600 ;
        RECT 66.480 65.450 70.330 65.600 ;
        RECT 59.130 65.000 59.430 65.450 ;
        RECT 70.030 65.000 70.330 65.450 ;
        RECT 59.130 64.850 62.980 65.000 ;
        RECT 66.480 64.850 70.330 65.000 ;
        RECT 59.130 64.400 59.430 64.850 ;
        RECT 70.030 64.400 70.330 64.850 ;
        RECT 59.130 64.250 62.980 64.400 ;
        RECT 66.480 64.250 70.330 64.400 ;
        RECT 59.130 63.800 59.430 64.250 ;
        RECT 70.030 63.800 70.330 64.250 ;
        RECT 59.130 63.650 62.980 63.800 ;
        RECT 66.480 63.650 70.330 63.800 ;
        RECT 59.130 63.200 59.430 63.650 ;
        RECT 70.030 63.200 70.330 63.650 ;
        RECT 59.130 63.050 62.980 63.200 ;
        RECT 66.480 63.050 70.330 63.200 ;
        RECT 59.130 62.600 59.430 63.050 ;
        RECT 70.030 62.600 70.330 63.050 ;
        RECT 59.130 62.450 62.980 62.600 ;
        RECT 66.480 62.450 70.330 62.600 ;
        RECT 59.130 62.000 59.430 62.450 ;
        RECT 70.030 62.000 70.330 62.450 ;
        RECT 59.130 61.450 62.930 62.000 ;
        RECT 46.530 61.400 62.930 61.450 ;
        RECT 66.530 61.450 70.330 62.000 ;
        RECT 70.780 61.450 70.930 69.650 ;
        RECT 71.380 61.450 71.530 69.650 ;
        RECT 71.980 61.450 72.130 69.650 ;
        RECT 72.580 61.450 72.730 69.650 ;
        RECT 73.180 61.450 73.330 69.650 ;
        RECT 73.780 61.450 73.930 69.650 ;
        RECT 74.380 61.450 75.080 78.550 ;
        RECT 75.530 70.350 75.680 78.550 ;
        RECT 76.130 70.350 76.280 78.550 ;
        RECT 76.730 70.350 76.880 78.550 ;
        RECT 77.330 70.350 77.480 78.550 ;
        RECT 77.930 70.350 78.080 78.550 ;
        RECT 78.530 70.350 78.680 78.550 ;
        RECT 79.130 78.000 82.930 78.550 ;
        RECT 86.530 78.550 102.930 78.600 ;
        RECT 86.530 78.000 90.330 78.550 ;
        RECT 79.130 77.550 79.430 78.000 ;
        RECT 90.030 77.550 90.330 78.000 ;
        RECT 79.130 77.400 82.980 77.550 ;
        RECT 86.480 77.400 90.330 77.550 ;
        RECT 79.130 76.950 79.430 77.400 ;
        RECT 90.030 76.950 90.330 77.400 ;
        RECT 79.130 76.800 82.980 76.950 ;
        RECT 86.480 76.800 90.330 76.950 ;
        RECT 79.130 76.350 79.430 76.800 ;
        RECT 90.030 76.350 90.330 76.800 ;
        RECT 79.130 76.200 82.980 76.350 ;
        RECT 86.480 76.200 90.330 76.350 ;
        RECT 79.130 75.750 79.430 76.200 ;
        RECT 90.030 75.750 90.330 76.200 ;
        RECT 79.130 75.600 82.980 75.750 ;
        RECT 86.480 75.600 90.330 75.750 ;
        RECT 79.130 75.150 79.430 75.600 ;
        RECT 90.030 75.150 90.330 75.600 ;
        RECT 79.130 75.000 82.980 75.150 ;
        RECT 86.480 75.000 90.330 75.150 ;
        RECT 79.130 74.550 79.430 75.000 ;
        RECT 90.030 74.550 90.330 75.000 ;
        RECT 79.130 74.400 82.980 74.550 ;
        RECT 86.480 74.400 90.330 74.550 ;
        RECT 79.130 73.950 79.430 74.400 ;
        RECT 90.030 73.950 90.330 74.400 ;
        RECT 79.130 73.800 82.980 73.950 ;
        RECT 86.480 73.800 90.330 73.950 ;
        RECT 79.130 73.350 79.430 73.800 ;
        RECT 90.030 73.350 90.330 73.800 ;
        RECT 79.130 73.200 82.980 73.350 ;
        RECT 86.480 73.200 90.330 73.350 ;
        RECT 79.130 72.750 79.430 73.200 ;
        RECT 79.130 72.600 82.980 72.750 ;
        RECT 79.130 72.150 79.430 72.600 ;
        RECT 79.130 72.000 82.980 72.150 ;
        RECT 79.130 71.550 79.430 72.000 ;
        RECT 79.130 71.400 82.980 71.550 ;
        RECT 79.130 70.950 79.430 71.400 ;
        RECT 79.130 70.800 82.980 70.950 ;
        RECT 79.130 70.350 79.430 70.800 ;
        RECT 75.530 61.450 75.680 69.650 ;
        RECT 76.130 61.450 76.280 69.650 ;
        RECT 76.730 61.450 76.880 69.650 ;
        RECT 77.330 61.450 77.480 69.650 ;
        RECT 77.930 61.450 78.080 69.650 ;
        RECT 78.530 61.450 78.680 69.650 ;
        RECT 79.130 69.200 79.430 69.650 ;
        RECT 79.130 69.050 82.980 69.200 ;
        RECT 79.130 68.600 79.430 69.050 ;
        RECT 79.130 68.450 82.980 68.600 ;
        RECT 79.130 68.000 79.430 68.450 ;
        RECT 79.130 67.850 82.980 68.000 ;
        RECT 79.130 67.400 79.430 67.850 ;
        RECT 79.130 67.250 82.980 67.400 ;
        RECT 79.130 66.800 79.430 67.250 ;
        RECT 83.830 66.800 85.630 73.200 ;
        RECT 90.030 72.750 90.330 73.200 ;
        RECT 86.480 72.600 90.330 72.750 ;
        RECT 90.030 72.150 90.330 72.600 ;
        RECT 86.480 72.000 90.330 72.150 ;
        RECT 90.030 71.550 90.330 72.000 ;
        RECT 86.480 71.400 90.330 71.550 ;
        RECT 90.030 70.950 90.330 71.400 ;
        RECT 86.480 70.800 90.330 70.950 ;
        RECT 90.030 70.350 90.330 70.800 ;
        RECT 90.780 70.350 90.930 78.550 ;
        RECT 91.380 70.350 91.530 78.550 ;
        RECT 91.980 70.350 92.130 78.550 ;
        RECT 92.580 70.350 92.730 78.550 ;
        RECT 93.180 70.350 93.330 78.550 ;
        RECT 93.780 70.350 93.930 78.550 ;
        RECT 90.030 69.200 90.330 69.650 ;
        RECT 86.480 69.050 90.330 69.200 ;
        RECT 90.030 68.600 90.330 69.050 ;
        RECT 86.480 68.450 90.330 68.600 ;
        RECT 90.030 68.000 90.330 68.450 ;
        RECT 86.480 67.850 90.330 68.000 ;
        RECT 90.030 67.400 90.330 67.850 ;
        RECT 86.480 67.250 90.330 67.400 ;
        RECT 90.030 66.800 90.330 67.250 ;
        RECT 79.130 66.650 82.980 66.800 ;
        RECT 86.480 66.650 90.330 66.800 ;
        RECT 79.130 66.200 79.430 66.650 ;
        RECT 90.030 66.200 90.330 66.650 ;
        RECT 79.130 66.050 82.980 66.200 ;
        RECT 86.480 66.050 90.330 66.200 ;
        RECT 79.130 65.600 79.430 66.050 ;
        RECT 90.030 65.600 90.330 66.050 ;
        RECT 79.130 65.450 82.980 65.600 ;
        RECT 86.480 65.450 90.330 65.600 ;
        RECT 79.130 65.000 79.430 65.450 ;
        RECT 90.030 65.000 90.330 65.450 ;
        RECT 79.130 64.850 82.980 65.000 ;
        RECT 86.480 64.850 90.330 65.000 ;
        RECT 79.130 64.400 79.430 64.850 ;
        RECT 90.030 64.400 90.330 64.850 ;
        RECT 79.130 64.250 82.980 64.400 ;
        RECT 86.480 64.250 90.330 64.400 ;
        RECT 79.130 63.800 79.430 64.250 ;
        RECT 90.030 63.800 90.330 64.250 ;
        RECT 79.130 63.650 82.980 63.800 ;
        RECT 86.480 63.650 90.330 63.800 ;
        RECT 79.130 63.200 79.430 63.650 ;
        RECT 90.030 63.200 90.330 63.650 ;
        RECT 79.130 63.050 82.980 63.200 ;
        RECT 86.480 63.050 90.330 63.200 ;
        RECT 79.130 62.600 79.430 63.050 ;
        RECT 90.030 62.600 90.330 63.050 ;
        RECT 79.130 62.450 82.980 62.600 ;
        RECT 86.480 62.450 90.330 62.600 ;
        RECT 79.130 62.000 79.430 62.450 ;
        RECT 90.030 62.000 90.330 62.450 ;
        RECT 79.130 61.450 82.930 62.000 ;
        RECT 66.530 61.400 82.930 61.450 ;
        RECT 86.530 61.450 90.330 62.000 ;
        RECT 90.780 61.450 90.930 69.650 ;
        RECT 91.380 61.450 91.530 69.650 ;
        RECT 91.980 61.450 92.130 69.650 ;
        RECT 92.580 61.450 92.730 69.650 ;
        RECT 93.180 61.450 93.330 69.650 ;
        RECT 93.780 61.450 93.930 69.650 ;
        RECT 94.380 61.450 95.080 78.550 ;
        RECT 95.530 70.350 95.680 78.550 ;
        RECT 96.130 70.350 96.280 78.550 ;
        RECT 96.730 70.350 96.880 78.550 ;
        RECT 97.330 70.350 97.480 78.550 ;
        RECT 97.930 70.350 98.080 78.550 ;
        RECT 98.530 70.350 98.680 78.550 ;
        RECT 99.130 78.000 102.930 78.550 ;
        RECT 99.130 77.550 99.430 78.000 ;
        RECT 99.130 77.400 102.980 77.550 ;
        RECT 99.130 76.950 99.430 77.400 ;
        RECT 99.130 76.800 102.980 76.950 ;
        RECT 99.130 76.350 99.430 76.800 ;
        RECT 99.130 76.200 102.980 76.350 ;
        RECT 99.130 75.750 99.430 76.200 ;
        RECT 99.130 75.600 102.980 75.750 ;
        RECT 99.130 75.150 99.430 75.600 ;
        RECT 99.130 75.000 102.980 75.150 ;
        RECT 99.130 74.550 99.430 75.000 ;
        RECT 99.130 74.400 102.980 74.550 ;
        RECT 99.130 73.950 99.430 74.400 ;
        RECT 99.130 73.800 102.980 73.950 ;
        RECT 99.130 73.350 99.430 73.800 ;
        RECT 99.130 73.200 102.980 73.350 ;
        RECT 99.130 72.750 99.430 73.200 ;
        RECT 99.130 72.600 102.980 72.750 ;
        RECT 99.130 72.150 99.430 72.600 ;
        RECT 99.130 72.000 102.980 72.150 ;
        RECT 99.130 71.550 99.430 72.000 ;
        RECT 99.130 71.400 102.980 71.550 ;
        RECT 99.130 70.950 99.430 71.400 ;
        RECT 99.130 70.800 102.980 70.950 ;
        RECT 99.130 70.350 99.430 70.800 ;
        RECT 95.530 61.450 95.680 69.650 ;
        RECT 96.130 61.450 96.280 69.650 ;
        RECT 96.730 61.450 96.880 69.650 ;
        RECT 97.330 61.450 97.480 69.650 ;
        RECT 97.930 61.450 98.080 69.650 ;
        RECT 98.530 61.450 98.680 69.650 ;
        RECT 99.130 69.200 99.430 69.650 ;
        RECT 99.130 69.050 102.980 69.200 ;
        RECT 99.130 68.600 99.430 69.050 ;
        RECT 99.130 68.450 102.980 68.600 ;
        RECT 99.130 68.000 99.430 68.450 ;
        RECT 99.130 67.850 102.980 68.000 ;
        RECT 99.130 67.400 99.430 67.850 ;
        RECT 99.130 67.250 102.980 67.400 ;
        RECT 99.130 66.800 99.430 67.250 ;
        RECT 103.830 66.800 104.730 73.200 ;
        RECT 109.850 70.130 111.850 71.405 ;
        RECT 99.130 66.650 102.980 66.800 ;
        RECT 99.130 66.200 99.430 66.650 ;
        RECT 99.130 66.050 102.980 66.200 ;
        RECT 99.130 65.600 99.430 66.050 ;
        RECT 99.130 65.450 102.980 65.600 ;
        RECT 99.130 65.000 99.430 65.450 ;
        RECT 99.130 64.850 102.980 65.000 ;
        RECT 99.130 64.400 99.430 64.850 ;
        RECT 99.130 64.250 102.980 64.400 ;
        RECT 99.130 63.800 99.430 64.250 ;
        RECT 99.130 63.650 102.980 63.800 ;
        RECT 99.130 63.200 99.430 63.650 ;
        RECT 99.130 63.050 102.980 63.200 ;
        RECT 99.130 62.600 99.430 63.050 ;
        RECT 99.130 62.450 102.980 62.600 ;
        RECT 99.130 62.000 99.430 62.450 ;
        RECT 99.130 61.450 102.930 62.000 ;
        RECT 86.530 61.400 102.930 61.450 ;
        RECT 9.630 60.900 19.830 61.400 ;
        RECT 29.630 60.900 39.830 61.400 ;
        RECT 49.630 60.900 59.830 61.400 ;
        RECT 69.630 60.900 79.830 61.400 ;
        RECT 89.630 60.900 99.830 61.400 ;
        RECT 11.530 59.100 17.930 60.900 ;
        RECT 31.530 59.100 37.930 60.900 ;
        RECT 51.530 59.100 57.930 60.900 ;
        RECT 71.530 59.100 77.930 60.900 ;
        RECT 91.530 59.100 97.930 60.900 ;
        RECT 9.630 58.600 19.830 59.100 ;
        RECT 29.630 58.600 39.830 59.100 ;
        RECT 49.630 58.600 59.830 59.100 ;
        RECT 69.630 58.600 79.830 59.100 ;
        RECT 89.630 58.600 99.830 59.100 ;
        RECT 6.530 58.550 22.930 58.600 ;
        RECT 6.530 58.000 10.330 58.550 ;
        RECT 10.030 57.550 10.330 58.000 ;
        RECT 6.480 57.400 10.330 57.550 ;
        RECT 10.030 56.950 10.330 57.400 ;
        RECT 6.480 56.800 10.330 56.950 ;
        RECT 10.030 56.350 10.330 56.800 ;
        RECT 6.480 56.200 10.330 56.350 ;
        RECT 10.030 55.750 10.330 56.200 ;
        RECT 6.480 55.600 10.330 55.750 ;
        RECT 10.030 55.150 10.330 55.600 ;
        RECT 6.480 55.000 10.330 55.150 ;
        RECT 10.030 54.550 10.330 55.000 ;
        RECT 6.480 54.400 10.330 54.550 ;
        RECT 10.030 53.950 10.330 54.400 ;
        RECT 6.480 53.800 10.330 53.950 ;
        RECT 10.030 53.350 10.330 53.800 ;
        RECT 6.480 53.200 10.330 53.350 ;
        RECT 4.730 46.800 5.630 53.200 ;
        RECT 10.030 52.750 10.330 53.200 ;
        RECT 6.480 52.600 10.330 52.750 ;
        RECT 10.030 52.150 10.330 52.600 ;
        RECT 6.480 52.000 10.330 52.150 ;
        RECT 10.030 51.550 10.330 52.000 ;
        RECT 6.480 51.400 10.330 51.550 ;
        RECT 10.030 50.950 10.330 51.400 ;
        RECT 6.480 50.800 10.330 50.950 ;
        RECT 10.030 50.350 10.330 50.800 ;
        RECT 10.780 50.350 10.930 58.550 ;
        RECT 11.380 50.350 11.530 58.550 ;
        RECT 11.980 50.350 12.130 58.550 ;
        RECT 12.580 50.350 12.730 58.550 ;
        RECT 13.180 50.350 13.330 58.550 ;
        RECT 13.780 50.350 13.930 58.550 ;
        RECT 10.030 49.200 10.330 49.650 ;
        RECT 6.480 49.050 10.330 49.200 ;
        RECT 10.030 48.600 10.330 49.050 ;
        RECT 6.480 48.450 10.330 48.600 ;
        RECT 10.030 48.000 10.330 48.450 ;
        RECT 6.480 47.850 10.330 48.000 ;
        RECT 10.030 47.400 10.330 47.850 ;
        RECT 6.480 47.250 10.330 47.400 ;
        RECT 10.030 46.800 10.330 47.250 ;
        RECT 6.480 46.650 10.330 46.800 ;
        RECT 10.030 46.200 10.330 46.650 ;
        RECT 6.480 46.050 10.330 46.200 ;
        RECT 10.030 45.600 10.330 46.050 ;
        RECT 6.480 45.450 10.330 45.600 ;
        RECT 10.030 45.000 10.330 45.450 ;
        RECT 6.480 44.850 10.330 45.000 ;
        RECT 10.030 44.400 10.330 44.850 ;
        RECT 6.480 44.250 10.330 44.400 ;
        RECT 10.030 43.800 10.330 44.250 ;
        RECT 6.480 43.650 10.330 43.800 ;
        RECT 10.030 43.200 10.330 43.650 ;
        RECT 6.480 43.050 10.330 43.200 ;
        RECT 10.030 42.600 10.330 43.050 ;
        RECT 6.480 42.450 10.330 42.600 ;
        RECT 10.030 42.000 10.330 42.450 ;
        RECT 6.530 41.450 10.330 42.000 ;
        RECT 10.780 41.450 10.930 49.650 ;
        RECT 11.380 41.450 11.530 49.650 ;
        RECT 11.980 41.450 12.130 49.650 ;
        RECT 12.580 41.450 12.730 49.650 ;
        RECT 13.180 41.450 13.330 49.650 ;
        RECT 13.780 41.450 13.930 49.650 ;
        RECT 14.380 41.450 15.080 58.550 ;
        RECT 15.530 50.350 15.680 58.550 ;
        RECT 16.130 50.350 16.280 58.550 ;
        RECT 16.730 50.350 16.880 58.550 ;
        RECT 17.330 50.350 17.480 58.550 ;
        RECT 17.930 50.350 18.080 58.550 ;
        RECT 18.530 50.350 18.680 58.550 ;
        RECT 19.130 58.000 22.930 58.550 ;
        RECT 26.530 58.550 42.930 58.600 ;
        RECT 26.530 58.000 30.330 58.550 ;
        RECT 19.130 57.550 19.430 58.000 ;
        RECT 30.030 57.550 30.330 58.000 ;
        RECT 19.130 57.400 22.980 57.550 ;
        RECT 26.480 57.400 30.330 57.550 ;
        RECT 19.130 56.950 19.430 57.400 ;
        RECT 30.030 56.950 30.330 57.400 ;
        RECT 19.130 56.800 22.980 56.950 ;
        RECT 26.480 56.800 30.330 56.950 ;
        RECT 19.130 56.350 19.430 56.800 ;
        RECT 30.030 56.350 30.330 56.800 ;
        RECT 19.130 56.200 22.980 56.350 ;
        RECT 26.480 56.200 30.330 56.350 ;
        RECT 19.130 55.750 19.430 56.200 ;
        RECT 30.030 55.750 30.330 56.200 ;
        RECT 19.130 55.600 22.980 55.750 ;
        RECT 26.480 55.600 30.330 55.750 ;
        RECT 19.130 55.150 19.430 55.600 ;
        RECT 30.030 55.150 30.330 55.600 ;
        RECT 19.130 55.000 22.980 55.150 ;
        RECT 26.480 55.000 30.330 55.150 ;
        RECT 19.130 54.550 19.430 55.000 ;
        RECT 30.030 54.550 30.330 55.000 ;
        RECT 19.130 54.400 22.980 54.550 ;
        RECT 26.480 54.400 30.330 54.550 ;
        RECT 19.130 53.950 19.430 54.400 ;
        RECT 30.030 53.950 30.330 54.400 ;
        RECT 19.130 53.800 22.980 53.950 ;
        RECT 26.480 53.800 30.330 53.950 ;
        RECT 19.130 53.350 19.430 53.800 ;
        RECT 30.030 53.350 30.330 53.800 ;
        RECT 19.130 53.200 22.980 53.350 ;
        RECT 26.480 53.200 30.330 53.350 ;
        RECT 19.130 52.750 19.430 53.200 ;
        RECT 19.130 52.600 22.980 52.750 ;
        RECT 19.130 52.150 19.430 52.600 ;
        RECT 19.130 52.000 22.980 52.150 ;
        RECT 19.130 51.550 19.430 52.000 ;
        RECT 19.130 51.400 22.980 51.550 ;
        RECT 19.130 50.950 19.430 51.400 ;
        RECT 19.130 50.800 22.980 50.950 ;
        RECT 19.130 50.350 19.430 50.800 ;
        RECT 15.530 41.450 15.680 49.650 ;
        RECT 16.130 41.450 16.280 49.650 ;
        RECT 16.730 41.450 16.880 49.650 ;
        RECT 17.330 41.450 17.480 49.650 ;
        RECT 17.930 41.450 18.080 49.650 ;
        RECT 18.530 41.450 18.680 49.650 ;
        RECT 19.130 49.200 19.430 49.650 ;
        RECT 19.130 49.050 22.980 49.200 ;
        RECT 19.130 48.600 19.430 49.050 ;
        RECT 19.130 48.450 22.980 48.600 ;
        RECT 19.130 48.000 19.430 48.450 ;
        RECT 19.130 47.850 22.980 48.000 ;
        RECT 19.130 47.400 19.430 47.850 ;
        RECT 19.130 47.250 22.980 47.400 ;
        RECT 19.130 46.800 19.430 47.250 ;
        RECT 23.830 46.800 25.630 53.200 ;
        RECT 30.030 52.750 30.330 53.200 ;
        RECT 26.480 52.600 30.330 52.750 ;
        RECT 30.030 52.150 30.330 52.600 ;
        RECT 26.480 52.000 30.330 52.150 ;
        RECT 30.030 51.550 30.330 52.000 ;
        RECT 26.480 51.400 30.330 51.550 ;
        RECT 30.030 50.950 30.330 51.400 ;
        RECT 26.480 50.800 30.330 50.950 ;
        RECT 30.030 50.350 30.330 50.800 ;
        RECT 30.780 50.350 30.930 58.550 ;
        RECT 31.380 50.350 31.530 58.550 ;
        RECT 31.980 50.350 32.130 58.550 ;
        RECT 32.580 50.350 32.730 58.550 ;
        RECT 33.180 50.350 33.330 58.550 ;
        RECT 33.780 50.350 33.930 58.550 ;
        RECT 30.030 49.200 30.330 49.650 ;
        RECT 26.480 49.050 30.330 49.200 ;
        RECT 30.030 48.600 30.330 49.050 ;
        RECT 26.480 48.450 30.330 48.600 ;
        RECT 30.030 48.000 30.330 48.450 ;
        RECT 26.480 47.850 30.330 48.000 ;
        RECT 30.030 47.400 30.330 47.850 ;
        RECT 26.480 47.250 30.330 47.400 ;
        RECT 30.030 46.800 30.330 47.250 ;
        RECT 19.130 46.650 22.980 46.800 ;
        RECT 26.480 46.650 30.330 46.800 ;
        RECT 19.130 46.200 19.430 46.650 ;
        RECT 30.030 46.200 30.330 46.650 ;
        RECT 19.130 46.050 22.980 46.200 ;
        RECT 26.480 46.050 30.330 46.200 ;
        RECT 19.130 45.600 19.430 46.050 ;
        RECT 30.030 45.600 30.330 46.050 ;
        RECT 19.130 45.450 22.980 45.600 ;
        RECT 26.480 45.450 30.330 45.600 ;
        RECT 19.130 45.000 19.430 45.450 ;
        RECT 30.030 45.000 30.330 45.450 ;
        RECT 19.130 44.850 22.980 45.000 ;
        RECT 26.480 44.850 30.330 45.000 ;
        RECT 19.130 44.400 19.430 44.850 ;
        RECT 30.030 44.400 30.330 44.850 ;
        RECT 19.130 44.250 22.980 44.400 ;
        RECT 26.480 44.250 30.330 44.400 ;
        RECT 19.130 43.800 19.430 44.250 ;
        RECT 30.030 43.800 30.330 44.250 ;
        RECT 19.130 43.650 22.980 43.800 ;
        RECT 26.480 43.650 30.330 43.800 ;
        RECT 19.130 43.200 19.430 43.650 ;
        RECT 30.030 43.200 30.330 43.650 ;
        RECT 19.130 43.050 22.980 43.200 ;
        RECT 26.480 43.050 30.330 43.200 ;
        RECT 19.130 42.600 19.430 43.050 ;
        RECT 30.030 42.600 30.330 43.050 ;
        RECT 19.130 42.450 22.980 42.600 ;
        RECT 26.480 42.450 30.330 42.600 ;
        RECT 19.130 42.000 19.430 42.450 ;
        RECT 30.030 42.000 30.330 42.450 ;
        RECT 19.130 41.450 22.930 42.000 ;
        RECT 6.530 41.400 22.930 41.450 ;
        RECT 26.530 41.450 30.330 42.000 ;
        RECT 30.780 41.450 30.930 49.650 ;
        RECT 31.380 41.450 31.530 49.650 ;
        RECT 31.980 41.450 32.130 49.650 ;
        RECT 32.580 41.450 32.730 49.650 ;
        RECT 33.180 41.450 33.330 49.650 ;
        RECT 33.780 41.450 33.930 49.650 ;
        RECT 34.380 41.450 35.080 58.550 ;
        RECT 35.530 50.350 35.680 58.550 ;
        RECT 36.130 50.350 36.280 58.550 ;
        RECT 36.730 50.350 36.880 58.550 ;
        RECT 37.330 50.350 37.480 58.550 ;
        RECT 37.930 50.350 38.080 58.550 ;
        RECT 38.530 50.350 38.680 58.550 ;
        RECT 39.130 58.000 42.930 58.550 ;
        RECT 46.530 58.550 62.930 58.600 ;
        RECT 46.530 58.000 50.330 58.550 ;
        RECT 39.130 57.550 39.430 58.000 ;
        RECT 50.030 57.550 50.330 58.000 ;
        RECT 39.130 57.400 42.980 57.550 ;
        RECT 46.480 57.400 50.330 57.550 ;
        RECT 39.130 56.950 39.430 57.400 ;
        RECT 50.030 56.950 50.330 57.400 ;
        RECT 39.130 56.800 42.980 56.950 ;
        RECT 46.480 56.800 50.330 56.950 ;
        RECT 39.130 56.350 39.430 56.800 ;
        RECT 50.030 56.350 50.330 56.800 ;
        RECT 39.130 56.200 42.980 56.350 ;
        RECT 46.480 56.200 50.330 56.350 ;
        RECT 39.130 55.750 39.430 56.200 ;
        RECT 50.030 55.750 50.330 56.200 ;
        RECT 39.130 55.600 42.980 55.750 ;
        RECT 46.480 55.600 50.330 55.750 ;
        RECT 39.130 55.150 39.430 55.600 ;
        RECT 50.030 55.150 50.330 55.600 ;
        RECT 39.130 55.000 42.980 55.150 ;
        RECT 46.480 55.000 50.330 55.150 ;
        RECT 39.130 54.550 39.430 55.000 ;
        RECT 50.030 54.550 50.330 55.000 ;
        RECT 39.130 54.400 42.980 54.550 ;
        RECT 46.480 54.400 50.330 54.550 ;
        RECT 39.130 53.950 39.430 54.400 ;
        RECT 50.030 53.950 50.330 54.400 ;
        RECT 39.130 53.800 42.980 53.950 ;
        RECT 46.480 53.800 50.330 53.950 ;
        RECT 39.130 53.350 39.430 53.800 ;
        RECT 50.030 53.350 50.330 53.800 ;
        RECT 39.130 53.200 42.980 53.350 ;
        RECT 46.480 53.200 50.330 53.350 ;
        RECT 39.130 52.750 39.430 53.200 ;
        RECT 39.130 52.600 42.980 52.750 ;
        RECT 39.130 52.150 39.430 52.600 ;
        RECT 39.130 52.000 42.980 52.150 ;
        RECT 39.130 51.550 39.430 52.000 ;
        RECT 39.130 51.400 42.980 51.550 ;
        RECT 39.130 50.950 39.430 51.400 ;
        RECT 39.130 50.800 42.980 50.950 ;
        RECT 39.130 50.350 39.430 50.800 ;
        RECT 35.530 41.450 35.680 49.650 ;
        RECT 36.130 41.450 36.280 49.650 ;
        RECT 36.730 41.450 36.880 49.650 ;
        RECT 37.330 41.450 37.480 49.650 ;
        RECT 37.930 41.450 38.080 49.650 ;
        RECT 38.530 41.450 38.680 49.650 ;
        RECT 39.130 49.200 39.430 49.650 ;
        RECT 39.130 49.050 42.980 49.200 ;
        RECT 39.130 48.600 39.430 49.050 ;
        RECT 39.130 48.450 42.980 48.600 ;
        RECT 39.130 48.000 39.430 48.450 ;
        RECT 39.130 47.850 42.980 48.000 ;
        RECT 39.130 47.400 39.430 47.850 ;
        RECT 39.130 47.250 42.980 47.400 ;
        RECT 39.130 46.800 39.430 47.250 ;
        RECT 43.830 46.800 45.630 53.200 ;
        RECT 50.030 52.750 50.330 53.200 ;
        RECT 46.480 52.600 50.330 52.750 ;
        RECT 50.030 52.150 50.330 52.600 ;
        RECT 46.480 52.000 50.330 52.150 ;
        RECT 50.030 51.550 50.330 52.000 ;
        RECT 46.480 51.400 50.330 51.550 ;
        RECT 50.030 50.950 50.330 51.400 ;
        RECT 46.480 50.800 50.330 50.950 ;
        RECT 50.030 50.350 50.330 50.800 ;
        RECT 50.780 50.350 50.930 58.550 ;
        RECT 51.380 50.350 51.530 58.550 ;
        RECT 51.980 50.350 52.130 58.550 ;
        RECT 52.580 50.350 52.730 58.550 ;
        RECT 53.180 50.350 53.330 58.550 ;
        RECT 53.780 50.350 53.930 58.550 ;
        RECT 50.030 49.200 50.330 49.650 ;
        RECT 46.480 49.050 50.330 49.200 ;
        RECT 50.030 48.600 50.330 49.050 ;
        RECT 46.480 48.450 50.330 48.600 ;
        RECT 50.030 48.000 50.330 48.450 ;
        RECT 46.480 47.850 50.330 48.000 ;
        RECT 50.030 47.400 50.330 47.850 ;
        RECT 46.480 47.250 50.330 47.400 ;
        RECT 50.030 46.800 50.330 47.250 ;
        RECT 39.130 46.650 42.980 46.800 ;
        RECT 46.480 46.650 50.330 46.800 ;
        RECT 39.130 46.200 39.430 46.650 ;
        RECT 50.030 46.200 50.330 46.650 ;
        RECT 39.130 46.050 42.980 46.200 ;
        RECT 46.480 46.050 50.330 46.200 ;
        RECT 39.130 45.600 39.430 46.050 ;
        RECT 50.030 45.600 50.330 46.050 ;
        RECT 39.130 45.450 42.980 45.600 ;
        RECT 46.480 45.450 50.330 45.600 ;
        RECT 39.130 45.000 39.430 45.450 ;
        RECT 50.030 45.000 50.330 45.450 ;
        RECT 39.130 44.850 42.980 45.000 ;
        RECT 46.480 44.850 50.330 45.000 ;
        RECT 39.130 44.400 39.430 44.850 ;
        RECT 50.030 44.400 50.330 44.850 ;
        RECT 39.130 44.250 42.980 44.400 ;
        RECT 46.480 44.250 50.330 44.400 ;
        RECT 39.130 43.800 39.430 44.250 ;
        RECT 50.030 43.800 50.330 44.250 ;
        RECT 39.130 43.650 42.980 43.800 ;
        RECT 46.480 43.650 50.330 43.800 ;
        RECT 39.130 43.200 39.430 43.650 ;
        RECT 50.030 43.200 50.330 43.650 ;
        RECT 39.130 43.050 42.980 43.200 ;
        RECT 46.480 43.050 50.330 43.200 ;
        RECT 39.130 42.600 39.430 43.050 ;
        RECT 50.030 42.600 50.330 43.050 ;
        RECT 39.130 42.450 42.980 42.600 ;
        RECT 46.480 42.450 50.330 42.600 ;
        RECT 39.130 42.000 39.430 42.450 ;
        RECT 50.030 42.000 50.330 42.450 ;
        RECT 39.130 41.450 42.930 42.000 ;
        RECT 26.530 41.400 42.930 41.450 ;
        RECT 46.530 41.450 50.330 42.000 ;
        RECT 50.780 41.450 50.930 49.650 ;
        RECT 51.380 41.450 51.530 49.650 ;
        RECT 51.980 41.450 52.130 49.650 ;
        RECT 52.580 41.450 52.730 49.650 ;
        RECT 53.180 41.450 53.330 49.650 ;
        RECT 53.780 41.450 53.930 49.650 ;
        RECT 54.380 41.450 55.080 58.550 ;
        RECT 55.530 50.350 55.680 58.550 ;
        RECT 56.130 50.350 56.280 58.550 ;
        RECT 56.730 50.350 56.880 58.550 ;
        RECT 57.330 50.350 57.480 58.550 ;
        RECT 57.930 50.350 58.080 58.550 ;
        RECT 58.530 50.350 58.680 58.550 ;
        RECT 59.130 58.000 62.930 58.550 ;
        RECT 66.530 58.550 82.930 58.600 ;
        RECT 66.530 58.000 70.330 58.550 ;
        RECT 59.130 57.550 59.430 58.000 ;
        RECT 70.030 57.550 70.330 58.000 ;
        RECT 59.130 57.400 62.980 57.550 ;
        RECT 66.480 57.400 70.330 57.550 ;
        RECT 59.130 56.950 59.430 57.400 ;
        RECT 70.030 56.950 70.330 57.400 ;
        RECT 59.130 56.800 62.980 56.950 ;
        RECT 66.480 56.800 70.330 56.950 ;
        RECT 59.130 56.350 59.430 56.800 ;
        RECT 70.030 56.350 70.330 56.800 ;
        RECT 59.130 56.200 62.980 56.350 ;
        RECT 66.480 56.200 70.330 56.350 ;
        RECT 59.130 55.750 59.430 56.200 ;
        RECT 70.030 55.750 70.330 56.200 ;
        RECT 59.130 55.600 62.980 55.750 ;
        RECT 66.480 55.600 70.330 55.750 ;
        RECT 59.130 55.150 59.430 55.600 ;
        RECT 70.030 55.150 70.330 55.600 ;
        RECT 59.130 55.000 62.980 55.150 ;
        RECT 66.480 55.000 70.330 55.150 ;
        RECT 59.130 54.550 59.430 55.000 ;
        RECT 70.030 54.550 70.330 55.000 ;
        RECT 59.130 54.400 62.980 54.550 ;
        RECT 66.480 54.400 70.330 54.550 ;
        RECT 59.130 53.950 59.430 54.400 ;
        RECT 70.030 53.950 70.330 54.400 ;
        RECT 59.130 53.800 62.980 53.950 ;
        RECT 66.480 53.800 70.330 53.950 ;
        RECT 59.130 53.350 59.430 53.800 ;
        RECT 70.030 53.350 70.330 53.800 ;
        RECT 59.130 53.200 62.980 53.350 ;
        RECT 66.480 53.200 70.330 53.350 ;
        RECT 59.130 52.750 59.430 53.200 ;
        RECT 59.130 52.600 62.980 52.750 ;
        RECT 59.130 52.150 59.430 52.600 ;
        RECT 59.130 52.000 62.980 52.150 ;
        RECT 59.130 51.550 59.430 52.000 ;
        RECT 59.130 51.400 62.980 51.550 ;
        RECT 59.130 50.950 59.430 51.400 ;
        RECT 59.130 50.800 62.980 50.950 ;
        RECT 59.130 50.350 59.430 50.800 ;
        RECT 55.530 41.450 55.680 49.650 ;
        RECT 56.130 41.450 56.280 49.650 ;
        RECT 56.730 41.450 56.880 49.650 ;
        RECT 57.330 41.450 57.480 49.650 ;
        RECT 57.930 41.450 58.080 49.650 ;
        RECT 58.530 41.450 58.680 49.650 ;
        RECT 59.130 49.200 59.430 49.650 ;
        RECT 59.130 49.050 62.980 49.200 ;
        RECT 59.130 48.600 59.430 49.050 ;
        RECT 59.130 48.450 62.980 48.600 ;
        RECT 59.130 48.000 59.430 48.450 ;
        RECT 59.130 47.850 62.980 48.000 ;
        RECT 59.130 47.400 59.430 47.850 ;
        RECT 59.130 47.250 62.980 47.400 ;
        RECT 59.130 46.800 59.430 47.250 ;
        RECT 63.830 46.800 65.630 53.200 ;
        RECT 70.030 52.750 70.330 53.200 ;
        RECT 66.480 52.600 70.330 52.750 ;
        RECT 70.030 52.150 70.330 52.600 ;
        RECT 66.480 52.000 70.330 52.150 ;
        RECT 70.030 51.550 70.330 52.000 ;
        RECT 66.480 51.400 70.330 51.550 ;
        RECT 70.030 50.950 70.330 51.400 ;
        RECT 66.480 50.800 70.330 50.950 ;
        RECT 70.030 50.350 70.330 50.800 ;
        RECT 70.780 50.350 70.930 58.550 ;
        RECT 71.380 50.350 71.530 58.550 ;
        RECT 71.980 50.350 72.130 58.550 ;
        RECT 72.580 50.350 72.730 58.550 ;
        RECT 73.180 50.350 73.330 58.550 ;
        RECT 73.780 50.350 73.930 58.550 ;
        RECT 70.030 49.200 70.330 49.650 ;
        RECT 66.480 49.050 70.330 49.200 ;
        RECT 70.030 48.600 70.330 49.050 ;
        RECT 66.480 48.450 70.330 48.600 ;
        RECT 70.030 48.000 70.330 48.450 ;
        RECT 66.480 47.850 70.330 48.000 ;
        RECT 70.030 47.400 70.330 47.850 ;
        RECT 66.480 47.250 70.330 47.400 ;
        RECT 70.030 46.800 70.330 47.250 ;
        RECT 59.130 46.650 62.980 46.800 ;
        RECT 66.480 46.650 70.330 46.800 ;
        RECT 59.130 46.200 59.430 46.650 ;
        RECT 70.030 46.200 70.330 46.650 ;
        RECT 59.130 46.050 62.980 46.200 ;
        RECT 66.480 46.050 70.330 46.200 ;
        RECT 59.130 45.600 59.430 46.050 ;
        RECT 70.030 45.600 70.330 46.050 ;
        RECT 59.130 45.450 62.980 45.600 ;
        RECT 66.480 45.450 70.330 45.600 ;
        RECT 59.130 45.000 59.430 45.450 ;
        RECT 70.030 45.000 70.330 45.450 ;
        RECT 59.130 44.850 62.980 45.000 ;
        RECT 66.480 44.850 70.330 45.000 ;
        RECT 59.130 44.400 59.430 44.850 ;
        RECT 70.030 44.400 70.330 44.850 ;
        RECT 59.130 44.250 62.980 44.400 ;
        RECT 66.480 44.250 70.330 44.400 ;
        RECT 59.130 43.800 59.430 44.250 ;
        RECT 70.030 43.800 70.330 44.250 ;
        RECT 59.130 43.650 62.980 43.800 ;
        RECT 66.480 43.650 70.330 43.800 ;
        RECT 59.130 43.200 59.430 43.650 ;
        RECT 70.030 43.200 70.330 43.650 ;
        RECT 59.130 43.050 62.980 43.200 ;
        RECT 66.480 43.050 70.330 43.200 ;
        RECT 59.130 42.600 59.430 43.050 ;
        RECT 70.030 42.600 70.330 43.050 ;
        RECT 59.130 42.450 62.980 42.600 ;
        RECT 66.480 42.450 70.330 42.600 ;
        RECT 59.130 42.000 59.430 42.450 ;
        RECT 70.030 42.000 70.330 42.450 ;
        RECT 59.130 41.450 62.930 42.000 ;
        RECT 46.530 41.400 62.930 41.450 ;
        RECT 66.530 41.450 70.330 42.000 ;
        RECT 70.780 41.450 70.930 49.650 ;
        RECT 71.380 41.450 71.530 49.650 ;
        RECT 71.980 41.450 72.130 49.650 ;
        RECT 72.580 41.450 72.730 49.650 ;
        RECT 73.180 41.450 73.330 49.650 ;
        RECT 73.780 41.450 73.930 49.650 ;
        RECT 74.380 41.450 75.080 58.550 ;
        RECT 75.530 50.350 75.680 58.550 ;
        RECT 76.130 50.350 76.280 58.550 ;
        RECT 76.730 50.350 76.880 58.550 ;
        RECT 77.330 50.350 77.480 58.550 ;
        RECT 77.930 50.350 78.080 58.550 ;
        RECT 78.530 50.350 78.680 58.550 ;
        RECT 79.130 58.000 82.930 58.550 ;
        RECT 86.530 58.550 102.930 58.600 ;
        RECT 86.530 58.000 90.330 58.550 ;
        RECT 79.130 57.550 79.430 58.000 ;
        RECT 90.030 57.550 90.330 58.000 ;
        RECT 79.130 57.400 82.980 57.550 ;
        RECT 86.480 57.400 90.330 57.550 ;
        RECT 79.130 56.950 79.430 57.400 ;
        RECT 90.030 56.950 90.330 57.400 ;
        RECT 79.130 56.800 82.980 56.950 ;
        RECT 86.480 56.800 90.330 56.950 ;
        RECT 79.130 56.350 79.430 56.800 ;
        RECT 90.030 56.350 90.330 56.800 ;
        RECT 79.130 56.200 82.980 56.350 ;
        RECT 86.480 56.200 90.330 56.350 ;
        RECT 79.130 55.750 79.430 56.200 ;
        RECT 90.030 55.750 90.330 56.200 ;
        RECT 79.130 55.600 82.980 55.750 ;
        RECT 86.480 55.600 90.330 55.750 ;
        RECT 79.130 55.150 79.430 55.600 ;
        RECT 90.030 55.150 90.330 55.600 ;
        RECT 79.130 55.000 82.980 55.150 ;
        RECT 86.480 55.000 90.330 55.150 ;
        RECT 79.130 54.550 79.430 55.000 ;
        RECT 90.030 54.550 90.330 55.000 ;
        RECT 79.130 54.400 82.980 54.550 ;
        RECT 86.480 54.400 90.330 54.550 ;
        RECT 79.130 53.950 79.430 54.400 ;
        RECT 90.030 53.950 90.330 54.400 ;
        RECT 79.130 53.800 82.980 53.950 ;
        RECT 86.480 53.800 90.330 53.950 ;
        RECT 79.130 53.350 79.430 53.800 ;
        RECT 90.030 53.350 90.330 53.800 ;
        RECT 79.130 53.200 82.980 53.350 ;
        RECT 86.480 53.200 90.330 53.350 ;
        RECT 79.130 52.750 79.430 53.200 ;
        RECT 79.130 52.600 82.980 52.750 ;
        RECT 79.130 52.150 79.430 52.600 ;
        RECT 79.130 52.000 82.980 52.150 ;
        RECT 79.130 51.550 79.430 52.000 ;
        RECT 79.130 51.400 82.980 51.550 ;
        RECT 79.130 50.950 79.430 51.400 ;
        RECT 79.130 50.800 82.980 50.950 ;
        RECT 79.130 50.350 79.430 50.800 ;
        RECT 75.530 41.450 75.680 49.650 ;
        RECT 76.130 41.450 76.280 49.650 ;
        RECT 76.730 41.450 76.880 49.650 ;
        RECT 77.330 41.450 77.480 49.650 ;
        RECT 77.930 41.450 78.080 49.650 ;
        RECT 78.530 41.450 78.680 49.650 ;
        RECT 79.130 49.200 79.430 49.650 ;
        RECT 79.130 49.050 82.980 49.200 ;
        RECT 79.130 48.600 79.430 49.050 ;
        RECT 79.130 48.450 82.980 48.600 ;
        RECT 79.130 48.000 79.430 48.450 ;
        RECT 79.130 47.850 82.980 48.000 ;
        RECT 79.130 47.400 79.430 47.850 ;
        RECT 79.130 47.250 82.980 47.400 ;
        RECT 79.130 46.800 79.430 47.250 ;
        RECT 83.830 46.800 85.630 53.200 ;
        RECT 90.030 52.750 90.330 53.200 ;
        RECT 86.480 52.600 90.330 52.750 ;
        RECT 90.030 52.150 90.330 52.600 ;
        RECT 86.480 52.000 90.330 52.150 ;
        RECT 90.030 51.550 90.330 52.000 ;
        RECT 86.480 51.400 90.330 51.550 ;
        RECT 90.030 50.950 90.330 51.400 ;
        RECT 86.480 50.800 90.330 50.950 ;
        RECT 90.030 50.350 90.330 50.800 ;
        RECT 90.780 50.350 90.930 58.550 ;
        RECT 91.380 50.350 91.530 58.550 ;
        RECT 91.980 50.350 92.130 58.550 ;
        RECT 92.580 50.350 92.730 58.550 ;
        RECT 93.180 50.350 93.330 58.550 ;
        RECT 93.780 50.350 93.930 58.550 ;
        RECT 90.030 49.200 90.330 49.650 ;
        RECT 86.480 49.050 90.330 49.200 ;
        RECT 90.030 48.600 90.330 49.050 ;
        RECT 86.480 48.450 90.330 48.600 ;
        RECT 90.030 48.000 90.330 48.450 ;
        RECT 86.480 47.850 90.330 48.000 ;
        RECT 90.030 47.400 90.330 47.850 ;
        RECT 86.480 47.250 90.330 47.400 ;
        RECT 90.030 46.800 90.330 47.250 ;
        RECT 79.130 46.650 82.980 46.800 ;
        RECT 86.480 46.650 90.330 46.800 ;
        RECT 79.130 46.200 79.430 46.650 ;
        RECT 90.030 46.200 90.330 46.650 ;
        RECT 79.130 46.050 82.980 46.200 ;
        RECT 86.480 46.050 90.330 46.200 ;
        RECT 79.130 45.600 79.430 46.050 ;
        RECT 90.030 45.600 90.330 46.050 ;
        RECT 79.130 45.450 82.980 45.600 ;
        RECT 86.480 45.450 90.330 45.600 ;
        RECT 79.130 45.000 79.430 45.450 ;
        RECT 90.030 45.000 90.330 45.450 ;
        RECT 79.130 44.850 82.980 45.000 ;
        RECT 86.480 44.850 90.330 45.000 ;
        RECT 79.130 44.400 79.430 44.850 ;
        RECT 90.030 44.400 90.330 44.850 ;
        RECT 79.130 44.250 82.980 44.400 ;
        RECT 86.480 44.250 90.330 44.400 ;
        RECT 79.130 43.800 79.430 44.250 ;
        RECT 90.030 43.800 90.330 44.250 ;
        RECT 79.130 43.650 82.980 43.800 ;
        RECT 86.480 43.650 90.330 43.800 ;
        RECT 79.130 43.200 79.430 43.650 ;
        RECT 90.030 43.200 90.330 43.650 ;
        RECT 79.130 43.050 82.980 43.200 ;
        RECT 86.480 43.050 90.330 43.200 ;
        RECT 79.130 42.600 79.430 43.050 ;
        RECT 90.030 42.600 90.330 43.050 ;
        RECT 79.130 42.450 82.980 42.600 ;
        RECT 86.480 42.450 90.330 42.600 ;
        RECT 79.130 42.000 79.430 42.450 ;
        RECT 90.030 42.000 90.330 42.450 ;
        RECT 79.130 41.450 82.930 42.000 ;
        RECT 66.530 41.400 82.930 41.450 ;
        RECT 86.530 41.450 90.330 42.000 ;
        RECT 90.780 41.450 90.930 49.650 ;
        RECT 91.380 41.450 91.530 49.650 ;
        RECT 91.980 41.450 92.130 49.650 ;
        RECT 92.580 41.450 92.730 49.650 ;
        RECT 93.180 41.450 93.330 49.650 ;
        RECT 93.780 41.450 93.930 49.650 ;
        RECT 94.380 41.450 95.080 58.550 ;
        RECT 95.530 50.350 95.680 58.550 ;
        RECT 96.130 50.350 96.280 58.550 ;
        RECT 96.730 50.350 96.880 58.550 ;
        RECT 97.330 50.350 97.480 58.550 ;
        RECT 97.930 50.350 98.080 58.550 ;
        RECT 98.530 50.350 98.680 58.550 ;
        RECT 99.130 58.000 102.930 58.550 ;
        RECT 99.130 57.550 99.430 58.000 ;
        RECT 99.130 57.400 102.980 57.550 ;
        RECT 99.130 56.950 99.430 57.400 ;
        RECT 99.130 56.800 102.980 56.950 ;
        RECT 99.130 56.350 99.430 56.800 ;
        RECT 99.130 56.200 102.980 56.350 ;
        RECT 99.130 55.750 99.430 56.200 ;
        RECT 99.130 55.600 102.980 55.750 ;
        RECT 99.130 55.150 99.430 55.600 ;
        RECT 99.130 55.000 102.980 55.150 ;
        RECT 99.130 54.550 99.430 55.000 ;
        RECT 99.130 54.400 102.980 54.550 ;
        RECT 99.130 53.950 99.430 54.400 ;
        RECT 99.130 53.800 102.980 53.950 ;
        RECT 99.130 53.350 99.430 53.800 ;
        RECT 99.130 53.200 102.980 53.350 ;
        RECT 99.130 52.750 99.430 53.200 ;
        RECT 99.130 52.600 102.980 52.750 ;
        RECT 99.130 52.150 99.430 52.600 ;
        RECT 99.130 52.000 102.980 52.150 ;
        RECT 99.130 51.550 99.430 52.000 ;
        RECT 99.130 51.400 102.980 51.550 ;
        RECT 99.130 50.950 99.430 51.400 ;
        RECT 99.130 50.800 102.980 50.950 ;
        RECT 99.130 50.350 99.430 50.800 ;
        RECT 95.530 41.450 95.680 49.650 ;
        RECT 96.130 41.450 96.280 49.650 ;
        RECT 96.730 41.450 96.880 49.650 ;
        RECT 97.330 41.450 97.480 49.650 ;
        RECT 97.930 41.450 98.080 49.650 ;
        RECT 98.530 41.450 98.680 49.650 ;
        RECT 99.130 49.200 99.430 49.650 ;
        RECT 99.130 49.050 102.980 49.200 ;
        RECT 99.130 48.600 99.430 49.050 ;
        RECT 99.130 48.450 102.980 48.600 ;
        RECT 99.130 48.000 99.430 48.450 ;
        RECT 99.130 47.850 102.980 48.000 ;
        RECT 99.130 47.400 99.430 47.850 ;
        RECT 99.130 47.250 102.980 47.400 ;
        RECT 99.130 46.800 99.430 47.250 ;
        RECT 103.830 46.800 104.730 53.200 ;
        RECT 109.850 50.310 111.850 51.585 ;
        RECT 99.130 46.650 102.980 46.800 ;
        RECT 99.130 46.200 99.430 46.650 ;
        RECT 99.130 46.050 102.980 46.200 ;
        RECT 99.130 45.600 99.430 46.050 ;
        RECT 99.130 45.450 102.980 45.600 ;
        RECT 99.130 45.000 99.430 45.450 ;
        RECT 99.130 44.850 102.980 45.000 ;
        RECT 99.130 44.400 99.430 44.850 ;
        RECT 99.130 44.250 102.980 44.400 ;
        RECT 99.130 43.800 99.430 44.250 ;
        RECT 99.130 43.650 102.980 43.800 ;
        RECT 99.130 43.200 99.430 43.650 ;
        RECT 99.130 43.050 102.980 43.200 ;
        RECT 99.130 42.600 99.430 43.050 ;
        RECT 99.130 42.450 102.980 42.600 ;
        RECT 99.130 42.000 99.430 42.450 ;
        RECT 99.130 41.450 102.930 42.000 ;
        RECT 86.530 41.400 102.930 41.450 ;
        RECT 9.630 40.900 19.830 41.400 ;
        RECT 29.630 40.900 39.830 41.400 ;
        RECT 49.630 40.900 59.830 41.400 ;
        RECT 69.630 40.900 79.830 41.400 ;
        RECT 89.630 40.900 99.830 41.400 ;
        RECT 11.530 39.100 17.930 40.900 ;
        RECT 31.530 39.100 37.930 40.900 ;
        RECT 51.530 39.100 57.930 40.900 ;
        RECT 71.530 39.100 77.930 40.900 ;
        RECT 91.530 39.100 97.930 40.900 ;
        RECT 9.630 38.600 19.830 39.100 ;
        RECT 29.630 38.600 39.830 39.100 ;
        RECT 49.630 38.600 59.830 39.100 ;
        RECT 69.630 38.600 79.830 39.100 ;
        RECT 89.630 38.600 99.830 39.100 ;
        RECT 6.530 38.550 22.930 38.600 ;
        RECT 6.530 38.000 10.330 38.550 ;
        RECT 10.030 37.550 10.330 38.000 ;
        RECT 6.480 37.400 10.330 37.550 ;
        RECT 10.030 36.950 10.330 37.400 ;
        RECT 6.480 36.800 10.330 36.950 ;
        RECT 10.030 36.350 10.330 36.800 ;
        RECT 6.480 36.200 10.330 36.350 ;
        RECT 10.030 35.750 10.330 36.200 ;
        RECT 6.480 35.600 10.330 35.750 ;
        RECT 10.030 35.150 10.330 35.600 ;
        RECT 6.480 35.000 10.330 35.150 ;
        RECT 10.030 34.550 10.330 35.000 ;
        RECT 6.480 34.400 10.330 34.550 ;
        RECT 10.030 33.950 10.330 34.400 ;
        RECT 6.480 33.800 10.330 33.950 ;
        RECT 10.030 33.350 10.330 33.800 ;
        RECT 6.480 33.200 10.330 33.350 ;
        RECT 4.730 26.800 5.630 33.200 ;
        RECT 10.030 32.750 10.330 33.200 ;
        RECT 6.480 32.600 10.330 32.750 ;
        RECT 10.030 32.150 10.330 32.600 ;
        RECT 6.480 32.000 10.330 32.150 ;
        RECT 10.030 31.550 10.330 32.000 ;
        RECT 6.480 31.400 10.330 31.550 ;
        RECT 10.030 30.950 10.330 31.400 ;
        RECT 6.480 30.800 10.330 30.950 ;
        RECT 10.030 30.350 10.330 30.800 ;
        RECT 10.780 30.350 10.930 38.550 ;
        RECT 11.380 30.350 11.530 38.550 ;
        RECT 11.980 30.350 12.130 38.550 ;
        RECT 12.580 30.350 12.730 38.550 ;
        RECT 13.180 30.350 13.330 38.550 ;
        RECT 13.780 30.350 13.930 38.550 ;
        RECT 10.030 29.200 10.330 29.650 ;
        RECT 6.480 29.050 10.330 29.200 ;
        RECT 10.030 28.600 10.330 29.050 ;
        RECT 6.480 28.450 10.330 28.600 ;
        RECT 10.030 28.000 10.330 28.450 ;
        RECT 6.480 27.850 10.330 28.000 ;
        RECT 10.030 27.400 10.330 27.850 ;
        RECT 6.480 27.250 10.330 27.400 ;
        RECT 10.030 26.800 10.330 27.250 ;
        RECT 6.480 26.650 10.330 26.800 ;
        RECT 10.030 26.200 10.330 26.650 ;
        RECT 6.480 26.050 10.330 26.200 ;
        RECT 10.030 25.600 10.330 26.050 ;
        RECT 6.480 25.450 10.330 25.600 ;
        RECT 10.030 25.000 10.330 25.450 ;
        RECT 6.480 24.850 10.330 25.000 ;
        RECT 10.030 24.400 10.330 24.850 ;
        RECT 6.480 24.250 10.330 24.400 ;
        RECT 10.030 23.800 10.330 24.250 ;
        RECT 6.480 23.650 10.330 23.800 ;
        RECT 10.030 23.200 10.330 23.650 ;
        RECT 6.480 23.050 10.330 23.200 ;
        RECT 10.030 22.600 10.330 23.050 ;
        RECT 6.480 22.450 10.330 22.600 ;
        RECT 10.030 22.000 10.330 22.450 ;
        RECT 6.530 21.450 10.330 22.000 ;
        RECT 10.780 21.450 10.930 29.650 ;
        RECT 11.380 21.450 11.530 29.650 ;
        RECT 11.980 21.450 12.130 29.650 ;
        RECT 12.580 21.450 12.730 29.650 ;
        RECT 13.180 21.450 13.330 29.650 ;
        RECT 13.780 21.450 13.930 29.650 ;
        RECT 14.380 21.450 15.080 38.550 ;
        RECT 15.530 30.350 15.680 38.550 ;
        RECT 16.130 30.350 16.280 38.550 ;
        RECT 16.730 30.350 16.880 38.550 ;
        RECT 17.330 30.350 17.480 38.550 ;
        RECT 17.930 30.350 18.080 38.550 ;
        RECT 18.530 30.350 18.680 38.550 ;
        RECT 19.130 38.000 22.930 38.550 ;
        RECT 26.530 38.550 42.930 38.600 ;
        RECT 26.530 38.000 30.330 38.550 ;
        RECT 19.130 37.550 19.430 38.000 ;
        RECT 30.030 37.550 30.330 38.000 ;
        RECT 19.130 37.400 22.980 37.550 ;
        RECT 26.480 37.400 30.330 37.550 ;
        RECT 19.130 36.950 19.430 37.400 ;
        RECT 30.030 36.950 30.330 37.400 ;
        RECT 19.130 36.800 22.980 36.950 ;
        RECT 26.480 36.800 30.330 36.950 ;
        RECT 19.130 36.350 19.430 36.800 ;
        RECT 30.030 36.350 30.330 36.800 ;
        RECT 19.130 36.200 22.980 36.350 ;
        RECT 26.480 36.200 30.330 36.350 ;
        RECT 19.130 35.750 19.430 36.200 ;
        RECT 30.030 35.750 30.330 36.200 ;
        RECT 19.130 35.600 22.980 35.750 ;
        RECT 26.480 35.600 30.330 35.750 ;
        RECT 19.130 35.150 19.430 35.600 ;
        RECT 30.030 35.150 30.330 35.600 ;
        RECT 19.130 35.000 22.980 35.150 ;
        RECT 26.480 35.000 30.330 35.150 ;
        RECT 19.130 34.550 19.430 35.000 ;
        RECT 30.030 34.550 30.330 35.000 ;
        RECT 19.130 34.400 22.980 34.550 ;
        RECT 26.480 34.400 30.330 34.550 ;
        RECT 19.130 33.950 19.430 34.400 ;
        RECT 30.030 33.950 30.330 34.400 ;
        RECT 19.130 33.800 22.980 33.950 ;
        RECT 26.480 33.800 30.330 33.950 ;
        RECT 19.130 33.350 19.430 33.800 ;
        RECT 30.030 33.350 30.330 33.800 ;
        RECT 19.130 33.200 22.980 33.350 ;
        RECT 26.480 33.200 30.330 33.350 ;
        RECT 19.130 32.750 19.430 33.200 ;
        RECT 19.130 32.600 22.980 32.750 ;
        RECT 19.130 32.150 19.430 32.600 ;
        RECT 19.130 32.000 22.980 32.150 ;
        RECT 19.130 31.550 19.430 32.000 ;
        RECT 19.130 31.400 22.980 31.550 ;
        RECT 19.130 30.950 19.430 31.400 ;
        RECT 19.130 30.800 22.980 30.950 ;
        RECT 19.130 30.350 19.430 30.800 ;
        RECT 15.530 21.450 15.680 29.650 ;
        RECT 16.130 21.450 16.280 29.650 ;
        RECT 16.730 21.450 16.880 29.650 ;
        RECT 17.330 21.450 17.480 29.650 ;
        RECT 17.930 21.450 18.080 29.650 ;
        RECT 18.530 21.450 18.680 29.650 ;
        RECT 19.130 29.200 19.430 29.650 ;
        RECT 19.130 29.050 22.980 29.200 ;
        RECT 19.130 28.600 19.430 29.050 ;
        RECT 19.130 28.450 22.980 28.600 ;
        RECT 19.130 28.000 19.430 28.450 ;
        RECT 19.130 27.850 22.980 28.000 ;
        RECT 19.130 27.400 19.430 27.850 ;
        RECT 19.130 27.250 22.980 27.400 ;
        RECT 19.130 26.800 19.430 27.250 ;
        RECT 23.830 26.800 25.630 33.200 ;
        RECT 30.030 32.750 30.330 33.200 ;
        RECT 26.480 32.600 30.330 32.750 ;
        RECT 30.030 32.150 30.330 32.600 ;
        RECT 26.480 32.000 30.330 32.150 ;
        RECT 30.030 31.550 30.330 32.000 ;
        RECT 26.480 31.400 30.330 31.550 ;
        RECT 30.030 30.950 30.330 31.400 ;
        RECT 26.480 30.800 30.330 30.950 ;
        RECT 30.030 30.350 30.330 30.800 ;
        RECT 30.780 30.350 30.930 38.550 ;
        RECT 31.380 30.350 31.530 38.550 ;
        RECT 31.980 30.350 32.130 38.550 ;
        RECT 32.580 30.350 32.730 38.550 ;
        RECT 33.180 30.350 33.330 38.550 ;
        RECT 33.780 30.350 33.930 38.550 ;
        RECT 30.030 29.200 30.330 29.650 ;
        RECT 26.480 29.050 30.330 29.200 ;
        RECT 30.030 28.600 30.330 29.050 ;
        RECT 26.480 28.450 30.330 28.600 ;
        RECT 30.030 28.000 30.330 28.450 ;
        RECT 26.480 27.850 30.330 28.000 ;
        RECT 30.030 27.400 30.330 27.850 ;
        RECT 26.480 27.250 30.330 27.400 ;
        RECT 30.030 26.800 30.330 27.250 ;
        RECT 19.130 26.650 22.980 26.800 ;
        RECT 26.480 26.650 30.330 26.800 ;
        RECT 19.130 26.200 19.430 26.650 ;
        RECT 30.030 26.200 30.330 26.650 ;
        RECT 19.130 26.050 22.980 26.200 ;
        RECT 26.480 26.050 30.330 26.200 ;
        RECT 19.130 25.600 19.430 26.050 ;
        RECT 30.030 25.600 30.330 26.050 ;
        RECT 19.130 25.450 22.980 25.600 ;
        RECT 26.480 25.450 30.330 25.600 ;
        RECT 19.130 25.000 19.430 25.450 ;
        RECT 30.030 25.000 30.330 25.450 ;
        RECT 19.130 24.850 22.980 25.000 ;
        RECT 26.480 24.850 30.330 25.000 ;
        RECT 19.130 24.400 19.430 24.850 ;
        RECT 30.030 24.400 30.330 24.850 ;
        RECT 19.130 24.250 22.980 24.400 ;
        RECT 26.480 24.250 30.330 24.400 ;
        RECT 19.130 23.800 19.430 24.250 ;
        RECT 30.030 23.800 30.330 24.250 ;
        RECT 19.130 23.650 22.980 23.800 ;
        RECT 26.480 23.650 30.330 23.800 ;
        RECT 19.130 23.200 19.430 23.650 ;
        RECT 30.030 23.200 30.330 23.650 ;
        RECT 19.130 23.050 22.980 23.200 ;
        RECT 26.480 23.050 30.330 23.200 ;
        RECT 19.130 22.600 19.430 23.050 ;
        RECT 30.030 22.600 30.330 23.050 ;
        RECT 19.130 22.450 22.980 22.600 ;
        RECT 26.480 22.450 30.330 22.600 ;
        RECT 19.130 22.000 19.430 22.450 ;
        RECT 30.030 22.000 30.330 22.450 ;
        RECT 19.130 21.450 22.930 22.000 ;
        RECT 6.530 21.400 22.930 21.450 ;
        RECT 26.530 21.450 30.330 22.000 ;
        RECT 30.780 21.450 30.930 29.650 ;
        RECT 31.380 21.450 31.530 29.650 ;
        RECT 31.980 21.450 32.130 29.650 ;
        RECT 32.580 21.450 32.730 29.650 ;
        RECT 33.180 21.450 33.330 29.650 ;
        RECT 33.780 21.450 33.930 29.650 ;
        RECT 34.380 21.450 35.080 38.550 ;
        RECT 35.530 30.350 35.680 38.550 ;
        RECT 36.130 30.350 36.280 38.550 ;
        RECT 36.730 30.350 36.880 38.550 ;
        RECT 37.330 30.350 37.480 38.550 ;
        RECT 37.930 30.350 38.080 38.550 ;
        RECT 38.530 30.350 38.680 38.550 ;
        RECT 39.130 38.000 42.930 38.550 ;
        RECT 46.530 38.550 62.930 38.600 ;
        RECT 46.530 38.000 50.330 38.550 ;
        RECT 39.130 37.550 39.430 38.000 ;
        RECT 50.030 37.550 50.330 38.000 ;
        RECT 39.130 37.400 42.980 37.550 ;
        RECT 46.480 37.400 50.330 37.550 ;
        RECT 39.130 36.950 39.430 37.400 ;
        RECT 50.030 36.950 50.330 37.400 ;
        RECT 39.130 36.800 42.980 36.950 ;
        RECT 46.480 36.800 50.330 36.950 ;
        RECT 39.130 36.350 39.430 36.800 ;
        RECT 50.030 36.350 50.330 36.800 ;
        RECT 39.130 36.200 42.980 36.350 ;
        RECT 46.480 36.200 50.330 36.350 ;
        RECT 39.130 35.750 39.430 36.200 ;
        RECT 50.030 35.750 50.330 36.200 ;
        RECT 39.130 35.600 42.980 35.750 ;
        RECT 46.480 35.600 50.330 35.750 ;
        RECT 39.130 35.150 39.430 35.600 ;
        RECT 50.030 35.150 50.330 35.600 ;
        RECT 39.130 35.000 42.980 35.150 ;
        RECT 46.480 35.000 50.330 35.150 ;
        RECT 39.130 34.550 39.430 35.000 ;
        RECT 50.030 34.550 50.330 35.000 ;
        RECT 39.130 34.400 42.980 34.550 ;
        RECT 46.480 34.400 50.330 34.550 ;
        RECT 39.130 33.950 39.430 34.400 ;
        RECT 50.030 33.950 50.330 34.400 ;
        RECT 39.130 33.800 42.980 33.950 ;
        RECT 46.480 33.800 50.330 33.950 ;
        RECT 39.130 33.350 39.430 33.800 ;
        RECT 50.030 33.350 50.330 33.800 ;
        RECT 39.130 33.200 42.980 33.350 ;
        RECT 46.480 33.200 50.330 33.350 ;
        RECT 39.130 32.750 39.430 33.200 ;
        RECT 39.130 32.600 42.980 32.750 ;
        RECT 39.130 32.150 39.430 32.600 ;
        RECT 39.130 32.000 42.980 32.150 ;
        RECT 39.130 31.550 39.430 32.000 ;
        RECT 39.130 31.400 42.980 31.550 ;
        RECT 39.130 30.950 39.430 31.400 ;
        RECT 39.130 30.800 42.980 30.950 ;
        RECT 39.130 30.350 39.430 30.800 ;
        RECT 35.530 21.450 35.680 29.650 ;
        RECT 36.130 21.450 36.280 29.650 ;
        RECT 36.730 21.450 36.880 29.650 ;
        RECT 37.330 21.450 37.480 29.650 ;
        RECT 37.930 21.450 38.080 29.650 ;
        RECT 38.530 21.450 38.680 29.650 ;
        RECT 39.130 29.200 39.430 29.650 ;
        RECT 39.130 29.050 42.980 29.200 ;
        RECT 39.130 28.600 39.430 29.050 ;
        RECT 39.130 28.450 42.980 28.600 ;
        RECT 39.130 28.000 39.430 28.450 ;
        RECT 39.130 27.850 42.980 28.000 ;
        RECT 39.130 27.400 39.430 27.850 ;
        RECT 39.130 27.250 42.980 27.400 ;
        RECT 39.130 26.800 39.430 27.250 ;
        RECT 43.830 26.800 45.630 33.200 ;
        RECT 50.030 32.750 50.330 33.200 ;
        RECT 46.480 32.600 50.330 32.750 ;
        RECT 50.030 32.150 50.330 32.600 ;
        RECT 46.480 32.000 50.330 32.150 ;
        RECT 50.030 31.550 50.330 32.000 ;
        RECT 46.480 31.400 50.330 31.550 ;
        RECT 50.030 30.950 50.330 31.400 ;
        RECT 46.480 30.800 50.330 30.950 ;
        RECT 50.030 30.350 50.330 30.800 ;
        RECT 50.780 30.350 50.930 38.550 ;
        RECT 51.380 30.350 51.530 38.550 ;
        RECT 51.980 30.350 52.130 38.550 ;
        RECT 52.580 30.350 52.730 38.550 ;
        RECT 53.180 30.350 53.330 38.550 ;
        RECT 53.780 30.350 53.930 38.550 ;
        RECT 50.030 29.200 50.330 29.650 ;
        RECT 46.480 29.050 50.330 29.200 ;
        RECT 50.030 28.600 50.330 29.050 ;
        RECT 46.480 28.450 50.330 28.600 ;
        RECT 50.030 28.000 50.330 28.450 ;
        RECT 46.480 27.850 50.330 28.000 ;
        RECT 50.030 27.400 50.330 27.850 ;
        RECT 46.480 27.250 50.330 27.400 ;
        RECT 50.030 26.800 50.330 27.250 ;
        RECT 39.130 26.650 42.980 26.800 ;
        RECT 46.480 26.650 50.330 26.800 ;
        RECT 39.130 26.200 39.430 26.650 ;
        RECT 50.030 26.200 50.330 26.650 ;
        RECT 39.130 26.050 42.980 26.200 ;
        RECT 46.480 26.050 50.330 26.200 ;
        RECT 39.130 25.600 39.430 26.050 ;
        RECT 50.030 25.600 50.330 26.050 ;
        RECT 39.130 25.450 42.980 25.600 ;
        RECT 46.480 25.450 50.330 25.600 ;
        RECT 39.130 25.000 39.430 25.450 ;
        RECT 50.030 25.000 50.330 25.450 ;
        RECT 39.130 24.850 42.980 25.000 ;
        RECT 46.480 24.850 50.330 25.000 ;
        RECT 39.130 24.400 39.430 24.850 ;
        RECT 50.030 24.400 50.330 24.850 ;
        RECT 39.130 24.250 42.980 24.400 ;
        RECT 46.480 24.250 50.330 24.400 ;
        RECT 39.130 23.800 39.430 24.250 ;
        RECT 50.030 23.800 50.330 24.250 ;
        RECT 39.130 23.650 42.980 23.800 ;
        RECT 46.480 23.650 50.330 23.800 ;
        RECT 39.130 23.200 39.430 23.650 ;
        RECT 50.030 23.200 50.330 23.650 ;
        RECT 39.130 23.050 42.980 23.200 ;
        RECT 46.480 23.050 50.330 23.200 ;
        RECT 39.130 22.600 39.430 23.050 ;
        RECT 50.030 22.600 50.330 23.050 ;
        RECT 39.130 22.450 42.980 22.600 ;
        RECT 46.480 22.450 50.330 22.600 ;
        RECT 39.130 22.000 39.430 22.450 ;
        RECT 50.030 22.000 50.330 22.450 ;
        RECT 39.130 21.450 42.930 22.000 ;
        RECT 26.530 21.400 42.930 21.450 ;
        RECT 46.530 21.450 50.330 22.000 ;
        RECT 50.780 21.450 50.930 29.650 ;
        RECT 51.380 21.450 51.530 29.650 ;
        RECT 51.980 21.450 52.130 29.650 ;
        RECT 52.580 21.450 52.730 29.650 ;
        RECT 53.180 21.450 53.330 29.650 ;
        RECT 53.780 21.450 53.930 29.650 ;
        RECT 54.380 21.450 55.080 38.550 ;
        RECT 55.530 30.350 55.680 38.550 ;
        RECT 56.130 30.350 56.280 38.550 ;
        RECT 56.730 30.350 56.880 38.550 ;
        RECT 57.330 30.350 57.480 38.550 ;
        RECT 57.930 30.350 58.080 38.550 ;
        RECT 58.530 30.350 58.680 38.550 ;
        RECT 59.130 38.000 62.930 38.550 ;
        RECT 66.530 38.550 82.930 38.600 ;
        RECT 66.530 38.000 70.330 38.550 ;
        RECT 59.130 37.550 59.430 38.000 ;
        RECT 70.030 37.550 70.330 38.000 ;
        RECT 59.130 37.400 62.980 37.550 ;
        RECT 66.480 37.400 70.330 37.550 ;
        RECT 59.130 36.950 59.430 37.400 ;
        RECT 70.030 36.950 70.330 37.400 ;
        RECT 59.130 36.800 62.980 36.950 ;
        RECT 66.480 36.800 70.330 36.950 ;
        RECT 59.130 36.350 59.430 36.800 ;
        RECT 70.030 36.350 70.330 36.800 ;
        RECT 59.130 36.200 62.980 36.350 ;
        RECT 66.480 36.200 70.330 36.350 ;
        RECT 59.130 35.750 59.430 36.200 ;
        RECT 70.030 35.750 70.330 36.200 ;
        RECT 59.130 35.600 62.980 35.750 ;
        RECT 66.480 35.600 70.330 35.750 ;
        RECT 59.130 35.150 59.430 35.600 ;
        RECT 70.030 35.150 70.330 35.600 ;
        RECT 59.130 35.000 62.980 35.150 ;
        RECT 66.480 35.000 70.330 35.150 ;
        RECT 59.130 34.550 59.430 35.000 ;
        RECT 70.030 34.550 70.330 35.000 ;
        RECT 59.130 34.400 62.980 34.550 ;
        RECT 66.480 34.400 70.330 34.550 ;
        RECT 59.130 33.950 59.430 34.400 ;
        RECT 70.030 33.950 70.330 34.400 ;
        RECT 59.130 33.800 62.980 33.950 ;
        RECT 66.480 33.800 70.330 33.950 ;
        RECT 59.130 33.350 59.430 33.800 ;
        RECT 70.030 33.350 70.330 33.800 ;
        RECT 59.130 33.200 62.980 33.350 ;
        RECT 66.480 33.200 70.330 33.350 ;
        RECT 59.130 32.750 59.430 33.200 ;
        RECT 59.130 32.600 62.980 32.750 ;
        RECT 59.130 32.150 59.430 32.600 ;
        RECT 59.130 32.000 62.980 32.150 ;
        RECT 59.130 31.550 59.430 32.000 ;
        RECT 59.130 31.400 62.980 31.550 ;
        RECT 59.130 30.950 59.430 31.400 ;
        RECT 59.130 30.800 62.980 30.950 ;
        RECT 59.130 30.350 59.430 30.800 ;
        RECT 55.530 21.450 55.680 29.650 ;
        RECT 56.130 21.450 56.280 29.650 ;
        RECT 56.730 21.450 56.880 29.650 ;
        RECT 57.330 21.450 57.480 29.650 ;
        RECT 57.930 21.450 58.080 29.650 ;
        RECT 58.530 21.450 58.680 29.650 ;
        RECT 59.130 29.200 59.430 29.650 ;
        RECT 59.130 29.050 62.980 29.200 ;
        RECT 59.130 28.600 59.430 29.050 ;
        RECT 59.130 28.450 62.980 28.600 ;
        RECT 59.130 28.000 59.430 28.450 ;
        RECT 59.130 27.850 62.980 28.000 ;
        RECT 59.130 27.400 59.430 27.850 ;
        RECT 59.130 27.250 62.980 27.400 ;
        RECT 59.130 26.800 59.430 27.250 ;
        RECT 63.830 26.800 65.630 33.200 ;
        RECT 70.030 32.750 70.330 33.200 ;
        RECT 66.480 32.600 70.330 32.750 ;
        RECT 70.030 32.150 70.330 32.600 ;
        RECT 66.480 32.000 70.330 32.150 ;
        RECT 70.030 31.550 70.330 32.000 ;
        RECT 66.480 31.400 70.330 31.550 ;
        RECT 70.030 30.950 70.330 31.400 ;
        RECT 66.480 30.800 70.330 30.950 ;
        RECT 70.030 30.350 70.330 30.800 ;
        RECT 70.780 30.350 70.930 38.550 ;
        RECT 71.380 30.350 71.530 38.550 ;
        RECT 71.980 30.350 72.130 38.550 ;
        RECT 72.580 30.350 72.730 38.550 ;
        RECT 73.180 30.350 73.330 38.550 ;
        RECT 73.780 30.350 73.930 38.550 ;
        RECT 70.030 29.200 70.330 29.650 ;
        RECT 66.480 29.050 70.330 29.200 ;
        RECT 70.030 28.600 70.330 29.050 ;
        RECT 66.480 28.450 70.330 28.600 ;
        RECT 70.030 28.000 70.330 28.450 ;
        RECT 66.480 27.850 70.330 28.000 ;
        RECT 70.030 27.400 70.330 27.850 ;
        RECT 66.480 27.250 70.330 27.400 ;
        RECT 70.030 26.800 70.330 27.250 ;
        RECT 59.130 26.650 62.980 26.800 ;
        RECT 66.480 26.650 70.330 26.800 ;
        RECT 59.130 26.200 59.430 26.650 ;
        RECT 70.030 26.200 70.330 26.650 ;
        RECT 59.130 26.050 62.980 26.200 ;
        RECT 66.480 26.050 70.330 26.200 ;
        RECT 59.130 25.600 59.430 26.050 ;
        RECT 70.030 25.600 70.330 26.050 ;
        RECT 59.130 25.450 62.980 25.600 ;
        RECT 66.480 25.450 70.330 25.600 ;
        RECT 59.130 25.000 59.430 25.450 ;
        RECT 70.030 25.000 70.330 25.450 ;
        RECT 59.130 24.850 62.980 25.000 ;
        RECT 66.480 24.850 70.330 25.000 ;
        RECT 59.130 24.400 59.430 24.850 ;
        RECT 70.030 24.400 70.330 24.850 ;
        RECT 59.130 24.250 62.980 24.400 ;
        RECT 66.480 24.250 70.330 24.400 ;
        RECT 59.130 23.800 59.430 24.250 ;
        RECT 70.030 23.800 70.330 24.250 ;
        RECT 59.130 23.650 62.980 23.800 ;
        RECT 66.480 23.650 70.330 23.800 ;
        RECT 59.130 23.200 59.430 23.650 ;
        RECT 70.030 23.200 70.330 23.650 ;
        RECT 59.130 23.050 62.980 23.200 ;
        RECT 66.480 23.050 70.330 23.200 ;
        RECT 59.130 22.600 59.430 23.050 ;
        RECT 70.030 22.600 70.330 23.050 ;
        RECT 59.130 22.450 62.980 22.600 ;
        RECT 66.480 22.450 70.330 22.600 ;
        RECT 59.130 22.000 59.430 22.450 ;
        RECT 70.030 22.000 70.330 22.450 ;
        RECT 59.130 21.450 62.930 22.000 ;
        RECT 46.530 21.400 62.930 21.450 ;
        RECT 66.530 21.450 70.330 22.000 ;
        RECT 70.780 21.450 70.930 29.650 ;
        RECT 71.380 21.450 71.530 29.650 ;
        RECT 71.980 21.450 72.130 29.650 ;
        RECT 72.580 21.450 72.730 29.650 ;
        RECT 73.180 21.450 73.330 29.650 ;
        RECT 73.780 21.450 73.930 29.650 ;
        RECT 74.380 21.450 75.080 38.550 ;
        RECT 75.530 30.350 75.680 38.550 ;
        RECT 76.130 30.350 76.280 38.550 ;
        RECT 76.730 30.350 76.880 38.550 ;
        RECT 77.330 30.350 77.480 38.550 ;
        RECT 77.930 30.350 78.080 38.550 ;
        RECT 78.530 30.350 78.680 38.550 ;
        RECT 79.130 38.000 82.930 38.550 ;
        RECT 86.530 38.550 102.930 38.600 ;
        RECT 86.530 38.000 90.330 38.550 ;
        RECT 79.130 37.550 79.430 38.000 ;
        RECT 90.030 37.550 90.330 38.000 ;
        RECT 79.130 37.400 82.980 37.550 ;
        RECT 86.480 37.400 90.330 37.550 ;
        RECT 79.130 36.950 79.430 37.400 ;
        RECT 90.030 36.950 90.330 37.400 ;
        RECT 79.130 36.800 82.980 36.950 ;
        RECT 86.480 36.800 90.330 36.950 ;
        RECT 79.130 36.350 79.430 36.800 ;
        RECT 90.030 36.350 90.330 36.800 ;
        RECT 79.130 36.200 82.980 36.350 ;
        RECT 86.480 36.200 90.330 36.350 ;
        RECT 79.130 35.750 79.430 36.200 ;
        RECT 90.030 35.750 90.330 36.200 ;
        RECT 79.130 35.600 82.980 35.750 ;
        RECT 86.480 35.600 90.330 35.750 ;
        RECT 79.130 35.150 79.430 35.600 ;
        RECT 90.030 35.150 90.330 35.600 ;
        RECT 79.130 35.000 82.980 35.150 ;
        RECT 86.480 35.000 90.330 35.150 ;
        RECT 79.130 34.550 79.430 35.000 ;
        RECT 90.030 34.550 90.330 35.000 ;
        RECT 79.130 34.400 82.980 34.550 ;
        RECT 86.480 34.400 90.330 34.550 ;
        RECT 79.130 33.950 79.430 34.400 ;
        RECT 90.030 33.950 90.330 34.400 ;
        RECT 79.130 33.800 82.980 33.950 ;
        RECT 86.480 33.800 90.330 33.950 ;
        RECT 79.130 33.350 79.430 33.800 ;
        RECT 90.030 33.350 90.330 33.800 ;
        RECT 79.130 33.200 82.980 33.350 ;
        RECT 86.480 33.200 90.330 33.350 ;
        RECT 79.130 32.750 79.430 33.200 ;
        RECT 79.130 32.600 82.980 32.750 ;
        RECT 79.130 32.150 79.430 32.600 ;
        RECT 79.130 32.000 82.980 32.150 ;
        RECT 79.130 31.550 79.430 32.000 ;
        RECT 79.130 31.400 82.980 31.550 ;
        RECT 79.130 30.950 79.430 31.400 ;
        RECT 79.130 30.800 82.980 30.950 ;
        RECT 79.130 30.350 79.430 30.800 ;
        RECT 75.530 21.450 75.680 29.650 ;
        RECT 76.130 21.450 76.280 29.650 ;
        RECT 76.730 21.450 76.880 29.650 ;
        RECT 77.330 21.450 77.480 29.650 ;
        RECT 77.930 21.450 78.080 29.650 ;
        RECT 78.530 21.450 78.680 29.650 ;
        RECT 79.130 29.200 79.430 29.650 ;
        RECT 79.130 29.050 82.980 29.200 ;
        RECT 79.130 28.600 79.430 29.050 ;
        RECT 79.130 28.450 82.980 28.600 ;
        RECT 79.130 28.000 79.430 28.450 ;
        RECT 79.130 27.850 82.980 28.000 ;
        RECT 79.130 27.400 79.430 27.850 ;
        RECT 79.130 27.250 82.980 27.400 ;
        RECT 79.130 26.800 79.430 27.250 ;
        RECT 83.830 26.800 85.630 33.200 ;
        RECT 90.030 32.750 90.330 33.200 ;
        RECT 86.480 32.600 90.330 32.750 ;
        RECT 90.030 32.150 90.330 32.600 ;
        RECT 86.480 32.000 90.330 32.150 ;
        RECT 90.030 31.550 90.330 32.000 ;
        RECT 86.480 31.400 90.330 31.550 ;
        RECT 90.030 30.950 90.330 31.400 ;
        RECT 86.480 30.800 90.330 30.950 ;
        RECT 90.030 30.350 90.330 30.800 ;
        RECT 90.780 30.350 90.930 38.550 ;
        RECT 91.380 30.350 91.530 38.550 ;
        RECT 91.980 30.350 92.130 38.550 ;
        RECT 92.580 30.350 92.730 38.550 ;
        RECT 93.180 30.350 93.330 38.550 ;
        RECT 93.780 30.350 93.930 38.550 ;
        RECT 90.030 29.200 90.330 29.650 ;
        RECT 86.480 29.050 90.330 29.200 ;
        RECT 90.030 28.600 90.330 29.050 ;
        RECT 86.480 28.450 90.330 28.600 ;
        RECT 90.030 28.000 90.330 28.450 ;
        RECT 86.480 27.850 90.330 28.000 ;
        RECT 90.030 27.400 90.330 27.850 ;
        RECT 86.480 27.250 90.330 27.400 ;
        RECT 90.030 26.800 90.330 27.250 ;
        RECT 79.130 26.650 82.980 26.800 ;
        RECT 86.480 26.650 90.330 26.800 ;
        RECT 79.130 26.200 79.430 26.650 ;
        RECT 90.030 26.200 90.330 26.650 ;
        RECT 79.130 26.050 82.980 26.200 ;
        RECT 86.480 26.050 90.330 26.200 ;
        RECT 79.130 25.600 79.430 26.050 ;
        RECT 90.030 25.600 90.330 26.050 ;
        RECT 79.130 25.450 82.980 25.600 ;
        RECT 86.480 25.450 90.330 25.600 ;
        RECT 79.130 25.000 79.430 25.450 ;
        RECT 90.030 25.000 90.330 25.450 ;
        RECT 79.130 24.850 82.980 25.000 ;
        RECT 86.480 24.850 90.330 25.000 ;
        RECT 79.130 24.400 79.430 24.850 ;
        RECT 90.030 24.400 90.330 24.850 ;
        RECT 79.130 24.250 82.980 24.400 ;
        RECT 86.480 24.250 90.330 24.400 ;
        RECT 79.130 23.800 79.430 24.250 ;
        RECT 90.030 23.800 90.330 24.250 ;
        RECT 79.130 23.650 82.980 23.800 ;
        RECT 86.480 23.650 90.330 23.800 ;
        RECT 79.130 23.200 79.430 23.650 ;
        RECT 90.030 23.200 90.330 23.650 ;
        RECT 79.130 23.050 82.980 23.200 ;
        RECT 86.480 23.050 90.330 23.200 ;
        RECT 79.130 22.600 79.430 23.050 ;
        RECT 90.030 22.600 90.330 23.050 ;
        RECT 79.130 22.450 82.980 22.600 ;
        RECT 86.480 22.450 90.330 22.600 ;
        RECT 79.130 22.000 79.430 22.450 ;
        RECT 90.030 22.000 90.330 22.450 ;
        RECT 79.130 21.450 82.930 22.000 ;
        RECT 66.530 21.400 82.930 21.450 ;
        RECT 86.530 21.450 90.330 22.000 ;
        RECT 90.780 21.450 90.930 29.650 ;
        RECT 91.380 21.450 91.530 29.650 ;
        RECT 91.980 21.450 92.130 29.650 ;
        RECT 92.580 21.450 92.730 29.650 ;
        RECT 93.180 21.450 93.330 29.650 ;
        RECT 93.780 21.450 93.930 29.650 ;
        RECT 94.380 21.450 95.080 38.550 ;
        RECT 95.530 30.350 95.680 38.550 ;
        RECT 96.130 30.350 96.280 38.550 ;
        RECT 96.730 30.350 96.880 38.550 ;
        RECT 97.330 30.350 97.480 38.550 ;
        RECT 97.930 30.350 98.080 38.550 ;
        RECT 98.530 30.350 98.680 38.550 ;
        RECT 99.130 38.000 102.930 38.550 ;
        RECT 99.130 37.550 99.430 38.000 ;
        RECT 99.130 37.400 102.980 37.550 ;
        RECT 99.130 36.950 99.430 37.400 ;
        RECT 99.130 36.800 102.980 36.950 ;
        RECT 99.130 36.350 99.430 36.800 ;
        RECT 99.130 36.200 102.980 36.350 ;
        RECT 99.130 35.750 99.430 36.200 ;
        RECT 99.130 35.600 102.980 35.750 ;
        RECT 99.130 35.150 99.430 35.600 ;
        RECT 99.130 35.000 102.980 35.150 ;
        RECT 99.130 34.550 99.430 35.000 ;
        RECT 99.130 34.400 102.980 34.550 ;
        RECT 99.130 33.950 99.430 34.400 ;
        RECT 99.130 33.800 102.980 33.950 ;
        RECT 99.130 33.350 99.430 33.800 ;
        RECT 99.130 33.200 102.980 33.350 ;
        RECT 99.130 32.750 99.430 33.200 ;
        RECT 99.130 32.600 102.980 32.750 ;
        RECT 99.130 32.150 99.430 32.600 ;
        RECT 99.130 32.000 102.980 32.150 ;
        RECT 99.130 31.550 99.430 32.000 ;
        RECT 99.130 31.400 102.980 31.550 ;
        RECT 99.130 30.950 99.430 31.400 ;
        RECT 99.130 30.800 102.980 30.950 ;
        RECT 99.130 30.350 99.430 30.800 ;
        RECT 95.530 21.450 95.680 29.650 ;
        RECT 96.130 21.450 96.280 29.650 ;
        RECT 96.730 21.450 96.880 29.650 ;
        RECT 97.330 21.450 97.480 29.650 ;
        RECT 97.930 21.450 98.080 29.650 ;
        RECT 98.530 21.450 98.680 29.650 ;
        RECT 99.130 29.200 99.430 29.650 ;
        RECT 99.130 29.050 102.980 29.200 ;
        RECT 99.130 28.600 99.430 29.050 ;
        RECT 99.130 28.450 102.980 28.600 ;
        RECT 99.130 28.000 99.430 28.450 ;
        RECT 99.130 27.850 102.980 28.000 ;
        RECT 99.130 27.400 99.430 27.850 ;
        RECT 99.130 27.250 102.980 27.400 ;
        RECT 99.130 26.800 99.430 27.250 ;
        RECT 103.830 26.800 104.730 33.200 ;
        RECT 109.850 30.250 111.850 31.525 ;
        RECT 99.130 26.650 102.980 26.800 ;
        RECT 99.130 26.200 99.430 26.650 ;
        RECT 99.130 26.050 102.980 26.200 ;
        RECT 99.130 25.600 99.430 26.050 ;
        RECT 99.130 25.450 102.980 25.600 ;
        RECT 99.130 25.000 99.430 25.450 ;
        RECT 99.130 24.850 102.980 25.000 ;
        RECT 99.130 24.400 99.430 24.850 ;
        RECT 99.130 24.250 102.980 24.400 ;
        RECT 99.130 23.800 99.430 24.250 ;
        RECT 99.130 23.650 102.980 23.800 ;
        RECT 99.130 23.200 99.430 23.650 ;
        RECT 99.130 23.050 102.980 23.200 ;
        RECT 99.130 22.600 99.430 23.050 ;
        RECT 99.130 22.450 102.980 22.600 ;
        RECT 99.130 22.000 99.430 22.450 ;
        RECT 99.130 21.450 102.930 22.000 ;
        RECT 86.530 21.400 102.930 21.450 ;
        RECT 9.630 20.900 19.830 21.400 ;
        RECT 29.630 20.900 39.830 21.400 ;
        RECT 49.630 20.900 59.830 21.400 ;
        RECT 69.630 20.900 79.830 21.400 ;
        RECT 89.630 20.900 99.830 21.400 ;
        RECT 11.530 19.100 17.930 20.900 ;
        RECT 31.530 19.100 37.930 20.900 ;
        RECT 51.530 19.100 57.930 20.900 ;
        RECT 71.530 19.100 77.930 20.900 ;
        RECT 91.530 19.100 97.930 20.900 ;
        RECT 9.630 18.600 19.830 19.100 ;
        RECT 29.630 18.600 39.830 19.100 ;
        RECT 49.630 18.600 59.830 19.100 ;
        RECT 69.630 18.600 79.830 19.100 ;
        RECT 89.630 18.600 99.830 19.100 ;
        RECT 6.530 18.550 22.930 18.600 ;
        RECT 6.530 18.000 10.330 18.550 ;
        RECT 10.030 17.550 10.330 18.000 ;
        RECT 6.480 17.400 10.330 17.550 ;
        RECT 10.030 16.950 10.330 17.400 ;
        RECT 6.480 16.800 10.330 16.950 ;
        RECT 10.030 16.350 10.330 16.800 ;
        RECT 6.480 16.200 10.330 16.350 ;
        RECT 10.030 15.750 10.330 16.200 ;
        RECT 6.480 15.600 10.330 15.750 ;
        RECT 10.030 15.150 10.330 15.600 ;
        RECT 6.480 15.000 10.330 15.150 ;
        RECT 10.030 14.550 10.330 15.000 ;
        RECT 6.480 14.400 10.330 14.550 ;
        RECT 10.030 13.950 10.330 14.400 ;
        RECT 6.480 13.800 10.330 13.950 ;
        RECT 10.030 13.350 10.330 13.800 ;
        RECT 6.480 13.200 10.330 13.350 ;
        RECT 4.730 6.800 5.630 13.200 ;
        RECT 10.030 12.750 10.330 13.200 ;
        RECT 6.480 12.600 10.330 12.750 ;
        RECT 10.030 12.150 10.330 12.600 ;
        RECT 6.480 12.000 10.330 12.150 ;
        RECT 10.030 11.550 10.330 12.000 ;
        RECT 6.480 11.400 10.330 11.550 ;
        RECT 10.030 10.950 10.330 11.400 ;
        RECT 6.480 10.800 10.330 10.950 ;
        RECT 10.030 10.350 10.330 10.800 ;
        RECT 10.780 10.350 10.930 18.550 ;
        RECT 11.380 10.350 11.530 18.550 ;
        RECT 11.980 10.350 12.130 18.550 ;
        RECT 12.580 10.350 12.730 18.550 ;
        RECT 13.180 10.350 13.330 18.550 ;
        RECT 13.780 10.350 13.930 18.550 ;
        RECT 10.030 9.200 10.330 9.650 ;
        RECT 6.480 9.050 10.330 9.200 ;
        RECT 10.030 8.600 10.330 9.050 ;
        RECT 6.480 8.450 10.330 8.600 ;
        RECT 10.030 8.000 10.330 8.450 ;
        RECT 6.480 7.850 10.330 8.000 ;
        RECT 10.030 7.400 10.330 7.850 ;
        RECT 6.480 7.250 10.330 7.400 ;
        RECT 10.030 6.800 10.330 7.250 ;
        RECT 6.480 6.650 10.330 6.800 ;
        RECT 10.030 6.200 10.330 6.650 ;
        RECT 6.480 6.050 10.330 6.200 ;
        RECT 10.030 5.600 10.330 6.050 ;
        RECT 6.480 5.450 10.330 5.600 ;
        RECT 10.030 5.000 10.330 5.450 ;
        RECT 6.480 4.850 10.330 5.000 ;
        RECT 10.030 4.400 10.330 4.850 ;
        RECT 6.480 4.250 10.330 4.400 ;
        RECT 10.030 3.800 10.330 4.250 ;
        RECT 6.480 3.650 10.330 3.800 ;
        RECT 10.030 3.200 10.330 3.650 ;
        RECT 6.480 3.050 10.330 3.200 ;
        RECT 10.030 2.600 10.330 3.050 ;
        RECT 6.480 2.450 10.330 2.600 ;
        RECT 10.030 2.000 10.330 2.450 ;
        RECT 6.530 1.450 10.330 2.000 ;
        RECT 10.780 1.450 10.930 9.650 ;
        RECT 11.380 1.450 11.530 9.650 ;
        RECT 11.980 1.450 12.130 9.650 ;
        RECT 12.580 1.450 12.730 9.650 ;
        RECT 13.180 1.450 13.330 9.650 ;
        RECT 13.780 1.450 13.930 9.650 ;
        RECT 14.380 1.450 15.080 18.550 ;
        RECT 15.530 10.350 15.680 18.550 ;
        RECT 16.130 10.350 16.280 18.550 ;
        RECT 16.730 10.350 16.880 18.550 ;
        RECT 17.330 10.350 17.480 18.550 ;
        RECT 17.930 10.350 18.080 18.550 ;
        RECT 18.530 10.350 18.680 18.550 ;
        RECT 19.130 18.000 22.930 18.550 ;
        RECT 26.530 18.550 42.930 18.600 ;
        RECT 26.530 18.000 30.330 18.550 ;
        RECT 19.130 17.550 19.430 18.000 ;
        RECT 30.030 17.550 30.330 18.000 ;
        RECT 19.130 17.400 22.980 17.550 ;
        RECT 26.480 17.400 30.330 17.550 ;
        RECT 19.130 16.950 19.430 17.400 ;
        RECT 30.030 16.950 30.330 17.400 ;
        RECT 19.130 16.800 22.980 16.950 ;
        RECT 26.480 16.800 30.330 16.950 ;
        RECT 19.130 16.350 19.430 16.800 ;
        RECT 30.030 16.350 30.330 16.800 ;
        RECT 19.130 16.200 22.980 16.350 ;
        RECT 26.480 16.200 30.330 16.350 ;
        RECT 19.130 15.750 19.430 16.200 ;
        RECT 30.030 15.750 30.330 16.200 ;
        RECT 19.130 15.600 22.980 15.750 ;
        RECT 26.480 15.600 30.330 15.750 ;
        RECT 19.130 15.150 19.430 15.600 ;
        RECT 30.030 15.150 30.330 15.600 ;
        RECT 19.130 15.000 22.980 15.150 ;
        RECT 26.480 15.000 30.330 15.150 ;
        RECT 19.130 14.550 19.430 15.000 ;
        RECT 30.030 14.550 30.330 15.000 ;
        RECT 19.130 14.400 22.980 14.550 ;
        RECT 26.480 14.400 30.330 14.550 ;
        RECT 19.130 13.950 19.430 14.400 ;
        RECT 30.030 13.950 30.330 14.400 ;
        RECT 19.130 13.800 22.980 13.950 ;
        RECT 26.480 13.800 30.330 13.950 ;
        RECT 19.130 13.350 19.430 13.800 ;
        RECT 30.030 13.350 30.330 13.800 ;
        RECT 19.130 13.200 22.980 13.350 ;
        RECT 26.480 13.200 30.330 13.350 ;
        RECT 19.130 12.750 19.430 13.200 ;
        RECT 19.130 12.600 22.980 12.750 ;
        RECT 19.130 12.150 19.430 12.600 ;
        RECT 19.130 12.000 22.980 12.150 ;
        RECT 19.130 11.550 19.430 12.000 ;
        RECT 19.130 11.400 22.980 11.550 ;
        RECT 19.130 10.950 19.430 11.400 ;
        RECT 19.130 10.800 22.980 10.950 ;
        RECT 19.130 10.350 19.430 10.800 ;
        RECT 15.530 1.450 15.680 9.650 ;
        RECT 16.130 1.450 16.280 9.650 ;
        RECT 16.730 1.450 16.880 9.650 ;
        RECT 17.330 1.450 17.480 9.650 ;
        RECT 17.930 1.450 18.080 9.650 ;
        RECT 18.530 1.450 18.680 9.650 ;
        RECT 19.130 9.200 19.430 9.650 ;
        RECT 19.130 9.050 22.980 9.200 ;
        RECT 19.130 8.600 19.430 9.050 ;
        RECT 19.130 8.450 22.980 8.600 ;
        RECT 19.130 8.000 19.430 8.450 ;
        RECT 19.130 7.850 22.980 8.000 ;
        RECT 19.130 7.400 19.430 7.850 ;
        RECT 19.130 7.250 22.980 7.400 ;
        RECT 19.130 6.800 19.430 7.250 ;
        RECT 23.830 6.800 25.630 13.200 ;
        RECT 30.030 12.750 30.330 13.200 ;
        RECT 26.480 12.600 30.330 12.750 ;
        RECT 30.030 12.150 30.330 12.600 ;
        RECT 26.480 12.000 30.330 12.150 ;
        RECT 30.030 11.550 30.330 12.000 ;
        RECT 26.480 11.400 30.330 11.550 ;
        RECT 30.030 10.950 30.330 11.400 ;
        RECT 26.480 10.800 30.330 10.950 ;
        RECT 30.030 10.350 30.330 10.800 ;
        RECT 30.780 10.350 30.930 18.550 ;
        RECT 31.380 10.350 31.530 18.550 ;
        RECT 31.980 10.350 32.130 18.550 ;
        RECT 32.580 10.350 32.730 18.550 ;
        RECT 33.180 10.350 33.330 18.550 ;
        RECT 33.780 10.350 33.930 18.550 ;
        RECT 30.030 9.200 30.330 9.650 ;
        RECT 26.480 9.050 30.330 9.200 ;
        RECT 30.030 8.600 30.330 9.050 ;
        RECT 26.480 8.450 30.330 8.600 ;
        RECT 30.030 8.000 30.330 8.450 ;
        RECT 26.480 7.850 30.330 8.000 ;
        RECT 30.030 7.400 30.330 7.850 ;
        RECT 26.480 7.250 30.330 7.400 ;
        RECT 30.030 6.800 30.330 7.250 ;
        RECT 19.130 6.650 22.980 6.800 ;
        RECT 26.480 6.650 30.330 6.800 ;
        RECT 19.130 6.200 19.430 6.650 ;
        RECT 30.030 6.200 30.330 6.650 ;
        RECT 19.130 6.050 22.980 6.200 ;
        RECT 26.480 6.050 30.330 6.200 ;
        RECT 19.130 5.600 19.430 6.050 ;
        RECT 30.030 5.600 30.330 6.050 ;
        RECT 19.130 5.450 22.980 5.600 ;
        RECT 26.480 5.450 30.330 5.600 ;
        RECT 19.130 5.000 19.430 5.450 ;
        RECT 30.030 5.000 30.330 5.450 ;
        RECT 19.130 4.850 22.980 5.000 ;
        RECT 26.480 4.850 30.330 5.000 ;
        RECT 19.130 4.400 19.430 4.850 ;
        RECT 30.030 4.400 30.330 4.850 ;
        RECT 19.130 4.250 22.980 4.400 ;
        RECT 26.480 4.250 30.330 4.400 ;
        RECT 19.130 3.800 19.430 4.250 ;
        RECT 30.030 3.800 30.330 4.250 ;
        RECT 19.130 3.650 22.980 3.800 ;
        RECT 26.480 3.650 30.330 3.800 ;
        RECT 19.130 3.200 19.430 3.650 ;
        RECT 30.030 3.200 30.330 3.650 ;
        RECT 19.130 3.050 22.980 3.200 ;
        RECT 26.480 3.050 30.330 3.200 ;
        RECT 19.130 2.600 19.430 3.050 ;
        RECT 30.030 2.600 30.330 3.050 ;
        RECT 19.130 2.450 22.980 2.600 ;
        RECT 26.480 2.450 30.330 2.600 ;
        RECT 19.130 2.000 19.430 2.450 ;
        RECT 30.030 2.000 30.330 2.450 ;
        RECT 19.130 1.450 22.930 2.000 ;
        RECT 6.530 1.400 22.930 1.450 ;
        RECT 26.530 1.450 30.330 2.000 ;
        RECT 30.780 1.450 30.930 9.650 ;
        RECT 31.380 1.450 31.530 9.650 ;
        RECT 31.980 1.450 32.130 9.650 ;
        RECT 32.580 1.450 32.730 9.650 ;
        RECT 33.180 1.450 33.330 9.650 ;
        RECT 33.780 1.450 33.930 9.650 ;
        RECT 34.380 1.450 35.080 18.550 ;
        RECT 35.530 10.350 35.680 18.550 ;
        RECT 36.130 10.350 36.280 18.550 ;
        RECT 36.730 10.350 36.880 18.550 ;
        RECT 37.330 10.350 37.480 18.550 ;
        RECT 37.930 10.350 38.080 18.550 ;
        RECT 38.530 10.350 38.680 18.550 ;
        RECT 39.130 18.000 42.930 18.550 ;
        RECT 46.530 18.550 62.930 18.600 ;
        RECT 46.530 18.000 50.330 18.550 ;
        RECT 39.130 17.550 39.430 18.000 ;
        RECT 50.030 17.550 50.330 18.000 ;
        RECT 39.130 17.400 42.980 17.550 ;
        RECT 46.480 17.400 50.330 17.550 ;
        RECT 39.130 16.950 39.430 17.400 ;
        RECT 50.030 16.950 50.330 17.400 ;
        RECT 39.130 16.800 42.980 16.950 ;
        RECT 46.480 16.800 50.330 16.950 ;
        RECT 39.130 16.350 39.430 16.800 ;
        RECT 50.030 16.350 50.330 16.800 ;
        RECT 39.130 16.200 42.980 16.350 ;
        RECT 46.480 16.200 50.330 16.350 ;
        RECT 39.130 15.750 39.430 16.200 ;
        RECT 50.030 15.750 50.330 16.200 ;
        RECT 39.130 15.600 42.980 15.750 ;
        RECT 46.480 15.600 50.330 15.750 ;
        RECT 39.130 15.150 39.430 15.600 ;
        RECT 50.030 15.150 50.330 15.600 ;
        RECT 39.130 15.000 42.980 15.150 ;
        RECT 46.480 15.000 50.330 15.150 ;
        RECT 39.130 14.550 39.430 15.000 ;
        RECT 50.030 14.550 50.330 15.000 ;
        RECT 39.130 14.400 42.980 14.550 ;
        RECT 46.480 14.400 50.330 14.550 ;
        RECT 39.130 13.950 39.430 14.400 ;
        RECT 50.030 13.950 50.330 14.400 ;
        RECT 39.130 13.800 42.980 13.950 ;
        RECT 46.480 13.800 50.330 13.950 ;
        RECT 39.130 13.350 39.430 13.800 ;
        RECT 50.030 13.350 50.330 13.800 ;
        RECT 39.130 13.200 42.980 13.350 ;
        RECT 46.480 13.200 50.330 13.350 ;
        RECT 39.130 12.750 39.430 13.200 ;
        RECT 39.130 12.600 42.980 12.750 ;
        RECT 39.130 12.150 39.430 12.600 ;
        RECT 39.130 12.000 42.980 12.150 ;
        RECT 39.130 11.550 39.430 12.000 ;
        RECT 39.130 11.400 42.980 11.550 ;
        RECT 39.130 10.950 39.430 11.400 ;
        RECT 39.130 10.800 42.980 10.950 ;
        RECT 39.130 10.350 39.430 10.800 ;
        RECT 35.530 1.450 35.680 9.650 ;
        RECT 36.130 1.450 36.280 9.650 ;
        RECT 36.730 1.450 36.880 9.650 ;
        RECT 37.330 1.450 37.480 9.650 ;
        RECT 37.930 1.450 38.080 9.650 ;
        RECT 38.530 1.450 38.680 9.650 ;
        RECT 39.130 9.200 39.430 9.650 ;
        RECT 39.130 9.050 42.980 9.200 ;
        RECT 39.130 8.600 39.430 9.050 ;
        RECT 39.130 8.450 42.980 8.600 ;
        RECT 39.130 8.000 39.430 8.450 ;
        RECT 39.130 7.850 42.980 8.000 ;
        RECT 39.130 7.400 39.430 7.850 ;
        RECT 39.130 7.250 42.980 7.400 ;
        RECT 39.130 6.800 39.430 7.250 ;
        RECT 43.830 6.800 45.630 13.200 ;
        RECT 50.030 12.750 50.330 13.200 ;
        RECT 46.480 12.600 50.330 12.750 ;
        RECT 50.030 12.150 50.330 12.600 ;
        RECT 46.480 12.000 50.330 12.150 ;
        RECT 50.030 11.550 50.330 12.000 ;
        RECT 46.480 11.400 50.330 11.550 ;
        RECT 50.030 10.950 50.330 11.400 ;
        RECT 46.480 10.800 50.330 10.950 ;
        RECT 50.030 10.350 50.330 10.800 ;
        RECT 50.780 10.350 50.930 18.550 ;
        RECT 51.380 10.350 51.530 18.550 ;
        RECT 51.980 10.350 52.130 18.550 ;
        RECT 52.580 10.350 52.730 18.550 ;
        RECT 53.180 10.350 53.330 18.550 ;
        RECT 53.780 10.350 53.930 18.550 ;
        RECT 50.030 9.200 50.330 9.650 ;
        RECT 46.480 9.050 50.330 9.200 ;
        RECT 50.030 8.600 50.330 9.050 ;
        RECT 46.480 8.450 50.330 8.600 ;
        RECT 50.030 8.000 50.330 8.450 ;
        RECT 46.480 7.850 50.330 8.000 ;
        RECT 50.030 7.400 50.330 7.850 ;
        RECT 46.480 7.250 50.330 7.400 ;
        RECT 50.030 6.800 50.330 7.250 ;
        RECT 39.130 6.650 42.980 6.800 ;
        RECT 46.480 6.650 50.330 6.800 ;
        RECT 39.130 6.200 39.430 6.650 ;
        RECT 50.030 6.200 50.330 6.650 ;
        RECT 39.130 6.050 42.980 6.200 ;
        RECT 46.480 6.050 50.330 6.200 ;
        RECT 39.130 5.600 39.430 6.050 ;
        RECT 50.030 5.600 50.330 6.050 ;
        RECT 39.130 5.450 42.980 5.600 ;
        RECT 46.480 5.450 50.330 5.600 ;
        RECT 39.130 5.000 39.430 5.450 ;
        RECT 50.030 5.000 50.330 5.450 ;
        RECT 39.130 4.850 42.980 5.000 ;
        RECT 46.480 4.850 50.330 5.000 ;
        RECT 39.130 4.400 39.430 4.850 ;
        RECT 50.030 4.400 50.330 4.850 ;
        RECT 39.130 4.250 42.980 4.400 ;
        RECT 46.480 4.250 50.330 4.400 ;
        RECT 39.130 3.800 39.430 4.250 ;
        RECT 50.030 3.800 50.330 4.250 ;
        RECT 39.130 3.650 42.980 3.800 ;
        RECT 46.480 3.650 50.330 3.800 ;
        RECT 39.130 3.200 39.430 3.650 ;
        RECT 50.030 3.200 50.330 3.650 ;
        RECT 39.130 3.050 42.980 3.200 ;
        RECT 46.480 3.050 50.330 3.200 ;
        RECT 39.130 2.600 39.430 3.050 ;
        RECT 50.030 2.600 50.330 3.050 ;
        RECT 39.130 2.450 42.980 2.600 ;
        RECT 46.480 2.450 50.330 2.600 ;
        RECT 39.130 2.000 39.430 2.450 ;
        RECT 50.030 2.000 50.330 2.450 ;
        RECT 39.130 1.450 42.930 2.000 ;
        RECT 26.530 1.400 42.930 1.450 ;
        RECT 46.530 1.450 50.330 2.000 ;
        RECT 50.780 1.450 50.930 9.650 ;
        RECT 51.380 1.450 51.530 9.650 ;
        RECT 51.980 1.450 52.130 9.650 ;
        RECT 52.580 1.450 52.730 9.650 ;
        RECT 53.180 1.450 53.330 9.650 ;
        RECT 53.780 1.450 53.930 9.650 ;
        RECT 54.380 1.450 55.080 18.550 ;
        RECT 55.530 10.350 55.680 18.550 ;
        RECT 56.130 10.350 56.280 18.550 ;
        RECT 56.730 10.350 56.880 18.550 ;
        RECT 57.330 10.350 57.480 18.550 ;
        RECT 57.930 10.350 58.080 18.550 ;
        RECT 58.530 10.350 58.680 18.550 ;
        RECT 59.130 18.000 62.930 18.550 ;
        RECT 66.530 18.550 82.930 18.600 ;
        RECT 66.530 18.000 70.330 18.550 ;
        RECT 59.130 17.550 59.430 18.000 ;
        RECT 70.030 17.550 70.330 18.000 ;
        RECT 59.130 17.400 62.980 17.550 ;
        RECT 66.480 17.400 70.330 17.550 ;
        RECT 59.130 16.950 59.430 17.400 ;
        RECT 70.030 16.950 70.330 17.400 ;
        RECT 59.130 16.800 62.980 16.950 ;
        RECT 66.480 16.800 70.330 16.950 ;
        RECT 59.130 16.350 59.430 16.800 ;
        RECT 70.030 16.350 70.330 16.800 ;
        RECT 59.130 16.200 62.980 16.350 ;
        RECT 66.480 16.200 70.330 16.350 ;
        RECT 59.130 15.750 59.430 16.200 ;
        RECT 70.030 15.750 70.330 16.200 ;
        RECT 59.130 15.600 62.980 15.750 ;
        RECT 66.480 15.600 70.330 15.750 ;
        RECT 59.130 15.150 59.430 15.600 ;
        RECT 70.030 15.150 70.330 15.600 ;
        RECT 59.130 15.000 62.980 15.150 ;
        RECT 66.480 15.000 70.330 15.150 ;
        RECT 59.130 14.550 59.430 15.000 ;
        RECT 70.030 14.550 70.330 15.000 ;
        RECT 59.130 14.400 62.980 14.550 ;
        RECT 66.480 14.400 70.330 14.550 ;
        RECT 59.130 13.950 59.430 14.400 ;
        RECT 70.030 13.950 70.330 14.400 ;
        RECT 59.130 13.800 62.980 13.950 ;
        RECT 66.480 13.800 70.330 13.950 ;
        RECT 59.130 13.350 59.430 13.800 ;
        RECT 70.030 13.350 70.330 13.800 ;
        RECT 59.130 13.200 62.980 13.350 ;
        RECT 66.480 13.200 70.330 13.350 ;
        RECT 59.130 12.750 59.430 13.200 ;
        RECT 59.130 12.600 62.980 12.750 ;
        RECT 59.130 12.150 59.430 12.600 ;
        RECT 59.130 12.000 62.980 12.150 ;
        RECT 59.130 11.550 59.430 12.000 ;
        RECT 59.130 11.400 62.980 11.550 ;
        RECT 59.130 10.950 59.430 11.400 ;
        RECT 59.130 10.800 62.980 10.950 ;
        RECT 59.130 10.350 59.430 10.800 ;
        RECT 55.530 1.450 55.680 9.650 ;
        RECT 56.130 1.450 56.280 9.650 ;
        RECT 56.730 1.450 56.880 9.650 ;
        RECT 57.330 1.450 57.480 9.650 ;
        RECT 57.930 1.450 58.080 9.650 ;
        RECT 58.530 1.450 58.680 9.650 ;
        RECT 59.130 9.200 59.430 9.650 ;
        RECT 59.130 9.050 62.980 9.200 ;
        RECT 59.130 8.600 59.430 9.050 ;
        RECT 59.130 8.450 62.980 8.600 ;
        RECT 59.130 8.000 59.430 8.450 ;
        RECT 59.130 7.850 62.980 8.000 ;
        RECT 59.130 7.400 59.430 7.850 ;
        RECT 59.130 7.250 62.980 7.400 ;
        RECT 59.130 6.800 59.430 7.250 ;
        RECT 63.830 6.800 65.630 13.200 ;
        RECT 70.030 12.750 70.330 13.200 ;
        RECT 66.480 12.600 70.330 12.750 ;
        RECT 70.030 12.150 70.330 12.600 ;
        RECT 66.480 12.000 70.330 12.150 ;
        RECT 70.030 11.550 70.330 12.000 ;
        RECT 66.480 11.400 70.330 11.550 ;
        RECT 70.030 10.950 70.330 11.400 ;
        RECT 66.480 10.800 70.330 10.950 ;
        RECT 70.030 10.350 70.330 10.800 ;
        RECT 70.780 10.350 70.930 18.550 ;
        RECT 71.380 10.350 71.530 18.550 ;
        RECT 71.980 10.350 72.130 18.550 ;
        RECT 72.580 10.350 72.730 18.550 ;
        RECT 73.180 10.350 73.330 18.550 ;
        RECT 73.780 10.350 73.930 18.550 ;
        RECT 70.030 9.200 70.330 9.650 ;
        RECT 66.480 9.050 70.330 9.200 ;
        RECT 70.030 8.600 70.330 9.050 ;
        RECT 66.480 8.450 70.330 8.600 ;
        RECT 70.030 8.000 70.330 8.450 ;
        RECT 66.480 7.850 70.330 8.000 ;
        RECT 70.030 7.400 70.330 7.850 ;
        RECT 66.480 7.250 70.330 7.400 ;
        RECT 70.030 6.800 70.330 7.250 ;
        RECT 59.130 6.650 62.980 6.800 ;
        RECT 66.480 6.650 70.330 6.800 ;
        RECT 59.130 6.200 59.430 6.650 ;
        RECT 70.030 6.200 70.330 6.650 ;
        RECT 59.130 6.050 62.980 6.200 ;
        RECT 66.480 6.050 70.330 6.200 ;
        RECT 59.130 5.600 59.430 6.050 ;
        RECT 70.030 5.600 70.330 6.050 ;
        RECT 59.130 5.450 62.980 5.600 ;
        RECT 66.480 5.450 70.330 5.600 ;
        RECT 59.130 5.000 59.430 5.450 ;
        RECT 70.030 5.000 70.330 5.450 ;
        RECT 59.130 4.850 62.980 5.000 ;
        RECT 66.480 4.850 70.330 5.000 ;
        RECT 59.130 4.400 59.430 4.850 ;
        RECT 70.030 4.400 70.330 4.850 ;
        RECT 59.130 4.250 62.980 4.400 ;
        RECT 66.480 4.250 70.330 4.400 ;
        RECT 59.130 3.800 59.430 4.250 ;
        RECT 70.030 3.800 70.330 4.250 ;
        RECT 59.130 3.650 62.980 3.800 ;
        RECT 66.480 3.650 70.330 3.800 ;
        RECT 59.130 3.200 59.430 3.650 ;
        RECT 70.030 3.200 70.330 3.650 ;
        RECT 59.130 3.050 62.980 3.200 ;
        RECT 66.480 3.050 70.330 3.200 ;
        RECT 59.130 2.600 59.430 3.050 ;
        RECT 70.030 2.600 70.330 3.050 ;
        RECT 59.130 2.450 62.980 2.600 ;
        RECT 66.480 2.450 70.330 2.600 ;
        RECT 59.130 2.000 59.430 2.450 ;
        RECT 70.030 2.000 70.330 2.450 ;
        RECT 59.130 1.450 62.930 2.000 ;
        RECT 46.530 1.400 62.930 1.450 ;
        RECT 66.530 1.450 70.330 2.000 ;
        RECT 70.780 1.450 70.930 9.650 ;
        RECT 71.380 1.450 71.530 9.650 ;
        RECT 71.980 1.450 72.130 9.650 ;
        RECT 72.580 1.450 72.730 9.650 ;
        RECT 73.180 1.450 73.330 9.650 ;
        RECT 73.780 1.450 73.930 9.650 ;
        RECT 74.380 1.450 75.080 18.550 ;
        RECT 75.530 10.350 75.680 18.550 ;
        RECT 76.130 10.350 76.280 18.550 ;
        RECT 76.730 10.350 76.880 18.550 ;
        RECT 77.330 10.350 77.480 18.550 ;
        RECT 77.930 10.350 78.080 18.550 ;
        RECT 78.530 10.350 78.680 18.550 ;
        RECT 79.130 18.000 82.930 18.550 ;
        RECT 86.530 18.550 102.930 18.600 ;
        RECT 86.530 18.000 90.330 18.550 ;
        RECT 79.130 17.550 79.430 18.000 ;
        RECT 90.030 17.550 90.330 18.000 ;
        RECT 79.130 17.400 82.980 17.550 ;
        RECT 86.480 17.400 90.330 17.550 ;
        RECT 79.130 16.950 79.430 17.400 ;
        RECT 90.030 16.950 90.330 17.400 ;
        RECT 79.130 16.800 82.980 16.950 ;
        RECT 86.480 16.800 90.330 16.950 ;
        RECT 79.130 16.350 79.430 16.800 ;
        RECT 90.030 16.350 90.330 16.800 ;
        RECT 79.130 16.200 82.980 16.350 ;
        RECT 86.480 16.200 90.330 16.350 ;
        RECT 79.130 15.750 79.430 16.200 ;
        RECT 90.030 15.750 90.330 16.200 ;
        RECT 79.130 15.600 82.980 15.750 ;
        RECT 86.480 15.600 90.330 15.750 ;
        RECT 79.130 15.150 79.430 15.600 ;
        RECT 90.030 15.150 90.330 15.600 ;
        RECT 79.130 15.000 82.980 15.150 ;
        RECT 86.480 15.000 90.330 15.150 ;
        RECT 79.130 14.550 79.430 15.000 ;
        RECT 90.030 14.550 90.330 15.000 ;
        RECT 79.130 14.400 82.980 14.550 ;
        RECT 86.480 14.400 90.330 14.550 ;
        RECT 79.130 13.950 79.430 14.400 ;
        RECT 90.030 13.950 90.330 14.400 ;
        RECT 79.130 13.800 82.980 13.950 ;
        RECT 86.480 13.800 90.330 13.950 ;
        RECT 79.130 13.350 79.430 13.800 ;
        RECT 90.030 13.350 90.330 13.800 ;
        RECT 79.130 13.200 82.980 13.350 ;
        RECT 86.480 13.200 90.330 13.350 ;
        RECT 79.130 12.750 79.430 13.200 ;
        RECT 79.130 12.600 82.980 12.750 ;
        RECT 79.130 12.150 79.430 12.600 ;
        RECT 79.130 12.000 82.980 12.150 ;
        RECT 79.130 11.550 79.430 12.000 ;
        RECT 79.130 11.400 82.980 11.550 ;
        RECT 79.130 10.950 79.430 11.400 ;
        RECT 79.130 10.800 82.980 10.950 ;
        RECT 79.130 10.350 79.430 10.800 ;
        RECT 75.530 1.450 75.680 9.650 ;
        RECT 76.130 1.450 76.280 9.650 ;
        RECT 76.730 1.450 76.880 9.650 ;
        RECT 77.330 1.450 77.480 9.650 ;
        RECT 77.930 1.450 78.080 9.650 ;
        RECT 78.530 1.450 78.680 9.650 ;
        RECT 79.130 9.200 79.430 9.650 ;
        RECT 79.130 9.050 82.980 9.200 ;
        RECT 79.130 8.600 79.430 9.050 ;
        RECT 79.130 8.450 82.980 8.600 ;
        RECT 79.130 8.000 79.430 8.450 ;
        RECT 79.130 7.850 82.980 8.000 ;
        RECT 79.130 7.400 79.430 7.850 ;
        RECT 79.130 7.250 82.980 7.400 ;
        RECT 79.130 6.800 79.430 7.250 ;
        RECT 83.830 6.800 85.630 13.200 ;
        RECT 90.030 12.750 90.330 13.200 ;
        RECT 86.480 12.600 90.330 12.750 ;
        RECT 90.030 12.150 90.330 12.600 ;
        RECT 86.480 12.000 90.330 12.150 ;
        RECT 90.030 11.550 90.330 12.000 ;
        RECT 86.480 11.400 90.330 11.550 ;
        RECT 90.030 10.950 90.330 11.400 ;
        RECT 86.480 10.800 90.330 10.950 ;
        RECT 90.030 10.350 90.330 10.800 ;
        RECT 90.780 10.350 90.930 18.550 ;
        RECT 91.380 10.350 91.530 18.550 ;
        RECT 91.980 10.350 92.130 18.550 ;
        RECT 92.580 10.350 92.730 18.550 ;
        RECT 93.180 10.350 93.330 18.550 ;
        RECT 93.780 10.350 93.930 18.550 ;
        RECT 90.030 9.200 90.330 9.650 ;
        RECT 86.480 9.050 90.330 9.200 ;
        RECT 90.030 8.600 90.330 9.050 ;
        RECT 86.480 8.450 90.330 8.600 ;
        RECT 90.030 8.000 90.330 8.450 ;
        RECT 86.480 7.850 90.330 8.000 ;
        RECT 90.030 7.400 90.330 7.850 ;
        RECT 86.480 7.250 90.330 7.400 ;
        RECT 90.030 6.800 90.330 7.250 ;
        RECT 79.130 6.650 82.980 6.800 ;
        RECT 86.480 6.650 90.330 6.800 ;
        RECT 79.130 6.200 79.430 6.650 ;
        RECT 90.030 6.200 90.330 6.650 ;
        RECT 79.130 6.050 82.980 6.200 ;
        RECT 86.480 6.050 90.330 6.200 ;
        RECT 79.130 5.600 79.430 6.050 ;
        RECT 90.030 5.600 90.330 6.050 ;
        RECT 79.130 5.450 82.980 5.600 ;
        RECT 86.480 5.450 90.330 5.600 ;
        RECT 79.130 5.000 79.430 5.450 ;
        RECT 90.030 5.000 90.330 5.450 ;
        RECT 79.130 4.850 82.980 5.000 ;
        RECT 86.480 4.850 90.330 5.000 ;
        RECT 79.130 4.400 79.430 4.850 ;
        RECT 90.030 4.400 90.330 4.850 ;
        RECT 79.130 4.250 82.980 4.400 ;
        RECT 86.480 4.250 90.330 4.400 ;
        RECT 79.130 3.800 79.430 4.250 ;
        RECT 90.030 3.800 90.330 4.250 ;
        RECT 79.130 3.650 82.980 3.800 ;
        RECT 86.480 3.650 90.330 3.800 ;
        RECT 79.130 3.200 79.430 3.650 ;
        RECT 90.030 3.200 90.330 3.650 ;
        RECT 79.130 3.050 82.980 3.200 ;
        RECT 86.480 3.050 90.330 3.200 ;
        RECT 79.130 2.600 79.430 3.050 ;
        RECT 90.030 2.600 90.330 3.050 ;
        RECT 79.130 2.450 82.980 2.600 ;
        RECT 86.480 2.450 90.330 2.600 ;
        RECT 79.130 2.000 79.430 2.450 ;
        RECT 90.030 2.000 90.330 2.450 ;
        RECT 79.130 1.450 82.930 2.000 ;
        RECT 66.530 1.400 82.930 1.450 ;
        RECT 86.530 1.450 90.330 2.000 ;
        RECT 90.780 1.450 90.930 9.650 ;
        RECT 91.380 1.450 91.530 9.650 ;
        RECT 91.980 1.450 92.130 9.650 ;
        RECT 92.580 1.450 92.730 9.650 ;
        RECT 93.180 1.450 93.330 9.650 ;
        RECT 93.780 1.450 93.930 9.650 ;
        RECT 94.380 1.450 95.080 18.550 ;
        RECT 95.530 10.350 95.680 18.550 ;
        RECT 96.130 10.350 96.280 18.550 ;
        RECT 96.730 10.350 96.880 18.550 ;
        RECT 97.330 10.350 97.480 18.550 ;
        RECT 97.930 10.350 98.080 18.550 ;
        RECT 98.530 10.350 98.680 18.550 ;
        RECT 99.130 18.000 102.930 18.550 ;
        RECT 99.130 17.550 99.430 18.000 ;
        RECT 99.130 17.400 102.980 17.550 ;
        RECT 99.130 16.950 99.430 17.400 ;
        RECT 99.130 16.800 102.980 16.950 ;
        RECT 99.130 16.350 99.430 16.800 ;
        RECT 99.130 16.200 102.980 16.350 ;
        RECT 99.130 15.750 99.430 16.200 ;
        RECT 99.130 15.600 102.980 15.750 ;
        RECT 99.130 15.150 99.430 15.600 ;
        RECT 99.130 15.000 102.980 15.150 ;
        RECT 99.130 14.550 99.430 15.000 ;
        RECT 99.130 14.400 102.980 14.550 ;
        RECT 99.130 13.950 99.430 14.400 ;
        RECT 99.130 13.800 102.980 13.950 ;
        RECT 99.130 13.350 99.430 13.800 ;
        RECT 99.130 13.200 102.980 13.350 ;
        RECT 99.130 12.750 99.430 13.200 ;
        RECT 99.130 12.600 102.980 12.750 ;
        RECT 99.130 12.150 99.430 12.600 ;
        RECT 99.130 12.000 102.980 12.150 ;
        RECT 99.130 11.550 99.430 12.000 ;
        RECT 99.130 11.400 102.980 11.550 ;
        RECT 99.130 10.950 99.430 11.400 ;
        RECT 99.130 10.800 102.980 10.950 ;
        RECT 99.130 10.350 99.430 10.800 ;
        RECT 95.530 1.450 95.680 9.650 ;
        RECT 96.130 1.450 96.280 9.650 ;
        RECT 96.730 1.450 96.880 9.650 ;
        RECT 97.330 1.450 97.480 9.650 ;
        RECT 97.930 1.450 98.080 9.650 ;
        RECT 98.530 1.450 98.680 9.650 ;
        RECT 99.130 9.200 99.430 9.650 ;
        RECT 99.130 9.050 102.980 9.200 ;
        RECT 99.130 8.600 99.430 9.050 ;
        RECT 99.130 8.450 102.980 8.600 ;
        RECT 99.130 8.000 99.430 8.450 ;
        RECT 99.130 7.850 102.980 8.000 ;
        RECT 99.130 7.400 99.430 7.850 ;
        RECT 99.130 7.250 102.980 7.400 ;
        RECT 99.130 6.800 99.430 7.250 ;
        RECT 103.830 6.800 104.730 13.200 ;
        RECT 109.850 10.250 111.850 11.525 ;
        RECT 99.130 6.650 102.980 6.800 ;
        RECT 99.130 6.200 99.430 6.650 ;
        RECT 99.130 6.050 102.980 6.200 ;
        RECT 99.130 5.600 99.430 6.050 ;
        RECT 99.130 5.450 102.980 5.600 ;
        RECT 99.130 5.000 99.430 5.450 ;
        RECT 99.130 4.850 102.980 5.000 ;
        RECT 99.130 4.400 99.430 4.850 ;
        RECT 99.130 4.250 102.980 4.400 ;
        RECT 99.130 3.800 99.430 4.250 ;
        RECT 99.130 3.650 102.980 3.800 ;
        RECT 99.130 3.200 99.430 3.650 ;
        RECT 99.130 3.050 102.980 3.200 ;
        RECT 99.130 2.600 99.430 3.050 ;
        RECT 99.130 2.450 102.980 2.600 ;
        RECT 99.130 2.000 99.430 2.450 ;
        RECT 99.130 1.450 102.930 2.000 ;
        RECT 86.530 1.400 102.930 1.450 ;
        RECT 9.630 0.900 19.830 1.400 ;
        RECT 29.630 0.900 39.830 1.400 ;
        RECT 49.630 0.900 59.830 1.400 ;
        RECT 69.630 0.900 79.830 1.400 ;
        RECT 89.630 0.900 99.830 1.400 ;
        RECT 11.530 0.000 17.930 0.900 ;
        RECT 31.530 0.000 37.930 0.900 ;
        RECT 51.530 0.000 57.930 0.900 ;
        RECT 71.530 0.000 77.930 0.900 ;
        RECT 91.530 0.000 97.930 0.900 ;
      LAYER via2 ;
        RECT 110.050 369.975 110.410 370.355 ;
        RECT 110.680 369.975 111.040 370.355 ;
        RECT 111.280 369.975 111.640 370.355 ;
        RECT 110.050 369.385 110.410 369.765 ;
        RECT 110.680 369.385 111.040 369.765 ;
        RECT 111.280 369.385 111.640 369.765 ;
        RECT 110.050 349.975 110.410 350.355 ;
        RECT 110.680 349.975 111.040 350.355 ;
        RECT 111.280 349.975 111.640 350.355 ;
        RECT 110.050 349.385 110.410 349.765 ;
        RECT 110.680 349.385 111.040 349.765 ;
        RECT 111.280 349.385 111.640 349.765 ;
        RECT 110.050 329.910 110.410 330.290 ;
        RECT 110.680 329.910 111.040 330.290 ;
        RECT 111.280 329.910 111.640 330.290 ;
        RECT 110.050 329.320 110.410 329.700 ;
        RECT 110.680 329.320 111.040 329.700 ;
        RECT 111.280 329.320 111.640 329.700 ;
        RECT 110.050 309.905 110.410 310.285 ;
        RECT 110.680 309.905 111.040 310.285 ;
        RECT 111.280 309.905 111.640 310.285 ;
        RECT 110.050 309.315 110.410 309.695 ;
        RECT 110.680 309.315 111.040 309.695 ;
        RECT 111.280 309.315 111.640 309.695 ;
        RECT 110.050 290.100 110.410 290.480 ;
        RECT 110.680 290.100 111.040 290.480 ;
        RECT 111.280 290.100 111.640 290.480 ;
        RECT 110.050 289.510 110.410 289.890 ;
        RECT 110.680 289.510 111.040 289.890 ;
        RECT 111.280 289.510 111.640 289.890 ;
        RECT 110.050 270.015 110.410 270.395 ;
        RECT 110.680 270.015 111.040 270.395 ;
        RECT 111.280 270.015 111.640 270.395 ;
        RECT 110.050 269.425 110.410 269.805 ;
        RECT 110.680 269.425 111.040 269.805 ;
        RECT 111.280 269.425 111.640 269.805 ;
        RECT 110.050 250.410 110.410 250.790 ;
        RECT 110.680 250.410 111.040 250.790 ;
        RECT 111.280 250.410 111.640 250.790 ;
        RECT 110.050 249.820 110.410 250.200 ;
        RECT 110.680 249.820 111.040 250.200 ;
        RECT 111.280 249.820 111.640 250.200 ;
        RECT 110.050 229.120 110.410 229.500 ;
        RECT 110.680 229.120 111.040 229.500 ;
        RECT 111.280 229.120 111.640 229.500 ;
        RECT 110.050 228.530 110.410 228.910 ;
        RECT 110.680 228.530 111.040 228.910 ;
        RECT 111.280 228.530 111.640 228.910 ;
        RECT 110.030 217.570 111.490 219.190 ;
        RECT 110.030 183.150 111.490 184.770 ;
        RECT 110.050 150.270 110.410 150.650 ;
        RECT 110.680 150.270 111.040 150.650 ;
        RECT 111.280 150.270 111.640 150.650 ;
        RECT 110.050 149.680 110.410 150.060 ;
        RECT 110.680 149.680 111.040 150.060 ;
        RECT 111.280 149.680 111.640 150.060 ;
        RECT 110.050 129.475 110.410 129.855 ;
        RECT 110.680 129.475 111.040 129.855 ;
        RECT 111.280 129.475 111.640 129.855 ;
        RECT 110.050 128.885 110.410 129.265 ;
        RECT 110.680 128.885 111.040 129.265 ;
        RECT 111.280 128.885 111.640 129.265 ;
        RECT 110.050 110.525 110.410 110.905 ;
        RECT 110.680 110.525 111.040 110.905 ;
        RECT 111.280 110.525 111.640 110.905 ;
        RECT 110.050 109.935 110.410 110.315 ;
        RECT 110.680 109.935 111.040 110.315 ;
        RECT 111.280 109.935 111.640 110.315 ;
        RECT 110.050 89.990 110.410 90.370 ;
        RECT 110.680 89.990 111.040 90.370 ;
        RECT 111.280 89.990 111.640 90.370 ;
        RECT 110.050 89.400 110.410 89.780 ;
        RECT 110.680 89.400 111.040 89.780 ;
        RECT 111.280 89.400 111.640 89.780 ;
        RECT 110.050 70.900 110.410 71.280 ;
        RECT 110.680 70.900 111.040 71.280 ;
        RECT 111.280 70.900 111.640 71.280 ;
        RECT 110.050 70.310 110.410 70.690 ;
        RECT 110.680 70.310 111.040 70.690 ;
        RECT 111.280 70.310 111.640 70.690 ;
        RECT 110.050 51.080 110.410 51.460 ;
        RECT 110.680 51.080 111.040 51.460 ;
        RECT 111.280 51.080 111.640 51.460 ;
        RECT 110.050 50.490 110.410 50.870 ;
        RECT 110.680 50.490 111.040 50.870 ;
        RECT 111.280 50.490 111.640 50.870 ;
        RECT 110.050 31.020 110.410 31.400 ;
        RECT 110.680 31.020 111.040 31.400 ;
        RECT 111.280 31.020 111.640 31.400 ;
        RECT 110.050 30.430 110.410 30.810 ;
        RECT 110.680 30.430 111.040 30.810 ;
        RECT 111.280 30.430 111.640 30.810 ;
        RECT 110.050 11.020 110.410 11.400 ;
        RECT 110.680 11.020 111.040 11.400 ;
        RECT 111.280 11.020 111.640 11.400 ;
        RECT 110.050 10.430 110.410 10.810 ;
        RECT 110.680 10.430 111.040 10.810 ;
        RECT 111.280 10.430 111.640 10.810 ;
      LAYER met3 ;
        RECT 109.850 369.205 111.850 370.480 ;
        RECT 109.850 349.205 111.850 350.480 ;
        RECT 109.850 329.140 111.850 330.415 ;
        RECT 109.850 309.135 111.850 310.410 ;
        RECT 109.850 289.330 111.850 290.605 ;
        RECT 109.850 269.245 111.850 270.520 ;
        RECT 109.850 249.640 111.850 250.915 ;
        RECT 109.850 228.350 111.850 229.625 ;
        RECT 109.850 217.400 111.850 219.350 ;
        RECT 109.850 182.980 111.850 184.930 ;
        RECT 109.850 149.500 111.850 150.775 ;
        RECT 109.850 128.705 111.850 129.980 ;
        RECT 109.850 109.755 111.850 111.030 ;
        RECT 109.850 89.220 111.850 90.495 ;
        RECT 109.850 70.130 111.850 71.405 ;
        RECT 109.850 50.310 111.850 51.585 ;
        RECT 109.850 30.250 111.850 31.525 ;
        RECT 109.850 10.250 111.850 11.525 ;
      LAYER via3 ;
        RECT 110.050 369.975 110.410 370.355 ;
        RECT 110.680 369.975 111.040 370.355 ;
        RECT 111.280 369.975 111.640 370.355 ;
        RECT 110.050 369.385 110.410 369.765 ;
        RECT 110.680 369.385 111.040 369.765 ;
        RECT 111.280 369.385 111.640 369.765 ;
        RECT 110.050 349.975 110.410 350.355 ;
        RECT 110.680 349.975 111.040 350.355 ;
        RECT 111.280 349.975 111.640 350.355 ;
        RECT 110.050 349.385 110.410 349.765 ;
        RECT 110.680 349.385 111.040 349.765 ;
        RECT 111.280 349.385 111.640 349.765 ;
        RECT 110.050 329.910 110.410 330.290 ;
        RECT 110.680 329.910 111.040 330.290 ;
        RECT 111.280 329.910 111.640 330.290 ;
        RECT 110.050 329.320 110.410 329.700 ;
        RECT 110.680 329.320 111.040 329.700 ;
        RECT 111.280 329.320 111.640 329.700 ;
        RECT 110.050 309.905 110.410 310.285 ;
        RECT 110.680 309.905 111.040 310.285 ;
        RECT 111.280 309.905 111.640 310.285 ;
        RECT 110.050 309.315 110.410 309.695 ;
        RECT 110.680 309.315 111.040 309.695 ;
        RECT 111.280 309.315 111.640 309.695 ;
        RECT 110.050 290.100 110.410 290.480 ;
        RECT 110.680 290.100 111.040 290.480 ;
        RECT 111.280 290.100 111.640 290.480 ;
        RECT 110.050 289.510 110.410 289.890 ;
        RECT 110.680 289.510 111.040 289.890 ;
        RECT 111.280 289.510 111.640 289.890 ;
        RECT 110.050 270.015 110.410 270.395 ;
        RECT 110.680 270.015 111.040 270.395 ;
        RECT 111.280 270.015 111.640 270.395 ;
        RECT 110.050 269.425 110.410 269.805 ;
        RECT 110.680 269.425 111.040 269.805 ;
        RECT 111.280 269.425 111.640 269.805 ;
        RECT 110.050 250.410 110.410 250.790 ;
        RECT 110.680 250.410 111.040 250.790 ;
        RECT 111.280 250.410 111.640 250.790 ;
        RECT 110.050 249.820 110.410 250.200 ;
        RECT 110.680 249.820 111.040 250.200 ;
        RECT 111.280 249.820 111.640 250.200 ;
        RECT 110.050 229.120 110.410 229.500 ;
        RECT 110.680 229.120 111.040 229.500 ;
        RECT 111.280 229.120 111.640 229.500 ;
        RECT 110.050 228.530 110.410 228.910 ;
        RECT 110.680 228.530 111.040 228.910 ;
        RECT 111.280 228.530 111.640 228.910 ;
        RECT 110.030 217.570 111.490 219.190 ;
        RECT 110.030 183.150 111.490 184.770 ;
        RECT 110.050 150.270 110.410 150.650 ;
        RECT 110.680 150.270 111.040 150.650 ;
        RECT 111.280 150.270 111.640 150.650 ;
        RECT 110.050 149.680 110.410 150.060 ;
        RECT 110.680 149.680 111.040 150.060 ;
        RECT 111.280 149.680 111.640 150.060 ;
        RECT 110.050 129.475 110.410 129.855 ;
        RECT 110.680 129.475 111.040 129.855 ;
        RECT 111.280 129.475 111.640 129.855 ;
        RECT 110.050 128.885 110.410 129.265 ;
        RECT 110.680 128.885 111.040 129.265 ;
        RECT 111.280 128.885 111.640 129.265 ;
        RECT 110.050 110.525 110.410 110.905 ;
        RECT 110.680 110.525 111.040 110.905 ;
        RECT 111.280 110.525 111.640 110.905 ;
        RECT 110.050 109.935 110.410 110.315 ;
        RECT 110.680 109.935 111.040 110.315 ;
        RECT 111.280 109.935 111.640 110.315 ;
        RECT 110.050 89.990 110.410 90.370 ;
        RECT 110.680 89.990 111.040 90.370 ;
        RECT 111.280 89.990 111.640 90.370 ;
        RECT 110.050 89.400 110.410 89.780 ;
        RECT 110.680 89.400 111.040 89.780 ;
        RECT 111.280 89.400 111.640 89.780 ;
        RECT 110.050 70.900 110.410 71.280 ;
        RECT 110.680 70.900 111.040 71.280 ;
        RECT 111.280 70.900 111.640 71.280 ;
        RECT 110.050 70.310 110.410 70.690 ;
        RECT 110.680 70.310 111.040 70.690 ;
        RECT 111.280 70.310 111.640 70.690 ;
        RECT 110.050 51.080 110.410 51.460 ;
        RECT 110.680 51.080 111.040 51.460 ;
        RECT 111.280 51.080 111.640 51.460 ;
        RECT 110.050 50.490 110.410 50.870 ;
        RECT 110.680 50.490 111.040 50.870 ;
        RECT 111.280 50.490 111.640 50.870 ;
        RECT 110.050 31.020 110.410 31.400 ;
        RECT 110.680 31.020 111.040 31.400 ;
        RECT 111.280 31.020 111.640 31.400 ;
        RECT 110.050 30.430 110.410 30.810 ;
        RECT 110.680 30.430 111.040 30.810 ;
        RECT 111.280 30.430 111.640 30.810 ;
        RECT 110.050 11.020 110.410 11.400 ;
        RECT 110.680 11.020 111.040 11.400 ;
        RECT 111.280 11.020 111.640 11.400 ;
        RECT 110.050 10.430 110.410 10.810 ;
        RECT 110.680 10.430 111.040 10.810 ;
        RECT 111.280 10.430 111.640 10.810 ;
      LAYER met4 ;
        RECT 109.850 0.000 111.850 380.000 ;
    END
  END vcm
  OBS
      LAYER pwell ;
        RECT 17.765 195.350 17.935 195.540 ;
        RECT 20.525 195.350 20.695 195.540 ;
        RECT 21.910 195.370 22.080 195.540 ;
        RECT 23.290 195.370 23.460 195.540 ;
        RECT 21.910 195.350 22.015 195.370 ;
        RECT 23.290 195.350 23.395 195.370 ;
        RECT 15.470 194.440 18.080 195.350 ;
        RECT 18.230 194.440 20.840 195.350 ;
        RECT 21.085 194.440 22.015 195.350 ;
        RECT 22.465 194.440 23.395 195.350 ;
        RECT 8.430 190.120 9.780 191.030 ;
        RECT 10.475 190.800 14.225 191.030 ;
        RECT 15.075 190.800 18.825 191.030 ;
        RECT 19.675 190.800 23.425 191.030 ;
        RECT 9.990 190.120 14.225 190.800 ;
        RECT 14.590 190.120 18.825 190.800 ;
        RECT 19.190 190.120 23.425 190.800 ;
        RECT 7.190 189.930 7.360 190.100 ;
        RECT 7.255 189.910 7.360 189.930 ;
        RECT 8.565 189.910 8.735 190.100 ;
        RECT 9.495 189.930 9.665 190.120 ;
        RECT 9.990 190.100 10.100 190.120 ;
        RECT 14.590 190.100 14.700 190.120 ;
        RECT 19.190 190.100 19.300 190.120 ;
        RECT 9.930 189.930 10.100 190.100 ;
        RECT 14.530 189.930 14.700 190.100 ;
        RECT 19.130 189.930 19.300 190.100 ;
        RECT 9.990 189.910 10.100 189.930 ;
        RECT 14.590 189.910 14.700 189.930 ;
        RECT 19.190 189.910 19.300 189.930 ;
        RECT 7.255 189.000 8.185 189.910 ;
        RECT 8.450 189.000 9.800 189.910 ;
        RECT 9.990 189.230 14.225 189.910 ;
        RECT 14.590 189.230 18.825 189.910 ;
        RECT 19.190 189.230 23.425 189.910 ;
        RECT 10.475 189.000 14.225 189.230 ;
        RECT 15.075 189.000 18.825 189.230 ;
        RECT 19.675 189.000 23.425 189.230 ;
        RECT 15.470 184.680 18.080 185.590 ;
        RECT 18.230 184.680 20.840 185.590 ;
        RECT 21.085 184.680 22.015 185.590 ;
        RECT 22.465 184.680 23.395 185.590 ;
        RECT 17.765 184.490 17.935 184.680 ;
        RECT 20.525 184.490 20.695 184.680 ;
        RECT 21.910 184.660 22.015 184.680 ;
        RECT 23.290 184.660 23.395 184.680 ;
        RECT 21.910 184.490 22.080 184.660 ;
        RECT 23.290 184.490 23.460 184.660 ;
      LAYER li1 ;
        RECT 8.250 196.115 8.980 196.645 ;
        RECT 10.960 196.115 11.135 196.185 ;
        RECT 8.250 195.945 11.135 196.115 ;
        RECT 12.695 195.980 13.425 196.680 ;
        RECT 8.810 193.450 8.980 195.450 ;
        RECT 10.960 195.390 11.135 195.945 ;
        RECT 10.965 193.440 11.135 195.390 ;
        RECT 13.190 193.445 13.360 195.980 ;
        RECT 14.425 194.730 14.755 194.910 ;
        RECT 16.060 194.720 16.230 195.200 ;
        RECT 16.900 194.720 17.070 195.200 ;
        RECT 17.740 194.720 17.910 195.200 ;
        RECT 16.060 194.550 17.070 194.720 ;
        RECT 17.275 194.550 17.910 194.720 ;
        RECT 18.820 194.720 18.990 195.200 ;
        RECT 19.660 194.720 19.830 195.200 ;
        RECT 20.500 194.720 20.670 195.200 ;
        RECT 18.820 194.550 19.830 194.720 ;
        RECT 20.035 194.550 20.670 194.720 ;
        RECT 21.175 194.570 21.505 195.200 ;
        RECT 22.555 194.570 22.885 195.200 ;
        RECT 14.500 194.180 14.865 194.350 ;
        RECT 16.060 194.010 16.555 194.550 ;
        RECT 17.275 194.380 17.445 194.550 ;
        RECT 16.945 194.210 17.445 194.380 ;
        RECT 16.060 193.840 17.070 194.010 ;
        RECT 16.060 192.990 16.230 193.840 ;
        RECT 16.900 192.990 17.070 193.840 ;
        RECT 17.275 193.970 17.445 194.210 ;
        RECT 17.615 194.140 17.995 194.380 ;
        RECT 18.820 194.010 19.315 194.550 ;
        RECT 20.035 194.380 20.205 194.550 ;
        RECT 19.705 194.210 20.205 194.380 ;
        RECT 17.275 193.800 17.990 193.970 ;
        RECT 17.660 192.990 17.990 193.800 ;
        RECT 18.820 193.840 19.830 194.010 ;
        RECT 18.820 192.990 18.990 193.840 ;
        RECT 19.660 192.990 19.830 193.840 ;
        RECT 20.035 193.970 20.205 194.210 ;
        RECT 20.375 194.140 20.755 194.380 ;
        RECT 21.175 193.970 21.405 194.570 ;
        RECT 22.555 194.380 22.785 194.570 ;
        RECT 21.575 194.140 22.785 194.380 ;
        RECT 22.955 194.145 23.315 194.380 ;
        RECT 22.955 194.140 23.285 194.145 ;
        RECT 22.555 193.970 22.785 194.140 ;
        RECT 20.035 193.800 20.750 193.970 ;
        RECT 20.420 192.990 20.750 193.800 ;
        RECT 21.175 192.990 21.505 193.970 ;
        RECT 22.555 192.990 22.885 193.970 ;
        RECT 8.940 191.500 9.270 192.480 ;
        RECT 9.890 192.055 10.330 192.480 ;
        RECT 9.890 191.885 10.885 192.055 ;
        RECT 9.035 190.900 9.205 191.500 ;
        RECT 9.375 191.070 9.710 191.340 ;
        RECT 9.890 191.010 10.380 191.715 ;
        RECT 10.550 191.340 10.885 191.885 ;
        RECT 11.055 191.690 11.325 192.480 ;
        RECT 11.495 192.055 11.745 192.480 ;
        RECT 11.495 191.860 12.300 192.055 ;
        RECT 11.055 191.510 11.780 191.690 ;
        RECT 10.550 191.010 10.960 191.340 ;
        RECT 11.130 191.010 11.780 191.510 ;
        RECT 11.950 191.340 12.300 191.860 ;
        RECT 12.470 191.690 12.720 192.480 ;
        RECT 12.890 192.055 13.160 192.480 ;
        RECT 12.890 191.860 13.715 192.055 ;
        RECT 12.470 191.510 13.195 191.690 ;
        RECT 11.950 191.010 12.375 191.340 ;
        RECT 12.545 191.010 13.195 191.510 ;
        RECT 13.365 191.340 13.715 191.860 ;
        RECT 13.885 191.715 14.320 192.480 ;
        RECT 14.490 192.055 14.930 192.480 ;
        RECT 14.490 191.885 15.485 192.055 ;
        RECT 13.885 191.510 14.980 191.715 ;
        RECT 13.365 191.010 13.790 191.340 ;
        RECT 13.960 191.010 14.980 191.510 ;
        RECT 15.150 191.340 15.485 191.885 ;
        RECT 15.655 191.690 15.925 192.480 ;
        RECT 16.095 192.055 16.345 192.480 ;
        RECT 16.095 191.860 16.900 192.055 ;
        RECT 15.655 191.510 16.380 191.690 ;
        RECT 15.150 191.010 15.560 191.340 ;
        RECT 15.730 191.010 16.380 191.510 ;
        RECT 16.550 191.340 16.900 191.860 ;
        RECT 17.070 191.690 17.320 192.480 ;
        RECT 17.490 192.055 17.760 192.480 ;
        RECT 17.490 191.860 18.315 192.055 ;
        RECT 17.070 191.510 17.795 191.690 ;
        RECT 16.550 191.010 16.975 191.340 ;
        RECT 17.145 191.010 17.795 191.510 ;
        RECT 17.965 191.340 18.315 191.860 ;
        RECT 18.485 191.715 18.920 192.480 ;
        RECT 19.090 192.055 19.530 192.480 ;
        RECT 19.090 191.885 20.085 192.055 ;
        RECT 18.485 191.510 19.580 191.715 ;
        RECT 17.965 191.010 18.390 191.340 ;
        RECT 18.560 191.010 19.580 191.510 ;
        RECT 19.750 191.340 20.085 191.885 ;
        RECT 20.255 191.690 20.525 192.480 ;
        RECT 20.695 192.055 20.945 192.480 ;
        RECT 20.695 191.860 21.500 192.055 ;
        RECT 20.255 191.510 20.980 191.690 ;
        RECT 19.750 191.010 20.160 191.340 ;
        RECT 20.330 191.010 20.980 191.510 ;
        RECT 21.150 191.340 21.500 191.860 ;
        RECT 21.670 191.690 21.920 192.480 ;
        RECT 22.090 192.055 22.360 192.480 ;
        RECT 22.090 191.860 22.915 192.055 ;
        RECT 21.670 191.510 22.395 191.690 ;
        RECT 21.150 191.010 21.575 191.340 ;
        RECT 21.745 191.010 22.395 191.510 ;
        RECT 22.565 191.340 22.915 191.860 ;
        RECT 23.085 191.510 23.520 192.480 ;
        RECT 22.565 191.010 22.990 191.340 ;
        RECT 8.510 190.270 9.205 190.900 ;
        RECT 10.550 190.840 10.885 191.010 ;
        RECT 11.130 190.840 11.325 191.010 ;
        RECT 11.950 190.840 12.300 191.010 ;
        RECT 12.545 190.840 12.720 191.010 ;
        RECT 13.365 190.840 13.715 191.010 ;
        RECT 13.960 190.840 14.320 191.010 ;
        RECT 15.150 190.840 15.485 191.010 ;
        RECT 15.730 190.840 15.925 191.010 ;
        RECT 16.550 190.840 16.900 191.010 ;
        RECT 17.145 190.840 17.320 191.010 ;
        RECT 17.965 190.840 18.315 191.010 ;
        RECT 18.560 190.840 18.920 191.010 ;
        RECT 19.750 190.840 20.085 191.010 ;
        RECT 20.330 190.840 20.525 191.010 ;
        RECT 21.150 190.840 21.500 191.010 ;
        RECT 21.745 190.840 21.920 191.010 ;
        RECT 22.565 190.840 22.915 191.010 ;
        RECT 23.160 190.840 23.520 191.510 ;
        RECT 9.890 190.670 10.885 190.840 ;
        RECT 9.890 190.270 10.330 190.670 ;
        RECT 11.055 190.270 11.325 190.840 ;
        RECT 11.495 190.670 12.300 190.840 ;
        RECT 11.495 190.270 11.745 190.670 ;
        RECT 12.470 190.270 12.720 190.840 ;
        RECT 12.890 190.670 13.715 190.840 ;
        RECT 12.890 190.270 13.160 190.670 ;
        RECT 13.885 190.270 14.320 190.840 ;
        RECT 14.490 190.670 15.485 190.840 ;
        RECT 14.490 190.270 14.930 190.670 ;
        RECT 15.655 190.270 15.925 190.840 ;
        RECT 16.095 190.670 16.900 190.840 ;
        RECT 16.095 190.270 16.345 190.670 ;
        RECT 17.070 190.270 17.320 190.840 ;
        RECT 17.490 190.670 18.315 190.840 ;
        RECT 17.490 190.270 17.760 190.670 ;
        RECT 18.485 190.270 18.920 190.840 ;
        RECT 19.090 190.670 20.085 190.840 ;
        RECT 19.090 190.270 19.530 190.670 ;
        RECT 20.255 190.270 20.525 190.840 ;
        RECT 20.695 190.670 21.500 190.840 ;
        RECT 20.695 190.270 20.945 190.670 ;
        RECT 21.670 190.270 21.920 190.840 ;
        RECT 22.090 190.670 22.915 190.840 ;
        RECT 22.090 190.270 22.360 190.670 ;
        RECT 23.085 190.270 23.520 190.840 ;
        RECT 7.765 189.130 8.095 189.760 ;
        RECT 7.865 188.940 8.095 189.130 ;
        RECT 9.025 189.130 9.720 189.760 ;
        RECT 9.890 189.360 10.330 189.760 ;
        RECT 9.890 189.190 10.885 189.360 ;
        RECT 11.055 189.190 11.325 189.760 ;
        RECT 11.495 189.360 11.745 189.760 ;
        RECT 11.495 189.190 12.300 189.360 ;
        RECT 12.470 189.190 12.720 189.760 ;
        RECT 12.890 189.360 13.160 189.760 ;
        RECT 12.890 189.190 13.715 189.360 ;
        RECT 13.885 189.190 14.320 189.760 ;
        RECT 14.490 189.360 14.930 189.760 ;
        RECT 14.490 189.190 15.485 189.360 ;
        RECT 15.655 189.190 15.925 189.760 ;
        RECT 16.095 189.360 16.345 189.760 ;
        RECT 16.095 189.190 16.900 189.360 ;
        RECT 17.070 189.190 17.320 189.760 ;
        RECT 17.490 189.360 17.760 189.760 ;
        RECT 17.490 189.190 18.315 189.360 ;
        RECT 18.485 189.190 18.920 189.760 ;
        RECT 19.090 189.360 19.530 189.760 ;
        RECT 19.090 189.190 20.085 189.360 ;
        RECT 20.255 189.190 20.525 189.760 ;
        RECT 20.695 189.360 20.945 189.760 ;
        RECT 20.695 189.190 21.500 189.360 ;
        RECT 21.670 189.190 21.920 189.760 ;
        RECT 22.090 189.360 22.360 189.760 ;
        RECT 22.090 189.190 22.915 189.360 ;
        RECT 23.085 189.190 23.520 189.760 ;
        RECT 8.520 188.940 8.855 188.960 ;
        RECT 7.865 188.725 8.855 188.940 ;
        RECT 7.865 188.530 8.095 188.725 ;
        RECT 8.520 188.690 8.855 188.725 ;
        RECT 9.025 188.530 9.195 189.130 ;
        RECT 10.550 189.020 10.885 189.190 ;
        RECT 11.130 189.020 11.325 189.190 ;
        RECT 11.950 189.020 12.300 189.190 ;
        RECT 12.545 189.020 12.720 189.190 ;
        RECT 13.365 189.020 13.715 189.190 ;
        RECT 13.960 189.020 14.320 189.190 ;
        RECT 15.150 189.020 15.485 189.190 ;
        RECT 15.730 189.020 15.925 189.190 ;
        RECT 16.550 189.020 16.900 189.190 ;
        RECT 17.145 189.020 17.320 189.190 ;
        RECT 17.965 189.020 18.315 189.190 ;
        RECT 18.560 189.020 18.920 189.190 ;
        RECT 19.750 189.020 20.085 189.190 ;
        RECT 20.330 189.020 20.525 189.190 ;
        RECT 21.150 189.020 21.500 189.190 ;
        RECT 21.745 189.020 21.920 189.190 ;
        RECT 22.565 189.020 22.915 189.190 ;
        RECT 9.365 188.690 9.700 188.940 ;
        RECT 7.765 187.550 8.095 188.530 ;
        RECT 8.960 187.550 9.290 188.530 ;
        RECT 9.890 188.315 10.380 189.020 ;
        RECT 10.550 188.690 10.960 189.020 ;
        RECT 10.550 188.145 10.885 188.690 ;
        RECT 11.130 188.520 11.780 189.020 ;
        RECT 9.890 187.975 10.885 188.145 ;
        RECT 11.055 188.340 11.780 188.520 ;
        RECT 11.950 188.690 12.375 189.020 ;
        RECT 9.890 187.550 10.330 187.975 ;
        RECT 11.055 187.550 11.325 188.340 ;
        RECT 11.950 188.170 12.300 188.690 ;
        RECT 12.545 188.520 13.195 189.020 ;
        RECT 11.495 187.975 12.300 188.170 ;
        RECT 12.470 188.340 13.195 188.520 ;
        RECT 13.365 188.690 13.790 189.020 ;
        RECT 11.495 187.550 11.745 187.975 ;
        RECT 12.470 187.550 12.720 188.340 ;
        RECT 13.365 188.170 13.715 188.690 ;
        RECT 13.960 188.520 14.980 189.020 ;
        RECT 12.890 187.975 13.715 188.170 ;
        RECT 13.885 188.315 14.980 188.520 ;
        RECT 15.150 188.690 15.560 189.020 ;
        RECT 12.890 187.550 13.160 187.975 ;
        RECT 13.885 187.550 14.320 188.315 ;
        RECT 15.150 188.145 15.485 188.690 ;
        RECT 15.730 188.520 16.380 189.020 ;
        RECT 14.490 187.975 15.485 188.145 ;
        RECT 15.655 188.340 16.380 188.520 ;
        RECT 16.550 188.690 16.975 189.020 ;
        RECT 14.490 187.550 14.930 187.975 ;
        RECT 15.655 187.550 15.925 188.340 ;
        RECT 16.550 188.170 16.900 188.690 ;
        RECT 17.145 188.520 17.795 189.020 ;
        RECT 16.095 187.975 16.900 188.170 ;
        RECT 17.070 188.340 17.795 188.520 ;
        RECT 17.965 188.690 18.390 189.020 ;
        RECT 16.095 187.550 16.345 187.975 ;
        RECT 17.070 187.550 17.320 188.340 ;
        RECT 17.965 188.170 18.315 188.690 ;
        RECT 18.560 188.520 19.580 189.020 ;
        RECT 17.490 187.975 18.315 188.170 ;
        RECT 18.485 188.315 19.580 188.520 ;
        RECT 19.750 188.690 20.160 189.020 ;
        RECT 17.490 187.550 17.760 187.975 ;
        RECT 18.485 187.550 18.920 188.315 ;
        RECT 19.750 188.145 20.085 188.690 ;
        RECT 20.330 188.520 20.980 189.020 ;
        RECT 19.090 187.975 20.085 188.145 ;
        RECT 20.255 188.340 20.980 188.520 ;
        RECT 21.150 188.690 21.575 189.020 ;
        RECT 19.090 187.550 19.530 187.975 ;
        RECT 20.255 187.550 20.525 188.340 ;
        RECT 21.150 188.170 21.500 188.690 ;
        RECT 21.745 188.520 22.395 189.020 ;
        RECT 20.695 187.975 21.500 188.170 ;
        RECT 21.670 188.340 22.395 188.520 ;
        RECT 22.565 188.690 22.990 189.020 ;
        RECT 20.695 187.550 20.945 187.975 ;
        RECT 21.670 187.550 21.920 188.340 ;
        RECT 22.565 188.170 22.915 188.690 ;
        RECT 23.160 188.520 23.520 189.190 ;
        RECT 22.090 187.975 22.915 188.170 ;
        RECT 22.090 187.550 22.360 187.975 ;
        RECT 23.085 187.550 23.520 188.520 ;
        RECT 8.400 185.935 8.695 186.875 ;
        RECT 9.785 185.145 9.955 186.585 ;
        RECT 9.730 184.605 9.955 185.145 ;
        RECT 11.365 185.145 11.535 186.585 ;
        RECT 12.185 186.275 12.355 186.585 ;
        RECT 12.180 185.145 12.355 186.275 ;
        RECT 11.365 184.605 11.590 185.145 ;
        RECT 12.115 184.605 12.355 185.145 ;
        RECT 12.975 184.190 13.145 186.585 ;
        RECT 13.765 185.145 13.935 186.585 ;
        RECT 16.060 186.190 16.230 187.040 ;
        RECT 16.900 186.190 17.070 187.040 ;
        RECT 17.660 186.230 17.990 187.040 ;
        RECT 16.060 186.020 17.070 186.190 ;
        RECT 17.275 186.060 17.990 186.230 ;
        RECT 18.820 186.190 18.990 187.040 ;
        RECT 19.660 186.190 19.830 187.040 ;
        RECT 20.420 186.230 20.750 187.040 ;
        RECT 14.420 185.690 14.760 185.860 ;
        RECT 16.060 185.480 16.555 186.020 ;
        RECT 17.275 185.820 17.445 186.060 ;
        RECT 18.820 186.020 19.830 186.190 ;
        RECT 20.035 186.060 20.750 186.230 ;
        RECT 21.175 186.060 21.505 187.040 ;
        RECT 22.555 186.060 22.885 187.040 ;
        RECT 16.945 185.650 17.445 185.820 ;
        RECT 17.615 185.650 17.995 185.890 ;
        RECT 17.275 185.480 17.445 185.650 ;
        RECT 18.820 185.480 19.315 186.020 ;
        RECT 20.035 185.820 20.205 186.060 ;
        RECT 19.705 185.650 20.205 185.820 ;
        RECT 20.375 185.650 20.755 185.890 ;
        RECT 20.035 185.480 20.205 185.650 ;
        RECT 16.060 185.310 17.070 185.480 ;
        RECT 17.275 185.310 17.910 185.480 ;
        RECT 13.765 184.640 14.000 185.145 ;
        RECT 14.565 184.935 14.780 185.290 ;
        RECT 16.060 184.830 16.230 185.310 ;
        RECT 16.900 184.830 17.070 185.310 ;
        RECT 17.740 184.830 17.910 185.310 ;
        RECT 18.820 185.310 19.830 185.480 ;
        RECT 20.035 185.310 20.670 185.480 ;
        RECT 18.820 184.830 18.990 185.310 ;
        RECT 19.660 184.830 19.830 185.310 ;
        RECT 20.500 184.830 20.670 185.310 ;
        RECT 21.175 185.460 21.405 186.060 ;
        RECT 22.555 185.890 22.785 186.060 ;
        RECT 21.575 185.650 22.785 185.890 ;
        RECT 22.955 185.655 23.305 185.890 ;
        RECT 22.955 185.650 23.285 185.655 ;
        RECT 22.555 185.460 22.785 185.650 ;
        RECT 21.175 184.830 21.505 185.460 ;
        RECT 22.555 184.830 22.885 185.460 ;
        RECT 13.765 184.190 14.395 184.640 ;
        RECT 12.690 183.515 13.425 184.190 ;
        RECT 13.760 183.535 14.495 184.190 ;
      LAYER mcon ;
        RECT 8.310 196.395 8.520 196.605 ;
        RECT 8.710 196.395 8.920 196.605 ;
        RECT 8.310 195.995 8.520 196.205 ;
        RECT 8.710 195.995 8.920 196.205 ;
        RECT 12.755 196.430 12.965 196.640 ;
        RECT 13.155 196.430 13.365 196.640 ;
        RECT 10.960 195.955 11.135 196.150 ;
        RECT 12.755 196.030 12.965 196.240 ;
        RECT 13.155 196.030 13.365 196.240 ;
        RECT 8.810 193.530 8.980 193.910 ;
        RECT 14.505 194.735 14.675 194.905 ;
        RECT 21.255 194.630 21.425 194.800 ;
        RECT 14.605 194.180 14.775 194.350 ;
        RECT 16.265 194.180 16.440 194.350 ;
        RECT 17.765 194.180 17.935 194.350 ;
        RECT 19.000 193.895 19.175 194.065 ;
        RECT 20.525 194.180 20.695 194.350 ;
        RECT 21.695 194.180 21.865 194.350 ;
        RECT 23.075 194.180 23.250 194.355 ;
        RECT 9.035 191.135 9.205 191.305 ;
        RECT 9.495 191.120 9.665 191.290 ;
        RECT 10.145 191.090 10.315 191.260 ;
        RECT 23.310 191.120 23.480 191.290 ;
        RECT 9.025 188.765 9.195 188.935 ;
        RECT 9.445 188.770 9.615 188.940 ;
        RECT 9.930 188.740 10.100 188.910 ;
        RECT 23.310 188.740 23.480 188.910 ;
        RECT 8.430 186.550 8.660 186.790 ;
        RECT 8.430 186.000 8.660 186.225 ;
        RECT 9.785 185.450 9.955 185.720 ;
        RECT 11.365 185.445 11.535 185.715 ;
        RECT 12.180 185.475 12.355 185.730 ;
        RECT 13.765 185.460 13.935 185.715 ;
        RECT 14.510 185.690 14.680 185.860 ;
        RECT 16.185 185.685 16.355 185.855 ;
        RECT 19.035 185.965 19.205 186.135 ;
        RECT 17.765 185.680 17.935 185.850 ;
        RECT 20.525 185.680 20.695 185.850 ;
        RECT 14.580 185.015 14.765 185.190 ;
        RECT 22.615 185.680 22.785 185.850 ;
        RECT 23.075 185.680 23.245 185.850 ;
        RECT 21.255 185.230 21.425 185.400 ;
        RECT 12.755 183.940 12.965 184.150 ;
        RECT 13.155 183.940 13.365 184.150 ;
        RECT 12.755 183.555 12.965 183.750 ;
        RECT 13.155 183.555 13.365 183.750 ;
        RECT 13.825 183.940 14.035 184.150 ;
        RECT 14.225 183.940 14.435 184.150 ;
        RECT 13.825 183.565 14.035 183.735 ;
        RECT 14.225 183.565 14.435 183.735 ;
      LAYER met1 ;
        RECT 8.250 196.165 8.980 196.645 ;
        RECT 10.835 196.165 11.195 196.180 ;
        RECT 8.250 195.945 11.195 196.165 ;
        RECT 12.695 195.980 13.425 196.680 ;
        RECT 10.835 195.925 11.195 195.945 ;
        RECT 14.445 194.910 14.750 194.935 ;
        RECT 14.445 194.730 16.850 194.910 ;
        RECT 14.445 194.705 14.750 194.730 ;
        RECT 14.500 194.145 16.505 194.380 ;
        RECT 7.475 193.850 7.845 193.905 ;
        RECT 8.775 193.850 9.010 193.970 ;
        RECT 16.710 193.860 16.850 194.730 ;
        RECT 18.075 194.600 21.485 194.830 ;
        RECT 17.615 194.380 17.935 194.400 ;
        RECT 18.075 194.380 18.250 194.600 ;
        RECT 20.460 194.380 20.780 194.390 ;
        RECT 23.050 194.385 23.310 194.425 ;
        RECT 17.615 194.150 18.250 194.380 ;
        RECT 20.375 194.150 21.925 194.380 ;
        RECT 17.615 194.140 17.935 194.150 ;
        RECT 20.460 194.130 20.780 194.150 ;
        RECT 23.040 194.145 23.310 194.385 ;
        RECT 18.960 193.860 19.205 194.125 ;
        RECT 23.050 194.105 23.310 194.145 ;
        RECT 7.475 193.585 9.010 193.850 ;
        RECT 16.705 193.685 19.205 193.860 ;
        RECT 8.775 193.470 9.010 193.585 ;
        RECT 18.040 191.670 18.300 191.770 ;
        RECT 9.465 191.525 18.300 191.670 ;
        RECT 9.005 191.050 9.235 191.375 ;
        RECT 9.465 191.060 9.705 191.525 ;
        RECT 18.040 191.450 18.300 191.525 ;
        RECT 9.025 190.920 9.235 191.050 ;
        RECT 10.095 191.010 10.380 191.375 ;
        RECT 23.260 191.045 23.520 191.365 ;
        RECT 10.095 190.920 10.315 191.010 ;
        RECT 9.025 190.775 10.315 190.920 ;
        RECT 17.585 189.445 17.905 189.485 ;
        RECT 9.370 189.270 17.905 189.445 ;
        RECT 8.995 188.540 9.225 189.255 ;
        RECT 9.370 188.690 9.700 189.270 ;
        RECT 17.585 189.225 17.905 189.270 ;
        RECT 9.900 188.540 10.160 188.975 ;
        RECT 23.260 188.665 23.520 188.985 ;
        RECT 8.995 188.400 10.160 188.540 ;
        RECT 8.400 185.750 8.695 186.875 ;
        RECT 16.660 186.325 19.205 186.500 ;
        RECT 8.400 185.420 11.600 185.750 ;
        RECT 12.080 185.425 14.020 185.760 ;
        RECT 14.335 185.655 16.475 185.890 ;
        RECT 8.400 185.415 8.695 185.420 ;
        RECT 9.725 185.415 11.600 185.420 ;
        RECT 16.660 185.345 16.875 186.325 ;
        RECT 19.030 186.165 19.205 186.325 ;
        RECT 17.735 185.880 18.230 185.910 ;
        RECT 19.005 185.905 19.240 186.165 ;
        RECT 17.615 185.650 18.230 185.880 ;
        RECT 14.845 185.290 16.875 185.345 ;
        RECT 14.550 185.170 16.875 185.290 ;
        RECT 18.050 185.430 18.230 185.650 ;
        RECT 20.375 185.890 20.780 185.900 ;
        RECT 20.375 185.650 22.845 185.890 ;
        RECT 20.375 185.640 20.780 185.650 ;
        RECT 23.045 185.615 23.305 185.935 ;
        RECT 18.050 185.190 21.485 185.430 ;
        RECT 14.550 185.115 14.935 185.170 ;
        RECT 14.550 184.955 14.795 185.115 ;
        RECT 12.690 183.245 13.425 184.190 ;
        RECT 13.760 183.535 14.495 184.190 ;
      LAYER via ;
        RECT 8.310 196.345 8.570 196.605 ;
        RECT 8.660 196.345 8.920 196.605 ;
        RECT 8.310 195.995 8.570 196.255 ;
        RECT 8.660 195.995 8.920 196.255 ;
        RECT 12.755 196.380 13.015 196.640 ;
        RECT 13.105 196.380 13.365 196.640 ;
        RECT 12.755 196.030 13.015 196.290 ;
        RECT 13.105 196.030 13.365 196.290 ;
        RECT 7.515 193.610 7.815 193.870 ;
        RECT 17.645 194.140 17.905 194.400 ;
        RECT 23.050 194.135 23.310 194.395 ;
        RECT 18.040 191.480 18.300 191.740 ;
        RECT 23.260 191.075 23.520 191.335 ;
        RECT 17.615 189.225 17.875 189.485 ;
        RECT 23.260 188.695 23.520 188.955 ;
        RECT 8.415 186.530 8.675 186.790 ;
        RECT 8.415 186.000 8.675 186.260 ;
        RECT 17.765 185.650 18.025 185.910 ;
        RECT 23.045 185.645 23.305 185.905 ;
        RECT 12.755 183.890 13.015 184.150 ;
        RECT 13.105 183.890 13.365 184.150 ;
        RECT 12.755 183.555 13.015 183.815 ;
        RECT 13.105 183.555 13.365 183.815 ;
        RECT 13.825 183.890 14.085 184.150 ;
        RECT 14.175 183.890 14.435 184.150 ;
        RECT 13.825 183.565 14.085 183.825 ;
        RECT 14.175 183.565 14.435 183.825 ;
      LAYER met2 ;
        RECT 8.250 198.880 11.990 199.700 ;
        RECT 8.250 198.870 11.980 198.880 ;
        RECT 7.055 195.845 7.845 196.665 ;
        RECT 8.250 195.945 8.980 198.870 ;
        RECT 16.760 198.775 17.510 199.595 ;
        RECT 16.760 198.770 17.500 198.775 ;
        RECT 7.475 193.585 7.845 195.845 ;
        RECT 8.400 185.935 8.695 195.945 ;
        RECT 12.690 182.380 13.425 196.680 ;
        RECT 13.755 196.265 14.495 196.660 ;
        RECT 13.760 183.535 14.495 196.265 ;
        RECT 16.760 195.845 17.495 198.770 ;
        RECT 17.615 194.140 17.935 194.400 ;
        RECT 17.685 189.485 17.840 194.140 ;
        RECT 23.050 194.105 23.520 194.425 ;
        RECT 18.040 191.450 18.300 191.770 ;
        RECT 17.585 189.225 17.905 189.485 ;
        RECT 18.100 185.925 18.245 191.450 ;
        RECT 23.260 191.045 23.520 194.105 ;
        RECT 23.260 185.935 23.520 188.985 ;
        RECT 17.680 185.630 18.245 185.925 ;
        RECT 23.045 185.615 23.520 185.935 ;
        RECT 12.675 182.375 13.425 182.380 ;
        RECT 12.675 181.955 13.445 182.375 ;
      LAYER via2 ;
        RECT 11.285 199.345 11.565 199.625 ;
        RECT 11.685 199.345 11.965 199.625 ;
        RECT 11.285 198.945 11.565 199.225 ;
        RECT 11.685 198.945 11.965 199.225 ;
        RECT 16.805 199.240 17.085 199.520 ;
        RECT 17.205 199.240 17.485 199.520 ;
        RECT 7.080 196.315 7.360 196.595 ;
        RECT 7.490 196.320 7.770 196.600 ;
        RECT 7.085 195.915 7.365 196.195 ;
        RECT 7.495 195.920 7.775 196.200 ;
        RECT 16.805 198.840 17.085 199.120 ;
        RECT 17.205 198.840 17.485 199.120 ;
        RECT 13.800 196.310 14.080 196.590 ;
        RECT 14.200 196.305 14.480 196.585 ;
        RECT 13.805 195.905 14.085 196.185 ;
        RECT 14.205 195.905 14.485 196.185 ;
        RECT 16.800 196.305 17.080 196.585 ;
        RECT 17.200 196.300 17.480 196.580 ;
        RECT 16.805 195.900 17.085 196.180 ;
        RECT 17.205 195.900 17.485 196.180 ;
        RECT 12.720 182.005 13.000 182.315 ;
        RECT 13.120 182.005 13.400 182.315 ;
      LAYER met3 ;
        RECT 4.730 378.750 9.130 380.000 ;
        RECT 11.530 379.150 17.930 380.000 ;
        RECT 20.330 378.750 29.130 380.000 ;
        RECT 31.530 379.150 37.930 380.000 ;
        RECT 40.330 378.750 49.130 380.000 ;
        RECT 51.530 379.150 57.930 380.000 ;
        RECT 60.330 378.750 69.130 380.000 ;
        RECT 71.530 379.150 77.930 380.000 ;
        RECT 80.330 378.750 89.130 380.000 ;
        RECT 91.530 379.150 97.930 380.000 ;
        RECT 100.330 378.750 104.730 380.000 ;
        RECT 4.730 375.600 104.730 378.750 ;
        RECT 4.730 366.800 5.580 373.200 ;
        RECT 5.980 364.400 23.480 375.600 ;
        RECT 23.880 366.800 25.580 373.200 ;
        RECT 25.980 364.400 43.480 375.600 ;
        RECT 43.880 366.800 45.580 373.200 ;
        RECT 45.980 364.400 63.480 375.600 ;
        RECT 63.880 366.800 65.580 373.200 ;
        RECT 65.980 364.400 83.480 375.600 ;
        RECT 83.880 366.800 85.580 373.200 ;
        RECT 85.980 364.400 103.480 375.600 ;
        RECT 103.880 366.800 104.730 373.200 ;
        RECT 4.730 361.250 104.730 364.400 ;
        RECT 4.730 358.750 9.130 361.250 ;
        RECT 11.530 359.150 17.930 360.850 ;
        RECT 20.330 358.750 29.130 361.250 ;
        RECT 31.530 359.150 37.930 360.850 ;
        RECT 40.330 358.750 49.130 361.250 ;
        RECT 51.530 359.150 57.930 360.850 ;
        RECT 60.330 358.750 69.130 361.250 ;
        RECT 71.530 359.150 77.930 360.850 ;
        RECT 80.330 358.750 89.130 361.250 ;
        RECT 91.530 359.150 97.930 360.850 ;
        RECT 100.330 358.750 104.730 361.250 ;
        RECT 4.730 355.600 104.730 358.750 ;
        RECT 4.730 346.800 5.580 353.200 ;
        RECT 5.980 344.400 23.480 355.600 ;
        RECT 23.880 346.800 25.580 353.200 ;
        RECT 25.980 344.400 43.480 355.600 ;
        RECT 43.880 346.800 45.580 353.200 ;
        RECT 45.980 344.400 63.480 355.600 ;
        RECT 63.880 346.800 65.580 353.200 ;
        RECT 65.980 344.400 83.480 355.600 ;
        RECT 83.880 346.800 85.580 353.200 ;
        RECT 85.980 344.400 103.480 355.600 ;
        RECT 103.880 346.800 104.730 353.200 ;
        RECT 4.730 341.250 104.730 344.400 ;
        RECT 4.730 338.750 9.130 341.250 ;
        RECT 11.530 339.150 17.930 340.850 ;
        RECT 20.330 338.750 29.130 341.250 ;
        RECT 31.530 339.150 37.930 340.850 ;
        RECT 40.330 338.750 49.130 341.250 ;
        RECT 51.530 339.150 57.930 340.850 ;
        RECT 60.330 338.750 69.130 341.250 ;
        RECT 71.530 339.150 77.930 340.850 ;
        RECT 80.330 338.750 89.130 341.250 ;
        RECT 91.530 339.150 97.930 340.850 ;
        RECT 100.330 338.750 104.730 341.250 ;
        RECT 4.730 335.600 104.730 338.750 ;
        RECT 4.730 326.800 5.580 333.200 ;
        RECT 5.980 324.400 23.480 335.600 ;
        RECT 23.880 326.800 25.580 333.200 ;
        RECT 25.980 324.400 43.480 335.600 ;
        RECT 43.880 326.800 45.580 333.200 ;
        RECT 45.980 324.400 63.480 335.600 ;
        RECT 63.880 326.800 65.580 333.200 ;
        RECT 65.980 324.400 83.480 335.600 ;
        RECT 83.880 326.800 85.580 333.200 ;
        RECT 85.980 324.400 103.480 335.600 ;
        RECT 103.880 326.800 104.730 333.200 ;
        RECT 4.730 321.250 104.730 324.400 ;
        RECT 4.730 318.750 9.130 321.250 ;
        RECT 11.530 319.150 17.930 320.850 ;
        RECT 20.330 318.750 29.130 321.250 ;
        RECT 31.530 319.150 37.930 320.850 ;
        RECT 40.330 318.750 49.130 321.250 ;
        RECT 51.530 319.150 57.930 320.850 ;
        RECT 60.330 318.750 69.130 321.250 ;
        RECT 71.530 319.150 77.930 320.850 ;
        RECT 80.330 318.750 89.130 321.250 ;
        RECT 91.530 319.150 97.930 320.850 ;
        RECT 100.330 318.750 104.730 321.250 ;
        RECT 4.730 315.600 104.730 318.750 ;
        RECT 4.730 306.800 5.580 313.200 ;
        RECT 5.980 304.400 23.480 315.600 ;
        RECT 23.880 306.800 25.580 313.200 ;
        RECT 25.980 304.400 43.480 315.600 ;
        RECT 43.880 306.800 45.580 313.200 ;
        RECT 45.980 304.400 63.480 315.600 ;
        RECT 63.880 306.800 65.580 313.200 ;
        RECT 65.980 304.400 83.480 315.600 ;
        RECT 83.880 306.800 85.580 313.200 ;
        RECT 85.980 304.400 103.480 315.600 ;
        RECT 103.880 306.800 104.730 313.200 ;
        RECT 4.730 301.250 104.730 304.400 ;
        RECT 4.730 298.750 9.130 301.250 ;
        RECT 11.530 299.150 17.930 300.850 ;
        RECT 20.330 298.750 29.130 301.250 ;
        RECT 31.530 299.150 37.930 300.850 ;
        RECT 40.330 298.750 49.130 301.250 ;
        RECT 51.530 299.150 57.930 300.850 ;
        RECT 60.330 298.750 69.130 301.250 ;
        RECT 71.530 299.150 77.930 300.850 ;
        RECT 80.330 298.750 89.130 301.250 ;
        RECT 91.530 299.150 97.930 300.850 ;
        RECT 100.330 298.750 104.730 301.250 ;
        RECT 4.730 295.600 104.730 298.750 ;
        RECT 4.730 286.800 5.580 293.200 ;
        RECT 5.980 284.400 23.480 295.600 ;
        RECT 23.880 286.800 25.580 293.200 ;
        RECT 25.980 284.400 43.480 295.600 ;
        RECT 43.880 286.800 45.580 293.200 ;
        RECT 45.980 284.400 63.480 295.600 ;
        RECT 63.880 286.800 65.580 293.200 ;
        RECT 65.980 284.400 83.480 295.600 ;
        RECT 83.880 286.800 85.580 293.200 ;
        RECT 85.980 284.400 103.480 295.600 ;
        RECT 103.880 286.800 104.730 293.200 ;
        RECT 4.730 281.250 104.730 284.400 ;
        RECT 4.730 278.750 9.130 281.250 ;
        RECT 11.530 279.150 17.930 280.850 ;
        RECT 20.330 278.750 29.130 281.250 ;
        RECT 31.530 279.150 37.930 280.850 ;
        RECT 40.330 278.750 49.130 281.250 ;
        RECT 51.530 279.150 57.930 280.850 ;
        RECT 60.330 278.750 69.130 281.250 ;
        RECT 71.530 279.150 77.930 280.850 ;
        RECT 80.330 278.750 89.130 281.250 ;
        RECT 91.530 279.150 97.930 280.850 ;
        RECT 100.330 278.750 104.730 281.250 ;
        RECT 4.730 275.600 104.730 278.750 ;
        RECT 4.730 266.800 5.580 273.200 ;
        RECT 5.980 264.400 23.480 275.600 ;
        RECT 23.880 266.800 25.580 273.200 ;
        RECT 25.980 264.400 43.480 275.600 ;
        RECT 43.880 266.800 45.580 273.200 ;
        RECT 45.980 264.400 63.480 275.600 ;
        RECT 63.880 266.800 65.580 273.200 ;
        RECT 65.980 264.400 83.480 275.600 ;
        RECT 83.880 266.800 85.580 273.200 ;
        RECT 85.980 264.400 103.480 275.600 ;
        RECT 103.880 266.800 104.730 273.200 ;
        RECT 4.730 261.250 104.730 264.400 ;
        RECT 4.730 258.750 9.130 261.250 ;
        RECT 11.530 259.150 17.930 260.850 ;
        RECT 20.330 258.750 29.130 261.250 ;
        RECT 31.530 259.150 37.930 260.850 ;
        RECT 40.330 258.750 49.130 261.250 ;
        RECT 51.530 259.150 57.930 260.850 ;
        RECT 60.330 258.750 69.130 261.250 ;
        RECT 71.530 259.150 77.930 260.850 ;
        RECT 80.330 258.750 89.130 261.250 ;
        RECT 91.530 259.150 97.930 260.850 ;
        RECT 100.330 258.750 104.730 261.250 ;
        RECT 4.730 255.600 104.730 258.750 ;
        RECT 4.730 246.800 5.580 253.200 ;
        RECT 5.980 244.400 23.480 255.600 ;
        RECT 23.880 246.800 25.580 253.200 ;
        RECT 25.980 244.400 43.480 255.600 ;
        RECT 43.880 246.800 45.580 253.200 ;
        RECT 45.980 244.400 63.480 255.600 ;
        RECT 63.880 246.800 65.580 253.200 ;
        RECT 65.980 244.400 83.480 255.600 ;
        RECT 83.880 246.800 85.580 253.200 ;
        RECT 85.980 244.400 103.480 255.600 ;
        RECT 103.880 246.800 104.730 253.200 ;
        RECT 4.730 241.250 104.730 244.400 ;
        RECT 4.730 238.750 9.130 241.250 ;
        RECT 11.530 239.150 17.930 240.850 ;
        RECT 20.330 238.750 29.130 241.250 ;
        RECT 31.530 239.150 37.930 240.850 ;
        RECT 40.330 238.750 49.130 241.250 ;
        RECT 51.530 239.150 57.930 240.850 ;
        RECT 60.330 238.750 69.130 241.250 ;
        RECT 71.530 239.150 77.930 240.850 ;
        RECT 80.330 238.750 89.130 241.250 ;
        RECT 91.530 239.150 97.930 240.850 ;
        RECT 100.330 238.750 104.730 241.250 ;
        RECT 4.730 235.600 104.730 238.750 ;
        RECT 4.730 226.800 5.580 233.200 ;
        RECT 5.980 224.400 23.480 235.600 ;
        RECT 23.880 226.800 25.580 233.200 ;
        RECT 25.980 224.400 43.480 235.600 ;
        RECT 43.880 226.800 45.580 233.200 ;
        RECT 45.980 224.400 63.480 235.600 ;
        RECT 63.880 226.800 65.580 233.200 ;
        RECT 65.980 224.400 83.480 235.600 ;
        RECT 83.880 226.800 85.580 233.200 ;
        RECT 85.980 224.400 103.480 235.600 ;
        RECT 103.880 226.800 104.730 233.200 ;
        RECT 4.730 221.250 104.730 224.400 ;
        RECT 4.730 220.000 9.130 221.250 ;
        RECT 11.530 220.000 17.930 220.850 ;
        RECT 20.330 220.000 29.130 221.250 ;
        RECT 31.530 220.000 37.930 220.850 ;
        RECT 40.330 220.000 49.130 221.250 ;
        RECT 51.530 220.000 57.930 220.850 ;
        RECT 60.330 220.000 69.130 221.250 ;
        RECT 71.530 220.000 77.930 220.850 ;
        RECT 80.330 220.000 89.130 221.250 ;
        RECT 91.530 220.000 97.930 220.850 ;
        RECT 100.330 220.000 104.730 221.250 ;
        RECT 11.240 198.875 12.005 199.700 ;
        RECT 16.760 198.770 21.725 199.600 ;
        RECT 13.445 196.665 17.510 196.670 ;
        RECT 7.055 195.845 17.510 196.665 ;
        RECT 12.675 182.375 13.440 182.380 ;
        RECT 12.675 181.955 13.445 182.375 ;
        RECT 11.530 159.150 17.930 160.000 ;
        RECT 31.530 159.150 37.930 160.000 ;
        RECT 51.530 159.150 57.930 160.000 ;
        RECT 71.530 159.150 77.930 160.000 ;
        RECT 91.530 159.150 97.930 160.000 ;
        RECT 4.730 146.800 5.580 153.200 ;
        RECT 23.880 146.800 25.580 153.200 ;
        RECT 43.880 146.800 45.580 153.200 ;
        RECT 63.880 146.800 65.580 153.200 ;
        RECT 83.880 146.800 85.580 153.200 ;
        RECT 103.880 146.800 104.730 153.200 ;
        RECT 11.530 139.150 17.930 140.850 ;
        RECT 31.530 139.150 37.930 140.850 ;
        RECT 51.530 139.150 57.930 140.850 ;
        RECT 71.530 139.150 77.930 140.850 ;
        RECT 91.530 139.150 97.930 140.850 ;
        RECT 4.730 126.800 5.580 133.200 ;
        RECT 23.880 126.800 25.580 133.200 ;
        RECT 43.880 126.800 45.580 133.200 ;
        RECT 63.880 126.800 65.580 133.200 ;
        RECT 83.880 126.800 85.580 133.200 ;
        RECT 103.880 126.800 104.730 133.200 ;
        RECT 11.530 119.150 17.930 120.850 ;
        RECT 31.530 119.150 37.930 120.850 ;
        RECT 51.530 119.150 57.930 120.850 ;
        RECT 71.530 119.150 77.930 120.850 ;
        RECT 91.530 119.150 97.930 120.850 ;
        RECT 4.730 106.800 5.580 113.200 ;
        RECT 23.880 106.800 25.580 113.200 ;
        RECT 43.880 106.800 45.580 113.200 ;
        RECT 63.880 106.800 65.580 113.200 ;
        RECT 83.880 106.800 85.580 113.200 ;
        RECT 103.880 106.800 104.730 113.200 ;
        RECT 11.530 99.150 17.930 100.850 ;
        RECT 31.530 99.150 37.930 100.850 ;
        RECT 51.530 99.150 57.930 100.850 ;
        RECT 71.530 99.150 77.930 100.850 ;
        RECT 91.530 99.150 97.930 100.850 ;
        RECT 4.730 86.800 5.580 93.200 ;
        RECT 23.880 86.800 25.580 93.200 ;
        RECT 43.880 86.800 45.580 93.200 ;
        RECT 63.880 86.800 65.580 93.200 ;
        RECT 83.880 86.800 85.580 93.200 ;
        RECT 103.880 86.800 104.730 93.200 ;
        RECT 11.530 79.150 17.930 80.850 ;
        RECT 31.530 79.150 37.930 80.850 ;
        RECT 51.530 79.150 57.930 80.850 ;
        RECT 71.530 79.150 77.930 80.850 ;
        RECT 91.530 79.150 97.930 80.850 ;
        RECT 4.730 66.800 5.580 73.200 ;
        RECT 23.880 66.800 25.580 73.200 ;
        RECT 43.880 66.800 45.580 73.200 ;
        RECT 63.880 66.800 65.580 73.200 ;
        RECT 83.880 66.800 85.580 73.200 ;
        RECT 103.880 66.800 104.730 73.200 ;
        RECT 11.530 59.150 17.930 60.850 ;
        RECT 31.530 59.150 37.930 60.850 ;
        RECT 51.530 59.150 57.930 60.850 ;
        RECT 71.530 59.150 77.930 60.850 ;
        RECT 91.530 59.150 97.930 60.850 ;
        RECT 4.730 46.800 5.580 53.200 ;
        RECT 23.880 46.800 25.580 53.200 ;
        RECT 43.880 46.800 45.580 53.200 ;
        RECT 63.880 46.800 65.580 53.200 ;
        RECT 83.880 46.800 85.580 53.200 ;
        RECT 103.880 46.800 104.730 53.200 ;
        RECT 11.530 39.150 17.930 40.850 ;
        RECT 31.530 39.150 37.930 40.850 ;
        RECT 51.530 39.150 57.930 40.850 ;
        RECT 71.530 39.150 77.930 40.850 ;
        RECT 91.530 39.150 97.930 40.850 ;
        RECT 4.730 26.800 5.580 33.200 ;
        RECT 23.880 26.800 25.580 33.200 ;
        RECT 43.880 26.800 45.580 33.200 ;
        RECT 63.880 26.800 65.580 33.200 ;
        RECT 83.880 26.800 85.580 33.200 ;
        RECT 103.880 26.800 104.730 33.200 ;
        RECT 11.530 19.150 17.930 20.850 ;
        RECT 31.530 19.150 37.930 20.850 ;
        RECT 51.530 19.150 57.930 20.850 ;
        RECT 71.530 19.150 77.930 20.850 ;
        RECT 91.530 19.150 97.930 20.850 ;
        RECT 4.730 6.800 5.580 13.200 ;
        RECT 23.880 6.800 25.580 13.200 ;
        RECT 43.880 6.800 45.580 13.200 ;
        RECT 63.880 6.800 65.580 13.200 ;
        RECT 83.880 6.800 85.580 13.200 ;
        RECT 103.880 6.800 104.730 13.200 ;
        RECT 11.530 0.000 17.930 0.850 ;
        RECT 31.530 0.000 37.930 0.850 ;
        RECT 51.530 0.000 57.930 0.850 ;
        RECT 71.530 0.000 77.930 0.850 ;
        RECT 91.530 0.000 97.930 0.850 ;
      LAYER via3 ;
        RECT 4.830 379.050 5.680 379.900 ;
        RECT 5.780 379.050 6.630 379.900 ;
        RECT 7.230 379.050 8.080 379.900 ;
        RECT 8.180 379.050 9.030 379.900 ;
        RECT 11.630 379.250 12.280 379.900 ;
        RECT 12.430 379.250 13.080 379.900 ;
        RECT 13.230 379.250 13.880 379.900 ;
        RECT 15.580 379.250 16.230 379.900 ;
        RECT 16.380 379.250 17.030 379.900 ;
        RECT 17.180 379.250 17.830 379.900 ;
        RECT 4.830 378.100 5.680 378.950 ;
        RECT 20.430 379.050 21.280 379.900 ;
        RECT 21.380 379.050 22.230 379.900 ;
        RECT 22.830 379.050 23.680 379.900 ;
        RECT 23.780 379.050 24.630 379.900 ;
        RECT 24.830 379.050 25.680 379.900 ;
        RECT 25.780 379.050 26.630 379.900 ;
        RECT 27.230 379.050 28.080 379.900 ;
        RECT 28.180 379.050 29.030 379.900 ;
        RECT 31.630 379.250 32.280 379.900 ;
        RECT 32.430 379.250 33.080 379.900 ;
        RECT 33.230 379.250 33.880 379.900 ;
        RECT 35.580 379.250 36.230 379.900 ;
        RECT 36.380 379.250 37.030 379.900 ;
        RECT 37.180 379.250 37.830 379.900 ;
        RECT 23.780 378.100 24.630 378.950 ;
        RECT 24.830 378.100 25.680 378.950 ;
        RECT 40.430 379.050 41.280 379.900 ;
        RECT 41.380 379.050 42.230 379.900 ;
        RECT 42.830 379.050 43.680 379.900 ;
        RECT 43.780 379.050 44.630 379.900 ;
        RECT 44.830 379.050 45.680 379.900 ;
        RECT 45.780 379.050 46.630 379.900 ;
        RECT 47.230 379.050 48.080 379.900 ;
        RECT 48.180 379.050 49.030 379.900 ;
        RECT 51.630 379.250 52.280 379.900 ;
        RECT 52.430 379.250 53.080 379.900 ;
        RECT 53.230 379.250 53.880 379.900 ;
        RECT 55.580 379.250 56.230 379.900 ;
        RECT 56.380 379.250 57.030 379.900 ;
        RECT 57.180 379.250 57.830 379.900 ;
        RECT 43.780 378.100 44.630 378.950 ;
        RECT 44.830 378.100 45.680 378.950 ;
        RECT 60.430 379.050 61.280 379.900 ;
        RECT 61.380 379.050 62.230 379.900 ;
        RECT 62.830 379.050 63.680 379.900 ;
        RECT 63.780 379.050 64.630 379.900 ;
        RECT 64.830 379.050 65.680 379.900 ;
        RECT 65.780 379.050 66.630 379.900 ;
        RECT 67.230 379.050 68.080 379.900 ;
        RECT 68.180 379.050 69.030 379.900 ;
        RECT 71.630 379.250 72.280 379.900 ;
        RECT 72.430 379.250 73.080 379.900 ;
        RECT 73.230 379.250 73.880 379.900 ;
        RECT 75.580 379.250 76.230 379.900 ;
        RECT 76.380 379.250 77.030 379.900 ;
        RECT 77.180 379.250 77.830 379.900 ;
        RECT 63.780 378.100 64.630 378.950 ;
        RECT 64.830 378.100 65.680 378.950 ;
        RECT 80.430 379.050 81.280 379.900 ;
        RECT 81.380 379.050 82.230 379.900 ;
        RECT 82.830 379.050 83.680 379.900 ;
        RECT 83.780 379.050 84.630 379.900 ;
        RECT 84.830 379.050 85.680 379.900 ;
        RECT 85.780 379.050 86.630 379.900 ;
        RECT 87.230 379.050 88.080 379.900 ;
        RECT 88.180 379.050 89.030 379.900 ;
        RECT 91.630 379.250 92.280 379.900 ;
        RECT 92.430 379.250 93.080 379.900 ;
        RECT 93.230 379.250 93.880 379.900 ;
        RECT 95.580 379.250 96.230 379.900 ;
        RECT 96.380 379.250 97.030 379.900 ;
        RECT 97.180 379.250 97.830 379.900 ;
        RECT 83.780 378.100 84.630 378.950 ;
        RECT 84.830 378.100 85.680 378.950 ;
        RECT 100.430 379.050 101.280 379.900 ;
        RECT 101.380 379.050 102.230 379.900 ;
        RECT 102.830 379.050 103.680 379.900 ;
        RECT 103.780 379.050 104.630 379.900 ;
        RECT 103.780 378.100 104.630 378.950 ;
        RECT 4.830 376.650 5.680 377.500 ;
        RECT 23.780 376.650 24.630 377.500 ;
        RECT 24.830 376.650 25.680 377.500 ;
        RECT 43.780 376.650 44.630 377.500 ;
        RECT 44.830 376.650 45.680 377.500 ;
        RECT 63.780 376.650 64.630 377.500 ;
        RECT 64.830 376.650 65.680 377.500 ;
        RECT 83.780 376.650 84.630 377.500 ;
        RECT 84.830 376.650 85.680 377.500 ;
        RECT 103.780 376.650 104.630 377.500 ;
        RECT 4.830 375.700 5.680 376.550 ;
        RECT 23.780 375.700 24.630 376.550 ;
        RECT 24.830 375.700 25.680 376.550 ;
        RECT 43.780 375.700 44.630 376.550 ;
        RECT 44.830 375.700 45.680 376.550 ;
        RECT 63.780 375.700 64.630 376.550 ;
        RECT 64.830 375.700 65.680 376.550 ;
        RECT 83.780 375.700 84.630 376.550 ;
        RECT 84.830 375.700 85.680 376.550 ;
        RECT 103.780 375.700 104.630 376.550 ;
        RECT 4.830 372.450 5.480 373.100 ;
        RECT 4.830 371.650 5.480 372.300 ;
        RECT 4.830 370.850 5.480 371.500 ;
        RECT 4.830 368.500 5.480 369.150 ;
        RECT 4.830 367.700 5.480 368.350 ;
        RECT 4.830 366.900 5.480 367.550 ;
        RECT 23.980 372.450 24.630 373.100 ;
        RECT 24.830 372.450 25.480 373.100 ;
        RECT 23.980 371.650 24.630 372.300 ;
        RECT 24.830 371.650 25.480 372.300 ;
        RECT 23.980 370.850 24.630 371.500 ;
        RECT 24.830 370.850 25.480 371.500 ;
        RECT 23.980 368.500 24.630 369.150 ;
        RECT 24.830 368.500 25.480 369.150 ;
        RECT 23.980 367.700 24.630 368.350 ;
        RECT 24.830 367.700 25.480 368.350 ;
        RECT 23.980 366.900 24.630 367.550 ;
        RECT 24.830 366.900 25.480 367.550 ;
        RECT 43.980 372.450 44.630 373.100 ;
        RECT 44.830 372.450 45.480 373.100 ;
        RECT 43.980 371.650 44.630 372.300 ;
        RECT 44.830 371.650 45.480 372.300 ;
        RECT 43.980 370.850 44.630 371.500 ;
        RECT 44.830 370.850 45.480 371.500 ;
        RECT 43.980 368.500 44.630 369.150 ;
        RECT 44.830 368.500 45.480 369.150 ;
        RECT 43.980 367.700 44.630 368.350 ;
        RECT 44.830 367.700 45.480 368.350 ;
        RECT 43.980 366.900 44.630 367.550 ;
        RECT 44.830 366.900 45.480 367.550 ;
        RECT 63.980 372.450 64.630 373.100 ;
        RECT 64.830 372.450 65.480 373.100 ;
        RECT 63.980 371.650 64.630 372.300 ;
        RECT 64.830 371.650 65.480 372.300 ;
        RECT 63.980 370.850 64.630 371.500 ;
        RECT 64.830 370.850 65.480 371.500 ;
        RECT 63.980 368.500 64.630 369.150 ;
        RECT 64.830 368.500 65.480 369.150 ;
        RECT 63.980 367.700 64.630 368.350 ;
        RECT 64.830 367.700 65.480 368.350 ;
        RECT 63.980 366.900 64.630 367.550 ;
        RECT 64.830 366.900 65.480 367.550 ;
        RECT 83.980 372.450 84.630 373.100 ;
        RECT 84.830 372.450 85.480 373.100 ;
        RECT 83.980 371.650 84.630 372.300 ;
        RECT 84.830 371.650 85.480 372.300 ;
        RECT 83.980 370.850 84.630 371.500 ;
        RECT 84.830 370.850 85.480 371.500 ;
        RECT 83.980 368.500 84.630 369.150 ;
        RECT 84.830 368.500 85.480 369.150 ;
        RECT 83.980 367.700 84.630 368.350 ;
        RECT 84.830 367.700 85.480 368.350 ;
        RECT 83.980 366.900 84.630 367.550 ;
        RECT 84.830 366.900 85.480 367.550 ;
        RECT 103.980 372.450 104.630 373.100 ;
        RECT 103.980 371.650 104.630 372.300 ;
        RECT 103.980 370.850 104.630 371.500 ;
        RECT 103.980 368.500 104.630 369.150 ;
        RECT 103.980 367.700 104.630 368.350 ;
        RECT 103.980 366.900 104.630 367.550 ;
        RECT 4.830 363.450 5.680 364.300 ;
        RECT 23.780 363.450 24.630 364.300 ;
        RECT 24.830 363.450 25.680 364.300 ;
        RECT 43.780 363.450 44.630 364.300 ;
        RECT 44.830 363.450 45.680 364.300 ;
        RECT 63.780 363.450 64.630 364.300 ;
        RECT 64.830 363.450 65.680 364.300 ;
        RECT 83.780 363.450 84.630 364.300 ;
        RECT 84.830 363.450 85.680 364.300 ;
        RECT 103.780 363.450 104.630 364.300 ;
        RECT 4.830 362.500 5.680 363.350 ;
        RECT 23.780 362.500 24.630 363.350 ;
        RECT 24.830 362.500 25.680 363.350 ;
        RECT 43.780 362.500 44.630 363.350 ;
        RECT 44.830 362.500 45.680 363.350 ;
        RECT 63.780 362.500 64.630 363.350 ;
        RECT 64.830 362.500 65.680 363.350 ;
        RECT 83.780 362.500 84.630 363.350 ;
        RECT 84.830 362.500 85.680 363.350 ;
        RECT 103.780 362.500 104.630 363.350 ;
        RECT 4.830 361.050 5.680 361.900 ;
        RECT 4.830 360.100 5.680 360.950 ;
        RECT 5.780 360.100 6.630 360.950 ;
        RECT 7.230 360.100 8.080 360.950 ;
        RECT 8.180 360.100 9.030 360.950 ;
        RECT 23.780 361.050 24.630 361.900 ;
        RECT 24.830 361.050 25.680 361.900 ;
        RECT 4.830 359.050 5.680 359.900 ;
        RECT 5.780 359.050 6.630 359.900 ;
        RECT 7.230 359.050 8.080 359.900 ;
        RECT 8.180 359.050 9.030 359.900 ;
        RECT 11.630 360.100 12.280 360.750 ;
        RECT 12.430 360.100 13.080 360.750 ;
        RECT 13.230 360.100 13.880 360.750 ;
        RECT 15.580 360.100 16.230 360.750 ;
        RECT 16.380 360.100 17.030 360.750 ;
        RECT 17.180 360.100 17.830 360.750 ;
        RECT 11.630 359.250 12.280 359.900 ;
        RECT 12.430 359.250 13.080 359.900 ;
        RECT 13.230 359.250 13.880 359.900 ;
        RECT 15.580 359.250 16.230 359.900 ;
        RECT 16.380 359.250 17.030 359.900 ;
        RECT 17.180 359.250 17.830 359.900 ;
        RECT 20.430 360.100 21.280 360.950 ;
        RECT 21.380 360.100 22.230 360.950 ;
        RECT 22.830 360.100 23.680 360.950 ;
        RECT 23.780 360.100 24.630 360.950 ;
        RECT 24.830 360.100 25.680 360.950 ;
        RECT 25.780 360.100 26.630 360.950 ;
        RECT 27.230 360.100 28.080 360.950 ;
        RECT 28.180 360.100 29.030 360.950 ;
        RECT 43.780 361.050 44.630 361.900 ;
        RECT 44.830 361.050 45.680 361.900 ;
        RECT 4.830 358.100 5.680 358.950 ;
        RECT 20.430 359.050 21.280 359.900 ;
        RECT 21.380 359.050 22.230 359.900 ;
        RECT 22.830 359.050 23.680 359.900 ;
        RECT 23.780 359.050 24.630 359.900 ;
        RECT 24.830 359.050 25.680 359.900 ;
        RECT 25.780 359.050 26.630 359.900 ;
        RECT 27.230 359.050 28.080 359.900 ;
        RECT 28.180 359.050 29.030 359.900 ;
        RECT 31.630 360.100 32.280 360.750 ;
        RECT 32.430 360.100 33.080 360.750 ;
        RECT 33.230 360.100 33.880 360.750 ;
        RECT 35.580 360.100 36.230 360.750 ;
        RECT 36.380 360.100 37.030 360.750 ;
        RECT 37.180 360.100 37.830 360.750 ;
        RECT 31.630 359.250 32.280 359.900 ;
        RECT 32.430 359.250 33.080 359.900 ;
        RECT 33.230 359.250 33.880 359.900 ;
        RECT 35.580 359.250 36.230 359.900 ;
        RECT 36.380 359.250 37.030 359.900 ;
        RECT 37.180 359.250 37.830 359.900 ;
        RECT 40.430 360.100 41.280 360.950 ;
        RECT 41.380 360.100 42.230 360.950 ;
        RECT 42.830 360.100 43.680 360.950 ;
        RECT 43.780 360.100 44.630 360.950 ;
        RECT 44.830 360.100 45.680 360.950 ;
        RECT 45.780 360.100 46.630 360.950 ;
        RECT 47.230 360.100 48.080 360.950 ;
        RECT 48.180 360.100 49.030 360.950 ;
        RECT 63.780 361.050 64.630 361.900 ;
        RECT 64.830 361.050 65.680 361.900 ;
        RECT 23.780 358.100 24.630 358.950 ;
        RECT 24.830 358.100 25.680 358.950 ;
        RECT 40.430 359.050 41.280 359.900 ;
        RECT 41.380 359.050 42.230 359.900 ;
        RECT 42.830 359.050 43.680 359.900 ;
        RECT 43.780 359.050 44.630 359.900 ;
        RECT 44.830 359.050 45.680 359.900 ;
        RECT 45.780 359.050 46.630 359.900 ;
        RECT 47.230 359.050 48.080 359.900 ;
        RECT 48.180 359.050 49.030 359.900 ;
        RECT 51.630 360.100 52.280 360.750 ;
        RECT 52.430 360.100 53.080 360.750 ;
        RECT 53.230 360.100 53.880 360.750 ;
        RECT 55.580 360.100 56.230 360.750 ;
        RECT 56.380 360.100 57.030 360.750 ;
        RECT 57.180 360.100 57.830 360.750 ;
        RECT 51.630 359.250 52.280 359.900 ;
        RECT 52.430 359.250 53.080 359.900 ;
        RECT 53.230 359.250 53.880 359.900 ;
        RECT 55.580 359.250 56.230 359.900 ;
        RECT 56.380 359.250 57.030 359.900 ;
        RECT 57.180 359.250 57.830 359.900 ;
        RECT 60.430 360.100 61.280 360.950 ;
        RECT 61.380 360.100 62.230 360.950 ;
        RECT 62.830 360.100 63.680 360.950 ;
        RECT 63.780 360.100 64.630 360.950 ;
        RECT 64.830 360.100 65.680 360.950 ;
        RECT 65.780 360.100 66.630 360.950 ;
        RECT 67.230 360.100 68.080 360.950 ;
        RECT 68.180 360.100 69.030 360.950 ;
        RECT 83.780 361.050 84.630 361.900 ;
        RECT 84.830 361.050 85.680 361.900 ;
        RECT 43.780 358.100 44.630 358.950 ;
        RECT 44.830 358.100 45.680 358.950 ;
        RECT 60.430 359.050 61.280 359.900 ;
        RECT 61.380 359.050 62.230 359.900 ;
        RECT 62.830 359.050 63.680 359.900 ;
        RECT 63.780 359.050 64.630 359.900 ;
        RECT 64.830 359.050 65.680 359.900 ;
        RECT 65.780 359.050 66.630 359.900 ;
        RECT 67.230 359.050 68.080 359.900 ;
        RECT 68.180 359.050 69.030 359.900 ;
        RECT 71.630 360.100 72.280 360.750 ;
        RECT 72.430 360.100 73.080 360.750 ;
        RECT 73.230 360.100 73.880 360.750 ;
        RECT 75.580 360.100 76.230 360.750 ;
        RECT 76.380 360.100 77.030 360.750 ;
        RECT 77.180 360.100 77.830 360.750 ;
        RECT 71.630 359.250 72.280 359.900 ;
        RECT 72.430 359.250 73.080 359.900 ;
        RECT 73.230 359.250 73.880 359.900 ;
        RECT 75.580 359.250 76.230 359.900 ;
        RECT 76.380 359.250 77.030 359.900 ;
        RECT 77.180 359.250 77.830 359.900 ;
        RECT 80.430 360.100 81.280 360.950 ;
        RECT 81.380 360.100 82.230 360.950 ;
        RECT 82.830 360.100 83.680 360.950 ;
        RECT 83.780 360.100 84.630 360.950 ;
        RECT 84.830 360.100 85.680 360.950 ;
        RECT 85.780 360.100 86.630 360.950 ;
        RECT 87.230 360.100 88.080 360.950 ;
        RECT 88.180 360.100 89.030 360.950 ;
        RECT 103.780 361.050 104.630 361.900 ;
        RECT 63.780 358.100 64.630 358.950 ;
        RECT 64.830 358.100 65.680 358.950 ;
        RECT 80.430 359.050 81.280 359.900 ;
        RECT 81.380 359.050 82.230 359.900 ;
        RECT 82.830 359.050 83.680 359.900 ;
        RECT 83.780 359.050 84.630 359.900 ;
        RECT 84.830 359.050 85.680 359.900 ;
        RECT 85.780 359.050 86.630 359.900 ;
        RECT 87.230 359.050 88.080 359.900 ;
        RECT 88.180 359.050 89.030 359.900 ;
        RECT 91.630 360.100 92.280 360.750 ;
        RECT 92.430 360.100 93.080 360.750 ;
        RECT 93.230 360.100 93.880 360.750 ;
        RECT 95.580 360.100 96.230 360.750 ;
        RECT 96.380 360.100 97.030 360.750 ;
        RECT 97.180 360.100 97.830 360.750 ;
        RECT 91.630 359.250 92.280 359.900 ;
        RECT 92.430 359.250 93.080 359.900 ;
        RECT 93.230 359.250 93.880 359.900 ;
        RECT 95.580 359.250 96.230 359.900 ;
        RECT 96.380 359.250 97.030 359.900 ;
        RECT 97.180 359.250 97.830 359.900 ;
        RECT 100.430 360.100 101.280 360.950 ;
        RECT 101.380 360.100 102.230 360.950 ;
        RECT 102.830 360.100 103.680 360.950 ;
        RECT 103.780 360.100 104.630 360.950 ;
        RECT 83.780 358.100 84.630 358.950 ;
        RECT 84.830 358.100 85.680 358.950 ;
        RECT 100.430 359.050 101.280 359.900 ;
        RECT 101.380 359.050 102.230 359.900 ;
        RECT 102.830 359.050 103.680 359.900 ;
        RECT 103.780 359.050 104.630 359.900 ;
        RECT 103.780 358.100 104.630 358.950 ;
        RECT 4.830 356.650 5.680 357.500 ;
        RECT 23.780 356.650 24.630 357.500 ;
        RECT 24.830 356.650 25.680 357.500 ;
        RECT 43.780 356.650 44.630 357.500 ;
        RECT 44.830 356.650 45.680 357.500 ;
        RECT 63.780 356.650 64.630 357.500 ;
        RECT 64.830 356.650 65.680 357.500 ;
        RECT 83.780 356.650 84.630 357.500 ;
        RECT 84.830 356.650 85.680 357.500 ;
        RECT 103.780 356.650 104.630 357.500 ;
        RECT 4.830 355.700 5.680 356.550 ;
        RECT 23.780 355.700 24.630 356.550 ;
        RECT 24.830 355.700 25.680 356.550 ;
        RECT 43.780 355.700 44.630 356.550 ;
        RECT 44.830 355.700 45.680 356.550 ;
        RECT 63.780 355.700 64.630 356.550 ;
        RECT 64.830 355.700 65.680 356.550 ;
        RECT 83.780 355.700 84.630 356.550 ;
        RECT 84.830 355.700 85.680 356.550 ;
        RECT 103.780 355.700 104.630 356.550 ;
        RECT 4.830 352.450 5.480 353.100 ;
        RECT 4.830 351.650 5.480 352.300 ;
        RECT 4.830 350.850 5.480 351.500 ;
        RECT 4.830 348.500 5.480 349.150 ;
        RECT 4.830 347.700 5.480 348.350 ;
        RECT 4.830 346.900 5.480 347.550 ;
        RECT 23.980 352.450 24.630 353.100 ;
        RECT 24.830 352.450 25.480 353.100 ;
        RECT 23.980 351.650 24.630 352.300 ;
        RECT 24.830 351.650 25.480 352.300 ;
        RECT 23.980 350.850 24.630 351.500 ;
        RECT 24.830 350.850 25.480 351.500 ;
        RECT 23.980 348.500 24.630 349.150 ;
        RECT 24.830 348.500 25.480 349.150 ;
        RECT 23.980 347.700 24.630 348.350 ;
        RECT 24.830 347.700 25.480 348.350 ;
        RECT 23.980 346.900 24.630 347.550 ;
        RECT 24.830 346.900 25.480 347.550 ;
        RECT 43.980 352.450 44.630 353.100 ;
        RECT 44.830 352.450 45.480 353.100 ;
        RECT 43.980 351.650 44.630 352.300 ;
        RECT 44.830 351.650 45.480 352.300 ;
        RECT 43.980 350.850 44.630 351.500 ;
        RECT 44.830 350.850 45.480 351.500 ;
        RECT 43.980 348.500 44.630 349.150 ;
        RECT 44.830 348.500 45.480 349.150 ;
        RECT 43.980 347.700 44.630 348.350 ;
        RECT 44.830 347.700 45.480 348.350 ;
        RECT 43.980 346.900 44.630 347.550 ;
        RECT 44.830 346.900 45.480 347.550 ;
        RECT 63.980 352.450 64.630 353.100 ;
        RECT 64.830 352.450 65.480 353.100 ;
        RECT 63.980 351.650 64.630 352.300 ;
        RECT 64.830 351.650 65.480 352.300 ;
        RECT 63.980 350.850 64.630 351.500 ;
        RECT 64.830 350.850 65.480 351.500 ;
        RECT 63.980 348.500 64.630 349.150 ;
        RECT 64.830 348.500 65.480 349.150 ;
        RECT 63.980 347.700 64.630 348.350 ;
        RECT 64.830 347.700 65.480 348.350 ;
        RECT 63.980 346.900 64.630 347.550 ;
        RECT 64.830 346.900 65.480 347.550 ;
        RECT 83.980 352.450 84.630 353.100 ;
        RECT 84.830 352.450 85.480 353.100 ;
        RECT 83.980 351.650 84.630 352.300 ;
        RECT 84.830 351.650 85.480 352.300 ;
        RECT 83.980 350.850 84.630 351.500 ;
        RECT 84.830 350.850 85.480 351.500 ;
        RECT 83.980 348.500 84.630 349.150 ;
        RECT 84.830 348.500 85.480 349.150 ;
        RECT 83.980 347.700 84.630 348.350 ;
        RECT 84.830 347.700 85.480 348.350 ;
        RECT 83.980 346.900 84.630 347.550 ;
        RECT 84.830 346.900 85.480 347.550 ;
        RECT 103.980 352.450 104.630 353.100 ;
        RECT 103.980 351.650 104.630 352.300 ;
        RECT 103.980 350.850 104.630 351.500 ;
        RECT 103.980 348.500 104.630 349.150 ;
        RECT 103.980 347.700 104.630 348.350 ;
        RECT 103.980 346.900 104.630 347.550 ;
        RECT 4.830 343.450 5.680 344.300 ;
        RECT 23.780 343.450 24.630 344.300 ;
        RECT 24.830 343.450 25.680 344.300 ;
        RECT 43.780 343.450 44.630 344.300 ;
        RECT 44.830 343.450 45.680 344.300 ;
        RECT 63.780 343.450 64.630 344.300 ;
        RECT 64.830 343.450 65.680 344.300 ;
        RECT 83.780 343.450 84.630 344.300 ;
        RECT 84.830 343.450 85.680 344.300 ;
        RECT 103.780 343.450 104.630 344.300 ;
        RECT 4.830 342.500 5.680 343.350 ;
        RECT 23.780 342.500 24.630 343.350 ;
        RECT 24.830 342.500 25.680 343.350 ;
        RECT 43.780 342.500 44.630 343.350 ;
        RECT 44.830 342.500 45.680 343.350 ;
        RECT 63.780 342.500 64.630 343.350 ;
        RECT 64.830 342.500 65.680 343.350 ;
        RECT 83.780 342.500 84.630 343.350 ;
        RECT 84.830 342.500 85.680 343.350 ;
        RECT 103.780 342.500 104.630 343.350 ;
        RECT 4.830 341.050 5.680 341.900 ;
        RECT 4.830 340.100 5.680 340.950 ;
        RECT 5.780 340.100 6.630 340.950 ;
        RECT 7.230 340.100 8.080 340.950 ;
        RECT 8.180 340.100 9.030 340.950 ;
        RECT 23.780 341.050 24.630 341.900 ;
        RECT 24.830 341.050 25.680 341.900 ;
        RECT 4.830 339.050 5.680 339.900 ;
        RECT 5.780 339.050 6.630 339.900 ;
        RECT 7.230 339.050 8.080 339.900 ;
        RECT 8.180 339.050 9.030 339.900 ;
        RECT 11.630 340.100 12.280 340.750 ;
        RECT 12.430 340.100 13.080 340.750 ;
        RECT 13.230 340.100 13.880 340.750 ;
        RECT 15.580 340.100 16.230 340.750 ;
        RECT 16.380 340.100 17.030 340.750 ;
        RECT 17.180 340.100 17.830 340.750 ;
        RECT 11.630 339.250 12.280 339.900 ;
        RECT 12.430 339.250 13.080 339.900 ;
        RECT 13.230 339.250 13.880 339.900 ;
        RECT 15.580 339.250 16.230 339.900 ;
        RECT 16.380 339.250 17.030 339.900 ;
        RECT 17.180 339.250 17.830 339.900 ;
        RECT 20.430 340.100 21.280 340.950 ;
        RECT 21.380 340.100 22.230 340.950 ;
        RECT 22.830 340.100 23.680 340.950 ;
        RECT 23.780 340.100 24.630 340.950 ;
        RECT 24.830 340.100 25.680 340.950 ;
        RECT 25.780 340.100 26.630 340.950 ;
        RECT 27.230 340.100 28.080 340.950 ;
        RECT 28.180 340.100 29.030 340.950 ;
        RECT 43.780 341.050 44.630 341.900 ;
        RECT 44.830 341.050 45.680 341.900 ;
        RECT 4.830 338.100 5.680 338.950 ;
        RECT 20.430 339.050 21.280 339.900 ;
        RECT 21.380 339.050 22.230 339.900 ;
        RECT 22.830 339.050 23.680 339.900 ;
        RECT 23.780 339.050 24.630 339.900 ;
        RECT 24.830 339.050 25.680 339.900 ;
        RECT 25.780 339.050 26.630 339.900 ;
        RECT 27.230 339.050 28.080 339.900 ;
        RECT 28.180 339.050 29.030 339.900 ;
        RECT 31.630 340.100 32.280 340.750 ;
        RECT 32.430 340.100 33.080 340.750 ;
        RECT 33.230 340.100 33.880 340.750 ;
        RECT 35.580 340.100 36.230 340.750 ;
        RECT 36.380 340.100 37.030 340.750 ;
        RECT 37.180 340.100 37.830 340.750 ;
        RECT 31.630 339.250 32.280 339.900 ;
        RECT 32.430 339.250 33.080 339.900 ;
        RECT 33.230 339.250 33.880 339.900 ;
        RECT 35.580 339.250 36.230 339.900 ;
        RECT 36.380 339.250 37.030 339.900 ;
        RECT 37.180 339.250 37.830 339.900 ;
        RECT 40.430 340.100 41.280 340.950 ;
        RECT 41.380 340.100 42.230 340.950 ;
        RECT 42.830 340.100 43.680 340.950 ;
        RECT 43.780 340.100 44.630 340.950 ;
        RECT 44.830 340.100 45.680 340.950 ;
        RECT 45.780 340.100 46.630 340.950 ;
        RECT 47.230 340.100 48.080 340.950 ;
        RECT 48.180 340.100 49.030 340.950 ;
        RECT 63.780 341.050 64.630 341.900 ;
        RECT 64.830 341.050 65.680 341.900 ;
        RECT 23.780 338.100 24.630 338.950 ;
        RECT 24.830 338.100 25.680 338.950 ;
        RECT 40.430 339.050 41.280 339.900 ;
        RECT 41.380 339.050 42.230 339.900 ;
        RECT 42.830 339.050 43.680 339.900 ;
        RECT 43.780 339.050 44.630 339.900 ;
        RECT 44.830 339.050 45.680 339.900 ;
        RECT 45.780 339.050 46.630 339.900 ;
        RECT 47.230 339.050 48.080 339.900 ;
        RECT 48.180 339.050 49.030 339.900 ;
        RECT 51.630 340.100 52.280 340.750 ;
        RECT 52.430 340.100 53.080 340.750 ;
        RECT 53.230 340.100 53.880 340.750 ;
        RECT 55.580 340.100 56.230 340.750 ;
        RECT 56.380 340.100 57.030 340.750 ;
        RECT 57.180 340.100 57.830 340.750 ;
        RECT 51.630 339.250 52.280 339.900 ;
        RECT 52.430 339.250 53.080 339.900 ;
        RECT 53.230 339.250 53.880 339.900 ;
        RECT 55.580 339.250 56.230 339.900 ;
        RECT 56.380 339.250 57.030 339.900 ;
        RECT 57.180 339.250 57.830 339.900 ;
        RECT 60.430 340.100 61.280 340.950 ;
        RECT 61.380 340.100 62.230 340.950 ;
        RECT 62.830 340.100 63.680 340.950 ;
        RECT 63.780 340.100 64.630 340.950 ;
        RECT 64.830 340.100 65.680 340.950 ;
        RECT 65.780 340.100 66.630 340.950 ;
        RECT 67.230 340.100 68.080 340.950 ;
        RECT 68.180 340.100 69.030 340.950 ;
        RECT 83.780 341.050 84.630 341.900 ;
        RECT 84.830 341.050 85.680 341.900 ;
        RECT 43.780 338.100 44.630 338.950 ;
        RECT 44.830 338.100 45.680 338.950 ;
        RECT 60.430 339.050 61.280 339.900 ;
        RECT 61.380 339.050 62.230 339.900 ;
        RECT 62.830 339.050 63.680 339.900 ;
        RECT 63.780 339.050 64.630 339.900 ;
        RECT 64.830 339.050 65.680 339.900 ;
        RECT 65.780 339.050 66.630 339.900 ;
        RECT 67.230 339.050 68.080 339.900 ;
        RECT 68.180 339.050 69.030 339.900 ;
        RECT 71.630 340.100 72.280 340.750 ;
        RECT 72.430 340.100 73.080 340.750 ;
        RECT 73.230 340.100 73.880 340.750 ;
        RECT 75.580 340.100 76.230 340.750 ;
        RECT 76.380 340.100 77.030 340.750 ;
        RECT 77.180 340.100 77.830 340.750 ;
        RECT 71.630 339.250 72.280 339.900 ;
        RECT 72.430 339.250 73.080 339.900 ;
        RECT 73.230 339.250 73.880 339.900 ;
        RECT 75.580 339.250 76.230 339.900 ;
        RECT 76.380 339.250 77.030 339.900 ;
        RECT 77.180 339.250 77.830 339.900 ;
        RECT 80.430 340.100 81.280 340.950 ;
        RECT 81.380 340.100 82.230 340.950 ;
        RECT 82.830 340.100 83.680 340.950 ;
        RECT 83.780 340.100 84.630 340.950 ;
        RECT 84.830 340.100 85.680 340.950 ;
        RECT 85.780 340.100 86.630 340.950 ;
        RECT 87.230 340.100 88.080 340.950 ;
        RECT 88.180 340.100 89.030 340.950 ;
        RECT 103.780 341.050 104.630 341.900 ;
        RECT 63.780 338.100 64.630 338.950 ;
        RECT 64.830 338.100 65.680 338.950 ;
        RECT 80.430 339.050 81.280 339.900 ;
        RECT 81.380 339.050 82.230 339.900 ;
        RECT 82.830 339.050 83.680 339.900 ;
        RECT 83.780 339.050 84.630 339.900 ;
        RECT 84.830 339.050 85.680 339.900 ;
        RECT 85.780 339.050 86.630 339.900 ;
        RECT 87.230 339.050 88.080 339.900 ;
        RECT 88.180 339.050 89.030 339.900 ;
        RECT 91.630 340.100 92.280 340.750 ;
        RECT 92.430 340.100 93.080 340.750 ;
        RECT 93.230 340.100 93.880 340.750 ;
        RECT 95.580 340.100 96.230 340.750 ;
        RECT 96.380 340.100 97.030 340.750 ;
        RECT 97.180 340.100 97.830 340.750 ;
        RECT 91.630 339.250 92.280 339.900 ;
        RECT 92.430 339.250 93.080 339.900 ;
        RECT 93.230 339.250 93.880 339.900 ;
        RECT 95.580 339.250 96.230 339.900 ;
        RECT 96.380 339.250 97.030 339.900 ;
        RECT 97.180 339.250 97.830 339.900 ;
        RECT 100.430 340.100 101.280 340.950 ;
        RECT 101.380 340.100 102.230 340.950 ;
        RECT 102.830 340.100 103.680 340.950 ;
        RECT 103.780 340.100 104.630 340.950 ;
        RECT 83.780 338.100 84.630 338.950 ;
        RECT 84.830 338.100 85.680 338.950 ;
        RECT 100.430 339.050 101.280 339.900 ;
        RECT 101.380 339.050 102.230 339.900 ;
        RECT 102.830 339.050 103.680 339.900 ;
        RECT 103.780 339.050 104.630 339.900 ;
        RECT 103.780 338.100 104.630 338.950 ;
        RECT 4.830 336.650 5.680 337.500 ;
        RECT 23.780 336.650 24.630 337.500 ;
        RECT 24.830 336.650 25.680 337.500 ;
        RECT 43.780 336.650 44.630 337.500 ;
        RECT 44.830 336.650 45.680 337.500 ;
        RECT 63.780 336.650 64.630 337.500 ;
        RECT 64.830 336.650 65.680 337.500 ;
        RECT 83.780 336.650 84.630 337.500 ;
        RECT 84.830 336.650 85.680 337.500 ;
        RECT 103.780 336.650 104.630 337.500 ;
        RECT 4.830 335.700 5.680 336.550 ;
        RECT 23.780 335.700 24.630 336.550 ;
        RECT 24.830 335.700 25.680 336.550 ;
        RECT 43.780 335.700 44.630 336.550 ;
        RECT 44.830 335.700 45.680 336.550 ;
        RECT 63.780 335.700 64.630 336.550 ;
        RECT 64.830 335.700 65.680 336.550 ;
        RECT 83.780 335.700 84.630 336.550 ;
        RECT 84.830 335.700 85.680 336.550 ;
        RECT 103.780 335.700 104.630 336.550 ;
        RECT 4.830 332.450 5.480 333.100 ;
        RECT 4.830 331.650 5.480 332.300 ;
        RECT 4.830 330.850 5.480 331.500 ;
        RECT 4.830 328.500 5.480 329.150 ;
        RECT 4.830 327.700 5.480 328.350 ;
        RECT 4.830 326.900 5.480 327.550 ;
        RECT 23.980 332.450 24.630 333.100 ;
        RECT 24.830 332.450 25.480 333.100 ;
        RECT 23.980 331.650 24.630 332.300 ;
        RECT 24.830 331.650 25.480 332.300 ;
        RECT 23.980 330.850 24.630 331.500 ;
        RECT 24.830 330.850 25.480 331.500 ;
        RECT 23.980 328.500 24.630 329.150 ;
        RECT 24.830 328.500 25.480 329.150 ;
        RECT 23.980 327.700 24.630 328.350 ;
        RECT 24.830 327.700 25.480 328.350 ;
        RECT 23.980 326.900 24.630 327.550 ;
        RECT 24.830 326.900 25.480 327.550 ;
        RECT 43.980 332.450 44.630 333.100 ;
        RECT 44.830 332.450 45.480 333.100 ;
        RECT 43.980 331.650 44.630 332.300 ;
        RECT 44.830 331.650 45.480 332.300 ;
        RECT 43.980 330.850 44.630 331.500 ;
        RECT 44.830 330.850 45.480 331.500 ;
        RECT 43.980 328.500 44.630 329.150 ;
        RECT 44.830 328.500 45.480 329.150 ;
        RECT 43.980 327.700 44.630 328.350 ;
        RECT 44.830 327.700 45.480 328.350 ;
        RECT 43.980 326.900 44.630 327.550 ;
        RECT 44.830 326.900 45.480 327.550 ;
        RECT 63.980 332.450 64.630 333.100 ;
        RECT 64.830 332.450 65.480 333.100 ;
        RECT 63.980 331.650 64.630 332.300 ;
        RECT 64.830 331.650 65.480 332.300 ;
        RECT 63.980 330.850 64.630 331.500 ;
        RECT 64.830 330.850 65.480 331.500 ;
        RECT 63.980 328.500 64.630 329.150 ;
        RECT 64.830 328.500 65.480 329.150 ;
        RECT 63.980 327.700 64.630 328.350 ;
        RECT 64.830 327.700 65.480 328.350 ;
        RECT 63.980 326.900 64.630 327.550 ;
        RECT 64.830 326.900 65.480 327.550 ;
        RECT 83.980 332.450 84.630 333.100 ;
        RECT 84.830 332.450 85.480 333.100 ;
        RECT 83.980 331.650 84.630 332.300 ;
        RECT 84.830 331.650 85.480 332.300 ;
        RECT 83.980 330.850 84.630 331.500 ;
        RECT 84.830 330.850 85.480 331.500 ;
        RECT 83.980 328.500 84.630 329.150 ;
        RECT 84.830 328.500 85.480 329.150 ;
        RECT 83.980 327.700 84.630 328.350 ;
        RECT 84.830 327.700 85.480 328.350 ;
        RECT 83.980 326.900 84.630 327.550 ;
        RECT 84.830 326.900 85.480 327.550 ;
        RECT 103.980 332.450 104.630 333.100 ;
        RECT 103.980 331.650 104.630 332.300 ;
        RECT 103.980 330.850 104.630 331.500 ;
        RECT 103.980 328.500 104.630 329.150 ;
        RECT 103.980 327.700 104.630 328.350 ;
        RECT 103.980 326.900 104.630 327.550 ;
        RECT 4.830 323.450 5.680 324.300 ;
        RECT 23.780 323.450 24.630 324.300 ;
        RECT 24.830 323.450 25.680 324.300 ;
        RECT 43.780 323.450 44.630 324.300 ;
        RECT 44.830 323.450 45.680 324.300 ;
        RECT 63.780 323.450 64.630 324.300 ;
        RECT 64.830 323.450 65.680 324.300 ;
        RECT 83.780 323.450 84.630 324.300 ;
        RECT 84.830 323.450 85.680 324.300 ;
        RECT 103.780 323.450 104.630 324.300 ;
        RECT 4.830 322.500 5.680 323.350 ;
        RECT 23.780 322.500 24.630 323.350 ;
        RECT 24.830 322.500 25.680 323.350 ;
        RECT 43.780 322.500 44.630 323.350 ;
        RECT 44.830 322.500 45.680 323.350 ;
        RECT 63.780 322.500 64.630 323.350 ;
        RECT 64.830 322.500 65.680 323.350 ;
        RECT 83.780 322.500 84.630 323.350 ;
        RECT 84.830 322.500 85.680 323.350 ;
        RECT 103.780 322.500 104.630 323.350 ;
        RECT 4.830 321.050 5.680 321.900 ;
        RECT 4.830 320.100 5.680 320.950 ;
        RECT 5.780 320.100 6.630 320.950 ;
        RECT 7.230 320.100 8.080 320.950 ;
        RECT 8.180 320.100 9.030 320.950 ;
        RECT 23.780 321.050 24.630 321.900 ;
        RECT 24.830 321.050 25.680 321.900 ;
        RECT 4.830 319.050 5.680 319.900 ;
        RECT 5.780 319.050 6.630 319.900 ;
        RECT 7.230 319.050 8.080 319.900 ;
        RECT 8.180 319.050 9.030 319.900 ;
        RECT 11.630 320.100 12.280 320.750 ;
        RECT 12.430 320.100 13.080 320.750 ;
        RECT 13.230 320.100 13.880 320.750 ;
        RECT 15.580 320.100 16.230 320.750 ;
        RECT 16.380 320.100 17.030 320.750 ;
        RECT 17.180 320.100 17.830 320.750 ;
        RECT 11.630 319.250 12.280 319.900 ;
        RECT 12.430 319.250 13.080 319.900 ;
        RECT 13.230 319.250 13.880 319.900 ;
        RECT 15.580 319.250 16.230 319.900 ;
        RECT 16.380 319.250 17.030 319.900 ;
        RECT 17.180 319.250 17.830 319.900 ;
        RECT 20.430 320.100 21.280 320.950 ;
        RECT 21.380 320.100 22.230 320.950 ;
        RECT 22.830 320.100 23.680 320.950 ;
        RECT 23.780 320.100 24.630 320.950 ;
        RECT 24.830 320.100 25.680 320.950 ;
        RECT 25.780 320.100 26.630 320.950 ;
        RECT 27.230 320.100 28.080 320.950 ;
        RECT 28.180 320.100 29.030 320.950 ;
        RECT 43.780 321.050 44.630 321.900 ;
        RECT 44.830 321.050 45.680 321.900 ;
        RECT 4.830 318.100 5.680 318.950 ;
        RECT 20.430 319.050 21.280 319.900 ;
        RECT 21.380 319.050 22.230 319.900 ;
        RECT 22.830 319.050 23.680 319.900 ;
        RECT 23.780 319.050 24.630 319.900 ;
        RECT 24.830 319.050 25.680 319.900 ;
        RECT 25.780 319.050 26.630 319.900 ;
        RECT 27.230 319.050 28.080 319.900 ;
        RECT 28.180 319.050 29.030 319.900 ;
        RECT 31.630 320.100 32.280 320.750 ;
        RECT 32.430 320.100 33.080 320.750 ;
        RECT 33.230 320.100 33.880 320.750 ;
        RECT 35.580 320.100 36.230 320.750 ;
        RECT 36.380 320.100 37.030 320.750 ;
        RECT 37.180 320.100 37.830 320.750 ;
        RECT 31.630 319.250 32.280 319.900 ;
        RECT 32.430 319.250 33.080 319.900 ;
        RECT 33.230 319.250 33.880 319.900 ;
        RECT 35.580 319.250 36.230 319.900 ;
        RECT 36.380 319.250 37.030 319.900 ;
        RECT 37.180 319.250 37.830 319.900 ;
        RECT 40.430 320.100 41.280 320.950 ;
        RECT 41.380 320.100 42.230 320.950 ;
        RECT 42.830 320.100 43.680 320.950 ;
        RECT 43.780 320.100 44.630 320.950 ;
        RECT 44.830 320.100 45.680 320.950 ;
        RECT 45.780 320.100 46.630 320.950 ;
        RECT 47.230 320.100 48.080 320.950 ;
        RECT 48.180 320.100 49.030 320.950 ;
        RECT 63.780 321.050 64.630 321.900 ;
        RECT 64.830 321.050 65.680 321.900 ;
        RECT 23.780 318.100 24.630 318.950 ;
        RECT 24.830 318.100 25.680 318.950 ;
        RECT 40.430 319.050 41.280 319.900 ;
        RECT 41.380 319.050 42.230 319.900 ;
        RECT 42.830 319.050 43.680 319.900 ;
        RECT 43.780 319.050 44.630 319.900 ;
        RECT 44.830 319.050 45.680 319.900 ;
        RECT 45.780 319.050 46.630 319.900 ;
        RECT 47.230 319.050 48.080 319.900 ;
        RECT 48.180 319.050 49.030 319.900 ;
        RECT 51.630 320.100 52.280 320.750 ;
        RECT 52.430 320.100 53.080 320.750 ;
        RECT 53.230 320.100 53.880 320.750 ;
        RECT 55.580 320.100 56.230 320.750 ;
        RECT 56.380 320.100 57.030 320.750 ;
        RECT 57.180 320.100 57.830 320.750 ;
        RECT 51.630 319.250 52.280 319.900 ;
        RECT 52.430 319.250 53.080 319.900 ;
        RECT 53.230 319.250 53.880 319.900 ;
        RECT 55.580 319.250 56.230 319.900 ;
        RECT 56.380 319.250 57.030 319.900 ;
        RECT 57.180 319.250 57.830 319.900 ;
        RECT 60.430 320.100 61.280 320.950 ;
        RECT 61.380 320.100 62.230 320.950 ;
        RECT 62.830 320.100 63.680 320.950 ;
        RECT 63.780 320.100 64.630 320.950 ;
        RECT 64.830 320.100 65.680 320.950 ;
        RECT 65.780 320.100 66.630 320.950 ;
        RECT 67.230 320.100 68.080 320.950 ;
        RECT 68.180 320.100 69.030 320.950 ;
        RECT 83.780 321.050 84.630 321.900 ;
        RECT 84.830 321.050 85.680 321.900 ;
        RECT 43.780 318.100 44.630 318.950 ;
        RECT 44.830 318.100 45.680 318.950 ;
        RECT 60.430 319.050 61.280 319.900 ;
        RECT 61.380 319.050 62.230 319.900 ;
        RECT 62.830 319.050 63.680 319.900 ;
        RECT 63.780 319.050 64.630 319.900 ;
        RECT 64.830 319.050 65.680 319.900 ;
        RECT 65.780 319.050 66.630 319.900 ;
        RECT 67.230 319.050 68.080 319.900 ;
        RECT 68.180 319.050 69.030 319.900 ;
        RECT 71.630 320.100 72.280 320.750 ;
        RECT 72.430 320.100 73.080 320.750 ;
        RECT 73.230 320.100 73.880 320.750 ;
        RECT 75.580 320.100 76.230 320.750 ;
        RECT 76.380 320.100 77.030 320.750 ;
        RECT 77.180 320.100 77.830 320.750 ;
        RECT 71.630 319.250 72.280 319.900 ;
        RECT 72.430 319.250 73.080 319.900 ;
        RECT 73.230 319.250 73.880 319.900 ;
        RECT 75.580 319.250 76.230 319.900 ;
        RECT 76.380 319.250 77.030 319.900 ;
        RECT 77.180 319.250 77.830 319.900 ;
        RECT 80.430 320.100 81.280 320.950 ;
        RECT 81.380 320.100 82.230 320.950 ;
        RECT 82.830 320.100 83.680 320.950 ;
        RECT 83.780 320.100 84.630 320.950 ;
        RECT 84.830 320.100 85.680 320.950 ;
        RECT 85.780 320.100 86.630 320.950 ;
        RECT 87.230 320.100 88.080 320.950 ;
        RECT 88.180 320.100 89.030 320.950 ;
        RECT 103.780 321.050 104.630 321.900 ;
        RECT 63.780 318.100 64.630 318.950 ;
        RECT 64.830 318.100 65.680 318.950 ;
        RECT 80.430 319.050 81.280 319.900 ;
        RECT 81.380 319.050 82.230 319.900 ;
        RECT 82.830 319.050 83.680 319.900 ;
        RECT 83.780 319.050 84.630 319.900 ;
        RECT 84.830 319.050 85.680 319.900 ;
        RECT 85.780 319.050 86.630 319.900 ;
        RECT 87.230 319.050 88.080 319.900 ;
        RECT 88.180 319.050 89.030 319.900 ;
        RECT 91.630 320.100 92.280 320.750 ;
        RECT 92.430 320.100 93.080 320.750 ;
        RECT 93.230 320.100 93.880 320.750 ;
        RECT 95.580 320.100 96.230 320.750 ;
        RECT 96.380 320.100 97.030 320.750 ;
        RECT 97.180 320.100 97.830 320.750 ;
        RECT 91.630 319.250 92.280 319.900 ;
        RECT 92.430 319.250 93.080 319.900 ;
        RECT 93.230 319.250 93.880 319.900 ;
        RECT 95.580 319.250 96.230 319.900 ;
        RECT 96.380 319.250 97.030 319.900 ;
        RECT 97.180 319.250 97.830 319.900 ;
        RECT 100.430 320.100 101.280 320.950 ;
        RECT 101.380 320.100 102.230 320.950 ;
        RECT 102.830 320.100 103.680 320.950 ;
        RECT 103.780 320.100 104.630 320.950 ;
        RECT 83.780 318.100 84.630 318.950 ;
        RECT 84.830 318.100 85.680 318.950 ;
        RECT 100.430 319.050 101.280 319.900 ;
        RECT 101.380 319.050 102.230 319.900 ;
        RECT 102.830 319.050 103.680 319.900 ;
        RECT 103.780 319.050 104.630 319.900 ;
        RECT 103.780 318.100 104.630 318.950 ;
        RECT 4.830 316.650 5.680 317.500 ;
        RECT 23.780 316.650 24.630 317.500 ;
        RECT 24.830 316.650 25.680 317.500 ;
        RECT 43.780 316.650 44.630 317.500 ;
        RECT 44.830 316.650 45.680 317.500 ;
        RECT 63.780 316.650 64.630 317.500 ;
        RECT 64.830 316.650 65.680 317.500 ;
        RECT 83.780 316.650 84.630 317.500 ;
        RECT 84.830 316.650 85.680 317.500 ;
        RECT 103.780 316.650 104.630 317.500 ;
        RECT 4.830 315.700 5.680 316.550 ;
        RECT 23.780 315.700 24.630 316.550 ;
        RECT 24.830 315.700 25.680 316.550 ;
        RECT 43.780 315.700 44.630 316.550 ;
        RECT 44.830 315.700 45.680 316.550 ;
        RECT 63.780 315.700 64.630 316.550 ;
        RECT 64.830 315.700 65.680 316.550 ;
        RECT 83.780 315.700 84.630 316.550 ;
        RECT 84.830 315.700 85.680 316.550 ;
        RECT 103.780 315.700 104.630 316.550 ;
        RECT 4.830 312.450 5.480 313.100 ;
        RECT 4.830 311.650 5.480 312.300 ;
        RECT 4.830 310.850 5.480 311.500 ;
        RECT 4.830 308.500 5.480 309.150 ;
        RECT 4.830 307.700 5.480 308.350 ;
        RECT 4.830 306.900 5.480 307.550 ;
        RECT 23.980 312.450 24.630 313.100 ;
        RECT 24.830 312.450 25.480 313.100 ;
        RECT 23.980 311.650 24.630 312.300 ;
        RECT 24.830 311.650 25.480 312.300 ;
        RECT 23.980 310.850 24.630 311.500 ;
        RECT 24.830 310.850 25.480 311.500 ;
        RECT 23.980 308.500 24.630 309.150 ;
        RECT 24.830 308.500 25.480 309.150 ;
        RECT 23.980 307.700 24.630 308.350 ;
        RECT 24.830 307.700 25.480 308.350 ;
        RECT 23.980 306.900 24.630 307.550 ;
        RECT 24.830 306.900 25.480 307.550 ;
        RECT 43.980 312.450 44.630 313.100 ;
        RECT 44.830 312.450 45.480 313.100 ;
        RECT 43.980 311.650 44.630 312.300 ;
        RECT 44.830 311.650 45.480 312.300 ;
        RECT 43.980 310.850 44.630 311.500 ;
        RECT 44.830 310.850 45.480 311.500 ;
        RECT 43.980 308.500 44.630 309.150 ;
        RECT 44.830 308.500 45.480 309.150 ;
        RECT 43.980 307.700 44.630 308.350 ;
        RECT 44.830 307.700 45.480 308.350 ;
        RECT 43.980 306.900 44.630 307.550 ;
        RECT 44.830 306.900 45.480 307.550 ;
        RECT 63.980 312.450 64.630 313.100 ;
        RECT 64.830 312.450 65.480 313.100 ;
        RECT 63.980 311.650 64.630 312.300 ;
        RECT 64.830 311.650 65.480 312.300 ;
        RECT 63.980 310.850 64.630 311.500 ;
        RECT 64.830 310.850 65.480 311.500 ;
        RECT 63.980 308.500 64.630 309.150 ;
        RECT 64.830 308.500 65.480 309.150 ;
        RECT 63.980 307.700 64.630 308.350 ;
        RECT 64.830 307.700 65.480 308.350 ;
        RECT 63.980 306.900 64.630 307.550 ;
        RECT 64.830 306.900 65.480 307.550 ;
        RECT 83.980 312.450 84.630 313.100 ;
        RECT 84.830 312.450 85.480 313.100 ;
        RECT 83.980 311.650 84.630 312.300 ;
        RECT 84.830 311.650 85.480 312.300 ;
        RECT 83.980 310.850 84.630 311.500 ;
        RECT 84.830 310.850 85.480 311.500 ;
        RECT 83.980 308.500 84.630 309.150 ;
        RECT 84.830 308.500 85.480 309.150 ;
        RECT 83.980 307.700 84.630 308.350 ;
        RECT 84.830 307.700 85.480 308.350 ;
        RECT 83.980 306.900 84.630 307.550 ;
        RECT 84.830 306.900 85.480 307.550 ;
        RECT 103.980 312.450 104.630 313.100 ;
        RECT 103.980 311.650 104.630 312.300 ;
        RECT 103.980 310.850 104.630 311.500 ;
        RECT 103.980 308.500 104.630 309.150 ;
        RECT 103.980 307.700 104.630 308.350 ;
        RECT 103.980 306.900 104.630 307.550 ;
        RECT 4.830 303.450 5.680 304.300 ;
        RECT 23.780 303.450 24.630 304.300 ;
        RECT 24.830 303.450 25.680 304.300 ;
        RECT 43.780 303.450 44.630 304.300 ;
        RECT 44.830 303.450 45.680 304.300 ;
        RECT 63.780 303.450 64.630 304.300 ;
        RECT 64.830 303.450 65.680 304.300 ;
        RECT 83.780 303.450 84.630 304.300 ;
        RECT 84.830 303.450 85.680 304.300 ;
        RECT 103.780 303.450 104.630 304.300 ;
        RECT 4.830 302.500 5.680 303.350 ;
        RECT 23.780 302.500 24.630 303.350 ;
        RECT 24.830 302.500 25.680 303.350 ;
        RECT 43.780 302.500 44.630 303.350 ;
        RECT 44.830 302.500 45.680 303.350 ;
        RECT 63.780 302.500 64.630 303.350 ;
        RECT 64.830 302.500 65.680 303.350 ;
        RECT 83.780 302.500 84.630 303.350 ;
        RECT 84.830 302.500 85.680 303.350 ;
        RECT 103.780 302.500 104.630 303.350 ;
        RECT 4.830 301.050 5.680 301.900 ;
        RECT 4.830 300.100 5.680 300.950 ;
        RECT 5.780 300.100 6.630 300.950 ;
        RECT 7.230 300.100 8.080 300.950 ;
        RECT 8.180 300.100 9.030 300.950 ;
        RECT 23.780 301.050 24.630 301.900 ;
        RECT 24.830 301.050 25.680 301.900 ;
        RECT 4.830 299.050 5.680 299.900 ;
        RECT 5.780 299.050 6.630 299.900 ;
        RECT 7.230 299.050 8.080 299.900 ;
        RECT 8.180 299.050 9.030 299.900 ;
        RECT 11.630 300.100 12.280 300.750 ;
        RECT 12.430 300.100 13.080 300.750 ;
        RECT 13.230 300.100 13.880 300.750 ;
        RECT 15.580 300.100 16.230 300.750 ;
        RECT 16.380 300.100 17.030 300.750 ;
        RECT 17.180 300.100 17.830 300.750 ;
        RECT 11.630 299.250 12.280 299.900 ;
        RECT 12.430 299.250 13.080 299.900 ;
        RECT 13.230 299.250 13.880 299.900 ;
        RECT 15.580 299.250 16.230 299.900 ;
        RECT 16.380 299.250 17.030 299.900 ;
        RECT 17.180 299.250 17.830 299.900 ;
        RECT 20.430 300.100 21.280 300.950 ;
        RECT 21.380 300.100 22.230 300.950 ;
        RECT 22.830 300.100 23.680 300.950 ;
        RECT 23.780 300.100 24.630 300.950 ;
        RECT 24.830 300.100 25.680 300.950 ;
        RECT 25.780 300.100 26.630 300.950 ;
        RECT 27.230 300.100 28.080 300.950 ;
        RECT 28.180 300.100 29.030 300.950 ;
        RECT 43.780 301.050 44.630 301.900 ;
        RECT 44.830 301.050 45.680 301.900 ;
        RECT 4.830 298.100 5.680 298.950 ;
        RECT 20.430 299.050 21.280 299.900 ;
        RECT 21.380 299.050 22.230 299.900 ;
        RECT 22.830 299.050 23.680 299.900 ;
        RECT 23.780 299.050 24.630 299.900 ;
        RECT 24.830 299.050 25.680 299.900 ;
        RECT 25.780 299.050 26.630 299.900 ;
        RECT 27.230 299.050 28.080 299.900 ;
        RECT 28.180 299.050 29.030 299.900 ;
        RECT 31.630 300.100 32.280 300.750 ;
        RECT 32.430 300.100 33.080 300.750 ;
        RECT 33.230 300.100 33.880 300.750 ;
        RECT 35.580 300.100 36.230 300.750 ;
        RECT 36.380 300.100 37.030 300.750 ;
        RECT 37.180 300.100 37.830 300.750 ;
        RECT 31.630 299.250 32.280 299.900 ;
        RECT 32.430 299.250 33.080 299.900 ;
        RECT 33.230 299.250 33.880 299.900 ;
        RECT 35.580 299.250 36.230 299.900 ;
        RECT 36.380 299.250 37.030 299.900 ;
        RECT 37.180 299.250 37.830 299.900 ;
        RECT 40.430 300.100 41.280 300.950 ;
        RECT 41.380 300.100 42.230 300.950 ;
        RECT 42.830 300.100 43.680 300.950 ;
        RECT 43.780 300.100 44.630 300.950 ;
        RECT 44.830 300.100 45.680 300.950 ;
        RECT 45.780 300.100 46.630 300.950 ;
        RECT 47.230 300.100 48.080 300.950 ;
        RECT 48.180 300.100 49.030 300.950 ;
        RECT 63.780 301.050 64.630 301.900 ;
        RECT 64.830 301.050 65.680 301.900 ;
        RECT 23.780 298.100 24.630 298.950 ;
        RECT 24.830 298.100 25.680 298.950 ;
        RECT 40.430 299.050 41.280 299.900 ;
        RECT 41.380 299.050 42.230 299.900 ;
        RECT 42.830 299.050 43.680 299.900 ;
        RECT 43.780 299.050 44.630 299.900 ;
        RECT 44.830 299.050 45.680 299.900 ;
        RECT 45.780 299.050 46.630 299.900 ;
        RECT 47.230 299.050 48.080 299.900 ;
        RECT 48.180 299.050 49.030 299.900 ;
        RECT 51.630 300.100 52.280 300.750 ;
        RECT 52.430 300.100 53.080 300.750 ;
        RECT 53.230 300.100 53.880 300.750 ;
        RECT 55.580 300.100 56.230 300.750 ;
        RECT 56.380 300.100 57.030 300.750 ;
        RECT 57.180 300.100 57.830 300.750 ;
        RECT 51.630 299.250 52.280 299.900 ;
        RECT 52.430 299.250 53.080 299.900 ;
        RECT 53.230 299.250 53.880 299.900 ;
        RECT 55.580 299.250 56.230 299.900 ;
        RECT 56.380 299.250 57.030 299.900 ;
        RECT 57.180 299.250 57.830 299.900 ;
        RECT 60.430 300.100 61.280 300.950 ;
        RECT 61.380 300.100 62.230 300.950 ;
        RECT 62.830 300.100 63.680 300.950 ;
        RECT 63.780 300.100 64.630 300.950 ;
        RECT 64.830 300.100 65.680 300.950 ;
        RECT 65.780 300.100 66.630 300.950 ;
        RECT 67.230 300.100 68.080 300.950 ;
        RECT 68.180 300.100 69.030 300.950 ;
        RECT 83.780 301.050 84.630 301.900 ;
        RECT 84.830 301.050 85.680 301.900 ;
        RECT 43.780 298.100 44.630 298.950 ;
        RECT 44.830 298.100 45.680 298.950 ;
        RECT 60.430 299.050 61.280 299.900 ;
        RECT 61.380 299.050 62.230 299.900 ;
        RECT 62.830 299.050 63.680 299.900 ;
        RECT 63.780 299.050 64.630 299.900 ;
        RECT 64.830 299.050 65.680 299.900 ;
        RECT 65.780 299.050 66.630 299.900 ;
        RECT 67.230 299.050 68.080 299.900 ;
        RECT 68.180 299.050 69.030 299.900 ;
        RECT 71.630 300.100 72.280 300.750 ;
        RECT 72.430 300.100 73.080 300.750 ;
        RECT 73.230 300.100 73.880 300.750 ;
        RECT 75.580 300.100 76.230 300.750 ;
        RECT 76.380 300.100 77.030 300.750 ;
        RECT 77.180 300.100 77.830 300.750 ;
        RECT 71.630 299.250 72.280 299.900 ;
        RECT 72.430 299.250 73.080 299.900 ;
        RECT 73.230 299.250 73.880 299.900 ;
        RECT 75.580 299.250 76.230 299.900 ;
        RECT 76.380 299.250 77.030 299.900 ;
        RECT 77.180 299.250 77.830 299.900 ;
        RECT 80.430 300.100 81.280 300.950 ;
        RECT 81.380 300.100 82.230 300.950 ;
        RECT 82.830 300.100 83.680 300.950 ;
        RECT 83.780 300.100 84.630 300.950 ;
        RECT 84.830 300.100 85.680 300.950 ;
        RECT 85.780 300.100 86.630 300.950 ;
        RECT 87.230 300.100 88.080 300.950 ;
        RECT 88.180 300.100 89.030 300.950 ;
        RECT 103.780 301.050 104.630 301.900 ;
        RECT 63.780 298.100 64.630 298.950 ;
        RECT 64.830 298.100 65.680 298.950 ;
        RECT 80.430 299.050 81.280 299.900 ;
        RECT 81.380 299.050 82.230 299.900 ;
        RECT 82.830 299.050 83.680 299.900 ;
        RECT 83.780 299.050 84.630 299.900 ;
        RECT 84.830 299.050 85.680 299.900 ;
        RECT 85.780 299.050 86.630 299.900 ;
        RECT 87.230 299.050 88.080 299.900 ;
        RECT 88.180 299.050 89.030 299.900 ;
        RECT 91.630 300.100 92.280 300.750 ;
        RECT 92.430 300.100 93.080 300.750 ;
        RECT 93.230 300.100 93.880 300.750 ;
        RECT 95.580 300.100 96.230 300.750 ;
        RECT 96.380 300.100 97.030 300.750 ;
        RECT 97.180 300.100 97.830 300.750 ;
        RECT 91.630 299.250 92.280 299.900 ;
        RECT 92.430 299.250 93.080 299.900 ;
        RECT 93.230 299.250 93.880 299.900 ;
        RECT 95.580 299.250 96.230 299.900 ;
        RECT 96.380 299.250 97.030 299.900 ;
        RECT 97.180 299.250 97.830 299.900 ;
        RECT 100.430 300.100 101.280 300.950 ;
        RECT 101.380 300.100 102.230 300.950 ;
        RECT 102.830 300.100 103.680 300.950 ;
        RECT 103.780 300.100 104.630 300.950 ;
        RECT 83.780 298.100 84.630 298.950 ;
        RECT 84.830 298.100 85.680 298.950 ;
        RECT 100.430 299.050 101.280 299.900 ;
        RECT 101.380 299.050 102.230 299.900 ;
        RECT 102.830 299.050 103.680 299.900 ;
        RECT 103.780 299.050 104.630 299.900 ;
        RECT 103.780 298.100 104.630 298.950 ;
        RECT 4.830 296.650 5.680 297.500 ;
        RECT 23.780 296.650 24.630 297.500 ;
        RECT 24.830 296.650 25.680 297.500 ;
        RECT 43.780 296.650 44.630 297.500 ;
        RECT 44.830 296.650 45.680 297.500 ;
        RECT 63.780 296.650 64.630 297.500 ;
        RECT 64.830 296.650 65.680 297.500 ;
        RECT 83.780 296.650 84.630 297.500 ;
        RECT 84.830 296.650 85.680 297.500 ;
        RECT 103.780 296.650 104.630 297.500 ;
        RECT 4.830 295.700 5.680 296.550 ;
        RECT 23.780 295.700 24.630 296.550 ;
        RECT 24.830 295.700 25.680 296.550 ;
        RECT 43.780 295.700 44.630 296.550 ;
        RECT 44.830 295.700 45.680 296.550 ;
        RECT 63.780 295.700 64.630 296.550 ;
        RECT 64.830 295.700 65.680 296.550 ;
        RECT 83.780 295.700 84.630 296.550 ;
        RECT 84.830 295.700 85.680 296.550 ;
        RECT 103.780 295.700 104.630 296.550 ;
        RECT 4.830 292.450 5.480 293.100 ;
        RECT 4.830 291.650 5.480 292.300 ;
        RECT 4.830 290.850 5.480 291.500 ;
        RECT 4.830 288.500 5.480 289.150 ;
        RECT 4.830 287.700 5.480 288.350 ;
        RECT 4.830 286.900 5.480 287.550 ;
        RECT 23.980 292.450 24.630 293.100 ;
        RECT 24.830 292.450 25.480 293.100 ;
        RECT 23.980 291.650 24.630 292.300 ;
        RECT 24.830 291.650 25.480 292.300 ;
        RECT 23.980 290.850 24.630 291.500 ;
        RECT 24.830 290.850 25.480 291.500 ;
        RECT 23.980 288.500 24.630 289.150 ;
        RECT 24.830 288.500 25.480 289.150 ;
        RECT 23.980 287.700 24.630 288.350 ;
        RECT 24.830 287.700 25.480 288.350 ;
        RECT 23.980 286.900 24.630 287.550 ;
        RECT 24.830 286.900 25.480 287.550 ;
        RECT 43.980 292.450 44.630 293.100 ;
        RECT 44.830 292.450 45.480 293.100 ;
        RECT 43.980 291.650 44.630 292.300 ;
        RECT 44.830 291.650 45.480 292.300 ;
        RECT 43.980 290.850 44.630 291.500 ;
        RECT 44.830 290.850 45.480 291.500 ;
        RECT 43.980 288.500 44.630 289.150 ;
        RECT 44.830 288.500 45.480 289.150 ;
        RECT 43.980 287.700 44.630 288.350 ;
        RECT 44.830 287.700 45.480 288.350 ;
        RECT 43.980 286.900 44.630 287.550 ;
        RECT 44.830 286.900 45.480 287.550 ;
        RECT 63.980 292.450 64.630 293.100 ;
        RECT 64.830 292.450 65.480 293.100 ;
        RECT 63.980 291.650 64.630 292.300 ;
        RECT 64.830 291.650 65.480 292.300 ;
        RECT 63.980 290.850 64.630 291.500 ;
        RECT 64.830 290.850 65.480 291.500 ;
        RECT 63.980 288.500 64.630 289.150 ;
        RECT 64.830 288.500 65.480 289.150 ;
        RECT 63.980 287.700 64.630 288.350 ;
        RECT 64.830 287.700 65.480 288.350 ;
        RECT 63.980 286.900 64.630 287.550 ;
        RECT 64.830 286.900 65.480 287.550 ;
        RECT 83.980 292.450 84.630 293.100 ;
        RECT 84.830 292.450 85.480 293.100 ;
        RECT 83.980 291.650 84.630 292.300 ;
        RECT 84.830 291.650 85.480 292.300 ;
        RECT 83.980 290.850 84.630 291.500 ;
        RECT 84.830 290.850 85.480 291.500 ;
        RECT 83.980 288.500 84.630 289.150 ;
        RECT 84.830 288.500 85.480 289.150 ;
        RECT 83.980 287.700 84.630 288.350 ;
        RECT 84.830 287.700 85.480 288.350 ;
        RECT 83.980 286.900 84.630 287.550 ;
        RECT 84.830 286.900 85.480 287.550 ;
        RECT 103.980 292.450 104.630 293.100 ;
        RECT 103.980 291.650 104.630 292.300 ;
        RECT 103.980 290.850 104.630 291.500 ;
        RECT 103.980 288.500 104.630 289.150 ;
        RECT 103.980 287.700 104.630 288.350 ;
        RECT 103.980 286.900 104.630 287.550 ;
        RECT 4.830 283.450 5.680 284.300 ;
        RECT 23.780 283.450 24.630 284.300 ;
        RECT 24.830 283.450 25.680 284.300 ;
        RECT 43.780 283.450 44.630 284.300 ;
        RECT 44.830 283.450 45.680 284.300 ;
        RECT 63.780 283.450 64.630 284.300 ;
        RECT 64.830 283.450 65.680 284.300 ;
        RECT 83.780 283.450 84.630 284.300 ;
        RECT 84.830 283.450 85.680 284.300 ;
        RECT 103.780 283.450 104.630 284.300 ;
        RECT 4.830 282.500 5.680 283.350 ;
        RECT 23.780 282.500 24.630 283.350 ;
        RECT 24.830 282.500 25.680 283.350 ;
        RECT 43.780 282.500 44.630 283.350 ;
        RECT 44.830 282.500 45.680 283.350 ;
        RECT 63.780 282.500 64.630 283.350 ;
        RECT 64.830 282.500 65.680 283.350 ;
        RECT 83.780 282.500 84.630 283.350 ;
        RECT 84.830 282.500 85.680 283.350 ;
        RECT 103.780 282.500 104.630 283.350 ;
        RECT 4.830 281.050 5.680 281.900 ;
        RECT 4.830 280.100 5.680 280.950 ;
        RECT 5.780 280.100 6.630 280.950 ;
        RECT 7.230 280.100 8.080 280.950 ;
        RECT 8.180 280.100 9.030 280.950 ;
        RECT 23.780 281.050 24.630 281.900 ;
        RECT 24.830 281.050 25.680 281.900 ;
        RECT 4.830 279.050 5.680 279.900 ;
        RECT 5.780 279.050 6.630 279.900 ;
        RECT 7.230 279.050 8.080 279.900 ;
        RECT 8.180 279.050 9.030 279.900 ;
        RECT 11.630 280.100 12.280 280.750 ;
        RECT 12.430 280.100 13.080 280.750 ;
        RECT 13.230 280.100 13.880 280.750 ;
        RECT 15.580 280.100 16.230 280.750 ;
        RECT 16.380 280.100 17.030 280.750 ;
        RECT 17.180 280.100 17.830 280.750 ;
        RECT 11.630 279.250 12.280 279.900 ;
        RECT 12.430 279.250 13.080 279.900 ;
        RECT 13.230 279.250 13.880 279.900 ;
        RECT 15.580 279.250 16.230 279.900 ;
        RECT 16.380 279.250 17.030 279.900 ;
        RECT 17.180 279.250 17.830 279.900 ;
        RECT 20.430 280.100 21.280 280.950 ;
        RECT 21.380 280.100 22.230 280.950 ;
        RECT 22.830 280.100 23.680 280.950 ;
        RECT 23.780 280.100 24.630 280.950 ;
        RECT 24.830 280.100 25.680 280.950 ;
        RECT 25.780 280.100 26.630 280.950 ;
        RECT 27.230 280.100 28.080 280.950 ;
        RECT 28.180 280.100 29.030 280.950 ;
        RECT 43.780 281.050 44.630 281.900 ;
        RECT 44.830 281.050 45.680 281.900 ;
        RECT 4.830 278.100 5.680 278.950 ;
        RECT 20.430 279.050 21.280 279.900 ;
        RECT 21.380 279.050 22.230 279.900 ;
        RECT 22.830 279.050 23.680 279.900 ;
        RECT 23.780 279.050 24.630 279.900 ;
        RECT 24.830 279.050 25.680 279.900 ;
        RECT 25.780 279.050 26.630 279.900 ;
        RECT 27.230 279.050 28.080 279.900 ;
        RECT 28.180 279.050 29.030 279.900 ;
        RECT 31.630 280.100 32.280 280.750 ;
        RECT 32.430 280.100 33.080 280.750 ;
        RECT 33.230 280.100 33.880 280.750 ;
        RECT 35.580 280.100 36.230 280.750 ;
        RECT 36.380 280.100 37.030 280.750 ;
        RECT 37.180 280.100 37.830 280.750 ;
        RECT 31.630 279.250 32.280 279.900 ;
        RECT 32.430 279.250 33.080 279.900 ;
        RECT 33.230 279.250 33.880 279.900 ;
        RECT 35.580 279.250 36.230 279.900 ;
        RECT 36.380 279.250 37.030 279.900 ;
        RECT 37.180 279.250 37.830 279.900 ;
        RECT 40.430 280.100 41.280 280.950 ;
        RECT 41.380 280.100 42.230 280.950 ;
        RECT 42.830 280.100 43.680 280.950 ;
        RECT 43.780 280.100 44.630 280.950 ;
        RECT 44.830 280.100 45.680 280.950 ;
        RECT 45.780 280.100 46.630 280.950 ;
        RECT 47.230 280.100 48.080 280.950 ;
        RECT 48.180 280.100 49.030 280.950 ;
        RECT 63.780 281.050 64.630 281.900 ;
        RECT 64.830 281.050 65.680 281.900 ;
        RECT 23.780 278.100 24.630 278.950 ;
        RECT 24.830 278.100 25.680 278.950 ;
        RECT 40.430 279.050 41.280 279.900 ;
        RECT 41.380 279.050 42.230 279.900 ;
        RECT 42.830 279.050 43.680 279.900 ;
        RECT 43.780 279.050 44.630 279.900 ;
        RECT 44.830 279.050 45.680 279.900 ;
        RECT 45.780 279.050 46.630 279.900 ;
        RECT 47.230 279.050 48.080 279.900 ;
        RECT 48.180 279.050 49.030 279.900 ;
        RECT 51.630 280.100 52.280 280.750 ;
        RECT 52.430 280.100 53.080 280.750 ;
        RECT 53.230 280.100 53.880 280.750 ;
        RECT 55.580 280.100 56.230 280.750 ;
        RECT 56.380 280.100 57.030 280.750 ;
        RECT 57.180 280.100 57.830 280.750 ;
        RECT 51.630 279.250 52.280 279.900 ;
        RECT 52.430 279.250 53.080 279.900 ;
        RECT 53.230 279.250 53.880 279.900 ;
        RECT 55.580 279.250 56.230 279.900 ;
        RECT 56.380 279.250 57.030 279.900 ;
        RECT 57.180 279.250 57.830 279.900 ;
        RECT 60.430 280.100 61.280 280.950 ;
        RECT 61.380 280.100 62.230 280.950 ;
        RECT 62.830 280.100 63.680 280.950 ;
        RECT 63.780 280.100 64.630 280.950 ;
        RECT 64.830 280.100 65.680 280.950 ;
        RECT 65.780 280.100 66.630 280.950 ;
        RECT 67.230 280.100 68.080 280.950 ;
        RECT 68.180 280.100 69.030 280.950 ;
        RECT 83.780 281.050 84.630 281.900 ;
        RECT 84.830 281.050 85.680 281.900 ;
        RECT 43.780 278.100 44.630 278.950 ;
        RECT 44.830 278.100 45.680 278.950 ;
        RECT 60.430 279.050 61.280 279.900 ;
        RECT 61.380 279.050 62.230 279.900 ;
        RECT 62.830 279.050 63.680 279.900 ;
        RECT 63.780 279.050 64.630 279.900 ;
        RECT 64.830 279.050 65.680 279.900 ;
        RECT 65.780 279.050 66.630 279.900 ;
        RECT 67.230 279.050 68.080 279.900 ;
        RECT 68.180 279.050 69.030 279.900 ;
        RECT 71.630 280.100 72.280 280.750 ;
        RECT 72.430 280.100 73.080 280.750 ;
        RECT 73.230 280.100 73.880 280.750 ;
        RECT 75.580 280.100 76.230 280.750 ;
        RECT 76.380 280.100 77.030 280.750 ;
        RECT 77.180 280.100 77.830 280.750 ;
        RECT 71.630 279.250 72.280 279.900 ;
        RECT 72.430 279.250 73.080 279.900 ;
        RECT 73.230 279.250 73.880 279.900 ;
        RECT 75.580 279.250 76.230 279.900 ;
        RECT 76.380 279.250 77.030 279.900 ;
        RECT 77.180 279.250 77.830 279.900 ;
        RECT 80.430 280.100 81.280 280.950 ;
        RECT 81.380 280.100 82.230 280.950 ;
        RECT 82.830 280.100 83.680 280.950 ;
        RECT 83.780 280.100 84.630 280.950 ;
        RECT 84.830 280.100 85.680 280.950 ;
        RECT 85.780 280.100 86.630 280.950 ;
        RECT 87.230 280.100 88.080 280.950 ;
        RECT 88.180 280.100 89.030 280.950 ;
        RECT 103.780 281.050 104.630 281.900 ;
        RECT 63.780 278.100 64.630 278.950 ;
        RECT 64.830 278.100 65.680 278.950 ;
        RECT 80.430 279.050 81.280 279.900 ;
        RECT 81.380 279.050 82.230 279.900 ;
        RECT 82.830 279.050 83.680 279.900 ;
        RECT 83.780 279.050 84.630 279.900 ;
        RECT 84.830 279.050 85.680 279.900 ;
        RECT 85.780 279.050 86.630 279.900 ;
        RECT 87.230 279.050 88.080 279.900 ;
        RECT 88.180 279.050 89.030 279.900 ;
        RECT 91.630 280.100 92.280 280.750 ;
        RECT 92.430 280.100 93.080 280.750 ;
        RECT 93.230 280.100 93.880 280.750 ;
        RECT 95.580 280.100 96.230 280.750 ;
        RECT 96.380 280.100 97.030 280.750 ;
        RECT 97.180 280.100 97.830 280.750 ;
        RECT 91.630 279.250 92.280 279.900 ;
        RECT 92.430 279.250 93.080 279.900 ;
        RECT 93.230 279.250 93.880 279.900 ;
        RECT 95.580 279.250 96.230 279.900 ;
        RECT 96.380 279.250 97.030 279.900 ;
        RECT 97.180 279.250 97.830 279.900 ;
        RECT 100.430 280.100 101.280 280.950 ;
        RECT 101.380 280.100 102.230 280.950 ;
        RECT 102.830 280.100 103.680 280.950 ;
        RECT 103.780 280.100 104.630 280.950 ;
        RECT 83.780 278.100 84.630 278.950 ;
        RECT 84.830 278.100 85.680 278.950 ;
        RECT 100.430 279.050 101.280 279.900 ;
        RECT 101.380 279.050 102.230 279.900 ;
        RECT 102.830 279.050 103.680 279.900 ;
        RECT 103.780 279.050 104.630 279.900 ;
        RECT 103.780 278.100 104.630 278.950 ;
        RECT 4.830 276.650 5.680 277.500 ;
        RECT 23.780 276.650 24.630 277.500 ;
        RECT 24.830 276.650 25.680 277.500 ;
        RECT 43.780 276.650 44.630 277.500 ;
        RECT 44.830 276.650 45.680 277.500 ;
        RECT 63.780 276.650 64.630 277.500 ;
        RECT 64.830 276.650 65.680 277.500 ;
        RECT 83.780 276.650 84.630 277.500 ;
        RECT 84.830 276.650 85.680 277.500 ;
        RECT 103.780 276.650 104.630 277.500 ;
        RECT 4.830 275.700 5.680 276.550 ;
        RECT 23.780 275.700 24.630 276.550 ;
        RECT 24.830 275.700 25.680 276.550 ;
        RECT 43.780 275.700 44.630 276.550 ;
        RECT 44.830 275.700 45.680 276.550 ;
        RECT 63.780 275.700 64.630 276.550 ;
        RECT 64.830 275.700 65.680 276.550 ;
        RECT 83.780 275.700 84.630 276.550 ;
        RECT 84.830 275.700 85.680 276.550 ;
        RECT 103.780 275.700 104.630 276.550 ;
        RECT 4.830 272.450 5.480 273.100 ;
        RECT 4.830 271.650 5.480 272.300 ;
        RECT 4.830 270.850 5.480 271.500 ;
        RECT 4.830 268.500 5.480 269.150 ;
        RECT 4.830 267.700 5.480 268.350 ;
        RECT 4.830 266.900 5.480 267.550 ;
        RECT 23.980 272.450 24.630 273.100 ;
        RECT 24.830 272.450 25.480 273.100 ;
        RECT 23.980 271.650 24.630 272.300 ;
        RECT 24.830 271.650 25.480 272.300 ;
        RECT 23.980 270.850 24.630 271.500 ;
        RECT 24.830 270.850 25.480 271.500 ;
        RECT 23.980 268.500 24.630 269.150 ;
        RECT 24.830 268.500 25.480 269.150 ;
        RECT 23.980 267.700 24.630 268.350 ;
        RECT 24.830 267.700 25.480 268.350 ;
        RECT 23.980 266.900 24.630 267.550 ;
        RECT 24.830 266.900 25.480 267.550 ;
        RECT 43.980 272.450 44.630 273.100 ;
        RECT 44.830 272.450 45.480 273.100 ;
        RECT 43.980 271.650 44.630 272.300 ;
        RECT 44.830 271.650 45.480 272.300 ;
        RECT 43.980 270.850 44.630 271.500 ;
        RECT 44.830 270.850 45.480 271.500 ;
        RECT 43.980 268.500 44.630 269.150 ;
        RECT 44.830 268.500 45.480 269.150 ;
        RECT 43.980 267.700 44.630 268.350 ;
        RECT 44.830 267.700 45.480 268.350 ;
        RECT 43.980 266.900 44.630 267.550 ;
        RECT 44.830 266.900 45.480 267.550 ;
        RECT 63.980 272.450 64.630 273.100 ;
        RECT 64.830 272.450 65.480 273.100 ;
        RECT 63.980 271.650 64.630 272.300 ;
        RECT 64.830 271.650 65.480 272.300 ;
        RECT 63.980 270.850 64.630 271.500 ;
        RECT 64.830 270.850 65.480 271.500 ;
        RECT 63.980 268.500 64.630 269.150 ;
        RECT 64.830 268.500 65.480 269.150 ;
        RECT 63.980 267.700 64.630 268.350 ;
        RECT 64.830 267.700 65.480 268.350 ;
        RECT 63.980 266.900 64.630 267.550 ;
        RECT 64.830 266.900 65.480 267.550 ;
        RECT 83.980 272.450 84.630 273.100 ;
        RECT 84.830 272.450 85.480 273.100 ;
        RECT 83.980 271.650 84.630 272.300 ;
        RECT 84.830 271.650 85.480 272.300 ;
        RECT 83.980 270.850 84.630 271.500 ;
        RECT 84.830 270.850 85.480 271.500 ;
        RECT 83.980 268.500 84.630 269.150 ;
        RECT 84.830 268.500 85.480 269.150 ;
        RECT 83.980 267.700 84.630 268.350 ;
        RECT 84.830 267.700 85.480 268.350 ;
        RECT 83.980 266.900 84.630 267.550 ;
        RECT 84.830 266.900 85.480 267.550 ;
        RECT 103.980 272.450 104.630 273.100 ;
        RECT 103.980 271.650 104.630 272.300 ;
        RECT 103.980 270.850 104.630 271.500 ;
        RECT 103.980 268.500 104.630 269.150 ;
        RECT 103.980 267.700 104.630 268.350 ;
        RECT 103.980 266.900 104.630 267.550 ;
        RECT 4.830 263.450 5.680 264.300 ;
        RECT 23.780 263.450 24.630 264.300 ;
        RECT 24.830 263.450 25.680 264.300 ;
        RECT 43.780 263.450 44.630 264.300 ;
        RECT 44.830 263.450 45.680 264.300 ;
        RECT 63.780 263.450 64.630 264.300 ;
        RECT 64.830 263.450 65.680 264.300 ;
        RECT 83.780 263.450 84.630 264.300 ;
        RECT 84.830 263.450 85.680 264.300 ;
        RECT 103.780 263.450 104.630 264.300 ;
        RECT 4.830 262.500 5.680 263.350 ;
        RECT 23.780 262.500 24.630 263.350 ;
        RECT 24.830 262.500 25.680 263.350 ;
        RECT 43.780 262.500 44.630 263.350 ;
        RECT 44.830 262.500 45.680 263.350 ;
        RECT 63.780 262.500 64.630 263.350 ;
        RECT 64.830 262.500 65.680 263.350 ;
        RECT 83.780 262.500 84.630 263.350 ;
        RECT 84.830 262.500 85.680 263.350 ;
        RECT 103.780 262.500 104.630 263.350 ;
        RECT 4.830 261.050 5.680 261.900 ;
        RECT 4.830 260.100 5.680 260.950 ;
        RECT 5.780 260.100 6.630 260.950 ;
        RECT 7.230 260.100 8.080 260.950 ;
        RECT 8.180 260.100 9.030 260.950 ;
        RECT 23.780 261.050 24.630 261.900 ;
        RECT 24.830 261.050 25.680 261.900 ;
        RECT 4.830 259.050 5.680 259.900 ;
        RECT 5.780 259.050 6.630 259.900 ;
        RECT 7.230 259.050 8.080 259.900 ;
        RECT 8.180 259.050 9.030 259.900 ;
        RECT 11.630 260.100 12.280 260.750 ;
        RECT 12.430 260.100 13.080 260.750 ;
        RECT 13.230 260.100 13.880 260.750 ;
        RECT 15.580 260.100 16.230 260.750 ;
        RECT 16.380 260.100 17.030 260.750 ;
        RECT 17.180 260.100 17.830 260.750 ;
        RECT 11.630 259.250 12.280 259.900 ;
        RECT 12.430 259.250 13.080 259.900 ;
        RECT 13.230 259.250 13.880 259.900 ;
        RECT 15.580 259.250 16.230 259.900 ;
        RECT 16.380 259.250 17.030 259.900 ;
        RECT 17.180 259.250 17.830 259.900 ;
        RECT 20.430 260.100 21.280 260.950 ;
        RECT 21.380 260.100 22.230 260.950 ;
        RECT 22.830 260.100 23.680 260.950 ;
        RECT 23.780 260.100 24.630 260.950 ;
        RECT 24.830 260.100 25.680 260.950 ;
        RECT 25.780 260.100 26.630 260.950 ;
        RECT 27.230 260.100 28.080 260.950 ;
        RECT 28.180 260.100 29.030 260.950 ;
        RECT 43.780 261.050 44.630 261.900 ;
        RECT 44.830 261.050 45.680 261.900 ;
        RECT 4.830 258.100 5.680 258.950 ;
        RECT 20.430 259.050 21.280 259.900 ;
        RECT 21.380 259.050 22.230 259.900 ;
        RECT 22.830 259.050 23.680 259.900 ;
        RECT 23.780 259.050 24.630 259.900 ;
        RECT 24.830 259.050 25.680 259.900 ;
        RECT 25.780 259.050 26.630 259.900 ;
        RECT 27.230 259.050 28.080 259.900 ;
        RECT 28.180 259.050 29.030 259.900 ;
        RECT 31.630 260.100 32.280 260.750 ;
        RECT 32.430 260.100 33.080 260.750 ;
        RECT 33.230 260.100 33.880 260.750 ;
        RECT 35.580 260.100 36.230 260.750 ;
        RECT 36.380 260.100 37.030 260.750 ;
        RECT 37.180 260.100 37.830 260.750 ;
        RECT 31.630 259.250 32.280 259.900 ;
        RECT 32.430 259.250 33.080 259.900 ;
        RECT 33.230 259.250 33.880 259.900 ;
        RECT 35.580 259.250 36.230 259.900 ;
        RECT 36.380 259.250 37.030 259.900 ;
        RECT 37.180 259.250 37.830 259.900 ;
        RECT 40.430 260.100 41.280 260.950 ;
        RECT 41.380 260.100 42.230 260.950 ;
        RECT 42.830 260.100 43.680 260.950 ;
        RECT 43.780 260.100 44.630 260.950 ;
        RECT 44.830 260.100 45.680 260.950 ;
        RECT 45.780 260.100 46.630 260.950 ;
        RECT 47.230 260.100 48.080 260.950 ;
        RECT 48.180 260.100 49.030 260.950 ;
        RECT 63.780 261.050 64.630 261.900 ;
        RECT 64.830 261.050 65.680 261.900 ;
        RECT 23.780 258.100 24.630 258.950 ;
        RECT 24.830 258.100 25.680 258.950 ;
        RECT 40.430 259.050 41.280 259.900 ;
        RECT 41.380 259.050 42.230 259.900 ;
        RECT 42.830 259.050 43.680 259.900 ;
        RECT 43.780 259.050 44.630 259.900 ;
        RECT 44.830 259.050 45.680 259.900 ;
        RECT 45.780 259.050 46.630 259.900 ;
        RECT 47.230 259.050 48.080 259.900 ;
        RECT 48.180 259.050 49.030 259.900 ;
        RECT 51.630 260.100 52.280 260.750 ;
        RECT 52.430 260.100 53.080 260.750 ;
        RECT 53.230 260.100 53.880 260.750 ;
        RECT 55.580 260.100 56.230 260.750 ;
        RECT 56.380 260.100 57.030 260.750 ;
        RECT 57.180 260.100 57.830 260.750 ;
        RECT 51.630 259.250 52.280 259.900 ;
        RECT 52.430 259.250 53.080 259.900 ;
        RECT 53.230 259.250 53.880 259.900 ;
        RECT 55.580 259.250 56.230 259.900 ;
        RECT 56.380 259.250 57.030 259.900 ;
        RECT 57.180 259.250 57.830 259.900 ;
        RECT 60.430 260.100 61.280 260.950 ;
        RECT 61.380 260.100 62.230 260.950 ;
        RECT 62.830 260.100 63.680 260.950 ;
        RECT 63.780 260.100 64.630 260.950 ;
        RECT 64.830 260.100 65.680 260.950 ;
        RECT 65.780 260.100 66.630 260.950 ;
        RECT 67.230 260.100 68.080 260.950 ;
        RECT 68.180 260.100 69.030 260.950 ;
        RECT 83.780 261.050 84.630 261.900 ;
        RECT 84.830 261.050 85.680 261.900 ;
        RECT 43.780 258.100 44.630 258.950 ;
        RECT 44.830 258.100 45.680 258.950 ;
        RECT 60.430 259.050 61.280 259.900 ;
        RECT 61.380 259.050 62.230 259.900 ;
        RECT 62.830 259.050 63.680 259.900 ;
        RECT 63.780 259.050 64.630 259.900 ;
        RECT 64.830 259.050 65.680 259.900 ;
        RECT 65.780 259.050 66.630 259.900 ;
        RECT 67.230 259.050 68.080 259.900 ;
        RECT 68.180 259.050 69.030 259.900 ;
        RECT 71.630 260.100 72.280 260.750 ;
        RECT 72.430 260.100 73.080 260.750 ;
        RECT 73.230 260.100 73.880 260.750 ;
        RECT 75.580 260.100 76.230 260.750 ;
        RECT 76.380 260.100 77.030 260.750 ;
        RECT 77.180 260.100 77.830 260.750 ;
        RECT 71.630 259.250 72.280 259.900 ;
        RECT 72.430 259.250 73.080 259.900 ;
        RECT 73.230 259.250 73.880 259.900 ;
        RECT 75.580 259.250 76.230 259.900 ;
        RECT 76.380 259.250 77.030 259.900 ;
        RECT 77.180 259.250 77.830 259.900 ;
        RECT 80.430 260.100 81.280 260.950 ;
        RECT 81.380 260.100 82.230 260.950 ;
        RECT 82.830 260.100 83.680 260.950 ;
        RECT 83.780 260.100 84.630 260.950 ;
        RECT 84.830 260.100 85.680 260.950 ;
        RECT 85.780 260.100 86.630 260.950 ;
        RECT 87.230 260.100 88.080 260.950 ;
        RECT 88.180 260.100 89.030 260.950 ;
        RECT 103.780 261.050 104.630 261.900 ;
        RECT 63.780 258.100 64.630 258.950 ;
        RECT 64.830 258.100 65.680 258.950 ;
        RECT 80.430 259.050 81.280 259.900 ;
        RECT 81.380 259.050 82.230 259.900 ;
        RECT 82.830 259.050 83.680 259.900 ;
        RECT 83.780 259.050 84.630 259.900 ;
        RECT 84.830 259.050 85.680 259.900 ;
        RECT 85.780 259.050 86.630 259.900 ;
        RECT 87.230 259.050 88.080 259.900 ;
        RECT 88.180 259.050 89.030 259.900 ;
        RECT 91.630 260.100 92.280 260.750 ;
        RECT 92.430 260.100 93.080 260.750 ;
        RECT 93.230 260.100 93.880 260.750 ;
        RECT 95.580 260.100 96.230 260.750 ;
        RECT 96.380 260.100 97.030 260.750 ;
        RECT 97.180 260.100 97.830 260.750 ;
        RECT 91.630 259.250 92.280 259.900 ;
        RECT 92.430 259.250 93.080 259.900 ;
        RECT 93.230 259.250 93.880 259.900 ;
        RECT 95.580 259.250 96.230 259.900 ;
        RECT 96.380 259.250 97.030 259.900 ;
        RECT 97.180 259.250 97.830 259.900 ;
        RECT 100.430 260.100 101.280 260.950 ;
        RECT 101.380 260.100 102.230 260.950 ;
        RECT 102.830 260.100 103.680 260.950 ;
        RECT 103.780 260.100 104.630 260.950 ;
        RECT 83.780 258.100 84.630 258.950 ;
        RECT 84.830 258.100 85.680 258.950 ;
        RECT 100.430 259.050 101.280 259.900 ;
        RECT 101.380 259.050 102.230 259.900 ;
        RECT 102.830 259.050 103.680 259.900 ;
        RECT 103.780 259.050 104.630 259.900 ;
        RECT 103.780 258.100 104.630 258.950 ;
        RECT 4.830 256.650 5.680 257.500 ;
        RECT 23.780 256.650 24.630 257.500 ;
        RECT 24.830 256.650 25.680 257.500 ;
        RECT 43.780 256.650 44.630 257.500 ;
        RECT 44.830 256.650 45.680 257.500 ;
        RECT 63.780 256.650 64.630 257.500 ;
        RECT 64.830 256.650 65.680 257.500 ;
        RECT 83.780 256.650 84.630 257.500 ;
        RECT 84.830 256.650 85.680 257.500 ;
        RECT 103.780 256.650 104.630 257.500 ;
        RECT 4.830 255.700 5.680 256.550 ;
        RECT 23.780 255.700 24.630 256.550 ;
        RECT 24.830 255.700 25.680 256.550 ;
        RECT 43.780 255.700 44.630 256.550 ;
        RECT 44.830 255.700 45.680 256.550 ;
        RECT 63.780 255.700 64.630 256.550 ;
        RECT 64.830 255.700 65.680 256.550 ;
        RECT 83.780 255.700 84.630 256.550 ;
        RECT 84.830 255.700 85.680 256.550 ;
        RECT 103.780 255.700 104.630 256.550 ;
        RECT 4.830 252.450 5.480 253.100 ;
        RECT 4.830 251.650 5.480 252.300 ;
        RECT 4.830 250.850 5.480 251.500 ;
        RECT 4.830 248.500 5.480 249.150 ;
        RECT 4.830 247.700 5.480 248.350 ;
        RECT 4.830 246.900 5.480 247.550 ;
        RECT 23.980 252.450 24.630 253.100 ;
        RECT 24.830 252.450 25.480 253.100 ;
        RECT 23.980 251.650 24.630 252.300 ;
        RECT 24.830 251.650 25.480 252.300 ;
        RECT 23.980 250.850 24.630 251.500 ;
        RECT 24.830 250.850 25.480 251.500 ;
        RECT 23.980 248.500 24.630 249.150 ;
        RECT 24.830 248.500 25.480 249.150 ;
        RECT 23.980 247.700 24.630 248.350 ;
        RECT 24.830 247.700 25.480 248.350 ;
        RECT 23.980 246.900 24.630 247.550 ;
        RECT 24.830 246.900 25.480 247.550 ;
        RECT 43.980 252.450 44.630 253.100 ;
        RECT 44.830 252.450 45.480 253.100 ;
        RECT 43.980 251.650 44.630 252.300 ;
        RECT 44.830 251.650 45.480 252.300 ;
        RECT 43.980 250.850 44.630 251.500 ;
        RECT 44.830 250.850 45.480 251.500 ;
        RECT 43.980 248.500 44.630 249.150 ;
        RECT 44.830 248.500 45.480 249.150 ;
        RECT 43.980 247.700 44.630 248.350 ;
        RECT 44.830 247.700 45.480 248.350 ;
        RECT 43.980 246.900 44.630 247.550 ;
        RECT 44.830 246.900 45.480 247.550 ;
        RECT 63.980 252.450 64.630 253.100 ;
        RECT 64.830 252.450 65.480 253.100 ;
        RECT 63.980 251.650 64.630 252.300 ;
        RECT 64.830 251.650 65.480 252.300 ;
        RECT 63.980 250.850 64.630 251.500 ;
        RECT 64.830 250.850 65.480 251.500 ;
        RECT 63.980 248.500 64.630 249.150 ;
        RECT 64.830 248.500 65.480 249.150 ;
        RECT 63.980 247.700 64.630 248.350 ;
        RECT 64.830 247.700 65.480 248.350 ;
        RECT 63.980 246.900 64.630 247.550 ;
        RECT 64.830 246.900 65.480 247.550 ;
        RECT 83.980 252.450 84.630 253.100 ;
        RECT 84.830 252.450 85.480 253.100 ;
        RECT 83.980 251.650 84.630 252.300 ;
        RECT 84.830 251.650 85.480 252.300 ;
        RECT 83.980 250.850 84.630 251.500 ;
        RECT 84.830 250.850 85.480 251.500 ;
        RECT 83.980 248.500 84.630 249.150 ;
        RECT 84.830 248.500 85.480 249.150 ;
        RECT 83.980 247.700 84.630 248.350 ;
        RECT 84.830 247.700 85.480 248.350 ;
        RECT 83.980 246.900 84.630 247.550 ;
        RECT 84.830 246.900 85.480 247.550 ;
        RECT 103.980 252.450 104.630 253.100 ;
        RECT 103.980 251.650 104.630 252.300 ;
        RECT 103.980 250.850 104.630 251.500 ;
        RECT 103.980 248.500 104.630 249.150 ;
        RECT 103.980 247.700 104.630 248.350 ;
        RECT 103.980 246.900 104.630 247.550 ;
        RECT 4.830 243.450 5.680 244.300 ;
        RECT 23.780 243.450 24.630 244.300 ;
        RECT 24.830 243.450 25.680 244.300 ;
        RECT 43.780 243.450 44.630 244.300 ;
        RECT 44.830 243.450 45.680 244.300 ;
        RECT 63.780 243.450 64.630 244.300 ;
        RECT 64.830 243.450 65.680 244.300 ;
        RECT 83.780 243.450 84.630 244.300 ;
        RECT 84.830 243.450 85.680 244.300 ;
        RECT 103.780 243.450 104.630 244.300 ;
        RECT 4.830 242.500 5.680 243.350 ;
        RECT 23.780 242.500 24.630 243.350 ;
        RECT 24.830 242.500 25.680 243.350 ;
        RECT 43.780 242.500 44.630 243.350 ;
        RECT 44.830 242.500 45.680 243.350 ;
        RECT 63.780 242.500 64.630 243.350 ;
        RECT 64.830 242.500 65.680 243.350 ;
        RECT 83.780 242.500 84.630 243.350 ;
        RECT 84.830 242.500 85.680 243.350 ;
        RECT 103.780 242.500 104.630 243.350 ;
        RECT 4.830 241.050 5.680 241.900 ;
        RECT 4.830 240.100 5.680 240.950 ;
        RECT 5.780 240.100 6.630 240.950 ;
        RECT 7.230 240.100 8.080 240.950 ;
        RECT 8.180 240.100 9.030 240.950 ;
        RECT 23.780 241.050 24.630 241.900 ;
        RECT 24.830 241.050 25.680 241.900 ;
        RECT 4.830 239.050 5.680 239.900 ;
        RECT 5.780 239.050 6.630 239.900 ;
        RECT 7.230 239.050 8.080 239.900 ;
        RECT 8.180 239.050 9.030 239.900 ;
        RECT 11.630 240.100 12.280 240.750 ;
        RECT 12.430 240.100 13.080 240.750 ;
        RECT 13.230 240.100 13.880 240.750 ;
        RECT 15.580 240.100 16.230 240.750 ;
        RECT 16.380 240.100 17.030 240.750 ;
        RECT 17.180 240.100 17.830 240.750 ;
        RECT 11.630 239.250 12.280 239.900 ;
        RECT 12.430 239.250 13.080 239.900 ;
        RECT 13.230 239.250 13.880 239.900 ;
        RECT 15.580 239.250 16.230 239.900 ;
        RECT 16.380 239.250 17.030 239.900 ;
        RECT 17.180 239.250 17.830 239.900 ;
        RECT 20.430 240.100 21.280 240.950 ;
        RECT 21.380 240.100 22.230 240.950 ;
        RECT 22.830 240.100 23.680 240.950 ;
        RECT 23.780 240.100 24.630 240.950 ;
        RECT 24.830 240.100 25.680 240.950 ;
        RECT 25.780 240.100 26.630 240.950 ;
        RECT 27.230 240.100 28.080 240.950 ;
        RECT 28.180 240.100 29.030 240.950 ;
        RECT 43.780 241.050 44.630 241.900 ;
        RECT 44.830 241.050 45.680 241.900 ;
        RECT 4.830 238.100 5.680 238.950 ;
        RECT 20.430 239.050 21.280 239.900 ;
        RECT 21.380 239.050 22.230 239.900 ;
        RECT 22.830 239.050 23.680 239.900 ;
        RECT 23.780 239.050 24.630 239.900 ;
        RECT 24.830 239.050 25.680 239.900 ;
        RECT 25.780 239.050 26.630 239.900 ;
        RECT 27.230 239.050 28.080 239.900 ;
        RECT 28.180 239.050 29.030 239.900 ;
        RECT 31.630 240.100 32.280 240.750 ;
        RECT 32.430 240.100 33.080 240.750 ;
        RECT 33.230 240.100 33.880 240.750 ;
        RECT 35.580 240.100 36.230 240.750 ;
        RECT 36.380 240.100 37.030 240.750 ;
        RECT 37.180 240.100 37.830 240.750 ;
        RECT 31.630 239.250 32.280 239.900 ;
        RECT 32.430 239.250 33.080 239.900 ;
        RECT 33.230 239.250 33.880 239.900 ;
        RECT 35.580 239.250 36.230 239.900 ;
        RECT 36.380 239.250 37.030 239.900 ;
        RECT 37.180 239.250 37.830 239.900 ;
        RECT 40.430 240.100 41.280 240.950 ;
        RECT 41.380 240.100 42.230 240.950 ;
        RECT 42.830 240.100 43.680 240.950 ;
        RECT 43.780 240.100 44.630 240.950 ;
        RECT 44.830 240.100 45.680 240.950 ;
        RECT 45.780 240.100 46.630 240.950 ;
        RECT 47.230 240.100 48.080 240.950 ;
        RECT 48.180 240.100 49.030 240.950 ;
        RECT 63.780 241.050 64.630 241.900 ;
        RECT 64.830 241.050 65.680 241.900 ;
        RECT 23.780 238.100 24.630 238.950 ;
        RECT 24.830 238.100 25.680 238.950 ;
        RECT 40.430 239.050 41.280 239.900 ;
        RECT 41.380 239.050 42.230 239.900 ;
        RECT 42.830 239.050 43.680 239.900 ;
        RECT 43.780 239.050 44.630 239.900 ;
        RECT 44.830 239.050 45.680 239.900 ;
        RECT 45.780 239.050 46.630 239.900 ;
        RECT 47.230 239.050 48.080 239.900 ;
        RECT 48.180 239.050 49.030 239.900 ;
        RECT 51.630 240.100 52.280 240.750 ;
        RECT 52.430 240.100 53.080 240.750 ;
        RECT 53.230 240.100 53.880 240.750 ;
        RECT 55.580 240.100 56.230 240.750 ;
        RECT 56.380 240.100 57.030 240.750 ;
        RECT 57.180 240.100 57.830 240.750 ;
        RECT 51.630 239.250 52.280 239.900 ;
        RECT 52.430 239.250 53.080 239.900 ;
        RECT 53.230 239.250 53.880 239.900 ;
        RECT 55.580 239.250 56.230 239.900 ;
        RECT 56.380 239.250 57.030 239.900 ;
        RECT 57.180 239.250 57.830 239.900 ;
        RECT 60.430 240.100 61.280 240.950 ;
        RECT 61.380 240.100 62.230 240.950 ;
        RECT 62.830 240.100 63.680 240.950 ;
        RECT 63.780 240.100 64.630 240.950 ;
        RECT 64.830 240.100 65.680 240.950 ;
        RECT 65.780 240.100 66.630 240.950 ;
        RECT 67.230 240.100 68.080 240.950 ;
        RECT 68.180 240.100 69.030 240.950 ;
        RECT 83.780 241.050 84.630 241.900 ;
        RECT 84.830 241.050 85.680 241.900 ;
        RECT 43.780 238.100 44.630 238.950 ;
        RECT 44.830 238.100 45.680 238.950 ;
        RECT 60.430 239.050 61.280 239.900 ;
        RECT 61.380 239.050 62.230 239.900 ;
        RECT 62.830 239.050 63.680 239.900 ;
        RECT 63.780 239.050 64.630 239.900 ;
        RECT 64.830 239.050 65.680 239.900 ;
        RECT 65.780 239.050 66.630 239.900 ;
        RECT 67.230 239.050 68.080 239.900 ;
        RECT 68.180 239.050 69.030 239.900 ;
        RECT 71.630 240.100 72.280 240.750 ;
        RECT 72.430 240.100 73.080 240.750 ;
        RECT 73.230 240.100 73.880 240.750 ;
        RECT 75.580 240.100 76.230 240.750 ;
        RECT 76.380 240.100 77.030 240.750 ;
        RECT 77.180 240.100 77.830 240.750 ;
        RECT 71.630 239.250 72.280 239.900 ;
        RECT 72.430 239.250 73.080 239.900 ;
        RECT 73.230 239.250 73.880 239.900 ;
        RECT 75.580 239.250 76.230 239.900 ;
        RECT 76.380 239.250 77.030 239.900 ;
        RECT 77.180 239.250 77.830 239.900 ;
        RECT 80.430 240.100 81.280 240.950 ;
        RECT 81.380 240.100 82.230 240.950 ;
        RECT 82.830 240.100 83.680 240.950 ;
        RECT 83.780 240.100 84.630 240.950 ;
        RECT 84.830 240.100 85.680 240.950 ;
        RECT 85.780 240.100 86.630 240.950 ;
        RECT 87.230 240.100 88.080 240.950 ;
        RECT 88.180 240.100 89.030 240.950 ;
        RECT 103.780 241.050 104.630 241.900 ;
        RECT 63.780 238.100 64.630 238.950 ;
        RECT 64.830 238.100 65.680 238.950 ;
        RECT 80.430 239.050 81.280 239.900 ;
        RECT 81.380 239.050 82.230 239.900 ;
        RECT 82.830 239.050 83.680 239.900 ;
        RECT 83.780 239.050 84.630 239.900 ;
        RECT 84.830 239.050 85.680 239.900 ;
        RECT 85.780 239.050 86.630 239.900 ;
        RECT 87.230 239.050 88.080 239.900 ;
        RECT 88.180 239.050 89.030 239.900 ;
        RECT 91.630 240.100 92.280 240.750 ;
        RECT 92.430 240.100 93.080 240.750 ;
        RECT 93.230 240.100 93.880 240.750 ;
        RECT 95.580 240.100 96.230 240.750 ;
        RECT 96.380 240.100 97.030 240.750 ;
        RECT 97.180 240.100 97.830 240.750 ;
        RECT 91.630 239.250 92.280 239.900 ;
        RECT 92.430 239.250 93.080 239.900 ;
        RECT 93.230 239.250 93.880 239.900 ;
        RECT 95.580 239.250 96.230 239.900 ;
        RECT 96.380 239.250 97.030 239.900 ;
        RECT 97.180 239.250 97.830 239.900 ;
        RECT 100.430 240.100 101.280 240.950 ;
        RECT 101.380 240.100 102.230 240.950 ;
        RECT 102.830 240.100 103.680 240.950 ;
        RECT 103.780 240.100 104.630 240.950 ;
        RECT 83.780 238.100 84.630 238.950 ;
        RECT 84.830 238.100 85.680 238.950 ;
        RECT 100.430 239.050 101.280 239.900 ;
        RECT 101.380 239.050 102.230 239.900 ;
        RECT 102.830 239.050 103.680 239.900 ;
        RECT 103.780 239.050 104.630 239.900 ;
        RECT 103.780 238.100 104.630 238.950 ;
        RECT 4.830 236.650 5.680 237.500 ;
        RECT 23.780 236.650 24.630 237.500 ;
        RECT 24.830 236.650 25.680 237.500 ;
        RECT 43.780 236.650 44.630 237.500 ;
        RECT 44.830 236.650 45.680 237.500 ;
        RECT 63.780 236.650 64.630 237.500 ;
        RECT 64.830 236.650 65.680 237.500 ;
        RECT 83.780 236.650 84.630 237.500 ;
        RECT 84.830 236.650 85.680 237.500 ;
        RECT 103.780 236.650 104.630 237.500 ;
        RECT 4.830 235.700 5.680 236.550 ;
        RECT 23.780 235.700 24.630 236.550 ;
        RECT 24.830 235.700 25.680 236.550 ;
        RECT 43.780 235.700 44.630 236.550 ;
        RECT 44.830 235.700 45.680 236.550 ;
        RECT 63.780 235.700 64.630 236.550 ;
        RECT 64.830 235.700 65.680 236.550 ;
        RECT 83.780 235.700 84.630 236.550 ;
        RECT 84.830 235.700 85.680 236.550 ;
        RECT 103.780 235.700 104.630 236.550 ;
        RECT 4.830 232.450 5.480 233.100 ;
        RECT 4.830 231.650 5.480 232.300 ;
        RECT 4.830 230.850 5.480 231.500 ;
        RECT 4.830 228.500 5.480 229.150 ;
        RECT 4.830 227.700 5.480 228.350 ;
        RECT 4.830 226.900 5.480 227.550 ;
        RECT 23.980 232.450 24.630 233.100 ;
        RECT 24.830 232.450 25.480 233.100 ;
        RECT 23.980 231.650 24.630 232.300 ;
        RECT 24.830 231.650 25.480 232.300 ;
        RECT 23.980 230.850 24.630 231.500 ;
        RECT 24.830 230.850 25.480 231.500 ;
        RECT 23.980 228.500 24.630 229.150 ;
        RECT 24.830 228.500 25.480 229.150 ;
        RECT 23.980 227.700 24.630 228.350 ;
        RECT 24.830 227.700 25.480 228.350 ;
        RECT 23.980 226.900 24.630 227.550 ;
        RECT 24.830 226.900 25.480 227.550 ;
        RECT 43.980 232.450 44.630 233.100 ;
        RECT 44.830 232.450 45.480 233.100 ;
        RECT 43.980 231.650 44.630 232.300 ;
        RECT 44.830 231.650 45.480 232.300 ;
        RECT 43.980 230.850 44.630 231.500 ;
        RECT 44.830 230.850 45.480 231.500 ;
        RECT 43.980 228.500 44.630 229.150 ;
        RECT 44.830 228.500 45.480 229.150 ;
        RECT 43.980 227.700 44.630 228.350 ;
        RECT 44.830 227.700 45.480 228.350 ;
        RECT 43.980 226.900 44.630 227.550 ;
        RECT 44.830 226.900 45.480 227.550 ;
        RECT 63.980 232.450 64.630 233.100 ;
        RECT 64.830 232.450 65.480 233.100 ;
        RECT 63.980 231.650 64.630 232.300 ;
        RECT 64.830 231.650 65.480 232.300 ;
        RECT 63.980 230.850 64.630 231.500 ;
        RECT 64.830 230.850 65.480 231.500 ;
        RECT 63.980 228.500 64.630 229.150 ;
        RECT 64.830 228.500 65.480 229.150 ;
        RECT 63.980 227.700 64.630 228.350 ;
        RECT 64.830 227.700 65.480 228.350 ;
        RECT 63.980 226.900 64.630 227.550 ;
        RECT 64.830 226.900 65.480 227.550 ;
        RECT 83.980 232.450 84.630 233.100 ;
        RECT 84.830 232.450 85.480 233.100 ;
        RECT 83.980 231.650 84.630 232.300 ;
        RECT 84.830 231.650 85.480 232.300 ;
        RECT 83.980 230.850 84.630 231.500 ;
        RECT 84.830 230.850 85.480 231.500 ;
        RECT 83.980 228.500 84.630 229.150 ;
        RECT 84.830 228.500 85.480 229.150 ;
        RECT 83.980 227.700 84.630 228.350 ;
        RECT 84.830 227.700 85.480 228.350 ;
        RECT 83.980 226.900 84.630 227.550 ;
        RECT 84.830 226.900 85.480 227.550 ;
        RECT 103.980 232.450 104.630 233.100 ;
        RECT 103.980 231.650 104.630 232.300 ;
        RECT 103.980 230.850 104.630 231.500 ;
        RECT 103.980 228.500 104.630 229.150 ;
        RECT 103.980 227.700 104.630 228.350 ;
        RECT 103.980 226.900 104.630 227.550 ;
        RECT 4.830 223.450 5.680 224.300 ;
        RECT 23.780 223.450 24.630 224.300 ;
        RECT 24.830 223.450 25.680 224.300 ;
        RECT 43.780 223.450 44.630 224.300 ;
        RECT 44.830 223.450 45.680 224.300 ;
        RECT 63.780 223.450 64.630 224.300 ;
        RECT 64.830 223.450 65.680 224.300 ;
        RECT 83.780 223.450 84.630 224.300 ;
        RECT 84.830 223.450 85.680 224.300 ;
        RECT 103.780 223.450 104.630 224.300 ;
        RECT 4.830 222.500 5.680 223.350 ;
        RECT 23.780 222.500 24.630 223.350 ;
        RECT 24.830 222.500 25.680 223.350 ;
        RECT 43.780 222.500 44.630 223.350 ;
        RECT 44.830 222.500 45.680 223.350 ;
        RECT 63.780 222.500 64.630 223.350 ;
        RECT 64.830 222.500 65.680 223.350 ;
        RECT 83.780 222.500 84.630 223.350 ;
        RECT 84.830 222.500 85.680 223.350 ;
        RECT 103.780 222.500 104.630 223.350 ;
        RECT 4.830 221.050 5.680 221.900 ;
        RECT 4.830 220.100 5.680 220.950 ;
        RECT 5.780 220.100 6.630 220.950 ;
        RECT 7.230 220.100 8.080 220.950 ;
        RECT 8.180 220.100 9.030 220.950 ;
        RECT 23.780 221.050 24.630 221.900 ;
        RECT 24.830 221.050 25.680 221.900 ;
        RECT 11.630 220.100 12.280 220.750 ;
        RECT 12.430 220.100 13.080 220.750 ;
        RECT 13.230 220.100 13.880 220.750 ;
        RECT 15.580 220.100 16.230 220.750 ;
        RECT 16.380 220.100 17.030 220.750 ;
        RECT 17.180 220.100 17.830 220.750 ;
        RECT 20.430 220.100 21.280 220.950 ;
        RECT 21.380 220.100 22.230 220.950 ;
        RECT 22.830 220.100 23.680 220.950 ;
        RECT 23.780 220.100 24.630 220.950 ;
        RECT 24.830 220.100 25.680 220.950 ;
        RECT 25.780 220.100 26.630 220.950 ;
        RECT 27.230 220.100 28.080 220.950 ;
        RECT 28.180 220.100 29.030 220.950 ;
        RECT 43.780 221.050 44.630 221.900 ;
        RECT 44.830 221.050 45.680 221.900 ;
        RECT 31.630 220.100 32.280 220.750 ;
        RECT 32.430 220.100 33.080 220.750 ;
        RECT 33.230 220.100 33.880 220.750 ;
        RECT 35.580 220.100 36.230 220.750 ;
        RECT 36.380 220.100 37.030 220.750 ;
        RECT 37.180 220.100 37.830 220.750 ;
        RECT 40.430 220.100 41.280 220.950 ;
        RECT 41.380 220.100 42.230 220.950 ;
        RECT 42.830 220.100 43.680 220.950 ;
        RECT 43.780 220.100 44.630 220.950 ;
        RECT 44.830 220.100 45.680 220.950 ;
        RECT 45.780 220.100 46.630 220.950 ;
        RECT 47.230 220.100 48.080 220.950 ;
        RECT 48.180 220.100 49.030 220.950 ;
        RECT 63.780 221.050 64.630 221.900 ;
        RECT 64.830 221.050 65.680 221.900 ;
        RECT 51.630 220.100 52.280 220.750 ;
        RECT 52.430 220.100 53.080 220.750 ;
        RECT 53.230 220.100 53.880 220.750 ;
        RECT 55.580 220.100 56.230 220.750 ;
        RECT 56.380 220.100 57.030 220.750 ;
        RECT 57.180 220.100 57.830 220.750 ;
        RECT 60.430 220.100 61.280 220.950 ;
        RECT 61.380 220.100 62.230 220.950 ;
        RECT 62.830 220.100 63.680 220.950 ;
        RECT 63.780 220.100 64.630 220.950 ;
        RECT 64.830 220.100 65.680 220.950 ;
        RECT 65.780 220.100 66.630 220.950 ;
        RECT 67.230 220.100 68.080 220.950 ;
        RECT 68.180 220.100 69.030 220.950 ;
        RECT 83.780 221.050 84.630 221.900 ;
        RECT 84.830 221.050 85.680 221.900 ;
        RECT 71.630 220.100 72.280 220.750 ;
        RECT 72.430 220.100 73.080 220.750 ;
        RECT 73.230 220.100 73.880 220.750 ;
        RECT 75.580 220.100 76.230 220.750 ;
        RECT 76.380 220.100 77.030 220.750 ;
        RECT 77.180 220.100 77.830 220.750 ;
        RECT 80.430 220.100 81.280 220.950 ;
        RECT 81.380 220.100 82.230 220.950 ;
        RECT 82.830 220.100 83.680 220.950 ;
        RECT 83.780 220.100 84.630 220.950 ;
        RECT 84.830 220.100 85.680 220.950 ;
        RECT 85.780 220.100 86.630 220.950 ;
        RECT 87.230 220.100 88.080 220.950 ;
        RECT 88.180 220.100 89.030 220.950 ;
        RECT 103.780 221.050 104.630 221.900 ;
        RECT 91.630 220.100 92.280 220.750 ;
        RECT 92.430 220.100 93.080 220.750 ;
        RECT 93.230 220.100 93.880 220.750 ;
        RECT 95.580 220.100 96.230 220.750 ;
        RECT 96.380 220.100 97.030 220.750 ;
        RECT 97.180 220.100 97.830 220.750 ;
        RECT 100.430 220.100 101.280 220.950 ;
        RECT 101.380 220.100 102.230 220.950 ;
        RECT 102.830 220.100 103.680 220.950 ;
        RECT 103.780 220.100 104.630 220.950 ;
        RECT 11.245 199.305 11.565 199.625 ;
        RECT 11.685 199.305 12.005 199.625 ;
        RECT 11.245 198.905 11.565 199.225 ;
        RECT 11.685 198.905 12.005 199.225 ;
        RECT 20.960 199.205 21.280 199.525 ;
        RECT 21.400 199.205 21.720 199.525 ;
        RECT 20.960 198.805 21.280 199.125 ;
        RECT 21.400 198.805 21.720 199.125 ;
        RECT 12.680 181.995 13.000 182.315 ;
        RECT 13.120 181.995 13.440 182.315 ;
        RECT 11.630 159.250 12.280 159.900 ;
        RECT 12.430 159.250 13.080 159.900 ;
        RECT 13.230 159.250 13.880 159.900 ;
        RECT 15.580 159.250 16.230 159.900 ;
        RECT 16.380 159.250 17.030 159.900 ;
        RECT 17.180 159.250 17.830 159.900 ;
        RECT 31.630 159.250 32.280 159.900 ;
        RECT 32.430 159.250 33.080 159.900 ;
        RECT 33.230 159.250 33.880 159.900 ;
        RECT 35.580 159.250 36.230 159.900 ;
        RECT 36.380 159.250 37.030 159.900 ;
        RECT 37.180 159.250 37.830 159.900 ;
        RECT 51.630 159.250 52.280 159.900 ;
        RECT 52.430 159.250 53.080 159.900 ;
        RECT 53.230 159.250 53.880 159.900 ;
        RECT 55.580 159.250 56.230 159.900 ;
        RECT 56.380 159.250 57.030 159.900 ;
        RECT 57.180 159.250 57.830 159.900 ;
        RECT 71.630 159.250 72.280 159.900 ;
        RECT 72.430 159.250 73.080 159.900 ;
        RECT 73.230 159.250 73.880 159.900 ;
        RECT 75.580 159.250 76.230 159.900 ;
        RECT 76.380 159.250 77.030 159.900 ;
        RECT 77.180 159.250 77.830 159.900 ;
        RECT 91.630 159.250 92.280 159.900 ;
        RECT 92.430 159.250 93.080 159.900 ;
        RECT 93.230 159.250 93.880 159.900 ;
        RECT 95.580 159.250 96.230 159.900 ;
        RECT 96.380 159.250 97.030 159.900 ;
        RECT 97.180 159.250 97.830 159.900 ;
        RECT 4.830 152.450 5.480 153.100 ;
        RECT 4.830 151.650 5.480 152.300 ;
        RECT 4.830 150.850 5.480 151.500 ;
        RECT 4.830 148.500 5.480 149.150 ;
        RECT 4.830 147.700 5.480 148.350 ;
        RECT 4.830 146.900 5.480 147.550 ;
        RECT 23.980 152.450 24.630 153.100 ;
        RECT 24.830 152.450 25.480 153.100 ;
        RECT 23.980 151.650 24.630 152.300 ;
        RECT 24.830 151.650 25.480 152.300 ;
        RECT 23.980 150.850 24.630 151.500 ;
        RECT 24.830 150.850 25.480 151.500 ;
        RECT 23.980 148.500 24.630 149.150 ;
        RECT 24.830 148.500 25.480 149.150 ;
        RECT 23.980 147.700 24.630 148.350 ;
        RECT 24.830 147.700 25.480 148.350 ;
        RECT 23.980 146.900 24.630 147.550 ;
        RECT 24.830 146.900 25.480 147.550 ;
        RECT 43.980 152.450 44.630 153.100 ;
        RECT 44.830 152.450 45.480 153.100 ;
        RECT 43.980 151.650 44.630 152.300 ;
        RECT 44.830 151.650 45.480 152.300 ;
        RECT 43.980 150.850 44.630 151.500 ;
        RECT 44.830 150.850 45.480 151.500 ;
        RECT 43.980 148.500 44.630 149.150 ;
        RECT 44.830 148.500 45.480 149.150 ;
        RECT 43.980 147.700 44.630 148.350 ;
        RECT 44.830 147.700 45.480 148.350 ;
        RECT 43.980 146.900 44.630 147.550 ;
        RECT 44.830 146.900 45.480 147.550 ;
        RECT 63.980 152.450 64.630 153.100 ;
        RECT 64.830 152.450 65.480 153.100 ;
        RECT 63.980 151.650 64.630 152.300 ;
        RECT 64.830 151.650 65.480 152.300 ;
        RECT 63.980 150.850 64.630 151.500 ;
        RECT 64.830 150.850 65.480 151.500 ;
        RECT 63.980 148.500 64.630 149.150 ;
        RECT 64.830 148.500 65.480 149.150 ;
        RECT 63.980 147.700 64.630 148.350 ;
        RECT 64.830 147.700 65.480 148.350 ;
        RECT 63.980 146.900 64.630 147.550 ;
        RECT 64.830 146.900 65.480 147.550 ;
        RECT 83.980 152.450 84.630 153.100 ;
        RECT 84.830 152.450 85.480 153.100 ;
        RECT 83.980 151.650 84.630 152.300 ;
        RECT 84.830 151.650 85.480 152.300 ;
        RECT 83.980 150.850 84.630 151.500 ;
        RECT 84.830 150.850 85.480 151.500 ;
        RECT 83.980 148.500 84.630 149.150 ;
        RECT 84.830 148.500 85.480 149.150 ;
        RECT 83.980 147.700 84.630 148.350 ;
        RECT 84.830 147.700 85.480 148.350 ;
        RECT 83.980 146.900 84.630 147.550 ;
        RECT 84.830 146.900 85.480 147.550 ;
        RECT 103.980 152.450 104.630 153.100 ;
        RECT 103.980 151.650 104.630 152.300 ;
        RECT 103.980 150.850 104.630 151.500 ;
        RECT 103.980 148.500 104.630 149.150 ;
        RECT 103.980 147.700 104.630 148.350 ;
        RECT 103.980 146.900 104.630 147.550 ;
        RECT 11.630 140.100 12.280 140.750 ;
        RECT 12.430 140.100 13.080 140.750 ;
        RECT 13.230 140.100 13.880 140.750 ;
        RECT 15.580 140.100 16.230 140.750 ;
        RECT 16.380 140.100 17.030 140.750 ;
        RECT 17.180 140.100 17.830 140.750 ;
        RECT 11.630 139.250 12.280 139.900 ;
        RECT 12.430 139.250 13.080 139.900 ;
        RECT 13.230 139.250 13.880 139.900 ;
        RECT 15.580 139.250 16.230 139.900 ;
        RECT 16.380 139.250 17.030 139.900 ;
        RECT 17.180 139.250 17.830 139.900 ;
        RECT 31.630 140.100 32.280 140.750 ;
        RECT 32.430 140.100 33.080 140.750 ;
        RECT 33.230 140.100 33.880 140.750 ;
        RECT 35.580 140.100 36.230 140.750 ;
        RECT 36.380 140.100 37.030 140.750 ;
        RECT 37.180 140.100 37.830 140.750 ;
        RECT 31.630 139.250 32.280 139.900 ;
        RECT 32.430 139.250 33.080 139.900 ;
        RECT 33.230 139.250 33.880 139.900 ;
        RECT 35.580 139.250 36.230 139.900 ;
        RECT 36.380 139.250 37.030 139.900 ;
        RECT 37.180 139.250 37.830 139.900 ;
        RECT 51.630 140.100 52.280 140.750 ;
        RECT 52.430 140.100 53.080 140.750 ;
        RECT 53.230 140.100 53.880 140.750 ;
        RECT 55.580 140.100 56.230 140.750 ;
        RECT 56.380 140.100 57.030 140.750 ;
        RECT 57.180 140.100 57.830 140.750 ;
        RECT 51.630 139.250 52.280 139.900 ;
        RECT 52.430 139.250 53.080 139.900 ;
        RECT 53.230 139.250 53.880 139.900 ;
        RECT 55.580 139.250 56.230 139.900 ;
        RECT 56.380 139.250 57.030 139.900 ;
        RECT 57.180 139.250 57.830 139.900 ;
        RECT 71.630 140.100 72.280 140.750 ;
        RECT 72.430 140.100 73.080 140.750 ;
        RECT 73.230 140.100 73.880 140.750 ;
        RECT 75.580 140.100 76.230 140.750 ;
        RECT 76.380 140.100 77.030 140.750 ;
        RECT 77.180 140.100 77.830 140.750 ;
        RECT 71.630 139.250 72.280 139.900 ;
        RECT 72.430 139.250 73.080 139.900 ;
        RECT 73.230 139.250 73.880 139.900 ;
        RECT 75.580 139.250 76.230 139.900 ;
        RECT 76.380 139.250 77.030 139.900 ;
        RECT 77.180 139.250 77.830 139.900 ;
        RECT 91.630 140.100 92.280 140.750 ;
        RECT 92.430 140.100 93.080 140.750 ;
        RECT 93.230 140.100 93.880 140.750 ;
        RECT 95.580 140.100 96.230 140.750 ;
        RECT 96.380 140.100 97.030 140.750 ;
        RECT 97.180 140.100 97.830 140.750 ;
        RECT 91.630 139.250 92.280 139.900 ;
        RECT 92.430 139.250 93.080 139.900 ;
        RECT 93.230 139.250 93.880 139.900 ;
        RECT 95.580 139.250 96.230 139.900 ;
        RECT 96.380 139.250 97.030 139.900 ;
        RECT 97.180 139.250 97.830 139.900 ;
        RECT 4.830 132.450 5.480 133.100 ;
        RECT 4.830 131.650 5.480 132.300 ;
        RECT 4.830 130.850 5.480 131.500 ;
        RECT 4.830 128.500 5.480 129.150 ;
        RECT 4.830 127.700 5.480 128.350 ;
        RECT 4.830 126.900 5.480 127.550 ;
        RECT 23.980 132.450 24.630 133.100 ;
        RECT 24.830 132.450 25.480 133.100 ;
        RECT 23.980 131.650 24.630 132.300 ;
        RECT 24.830 131.650 25.480 132.300 ;
        RECT 23.980 130.850 24.630 131.500 ;
        RECT 24.830 130.850 25.480 131.500 ;
        RECT 23.980 128.500 24.630 129.150 ;
        RECT 24.830 128.500 25.480 129.150 ;
        RECT 23.980 127.700 24.630 128.350 ;
        RECT 24.830 127.700 25.480 128.350 ;
        RECT 23.980 126.900 24.630 127.550 ;
        RECT 24.830 126.900 25.480 127.550 ;
        RECT 43.980 132.450 44.630 133.100 ;
        RECT 44.830 132.450 45.480 133.100 ;
        RECT 43.980 131.650 44.630 132.300 ;
        RECT 44.830 131.650 45.480 132.300 ;
        RECT 43.980 130.850 44.630 131.500 ;
        RECT 44.830 130.850 45.480 131.500 ;
        RECT 43.980 128.500 44.630 129.150 ;
        RECT 44.830 128.500 45.480 129.150 ;
        RECT 43.980 127.700 44.630 128.350 ;
        RECT 44.830 127.700 45.480 128.350 ;
        RECT 43.980 126.900 44.630 127.550 ;
        RECT 44.830 126.900 45.480 127.550 ;
        RECT 63.980 132.450 64.630 133.100 ;
        RECT 64.830 132.450 65.480 133.100 ;
        RECT 63.980 131.650 64.630 132.300 ;
        RECT 64.830 131.650 65.480 132.300 ;
        RECT 63.980 130.850 64.630 131.500 ;
        RECT 64.830 130.850 65.480 131.500 ;
        RECT 63.980 128.500 64.630 129.150 ;
        RECT 64.830 128.500 65.480 129.150 ;
        RECT 63.980 127.700 64.630 128.350 ;
        RECT 64.830 127.700 65.480 128.350 ;
        RECT 63.980 126.900 64.630 127.550 ;
        RECT 64.830 126.900 65.480 127.550 ;
        RECT 83.980 132.450 84.630 133.100 ;
        RECT 84.830 132.450 85.480 133.100 ;
        RECT 83.980 131.650 84.630 132.300 ;
        RECT 84.830 131.650 85.480 132.300 ;
        RECT 83.980 130.850 84.630 131.500 ;
        RECT 84.830 130.850 85.480 131.500 ;
        RECT 83.980 128.500 84.630 129.150 ;
        RECT 84.830 128.500 85.480 129.150 ;
        RECT 83.980 127.700 84.630 128.350 ;
        RECT 84.830 127.700 85.480 128.350 ;
        RECT 83.980 126.900 84.630 127.550 ;
        RECT 84.830 126.900 85.480 127.550 ;
        RECT 103.980 132.450 104.630 133.100 ;
        RECT 103.980 131.650 104.630 132.300 ;
        RECT 103.980 130.850 104.630 131.500 ;
        RECT 103.980 128.500 104.630 129.150 ;
        RECT 103.980 127.700 104.630 128.350 ;
        RECT 103.980 126.900 104.630 127.550 ;
        RECT 11.630 120.100 12.280 120.750 ;
        RECT 12.430 120.100 13.080 120.750 ;
        RECT 13.230 120.100 13.880 120.750 ;
        RECT 15.580 120.100 16.230 120.750 ;
        RECT 16.380 120.100 17.030 120.750 ;
        RECT 17.180 120.100 17.830 120.750 ;
        RECT 11.630 119.250 12.280 119.900 ;
        RECT 12.430 119.250 13.080 119.900 ;
        RECT 13.230 119.250 13.880 119.900 ;
        RECT 15.580 119.250 16.230 119.900 ;
        RECT 16.380 119.250 17.030 119.900 ;
        RECT 17.180 119.250 17.830 119.900 ;
        RECT 31.630 120.100 32.280 120.750 ;
        RECT 32.430 120.100 33.080 120.750 ;
        RECT 33.230 120.100 33.880 120.750 ;
        RECT 35.580 120.100 36.230 120.750 ;
        RECT 36.380 120.100 37.030 120.750 ;
        RECT 37.180 120.100 37.830 120.750 ;
        RECT 31.630 119.250 32.280 119.900 ;
        RECT 32.430 119.250 33.080 119.900 ;
        RECT 33.230 119.250 33.880 119.900 ;
        RECT 35.580 119.250 36.230 119.900 ;
        RECT 36.380 119.250 37.030 119.900 ;
        RECT 37.180 119.250 37.830 119.900 ;
        RECT 51.630 120.100 52.280 120.750 ;
        RECT 52.430 120.100 53.080 120.750 ;
        RECT 53.230 120.100 53.880 120.750 ;
        RECT 55.580 120.100 56.230 120.750 ;
        RECT 56.380 120.100 57.030 120.750 ;
        RECT 57.180 120.100 57.830 120.750 ;
        RECT 51.630 119.250 52.280 119.900 ;
        RECT 52.430 119.250 53.080 119.900 ;
        RECT 53.230 119.250 53.880 119.900 ;
        RECT 55.580 119.250 56.230 119.900 ;
        RECT 56.380 119.250 57.030 119.900 ;
        RECT 57.180 119.250 57.830 119.900 ;
        RECT 71.630 120.100 72.280 120.750 ;
        RECT 72.430 120.100 73.080 120.750 ;
        RECT 73.230 120.100 73.880 120.750 ;
        RECT 75.580 120.100 76.230 120.750 ;
        RECT 76.380 120.100 77.030 120.750 ;
        RECT 77.180 120.100 77.830 120.750 ;
        RECT 71.630 119.250 72.280 119.900 ;
        RECT 72.430 119.250 73.080 119.900 ;
        RECT 73.230 119.250 73.880 119.900 ;
        RECT 75.580 119.250 76.230 119.900 ;
        RECT 76.380 119.250 77.030 119.900 ;
        RECT 77.180 119.250 77.830 119.900 ;
        RECT 91.630 120.100 92.280 120.750 ;
        RECT 92.430 120.100 93.080 120.750 ;
        RECT 93.230 120.100 93.880 120.750 ;
        RECT 95.580 120.100 96.230 120.750 ;
        RECT 96.380 120.100 97.030 120.750 ;
        RECT 97.180 120.100 97.830 120.750 ;
        RECT 91.630 119.250 92.280 119.900 ;
        RECT 92.430 119.250 93.080 119.900 ;
        RECT 93.230 119.250 93.880 119.900 ;
        RECT 95.580 119.250 96.230 119.900 ;
        RECT 96.380 119.250 97.030 119.900 ;
        RECT 97.180 119.250 97.830 119.900 ;
        RECT 4.830 112.450 5.480 113.100 ;
        RECT 4.830 111.650 5.480 112.300 ;
        RECT 4.830 110.850 5.480 111.500 ;
        RECT 4.830 108.500 5.480 109.150 ;
        RECT 4.830 107.700 5.480 108.350 ;
        RECT 4.830 106.900 5.480 107.550 ;
        RECT 23.980 112.450 24.630 113.100 ;
        RECT 24.830 112.450 25.480 113.100 ;
        RECT 23.980 111.650 24.630 112.300 ;
        RECT 24.830 111.650 25.480 112.300 ;
        RECT 23.980 110.850 24.630 111.500 ;
        RECT 24.830 110.850 25.480 111.500 ;
        RECT 23.980 108.500 24.630 109.150 ;
        RECT 24.830 108.500 25.480 109.150 ;
        RECT 23.980 107.700 24.630 108.350 ;
        RECT 24.830 107.700 25.480 108.350 ;
        RECT 23.980 106.900 24.630 107.550 ;
        RECT 24.830 106.900 25.480 107.550 ;
        RECT 43.980 112.450 44.630 113.100 ;
        RECT 44.830 112.450 45.480 113.100 ;
        RECT 43.980 111.650 44.630 112.300 ;
        RECT 44.830 111.650 45.480 112.300 ;
        RECT 43.980 110.850 44.630 111.500 ;
        RECT 44.830 110.850 45.480 111.500 ;
        RECT 43.980 108.500 44.630 109.150 ;
        RECT 44.830 108.500 45.480 109.150 ;
        RECT 43.980 107.700 44.630 108.350 ;
        RECT 44.830 107.700 45.480 108.350 ;
        RECT 43.980 106.900 44.630 107.550 ;
        RECT 44.830 106.900 45.480 107.550 ;
        RECT 63.980 112.450 64.630 113.100 ;
        RECT 64.830 112.450 65.480 113.100 ;
        RECT 63.980 111.650 64.630 112.300 ;
        RECT 64.830 111.650 65.480 112.300 ;
        RECT 63.980 110.850 64.630 111.500 ;
        RECT 64.830 110.850 65.480 111.500 ;
        RECT 63.980 108.500 64.630 109.150 ;
        RECT 64.830 108.500 65.480 109.150 ;
        RECT 63.980 107.700 64.630 108.350 ;
        RECT 64.830 107.700 65.480 108.350 ;
        RECT 63.980 106.900 64.630 107.550 ;
        RECT 64.830 106.900 65.480 107.550 ;
        RECT 83.980 112.450 84.630 113.100 ;
        RECT 84.830 112.450 85.480 113.100 ;
        RECT 83.980 111.650 84.630 112.300 ;
        RECT 84.830 111.650 85.480 112.300 ;
        RECT 83.980 110.850 84.630 111.500 ;
        RECT 84.830 110.850 85.480 111.500 ;
        RECT 83.980 108.500 84.630 109.150 ;
        RECT 84.830 108.500 85.480 109.150 ;
        RECT 83.980 107.700 84.630 108.350 ;
        RECT 84.830 107.700 85.480 108.350 ;
        RECT 83.980 106.900 84.630 107.550 ;
        RECT 84.830 106.900 85.480 107.550 ;
        RECT 103.980 112.450 104.630 113.100 ;
        RECT 103.980 111.650 104.630 112.300 ;
        RECT 103.980 110.850 104.630 111.500 ;
        RECT 103.980 108.500 104.630 109.150 ;
        RECT 103.980 107.700 104.630 108.350 ;
        RECT 103.980 106.900 104.630 107.550 ;
        RECT 11.630 100.100 12.280 100.750 ;
        RECT 12.430 100.100 13.080 100.750 ;
        RECT 13.230 100.100 13.880 100.750 ;
        RECT 15.580 100.100 16.230 100.750 ;
        RECT 16.380 100.100 17.030 100.750 ;
        RECT 17.180 100.100 17.830 100.750 ;
        RECT 11.630 99.250 12.280 99.900 ;
        RECT 12.430 99.250 13.080 99.900 ;
        RECT 13.230 99.250 13.880 99.900 ;
        RECT 15.580 99.250 16.230 99.900 ;
        RECT 16.380 99.250 17.030 99.900 ;
        RECT 17.180 99.250 17.830 99.900 ;
        RECT 31.630 100.100 32.280 100.750 ;
        RECT 32.430 100.100 33.080 100.750 ;
        RECT 33.230 100.100 33.880 100.750 ;
        RECT 35.580 100.100 36.230 100.750 ;
        RECT 36.380 100.100 37.030 100.750 ;
        RECT 37.180 100.100 37.830 100.750 ;
        RECT 31.630 99.250 32.280 99.900 ;
        RECT 32.430 99.250 33.080 99.900 ;
        RECT 33.230 99.250 33.880 99.900 ;
        RECT 35.580 99.250 36.230 99.900 ;
        RECT 36.380 99.250 37.030 99.900 ;
        RECT 37.180 99.250 37.830 99.900 ;
        RECT 51.630 100.100 52.280 100.750 ;
        RECT 52.430 100.100 53.080 100.750 ;
        RECT 53.230 100.100 53.880 100.750 ;
        RECT 55.580 100.100 56.230 100.750 ;
        RECT 56.380 100.100 57.030 100.750 ;
        RECT 57.180 100.100 57.830 100.750 ;
        RECT 51.630 99.250 52.280 99.900 ;
        RECT 52.430 99.250 53.080 99.900 ;
        RECT 53.230 99.250 53.880 99.900 ;
        RECT 55.580 99.250 56.230 99.900 ;
        RECT 56.380 99.250 57.030 99.900 ;
        RECT 57.180 99.250 57.830 99.900 ;
        RECT 71.630 100.100 72.280 100.750 ;
        RECT 72.430 100.100 73.080 100.750 ;
        RECT 73.230 100.100 73.880 100.750 ;
        RECT 75.580 100.100 76.230 100.750 ;
        RECT 76.380 100.100 77.030 100.750 ;
        RECT 77.180 100.100 77.830 100.750 ;
        RECT 71.630 99.250 72.280 99.900 ;
        RECT 72.430 99.250 73.080 99.900 ;
        RECT 73.230 99.250 73.880 99.900 ;
        RECT 75.580 99.250 76.230 99.900 ;
        RECT 76.380 99.250 77.030 99.900 ;
        RECT 77.180 99.250 77.830 99.900 ;
        RECT 91.630 100.100 92.280 100.750 ;
        RECT 92.430 100.100 93.080 100.750 ;
        RECT 93.230 100.100 93.880 100.750 ;
        RECT 95.580 100.100 96.230 100.750 ;
        RECT 96.380 100.100 97.030 100.750 ;
        RECT 97.180 100.100 97.830 100.750 ;
        RECT 91.630 99.250 92.280 99.900 ;
        RECT 92.430 99.250 93.080 99.900 ;
        RECT 93.230 99.250 93.880 99.900 ;
        RECT 95.580 99.250 96.230 99.900 ;
        RECT 96.380 99.250 97.030 99.900 ;
        RECT 97.180 99.250 97.830 99.900 ;
        RECT 4.830 92.450 5.480 93.100 ;
        RECT 4.830 91.650 5.480 92.300 ;
        RECT 4.830 90.850 5.480 91.500 ;
        RECT 4.830 88.500 5.480 89.150 ;
        RECT 4.830 87.700 5.480 88.350 ;
        RECT 4.830 86.900 5.480 87.550 ;
        RECT 23.980 92.450 24.630 93.100 ;
        RECT 24.830 92.450 25.480 93.100 ;
        RECT 23.980 91.650 24.630 92.300 ;
        RECT 24.830 91.650 25.480 92.300 ;
        RECT 23.980 90.850 24.630 91.500 ;
        RECT 24.830 90.850 25.480 91.500 ;
        RECT 23.980 88.500 24.630 89.150 ;
        RECT 24.830 88.500 25.480 89.150 ;
        RECT 23.980 87.700 24.630 88.350 ;
        RECT 24.830 87.700 25.480 88.350 ;
        RECT 23.980 86.900 24.630 87.550 ;
        RECT 24.830 86.900 25.480 87.550 ;
        RECT 43.980 92.450 44.630 93.100 ;
        RECT 44.830 92.450 45.480 93.100 ;
        RECT 43.980 91.650 44.630 92.300 ;
        RECT 44.830 91.650 45.480 92.300 ;
        RECT 43.980 90.850 44.630 91.500 ;
        RECT 44.830 90.850 45.480 91.500 ;
        RECT 43.980 88.500 44.630 89.150 ;
        RECT 44.830 88.500 45.480 89.150 ;
        RECT 43.980 87.700 44.630 88.350 ;
        RECT 44.830 87.700 45.480 88.350 ;
        RECT 43.980 86.900 44.630 87.550 ;
        RECT 44.830 86.900 45.480 87.550 ;
        RECT 63.980 92.450 64.630 93.100 ;
        RECT 64.830 92.450 65.480 93.100 ;
        RECT 63.980 91.650 64.630 92.300 ;
        RECT 64.830 91.650 65.480 92.300 ;
        RECT 63.980 90.850 64.630 91.500 ;
        RECT 64.830 90.850 65.480 91.500 ;
        RECT 63.980 88.500 64.630 89.150 ;
        RECT 64.830 88.500 65.480 89.150 ;
        RECT 63.980 87.700 64.630 88.350 ;
        RECT 64.830 87.700 65.480 88.350 ;
        RECT 63.980 86.900 64.630 87.550 ;
        RECT 64.830 86.900 65.480 87.550 ;
        RECT 83.980 92.450 84.630 93.100 ;
        RECT 84.830 92.450 85.480 93.100 ;
        RECT 83.980 91.650 84.630 92.300 ;
        RECT 84.830 91.650 85.480 92.300 ;
        RECT 83.980 90.850 84.630 91.500 ;
        RECT 84.830 90.850 85.480 91.500 ;
        RECT 83.980 88.500 84.630 89.150 ;
        RECT 84.830 88.500 85.480 89.150 ;
        RECT 83.980 87.700 84.630 88.350 ;
        RECT 84.830 87.700 85.480 88.350 ;
        RECT 83.980 86.900 84.630 87.550 ;
        RECT 84.830 86.900 85.480 87.550 ;
        RECT 103.980 92.450 104.630 93.100 ;
        RECT 103.980 91.650 104.630 92.300 ;
        RECT 103.980 90.850 104.630 91.500 ;
        RECT 103.980 88.500 104.630 89.150 ;
        RECT 103.980 87.700 104.630 88.350 ;
        RECT 103.980 86.900 104.630 87.550 ;
        RECT 11.630 80.100 12.280 80.750 ;
        RECT 12.430 80.100 13.080 80.750 ;
        RECT 13.230 80.100 13.880 80.750 ;
        RECT 15.580 80.100 16.230 80.750 ;
        RECT 16.380 80.100 17.030 80.750 ;
        RECT 17.180 80.100 17.830 80.750 ;
        RECT 11.630 79.250 12.280 79.900 ;
        RECT 12.430 79.250 13.080 79.900 ;
        RECT 13.230 79.250 13.880 79.900 ;
        RECT 15.580 79.250 16.230 79.900 ;
        RECT 16.380 79.250 17.030 79.900 ;
        RECT 17.180 79.250 17.830 79.900 ;
        RECT 31.630 80.100 32.280 80.750 ;
        RECT 32.430 80.100 33.080 80.750 ;
        RECT 33.230 80.100 33.880 80.750 ;
        RECT 35.580 80.100 36.230 80.750 ;
        RECT 36.380 80.100 37.030 80.750 ;
        RECT 37.180 80.100 37.830 80.750 ;
        RECT 31.630 79.250 32.280 79.900 ;
        RECT 32.430 79.250 33.080 79.900 ;
        RECT 33.230 79.250 33.880 79.900 ;
        RECT 35.580 79.250 36.230 79.900 ;
        RECT 36.380 79.250 37.030 79.900 ;
        RECT 37.180 79.250 37.830 79.900 ;
        RECT 51.630 80.100 52.280 80.750 ;
        RECT 52.430 80.100 53.080 80.750 ;
        RECT 53.230 80.100 53.880 80.750 ;
        RECT 55.580 80.100 56.230 80.750 ;
        RECT 56.380 80.100 57.030 80.750 ;
        RECT 57.180 80.100 57.830 80.750 ;
        RECT 51.630 79.250 52.280 79.900 ;
        RECT 52.430 79.250 53.080 79.900 ;
        RECT 53.230 79.250 53.880 79.900 ;
        RECT 55.580 79.250 56.230 79.900 ;
        RECT 56.380 79.250 57.030 79.900 ;
        RECT 57.180 79.250 57.830 79.900 ;
        RECT 71.630 80.100 72.280 80.750 ;
        RECT 72.430 80.100 73.080 80.750 ;
        RECT 73.230 80.100 73.880 80.750 ;
        RECT 75.580 80.100 76.230 80.750 ;
        RECT 76.380 80.100 77.030 80.750 ;
        RECT 77.180 80.100 77.830 80.750 ;
        RECT 71.630 79.250 72.280 79.900 ;
        RECT 72.430 79.250 73.080 79.900 ;
        RECT 73.230 79.250 73.880 79.900 ;
        RECT 75.580 79.250 76.230 79.900 ;
        RECT 76.380 79.250 77.030 79.900 ;
        RECT 77.180 79.250 77.830 79.900 ;
        RECT 91.630 80.100 92.280 80.750 ;
        RECT 92.430 80.100 93.080 80.750 ;
        RECT 93.230 80.100 93.880 80.750 ;
        RECT 95.580 80.100 96.230 80.750 ;
        RECT 96.380 80.100 97.030 80.750 ;
        RECT 97.180 80.100 97.830 80.750 ;
        RECT 91.630 79.250 92.280 79.900 ;
        RECT 92.430 79.250 93.080 79.900 ;
        RECT 93.230 79.250 93.880 79.900 ;
        RECT 95.580 79.250 96.230 79.900 ;
        RECT 96.380 79.250 97.030 79.900 ;
        RECT 97.180 79.250 97.830 79.900 ;
        RECT 4.830 72.450 5.480 73.100 ;
        RECT 4.830 71.650 5.480 72.300 ;
        RECT 4.830 70.850 5.480 71.500 ;
        RECT 4.830 68.500 5.480 69.150 ;
        RECT 4.830 67.700 5.480 68.350 ;
        RECT 4.830 66.900 5.480 67.550 ;
        RECT 23.980 72.450 24.630 73.100 ;
        RECT 24.830 72.450 25.480 73.100 ;
        RECT 23.980 71.650 24.630 72.300 ;
        RECT 24.830 71.650 25.480 72.300 ;
        RECT 23.980 70.850 24.630 71.500 ;
        RECT 24.830 70.850 25.480 71.500 ;
        RECT 23.980 68.500 24.630 69.150 ;
        RECT 24.830 68.500 25.480 69.150 ;
        RECT 23.980 67.700 24.630 68.350 ;
        RECT 24.830 67.700 25.480 68.350 ;
        RECT 23.980 66.900 24.630 67.550 ;
        RECT 24.830 66.900 25.480 67.550 ;
        RECT 43.980 72.450 44.630 73.100 ;
        RECT 44.830 72.450 45.480 73.100 ;
        RECT 43.980 71.650 44.630 72.300 ;
        RECT 44.830 71.650 45.480 72.300 ;
        RECT 43.980 70.850 44.630 71.500 ;
        RECT 44.830 70.850 45.480 71.500 ;
        RECT 43.980 68.500 44.630 69.150 ;
        RECT 44.830 68.500 45.480 69.150 ;
        RECT 43.980 67.700 44.630 68.350 ;
        RECT 44.830 67.700 45.480 68.350 ;
        RECT 43.980 66.900 44.630 67.550 ;
        RECT 44.830 66.900 45.480 67.550 ;
        RECT 63.980 72.450 64.630 73.100 ;
        RECT 64.830 72.450 65.480 73.100 ;
        RECT 63.980 71.650 64.630 72.300 ;
        RECT 64.830 71.650 65.480 72.300 ;
        RECT 63.980 70.850 64.630 71.500 ;
        RECT 64.830 70.850 65.480 71.500 ;
        RECT 63.980 68.500 64.630 69.150 ;
        RECT 64.830 68.500 65.480 69.150 ;
        RECT 63.980 67.700 64.630 68.350 ;
        RECT 64.830 67.700 65.480 68.350 ;
        RECT 63.980 66.900 64.630 67.550 ;
        RECT 64.830 66.900 65.480 67.550 ;
        RECT 83.980 72.450 84.630 73.100 ;
        RECT 84.830 72.450 85.480 73.100 ;
        RECT 83.980 71.650 84.630 72.300 ;
        RECT 84.830 71.650 85.480 72.300 ;
        RECT 83.980 70.850 84.630 71.500 ;
        RECT 84.830 70.850 85.480 71.500 ;
        RECT 83.980 68.500 84.630 69.150 ;
        RECT 84.830 68.500 85.480 69.150 ;
        RECT 83.980 67.700 84.630 68.350 ;
        RECT 84.830 67.700 85.480 68.350 ;
        RECT 83.980 66.900 84.630 67.550 ;
        RECT 84.830 66.900 85.480 67.550 ;
        RECT 103.980 72.450 104.630 73.100 ;
        RECT 103.980 71.650 104.630 72.300 ;
        RECT 103.980 70.850 104.630 71.500 ;
        RECT 103.980 68.500 104.630 69.150 ;
        RECT 103.980 67.700 104.630 68.350 ;
        RECT 103.980 66.900 104.630 67.550 ;
        RECT 11.630 60.100 12.280 60.750 ;
        RECT 12.430 60.100 13.080 60.750 ;
        RECT 13.230 60.100 13.880 60.750 ;
        RECT 15.580 60.100 16.230 60.750 ;
        RECT 16.380 60.100 17.030 60.750 ;
        RECT 17.180 60.100 17.830 60.750 ;
        RECT 11.630 59.250 12.280 59.900 ;
        RECT 12.430 59.250 13.080 59.900 ;
        RECT 13.230 59.250 13.880 59.900 ;
        RECT 15.580 59.250 16.230 59.900 ;
        RECT 16.380 59.250 17.030 59.900 ;
        RECT 17.180 59.250 17.830 59.900 ;
        RECT 31.630 60.100 32.280 60.750 ;
        RECT 32.430 60.100 33.080 60.750 ;
        RECT 33.230 60.100 33.880 60.750 ;
        RECT 35.580 60.100 36.230 60.750 ;
        RECT 36.380 60.100 37.030 60.750 ;
        RECT 37.180 60.100 37.830 60.750 ;
        RECT 31.630 59.250 32.280 59.900 ;
        RECT 32.430 59.250 33.080 59.900 ;
        RECT 33.230 59.250 33.880 59.900 ;
        RECT 35.580 59.250 36.230 59.900 ;
        RECT 36.380 59.250 37.030 59.900 ;
        RECT 37.180 59.250 37.830 59.900 ;
        RECT 51.630 60.100 52.280 60.750 ;
        RECT 52.430 60.100 53.080 60.750 ;
        RECT 53.230 60.100 53.880 60.750 ;
        RECT 55.580 60.100 56.230 60.750 ;
        RECT 56.380 60.100 57.030 60.750 ;
        RECT 57.180 60.100 57.830 60.750 ;
        RECT 51.630 59.250 52.280 59.900 ;
        RECT 52.430 59.250 53.080 59.900 ;
        RECT 53.230 59.250 53.880 59.900 ;
        RECT 55.580 59.250 56.230 59.900 ;
        RECT 56.380 59.250 57.030 59.900 ;
        RECT 57.180 59.250 57.830 59.900 ;
        RECT 71.630 60.100 72.280 60.750 ;
        RECT 72.430 60.100 73.080 60.750 ;
        RECT 73.230 60.100 73.880 60.750 ;
        RECT 75.580 60.100 76.230 60.750 ;
        RECT 76.380 60.100 77.030 60.750 ;
        RECT 77.180 60.100 77.830 60.750 ;
        RECT 71.630 59.250 72.280 59.900 ;
        RECT 72.430 59.250 73.080 59.900 ;
        RECT 73.230 59.250 73.880 59.900 ;
        RECT 75.580 59.250 76.230 59.900 ;
        RECT 76.380 59.250 77.030 59.900 ;
        RECT 77.180 59.250 77.830 59.900 ;
        RECT 91.630 60.100 92.280 60.750 ;
        RECT 92.430 60.100 93.080 60.750 ;
        RECT 93.230 60.100 93.880 60.750 ;
        RECT 95.580 60.100 96.230 60.750 ;
        RECT 96.380 60.100 97.030 60.750 ;
        RECT 97.180 60.100 97.830 60.750 ;
        RECT 91.630 59.250 92.280 59.900 ;
        RECT 92.430 59.250 93.080 59.900 ;
        RECT 93.230 59.250 93.880 59.900 ;
        RECT 95.580 59.250 96.230 59.900 ;
        RECT 96.380 59.250 97.030 59.900 ;
        RECT 97.180 59.250 97.830 59.900 ;
        RECT 4.830 52.450 5.480 53.100 ;
        RECT 4.830 51.650 5.480 52.300 ;
        RECT 4.830 50.850 5.480 51.500 ;
        RECT 4.830 48.500 5.480 49.150 ;
        RECT 4.830 47.700 5.480 48.350 ;
        RECT 4.830 46.900 5.480 47.550 ;
        RECT 23.980 52.450 24.630 53.100 ;
        RECT 24.830 52.450 25.480 53.100 ;
        RECT 23.980 51.650 24.630 52.300 ;
        RECT 24.830 51.650 25.480 52.300 ;
        RECT 23.980 50.850 24.630 51.500 ;
        RECT 24.830 50.850 25.480 51.500 ;
        RECT 23.980 48.500 24.630 49.150 ;
        RECT 24.830 48.500 25.480 49.150 ;
        RECT 23.980 47.700 24.630 48.350 ;
        RECT 24.830 47.700 25.480 48.350 ;
        RECT 23.980 46.900 24.630 47.550 ;
        RECT 24.830 46.900 25.480 47.550 ;
        RECT 43.980 52.450 44.630 53.100 ;
        RECT 44.830 52.450 45.480 53.100 ;
        RECT 43.980 51.650 44.630 52.300 ;
        RECT 44.830 51.650 45.480 52.300 ;
        RECT 43.980 50.850 44.630 51.500 ;
        RECT 44.830 50.850 45.480 51.500 ;
        RECT 43.980 48.500 44.630 49.150 ;
        RECT 44.830 48.500 45.480 49.150 ;
        RECT 43.980 47.700 44.630 48.350 ;
        RECT 44.830 47.700 45.480 48.350 ;
        RECT 43.980 46.900 44.630 47.550 ;
        RECT 44.830 46.900 45.480 47.550 ;
        RECT 63.980 52.450 64.630 53.100 ;
        RECT 64.830 52.450 65.480 53.100 ;
        RECT 63.980 51.650 64.630 52.300 ;
        RECT 64.830 51.650 65.480 52.300 ;
        RECT 63.980 50.850 64.630 51.500 ;
        RECT 64.830 50.850 65.480 51.500 ;
        RECT 63.980 48.500 64.630 49.150 ;
        RECT 64.830 48.500 65.480 49.150 ;
        RECT 63.980 47.700 64.630 48.350 ;
        RECT 64.830 47.700 65.480 48.350 ;
        RECT 63.980 46.900 64.630 47.550 ;
        RECT 64.830 46.900 65.480 47.550 ;
        RECT 83.980 52.450 84.630 53.100 ;
        RECT 84.830 52.450 85.480 53.100 ;
        RECT 83.980 51.650 84.630 52.300 ;
        RECT 84.830 51.650 85.480 52.300 ;
        RECT 83.980 50.850 84.630 51.500 ;
        RECT 84.830 50.850 85.480 51.500 ;
        RECT 83.980 48.500 84.630 49.150 ;
        RECT 84.830 48.500 85.480 49.150 ;
        RECT 83.980 47.700 84.630 48.350 ;
        RECT 84.830 47.700 85.480 48.350 ;
        RECT 83.980 46.900 84.630 47.550 ;
        RECT 84.830 46.900 85.480 47.550 ;
        RECT 103.980 52.450 104.630 53.100 ;
        RECT 103.980 51.650 104.630 52.300 ;
        RECT 103.980 50.850 104.630 51.500 ;
        RECT 103.980 48.500 104.630 49.150 ;
        RECT 103.980 47.700 104.630 48.350 ;
        RECT 103.980 46.900 104.630 47.550 ;
        RECT 11.630 40.100 12.280 40.750 ;
        RECT 12.430 40.100 13.080 40.750 ;
        RECT 13.230 40.100 13.880 40.750 ;
        RECT 15.580 40.100 16.230 40.750 ;
        RECT 16.380 40.100 17.030 40.750 ;
        RECT 17.180 40.100 17.830 40.750 ;
        RECT 11.630 39.250 12.280 39.900 ;
        RECT 12.430 39.250 13.080 39.900 ;
        RECT 13.230 39.250 13.880 39.900 ;
        RECT 15.580 39.250 16.230 39.900 ;
        RECT 16.380 39.250 17.030 39.900 ;
        RECT 17.180 39.250 17.830 39.900 ;
        RECT 31.630 40.100 32.280 40.750 ;
        RECT 32.430 40.100 33.080 40.750 ;
        RECT 33.230 40.100 33.880 40.750 ;
        RECT 35.580 40.100 36.230 40.750 ;
        RECT 36.380 40.100 37.030 40.750 ;
        RECT 37.180 40.100 37.830 40.750 ;
        RECT 31.630 39.250 32.280 39.900 ;
        RECT 32.430 39.250 33.080 39.900 ;
        RECT 33.230 39.250 33.880 39.900 ;
        RECT 35.580 39.250 36.230 39.900 ;
        RECT 36.380 39.250 37.030 39.900 ;
        RECT 37.180 39.250 37.830 39.900 ;
        RECT 51.630 40.100 52.280 40.750 ;
        RECT 52.430 40.100 53.080 40.750 ;
        RECT 53.230 40.100 53.880 40.750 ;
        RECT 55.580 40.100 56.230 40.750 ;
        RECT 56.380 40.100 57.030 40.750 ;
        RECT 57.180 40.100 57.830 40.750 ;
        RECT 51.630 39.250 52.280 39.900 ;
        RECT 52.430 39.250 53.080 39.900 ;
        RECT 53.230 39.250 53.880 39.900 ;
        RECT 55.580 39.250 56.230 39.900 ;
        RECT 56.380 39.250 57.030 39.900 ;
        RECT 57.180 39.250 57.830 39.900 ;
        RECT 71.630 40.100 72.280 40.750 ;
        RECT 72.430 40.100 73.080 40.750 ;
        RECT 73.230 40.100 73.880 40.750 ;
        RECT 75.580 40.100 76.230 40.750 ;
        RECT 76.380 40.100 77.030 40.750 ;
        RECT 77.180 40.100 77.830 40.750 ;
        RECT 71.630 39.250 72.280 39.900 ;
        RECT 72.430 39.250 73.080 39.900 ;
        RECT 73.230 39.250 73.880 39.900 ;
        RECT 75.580 39.250 76.230 39.900 ;
        RECT 76.380 39.250 77.030 39.900 ;
        RECT 77.180 39.250 77.830 39.900 ;
        RECT 91.630 40.100 92.280 40.750 ;
        RECT 92.430 40.100 93.080 40.750 ;
        RECT 93.230 40.100 93.880 40.750 ;
        RECT 95.580 40.100 96.230 40.750 ;
        RECT 96.380 40.100 97.030 40.750 ;
        RECT 97.180 40.100 97.830 40.750 ;
        RECT 91.630 39.250 92.280 39.900 ;
        RECT 92.430 39.250 93.080 39.900 ;
        RECT 93.230 39.250 93.880 39.900 ;
        RECT 95.580 39.250 96.230 39.900 ;
        RECT 96.380 39.250 97.030 39.900 ;
        RECT 97.180 39.250 97.830 39.900 ;
        RECT 4.830 32.450 5.480 33.100 ;
        RECT 4.830 31.650 5.480 32.300 ;
        RECT 4.830 30.850 5.480 31.500 ;
        RECT 4.830 28.500 5.480 29.150 ;
        RECT 4.830 27.700 5.480 28.350 ;
        RECT 4.830 26.900 5.480 27.550 ;
        RECT 23.980 32.450 24.630 33.100 ;
        RECT 24.830 32.450 25.480 33.100 ;
        RECT 23.980 31.650 24.630 32.300 ;
        RECT 24.830 31.650 25.480 32.300 ;
        RECT 23.980 30.850 24.630 31.500 ;
        RECT 24.830 30.850 25.480 31.500 ;
        RECT 23.980 28.500 24.630 29.150 ;
        RECT 24.830 28.500 25.480 29.150 ;
        RECT 23.980 27.700 24.630 28.350 ;
        RECT 24.830 27.700 25.480 28.350 ;
        RECT 23.980 26.900 24.630 27.550 ;
        RECT 24.830 26.900 25.480 27.550 ;
        RECT 43.980 32.450 44.630 33.100 ;
        RECT 44.830 32.450 45.480 33.100 ;
        RECT 43.980 31.650 44.630 32.300 ;
        RECT 44.830 31.650 45.480 32.300 ;
        RECT 43.980 30.850 44.630 31.500 ;
        RECT 44.830 30.850 45.480 31.500 ;
        RECT 43.980 28.500 44.630 29.150 ;
        RECT 44.830 28.500 45.480 29.150 ;
        RECT 43.980 27.700 44.630 28.350 ;
        RECT 44.830 27.700 45.480 28.350 ;
        RECT 43.980 26.900 44.630 27.550 ;
        RECT 44.830 26.900 45.480 27.550 ;
        RECT 63.980 32.450 64.630 33.100 ;
        RECT 64.830 32.450 65.480 33.100 ;
        RECT 63.980 31.650 64.630 32.300 ;
        RECT 64.830 31.650 65.480 32.300 ;
        RECT 63.980 30.850 64.630 31.500 ;
        RECT 64.830 30.850 65.480 31.500 ;
        RECT 63.980 28.500 64.630 29.150 ;
        RECT 64.830 28.500 65.480 29.150 ;
        RECT 63.980 27.700 64.630 28.350 ;
        RECT 64.830 27.700 65.480 28.350 ;
        RECT 63.980 26.900 64.630 27.550 ;
        RECT 64.830 26.900 65.480 27.550 ;
        RECT 83.980 32.450 84.630 33.100 ;
        RECT 84.830 32.450 85.480 33.100 ;
        RECT 83.980 31.650 84.630 32.300 ;
        RECT 84.830 31.650 85.480 32.300 ;
        RECT 83.980 30.850 84.630 31.500 ;
        RECT 84.830 30.850 85.480 31.500 ;
        RECT 83.980 28.500 84.630 29.150 ;
        RECT 84.830 28.500 85.480 29.150 ;
        RECT 83.980 27.700 84.630 28.350 ;
        RECT 84.830 27.700 85.480 28.350 ;
        RECT 83.980 26.900 84.630 27.550 ;
        RECT 84.830 26.900 85.480 27.550 ;
        RECT 103.980 32.450 104.630 33.100 ;
        RECT 103.980 31.650 104.630 32.300 ;
        RECT 103.980 30.850 104.630 31.500 ;
        RECT 103.980 28.500 104.630 29.150 ;
        RECT 103.980 27.700 104.630 28.350 ;
        RECT 103.980 26.900 104.630 27.550 ;
        RECT 11.630 20.100 12.280 20.750 ;
        RECT 12.430 20.100 13.080 20.750 ;
        RECT 13.230 20.100 13.880 20.750 ;
        RECT 15.580 20.100 16.230 20.750 ;
        RECT 16.380 20.100 17.030 20.750 ;
        RECT 17.180 20.100 17.830 20.750 ;
        RECT 11.630 19.250 12.280 19.900 ;
        RECT 12.430 19.250 13.080 19.900 ;
        RECT 13.230 19.250 13.880 19.900 ;
        RECT 15.580 19.250 16.230 19.900 ;
        RECT 16.380 19.250 17.030 19.900 ;
        RECT 17.180 19.250 17.830 19.900 ;
        RECT 31.630 20.100 32.280 20.750 ;
        RECT 32.430 20.100 33.080 20.750 ;
        RECT 33.230 20.100 33.880 20.750 ;
        RECT 35.580 20.100 36.230 20.750 ;
        RECT 36.380 20.100 37.030 20.750 ;
        RECT 37.180 20.100 37.830 20.750 ;
        RECT 31.630 19.250 32.280 19.900 ;
        RECT 32.430 19.250 33.080 19.900 ;
        RECT 33.230 19.250 33.880 19.900 ;
        RECT 35.580 19.250 36.230 19.900 ;
        RECT 36.380 19.250 37.030 19.900 ;
        RECT 37.180 19.250 37.830 19.900 ;
        RECT 51.630 20.100 52.280 20.750 ;
        RECT 52.430 20.100 53.080 20.750 ;
        RECT 53.230 20.100 53.880 20.750 ;
        RECT 55.580 20.100 56.230 20.750 ;
        RECT 56.380 20.100 57.030 20.750 ;
        RECT 57.180 20.100 57.830 20.750 ;
        RECT 51.630 19.250 52.280 19.900 ;
        RECT 52.430 19.250 53.080 19.900 ;
        RECT 53.230 19.250 53.880 19.900 ;
        RECT 55.580 19.250 56.230 19.900 ;
        RECT 56.380 19.250 57.030 19.900 ;
        RECT 57.180 19.250 57.830 19.900 ;
        RECT 71.630 20.100 72.280 20.750 ;
        RECT 72.430 20.100 73.080 20.750 ;
        RECT 73.230 20.100 73.880 20.750 ;
        RECT 75.580 20.100 76.230 20.750 ;
        RECT 76.380 20.100 77.030 20.750 ;
        RECT 77.180 20.100 77.830 20.750 ;
        RECT 71.630 19.250 72.280 19.900 ;
        RECT 72.430 19.250 73.080 19.900 ;
        RECT 73.230 19.250 73.880 19.900 ;
        RECT 75.580 19.250 76.230 19.900 ;
        RECT 76.380 19.250 77.030 19.900 ;
        RECT 77.180 19.250 77.830 19.900 ;
        RECT 91.630 20.100 92.280 20.750 ;
        RECT 92.430 20.100 93.080 20.750 ;
        RECT 93.230 20.100 93.880 20.750 ;
        RECT 95.580 20.100 96.230 20.750 ;
        RECT 96.380 20.100 97.030 20.750 ;
        RECT 97.180 20.100 97.830 20.750 ;
        RECT 91.630 19.250 92.280 19.900 ;
        RECT 92.430 19.250 93.080 19.900 ;
        RECT 93.230 19.250 93.880 19.900 ;
        RECT 95.580 19.250 96.230 19.900 ;
        RECT 96.380 19.250 97.030 19.900 ;
        RECT 97.180 19.250 97.830 19.900 ;
        RECT 4.830 12.450 5.480 13.100 ;
        RECT 4.830 11.650 5.480 12.300 ;
        RECT 4.830 10.850 5.480 11.500 ;
        RECT 4.830 8.500 5.480 9.150 ;
        RECT 4.830 7.700 5.480 8.350 ;
        RECT 4.830 6.900 5.480 7.550 ;
        RECT 23.980 12.450 24.630 13.100 ;
        RECT 24.830 12.450 25.480 13.100 ;
        RECT 23.980 11.650 24.630 12.300 ;
        RECT 24.830 11.650 25.480 12.300 ;
        RECT 23.980 10.850 24.630 11.500 ;
        RECT 24.830 10.850 25.480 11.500 ;
        RECT 23.980 8.500 24.630 9.150 ;
        RECT 24.830 8.500 25.480 9.150 ;
        RECT 23.980 7.700 24.630 8.350 ;
        RECT 24.830 7.700 25.480 8.350 ;
        RECT 23.980 6.900 24.630 7.550 ;
        RECT 24.830 6.900 25.480 7.550 ;
        RECT 43.980 12.450 44.630 13.100 ;
        RECT 44.830 12.450 45.480 13.100 ;
        RECT 43.980 11.650 44.630 12.300 ;
        RECT 44.830 11.650 45.480 12.300 ;
        RECT 43.980 10.850 44.630 11.500 ;
        RECT 44.830 10.850 45.480 11.500 ;
        RECT 43.980 8.500 44.630 9.150 ;
        RECT 44.830 8.500 45.480 9.150 ;
        RECT 43.980 7.700 44.630 8.350 ;
        RECT 44.830 7.700 45.480 8.350 ;
        RECT 43.980 6.900 44.630 7.550 ;
        RECT 44.830 6.900 45.480 7.550 ;
        RECT 63.980 12.450 64.630 13.100 ;
        RECT 64.830 12.450 65.480 13.100 ;
        RECT 63.980 11.650 64.630 12.300 ;
        RECT 64.830 11.650 65.480 12.300 ;
        RECT 63.980 10.850 64.630 11.500 ;
        RECT 64.830 10.850 65.480 11.500 ;
        RECT 63.980 8.500 64.630 9.150 ;
        RECT 64.830 8.500 65.480 9.150 ;
        RECT 63.980 7.700 64.630 8.350 ;
        RECT 64.830 7.700 65.480 8.350 ;
        RECT 63.980 6.900 64.630 7.550 ;
        RECT 64.830 6.900 65.480 7.550 ;
        RECT 83.980 12.450 84.630 13.100 ;
        RECT 84.830 12.450 85.480 13.100 ;
        RECT 83.980 11.650 84.630 12.300 ;
        RECT 84.830 11.650 85.480 12.300 ;
        RECT 83.980 10.850 84.630 11.500 ;
        RECT 84.830 10.850 85.480 11.500 ;
        RECT 83.980 8.500 84.630 9.150 ;
        RECT 84.830 8.500 85.480 9.150 ;
        RECT 83.980 7.700 84.630 8.350 ;
        RECT 84.830 7.700 85.480 8.350 ;
        RECT 83.980 6.900 84.630 7.550 ;
        RECT 84.830 6.900 85.480 7.550 ;
        RECT 103.980 12.450 104.630 13.100 ;
        RECT 103.980 11.650 104.630 12.300 ;
        RECT 103.980 10.850 104.630 11.500 ;
        RECT 103.980 8.500 104.630 9.150 ;
        RECT 103.980 7.700 104.630 8.350 ;
        RECT 103.980 6.900 104.630 7.550 ;
        RECT 11.630 0.100 12.280 0.750 ;
        RECT 12.430 0.100 13.080 0.750 ;
        RECT 13.230 0.100 13.880 0.750 ;
        RECT 15.580 0.100 16.230 0.750 ;
        RECT 16.380 0.100 17.030 0.750 ;
        RECT 17.180 0.100 17.830 0.750 ;
        RECT 31.630 0.100 32.280 0.750 ;
        RECT 32.430 0.100 33.080 0.750 ;
        RECT 33.230 0.100 33.880 0.750 ;
        RECT 35.580 0.100 36.230 0.750 ;
        RECT 36.380 0.100 37.030 0.750 ;
        RECT 37.180 0.100 37.830 0.750 ;
        RECT 51.630 0.100 52.280 0.750 ;
        RECT 52.430 0.100 53.080 0.750 ;
        RECT 53.230 0.100 53.880 0.750 ;
        RECT 55.580 0.100 56.230 0.750 ;
        RECT 56.380 0.100 57.030 0.750 ;
        RECT 57.180 0.100 57.830 0.750 ;
        RECT 71.630 0.100 72.280 0.750 ;
        RECT 72.430 0.100 73.080 0.750 ;
        RECT 73.230 0.100 73.880 0.750 ;
        RECT 75.580 0.100 76.230 0.750 ;
        RECT 76.380 0.100 77.030 0.750 ;
        RECT 77.180 0.100 77.830 0.750 ;
        RECT 91.630 0.100 92.280 0.750 ;
        RECT 92.430 0.100 93.080 0.750 ;
        RECT 93.230 0.100 93.880 0.750 ;
        RECT 95.580 0.100 96.230 0.750 ;
        RECT 96.380 0.100 97.030 0.750 ;
        RECT 97.180 0.100 97.830 0.750 ;
      LAYER met4 ;
        RECT 4.730 378.950 9.130 380.000 ;
        RECT 4.730 375.600 5.780 378.950 ;
        RECT 11.530 378.550 17.930 380.000 ;
        RECT 20.330 378.950 29.130 380.000 ;
        RECT 6.180 373.200 23.280 378.550 ;
        RECT 23.680 375.600 25.780 378.950 ;
        RECT 31.530 378.550 37.930 380.000 ;
        RECT 40.330 378.950 49.130 380.000 ;
        RECT 26.180 373.200 43.280 378.550 ;
        RECT 43.680 375.600 45.780 378.950 ;
        RECT 51.530 378.550 57.930 380.000 ;
        RECT 60.330 378.950 69.130 380.000 ;
        RECT 46.180 373.200 63.280 378.550 ;
        RECT 63.680 375.600 65.780 378.950 ;
        RECT 71.530 378.550 77.930 380.000 ;
        RECT 80.330 378.950 89.130 380.000 ;
        RECT 66.180 373.200 83.280 378.550 ;
        RECT 83.680 375.600 85.780 378.950 ;
        RECT 91.530 378.550 97.930 380.000 ;
        RECT 100.330 378.950 104.730 380.000 ;
        RECT 86.180 373.200 103.280 378.550 ;
        RECT 103.680 375.600 104.730 378.950 ;
        RECT 4.730 366.800 104.730 373.200 ;
        RECT 4.730 361.050 5.780 364.400 ;
        RECT 6.180 361.450 23.280 366.800 ;
        RECT 4.730 358.950 9.130 361.050 ;
        RECT 4.730 355.600 5.780 358.950 ;
        RECT 11.530 358.550 17.930 361.450 ;
        RECT 23.680 361.050 25.780 364.400 ;
        RECT 26.180 361.450 43.280 366.800 ;
        RECT 20.330 358.950 29.130 361.050 ;
        RECT 6.180 353.200 23.280 358.550 ;
        RECT 23.680 355.600 25.780 358.950 ;
        RECT 31.530 358.550 37.930 361.450 ;
        RECT 43.680 361.050 45.780 364.400 ;
        RECT 46.180 361.450 63.280 366.800 ;
        RECT 40.330 358.950 49.130 361.050 ;
        RECT 26.180 353.200 43.280 358.550 ;
        RECT 43.680 355.600 45.780 358.950 ;
        RECT 51.530 358.550 57.930 361.450 ;
        RECT 63.680 361.050 65.780 364.400 ;
        RECT 66.180 361.450 83.280 366.800 ;
        RECT 60.330 358.950 69.130 361.050 ;
        RECT 46.180 353.200 63.280 358.550 ;
        RECT 63.680 355.600 65.780 358.950 ;
        RECT 71.530 358.550 77.930 361.450 ;
        RECT 83.680 361.050 85.780 364.400 ;
        RECT 86.180 361.450 103.280 366.800 ;
        RECT 80.330 358.950 89.130 361.050 ;
        RECT 66.180 353.200 83.280 358.550 ;
        RECT 83.680 355.600 85.780 358.950 ;
        RECT 91.530 358.550 97.930 361.450 ;
        RECT 103.680 361.050 104.730 364.400 ;
        RECT 100.330 358.950 104.730 361.050 ;
        RECT 86.180 353.200 103.280 358.550 ;
        RECT 103.680 355.600 104.730 358.950 ;
        RECT 4.730 346.800 104.730 353.200 ;
        RECT 4.730 341.050 5.780 344.400 ;
        RECT 6.180 341.450 23.280 346.800 ;
        RECT 4.730 338.950 9.130 341.050 ;
        RECT 4.730 335.600 5.780 338.950 ;
        RECT 11.530 338.550 17.930 341.450 ;
        RECT 23.680 341.050 25.780 344.400 ;
        RECT 26.180 341.450 43.280 346.800 ;
        RECT 20.330 338.950 29.130 341.050 ;
        RECT 6.180 333.200 23.280 338.550 ;
        RECT 23.680 335.600 25.780 338.950 ;
        RECT 31.530 338.550 37.930 341.450 ;
        RECT 43.680 341.050 45.780 344.400 ;
        RECT 46.180 341.450 63.280 346.800 ;
        RECT 40.330 338.950 49.130 341.050 ;
        RECT 26.180 333.200 43.280 338.550 ;
        RECT 43.680 335.600 45.780 338.950 ;
        RECT 51.530 338.550 57.930 341.450 ;
        RECT 63.680 341.050 65.780 344.400 ;
        RECT 66.180 341.450 83.280 346.800 ;
        RECT 60.330 338.950 69.130 341.050 ;
        RECT 46.180 333.200 63.280 338.550 ;
        RECT 63.680 335.600 65.780 338.950 ;
        RECT 71.530 338.550 77.930 341.450 ;
        RECT 83.680 341.050 85.780 344.400 ;
        RECT 86.180 341.450 103.280 346.800 ;
        RECT 80.330 338.950 89.130 341.050 ;
        RECT 66.180 333.200 83.280 338.550 ;
        RECT 83.680 335.600 85.780 338.950 ;
        RECT 91.530 338.550 97.930 341.450 ;
        RECT 103.680 341.050 104.730 344.400 ;
        RECT 100.330 338.950 104.730 341.050 ;
        RECT 86.180 333.200 103.280 338.550 ;
        RECT 103.680 335.600 104.730 338.950 ;
        RECT 4.730 326.800 104.730 333.200 ;
        RECT 4.730 321.050 5.780 324.400 ;
        RECT 6.180 321.450 23.280 326.800 ;
        RECT 4.730 318.950 9.130 321.050 ;
        RECT 4.730 315.600 5.780 318.950 ;
        RECT 11.530 318.550 17.930 321.450 ;
        RECT 23.680 321.050 25.780 324.400 ;
        RECT 26.180 321.450 43.280 326.800 ;
        RECT 20.330 318.950 29.130 321.050 ;
        RECT 6.180 313.200 23.280 318.550 ;
        RECT 23.680 315.600 25.780 318.950 ;
        RECT 31.530 318.550 37.930 321.450 ;
        RECT 43.680 321.050 45.780 324.400 ;
        RECT 46.180 321.450 63.280 326.800 ;
        RECT 40.330 318.950 49.130 321.050 ;
        RECT 26.180 313.200 43.280 318.550 ;
        RECT 43.680 315.600 45.780 318.950 ;
        RECT 51.530 318.550 57.930 321.450 ;
        RECT 63.680 321.050 65.780 324.400 ;
        RECT 66.180 321.450 83.280 326.800 ;
        RECT 60.330 318.950 69.130 321.050 ;
        RECT 46.180 313.200 63.280 318.550 ;
        RECT 63.680 315.600 65.780 318.950 ;
        RECT 71.530 318.550 77.930 321.450 ;
        RECT 83.680 321.050 85.780 324.400 ;
        RECT 86.180 321.450 103.280 326.800 ;
        RECT 80.330 318.950 89.130 321.050 ;
        RECT 66.180 313.200 83.280 318.550 ;
        RECT 83.680 315.600 85.780 318.950 ;
        RECT 91.530 318.550 97.930 321.450 ;
        RECT 103.680 321.050 104.730 324.400 ;
        RECT 100.330 318.950 104.730 321.050 ;
        RECT 86.180 313.200 103.280 318.550 ;
        RECT 103.680 315.600 104.730 318.950 ;
        RECT 4.730 306.800 104.730 313.200 ;
        RECT 4.730 301.050 5.780 304.400 ;
        RECT 6.180 301.450 23.280 306.800 ;
        RECT 4.730 298.950 9.130 301.050 ;
        RECT 4.730 295.600 5.780 298.950 ;
        RECT 11.530 298.550 17.930 301.450 ;
        RECT 23.680 301.050 25.780 304.400 ;
        RECT 26.180 301.450 43.280 306.800 ;
        RECT 20.330 298.950 29.130 301.050 ;
        RECT 6.180 293.200 23.280 298.550 ;
        RECT 23.680 295.600 25.780 298.950 ;
        RECT 31.530 298.550 37.930 301.450 ;
        RECT 43.680 301.050 45.780 304.400 ;
        RECT 46.180 301.450 63.280 306.800 ;
        RECT 40.330 298.950 49.130 301.050 ;
        RECT 26.180 293.200 43.280 298.550 ;
        RECT 43.680 295.600 45.780 298.950 ;
        RECT 51.530 298.550 57.930 301.450 ;
        RECT 63.680 301.050 65.780 304.400 ;
        RECT 66.180 301.450 83.280 306.800 ;
        RECT 60.330 298.950 69.130 301.050 ;
        RECT 46.180 293.200 63.280 298.550 ;
        RECT 63.680 295.600 65.780 298.950 ;
        RECT 71.530 298.550 77.930 301.450 ;
        RECT 83.680 301.050 85.780 304.400 ;
        RECT 86.180 301.450 103.280 306.800 ;
        RECT 80.330 298.950 89.130 301.050 ;
        RECT 66.180 293.200 83.280 298.550 ;
        RECT 83.680 295.600 85.780 298.950 ;
        RECT 91.530 298.550 97.930 301.450 ;
        RECT 103.680 301.050 104.730 304.400 ;
        RECT 100.330 298.950 104.730 301.050 ;
        RECT 86.180 293.200 103.280 298.550 ;
        RECT 103.680 295.600 104.730 298.950 ;
        RECT 4.730 286.800 104.730 293.200 ;
        RECT 4.730 281.050 5.780 284.400 ;
        RECT 6.180 281.450 23.280 286.800 ;
        RECT 4.730 278.950 9.130 281.050 ;
        RECT 4.730 275.600 5.780 278.950 ;
        RECT 11.530 278.550 17.930 281.450 ;
        RECT 23.680 281.050 25.780 284.400 ;
        RECT 26.180 281.450 43.280 286.800 ;
        RECT 20.330 278.950 29.130 281.050 ;
        RECT 6.180 273.200 23.280 278.550 ;
        RECT 23.680 275.600 25.780 278.950 ;
        RECT 31.530 278.550 37.930 281.450 ;
        RECT 43.680 281.050 45.780 284.400 ;
        RECT 46.180 281.450 63.280 286.800 ;
        RECT 40.330 278.950 49.130 281.050 ;
        RECT 26.180 273.200 43.280 278.550 ;
        RECT 43.680 275.600 45.780 278.950 ;
        RECT 51.530 278.550 57.930 281.450 ;
        RECT 63.680 281.050 65.780 284.400 ;
        RECT 66.180 281.450 83.280 286.800 ;
        RECT 60.330 278.950 69.130 281.050 ;
        RECT 46.180 273.200 63.280 278.550 ;
        RECT 63.680 275.600 65.780 278.950 ;
        RECT 71.530 278.550 77.930 281.450 ;
        RECT 83.680 281.050 85.780 284.400 ;
        RECT 86.180 281.450 103.280 286.800 ;
        RECT 80.330 278.950 89.130 281.050 ;
        RECT 66.180 273.200 83.280 278.550 ;
        RECT 83.680 275.600 85.780 278.950 ;
        RECT 91.530 278.550 97.930 281.450 ;
        RECT 103.680 281.050 104.730 284.400 ;
        RECT 100.330 278.950 104.730 281.050 ;
        RECT 86.180 273.200 103.280 278.550 ;
        RECT 103.680 275.600 104.730 278.950 ;
        RECT 4.730 266.800 104.730 273.200 ;
        RECT 4.730 261.050 5.780 264.400 ;
        RECT 6.180 261.450 23.280 266.800 ;
        RECT 4.730 258.950 9.130 261.050 ;
        RECT 4.730 255.600 5.780 258.950 ;
        RECT 11.530 258.550 17.930 261.450 ;
        RECT 23.680 261.050 25.780 264.400 ;
        RECT 26.180 261.450 43.280 266.800 ;
        RECT 20.330 258.950 29.130 261.050 ;
        RECT 6.180 253.200 23.280 258.550 ;
        RECT 23.680 255.600 25.780 258.950 ;
        RECT 31.530 258.550 37.930 261.450 ;
        RECT 43.680 261.050 45.780 264.400 ;
        RECT 46.180 261.450 63.280 266.800 ;
        RECT 40.330 258.950 49.130 261.050 ;
        RECT 26.180 253.200 43.280 258.550 ;
        RECT 43.680 255.600 45.780 258.950 ;
        RECT 51.530 258.550 57.930 261.450 ;
        RECT 63.680 261.050 65.780 264.400 ;
        RECT 66.180 261.450 83.280 266.800 ;
        RECT 60.330 258.950 69.130 261.050 ;
        RECT 46.180 253.200 63.280 258.550 ;
        RECT 63.680 255.600 65.780 258.950 ;
        RECT 71.530 258.550 77.930 261.450 ;
        RECT 83.680 261.050 85.780 264.400 ;
        RECT 86.180 261.450 103.280 266.800 ;
        RECT 80.330 258.950 89.130 261.050 ;
        RECT 66.180 253.200 83.280 258.550 ;
        RECT 83.680 255.600 85.780 258.950 ;
        RECT 91.530 258.550 97.930 261.450 ;
        RECT 103.680 261.050 104.730 264.400 ;
        RECT 100.330 258.950 104.730 261.050 ;
        RECT 86.180 253.200 103.280 258.550 ;
        RECT 103.680 255.600 104.730 258.950 ;
        RECT 4.730 246.800 104.730 253.200 ;
        RECT 4.730 241.050 5.780 244.400 ;
        RECT 6.180 241.450 23.280 246.800 ;
        RECT 4.730 238.950 9.130 241.050 ;
        RECT 4.730 235.600 5.780 238.950 ;
        RECT 11.530 238.550 17.930 241.450 ;
        RECT 23.680 241.050 25.780 244.400 ;
        RECT 26.180 241.450 43.280 246.800 ;
        RECT 20.330 238.950 29.130 241.050 ;
        RECT 6.180 233.200 23.280 238.550 ;
        RECT 23.680 235.600 25.780 238.950 ;
        RECT 31.530 238.550 37.930 241.450 ;
        RECT 43.680 241.050 45.780 244.400 ;
        RECT 46.180 241.450 63.280 246.800 ;
        RECT 40.330 238.950 49.130 241.050 ;
        RECT 26.180 233.200 43.280 238.550 ;
        RECT 43.680 235.600 45.780 238.950 ;
        RECT 51.530 238.550 57.930 241.450 ;
        RECT 63.680 241.050 65.780 244.400 ;
        RECT 66.180 241.450 83.280 246.800 ;
        RECT 60.330 238.950 69.130 241.050 ;
        RECT 46.180 233.200 63.280 238.550 ;
        RECT 63.680 235.600 65.780 238.950 ;
        RECT 71.530 238.550 77.930 241.450 ;
        RECT 83.680 241.050 85.780 244.400 ;
        RECT 86.180 241.450 103.280 246.800 ;
        RECT 80.330 238.950 89.130 241.050 ;
        RECT 66.180 233.200 83.280 238.550 ;
        RECT 83.680 235.600 85.780 238.950 ;
        RECT 91.530 238.550 97.930 241.450 ;
        RECT 103.680 241.050 104.730 244.400 ;
        RECT 100.330 238.950 104.730 241.050 ;
        RECT 86.180 233.200 103.280 238.550 ;
        RECT 103.680 235.600 104.730 238.950 ;
        RECT 4.730 226.800 104.730 233.200 ;
        RECT 4.730 221.050 5.780 224.400 ;
        RECT 6.180 221.450 23.280 226.800 ;
        RECT 4.730 220.000 9.130 221.050 ;
        RECT 11.530 220.000 17.930 221.450 ;
        RECT 23.680 221.050 25.780 224.400 ;
        RECT 26.180 221.450 43.280 226.800 ;
        RECT 20.330 220.000 29.130 221.050 ;
        RECT 31.530 220.000 37.930 221.450 ;
        RECT 43.680 221.050 45.780 224.400 ;
        RECT 46.180 221.450 63.280 226.800 ;
        RECT 40.330 220.000 49.130 221.050 ;
        RECT 51.530 220.000 57.930 221.450 ;
        RECT 63.680 221.050 65.780 224.400 ;
        RECT 66.180 221.450 83.280 226.800 ;
        RECT 60.330 220.000 69.130 221.050 ;
        RECT 71.530 220.000 77.930 221.450 ;
        RECT 83.680 221.050 85.780 224.400 ;
        RECT 86.180 221.450 103.280 226.800 ;
        RECT 80.330 220.000 89.130 221.050 ;
        RECT 91.530 220.000 97.930 221.450 ;
        RECT 103.680 221.050 104.730 224.400 ;
        RECT 100.330 220.000 104.730 221.050 ;
        RECT 11.530 199.710 14.340 220.000 ;
        RECT 11.230 198.875 14.340 199.710 ;
        RECT 11.530 198.870 14.340 198.875 ;
        RECT 20.595 198.770 22.450 220.000 ;
        RECT 11.530 160.000 13.690 182.380 ;
        RECT 11.530 158.550 17.930 160.000 ;
        RECT 31.530 158.550 37.930 160.000 ;
        RECT 51.530 158.550 57.930 160.000 ;
        RECT 71.530 158.550 77.930 160.000 ;
        RECT 91.530 158.550 97.930 160.000 ;
        RECT 6.180 153.200 23.280 158.550 ;
        RECT 26.180 153.200 43.280 158.550 ;
        RECT 46.180 153.200 63.280 158.550 ;
        RECT 66.180 153.200 83.280 158.550 ;
        RECT 86.180 153.200 103.280 158.550 ;
        RECT 4.730 146.800 104.730 153.200 ;
        RECT 6.180 141.450 23.280 146.800 ;
        RECT 26.180 141.450 43.280 146.800 ;
        RECT 46.180 141.450 63.280 146.800 ;
        RECT 66.180 141.450 83.280 146.800 ;
        RECT 86.180 141.450 103.280 146.800 ;
        RECT 11.530 138.550 17.930 141.450 ;
        RECT 31.530 138.550 37.930 141.450 ;
        RECT 51.530 138.550 57.930 141.450 ;
        RECT 71.530 138.550 77.930 141.450 ;
        RECT 91.530 138.550 97.930 141.450 ;
        RECT 6.180 133.200 23.280 138.550 ;
        RECT 26.180 133.200 43.280 138.550 ;
        RECT 46.180 133.200 63.280 138.550 ;
        RECT 66.180 133.200 83.280 138.550 ;
        RECT 86.180 133.200 103.280 138.550 ;
        RECT 4.730 126.800 104.730 133.200 ;
        RECT 6.180 121.450 23.280 126.800 ;
        RECT 26.180 121.450 43.280 126.800 ;
        RECT 46.180 121.450 63.280 126.800 ;
        RECT 66.180 121.450 83.280 126.800 ;
        RECT 86.180 121.450 103.280 126.800 ;
        RECT 11.530 118.550 17.930 121.450 ;
        RECT 31.530 118.550 37.930 121.450 ;
        RECT 51.530 118.550 57.930 121.450 ;
        RECT 71.530 118.550 77.930 121.450 ;
        RECT 91.530 118.550 97.930 121.450 ;
        RECT 6.180 113.200 23.280 118.550 ;
        RECT 26.180 113.200 43.280 118.550 ;
        RECT 46.180 113.200 63.280 118.550 ;
        RECT 66.180 113.200 83.280 118.550 ;
        RECT 86.180 113.200 103.280 118.550 ;
        RECT 4.730 106.800 104.730 113.200 ;
        RECT 6.180 101.450 23.280 106.800 ;
        RECT 26.180 101.450 43.280 106.800 ;
        RECT 46.180 101.450 63.280 106.800 ;
        RECT 66.180 101.450 83.280 106.800 ;
        RECT 86.180 101.450 103.280 106.800 ;
        RECT 11.530 98.550 17.930 101.450 ;
        RECT 31.530 98.550 37.930 101.450 ;
        RECT 51.530 98.550 57.930 101.450 ;
        RECT 71.530 98.550 77.930 101.450 ;
        RECT 91.530 98.550 97.930 101.450 ;
        RECT 6.180 93.200 23.280 98.550 ;
        RECT 26.180 93.200 43.280 98.550 ;
        RECT 46.180 93.200 63.280 98.550 ;
        RECT 66.180 93.200 83.280 98.550 ;
        RECT 86.180 93.200 103.280 98.550 ;
        RECT 4.730 86.800 104.730 93.200 ;
        RECT 6.180 81.450 23.280 86.800 ;
        RECT 26.180 81.450 43.280 86.800 ;
        RECT 46.180 81.450 63.280 86.800 ;
        RECT 66.180 81.450 83.280 86.800 ;
        RECT 86.180 81.450 103.280 86.800 ;
        RECT 11.530 78.550 17.930 81.450 ;
        RECT 31.530 78.550 37.930 81.450 ;
        RECT 51.530 78.550 57.930 81.450 ;
        RECT 71.530 78.550 77.930 81.450 ;
        RECT 91.530 78.550 97.930 81.450 ;
        RECT 6.180 73.200 23.280 78.550 ;
        RECT 26.180 73.200 43.280 78.550 ;
        RECT 46.180 73.200 63.280 78.550 ;
        RECT 66.180 73.200 83.280 78.550 ;
        RECT 86.180 73.200 103.280 78.550 ;
        RECT 4.730 66.800 104.730 73.200 ;
        RECT 6.180 61.450 23.280 66.800 ;
        RECT 26.180 61.450 43.280 66.800 ;
        RECT 46.180 61.450 63.280 66.800 ;
        RECT 66.180 61.450 83.280 66.800 ;
        RECT 86.180 61.450 103.280 66.800 ;
        RECT 11.530 58.550 17.930 61.450 ;
        RECT 31.530 58.550 37.930 61.450 ;
        RECT 51.530 58.550 57.930 61.450 ;
        RECT 71.530 58.550 77.930 61.450 ;
        RECT 91.530 58.550 97.930 61.450 ;
        RECT 6.180 53.200 23.280 58.550 ;
        RECT 26.180 53.200 43.280 58.550 ;
        RECT 46.180 53.200 63.280 58.550 ;
        RECT 66.180 53.200 83.280 58.550 ;
        RECT 86.180 53.200 103.280 58.550 ;
        RECT 4.730 46.800 104.730 53.200 ;
        RECT 6.180 41.450 23.280 46.800 ;
        RECT 26.180 41.450 43.280 46.800 ;
        RECT 46.180 41.450 63.280 46.800 ;
        RECT 66.180 41.450 83.280 46.800 ;
        RECT 86.180 41.450 103.280 46.800 ;
        RECT 11.530 38.550 17.930 41.450 ;
        RECT 31.530 38.550 37.930 41.450 ;
        RECT 51.530 38.550 57.930 41.450 ;
        RECT 71.530 38.550 77.930 41.450 ;
        RECT 91.530 38.550 97.930 41.450 ;
        RECT 6.180 33.200 23.280 38.550 ;
        RECT 26.180 33.200 43.280 38.550 ;
        RECT 46.180 33.200 63.280 38.550 ;
        RECT 66.180 33.200 83.280 38.550 ;
        RECT 86.180 33.200 103.280 38.550 ;
        RECT 4.730 26.800 104.730 33.200 ;
        RECT 6.180 21.450 23.280 26.800 ;
        RECT 26.180 21.450 43.280 26.800 ;
        RECT 46.180 21.450 63.280 26.800 ;
        RECT 66.180 21.450 83.280 26.800 ;
        RECT 86.180 21.450 103.280 26.800 ;
        RECT 11.530 18.550 17.930 21.450 ;
        RECT 31.530 18.550 37.930 21.450 ;
        RECT 51.530 18.550 57.930 21.450 ;
        RECT 71.530 18.550 77.930 21.450 ;
        RECT 91.530 18.550 97.930 21.450 ;
        RECT 6.180 13.200 23.280 18.550 ;
        RECT 26.180 13.200 43.280 18.550 ;
        RECT 46.180 13.200 63.280 18.550 ;
        RECT 66.180 13.200 83.280 18.550 ;
        RECT 86.180 13.200 103.280 18.550 ;
        RECT 4.730 6.800 104.730 13.200 ;
        RECT 6.180 1.450 23.280 6.800 ;
        RECT 26.180 1.450 43.280 6.800 ;
        RECT 46.180 1.450 63.280 6.800 ;
        RECT 66.180 1.450 83.280 6.800 ;
        RECT 86.180 1.450 103.280 6.800 ;
        RECT 11.530 0.000 17.930 1.450 ;
        RECT 31.530 0.000 37.930 1.450 ;
        RECT 51.530 0.000 57.930 1.450 ;
        RECT 71.530 0.000 77.930 1.450 ;
        RECT 91.530 0.000 97.930 1.450 ;
  END
END adc_vcm_generator
END LIBRARY

